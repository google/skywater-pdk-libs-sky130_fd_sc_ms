* File: sky130_fd_sc_ms__sdfsbp_2.pxi.spice
* Created: Wed Sep  2 12:31:01 2020
* 
x_PM_SKY130_FD_SC_MS__SDFSBP_2%A_27_74# N_A_27_74#_M1044_s N_A_27_74#_M1009_s
+ N_A_27_74#_M1037_g N_A_27_74#_M1027_g N_A_27_74#_c_357_n N_A_27_74#_c_358_n
+ N_A_27_74#_c_365_n N_A_27_74#_c_359_n N_A_27_74#_c_360_n N_A_27_74#_c_366_n
+ N_A_27_74#_c_361_n N_A_27_74#_c_367_n N_A_27_74#_c_368_n N_A_27_74#_c_369_n
+ N_A_27_74#_c_362_n PM_SKY130_FD_SC_MS__SDFSBP_2%A_27_74#
x_PM_SKY130_FD_SC_MS__SDFSBP_2%SCE N_SCE_M1044_g N_SCE_M1009_g N_SCE_M1007_g
+ N_SCE_M1017_g N_SCE_c_435_n N_SCE_c_436_n N_SCE_c_437_n N_SCE_c_438_n SCE
+ N_SCE_c_439_n N_SCE_c_440_n N_SCE_c_441_n PM_SKY130_FD_SC_MS__SDFSBP_2%SCE
x_PM_SKY130_FD_SC_MS__SDFSBP_2%D N_D_c_512_n N_D_M1033_g N_D_M1038_g N_D_c_514_n
+ D D N_D_c_516_n N_D_c_517_n PM_SKY130_FD_SC_MS__SDFSBP_2%D
x_PM_SKY130_FD_SC_MS__SDFSBP_2%SCD N_SCD_M1041_g N_SCD_c_565_n N_SCD_c_566_n
+ N_SCD_M1015_g N_SCD_c_559_n N_SCD_c_560_n N_SCD_c_561_n SCD N_SCD_c_563_n
+ PM_SKY130_FD_SC_MS__SDFSBP_2%SCD
x_PM_SKY130_FD_SC_MS__SDFSBP_2%CLK N_CLK_M1036_g N_CLK_c_610_n N_CLK_M1043_g CLK
+ N_CLK_c_612_n PM_SKY130_FD_SC_MS__SDFSBP_2%CLK
x_PM_SKY130_FD_SC_MS__SDFSBP_2%A_871_74# N_A_871_74#_M1035_d N_A_871_74#_M1046_d
+ N_A_871_74#_M1006_g N_A_871_74#_c_646_n N_A_871_74#_c_647_n
+ N_A_871_74#_M1026_g N_A_871_74#_M1032_g N_A_871_74#_M1039_g
+ N_A_871_74#_c_651_n N_A_871_74#_c_652_n N_A_871_74#_c_653_n
+ N_A_871_74#_M1010_g N_A_871_74#_c_671_n N_A_871_74#_c_655_n
+ N_A_871_74#_c_672_n N_A_871_74#_c_656_n N_A_871_74#_c_657_n
+ N_A_871_74#_c_673_n N_A_871_74#_c_674_n N_A_871_74#_c_658_n
+ N_A_871_74#_c_659_n N_A_871_74#_c_660_n N_A_871_74#_c_661_n
+ N_A_871_74#_c_678_n N_A_871_74#_c_679_n N_A_871_74#_c_680_n
+ N_A_871_74#_c_681_n N_A_871_74#_c_682_n N_A_871_74#_c_683_n
+ N_A_871_74#_c_684_n N_A_871_74#_c_685_n N_A_871_74#_c_662_n
+ N_A_871_74#_c_663_n N_A_871_74#_c_664_n N_A_871_74#_c_665_n
+ N_A_871_74#_c_666_n N_A_871_74#_c_687_n N_A_871_74#_c_667_n
+ N_A_871_74#_c_668_n PM_SKY130_FD_SC_MS__SDFSBP_2%A_871_74#
x_PM_SKY130_FD_SC_MS__SDFSBP_2%A_1252_376# N_A_1252_376#_M1013_s
+ N_A_1252_376#_M1042_d N_A_1252_376#_M1030_g N_A_1252_376#_c_911_n
+ N_A_1252_376#_c_912_n N_A_1252_376#_c_904_n N_A_1252_376#_M1024_g
+ N_A_1252_376#_c_913_n N_A_1252_376#_c_914_n N_A_1252_376#_c_905_n
+ N_A_1252_376#_c_906_n N_A_1252_376#_c_907_n N_A_1252_376#_c_915_n
+ N_A_1252_376#_c_916_n N_A_1252_376#_c_908_n N_A_1252_376#_c_909_n
+ PM_SKY130_FD_SC_MS__SDFSBP_2%A_1252_376#
x_PM_SKY130_FD_SC_MS__SDFSBP_2%A_1069_81# N_A_1069_81#_M1019_d
+ N_A_1069_81#_M1006_d N_A_1069_81#_M1042_g N_A_1069_81#_M1013_g
+ N_A_1069_81#_c_992_n N_A_1069_81#_M1003_g N_A_1069_81#_M1005_g
+ N_A_1069_81#_c_994_n N_A_1069_81#_M1048_g N_A_1069_81#_M1011_g
+ N_A_1069_81#_c_997_n N_A_1069_81#_c_998_n N_A_1069_81#_c_999_n
+ N_A_1069_81#_c_1029_n N_A_1069_81#_c_1033_n N_A_1069_81#_c_1000_n
+ N_A_1069_81#_c_1001_n N_A_1069_81#_c_1002_n N_A_1069_81#_c_1003_n
+ N_A_1069_81#_c_1004_n N_A_1069_81#_c_1005_n N_A_1069_81#_c_1006_n
+ N_A_1069_81#_c_1013_n N_A_1069_81#_c_1007_n N_A_1069_81#_c_1008_n
+ N_A_1069_81#_c_1009_n PM_SKY130_FD_SC_MS__SDFSBP_2%A_1069_81#
x_PM_SKY130_FD_SC_MS__SDFSBP_2%SET_B N_SET_B_M1034_g N_SET_B_M1014_g
+ N_SET_B_M1021_g N_SET_B_M1018_g N_SET_B_c_1171_n N_SET_B_c_1182_n
+ N_SET_B_c_1172_n N_SET_B_c_1173_n N_SET_B_c_1174_n SET_B N_SET_B_c_1176_n
+ N_SET_B_c_1177_n N_SET_B_c_1178_n PM_SKY130_FD_SC_MS__SDFSBP_2%SET_B
x_PM_SKY130_FD_SC_MS__SDFSBP_2%A_619_368# N_A_619_368#_M1043_s
+ N_A_619_368#_M1036_s N_A_619_368#_M1035_g N_A_619_368#_M1046_g
+ N_A_619_368#_c_1312_n N_A_619_368#_c_1330_n N_A_619_368#_c_1313_n
+ N_A_619_368#_c_1314_n N_A_619_368#_c_1331_n N_A_619_368#_c_1332_n
+ N_A_619_368#_c_1315_n N_A_619_368#_M1019_g N_A_619_368#_M1002_g
+ N_A_619_368#_c_1334_n N_A_619_368#_c_1335_n N_A_619_368#_c_1336_n
+ N_A_619_368#_M1028_g N_A_619_368#_c_1337_n N_A_619_368#_c_1338_n
+ N_A_619_368#_c_1339_n N_A_619_368#_M1031_g N_A_619_368#_c_1340_n
+ N_A_619_368#_c_1341_n N_A_619_368#_c_1342_n N_A_619_368#_c_1343_n
+ N_A_619_368#_c_1316_n N_A_619_368#_c_1317_n N_A_619_368#_c_1318_n
+ N_A_619_368#_M1008_g N_A_619_368#_c_1319_n N_A_619_368#_c_1320_n
+ N_A_619_368#_c_1321_n N_A_619_368#_c_1348_n N_A_619_368#_c_1349_n
+ N_A_619_368#_c_1322_n N_A_619_368#_c_1323_n N_A_619_368#_c_1324_n
+ N_A_619_368#_c_1350_n N_A_619_368#_c_1325_n N_A_619_368#_c_1352_n
+ N_A_619_368#_c_1326_n N_A_619_368#_c_1353_n N_A_619_368#_c_1327_n
+ N_A_619_368#_c_1328_n N_A_619_368#_c_1355_n
+ PM_SKY130_FD_SC_MS__SDFSBP_2%A_619_368#
x_PM_SKY130_FD_SC_MS__SDFSBP_2%A_2513_258# N_A_2513_258#_M1040_d
+ N_A_2513_258#_M1045_s N_A_2513_258#_M1016_g N_A_2513_258#_M1020_g
+ N_A_2513_258#_c_1574_n N_A_2513_258#_c_1584_n N_A_2513_258#_c_1575_n
+ N_A_2513_258#_c_1576_n N_A_2513_258#_c_1577_n N_A_2513_258#_c_1578_n
+ N_A_2513_258#_c_1579_n N_A_2513_258#_c_1580_n N_A_2513_258#_c_1581_n
+ N_A_2513_258#_c_1587_n PM_SKY130_FD_SC_MS__SDFSBP_2%A_2513_258#
x_PM_SKY130_FD_SC_MS__SDFSBP_2%A_2067_74# N_A_2067_74#_M1032_s
+ N_A_2067_74#_M1008_s N_A_2067_74#_M1028_d N_A_2067_74#_M1010_d
+ N_A_2067_74#_M1018_d N_A_2067_74#_M1040_g N_A_2067_74#_c_1670_n
+ N_A_2067_74#_c_1689_n N_A_2067_74#_c_1690_n N_A_2067_74#_M1045_g
+ N_A_2067_74#_M1023_g N_A_2067_74#_M1004_g N_A_2067_74#_c_1673_n
+ N_A_2067_74#_M1025_g N_A_2067_74#_M1029_g N_A_2067_74#_c_1676_n
+ N_A_2067_74#_M1000_g N_A_2067_74#_M1012_g N_A_2067_74#_c_1679_n
+ N_A_2067_74#_c_1680_n N_A_2067_74#_c_1681_n N_A_2067_74#_c_1682_n
+ N_A_2067_74#_c_1719_n N_A_2067_74#_c_1695_n N_A_2067_74#_c_1720_n
+ N_A_2067_74#_c_1683_n N_A_2067_74#_c_1754_n N_A_2067_74#_c_1684_n
+ N_A_2067_74#_c_1696_n N_A_2067_74#_c_1697_n N_A_2067_74#_c_1698_n
+ N_A_2067_74#_c_1699_n N_A_2067_74#_c_1685_n N_A_2067_74#_c_1686_n
+ N_A_2067_74#_c_1687_n N_A_2067_74#_c_1701_n N_A_2067_74#_c_1688_n
+ PM_SKY130_FD_SC_MS__SDFSBP_2%A_2067_74#
x_PM_SKY130_FD_SC_MS__SDFSBP_2%A_3177_368# N_A_3177_368#_M1012_s
+ N_A_3177_368#_M1000_s N_A_3177_368#_M1047_g N_A_3177_368#_M1001_g
+ N_A_3177_368#_M1049_g N_A_3177_368#_M1022_g N_A_3177_368#_c_1892_n
+ N_A_3177_368#_c_1893_n N_A_3177_368#_c_1894_n N_A_3177_368#_c_1895_n
+ N_A_3177_368#_c_1896_n PM_SKY130_FD_SC_MS__SDFSBP_2%A_3177_368#
x_PM_SKY130_FD_SC_MS__SDFSBP_2%VPWR N_VPWR_M1009_d N_VPWR_M1041_d N_VPWR_M1036_d
+ N_VPWR_M1030_d N_VPWR_M1034_d N_VPWR_M1003_s N_VPWR_M1016_d N_VPWR_M1045_d
+ N_VPWR_M1029_s N_VPWR_M1000_d N_VPWR_M1049_s N_VPWR_c_1957_n N_VPWR_c_1958_n
+ N_VPWR_c_1959_n N_VPWR_c_1960_n N_VPWR_c_1961_n N_VPWR_c_1962_n
+ N_VPWR_c_1963_n N_VPWR_c_1964_n N_VPWR_c_1965_n N_VPWR_c_1966_n
+ N_VPWR_c_1967_n N_VPWR_c_1968_n N_VPWR_c_1969_n N_VPWR_c_1970_n
+ N_VPWR_c_1971_n N_VPWR_c_1972_n N_VPWR_c_1973_n N_VPWR_c_1974_n
+ N_VPWR_c_1975_n N_VPWR_c_1976_n VPWR N_VPWR_c_1977_n N_VPWR_c_1978_n
+ N_VPWR_c_1979_n N_VPWR_c_1980_n N_VPWR_c_1981_n N_VPWR_c_1982_n
+ N_VPWR_c_1983_n N_VPWR_c_1984_n N_VPWR_c_1985_n N_VPWR_c_1986_n
+ N_VPWR_c_1987_n N_VPWR_c_1988_n N_VPWR_c_1956_n
+ PM_SKY130_FD_SC_MS__SDFSBP_2%VPWR
x_PM_SKY130_FD_SC_MS__SDFSBP_2%A_307_74# N_A_307_74#_M1038_d N_A_307_74#_M1019_s
+ N_A_307_74#_M1033_d N_A_307_74#_M1006_s N_A_307_74#_c_2157_n
+ N_A_307_74#_c_2154_n N_A_307_74#_c_2159_n N_A_307_74#_c_2160_n
+ N_A_307_74#_c_2161_n N_A_307_74#_c_2177_n N_A_307_74#_c_2195_n
+ N_A_307_74#_c_2197_n N_A_307_74#_c_2155_n N_A_307_74#_c_2162_n
+ N_A_307_74#_c_2156_n PM_SKY130_FD_SC_MS__SDFSBP_2%A_307_74#
x_PM_SKY130_FD_SC_MS__SDFSBP_2%A_1789_424# N_A_1789_424#_M1003_d
+ N_A_1789_424#_M1048_d N_A_1789_424#_M1031_s N_A_1789_424#_c_2275_n
+ N_A_1789_424#_c_2269_n N_A_1789_424#_c_2278_n N_A_1789_424#_c_2270_n
+ N_A_1789_424#_c_2271_n N_A_1789_424#_c_2272_n N_A_1789_424#_c_2273_n
+ PM_SKY130_FD_SC_MS__SDFSBP_2%A_1789_424#
x_PM_SKY130_FD_SC_MS__SDFSBP_2%A_2277_455# N_A_2277_455#_M1010_s
+ N_A_2277_455#_M1016_s N_A_2277_455#_c_2317_n N_A_2277_455#_c_2318_n
+ N_A_2277_455#_c_2319_n N_A_2277_455#_c_2320_n
+ PM_SKY130_FD_SC_MS__SDFSBP_2%A_2277_455#
x_PM_SKY130_FD_SC_MS__SDFSBP_2%Q_N N_Q_N_M1023_d N_Q_N_M1004_d N_Q_N_c_2349_n
+ Q_N Q_N Q_N N_Q_N_c_2350_n Q_N PM_SKY130_FD_SC_MS__SDFSBP_2%Q_N
x_PM_SKY130_FD_SC_MS__SDFSBP_2%Q N_Q_M1001_s N_Q_M1047_d N_Q_c_2378_n
+ N_Q_c_2379_n N_Q_c_2375_n Q Q Q PM_SKY130_FD_SC_MS__SDFSBP_2%Q
x_PM_SKY130_FD_SC_MS__SDFSBP_2%VGND N_VGND_M1044_d N_VGND_M1015_d N_VGND_M1043_d
+ N_VGND_M1024_d N_VGND_M1014_d N_VGND_M1005_d N_VGND_M1021_d N_VGND_M1023_s
+ N_VGND_M1025_s N_VGND_M1012_d N_VGND_M1022_d N_VGND_c_2406_n N_VGND_c_2407_n
+ N_VGND_c_2408_n N_VGND_c_2409_n N_VGND_c_2410_n N_VGND_c_2411_n
+ N_VGND_c_2412_n N_VGND_c_2413_n N_VGND_c_2414_n N_VGND_c_2415_n
+ N_VGND_c_2416_n N_VGND_c_2417_n N_VGND_c_2418_n N_VGND_c_2419_n
+ N_VGND_c_2420_n N_VGND_c_2421_n N_VGND_c_2422_n N_VGND_c_2423_n
+ N_VGND_c_2424_n N_VGND_c_2425_n N_VGND_c_2426_n N_VGND_c_2427_n VGND
+ N_VGND_c_2428_n N_VGND_c_2429_n N_VGND_c_2430_n N_VGND_c_2431_n
+ N_VGND_c_2432_n N_VGND_c_2433_n N_VGND_c_2434_n N_VGND_c_2435_n
+ N_VGND_c_2436_n N_VGND_c_2437_n N_VGND_c_2438_n N_VGND_c_2439_n
+ PM_SKY130_FD_SC_MS__SDFSBP_2%VGND
x_PM_SKY130_FD_SC_MS__SDFSBP_2%A_1794_74# N_A_1794_74#_M1005_s
+ N_A_1794_74#_M1011_s N_A_1794_74#_M1039_d N_A_1794_74#_c_2593_n
+ N_A_1794_74#_c_2594_n N_A_1794_74#_c_2595_n N_A_1794_74#_c_2603_n
+ N_A_1794_74#_c_2596_n N_A_1794_74#_c_2597_n N_A_1794_74#_c_2598_n
+ PM_SKY130_FD_SC_MS__SDFSBP_2%A_1794_74#
cc_1 VNB N_A_27_74#_c_357_n 0.0250407f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_2 VNB N_A_27_74#_c_358_n 0.0202447f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.97
cc_3 VNB N_A_27_74#_c_359_n 0.00761332f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.065
cc_4 VNB N_A_27_74#_c_360_n 0.0300878f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.065
cc_5 VNB N_A_27_74#_c_361_n 0.0219083f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=1.065
cc_6 VNB N_A_27_74#_c_362_n 0.0178945f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=0.9
cc_7 VNB N_SCE_M1044_g 0.0623069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_SCE_c_435_n 0.0331355f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.23
cc_9 VNB N_SCE_c_436_n 0.00270489f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=2.465
cc_10 VNB N_SCE_c_437_n 0.0319263f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=2.465
cc_11 VNB N_SCE_c_438_n 0.00219979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_SCE_c_439_n 0.0798121f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=2.055
cc_13 VNB N_SCE_c_440_n 0.00307321f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=1.975
cc_14 VNB N_SCE_c_441_n 0.0216104f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=1.975
cc_15 VNB N_D_c_512_n 0.00539996f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=0.37
cc_16 VNB N_D_M1033_g 0.00813295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_D_c_514_n 0.0190815f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=2.14
cc_18 VNB D 0.00579289f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=2.64
cc_19 VNB N_D_c_516_n 0.0316793f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_20 VNB N_D_c_517_n 0.0221915f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.23
cc_21 VNB N_SCD_M1015_g 0.0227695f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=0.58
cc_22 VNB N_SCD_c_559_n 0.0189523f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=2.64
cc_23 VNB N_SCD_c_560_n 0.00249185f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=0.9
cc_24 VNB N_SCD_c_561_n 0.0251837f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=0.58
cc_25 VNB SCD 0.00682024f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_26 VNB N_SCD_c_563_n 0.0246471f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.97
cc_27 VNB N_CLK_M1036_g 0.00768081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_CLK_c_610_n 0.0194708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB CLK 0.00951065f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=0.58
cc_30 VNB N_CLK_c_612_n 0.0566906f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=0.9
cc_31 VNB N_A_871_74#_c_646_n 0.0346908f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=2.64
cc_32 VNB N_A_871_74#_c_647_n 0.0157874f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=2.64
cc_33 VNB N_A_871_74#_M1026_g 0.0207425f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=0.58
cc_34 VNB N_A_871_74#_M1032_g 0.0204977f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.97
cc_35 VNB N_A_871_74#_M1039_g 0.0284098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_871_74#_c_651_n 0.028453f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.065
cc_37 VNB N_A_871_74#_c_652_n 0.0466008f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.065
cc_38 VNB N_A_871_74#_c_653_n 0.0332744f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.065
cc_39 VNB N_A_871_74#_M1010_g 0.00269371f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=1.065
cc_40 VNB N_A_871_74#_c_655_n 0.00620399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_871_74#_c_656_n 0.0173245f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=2.14
cc_42 VNB N_A_871_74#_c_657_n 0.00279267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_871_74#_c_658_n 0.00319375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_871_74#_c_659_n 0.0172406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_871_74#_c_660_n 0.00181342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_871_74#_c_661_n 0.0689707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_871_74#_c_662_n 0.00513279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_871_74#_c_663_n 0.00422606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_871_74#_c_664_n 2.07961e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_871_74#_c_665_n 0.00317624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_871_74#_c_666_n 0.00914437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_871_74#_c_667_n 0.0200525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_871_74#_c_668_n 0.0263125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1252_376#_c_904_n 0.0167981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1252_376#_c_905_n 0.0137517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1252_376#_c_906_n 0.00892759f $X=-0.19 $Y=-0.245 $X2=0.98
+ $Y2=1.065
cc_57 VNB N_A_1252_376#_c_907_n 0.00356983f $X=-0.19 $Y=-0.245 $X2=0.265
+ $Y2=1.065
cc_58 VNB N_A_1252_376#_c_908_n 0.0230627f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=1.975
cc_59 VNB N_A_1252_376#_c_909_n 0.0502327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1069_81#_M1042_g 0.00122075f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=0.58
cc_61 VNB N_A_1069_81#_M1013_g 0.034972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1069_81#_c_992_n 0.0250974f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=0.58
cc_63 VNB N_A_1069_81#_M1003_g 0.0181656f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.97
cc_64 VNB N_A_1069_81#_c_994_n 0.00951082f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=1.065
cc_65 VNB N_A_1069_81#_M1048_g 0.0155475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1069_81#_M1011_g 0.0215209f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=2.055
cc_67 VNB N_A_1069_81#_c_997_n 0.015267f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=1.975
cc_68 VNB N_A_1069_81#_c_998_n 0.0179261f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=1.975
cc_69 VNB N_A_1069_81#_c_999_n 0.00574168f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=2.055
cc_70 VNB N_A_1069_81#_c_1000_n 0.00683698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1069_81#_c_1001_n 0.0100682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1069_81#_c_1002_n 0.00368108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1069_81#_c_1003_n 0.00596292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1069_81#_c_1004_n 0.0124499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1069_81#_c_1005_n 0.00977247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1069_81#_c_1006_n 0.0449671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1069_81#_c_1007_n 0.0115114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1069_81#_c_1008_n 0.00148462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1069_81#_c_1009_n 0.0540624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_SET_B_M1014_g 0.0580087f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=0.9
cc_81 VNB N_SET_B_M1021_g 0.0375934f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=2.64
cc_82 VNB N_SET_B_c_1171_n 0.0107422f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.97
cc_83 VNB N_SET_B_c_1172_n 0.0186488f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=2.465
cc_84 VNB N_SET_B_c_1173_n 0.00371196f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=2.465
cc_85 VNB N_SET_B_c_1174_n 0.00210148f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.065
cc_86 VNB SET_B 6.21758e-19 $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.065
cc_87 VNB N_SET_B_c_1176_n 0.0138031f $X=-0.19 $Y=-0.245 $X2=0.465 $Y2=2.055
cc_88 VNB N_SET_B_c_1177_n 0.00454843f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=1.065
cc_89 VNB N_SET_B_c_1178_n 0.0145598f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=1.975
cc_90 VNB N_A_619_368#_M1035_g 0.0274744f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=0.58
cc_91 VNB N_A_619_368#_c_1312_n 0.0166547f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_92 VNB N_A_619_368#_c_1313_n 0.0316114f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.97
cc_93 VNB N_A_619_368#_c_1314_n 0.0104746f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=2.14
cc_94 VNB N_A_619_368#_c_1315_n 0.0184603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_619_368#_c_1316_n 0.0235315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_619_368#_c_1317_n 0.0186956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_619_368#_c_1318_n 0.0222303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_619_368#_c_1319_n 0.0127729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_619_368#_c_1320_n 0.019625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_619_368#_c_1321_n 0.00936606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_619_368#_c_1322_n 0.0563283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_619_368#_c_1323_n 0.00824969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_619_368#_c_1324_n 0.00225483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_619_368#_c_1325_n 0.00368583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_619_368#_c_1326_n 0.00775223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_619_368#_c_1327_n 0.00164982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_619_368#_c_1328_n 0.00823064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_2513_258#_M1020_g 0.0355334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_2513_258#_c_1574_n 0.0131618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_2513_258#_c_1575_n 9.9353e-19 $X=-0.19 $Y=-0.245 $X2=0.275
+ $Y2=2.465
cc_111 VNB N_A_2513_258#_c_1576_n 0.0163581f $X=-0.19 $Y=-0.245 $X2=0.3
+ $Y2=2.465
cc_112 VNB N_A_2513_258#_c_1577_n 0.02419f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=1.065
cc_113 VNB N_A_2513_258#_c_1578_n 0.00837366f $X=-0.19 $Y=-0.245 $X2=0.98
+ $Y2=1.065
cc_114 VNB N_A_2513_258#_c_1579_n 0.0101585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_2513_258#_c_1580_n 0.00752831f $X=-0.19 $Y=-0.245 $X2=0.265
+ $Y2=1.065
cc_116 VNB N_A_2513_258#_c_1581_n 0.0155466f $X=-0.19 $Y=-0.245 $X2=0.275
+ $Y2=2.055
cc_117 VNB N_A_2067_74#_M1040_g 0.0460555f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.23
cc_118 VNB N_A_2067_74#_c_1670_n 0.0471136f $X=-0.19 $Y=-0.245 $X2=0.275
+ $Y2=2.14
cc_119 VNB N_A_2067_74#_M1023_g 0.0228116f $X=-0.19 $Y=-0.245 $X2=0.465
+ $Y2=2.055
cc_120 VNB N_A_2067_74#_M1004_g 0.0122279f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=1.975
cc_121 VNB N_A_2067_74#_c_1673_n 0.0102776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_2067_74#_M1025_g 0.0233211f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=0.9
cc_123 VNB N_A_2067_74#_M1029_g 0.0136295f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=2.14
cc_124 VNB N_A_2067_74#_c_1676_n 0.058445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_2067_74#_M1000_g 0.0124376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_A_2067_74#_M1012_g 0.0258629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_A_2067_74#_c_1679_n 0.0103217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_2067_74#_c_1680_n 0.00286548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_A_2067_74#_c_1681_n 0.00286548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_A_2067_74#_c_1682_n 0.00437802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_A_2067_74#_c_1683_n 0.00783755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_A_2067_74#_c_1684_n 0.0118908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_A_2067_74#_c_1685_n 8.34101e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_A_2067_74#_c_1686_n 0.0137219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_A_2067_74#_c_1687_n 0.00231564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_A_2067_74#_c_1688_n 0.00535782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_A_3177_368#_M1047_g 0.00169308f $X=-0.19 $Y=-0.245 $X2=1.07
+ $Y2=0.58
cc_138 VNB N_A_3177_368#_M1001_g 0.0228691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_A_3177_368#_M1049_g 0.00231818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_A_3177_368#_M1022_g 0.0260188f $X=-0.19 $Y=-0.245 $X2=0.275
+ $Y2=2.465
cc_141 VNB N_A_3177_368#_c_1892_n 0.0120685f $X=-0.19 $Y=-0.245 $X2=0.98
+ $Y2=1.065
cc_142 VNB N_A_3177_368#_c_1893_n 5.42215e-19 $X=-0.19 $Y=-0.245 $X2=1.775
+ $Y2=2.055
cc_143 VNB N_A_3177_368#_c_1894_n 0.00904052f $X=-0.19 $Y=-0.245 $X2=1.94
+ $Y2=1.975
cc_144 VNB N_A_3177_368#_c_1895_n 0.00280955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_A_3177_368#_c_1896_n 0.0662175f $X=-0.19 $Y=-0.245 $X2=1.94
+ $Y2=1.975
cc_146 VNB N_VPWR_c_1956_n 0.740851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_A_307_74#_c_2154_n 0.00882071f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.23
cc_148 VNB N_A_307_74#_c_2155_n 0.0035679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_A_307_74#_c_2156_n 0.00556247f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=0.9
cc_150 VNB N_Q_N_c_2349_n 0.00204548f $X=-0.19 $Y=-0.245 $X2=1.07 $Y2=0.58
cc_151 VNB N_Q_N_c_2350_n 0.00257348f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=2.465
cc_152 VNB N_Q_c_2375_n 0.00141953f $X=-0.19 $Y=-0.245 $X2=0.265 $Y2=0.58
cc_153 VNB Q 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_154 VNB Q 0.00429087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2406_n 0.00723643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2407_n 0.00970665f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=0.9
cc_157 VNB N_VGND_c_2408_n 0.0054384f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=2.14
cc_158 VNB N_VGND_c_2409_n 0.0152393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_2410_n 0.00953882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_2411_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_VGND_c_2412_n 0.00860026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VNB N_VGND_c_2413_n 0.0144665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_VGND_c_2414_n 0.0217072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VNB N_VGND_c_2415_n 0.0146831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_VGND_c_2416_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_VGND_c_2417_n 0.0505285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_VGND_c_2418_n 0.0506538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_VGND_c_2419_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_169 VNB N_VGND_c_2420_n 0.0271172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_170 VNB N_VGND_c_2421_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_VGND_c_2422_n 0.0911645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_172 VNB N_VGND_c_2423_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_173 VNB N_VGND_c_2424_n 0.0215588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_174 VNB N_VGND_c_2425_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_175 VNB N_VGND_c_2426_n 0.0199954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_176 VNB N_VGND_c_2427_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_177 VNB N_VGND_c_2428_n 0.0189171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_178 VNB N_VGND_c_2429_n 0.018606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_179 VNB N_VGND_c_2430_n 0.0671019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_180 VNB N_VGND_c_2431_n 0.0306291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_181 VNB N_VGND_c_2432_n 0.0231281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_182 VNB N_VGND_c_2433_n 0.0192531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_183 VNB N_VGND_c_2434_n 0.00760052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_184 VNB N_VGND_c_2435_n 0.00615422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_185 VNB N_VGND_c_2436_n 0.00644364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_186 VNB N_VGND_c_2437_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_187 VNB N_VGND_c_2438_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_188 VNB N_VGND_c_2439_n 0.99539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_189 VNB N_A_1794_74#_c_2593_n 0.00270668f $X=-0.19 $Y=-0.245 $X2=2.015
+ $Y2=2.64
cc_190 VNB N_A_1794_74#_c_2594_n 0.00449539f $X=-0.19 $Y=-0.245 $X2=0.265
+ $Y2=0.9
cc_191 VNB N_A_1794_74#_c_2595_n 4.59673e-19 $X=-0.19 $Y=-0.245 $X2=0.265
+ $Y2=0.58
cc_192 VNB N_A_1794_74#_c_2596_n 0.00313507f $X=-0.19 $Y=-0.245 $X2=0.275
+ $Y2=2.14
cc_193 VNB N_A_1794_74#_c_2597_n 0.00251555f $X=-0.19 $Y=-0.245 $X2=0.275
+ $Y2=2.465
cc_194 VNB N_A_1794_74#_c_2598_n 0.0118588f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=2.465
cc_195 VPB N_A_27_74#_M1027_g 0.0242712f $X=-0.19 $Y=1.66 $X2=2.015 $Y2=2.64
cc_196 VPB N_A_27_74#_c_358_n 0.0147344f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.97
cc_197 VPB N_A_27_74#_c_365_n 0.0376841f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=2.465
cc_198 VPB N_A_27_74#_c_366_n 0.0226472f $X=-0.19 $Y=1.66 $X2=1.775 $Y2=2.055
cc_199 VPB N_A_27_74#_c_367_n 0.0146808f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=2.055
cc_200 VPB N_A_27_74#_c_368_n 0.00434281f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=1.975
cc_201 VPB N_A_27_74#_c_369_n 0.0335867f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=1.975
cc_202 VPB N_SCE_M1009_g 0.0509437f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.9
cc_203 VPB N_SCE_M1007_g 0.0397602f $X=-0.19 $Y=1.66 $X2=2.015 $Y2=2.64
cc_204 VPB N_SCE_c_437_n 0.0205042f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=2.465
cc_205 VPB N_D_M1033_g 0.0530383f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_SCD_M1041_g 0.0376738f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_SCD_c_565_n 0.025822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_SCD_c_566_n 0.00933483f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_SCD_c_560_n 0.0094824f $X=-0.19 $Y=1.66 $X2=0.265 $Y2=0.9
cc_210 VPB N_CLK_M1036_g 0.0282941f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_871_74#_M1006_g 0.0332501f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.58
cc_212 VPB N_A_871_74#_M1010_g 0.0487799f $X=-0.19 $Y=1.66 $X2=0.265 $Y2=1.065
cc_213 VPB N_A_871_74#_c_671_n 0.017836f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=1.975
cc_214 VPB N_A_871_74#_c_672_n 0.00349515f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=1.975
cc_215 VPB N_A_871_74#_c_673_n 0.0217529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_871_74#_c_674_n 0.00388103f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_871_74#_c_658_n 0.00209765f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_871_74#_c_659_n 0.0105641f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_871_74#_c_660_n 0.00588447f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_871_74#_c_678_n 0.00281843f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_871_74#_c_679_n 0.0116167f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_871_74#_c_680_n 0.00424643f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_871_74#_c_681_n 0.0158111f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_871_74#_c_682_n 0.00260538f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_871_74#_c_683_n 0.00310194f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_871_74#_c_684_n 0.0138834f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_871_74#_c_685_n 4.80289e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_871_74#_c_662_n 0.0077675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_871_74#_c_687_n 9.12633e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_1252_376#_M1030_g 0.0332882f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.58
cc_231 VPB N_A_1252_376#_c_911_n 0.012809f $X=-0.19 $Y=1.66 $X2=2.015 $Y2=2.64
cc_232 VPB N_A_1252_376#_c_912_n 0.0123547f $X=-0.19 $Y=1.66 $X2=2.015 $Y2=2.64
cc_233 VPB N_A_1252_376#_c_913_n 0.0122171f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.23
cc_234 VPB N_A_1252_376#_c_914_n 0.0357008f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=2.465
cc_235 VPB N_A_1252_376#_c_915_n 0.00675698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_1252_376#_c_916_n 0.00243407f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.065
cc_237 VPB N_A_1252_376#_c_908_n 0.00261721f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=1.975
cc_238 VPB N_A_1069_81#_M1042_g 0.0516506f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.58
cc_239 VPB N_A_1069_81#_M1003_g 0.0362558f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.97
cc_240 VPB N_A_1069_81#_M1048_g 0.0397596f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_A_1069_81#_c_1013_n 0.00824141f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_A_1069_81#_c_1007_n 0.0108554f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_SET_B_M1034_g 0.0397755f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_SET_B_M1018_g 0.0496978f $X=-0.19 $Y=1.66 $X2=0.265 $Y2=0.58
cc_245 VPB N_SET_B_c_1171_n 0.0079736f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.97
cc_246 VPB N_SET_B_c_1182_n 0.0130201f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=2.14
cc_247 VPB N_SET_B_c_1172_n 0.0112351f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=2.465
cc_248 VPB N_SET_B_c_1173_n 0.0024764f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=2.465
cc_249 VPB N_SET_B_c_1174_n 0.00529978f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.065
cc_250 VPB SET_B 6.00473e-19 $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.065
cc_251 VPB N_SET_B_c_1177_n 0.00391415f $X=-0.19 $Y=1.66 $X2=0.265 $Y2=1.065
cc_252 VPB N_SET_B_c_1178_n 0.0196655f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=1.975
cc_253 VPB N_A_619_368#_M1046_g 0.0247851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_A_619_368#_c_1330_n 0.0757111f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.23
cc_255 VPB N_A_619_368#_c_1331_n 0.0600669f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=2.465
cc_256 VPB N_A_619_368#_c_1332_n 0.0123872f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=2.465
cc_257 VPB N_A_619_368#_M1002_g 0.0388891f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_A_619_368#_c_1334_n 0.210354f $X=-0.19 $Y=1.66 $X2=0.465 $Y2=2.055
cc_259 VPB N_A_619_368#_c_1335_n 0.0738062f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=1.975
cc_260 VPB N_A_619_368#_c_1336_n 0.0157699f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=1.975
cc_261 VPB N_A_619_368#_c_1337_n 0.0121871f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=2.055
cc_262 VPB N_A_619_368#_c_1338_n 0.0107697f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_A_619_368#_c_1339_n 0.0159298f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.065
cc_264 VPB N_A_619_368#_c_1340_n 0.0260476f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=1.975
cc_265 VPB N_A_619_368#_c_1341_n 0.057228f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_A_619_368#_c_1342_n 0.0711477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_A_619_368#_c_1343_n 0.0122279f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_A_619_368#_c_1317_n 0.071851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_A_619_368#_c_1319_n 0.00101684f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_A_619_368#_c_1320_n 0.00682721f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_A_619_368#_c_1321_n 6.04262e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_A_619_368#_c_1348_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_A_619_368#_c_1349_n 0.00637368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_A_619_368#_c_1350_n 0.00773831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_A_619_368#_c_1325_n 0.00170449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_A_619_368#_c_1352_n 0.0402381f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_A_619_368#_c_1353_n 0.0113817f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_A_619_368#_c_1328_n 0.027905f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_A_619_368#_c_1355_n 0.00113419f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_A_2513_258#_M1016_g 0.0457138f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.58
cc_281 VPB N_A_2513_258#_c_1574_n 0.00827326f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_A_2513_258#_c_1584_n 0.0153617f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.23
cc_283 VPB N_A_2513_258#_c_1575_n 0.00137888f $X=-0.19 $Y=1.66 $X2=0.275
+ $Y2=2.465
cc_284 VPB N_A_2513_258#_c_1580_n 0.0114425f $X=-0.19 $Y=1.66 $X2=0.265
+ $Y2=1.065
cc_285 VPB N_A_2513_258#_c_1587_n 0.00686537f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_286 VPB N_A_2067_74#_c_1689_n 0.0251978f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=2.465
cc_287 VPB N_A_2067_74#_c_1690_n 0.0225675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_288 VPB N_A_2067_74#_M1045_g 0.0251815f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.065
cc_289 VPB N_A_2067_74#_M1004_g 0.0238838f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=1.975
cc_290 VPB N_A_2067_74#_M1029_g 0.025985f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=2.14
cc_291 VPB N_A_2067_74#_M1000_g 0.026762f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_292 VPB N_A_2067_74#_c_1695_n 0.0093495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_293 VPB N_A_2067_74#_c_1696_n 0.00234531f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_294 VPB N_A_2067_74#_c_1697_n 0.0152136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_295 VPB N_A_2067_74#_c_1698_n 0.0103269f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_296 VPB N_A_2067_74#_c_1699_n 0.00884139f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_297 VPB N_A_2067_74#_c_1686_n 0.0363227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_298 VPB N_A_2067_74#_c_1701_n 0.006122f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_299 VPB N_A_2067_74#_c_1688_n 0.00248742f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_300 VPB N_A_3177_368#_M1047_g 0.0239925f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.58
cc_301 VPB N_A_3177_368#_M1049_g 0.0274022f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_302 VPB N_A_3177_368#_c_1893_n 0.0154468f $X=-0.19 $Y=1.66 $X2=1.775
+ $Y2=2.055
cc_303 VPB N_VPWR_c_1957_n 0.00893346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_304 VPB N_VPWR_c_1958_n 0.0121232f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=0.9
cc_305 VPB N_VPWR_c_1959_n 0.00693022f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_306 VPB N_VPWR_c_1960_n 0.0313096f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_307 VPB N_VPWR_c_1961_n 0.0111242f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_308 VPB N_VPWR_c_1962_n 0.00521506f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_309 VPB N_VPWR_c_1963_n 0.00979595f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_310 VPB N_VPWR_c_1964_n 0.0127208f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_311 VPB N_VPWR_c_1965_n 0.0263703f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_312 VPB N_VPWR_c_1966_n 0.0156914f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_313 VPB N_VPWR_c_1967_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_314 VPB N_VPWR_c_1968_n 0.0644823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_315 VPB N_VPWR_c_1969_n 0.020354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_316 VPB N_VPWR_c_1970_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_317 VPB N_VPWR_c_1971_n 0.0794393f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_318 VPB N_VPWR_c_1972_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_319 VPB N_VPWR_c_1973_n 0.0380992f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_320 VPB N_VPWR_c_1974_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_321 VPB N_VPWR_c_1975_n 0.0184862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_322 VPB N_VPWR_c_1976_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_323 VPB N_VPWR_c_1977_n 0.0193973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_324 VPB N_VPWR_c_1978_n 0.0448083f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_325 VPB N_VPWR_c_1979_n 0.0507274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_326 VPB N_VPWR_c_1980_n 0.0227335f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_327 VPB N_VPWR_c_1981_n 0.0203698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_328 VPB N_VPWR_c_1982_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_329 VPB N_VPWR_c_1983_n 0.00651209f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_330 VPB N_VPWR_c_1984_n 0.0214164f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_331 VPB N_VPWR_c_1985_n 0.0200392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_332 VPB N_VPWR_c_1986_n 0.00763133f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_333 VPB N_VPWR_c_1987_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_334 VPB N_VPWR_c_1988_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_335 VPB N_VPWR_c_1956_n 0.150001f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_336 VPB N_A_307_74#_c_2157_n 0.00824485f $X=-0.19 $Y=1.66 $X2=0.265 $Y2=0.58
cc_337 VPB N_A_307_74#_c_2154_n 0.0147808f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.23
cc_338 VPB N_A_307_74#_c_2159_n 0.0121196f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.97
cc_339 VPB N_A_307_74#_c_2160_n 0.00312412f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=2.465
cc_340 VPB N_A_307_74#_c_2161_n 0.00653294f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.065
cc_341 VPB N_A_307_74#_c_2162_n 0.0102155f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.065
cc_342 VPB N_A_307_74#_c_2156_n 0.00306764f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=0.9
cc_343 VPB N_A_1789_424#_c_2269_n 0.00217381f $X=-0.19 $Y=1.66 $X2=0.265 $Y2=0.9
cc_344 VPB N_A_1789_424#_c_2270_n 0.00623414f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_345 VPB N_A_1789_424#_c_2271_n 0.00160153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_346 VPB N_A_1789_424#_c_2272_n 0.00407868f $X=-0.19 $Y=1.66 $X2=0.275
+ $Y2=2.14
cc_347 VPB N_A_1789_424#_c_2273_n 0.0102478f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_348 VPB N_A_2277_455#_c_2317_n 0.00752457f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.58
cc_349 VPB N_A_2277_455#_c_2318_n 0.0144652f $X=-0.19 $Y=1.66 $X2=2.015 $Y2=2.64
cc_350 VPB N_A_2277_455#_c_2319_n 0.00404548f $X=-0.19 $Y=1.66 $X2=2.015
+ $Y2=2.64
cc_351 VPB N_A_2277_455#_c_2320_n 0.00577049f $X=-0.19 $Y=1.66 $X2=0.265
+ $Y2=0.58
cc_352 VPB N_Q_N_c_2349_n 0.0039248f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.58
cc_353 VPB N_Q_c_2378_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.07 $Y2=0.58
cc_354 VPB N_Q_c_2379_n 0.00447264f $X=-0.19 $Y=1.66 $X2=0.265 $Y2=0.9
cc_355 VPB N_Q_c_2375_n 0.0010488f $X=-0.19 $Y=1.66 $X2=0.265 $Y2=0.58
cc_356 N_A_27_74#_c_357_n N_SCE_M1044_g 0.011453f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_357 N_A_27_74#_c_358_n N_SCE_M1044_g 0.00547238f $X=0.17 $Y=1.97 $X2=0 $Y2=0
cc_358 N_A_27_74#_c_359_n N_SCE_M1044_g 0.0146918f $X=0.98 $Y=1.065 $X2=0 $Y2=0
cc_359 N_A_27_74#_c_360_n N_SCE_M1044_g 0.0176381f $X=0.98 $Y=1.065 $X2=0 $Y2=0
cc_360 N_A_27_74#_c_361_n N_SCE_M1044_g 0.00812645f $X=0.265 $Y=1.065 $X2=0
+ $Y2=0
cc_361 N_A_27_74#_c_362_n N_SCE_M1044_g 0.0119253f $X=0.98 $Y=0.9 $X2=0 $Y2=0
cc_362 N_A_27_74#_c_358_n N_SCE_M1009_g 0.00413205f $X=0.17 $Y=1.97 $X2=0 $Y2=0
cc_363 N_A_27_74#_c_365_n N_SCE_M1009_g 0.0153596f $X=0.3 $Y=2.465 $X2=0 $Y2=0
cc_364 N_A_27_74#_c_366_n N_SCE_M1009_g 0.0132272f $X=1.775 $Y=2.055 $X2=0 $Y2=0
cc_365 N_A_27_74#_c_367_n N_SCE_M1009_g 0.00446031f $X=0.275 $Y=2.055 $X2=0
+ $Y2=0
cc_366 N_A_27_74#_c_365_n N_SCE_M1007_g 9.63487e-19 $X=0.3 $Y=2.465 $X2=0 $Y2=0
cc_367 N_A_27_74#_c_366_n N_SCE_M1007_g 0.0164772f $X=1.775 $Y=2.055 $X2=0 $Y2=0
cc_368 N_A_27_74#_c_366_n N_SCE_c_435_n 0.0272489f $X=1.775 $Y=2.055 $X2=0 $Y2=0
cc_369 N_A_27_74#_c_368_n N_SCE_c_435_n 0.0194177f $X=1.94 $Y=1.975 $X2=0 $Y2=0
cc_370 N_A_27_74#_c_369_n N_SCE_c_435_n 0.00140807f $X=1.94 $Y=1.975 $X2=0 $Y2=0
cc_371 N_A_27_74#_c_358_n N_SCE_c_436_n 0.0317203f $X=0.17 $Y=1.97 $X2=0 $Y2=0
cc_372 N_A_27_74#_c_359_n N_SCE_c_436_n 0.0563109f $X=0.98 $Y=1.065 $X2=0 $Y2=0
cc_373 N_A_27_74#_c_360_n N_SCE_c_436_n 0.00277723f $X=0.98 $Y=1.065 $X2=0 $Y2=0
cc_374 N_A_27_74#_c_366_n N_SCE_c_436_n 0.0460993f $X=1.775 $Y=2.055 $X2=0 $Y2=0
cc_375 N_A_27_74#_c_361_n N_SCE_c_436_n 0.00161902f $X=0.265 $Y=1.065 $X2=0
+ $Y2=0
cc_376 N_A_27_74#_c_367_n N_SCE_c_436_n 0.00328312f $X=0.275 $Y=2.055 $X2=0
+ $Y2=0
cc_377 N_A_27_74#_c_358_n N_SCE_c_437_n 0.00871649f $X=0.17 $Y=1.97 $X2=0 $Y2=0
cc_378 N_A_27_74#_c_359_n N_SCE_c_437_n 0.00180003f $X=0.98 $Y=1.065 $X2=0 $Y2=0
cc_379 N_A_27_74#_c_360_n N_SCE_c_437_n 0.0153046f $X=0.98 $Y=1.065 $X2=0 $Y2=0
cc_380 N_A_27_74#_c_366_n N_SCE_c_437_n 0.00313888f $X=1.775 $Y=2.055 $X2=0
+ $Y2=0
cc_381 N_A_27_74#_c_361_n N_SCE_c_437_n 2.0611e-19 $X=0.265 $Y=1.065 $X2=0 $Y2=0
cc_382 N_A_27_74#_c_367_n N_SCE_c_437_n 7.36532e-19 $X=0.275 $Y=2.055 $X2=0
+ $Y2=0
cc_383 N_A_27_74#_c_369_n N_SCE_c_439_n 0.007769f $X=1.94 $Y=1.975 $X2=0 $Y2=0
cc_384 N_A_27_74#_M1027_g N_D_M1033_g 0.0116574f $X=2.015 $Y=2.64 $X2=0 $Y2=0
cc_385 N_A_27_74#_c_366_n N_D_M1033_g 0.0172611f $X=1.775 $Y=2.055 $X2=0 $Y2=0
cc_386 N_A_27_74#_c_368_n N_D_M1033_g 0.00116992f $X=1.94 $Y=1.975 $X2=0 $Y2=0
cc_387 N_A_27_74#_c_369_n N_D_M1033_g 0.0183745f $X=1.94 $Y=1.975 $X2=0 $Y2=0
cc_388 N_A_27_74#_c_359_n D 0.0201653f $X=0.98 $Y=1.065 $X2=0 $Y2=0
cc_389 N_A_27_74#_c_360_n D 4.18339e-19 $X=0.98 $Y=1.065 $X2=0 $Y2=0
cc_390 N_A_27_74#_c_362_n D 0.00225318f $X=0.98 $Y=0.9 $X2=0 $Y2=0
cc_391 N_A_27_74#_c_359_n N_D_c_516_n 0.00120526f $X=0.98 $Y=1.065 $X2=0 $Y2=0
cc_392 N_A_27_74#_c_360_n N_D_c_516_n 0.0255527f $X=0.98 $Y=1.065 $X2=0 $Y2=0
cc_393 N_A_27_74#_c_362_n N_D_c_517_n 0.0255527f $X=0.98 $Y=0.9 $X2=0 $Y2=0
cc_394 N_A_27_74#_M1027_g N_SCD_M1041_g 0.0340337f $X=2.015 $Y=2.64 $X2=0 $Y2=0
cc_395 N_A_27_74#_c_368_n N_SCD_c_566_n 0.00128345f $X=1.94 $Y=1.975 $X2=0 $Y2=0
cc_396 N_A_27_74#_c_369_n N_SCD_c_566_n 0.0340337f $X=1.94 $Y=1.975 $X2=0 $Y2=0
cc_397 N_A_27_74#_c_365_n N_VPWR_c_1957_n 0.0268536f $X=0.3 $Y=2.465 $X2=0 $Y2=0
cc_398 N_A_27_74#_c_366_n N_VPWR_c_1957_n 0.0274627f $X=1.775 $Y=2.055 $X2=0
+ $Y2=0
cc_399 N_A_27_74#_M1027_g N_VPWR_c_1958_n 0.00147831f $X=2.015 $Y=2.64 $X2=0
+ $Y2=0
cc_400 N_A_27_74#_c_365_n N_VPWR_c_1977_n 0.01678f $X=0.3 $Y=2.465 $X2=0 $Y2=0
cc_401 N_A_27_74#_M1027_g N_VPWR_c_1978_n 0.005209f $X=2.015 $Y=2.64 $X2=0 $Y2=0
cc_402 N_A_27_74#_M1027_g N_VPWR_c_1956_n 0.00537464f $X=2.015 $Y=2.64 $X2=0
+ $Y2=0
cc_403 N_A_27_74#_c_365_n N_VPWR_c_1956_n 0.0138209f $X=0.3 $Y=2.465 $X2=0 $Y2=0
cc_404 N_A_27_74#_M1027_g N_A_307_74#_c_2157_n 0.00956751f $X=2.015 $Y=2.64
+ $X2=0 $Y2=0
cc_405 N_A_27_74#_c_368_n N_A_307_74#_c_2157_n 0.0106621f $X=1.94 $Y=1.975 $X2=0
+ $Y2=0
cc_406 N_A_27_74#_c_368_n N_A_307_74#_c_2154_n 0.0128835f $X=1.94 $Y=1.975 $X2=0
+ $Y2=0
cc_407 N_A_27_74#_c_369_n N_A_307_74#_c_2154_n 0.00188419f $X=1.94 $Y=1.975
+ $X2=0 $Y2=0
cc_408 N_A_27_74#_M1027_g N_A_307_74#_c_2161_n 0.0109565f $X=2.015 $Y=2.64 $X2=0
+ $Y2=0
cc_409 N_A_27_74#_c_366_n N_A_307_74#_c_2161_n 0.0225281f $X=1.775 $Y=2.055
+ $X2=0 $Y2=0
cc_410 N_A_27_74#_c_368_n N_A_307_74#_c_2161_n 0.0150159f $X=1.94 $Y=1.975 $X2=0
+ $Y2=0
cc_411 N_A_27_74#_c_369_n N_A_307_74#_c_2161_n 0.00117194f $X=1.94 $Y=1.975
+ $X2=0 $Y2=0
cc_412 N_A_27_74#_c_357_n N_VGND_c_2406_n 0.0133638f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_413 N_A_27_74#_c_359_n N_VGND_c_2406_n 0.0255027f $X=0.98 $Y=1.065 $X2=0
+ $Y2=0
cc_414 N_A_27_74#_c_360_n N_VGND_c_2406_n 0.0038848f $X=0.98 $Y=1.065 $X2=0
+ $Y2=0
cc_415 N_A_27_74#_c_362_n N_VGND_c_2406_n 0.00981126f $X=0.98 $Y=0.9 $X2=0 $Y2=0
cc_416 N_A_27_74#_c_362_n N_VGND_c_2418_n 0.00383152f $X=0.98 $Y=0.9 $X2=0 $Y2=0
cc_417 N_A_27_74#_c_357_n N_VGND_c_2428_n 0.0159025f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_418 N_A_27_74#_c_357_n N_VGND_c_2439_n 0.0131064f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_419 N_A_27_74#_c_362_n N_VGND_c_2439_n 0.0075725f $X=0.98 $Y=0.9 $X2=0 $Y2=0
cc_420 N_SCE_c_435_n N_D_c_512_n 0.00445951f $X=1.965 $Y=1.485 $X2=-0.19
+ $Y2=-0.245
cc_421 N_SCE_c_437_n N_D_c_512_n 0.00828205f $X=0.92 $Y=1.635 $X2=-0.19
+ $Y2=-0.245
cc_422 N_SCE_c_435_n N_D_M1033_g 0.00429479f $X=1.965 $Y=1.485 $X2=0 $Y2=0
cc_423 N_SCE_c_437_n N_D_M1033_g 0.078215f $X=0.92 $Y=1.635 $X2=0 $Y2=0
cc_424 N_SCE_c_438_n N_D_M1033_g 0.0014191f $X=1.085 $Y=1.6 $X2=0 $Y2=0
cc_425 N_SCE_c_435_n N_D_c_514_n 0.00572304f $X=1.965 $Y=1.485 $X2=0 $Y2=0
cc_426 N_SCE_c_439_n N_D_c_514_n 0.00964743f $X=2.13 $Y=1.065 $X2=0 $Y2=0
cc_427 N_SCE_c_440_n N_D_c_514_n 9.50384e-19 $X=2.13 $Y=1.065 $X2=0 $Y2=0
cc_428 N_SCE_c_435_n D 0.0324073f $X=1.965 $Y=1.485 $X2=0 $Y2=0
cc_429 N_SCE_c_439_n D 0.00220222f $X=2.13 $Y=1.065 $X2=0 $Y2=0
cc_430 N_SCE_c_440_n D 0.0265741f $X=2.13 $Y=1.065 $X2=0 $Y2=0
cc_431 N_SCE_c_441_n D 0.00241363f $X=2.22 $Y=0.9 $X2=0 $Y2=0
cc_432 N_SCE_c_435_n N_D_c_516_n 0.00126891f $X=1.965 $Y=1.485 $X2=0 $Y2=0
cc_433 N_SCE_c_439_n N_D_c_516_n 0.0170267f $X=2.13 $Y=1.065 $X2=0 $Y2=0
cc_434 N_SCE_c_440_n N_D_c_516_n 3.60471e-19 $X=2.13 $Y=1.065 $X2=0 $Y2=0
cc_435 N_SCE_c_439_n N_SCD_c_566_n 0.00945859f $X=2.13 $Y=1.065 $X2=0 $Y2=0
cc_436 N_SCE_c_441_n N_SCD_M1015_g 0.0341499f $X=2.22 $Y=0.9 $X2=0 $Y2=0
cc_437 N_SCE_c_439_n N_SCD_c_559_n 0.0341499f $X=2.13 $Y=1.065 $X2=0 $Y2=0
cc_438 N_SCE_c_439_n SCD 5.07628e-19 $X=2.13 $Y=1.065 $X2=0 $Y2=0
cc_439 N_SCE_M1009_g N_VPWR_c_1957_n 0.00343158f $X=0.525 $Y=2.64 $X2=0 $Y2=0
cc_440 N_SCE_M1007_g N_VPWR_c_1957_n 0.0170614f $X=1.025 $Y=2.64 $X2=0 $Y2=0
cc_441 N_SCE_M1009_g N_VPWR_c_1977_n 0.005209f $X=0.525 $Y=2.64 $X2=0 $Y2=0
cc_442 N_SCE_M1007_g N_VPWR_c_1978_n 0.00460063f $X=1.025 $Y=2.64 $X2=0 $Y2=0
cc_443 N_SCE_M1009_g N_VPWR_c_1956_n 0.00985891f $X=0.525 $Y=2.64 $X2=0 $Y2=0
cc_444 N_SCE_M1007_g N_VPWR_c_1956_n 0.00908371f $X=1.025 $Y=2.64 $X2=0 $Y2=0
cc_445 N_SCE_c_435_n N_A_307_74#_c_2154_n 0.0129498f $X=1.965 $Y=1.485 $X2=0
+ $Y2=0
cc_446 N_SCE_c_439_n N_A_307_74#_c_2154_n 0.0142897f $X=2.13 $Y=1.065 $X2=0
+ $Y2=0
cc_447 N_SCE_c_440_n N_A_307_74#_c_2154_n 0.0356688f $X=2.13 $Y=1.065 $X2=0
+ $Y2=0
cc_448 N_SCE_c_441_n N_A_307_74#_c_2154_n 0.00470988f $X=2.22 $Y=0.9 $X2=0 $Y2=0
cc_449 N_SCE_M1007_g N_A_307_74#_c_2161_n 0.00189358f $X=1.025 $Y=2.64 $X2=0
+ $Y2=0
cc_450 N_SCE_c_439_n N_A_307_74#_c_2177_n 0.00233988f $X=2.13 $Y=1.065 $X2=0
+ $Y2=0
cc_451 N_SCE_c_440_n N_A_307_74#_c_2177_n 0.0260811f $X=2.13 $Y=1.065 $X2=0
+ $Y2=0
cc_452 N_SCE_c_441_n N_A_307_74#_c_2177_n 0.0150729f $X=2.22 $Y=0.9 $X2=0 $Y2=0
cc_453 N_SCE_M1044_g N_VGND_c_2406_n 0.00540268f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_454 N_SCE_c_441_n N_VGND_c_2407_n 0.00144244f $X=2.22 $Y=0.9 $X2=0 $Y2=0
cc_455 N_SCE_c_441_n N_VGND_c_2418_n 0.00314477f $X=2.22 $Y=0.9 $X2=0 $Y2=0
cc_456 N_SCE_M1044_g N_VGND_c_2428_n 0.00434272f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_457 N_SCE_M1044_g N_VGND_c_2439_n 0.00825006f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_458 N_SCE_c_441_n N_VGND_c_2439_n 0.00395526f $X=2.22 $Y=0.9 $X2=0 $Y2=0
cc_459 N_D_M1033_g N_VPWR_c_1957_n 0.00244273f $X=1.445 $Y=2.64 $X2=0 $Y2=0
cc_460 N_D_M1033_g N_VPWR_c_1978_n 0.005209f $X=1.445 $Y=2.64 $X2=0 $Y2=0
cc_461 N_D_M1033_g N_VPWR_c_1956_n 0.00984319f $X=1.445 $Y=2.64 $X2=0 $Y2=0
cc_462 D N_A_307_74#_M1038_d 0.00795735f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_463 D N_A_307_74#_c_2154_n 0.00450433f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_464 N_D_M1033_g N_A_307_74#_c_2161_n 0.0135292f $X=1.445 $Y=2.64 $X2=0 $Y2=0
cc_465 D N_A_307_74#_c_2177_n 0.0246293f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_466 N_D_c_517_n N_A_307_74#_c_2177_n 0.00242613f $X=1.55 $Y=0.9 $X2=0 $Y2=0
cc_467 D N_VGND_c_2406_n 0.0100693f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_468 N_D_c_517_n N_VGND_c_2406_n 0.00163952f $X=1.55 $Y=0.9 $X2=0 $Y2=0
cc_469 D N_VGND_c_2418_n 0.0118305f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_470 N_D_c_517_n N_VGND_c_2418_n 0.00304348f $X=1.55 $Y=0.9 $X2=0 $Y2=0
cc_471 D N_VGND_c_2439_n 0.0134831f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_472 N_D_c_517_n N_VGND_c_2439_n 0.00375359f $X=1.55 $Y=0.9 $X2=0 $Y2=0
cc_473 N_SCD_c_560_n N_CLK_M1036_g 0.00609219f $X=2.79 $Y=1.81 $X2=0 $Y2=0
cc_474 N_SCD_c_561_n N_CLK_M1036_g 0.0108696f $X=2.925 $Y=1.62 $X2=0 $Y2=0
cc_475 N_SCD_c_563_n N_CLK_c_610_n 0.00312834f $X=2.97 $Y=1.115 $X2=0 $Y2=0
cc_476 N_SCD_c_559_n N_CLK_c_612_n 0.0108696f $X=2.925 $Y=1.41 $X2=0 $Y2=0
cc_477 SCD N_CLK_c_612_n 0.00259806f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_478 N_SCD_M1015_g N_A_619_368#_c_1323_n 0.00509351f $X=2.79 $Y=0.58 $X2=0
+ $Y2=0
cc_479 N_SCD_c_559_n N_A_619_368#_c_1324_n 8.82504e-19 $X=2.925 $Y=1.41 $X2=0
+ $Y2=0
cc_480 N_SCD_c_560_n N_A_619_368#_c_1324_n 9.07157e-19 $X=2.79 $Y=1.81 $X2=0
+ $Y2=0
cc_481 N_SCD_M1041_g N_A_619_368#_c_1353_n 9.69705e-19 $X=2.435 $Y=2.64 $X2=0
+ $Y2=0
cc_482 N_SCD_c_560_n N_A_619_368#_c_1353_n 0.00224001f $X=2.79 $Y=1.81 $X2=0
+ $Y2=0
cc_483 N_SCD_c_561_n N_A_619_368#_c_1353_n 0.0015818f $X=2.925 $Y=1.62 $X2=0
+ $Y2=0
cc_484 SCD N_A_619_368#_c_1353_n 0.011212f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_485 SCD N_A_619_368#_c_1327_n 0.0526178f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_486 N_SCD_c_563_n N_A_619_368#_c_1327_n 4.41357e-19 $X=2.97 $Y=1.115 $X2=0
+ $Y2=0
cc_487 N_SCD_M1041_g N_VPWR_c_1958_n 0.0118374f $X=2.435 $Y=2.64 $X2=0 $Y2=0
cc_488 N_SCD_c_565_n N_VPWR_c_1958_n 5.1142e-19 $X=2.715 $Y=1.885 $X2=0 $Y2=0
cc_489 N_SCD_M1041_g N_VPWR_c_1978_n 0.00460063f $X=2.435 $Y=2.64 $X2=0 $Y2=0
cc_490 N_SCD_M1041_g N_VPWR_c_1956_n 0.00463131f $X=2.435 $Y=2.64 $X2=0 $Y2=0
cc_491 N_SCD_M1041_g N_A_307_74#_c_2157_n 0.0113443f $X=2.435 $Y=2.64 $X2=0
+ $Y2=0
cc_492 N_SCD_M1041_g N_A_307_74#_c_2154_n 0.0121985f $X=2.435 $Y=2.64 $X2=0
+ $Y2=0
cc_493 N_SCD_c_565_n N_A_307_74#_c_2154_n 0.00921263f $X=2.715 $Y=1.885 $X2=0
+ $Y2=0
cc_494 N_SCD_c_566_n N_A_307_74#_c_2154_n 0.00396493f $X=2.525 $Y=1.885 $X2=0
+ $Y2=0
cc_495 N_SCD_M1015_g N_A_307_74#_c_2154_n 0.0167474f $X=2.79 $Y=0.58 $X2=0 $Y2=0
cc_496 SCD N_A_307_74#_c_2154_n 0.0511176f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_497 N_SCD_c_565_n N_A_307_74#_c_2159_n 0.00737458f $X=2.715 $Y=1.885 $X2=0
+ $Y2=0
cc_498 N_SCD_c_561_n N_A_307_74#_c_2159_n 0.00511032f $X=2.925 $Y=1.62 $X2=0
+ $Y2=0
cc_499 N_SCD_M1041_g N_A_307_74#_c_2161_n 0.00174384f $X=2.435 $Y=2.64 $X2=0
+ $Y2=0
cc_500 N_SCD_M1015_g N_A_307_74#_c_2177_n 0.00177354f $X=2.79 $Y=0.58 $X2=0
+ $Y2=0
cc_501 N_SCD_M1041_g N_A_307_74#_c_2195_n 0.00630972f $X=2.435 $Y=2.64 $X2=0
+ $Y2=0
cc_502 N_SCD_M1015_g N_VGND_c_2407_n 0.0117409f $X=2.79 $Y=0.58 $X2=0 $Y2=0
cc_503 SCD N_VGND_c_2407_n 0.026063f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_504 N_SCD_c_563_n N_VGND_c_2407_n 0.0070747f $X=2.97 $Y=1.115 $X2=0 $Y2=0
cc_505 N_SCD_M1015_g N_VGND_c_2418_n 0.00383152f $X=2.79 $Y=0.58 $X2=0 $Y2=0
cc_506 N_SCD_M1015_g N_VGND_c_2439_n 0.0075725f $X=2.79 $Y=0.58 $X2=0 $Y2=0
cc_507 N_CLK_c_610_n N_A_619_368#_M1035_g 0.0188406f $X=3.78 $Y=1.22 $X2=0 $Y2=0
cc_508 CLK N_A_619_368#_M1035_g 0.0070177f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_509 N_CLK_c_612_n N_A_619_368#_M1035_g 0.0207024f $X=3.83 $Y=1.385 $X2=0
+ $Y2=0
cc_510 N_CLK_M1036_g N_A_619_368#_c_1319_n 0.0187125f $X=3.465 $Y=2.4 $X2=0
+ $Y2=0
cc_511 N_CLK_c_610_n N_A_619_368#_c_1323_n 6.69491e-19 $X=3.78 $Y=1.22 $X2=0
+ $Y2=0
cc_512 N_CLK_M1036_g N_A_619_368#_c_1324_n 0.0114872f $X=3.465 $Y=2.4 $X2=0
+ $Y2=0
cc_513 N_CLK_c_610_n N_A_619_368#_c_1324_n 0.00417982f $X=3.78 $Y=1.22 $X2=0
+ $Y2=0
cc_514 CLK N_A_619_368#_c_1324_n 0.0273382f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_515 N_CLK_c_612_n N_A_619_368#_c_1324_n 0.0152232f $X=3.83 $Y=1.385 $X2=0
+ $Y2=0
cc_516 N_CLK_M1036_g N_A_619_368#_c_1350_n 0.00408099f $X=3.465 $Y=2.4 $X2=0
+ $Y2=0
cc_517 CLK N_A_619_368#_c_1350_n 0.0289811f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_518 N_CLK_c_612_n N_A_619_368#_c_1350_n 0.0121116f $X=3.83 $Y=1.385 $X2=0
+ $Y2=0
cc_519 CLK N_A_619_368#_c_1325_n 0.0147056f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_520 N_CLK_M1036_g N_A_619_368#_c_1353_n 0.0125809f $X=3.465 $Y=2.4 $X2=0
+ $Y2=0
cc_521 N_CLK_c_612_n N_A_619_368#_c_1327_n 0.00440274f $X=3.83 $Y=1.385 $X2=0
+ $Y2=0
cc_522 N_CLK_M1036_g N_VPWR_c_1958_n 0.0114478f $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_523 N_CLK_M1036_g N_VPWR_c_1984_n 0.00460063f $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_524 N_CLK_M1036_g N_VPWR_c_1985_n 0.0245701f $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_525 N_CLK_M1036_g N_VPWR_c_1956_n 0.00466809f $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_526 N_CLK_M1036_g N_A_307_74#_c_2159_n 0.0156099f $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_527 N_CLK_M1036_g N_A_307_74#_c_2197_n 0.0046836f $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_528 N_CLK_c_610_n N_VGND_c_2407_n 0.00224794f $X=3.78 $Y=1.22 $X2=0 $Y2=0
cc_529 N_CLK_c_610_n N_VGND_c_2408_n 0.0118636f $X=3.78 $Y=1.22 $X2=0 $Y2=0
cc_530 CLK N_VGND_c_2408_n 0.0254134f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_531 N_CLK_c_612_n N_VGND_c_2408_n 8.35753e-19 $X=3.83 $Y=1.385 $X2=0 $Y2=0
cc_532 N_CLK_c_610_n N_VGND_c_2429_n 0.00383152f $X=3.78 $Y=1.22 $X2=0 $Y2=0
cc_533 N_CLK_c_610_n N_VGND_c_2439_n 0.00762539f $X=3.78 $Y=1.22 $X2=0 $Y2=0
cc_534 N_A_871_74#_c_660_n N_A_1252_376#_M1030_g 0.0082472f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_535 N_A_871_74#_c_678_n N_A_1252_376#_M1030_g 0.00256901f $X=6.155 $Y=2.905
+ $X2=0 $Y2=0
cc_536 N_A_871_74#_c_679_n N_A_1252_376#_M1030_g 0.0148939f $X=7.155 $Y=2.25
+ $X2=0 $Y2=0
cc_537 N_A_871_74#_c_687_n N_A_1252_376#_M1030_g 0.00434701f $X=6.187 $Y=2.25
+ $X2=0 $Y2=0
cc_538 N_A_871_74#_c_679_n N_A_1252_376#_c_911_n 0.0134562f $X=7.155 $Y=2.25
+ $X2=0 $Y2=0
cc_539 N_A_871_74#_c_671_n N_A_1252_376#_c_912_n 7.74578e-19 $X=5.395 $Y=1.96
+ $X2=0 $Y2=0
cc_540 N_A_871_74#_c_660_n N_A_1252_376#_c_912_n 0.00740993f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_541 N_A_871_74#_c_661_n N_A_1252_376#_c_912_n 0.00704054f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_542 N_A_871_74#_M1026_g N_A_1252_376#_c_904_n 0.0214745f $X=6.295 $Y=0.615
+ $X2=0 $Y2=0
cc_543 N_A_871_74#_c_660_n N_A_1252_376#_c_913_n 0.0123703f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_544 N_A_871_74#_c_679_n N_A_1252_376#_c_913_n 0.053889f $X=7.155 $Y=2.25
+ $X2=0 $Y2=0
cc_545 N_A_871_74#_c_660_n N_A_1252_376#_c_914_n 0.00209505f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_546 N_A_871_74#_c_681_n N_A_1252_376#_c_915_n 0.0226769f $X=7.995 $Y=2.99
+ $X2=0 $Y2=0
cc_547 N_A_871_74#_c_683_n N_A_1252_376#_c_915_n 0.0325867f $X=8.08 $Y=2.905
+ $X2=0 $Y2=0
cc_548 N_A_871_74#_c_679_n N_A_1252_376#_c_916_n 0.0128468f $X=7.155 $Y=2.25
+ $X2=0 $Y2=0
cc_549 N_A_871_74#_c_683_n N_A_1252_376#_c_916_n 0.00323174f $X=8.08 $Y=2.905
+ $X2=0 $Y2=0
cc_550 N_A_871_74#_c_685_n N_A_1252_376#_c_916_n 0.00813475f $X=8.165 $Y=2.135
+ $X2=0 $Y2=0
cc_551 N_A_871_74#_c_660_n N_A_1252_376#_c_908_n 0.00205641f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_552 N_A_871_74#_c_661_n N_A_1252_376#_c_909_n 0.0337032f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_553 N_A_871_74#_c_656_n N_A_1069_81#_M1019_d 4.5412e-19 $X=5.39 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_554 N_A_871_74#_c_666_n N_A_1069_81#_M1019_d 0.00650998f $X=5.395 $Y=1.29
+ $X2=-0.19 $Y2=-0.245
cc_555 N_A_871_74#_c_679_n N_A_1069_81#_M1042_g 0.00415215f $X=7.155 $Y=2.25
+ $X2=0 $Y2=0
cc_556 N_A_871_74#_c_680_n N_A_1069_81#_M1042_g 0.0122168f $X=7.24 $Y=2.905
+ $X2=0 $Y2=0
cc_557 N_A_871_74#_c_681_n N_A_1069_81#_M1042_g 0.00396457f $X=7.995 $Y=2.99
+ $X2=0 $Y2=0
cc_558 N_A_871_74#_c_683_n N_A_1069_81#_M1042_g 6.46673e-19 $X=8.08 $Y=2.905
+ $X2=0 $Y2=0
cc_559 N_A_871_74#_c_667_n N_A_1069_81#_M1003_g 0.00918793f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_560 N_A_871_74#_c_667_n N_A_1069_81#_c_994_n 0.00550305f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_561 N_A_871_74#_c_667_n N_A_1069_81#_M1048_g 0.00827881f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_562 N_A_871_74#_M1032_g N_A_1069_81#_M1011_g 0.0112306f $X=10.26 $Y=0.69
+ $X2=0 $Y2=0
cc_563 N_A_871_74#_c_664_n N_A_1069_81#_M1011_g 6.92746e-19 $X=10.545 $Y=1.365
+ $X2=0 $Y2=0
cc_564 N_A_871_74#_c_667_n N_A_1069_81#_c_997_n 0.00404676f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_565 N_A_871_74#_c_652_n N_A_1069_81#_c_999_n 0.0180937f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_566 N_A_871_74#_c_667_n N_A_1069_81#_c_999_n 0.00373591f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_567 N_A_871_74#_c_646_n N_A_1069_81#_c_1029_n 0.00361747f $X=6.02 $Y=1.365
+ $X2=0 $Y2=0
cc_568 N_A_871_74#_M1026_g N_A_1069_81#_c_1029_n 0.021861f $X=6.295 $Y=0.615
+ $X2=0 $Y2=0
cc_569 N_A_871_74#_c_660_n N_A_1069_81#_c_1029_n 0.0166876f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_570 N_A_871_74#_c_661_n N_A_1069_81#_c_1029_n 0.00318891f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_571 N_A_871_74#_c_666_n N_A_1069_81#_c_1033_n 0.0268483f $X=5.395 $Y=1.29
+ $X2=0 $Y2=0
cc_572 N_A_871_74#_M1026_g N_A_1069_81#_c_1000_n 0.00554569f $X=6.295 $Y=0.615
+ $X2=0 $Y2=0
cc_573 N_A_871_74#_c_660_n N_A_1069_81#_c_1000_n 0.0310926f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_574 N_A_871_74#_c_660_n N_A_1069_81#_c_1002_n 0.0140103f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_575 N_A_871_74#_c_661_n N_A_1069_81#_c_1002_n 0.00181486f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_576 N_A_871_74#_c_679_n N_A_1069_81#_c_1002_n 0.00555233f $X=7.155 $Y=2.25
+ $X2=0 $Y2=0
cc_577 N_A_871_74#_c_663_n N_A_1069_81#_c_1004_n 0.00180199f $X=8.565 $Y=1.43
+ $X2=0 $Y2=0
cc_578 N_A_871_74#_c_663_n N_A_1069_81#_c_1005_n 0.0140773f $X=8.565 $Y=1.43
+ $X2=0 $Y2=0
cc_579 N_A_871_74#_c_667_n N_A_1069_81#_c_1005_n 0.0208175f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_580 N_A_871_74#_c_663_n N_A_1069_81#_c_1006_n 8.79449e-19 $X=8.565 $Y=1.43
+ $X2=0 $Y2=0
cc_581 N_A_871_74#_c_667_n N_A_1069_81#_c_1006_n 0.0141435f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_582 N_A_871_74#_M1006_g N_A_1069_81#_c_1013_n 3.32654e-19 $X=5.43 $Y=2.525
+ $X2=0 $Y2=0
cc_583 N_A_871_74#_c_673_n N_A_1069_81#_c_1013_n 0.0232943f $X=6.07 $Y=2.99
+ $X2=0 $Y2=0
cc_584 N_A_871_74#_c_658_n N_A_1069_81#_c_1013_n 9.31843e-19 $X=5.395 $Y=1.455
+ $X2=0 $Y2=0
cc_585 N_A_871_74#_M1006_g N_A_1069_81#_c_1007_n 0.00645636f $X=5.43 $Y=2.525
+ $X2=0 $Y2=0
cc_586 N_A_871_74#_c_646_n N_A_1069_81#_c_1007_n 0.0145736f $X=6.02 $Y=1.365
+ $X2=0 $Y2=0
cc_587 N_A_871_74#_M1026_g N_A_1069_81#_c_1007_n 0.00324964f $X=6.295 $Y=0.615
+ $X2=0 $Y2=0
cc_588 N_A_871_74#_c_659_n N_A_1069_81#_c_1007_n 0.00788192f $X=5.395 $Y=1.455
+ $X2=0 $Y2=0
cc_589 N_A_871_74#_c_660_n N_A_1069_81#_c_1007_n 0.0890046f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_590 N_A_871_74#_c_661_n N_A_1069_81#_c_1007_n 0.00856636f $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_591 N_A_871_74#_c_666_n N_A_1069_81#_c_1007_n 0.0864367f $X=5.395 $Y=1.29
+ $X2=0 $Y2=0
cc_592 N_A_871_74#_c_687_n N_A_1069_81#_c_1007_n 0.0129429f $X=6.187 $Y=2.25
+ $X2=0 $Y2=0
cc_593 N_A_871_74#_c_681_n N_SET_B_M1034_g 0.00245855f $X=7.995 $Y=2.99 $X2=0
+ $Y2=0
cc_594 N_A_871_74#_c_683_n N_SET_B_M1034_g 0.0194795f $X=8.08 $Y=2.905 $X2=0
+ $Y2=0
cc_595 N_A_871_74#_c_685_n N_SET_B_M1034_g 0.00746389f $X=8.165 $Y=2.135 $X2=0
+ $Y2=0
cc_596 N_A_871_74#_c_662_n N_SET_B_M1034_g 0.00340414f $X=8.48 $Y=2.05 $X2=0
+ $Y2=0
cc_597 N_A_871_74#_c_662_n N_SET_B_M1014_g 0.00120161f $X=8.48 $Y=2.05 $X2=0
+ $Y2=0
cc_598 N_A_871_74#_c_663_n N_SET_B_M1014_g 0.00634353f $X=8.565 $Y=1.43 $X2=0
+ $Y2=0
cc_599 N_A_871_74#_c_651_n N_SET_B_c_1172_n 0.00307898f $X=11.18 $Y=1.41 $X2=0
+ $Y2=0
cc_600 N_A_871_74#_c_652_n N_SET_B_c_1172_n 0.00454536f $X=10.835 $Y=1.41 $X2=0
+ $Y2=0
cc_601 N_A_871_74#_c_653_n N_SET_B_c_1172_n 0.0108908f $X=11.67 $Y=1.545 $X2=0
+ $Y2=0
cc_602 N_A_871_74#_M1010_g N_SET_B_c_1172_n 0.00129463f $X=11.76 $Y=2.485 $X2=0
+ $Y2=0
cc_603 N_A_871_74#_c_684_n N_SET_B_c_1172_n 0.00699781f $X=8.395 $Y=2.135 $X2=0
+ $Y2=0
cc_604 N_A_871_74#_c_685_n N_SET_B_c_1172_n 6.08327e-19 $X=8.165 $Y=2.135 $X2=0
+ $Y2=0
cc_605 N_A_871_74#_c_662_n N_SET_B_c_1172_n 0.0184668f $X=8.48 $Y=2.05 $X2=0
+ $Y2=0
cc_606 N_A_871_74#_c_664_n N_SET_B_c_1172_n 0.024823f $X=10.545 $Y=1.365 $X2=0
+ $Y2=0
cc_607 N_A_871_74#_c_667_n N_SET_B_c_1172_n 0.0532159f $X=10.38 $Y=1.365 $X2=0
+ $Y2=0
cc_608 N_A_871_74#_c_668_n N_SET_B_c_1172_n 0.00257296f $X=11.39 $Y=1.41 $X2=0
+ $Y2=0
cc_609 N_A_871_74#_c_685_n N_SET_B_c_1173_n 4.33107e-19 $X=8.165 $Y=2.135 $X2=0
+ $Y2=0
cc_610 N_A_871_74#_c_662_n N_SET_B_c_1173_n 4.56685e-19 $X=8.48 $Y=2.05 $X2=0
+ $Y2=0
cc_611 N_A_871_74#_c_684_n N_SET_B_c_1174_n 0.00418019f $X=8.395 $Y=2.135 $X2=0
+ $Y2=0
cc_612 N_A_871_74#_c_685_n N_SET_B_c_1174_n 0.0129383f $X=8.165 $Y=2.135 $X2=0
+ $Y2=0
cc_613 N_A_871_74#_c_662_n N_SET_B_c_1174_n 0.0235365f $X=8.48 $Y=2.05 $X2=0
+ $Y2=0
cc_614 N_A_871_74#_c_684_n N_SET_B_c_1178_n 0.00157943f $X=8.395 $Y=2.135 $X2=0
+ $Y2=0
cc_615 N_A_871_74#_c_685_n N_SET_B_c_1178_n 0.00245159f $X=8.165 $Y=2.135 $X2=0
+ $Y2=0
cc_616 N_A_871_74#_c_662_n N_SET_B_c_1178_n 0.00142596f $X=8.48 $Y=2.05 $X2=0
+ $Y2=0
cc_617 N_A_871_74#_c_655_n N_A_619_368#_M1035_g 0.00716152f $X=4.495 $Y=0.505
+ $X2=0 $Y2=0
cc_618 N_A_871_74#_c_657_n N_A_619_368#_M1035_g 0.00462516f $X=4.66 $Y=0.34
+ $X2=0 $Y2=0
cc_619 N_A_871_74#_c_674_n N_A_619_368#_M1046_g 0.00149128f $X=4.72 $Y=2.99
+ $X2=0 $Y2=0
cc_620 N_A_871_74#_c_647_n N_A_619_368#_c_1312_n 0.00865427f $X=5.56 $Y=1.365
+ $X2=0 $Y2=0
cc_621 N_A_871_74#_c_658_n N_A_619_368#_c_1312_n 3.40049e-19 $X=5.395 $Y=1.455
+ $X2=0 $Y2=0
cc_622 N_A_871_74#_c_666_n N_A_619_368#_c_1312_n 7.18595e-19 $X=5.395 $Y=1.29
+ $X2=0 $Y2=0
cc_623 N_A_871_74#_M1006_g N_A_619_368#_c_1330_n 0.0192695f $X=5.43 $Y=2.525
+ $X2=0 $Y2=0
cc_624 N_A_871_74#_c_671_n N_A_619_368#_c_1330_n 0.00865427f $X=5.395 $Y=1.96
+ $X2=0 $Y2=0
cc_625 N_A_871_74#_c_672_n N_A_619_368#_c_1330_n 0.00716202f $X=4.555 $Y=2.725
+ $X2=0 $Y2=0
cc_626 N_A_871_74#_c_673_n N_A_619_368#_c_1330_n 0.0115238f $X=6.07 $Y=2.99
+ $X2=0 $Y2=0
cc_627 N_A_871_74#_c_647_n N_A_619_368#_c_1313_n 0.00655065f $X=5.56 $Y=1.365
+ $X2=0 $Y2=0
cc_628 N_A_871_74#_c_658_n N_A_619_368#_c_1313_n 8.57179e-19 $X=5.395 $Y=1.455
+ $X2=0 $Y2=0
cc_629 N_A_871_74#_c_661_n N_A_619_368#_c_1313_n 8.21735e-19 $X=6.185 $Y=1.135
+ $X2=0 $Y2=0
cc_630 N_A_871_74#_c_655_n N_A_619_368#_c_1314_n 0.00120198f $X=4.495 $Y=0.505
+ $X2=0 $Y2=0
cc_631 N_A_871_74#_c_656_n N_A_619_368#_c_1314_n 0.00410477f $X=5.39 $Y=0.34
+ $X2=0 $Y2=0
cc_632 N_A_871_74#_M1006_g N_A_619_368#_c_1331_n 0.0105864f $X=5.43 $Y=2.525
+ $X2=0 $Y2=0
cc_633 N_A_871_74#_c_673_n N_A_619_368#_c_1331_n 0.0142547f $X=6.07 $Y=2.99
+ $X2=0 $Y2=0
cc_634 N_A_871_74#_c_655_n N_A_619_368#_c_1315_n 0.00417367f $X=4.495 $Y=0.505
+ $X2=0 $Y2=0
cc_635 N_A_871_74#_c_656_n N_A_619_368#_c_1315_n 0.0163078f $X=5.39 $Y=0.34
+ $X2=0 $Y2=0
cc_636 N_A_871_74#_c_666_n N_A_619_368#_c_1315_n 0.013812f $X=5.395 $Y=1.29
+ $X2=0 $Y2=0
cc_637 N_A_871_74#_M1006_g N_A_619_368#_M1002_g 0.0109264f $X=5.43 $Y=2.525
+ $X2=0 $Y2=0
cc_638 N_A_871_74#_c_673_n N_A_619_368#_M1002_g 0.017774f $X=6.07 $Y=2.99 $X2=0
+ $Y2=0
cc_639 N_A_871_74#_c_678_n N_A_619_368#_M1002_g 0.00617239f $X=6.155 $Y=2.905
+ $X2=0 $Y2=0
cc_640 N_A_871_74#_c_687_n N_A_619_368#_M1002_g 0.00108428f $X=6.187 $Y=2.25
+ $X2=0 $Y2=0
cc_641 N_A_871_74#_c_673_n N_A_619_368#_c_1334_n 0.00458792f $X=6.07 $Y=2.99
+ $X2=0 $Y2=0
cc_642 N_A_871_74#_c_681_n N_A_619_368#_c_1334_n 0.0139183f $X=7.995 $Y=2.99
+ $X2=0 $Y2=0
cc_643 N_A_871_74#_c_682_n N_A_619_368#_c_1334_n 0.00420304f $X=7.325 $Y=2.99
+ $X2=0 $Y2=0
cc_644 N_A_871_74#_c_683_n N_A_619_368#_c_1335_n 0.0031126f $X=8.08 $Y=2.905
+ $X2=0 $Y2=0
cc_645 N_A_871_74#_c_684_n N_A_619_368#_c_1335_n 0.00356641f $X=8.395 $Y=2.135
+ $X2=0 $Y2=0
cc_646 N_A_871_74#_c_652_n N_A_619_368#_c_1337_n 0.0148136f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_647 N_A_871_74#_c_652_n N_A_619_368#_c_1338_n 0.00314865f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_648 N_A_871_74#_M1010_g N_A_619_368#_c_1340_n 0.0248224f $X=11.76 $Y=2.485
+ $X2=0 $Y2=0
cc_649 N_A_871_74#_c_668_n N_A_619_368#_c_1340_n 0.0148136f $X=11.39 $Y=1.41
+ $X2=0 $Y2=0
cc_650 N_A_871_74#_M1010_g N_A_619_368#_c_1342_n 0.0088468f $X=11.76 $Y=2.485
+ $X2=0 $Y2=0
cc_651 N_A_871_74#_c_653_n N_A_619_368#_c_1317_n 0.0379689f $X=11.67 $Y=1.545
+ $X2=0 $Y2=0
cc_652 N_A_871_74#_c_655_n N_A_619_368#_c_1320_n 0.00154941f $X=4.495 $Y=0.505
+ $X2=0 $Y2=0
cc_653 N_A_871_74#_c_658_n N_A_619_368#_c_1321_n 3.40049e-19 $X=5.395 $Y=1.455
+ $X2=0 $Y2=0
cc_654 N_A_871_74#_c_659_n N_A_619_368#_c_1321_n 0.00865427f $X=5.395 $Y=1.455
+ $X2=0 $Y2=0
cc_655 N_A_871_74#_c_651_n N_A_619_368#_c_1349_n 0.0148136f $X=11.18 $Y=1.41
+ $X2=0 $Y2=0
cc_656 N_A_871_74#_c_653_n N_A_619_368#_c_1322_n 0.00719229f $X=11.67 $Y=1.545
+ $X2=0 $Y2=0
cc_657 N_A_871_74#_c_668_n N_A_619_368#_c_1322_n 0.00115082f $X=11.39 $Y=1.41
+ $X2=0 $Y2=0
cc_658 N_A_871_74#_M1046_d N_A_619_368#_c_1350_n 0.00354757f $X=4.385 $Y=1.84
+ $X2=0 $Y2=0
cc_659 N_A_871_74#_c_655_n N_A_619_368#_c_1325_n 0.0130668f $X=4.495 $Y=0.505
+ $X2=0 $Y2=0
cc_660 N_A_871_74#_c_652_n N_A_619_368#_c_1352_n 0.015083f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_661 N_A_871_74#_M1010_g N_A_619_368#_c_1352_n 0.0122f $X=11.76 $Y=2.485 $X2=0
+ $Y2=0
cc_662 N_A_871_74#_c_664_n N_A_619_368#_c_1352_n 0.0651024f $X=10.545 $Y=1.365
+ $X2=0 $Y2=0
cc_663 N_A_871_74#_c_667_n N_A_619_368#_c_1352_n 0.0757222f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_664 N_A_871_74#_c_653_n N_A_619_368#_c_1326_n 0.00963508f $X=11.67 $Y=1.545
+ $X2=0 $Y2=0
cc_665 N_A_871_74#_M1010_g N_A_619_368#_c_1326_n 0.00312843f $X=11.76 $Y=2.485
+ $X2=0 $Y2=0
cc_666 N_A_871_74#_c_665_n N_A_619_368#_c_1326_n 0.0163715f $X=11.225 $Y=1.365
+ $X2=0 $Y2=0
cc_667 N_A_871_74#_c_668_n N_A_619_368#_c_1326_n 0.0016069f $X=11.39 $Y=1.41
+ $X2=0 $Y2=0
cc_668 N_A_871_74#_c_662_n N_A_619_368#_c_1328_n 0.00575281f $X=8.48 $Y=2.05
+ $X2=0 $Y2=0
cc_669 N_A_871_74#_c_667_n N_A_619_368#_c_1328_n 0.00273126f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_670 N_A_871_74#_c_662_n N_A_619_368#_c_1355_n 0.020865f $X=8.48 $Y=2.05 $X2=0
+ $Y2=0
cc_671 N_A_871_74#_c_667_n N_A_619_368#_c_1355_n 0.0204754f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_672 N_A_871_74#_M1010_g N_A_2067_74#_c_1695_n 0.0112991f $X=11.76 $Y=2.485
+ $X2=0 $Y2=0
cc_673 N_A_871_74#_M1039_g N_A_2067_74#_c_1683_n 0.0108721f $X=10.76 $Y=0.69
+ $X2=0 $Y2=0
cc_674 N_A_871_74#_c_651_n N_A_2067_74#_c_1683_n 0.0127999f $X=11.18 $Y=1.41
+ $X2=0 $Y2=0
cc_675 N_A_871_74#_c_665_n N_A_2067_74#_c_1683_n 0.0484336f $X=11.225 $Y=1.365
+ $X2=0 $Y2=0
cc_676 N_A_871_74#_M1039_g N_A_2067_74#_c_1684_n 0.00325302f $X=10.76 $Y=0.69
+ $X2=0 $Y2=0
cc_677 N_A_871_74#_c_653_n N_A_2067_74#_c_1684_n 0.00296879f $X=11.67 $Y=1.545
+ $X2=0 $Y2=0
cc_678 N_A_871_74#_c_665_n N_A_2067_74#_c_1684_n 7.314e-19 $X=11.225 $Y=1.365
+ $X2=0 $Y2=0
cc_679 N_A_871_74#_c_668_n N_A_2067_74#_c_1684_n 2.19145e-19 $X=11.39 $Y=1.41
+ $X2=0 $Y2=0
cc_680 N_A_871_74#_M1010_g N_A_2067_74#_c_1696_n 0.00622574f $X=11.76 $Y=2.485
+ $X2=0 $Y2=0
cc_681 N_A_871_74#_M1032_g N_A_2067_74#_c_1687_n 0.00233014f $X=10.26 $Y=0.69
+ $X2=0 $Y2=0
cc_682 N_A_871_74#_M1039_g N_A_2067_74#_c_1687_n 0.00694931f $X=10.76 $Y=0.69
+ $X2=0 $Y2=0
cc_683 N_A_871_74#_c_652_n N_A_2067_74#_c_1687_n 0.00409869f $X=10.835 $Y=1.41
+ $X2=0 $Y2=0
cc_684 N_A_871_74#_c_664_n N_A_2067_74#_c_1687_n 0.0257498f $X=10.545 $Y=1.365
+ $X2=0 $Y2=0
cc_685 N_A_871_74#_M1010_g N_A_2067_74#_c_1701_n 0.00710453f $X=11.76 $Y=2.485
+ $X2=0 $Y2=0
cc_686 N_A_871_74#_c_653_n N_A_2067_74#_c_1688_n 4.20992e-19 $X=11.67 $Y=1.545
+ $X2=0 $Y2=0
cc_687 N_A_871_74#_M1010_g N_A_2067_74#_c_1688_n 0.00100497f $X=11.76 $Y=2.485
+ $X2=0 $Y2=0
cc_688 N_A_871_74#_c_679_n N_VPWR_M1030_d 0.0123722f $X=7.155 $Y=2.25 $X2=0
+ $Y2=0
cc_689 N_A_871_74#_c_680_n N_VPWR_M1030_d 0.0118144f $X=7.24 $Y=2.905 $X2=0
+ $Y2=0
cc_690 N_A_871_74#_c_683_n N_VPWR_M1034_d 0.00453281f $X=8.08 $Y=2.905 $X2=0
+ $Y2=0
cc_691 N_A_871_74#_c_673_n N_VPWR_c_1959_n 0.0156599f $X=6.07 $Y=2.99 $X2=0
+ $Y2=0
cc_692 N_A_871_74#_c_678_n N_VPWR_c_1959_n 0.0228376f $X=6.155 $Y=2.905 $X2=0
+ $Y2=0
cc_693 N_A_871_74#_c_679_n N_VPWR_c_1959_n 0.0418307f $X=7.155 $Y=2.25 $X2=0
+ $Y2=0
cc_694 N_A_871_74#_c_680_n N_VPWR_c_1959_n 0.0324324f $X=7.24 $Y=2.905 $X2=0
+ $Y2=0
cc_695 N_A_871_74#_c_682_n N_VPWR_c_1959_n 0.0156604f $X=7.325 $Y=2.99 $X2=0
+ $Y2=0
cc_696 N_A_871_74#_c_681_n N_VPWR_c_1960_n 0.0546768f $X=7.995 $Y=2.99 $X2=0
+ $Y2=0
cc_697 N_A_871_74#_c_682_n N_VPWR_c_1960_n 0.0115893f $X=7.325 $Y=2.99 $X2=0
+ $Y2=0
cc_698 N_A_871_74#_c_681_n N_VPWR_c_1961_n 0.0150384f $X=7.995 $Y=2.99 $X2=0
+ $Y2=0
cc_699 N_A_871_74#_c_683_n N_VPWR_c_1961_n 0.0398049f $X=8.08 $Y=2.905 $X2=0
+ $Y2=0
cc_700 N_A_871_74#_c_684_n N_VPWR_c_1961_n 0.0203752f $X=8.395 $Y=2.135 $X2=0
+ $Y2=0
cc_701 N_A_871_74#_c_673_n N_VPWR_c_1979_n 0.0975191f $X=6.07 $Y=2.99 $X2=0
+ $Y2=0
cc_702 N_A_871_74#_c_674_n N_VPWR_c_1979_n 0.0234498f $X=4.72 $Y=2.99 $X2=0
+ $Y2=0
cc_703 N_A_871_74#_c_674_n N_VPWR_c_1985_n 0.0125561f $X=4.72 $Y=2.99 $X2=0
+ $Y2=0
cc_704 N_A_871_74#_c_673_n N_VPWR_c_1956_n 0.0511446f $X=6.07 $Y=2.99 $X2=0
+ $Y2=0
cc_705 N_A_871_74#_c_674_n N_VPWR_c_1956_n 0.0127907f $X=4.72 $Y=2.99 $X2=0
+ $Y2=0
cc_706 N_A_871_74#_c_681_n N_VPWR_c_1956_n 0.028344f $X=7.995 $Y=2.99 $X2=0
+ $Y2=0
cc_707 N_A_871_74#_c_682_n N_VPWR_c_1956_n 0.00583135f $X=7.325 $Y=2.99 $X2=0
+ $Y2=0
cc_708 N_A_871_74#_c_656_n N_A_307_74#_M1019_s 0.00224741f $X=5.39 $Y=0.34 $X2=0
+ $Y2=0
cc_709 N_A_871_74#_M1046_d N_A_307_74#_c_2160_n 0.00548347f $X=4.385 $Y=1.84
+ $X2=0 $Y2=0
cc_710 N_A_871_74#_c_672_n N_A_307_74#_c_2160_n 0.0223808f $X=4.555 $Y=2.725
+ $X2=0 $Y2=0
cc_711 N_A_871_74#_c_673_n N_A_307_74#_c_2160_n 0.00442331f $X=6.07 $Y=2.99
+ $X2=0 $Y2=0
cc_712 N_A_871_74#_c_655_n N_A_307_74#_c_2155_n 0.0273357f $X=4.495 $Y=0.505
+ $X2=0 $Y2=0
cc_713 N_A_871_74#_c_656_n N_A_307_74#_c_2155_n 0.0199805f $X=5.39 $Y=0.34 $X2=0
+ $Y2=0
cc_714 N_A_871_74#_c_666_n N_A_307_74#_c_2155_n 0.0100954f $X=5.395 $Y=1.29
+ $X2=0 $Y2=0
cc_715 N_A_871_74#_M1006_g N_A_307_74#_c_2162_n 0.0116109f $X=5.43 $Y=2.525
+ $X2=0 $Y2=0
cc_716 N_A_871_74#_c_671_n N_A_307_74#_c_2162_n 8.40494e-19 $X=5.395 $Y=1.96
+ $X2=0 $Y2=0
cc_717 N_A_871_74#_c_672_n N_A_307_74#_c_2162_n 0.0215555f $X=4.555 $Y=2.725
+ $X2=0 $Y2=0
cc_718 N_A_871_74#_c_673_n N_A_307_74#_c_2162_n 0.0344759f $X=6.07 $Y=2.99 $X2=0
+ $Y2=0
cc_719 N_A_871_74#_c_658_n N_A_307_74#_c_2162_n 0.012049f $X=5.395 $Y=1.455
+ $X2=0 $Y2=0
cc_720 N_A_871_74#_M1006_g N_A_307_74#_c_2156_n 0.00117754f $X=5.43 $Y=2.525
+ $X2=0 $Y2=0
cc_721 N_A_871_74#_c_647_n N_A_307_74#_c_2156_n 0.00447757f $X=5.56 $Y=1.365
+ $X2=0 $Y2=0
cc_722 N_A_871_74#_c_658_n N_A_307_74#_c_2156_n 0.0502424f $X=5.395 $Y=1.455
+ $X2=0 $Y2=0
cc_723 N_A_871_74#_c_666_n N_A_307_74#_c_2156_n 0.0181764f $X=5.395 $Y=1.29
+ $X2=0 $Y2=0
cc_724 N_A_871_74#_c_678_n A_1204_463# 0.00145959f $X=6.155 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_725 N_A_871_74#_c_684_n N_A_1789_424#_c_2273_n 0.00491328f $X=8.395 $Y=2.135
+ $X2=0 $Y2=0
cc_726 N_A_871_74#_M1010_g N_A_2277_455#_c_2317_n 0.00317116f $X=11.76 $Y=2.485
+ $X2=0 $Y2=0
cc_727 N_A_871_74#_M1010_g N_A_2277_455#_c_2318_n 0.00235121f $X=11.76 $Y=2.485
+ $X2=0 $Y2=0
cc_728 N_A_871_74#_c_657_n N_VGND_c_2408_n 0.011924f $X=4.66 $Y=0.34 $X2=0 $Y2=0
cc_729 N_A_871_74#_M1032_g N_VGND_c_2411_n 3.12362e-19 $X=10.26 $Y=0.69 $X2=0
+ $Y2=0
cc_730 N_A_871_74#_M1032_g N_VGND_c_2422_n 0.00278247f $X=10.26 $Y=0.69 $X2=0
+ $Y2=0
cc_731 N_A_871_74#_M1039_g N_VGND_c_2422_n 0.00278271f $X=10.76 $Y=0.69 $X2=0
+ $Y2=0
cc_732 N_A_871_74#_M1026_g N_VGND_c_2430_n 0.00405757f $X=6.295 $Y=0.615 $X2=0
+ $Y2=0
cc_733 N_A_871_74#_c_656_n N_VGND_c_2430_n 0.0591538f $X=5.39 $Y=0.34 $X2=0
+ $Y2=0
cc_734 N_A_871_74#_c_657_n N_VGND_c_2430_n 0.0235688f $X=4.66 $Y=0.34 $X2=0
+ $Y2=0
cc_735 N_A_871_74#_M1026_g N_VGND_c_2439_n 0.00534666f $X=6.295 $Y=0.615 $X2=0
+ $Y2=0
cc_736 N_A_871_74#_M1032_g N_VGND_c_2439_n 0.00354182f $X=10.26 $Y=0.69 $X2=0
+ $Y2=0
cc_737 N_A_871_74#_M1039_g N_VGND_c_2439_n 0.00358176f $X=10.76 $Y=0.69 $X2=0
+ $Y2=0
cc_738 N_A_871_74#_c_656_n N_VGND_c_2439_n 0.0340476f $X=5.39 $Y=0.34 $X2=0
+ $Y2=0
cc_739 N_A_871_74#_c_657_n N_VGND_c_2439_n 0.0127152f $X=4.66 $Y=0.34 $X2=0
+ $Y2=0
cc_740 N_A_871_74#_M1032_g N_A_1794_74#_c_2594_n 0.00556597f $X=10.26 $Y=0.69
+ $X2=0 $Y2=0
cc_741 N_A_871_74#_M1039_g N_A_1794_74#_c_2594_n 6.97072e-19 $X=10.76 $Y=0.69
+ $X2=0 $Y2=0
cc_742 N_A_871_74#_c_667_n N_A_1794_74#_c_2594_n 0.0650467f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_743 N_A_871_74#_c_667_n N_A_1794_74#_c_2595_n 0.0189433f $X=10.38 $Y=1.365
+ $X2=0 $Y2=0
cc_744 N_A_871_74#_M1032_g N_A_1794_74#_c_2603_n 0.007555f $X=10.26 $Y=0.69
+ $X2=0 $Y2=0
cc_745 N_A_871_74#_M1039_g N_A_1794_74#_c_2603_n 6.40354e-19 $X=10.76 $Y=0.69
+ $X2=0 $Y2=0
cc_746 N_A_871_74#_M1032_g N_A_1794_74#_c_2596_n 0.0104037f $X=10.26 $Y=0.69
+ $X2=0 $Y2=0
cc_747 N_A_871_74#_M1039_g N_A_1794_74#_c_2596_n 0.0112187f $X=10.76 $Y=0.69
+ $X2=0 $Y2=0
cc_748 N_A_871_74#_M1032_g N_A_1794_74#_c_2597_n 0.00155275f $X=10.26 $Y=0.69
+ $X2=0 $Y2=0
cc_749 N_A_871_74#_M1039_g N_A_1794_74#_c_2598_n 0.00165289f $X=10.76 $Y=0.69
+ $X2=0 $Y2=0
cc_750 N_A_1252_376#_c_913_n N_A_1069_81#_M1042_g 0.0199539f $X=7.495 $Y=1.865
+ $X2=0 $Y2=0
cc_751 N_A_1252_376#_c_914_n N_A_1069_81#_M1042_g 0.00815395f $X=6.8 $Y=1.865
+ $X2=0 $Y2=0
cc_752 N_A_1252_376#_c_915_n N_A_1069_81#_M1042_g 0.00601197f $X=7.66 $Y=2.515
+ $X2=0 $Y2=0
cc_753 N_A_1252_376#_c_916_n N_A_1069_81#_M1042_g 0.0104416f $X=7.66 $Y=2.295
+ $X2=0 $Y2=0
cc_754 N_A_1252_376#_c_905_n N_A_1069_81#_M1013_g 0.0056748f $X=7.38 $Y=0.955
+ $X2=0 $Y2=0
cc_755 N_A_1252_376#_c_906_n N_A_1069_81#_M1013_g 0.0116694f $X=7.545 $Y=0.58
+ $X2=0 $Y2=0
cc_756 N_A_1252_376#_c_907_n N_A_1069_81#_M1013_g 8.40065e-19 $X=6.98 $Y=0.955
+ $X2=0 $Y2=0
cc_757 N_A_1252_376#_c_909_n N_A_1069_81#_M1013_g 0.00473478f $X=6.89 $Y=1.1
+ $X2=0 $Y2=0
cc_758 N_A_1252_376#_c_904_n N_A_1069_81#_c_1029_n 0.0113068f $X=6.685 $Y=0.935
+ $X2=0 $Y2=0
cc_759 N_A_1252_376#_c_904_n N_A_1069_81#_c_1000_n 0.00436872f $X=6.685 $Y=0.935
+ $X2=0 $Y2=0
cc_760 N_A_1252_376#_c_907_n N_A_1069_81#_c_1000_n 0.0261072f $X=6.98 $Y=0.955
+ $X2=0 $Y2=0
cc_761 N_A_1252_376#_c_909_n N_A_1069_81#_c_1000_n 0.00911922f $X=6.89 $Y=1.1
+ $X2=0 $Y2=0
cc_762 N_A_1252_376#_c_913_n N_A_1069_81#_c_1001_n 0.0532877f $X=7.495 $Y=1.865
+ $X2=0 $Y2=0
cc_763 N_A_1252_376#_c_914_n N_A_1069_81#_c_1001_n 0.00180482f $X=6.8 $Y=1.865
+ $X2=0 $Y2=0
cc_764 N_A_1252_376#_c_905_n N_A_1069_81#_c_1001_n 0.00950459f $X=7.38 $Y=0.955
+ $X2=0 $Y2=0
cc_765 N_A_1252_376#_c_907_n N_A_1069_81#_c_1001_n 0.0243532f $X=6.98 $Y=0.955
+ $X2=0 $Y2=0
cc_766 N_A_1252_376#_c_908_n N_A_1069_81#_c_1001_n 0.0113822f $X=6.8 $Y=1.7
+ $X2=0 $Y2=0
cc_767 N_A_1252_376#_c_909_n N_A_1069_81#_c_1001_n 0.00787396f $X=6.89 $Y=1.1
+ $X2=0 $Y2=0
cc_768 N_A_1252_376#_c_911_n N_A_1069_81#_c_1002_n 0.00342884f $X=6.635 $Y=1.955
+ $X2=0 $Y2=0
cc_769 N_A_1252_376#_c_913_n N_A_1069_81#_c_1002_n 8.29766e-19 $X=7.495 $Y=1.865
+ $X2=0 $Y2=0
cc_770 N_A_1252_376#_c_905_n N_A_1069_81#_c_1003_n 0.00352223f $X=7.38 $Y=0.955
+ $X2=0 $Y2=0
cc_771 N_A_1252_376#_c_905_n N_A_1069_81#_c_1004_n 0.011024f $X=7.38 $Y=0.955
+ $X2=0 $Y2=0
cc_772 N_A_1252_376#_c_912_n N_A_1069_81#_c_1007_n 0.00123299f $X=6.44 $Y=1.955
+ $X2=0 $Y2=0
cc_773 N_A_1252_376#_c_913_n N_A_1069_81#_c_1008_n 0.0251552f $X=7.495 $Y=1.865
+ $X2=0 $Y2=0
cc_774 N_A_1252_376#_c_905_n N_A_1069_81#_c_1008_n 0.0260001f $X=7.38 $Y=0.955
+ $X2=0 $Y2=0
cc_775 N_A_1252_376#_c_907_n N_A_1069_81#_c_1008_n 9.46074e-19 $X=6.98 $Y=0.955
+ $X2=0 $Y2=0
cc_776 N_A_1252_376#_c_908_n N_A_1069_81#_c_1008_n 8.62215e-19 $X=6.8 $Y=1.7
+ $X2=0 $Y2=0
cc_777 N_A_1252_376#_c_909_n N_A_1069_81#_c_1008_n 3.37949e-19 $X=6.89 $Y=1.1
+ $X2=0 $Y2=0
cc_778 N_A_1252_376#_c_913_n N_A_1069_81#_c_1009_n 0.00102424f $X=7.495 $Y=1.865
+ $X2=0 $Y2=0
cc_779 N_A_1252_376#_c_905_n N_A_1069_81#_c_1009_n 0.00902757f $X=7.38 $Y=0.955
+ $X2=0 $Y2=0
cc_780 N_A_1252_376#_c_907_n N_A_1069_81#_c_1009_n 4.25533e-19 $X=6.98 $Y=0.955
+ $X2=0 $Y2=0
cc_781 N_A_1252_376#_c_908_n N_A_1069_81#_c_1009_n 0.0170764f $X=6.8 $Y=1.7
+ $X2=0 $Y2=0
cc_782 N_A_1252_376#_c_909_n N_A_1069_81#_c_1009_n 0.0072023f $X=6.89 $Y=1.1
+ $X2=0 $Y2=0
cc_783 N_A_1252_376#_c_915_n N_SET_B_M1034_g 0.00376229f $X=7.66 $Y=2.515 $X2=0
+ $Y2=0
cc_784 N_A_1252_376#_c_916_n N_SET_B_M1034_g 0.00293398f $X=7.66 $Y=2.295 $X2=0
+ $Y2=0
cc_785 N_A_1252_376#_c_906_n N_SET_B_M1014_g 0.00187295f $X=7.545 $Y=0.58 $X2=0
+ $Y2=0
cc_786 N_A_1252_376#_c_913_n N_SET_B_c_1173_n 0.00142282f $X=7.495 $Y=1.865
+ $X2=0 $Y2=0
cc_787 N_A_1252_376#_c_915_n N_SET_B_c_1173_n 0.00185005f $X=7.66 $Y=2.515 $X2=0
+ $Y2=0
cc_788 N_A_1252_376#_c_913_n N_SET_B_c_1174_n 0.0122254f $X=7.495 $Y=1.865 $X2=0
+ $Y2=0
cc_789 N_A_1252_376#_c_913_n N_SET_B_c_1178_n 0.00361742f $X=7.495 $Y=1.865
+ $X2=0 $Y2=0
cc_790 N_A_1252_376#_M1030_g N_A_619_368#_M1002_g 0.0310413f $X=6.35 $Y=2.525
+ $X2=0 $Y2=0
cc_791 N_A_1252_376#_M1030_g N_A_619_368#_c_1334_n 0.0123711f $X=6.35 $Y=2.525
+ $X2=0 $Y2=0
cc_792 N_A_1252_376#_M1030_g N_VPWR_c_1959_n 0.0129635f $X=6.35 $Y=2.525 $X2=0
+ $Y2=0
cc_793 N_A_1252_376#_M1030_g N_VPWR_c_1956_n 9.455e-19 $X=6.35 $Y=2.525 $X2=0
+ $Y2=0
cc_794 N_A_1252_376#_c_904_n N_VGND_c_2409_n 0.00545418f $X=6.685 $Y=0.935 $X2=0
+ $Y2=0
cc_795 N_A_1252_376#_c_906_n N_VGND_c_2409_n 0.0236236f $X=7.545 $Y=0.58 $X2=0
+ $Y2=0
cc_796 N_A_1252_376#_c_907_n N_VGND_c_2409_n 0.0287015f $X=6.98 $Y=0.955 $X2=0
+ $Y2=0
cc_797 N_A_1252_376#_c_909_n N_VGND_c_2409_n 0.00217452f $X=6.89 $Y=1.1 $X2=0
+ $Y2=0
cc_798 N_A_1252_376#_c_906_n N_VGND_c_2410_n 0.0104546f $X=7.545 $Y=0.58 $X2=0
+ $Y2=0
cc_799 N_A_1252_376#_c_904_n N_VGND_c_2430_n 0.00518115f $X=6.685 $Y=0.935 $X2=0
+ $Y2=0
cc_800 N_A_1252_376#_c_906_n N_VGND_c_2431_n 0.0145794f $X=7.545 $Y=0.58 $X2=0
+ $Y2=0
cc_801 N_A_1252_376#_c_904_n N_VGND_c_2439_n 0.00534666f $X=6.685 $Y=0.935 $X2=0
+ $Y2=0
cc_802 N_A_1252_376#_c_906_n N_VGND_c_2439_n 0.0120044f $X=7.545 $Y=0.58 $X2=0
+ $Y2=0
cc_803 N_A_1069_81#_M1042_g N_SET_B_M1034_g 0.0158048f $X=7.435 $Y=2.525 $X2=0
+ $Y2=0
cc_804 N_A_1069_81#_M1013_g N_SET_B_M1014_g 0.0537337f $X=7.76 $Y=0.58 $X2=0
+ $Y2=0
cc_805 N_A_1069_81#_c_1004_n N_SET_B_M1014_g 0.00531188f $X=8.05 $Y=1.037 $X2=0
+ $Y2=0
cc_806 N_A_1069_81#_c_1005_n N_SET_B_M1014_g 0.0172588f $X=8.695 $Y=1.065 $X2=0
+ $Y2=0
cc_807 N_A_1069_81#_c_1006_n N_SET_B_M1014_g 0.0140045f $X=8.695 $Y=1.065 $X2=0
+ $Y2=0
cc_808 N_A_1069_81#_c_1008_n N_SET_B_M1014_g 0.00108273f $X=7.51 $Y=1.295 $X2=0
+ $Y2=0
cc_809 N_A_1069_81#_c_1009_n N_SET_B_M1014_g 0.00736022f $X=7.52 $Y=1.375 $X2=0
+ $Y2=0
cc_810 N_A_1069_81#_M1003_g N_SET_B_c_1172_n 0.00307941f $X=9.365 $Y=2.54 $X2=0
+ $Y2=0
cc_811 N_A_1069_81#_M1048_g N_SET_B_c_1172_n 0.0037079f $X=9.815 $Y=2.54 $X2=0
+ $Y2=0
cc_812 N_A_1069_81#_c_1005_n N_SET_B_c_1172_n 0.00863597f $X=8.695 $Y=1.065
+ $X2=0 $Y2=0
cc_813 N_A_1069_81#_c_1003_n N_SET_B_c_1173_n 0.00409741f $X=7.88 $Y=1.295 $X2=0
+ $Y2=0
cc_814 N_A_1069_81#_c_1004_n N_SET_B_c_1173_n 0.00414232f $X=8.05 $Y=1.037 $X2=0
+ $Y2=0
cc_815 N_A_1069_81#_c_1005_n N_SET_B_c_1173_n 3.14556e-19 $X=8.695 $Y=1.065
+ $X2=0 $Y2=0
cc_816 N_A_1069_81#_c_1008_n N_SET_B_c_1173_n 4.88841e-19 $X=7.51 $Y=1.295 $X2=0
+ $Y2=0
cc_817 N_A_1069_81#_c_1009_n N_SET_B_c_1173_n 0.00312846f $X=7.52 $Y=1.375 $X2=0
+ $Y2=0
cc_818 N_A_1069_81#_M1042_g N_SET_B_c_1174_n 3.68151e-19 $X=7.435 $Y=2.525 $X2=0
+ $Y2=0
cc_819 N_A_1069_81#_c_1003_n N_SET_B_c_1174_n 0.0029943f $X=7.88 $Y=1.295 $X2=0
+ $Y2=0
cc_820 N_A_1069_81#_c_1004_n N_SET_B_c_1174_n 0.0116033f $X=8.05 $Y=1.037 $X2=0
+ $Y2=0
cc_821 N_A_1069_81#_c_1005_n N_SET_B_c_1174_n 0.00565821f $X=8.695 $Y=1.065
+ $X2=0 $Y2=0
cc_822 N_A_1069_81#_c_1008_n N_SET_B_c_1174_n 9.69441e-19 $X=7.51 $Y=1.295 $X2=0
+ $Y2=0
cc_823 N_A_1069_81#_c_1009_n N_SET_B_c_1174_n 0.00262295f $X=7.52 $Y=1.375 $X2=0
+ $Y2=0
cc_824 N_A_1069_81#_c_1004_n N_SET_B_c_1178_n 0.00294508f $X=8.05 $Y=1.037 $X2=0
+ $Y2=0
cc_825 N_A_1069_81#_c_1005_n N_SET_B_c_1178_n 4.50247e-19 $X=8.695 $Y=1.065
+ $X2=0 $Y2=0
cc_826 N_A_1069_81#_c_1009_n N_SET_B_c_1178_n 0.0158048f $X=7.52 $Y=1.375 $X2=0
+ $Y2=0
cc_827 N_A_1069_81#_c_1013_n N_A_619_368#_M1002_g 0.0072187f $X=5.705 $Y=2.515
+ $X2=0 $Y2=0
cc_828 N_A_1069_81#_c_1007_n N_A_619_368#_M1002_g 0.00371987f $X=5.72 $Y=2.295
+ $X2=0 $Y2=0
cc_829 N_A_1069_81#_M1042_g N_A_619_368#_c_1334_n 0.0105864f $X=7.435 $Y=2.525
+ $X2=0 $Y2=0
cc_830 N_A_1069_81#_M1003_g N_A_619_368#_c_1335_n 0.01921f $X=9.365 $Y=2.54
+ $X2=0 $Y2=0
cc_831 N_A_1069_81#_M1048_g N_A_619_368#_c_1338_n 0.025519f $X=9.815 $Y=2.54
+ $X2=0 $Y2=0
cc_832 N_A_1069_81#_M1003_g N_A_619_368#_c_1352_n 0.0108793f $X=9.365 $Y=2.54
+ $X2=0 $Y2=0
cc_833 N_A_1069_81#_c_994_n N_A_619_368#_c_1352_n 4.15884e-19 $X=9.725 $Y=1.31
+ $X2=0 $Y2=0
cc_834 N_A_1069_81#_M1048_g N_A_619_368#_c_1352_n 0.0134026f $X=9.815 $Y=2.54
+ $X2=0 $Y2=0
cc_835 N_A_1069_81#_M1003_g N_A_619_368#_c_1328_n 0.0213157f $X=9.365 $Y=2.54
+ $X2=0 $Y2=0
cc_836 N_A_1069_81#_c_1006_n N_A_619_368#_c_1328_n 0.010169f $X=8.695 $Y=1.065
+ $X2=0 $Y2=0
cc_837 N_A_1069_81#_M1003_g N_A_619_368#_c_1355_n 7.57277e-19 $X=9.365 $Y=2.54
+ $X2=0 $Y2=0
cc_838 N_A_1069_81#_M1048_g N_A_2067_74#_c_1719_n 2.228e-19 $X=9.815 $Y=2.54
+ $X2=0 $Y2=0
cc_839 N_A_1069_81#_M1048_g N_A_2067_74#_c_1720_n 3.22747e-19 $X=9.815 $Y=2.54
+ $X2=0 $Y2=0
cc_840 N_A_1069_81#_M1003_g N_VPWR_c_1962_n 0.0111192f $X=9.365 $Y=2.54 $X2=0
+ $Y2=0
cc_841 N_A_1069_81#_M1048_g N_VPWR_c_1962_n 0.00169232f $X=9.815 $Y=2.54 $X2=0
+ $Y2=0
cc_842 N_A_1069_81#_M1003_g N_VPWR_c_1969_n 0.00460063f $X=9.365 $Y=2.54 $X2=0
+ $Y2=0
cc_843 N_A_1069_81#_M1048_g N_VPWR_c_1971_n 0.00517089f $X=9.815 $Y=2.54 $X2=0
+ $Y2=0
cc_844 N_A_1069_81#_M1003_g N_VPWR_c_1956_n 0.00909806f $X=9.365 $Y=2.54 $X2=0
+ $Y2=0
cc_845 N_A_1069_81#_M1048_g N_VPWR_c_1956_n 0.00977588f $X=9.815 $Y=2.54 $X2=0
+ $Y2=0
cc_846 N_A_1069_81#_c_1013_n N_A_307_74#_c_2162_n 0.0182846f $X=5.705 $Y=2.515
+ $X2=0 $Y2=0
cc_847 N_A_1069_81#_c_1007_n N_A_307_74#_c_2162_n 0.00725666f $X=5.72 $Y=2.295
+ $X2=0 $Y2=0
cc_848 N_A_1069_81#_c_1007_n N_A_307_74#_c_2156_n 0.00342338f $X=5.72 $Y=2.295
+ $X2=0 $Y2=0
cc_849 N_A_1069_81#_M1003_g N_A_1789_424#_c_2275_n 0.0147908f $X=9.365 $Y=2.54
+ $X2=0 $Y2=0
cc_850 N_A_1069_81#_M1048_g N_A_1789_424#_c_2275_n 0.0134082f $X=9.815 $Y=2.54
+ $X2=0 $Y2=0
cc_851 N_A_1069_81#_M1048_g N_A_1789_424#_c_2269_n 0.00169334f $X=9.815 $Y=2.54
+ $X2=0 $Y2=0
cc_852 N_A_1069_81#_M1003_g N_A_1789_424#_c_2278_n 6.7008e-19 $X=9.365 $Y=2.54
+ $X2=0 $Y2=0
cc_853 N_A_1069_81#_M1048_g N_A_1789_424#_c_2278_n 0.00992722f $X=9.815 $Y=2.54
+ $X2=0 $Y2=0
cc_854 N_A_1069_81#_M1048_g N_A_1789_424#_c_2271_n 0.00347836f $X=9.815 $Y=2.54
+ $X2=0 $Y2=0
cc_855 N_A_1069_81#_M1003_g N_A_1789_424#_c_2273_n 0.00103604f $X=9.365 $Y=2.54
+ $X2=0 $Y2=0
cc_856 N_A_1069_81#_M1013_g N_VGND_c_2409_n 0.00342558f $X=7.76 $Y=0.58 $X2=0
+ $Y2=0
cc_857 N_A_1069_81#_M1013_g N_VGND_c_2410_n 0.00149517f $X=7.76 $Y=0.58 $X2=0
+ $Y2=0
cc_858 N_A_1069_81#_c_1005_n N_VGND_c_2410_n 0.0209685f $X=8.695 $Y=1.065 $X2=0
+ $Y2=0
cc_859 N_A_1069_81#_M1011_g N_VGND_c_2411_n 0.00973428f $X=9.83 $Y=0.69 $X2=0
+ $Y2=0
cc_860 N_A_1069_81#_c_998_n N_VGND_c_2411_n 0.0115887f $X=9.365 $Y=1.085 $X2=0
+ $Y2=0
cc_861 N_A_1069_81#_c_998_n N_VGND_c_2420_n 0.00444681f $X=9.365 $Y=1.085 $X2=0
+ $Y2=0
cc_862 N_A_1069_81#_M1011_g N_VGND_c_2422_n 0.00383152f $X=9.83 $Y=0.69 $X2=0
+ $Y2=0
cc_863 N_A_1069_81#_c_1029_n N_VGND_c_2430_n 0.0182889f $X=6.475 $Y=0.635 $X2=0
+ $Y2=0
cc_864 N_A_1069_81#_c_1033_n N_VGND_c_2430_n 0.00491805f $X=5.9 $Y=0.635 $X2=0
+ $Y2=0
cc_865 N_A_1069_81#_M1013_g N_VGND_c_2431_n 0.00434272f $X=7.76 $Y=0.58 $X2=0
+ $Y2=0
cc_866 N_A_1069_81#_M1013_g N_VGND_c_2439_n 0.00825979f $X=7.76 $Y=0.58 $X2=0
+ $Y2=0
cc_867 N_A_1069_81#_M1011_g N_VGND_c_2439_n 0.00757637f $X=9.83 $Y=0.69 $X2=0
+ $Y2=0
cc_868 N_A_1069_81#_c_998_n N_VGND_c_2439_n 0.00882517f $X=9.365 $Y=1.085 $X2=0
+ $Y2=0
cc_869 N_A_1069_81#_c_1029_n N_VGND_c_2439_n 0.0246945f $X=6.475 $Y=0.635 $X2=0
+ $Y2=0
cc_870 N_A_1069_81#_c_1033_n N_VGND_c_2439_n 0.00580745f $X=5.9 $Y=0.635 $X2=0
+ $Y2=0
cc_871 N_A_1069_81#_c_1029_n A_1274_81# 0.00374924f $X=6.475 $Y=0.635 $X2=-0.19
+ $Y2=-0.245
cc_872 N_A_1069_81#_c_1000_n A_1274_81# 3.0566e-19 $X=6.56 $Y=1.395 $X2=-0.19
+ $Y2=-0.245
cc_873 N_A_1069_81#_c_998_n N_A_1794_74#_c_2593_n 4.57511e-19 $X=9.365 $Y=1.085
+ $X2=0 $Y2=0
cc_874 N_A_1069_81#_c_1005_n N_A_1794_74#_c_2593_n 0.00836125f $X=8.695 $Y=1.065
+ $X2=0 $Y2=0
cc_875 N_A_1069_81#_c_1006_n N_A_1794_74#_c_2593_n 3.95109e-19 $X=8.695 $Y=1.065
+ $X2=0 $Y2=0
cc_876 N_A_1069_81#_c_994_n N_A_1794_74#_c_2594_n 0.00286179f $X=9.725 $Y=1.31
+ $X2=0 $Y2=0
cc_877 N_A_1069_81#_M1011_g N_A_1794_74#_c_2594_n 0.0142903f $X=9.83 $Y=0.69
+ $X2=0 $Y2=0
cc_878 N_A_1069_81#_c_997_n N_A_1794_74#_c_2594_n 0.00494339f $X=9.365 $Y=1.16
+ $X2=0 $Y2=0
cc_879 N_A_1069_81#_c_998_n N_A_1794_74#_c_2594_n 0.00947016f $X=9.365 $Y=1.085
+ $X2=0 $Y2=0
cc_880 N_A_1069_81#_c_992_n N_A_1794_74#_c_2595_n 0.00940114f $X=9.275 $Y=1.16
+ $X2=0 $Y2=0
cc_881 N_A_1069_81#_c_1005_n N_A_1794_74#_c_2595_n 0.0146575f $X=8.695 $Y=1.065
+ $X2=0 $Y2=0
cc_882 N_A_1069_81#_c_1006_n N_A_1794_74#_c_2595_n 3.57917e-19 $X=8.695 $Y=1.065
+ $X2=0 $Y2=0
cc_883 N_A_1069_81#_M1011_g N_A_1794_74#_c_2597_n 9.48753e-19 $X=9.83 $Y=0.69
+ $X2=0 $Y2=0
cc_884 N_SET_B_M1034_g N_A_619_368#_c_1334_n 0.0110759f $X=7.985 $Y=2.525 $X2=0
+ $Y2=0
cc_885 N_SET_B_c_1172_n N_A_619_368#_c_1316_n 0.00259421f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_886 N_SET_B_c_1172_n N_A_619_368#_c_1317_n 0.00188206f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_887 N_SET_B_c_1172_n N_A_619_368#_c_1322_n 0.00334987f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_888 N_SET_B_c_1172_n N_A_619_368#_c_1352_n 0.0734209f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_889 N_SET_B_c_1172_n N_A_619_368#_c_1326_n 0.0166357f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_890 N_SET_B_M1034_g N_A_619_368#_c_1328_n 0.0107311f $X=7.985 $Y=2.525 $X2=0
+ $Y2=0
cc_891 N_SET_B_c_1172_n N_A_619_368#_c_1328_n 0.00260077f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_892 N_SET_B_c_1178_n N_A_619_368#_c_1328_n 0.00509006f $X=8.06 $Y=1.715 $X2=0
+ $Y2=0
cc_893 N_SET_B_c_1172_n N_A_619_368#_c_1355_n 0.0149981f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_894 N_SET_B_M1018_g N_A_2513_258#_M1016_g 0.0343422f $X=13.25 $Y=2.75 $X2=0
+ $Y2=0
cc_895 N_SET_B_c_1182_n N_A_2513_258#_M1016_g 5.67665e-19 $X=13.27 $Y=1.97 $X2=0
+ $Y2=0
cc_896 N_SET_B_c_1177_n N_A_2513_258#_M1016_g 2.00699e-19 $X=13.27 $Y=1.465
+ $X2=0 $Y2=0
cc_897 N_SET_B_M1021_g N_A_2513_258#_M1020_g 0.057484f $X=13.21 $Y=0.58 $X2=0
+ $Y2=0
cc_898 N_SET_B_c_1171_n N_A_2513_258#_c_1574_n 0.0139984f $X=13.27 $Y=1.805
+ $X2=0 $Y2=0
cc_899 N_SET_B_c_1172_n N_A_2513_258#_c_1574_n 0.0013891f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_900 SET_B N_A_2513_258#_c_1574_n 0.00137814f $X=13.115 $Y=1.58 $X2=0 $Y2=0
cc_901 N_SET_B_c_1182_n N_A_2513_258#_c_1584_n 0.0139984f $X=13.27 $Y=1.97 $X2=0
+ $Y2=0
cc_902 N_SET_B_M1021_g N_A_2513_258#_c_1575_n 0.00109112f $X=13.21 $Y=0.58 $X2=0
+ $Y2=0
cc_903 N_SET_B_c_1172_n N_A_2513_258#_c_1575_n 0.0304377f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_904 SET_B N_A_2513_258#_c_1575_n 0.00262339f $X=13.115 $Y=1.58 $X2=0 $Y2=0
cc_905 N_SET_B_c_1176_n N_A_2513_258#_c_1575_n 8.82895e-19 $X=13.27 $Y=1.465
+ $X2=0 $Y2=0
cc_906 N_SET_B_c_1177_n N_A_2513_258#_c_1575_n 0.0453809f $X=13.27 $Y=1.465
+ $X2=0 $Y2=0
cc_907 N_SET_B_c_1176_n N_A_2513_258#_c_1576_n 0.0139984f $X=13.27 $Y=1.465
+ $X2=0 $Y2=0
cc_908 N_SET_B_c_1177_n N_A_2513_258#_c_1576_n 0.00347086f $X=13.27 $Y=1.465
+ $X2=0 $Y2=0
cc_909 N_SET_B_M1021_g N_A_2513_258#_c_1577_n 0.0144047f $X=13.21 $Y=0.58 $X2=0
+ $Y2=0
cc_910 N_SET_B_c_1172_n N_A_2513_258#_c_1577_n 0.00543614f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_911 SET_B N_A_2513_258#_c_1577_n 0.00220758f $X=13.115 $Y=1.58 $X2=0 $Y2=0
cc_912 N_SET_B_c_1176_n N_A_2513_258#_c_1577_n 0.00469569f $X=13.27 $Y=1.465
+ $X2=0 $Y2=0
cc_913 N_SET_B_c_1177_n N_A_2513_258#_c_1577_n 0.0264703f $X=13.27 $Y=1.465
+ $X2=0 $Y2=0
cc_914 N_SET_B_M1021_g N_A_2513_258#_c_1579_n 9.27178e-19 $X=13.21 $Y=0.58 $X2=0
+ $Y2=0
cc_915 N_SET_B_M1018_g N_A_2513_258#_c_1587_n 9.64169e-19 $X=13.25 $Y=2.75 $X2=0
+ $Y2=0
cc_916 N_SET_B_M1021_g N_A_2067_74#_M1040_g 0.0275785f $X=13.21 $Y=0.58 $X2=0
+ $Y2=0
cc_917 N_SET_B_c_1176_n N_A_2067_74#_c_1679_n 0.0214924f $X=13.27 $Y=1.465 $X2=0
+ $Y2=0
cc_918 N_SET_B_c_1177_n N_A_2067_74#_c_1679_n 0.00245749f $X=13.27 $Y=1.465
+ $X2=0 $Y2=0
cc_919 N_SET_B_c_1172_n N_A_2067_74#_c_1695_n 0.00657317f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_920 N_SET_B_c_1172_n N_A_2067_74#_c_1720_n 0.00145175f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_921 N_SET_B_c_1172_n N_A_2067_74#_c_1684_n 0.00295306f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_922 N_SET_B_M1018_g N_A_2067_74#_c_1697_n 0.0128631f $X=13.25 $Y=2.75 $X2=0
+ $Y2=0
cc_923 N_SET_B_c_1182_n N_A_2067_74#_c_1697_n 0.00143802f $X=13.27 $Y=1.97 $X2=0
+ $Y2=0
cc_924 N_SET_B_c_1172_n N_A_2067_74#_c_1697_n 0.0135949f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_925 SET_B N_A_2067_74#_c_1697_n 0.00238877f $X=13.115 $Y=1.58 $X2=0 $Y2=0
cc_926 N_SET_B_c_1177_n N_A_2067_74#_c_1697_n 0.0261515f $X=13.27 $Y=1.465 $X2=0
+ $Y2=0
cc_927 N_SET_B_M1018_g N_A_2067_74#_c_1698_n 0.0155046f $X=13.25 $Y=2.75 $X2=0
+ $Y2=0
cc_928 N_SET_B_M1018_g N_A_2067_74#_c_1699_n 0.0030803f $X=13.25 $Y=2.75 $X2=0
+ $Y2=0
cc_929 N_SET_B_c_1182_n N_A_2067_74#_c_1699_n 0.00246686f $X=13.27 $Y=1.97 $X2=0
+ $Y2=0
cc_930 N_SET_B_M1018_g N_A_2067_74#_c_1685_n 0.00106241f $X=13.25 $Y=2.75 $X2=0
+ $Y2=0
cc_931 SET_B N_A_2067_74#_c_1685_n 0.00131157f $X=13.115 $Y=1.58 $X2=0 $Y2=0
cc_932 N_SET_B_c_1176_n N_A_2067_74#_c_1685_n 8.41851e-19 $X=13.27 $Y=1.465
+ $X2=0 $Y2=0
cc_933 N_SET_B_c_1177_n N_A_2067_74#_c_1685_n 0.0411607f $X=13.27 $Y=1.465 $X2=0
+ $Y2=0
cc_934 N_SET_B_M1018_g N_A_2067_74#_c_1686_n 0.0146339f $X=13.25 $Y=2.75 $X2=0
+ $Y2=0
cc_935 N_SET_B_c_1171_n N_A_2067_74#_c_1686_n 0.0214924f $X=13.27 $Y=1.805 $X2=0
+ $Y2=0
cc_936 N_SET_B_c_1172_n N_A_2067_74#_c_1701_n 0.00914033f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_937 N_SET_B_c_1172_n N_A_2067_74#_c_1688_n 0.0224912f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_938 N_SET_B_M1034_g N_VPWR_c_1961_n 0.0016907f $X=7.985 $Y=2.525 $X2=0 $Y2=0
cc_939 N_SET_B_M1018_g N_VPWR_c_1963_n 0.0030528f $X=13.25 $Y=2.75 $X2=0 $Y2=0
cc_940 N_SET_B_M1018_g N_VPWR_c_1973_n 0.005209f $X=13.25 $Y=2.75 $X2=0 $Y2=0
cc_941 N_SET_B_M1018_g N_VPWR_c_1956_n 0.00987509f $X=13.25 $Y=2.75 $X2=0 $Y2=0
cc_942 N_SET_B_c_1172_n N_A_1789_424#_c_2275_n 0.00328854f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_943 N_SET_B_c_1172_n N_A_1789_424#_c_2269_n 0.00159688f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_944 N_SET_B_c_1172_n N_A_1789_424#_c_2273_n 0.00197494f $X=13.055 $Y=1.665
+ $X2=0 $Y2=0
cc_945 N_SET_B_M1014_g N_VGND_c_2410_n 0.0109278f $X=8.15 $Y=0.58 $X2=0 $Y2=0
cc_946 N_SET_B_M1021_g N_VGND_c_2412_n 0.0125621f $X=13.21 $Y=0.58 $X2=0 $Y2=0
cc_947 N_SET_B_M1021_g N_VGND_c_2422_n 0.00383152f $X=13.21 $Y=0.58 $X2=0 $Y2=0
cc_948 N_SET_B_M1014_g N_VGND_c_2431_n 0.00383152f $X=8.15 $Y=0.58 $X2=0 $Y2=0
cc_949 N_SET_B_M1014_g N_VGND_c_2439_n 0.0075725f $X=8.15 $Y=0.58 $X2=0 $Y2=0
cc_950 N_SET_B_M1021_g N_VGND_c_2439_n 0.0075725f $X=13.21 $Y=0.58 $X2=0 $Y2=0
cc_951 N_A_619_368#_c_1317_n N_A_2513_258#_M1016_g 0.0298674f $X=12.28 $Y=3.065
+ $X2=0 $Y2=0
cc_952 N_A_619_368#_c_1316_n N_A_2513_258#_M1020_g 0.00691527f $X=12.28 $Y=1.23
+ $X2=0 $Y2=0
cc_953 N_A_619_368#_c_1318_n N_A_2513_258#_M1020_g 0.0445874f $X=12.43 $Y=0.9
+ $X2=0 $Y2=0
cc_954 N_A_619_368#_c_1316_n N_A_2513_258#_c_1575_n 5.5693e-19 $X=12.28 $Y=1.23
+ $X2=0 $Y2=0
cc_955 N_A_619_368#_c_1317_n N_A_2513_258#_c_1575_n 8.7256e-19 $X=12.28 $Y=3.065
+ $X2=0 $Y2=0
cc_956 N_A_619_368#_c_1317_n N_A_2513_258#_c_1576_n 0.0424432f $X=12.28 $Y=3.065
+ $X2=0 $Y2=0
cc_957 N_A_619_368#_c_1316_n N_A_2513_258#_c_1578_n 0.00113941f $X=12.28 $Y=1.23
+ $X2=0 $Y2=0
cc_958 N_A_619_368#_c_1336_n N_A_2067_74#_c_1719_n 0.00713358f $X=10.265
+ $Y=2.045 $X2=0 $Y2=0
cc_959 N_A_619_368#_c_1337_n N_A_2067_74#_c_1695_n 3.96713e-19 $X=10.625 $Y=1.97
+ $X2=0 $Y2=0
cc_960 N_A_619_368#_c_1339_n N_A_2067_74#_c_1695_n 0.0140765f $X=10.715 $Y=2.045
+ $X2=0 $Y2=0
cc_961 N_A_619_368#_c_1340_n N_A_2067_74#_c_1695_n 0.00743694f $X=11.16 $Y=1.97
+ $X2=0 $Y2=0
cc_962 N_A_619_368#_c_1341_n N_A_2067_74#_c_1695_n 0.0136066f $X=11.235 $Y=3.065
+ $X2=0 $Y2=0
cc_963 N_A_619_368#_c_1349_n N_A_2067_74#_c_1695_n 0.00155547f $X=10.715 $Y=1.97
+ $X2=0 $Y2=0
cc_964 N_A_619_368#_c_1352_n N_A_2067_74#_c_1695_n 0.0845967f $X=11.72 $Y=1.785
+ $X2=0 $Y2=0
cc_965 N_A_619_368#_c_1336_n N_A_2067_74#_c_1720_n 0.00433521f $X=10.265
+ $Y=2.045 $X2=0 $Y2=0
cc_966 N_A_619_368#_c_1337_n N_A_2067_74#_c_1720_n 0.00402515f $X=10.625 $Y=1.97
+ $X2=0 $Y2=0
cc_967 N_A_619_368#_c_1338_n N_A_2067_74#_c_1720_n 3.37521e-19 $X=10.355 $Y=1.97
+ $X2=0 $Y2=0
cc_968 N_A_619_368#_c_1352_n N_A_2067_74#_c_1720_n 0.0184869f $X=11.72 $Y=1.785
+ $X2=0 $Y2=0
cc_969 N_A_619_368#_c_1318_n N_A_2067_74#_c_1754_n 0.00697999f $X=12.43 $Y=0.9
+ $X2=0 $Y2=0
cc_970 N_A_619_368#_c_1322_n N_A_2067_74#_c_1754_n 0.00936164f $X=12.205
+ $Y=1.065 $X2=0 $Y2=0
cc_971 N_A_619_368#_c_1326_n N_A_2067_74#_c_1754_n 0.0270286f $X=11.885 $Y=1.065
+ $X2=0 $Y2=0
cc_972 N_A_619_368#_c_1322_n N_A_2067_74#_c_1684_n 0.00342686f $X=12.205
+ $Y=1.065 $X2=0 $Y2=0
cc_973 N_A_619_368#_c_1352_n N_A_2067_74#_c_1684_n 0.00260498f $X=11.72 $Y=1.785
+ $X2=0 $Y2=0
cc_974 N_A_619_368#_c_1326_n N_A_2067_74#_c_1684_n 0.00977037f $X=11.885
+ $Y=1.065 $X2=0 $Y2=0
cc_975 N_A_619_368#_c_1317_n N_A_2067_74#_c_1696_n 0.0118527f $X=12.28 $Y=3.065
+ $X2=0 $Y2=0
cc_976 N_A_619_368#_c_1317_n N_A_2067_74#_c_1697_n 5.21162e-19 $X=12.28 $Y=3.065
+ $X2=0 $Y2=0
cc_977 N_A_619_368#_c_1341_n N_A_2067_74#_c_1701_n 8.69551e-19 $X=11.235
+ $Y=3.065 $X2=0 $Y2=0
cc_978 N_A_619_368#_c_1317_n N_A_2067_74#_c_1701_n 0.013226f $X=12.28 $Y=3.065
+ $X2=0 $Y2=0
cc_979 N_A_619_368#_c_1352_n N_A_2067_74#_c_1701_n 0.0197333f $X=11.72 $Y=1.785
+ $X2=0 $Y2=0
cc_980 N_A_619_368#_c_1316_n N_A_2067_74#_c_1688_n 0.01572f $X=12.28 $Y=1.23
+ $X2=0 $Y2=0
cc_981 N_A_619_368#_c_1317_n N_A_2067_74#_c_1688_n 0.0183062f $X=12.28 $Y=3.065
+ $X2=0 $Y2=0
cc_982 N_A_619_368#_c_1318_n N_A_2067_74#_c_1688_n 0.00528607f $X=12.43 $Y=0.9
+ $X2=0 $Y2=0
cc_983 N_A_619_368#_c_1352_n N_A_2067_74#_c_1688_n 0.0133324f $X=11.72 $Y=1.785
+ $X2=0 $Y2=0
cc_984 N_A_619_368#_c_1326_n N_A_2067_74#_c_1688_n 0.0582461f $X=11.885 $Y=1.065
+ $X2=0 $Y2=0
cc_985 N_A_619_368#_c_1350_n N_VPWR_M1036_d 0.00803991f $X=4.39 $Y=1.875 $X2=0
+ $Y2=0
cc_986 N_A_619_368#_M1002_g N_VPWR_c_1959_n 8.89341e-19 $X=5.93 $Y=2.525 $X2=0
+ $Y2=0
cc_987 N_A_619_368#_c_1334_n N_VPWR_c_1959_n 0.0390231f $X=8.72 $Y=3.15 $X2=0
+ $Y2=0
cc_988 N_A_619_368#_c_1334_n N_VPWR_c_1960_n 0.0322942f $X=8.72 $Y=3.15 $X2=0
+ $Y2=0
cc_989 N_A_619_368#_c_1334_n N_VPWR_c_1961_n 0.0244708f $X=8.72 $Y=3.15 $X2=0
+ $Y2=0
cc_990 N_A_619_368#_c_1335_n N_VPWR_c_1961_n 0.0129384f $X=8.795 $Y=3.075 $X2=0
+ $Y2=0
cc_991 N_A_619_368#_c_1334_n N_VPWR_c_1962_n 0.0020984f $X=8.72 $Y=3.15 $X2=0
+ $Y2=0
cc_992 N_A_619_368#_c_1335_n N_VPWR_c_1962_n 6.04219e-19 $X=8.795 $Y=3.075 $X2=0
+ $Y2=0
cc_993 N_A_619_368#_c_1317_n N_VPWR_c_1963_n 0.00189459f $X=12.28 $Y=3.065 $X2=0
+ $Y2=0
cc_994 N_A_619_368#_c_1334_n N_VPWR_c_1969_n 0.00796123f $X=8.72 $Y=3.15 $X2=0
+ $Y2=0
cc_995 N_A_619_368#_c_1336_n N_VPWR_c_1971_n 0.00333926f $X=10.265 $Y=2.045
+ $X2=0 $Y2=0
cc_996 N_A_619_368#_c_1339_n N_VPWR_c_1971_n 0.00333896f $X=10.715 $Y=2.045
+ $X2=0 $Y2=0
cc_997 N_A_619_368#_c_1343_n N_VPWR_c_1971_n 0.0286449f $X=11.31 $Y=3.14 $X2=0
+ $Y2=0
cc_998 N_A_619_368#_M1046_g N_VPWR_c_1979_n 0.0050621f $X=4.295 $Y=2.4 $X2=0
+ $Y2=0
cc_999 N_A_619_368#_c_1332_n N_VPWR_c_1979_n 0.0376458f $X=4.925 $Y=3.15 $X2=0
+ $Y2=0
cc_1000 N_A_619_368#_M1046_g N_VPWR_c_1985_n 0.00790916f $X=4.295 $Y=2.4 $X2=0
+ $Y2=0
cc_1001 N_A_619_368#_c_1332_n N_VPWR_c_1985_n 0.00232174f $X=4.925 $Y=3.15 $X2=0
+ $Y2=0
cc_1002 N_A_619_368#_M1046_g N_VPWR_c_1956_n 0.00995335f $X=4.295 $Y=2.4 $X2=0
+ $Y2=0
cc_1003 N_A_619_368#_c_1331_n N_VPWR_c_1956_n 0.0215278f $X=5.84 $Y=3.15 $X2=0
+ $Y2=0
cc_1004 N_A_619_368#_c_1332_n N_VPWR_c_1956_n 0.00600227f $X=4.925 $Y=3.15 $X2=0
+ $Y2=0
cc_1005 N_A_619_368#_c_1334_n N_VPWR_c_1956_n 0.0672811f $X=8.72 $Y=3.15 $X2=0
+ $Y2=0
cc_1006 N_A_619_368#_c_1336_n N_VPWR_c_1956_n 0.00422798f $X=10.265 $Y=2.045
+ $X2=0 $Y2=0
cc_1007 N_A_619_368#_c_1339_n N_VPWR_c_1956_n 0.00423488f $X=10.715 $Y=2.045
+ $X2=0 $Y2=0
cc_1008 N_A_619_368#_c_1342_n N_VPWR_c_1956_n 0.0290163f $X=12.205 $Y=3.14 $X2=0
+ $Y2=0
cc_1009 N_A_619_368#_c_1343_n N_VPWR_c_1956_n 0.0114038f $X=11.31 $Y=3.14 $X2=0
+ $Y2=0
cc_1010 N_A_619_368#_c_1348_n N_VPWR_c_1956_n 0.00445015f $X=5.93 $Y=3.15 $X2=0
+ $Y2=0
cc_1011 N_A_619_368#_c_1353_n N_A_307_74#_c_2154_n 0.0143692f $X=3.545 $Y=1.965
+ $X2=0 $Y2=0
cc_1012 N_A_619_368#_M1036_s N_A_307_74#_c_2159_n 0.00779918f $X=3.095 $Y=1.84
+ $X2=0 $Y2=0
cc_1013 N_A_619_368#_c_1350_n N_A_307_74#_c_2159_n 0.00476087f $X=4.39 $Y=1.875
+ $X2=0 $Y2=0
cc_1014 N_A_619_368#_c_1353_n N_A_307_74#_c_2159_n 0.0308023f $X=3.545 $Y=1.965
+ $X2=0 $Y2=0
cc_1015 N_A_619_368#_M1046_g N_A_307_74#_c_2160_n 0.0183131f $X=4.295 $Y=2.4
+ $X2=0 $Y2=0
cc_1016 N_A_619_368#_c_1330_n N_A_307_74#_c_2160_n 0.013162f $X=4.85 $Y=3.075
+ $X2=0 $Y2=0
cc_1017 N_A_619_368#_c_1320_n N_A_307_74#_c_2160_n 7.95206e-19 $X=4.775 $Y=1.515
+ $X2=0 $Y2=0
cc_1018 N_A_619_368#_c_1350_n N_A_307_74#_c_2160_n 0.0537833f $X=4.39 $Y=1.875
+ $X2=0 $Y2=0
cc_1019 N_A_619_368#_M1046_g N_A_307_74#_c_2197_n 0.00374807f $X=4.295 $Y=2.4
+ $X2=0 $Y2=0
cc_1020 N_A_619_368#_c_1350_n N_A_307_74#_c_2197_n 0.0129609f $X=4.39 $Y=1.875
+ $X2=0 $Y2=0
cc_1021 N_A_619_368#_c_1353_n N_A_307_74#_c_2197_n 6.86671e-19 $X=3.545 $Y=1.965
+ $X2=0 $Y2=0
cc_1022 N_A_619_368#_c_1313_n N_A_307_74#_c_2155_n 0.00547833f $X=5.195 $Y=0.975
+ $X2=0 $Y2=0
cc_1023 N_A_619_368#_c_1315_n N_A_307_74#_c_2155_n 0.00434355f $X=5.27 $Y=0.9
+ $X2=0 $Y2=0
cc_1024 N_A_619_368#_M1046_g N_A_307_74#_c_2162_n 9.57396e-19 $X=4.295 $Y=2.4
+ $X2=0 $Y2=0
cc_1025 N_A_619_368#_c_1330_n N_A_307_74#_c_2162_n 0.0176353f $X=4.85 $Y=3.075
+ $X2=0 $Y2=0
cc_1026 N_A_619_368#_M1002_g N_A_307_74#_c_2162_n 2.26734e-19 $X=5.93 $Y=2.525
+ $X2=0 $Y2=0
cc_1027 N_A_619_368#_M1035_g N_A_307_74#_c_2156_n 0.00150815f $X=4.28 $Y=0.74
+ $X2=0 $Y2=0
cc_1028 N_A_619_368#_M1046_g N_A_307_74#_c_2156_n 9.70488e-19 $X=4.295 $Y=2.4
+ $X2=0 $Y2=0
cc_1029 N_A_619_368#_c_1312_n N_A_307_74#_c_2156_n 0.00891258f $X=4.85 $Y=1.35
+ $X2=0 $Y2=0
cc_1030 N_A_619_368#_c_1330_n N_A_307_74#_c_2156_n 0.0105447f $X=4.85 $Y=3.075
+ $X2=0 $Y2=0
cc_1031 N_A_619_368#_c_1313_n N_A_307_74#_c_2156_n 0.0101656f $X=5.195 $Y=0.975
+ $X2=0 $Y2=0
cc_1032 N_A_619_368#_c_1314_n N_A_307_74#_c_2156_n 0.00285843f $X=4.925 $Y=0.975
+ $X2=0 $Y2=0
cc_1033 N_A_619_368#_c_1321_n N_A_307_74#_c_2156_n 0.00807793f $X=4.85 $Y=1.515
+ $X2=0 $Y2=0
cc_1034 N_A_619_368#_c_1350_n N_A_307_74#_c_2156_n 0.0137141f $X=4.39 $Y=1.875
+ $X2=0 $Y2=0
cc_1035 N_A_619_368#_c_1325_n N_A_307_74#_c_2156_n 0.0317952f $X=4.555 $Y=1.515
+ $X2=0 $Y2=0
cc_1036 N_A_619_368#_c_1352_n N_A_1789_424#_c_2275_n 0.0254537f $X=11.72
+ $Y=1.785 $X2=0 $Y2=0
cc_1037 N_A_619_368#_c_1352_n N_A_1789_424#_c_2269_n 0.0149891f $X=11.72
+ $Y=1.785 $X2=0 $Y2=0
cc_1038 N_A_619_368#_c_1336_n N_A_1789_424#_c_2270_n 0.0139927f $X=10.265
+ $Y=2.045 $X2=0 $Y2=0
cc_1039 N_A_619_368#_c_1339_n N_A_1789_424#_c_2270_n 0.0136253f $X=10.715
+ $Y=2.045 $X2=0 $Y2=0
cc_1040 N_A_619_368#_c_1341_n N_A_1789_424#_c_2270_n 0.00229358f $X=11.235
+ $Y=3.065 $X2=0 $Y2=0
cc_1041 N_A_619_368#_c_1336_n N_A_1789_424#_c_2272_n 7.36854e-19 $X=10.265
+ $Y=2.045 $X2=0 $Y2=0
cc_1042 N_A_619_368#_c_1339_n N_A_1789_424#_c_2272_n 0.00835326f $X=10.715
+ $Y=2.045 $X2=0 $Y2=0
cc_1043 N_A_619_368#_c_1340_n N_A_1789_424#_c_2272_n 9.46521e-19 $X=11.16
+ $Y=1.97 $X2=0 $Y2=0
cc_1044 N_A_619_368#_c_1341_n N_A_1789_424#_c_2272_n 0.00529022f $X=11.235
+ $Y=3.065 $X2=0 $Y2=0
cc_1045 N_A_619_368#_c_1335_n N_A_1789_424#_c_2273_n 0.0126169f $X=8.795
+ $Y=3.075 $X2=0 $Y2=0
cc_1046 N_A_619_368#_c_1352_n N_A_1789_424#_c_2273_n 0.00920624f $X=11.72
+ $Y=1.785 $X2=0 $Y2=0
cc_1047 N_A_619_368#_c_1328_n N_A_1789_424#_c_2273_n 0.00326139f $X=8.9 $Y=1.795
+ $X2=0 $Y2=0
cc_1048 N_A_619_368#_c_1355_n N_A_1789_424#_c_2273_n 0.0108129f $X=9.065
+ $Y=1.822 $X2=0 $Y2=0
cc_1049 N_A_619_368#_c_1341_n N_A_2277_455#_c_2317_n 0.00568213f $X=11.235
+ $Y=3.065 $X2=0 $Y2=0
cc_1050 N_A_619_368#_c_1317_n N_A_2277_455#_c_2317_n 0.00160564f $X=12.28
+ $Y=3.065 $X2=0 $Y2=0
cc_1051 N_A_619_368#_c_1342_n N_A_2277_455#_c_2318_n 0.00874016f $X=12.205
+ $Y=3.14 $X2=0 $Y2=0
cc_1052 N_A_619_368#_c_1317_n N_A_2277_455#_c_2318_n 0.0120677f $X=12.28
+ $Y=3.065 $X2=0 $Y2=0
cc_1053 N_A_619_368#_c_1341_n N_A_2277_455#_c_2319_n 0.00422063f $X=11.235
+ $Y=3.065 $X2=0 $Y2=0
cc_1054 N_A_619_368#_c_1342_n N_A_2277_455#_c_2319_n 0.00545232f $X=12.205
+ $Y=3.14 $X2=0 $Y2=0
cc_1055 N_A_619_368#_c_1317_n N_A_2277_455#_c_2320_n 0.00645514f $X=12.28
+ $Y=3.065 $X2=0 $Y2=0
cc_1056 N_A_619_368#_c_1323_n N_VGND_c_2407_n 0.0316927f $X=3.565 $Y=0.505 $X2=0
+ $Y2=0
cc_1057 N_A_619_368#_M1035_g N_VGND_c_2408_n 0.00470925f $X=4.28 $Y=0.74 $X2=0
+ $Y2=0
cc_1058 N_A_619_368#_c_1323_n N_VGND_c_2408_n 0.025141f $X=3.565 $Y=0.505 $X2=0
+ $Y2=0
cc_1059 N_A_619_368#_c_1318_n N_VGND_c_2422_n 0.0042336f $X=12.43 $Y=0.9 $X2=0
+ $Y2=0
cc_1060 N_A_619_368#_c_1323_n N_VGND_c_2429_n 0.0126849f $X=3.565 $Y=0.505 $X2=0
+ $Y2=0
cc_1061 N_A_619_368#_M1035_g N_VGND_c_2430_n 0.00430908f $X=4.28 $Y=0.74 $X2=0
+ $Y2=0
cc_1062 N_A_619_368#_c_1315_n N_VGND_c_2430_n 9.15902e-19 $X=5.27 $Y=0.9 $X2=0
+ $Y2=0
cc_1063 N_A_619_368#_M1035_g N_VGND_c_2439_n 0.00821169f $X=4.28 $Y=0.74 $X2=0
+ $Y2=0
cc_1064 N_A_619_368#_c_1318_n N_VGND_c_2439_n 0.0078709f $X=12.43 $Y=0.9 $X2=0
+ $Y2=0
cc_1065 N_A_619_368#_c_1323_n N_VGND_c_2439_n 0.0101411f $X=3.565 $Y=0.505 $X2=0
+ $Y2=0
cc_1066 N_A_2513_258#_c_1577_n N_A_2067_74#_M1040_g 0.0115126f $X=13.77 $Y=1.045
+ $X2=0 $Y2=0
cc_1067 N_A_2513_258#_c_1579_n N_A_2067_74#_M1040_g 0.0125515f $X=13.935 $Y=0.58
+ $X2=0 $Y2=0
cc_1068 N_A_2513_258#_c_1580_n N_A_2067_74#_M1040_g 0.00477786f $X=14.23 $Y=2.48
+ $X2=0 $Y2=0
cc_1069 N_A_2513_258#_c_1581_n N_A_2067_74#_M1040_g 0.00461905f $X=14.042
+ $Y=1.045 $X2=0 $Y2=0
cc_1070 N_A_2513_258#_c_1580_n N_A_2067_74#_c_1670_n 0.0153375f $X=14.23 $Y=2.48
+ $X2=0 $Y2=0
cc_1071 N_A_2513_258#_c_1580_n N_A_2067_74#_c_1689_n 0.00918623f $X=14.23
+ $Y=2.48 $X2=0 $Y2=0
cc_1072 N_A_2513_258#_c_1587_n N_A_2067_74#_c_1690_n 0.00865699f $X=14.23
+ $Y=2.695 $X2=0 $Y2=0
cc_1073 N_A_2513_258#_c_1580_n N_A_2067_74#_M1045_g 0.00654001f $X=14.23 $Y=2.48
+ $X2=0 $Y2=0
cc_1074 N_A_2513_258#_c_1587_n N_A_2067_74#_M1045_g 0.0110144f $X=14.23 $Y=2.695
+ $X2=0 $Y2=0
cc_1075 N_A_2513_258#_c_1579_n N_A_2067_74#_M1023_g 0.00441492f $X=13.935
+ $Y=0.58 $X2=0 $Y2=0
cc_1076 N_A_2513_258#_c_1580_n N_A_2067_74#_M1023_g 0.0029433f $X=14.23 $Y=2.48
+ $X2=0 $Y2=0
cc_1077 N_A_2513_258#_c_1581_n N_A_2067_74#_M1023_g 0.00323313f $X=14.042
+ $Y=1.045 $X2=0 $Y2=0
cc_1078 N_A_2513_258#_c_1580_n N_A_2067_74#_M1004_g 0.00713224f $X=14.23 $Y=2.48
+ $X2=0 $Y2=0
cc_1079 N_A_2513_258#_c_1581_n N_A_2067_74#_c_1679_n 0.0080581f $X=14.042
+ $Y=1.045 $X2=0 $Y2=0
cc_1080 N_A_2513_258#_M1020_g N_A_2067_74#_c_1754_n 0.00165231f $X=12.82 $Y=0.58
+ $X2=0 $Y2=0
cc_1081 N_A_2513_258#_M1016_g N_A_2067_74#_c_1696_n 0.00105371f $X=12.8 $Y=2.75
+ $X2=0 $Y2=0
cc_1082 N_A_2513_258#_M1016_g N_A_2067_74#_c_1697_n 0.0164508f $X=12.8 $Y=2.75
+ $X2=0 $Y2=0
cc_1083 N_A_2513_258#_c_1584_n N_A_2067_74#_c_1697_n 9.90657e-19 $X=12.73
+ $Y=1.96 $X2=0 $Y2=0
cc_1084 N_A_2513_258#_c_1575_n N_A_2067_74#_c_1697_n 0.0231756f $X=12.73
+ $Y=1.455 $X2=0 $Y2=0
cc_1085 N_A_2513_258#_M1016_g N_A_2067_74#_c_1698_n 0.00114505f $X=12.8 $Y=2.75
+ $X2=0 $Y2=0
cc_1086 N_A_2513_258#_c_1580_n N_A_2067_74#_c_1698_n 0.00614772f $X=14.23
+ $Y=2.48 $X2=0 $Y2=0
cc_1087 N_A_2513_258#_c_1587_n N_A_2067_74#_c_1698_n 0.0296213f $X=14.23
+ $Y=2.695 $X2=0 $Y2=0
cc_1088 N_A_2513_258#_c_1580_n N_A_2067_74#_c_1699_n 0.0128267f $X=14.23 $Y=2.48
+ $X2=0 $Y2=0
cc_1089 N_A_2513_258#_c_1587_n N_A_2067_74#_c_1699_n 0.00797082f $X=14.23
+ $Y=2.695 $X2=0 $Y2=0
cc_1090 N_A_2513_258#_c_1577_n N_A_2067_74#_c_1685_n 0.00941168f $X=13.77
+ $Y=1.045 $X2=0 $Y2=0
cc_1091 N_A_2513_258#_c_1580_n N_A_2067_74#_c_1685_n 0.062535f $X=14.23 $Y=2.48
+ $X2=0 $Y2=0
cc_1092 N_A_2513_258#_c_1581_n N_A_2067_74#_c_1685_n 0.0180767f $X=14.042
+ $Y=1.045 $X2=0 $Y2=0
cc_1093 N_A_2513_258#_c_1580_n N_A_2067_74#_c_1686_n 0.0118829f $X=14.23 $Y=2.48
+ $X2=0 $Y2=0
cc_1094 N_A_2513_258#_M1016_g N_A_2067_74#_c_1688_n 0.00372173f $X=12.8 $Y=2.75
+ $X2=0 $Y2=0
cc_1095 N_A_2513_258#_M1020_g N_A_2067_74#_c_1688_n 0.00178906f $X=12.82 $Y=0.58
+ $X2=0 $Y2=0
cc_1096 N_A_2513_258#_c_1575_n N_A_2067_74#_c_1688_n 0.0605029f $X=12.73
+ $Y=1.455 $X2=0 $Y2=0
cc_1097 N_A_2513_258#_c_1576_n N_A_2067_74#_c_1688_n 0.0033491f $X=12.73
+ $Y=1.455 $X2=0 $Y2=0
cc_1098 N_A_2513_258#_c_1578_n N_A_2067_74#_c_1688_n 0.0137215f $X=12.895
+ $Y=1.045 $X2=0 $Y2=0
cc_1099 N_A_2513_258#_M1016_g N_VPWR_c_1963_n 0.00181319f $X=12.8 $Y=2.75 $X2=0
+ $Y2=0
cc_1100 N_A_2513_258#_c_1580_n N_VPWR_c_1964_n 0.0476064f $X=14.23 $Y=2.48 $X2=0
+ $Y2=0
cc_1101 N_A_2513_258#_c_1587_n N_VPWR_c_1964_n 0.0325137f $X=14.23 $Y=2.695
+ $X2=0 $Y2=0
cc_1102 N_A_2513_258#_M1016_g N_VPWR_c_1971_n 0.0051767f $X=12.8 $Y=2.75 $X2=0
+ $Y2=0
cc_1103 N_A_2513_258#_c_1587_n N_VPWR_c_1973_n 0.0145493f $X=14.23 $Y=2.695
+ $X2=0 $Y2=0
cc_1104 N_A_2513_258#_M1016_g N_VPWR_c_1956_n 0.00978534f $X=12.8 $Y=2.75 $X2=0
+ $Y2=0
cc_1105 N_A_2513_258#_c_1587_n N_VPWR_c_1956_n 0.0153061f $X=14.23 $Y=2.695
+ $X2=0 $Y2=0
cc_1106 N_A_2513_258#_M1016_g N_A_2277_455#_c_2318_n 0.0037636f $X=12.8 $Y=2.75
+ $X2=0 $Y2=0
cc_1107 N_A_2513_258#_M1016_g N_A_2277_455#_c_2320_n 0.00521172f $X=12.8 $Y=2.75
+ $X2=0 $Y2=0
cc_1108 N_A_2513_258#_c_1580_n N_Q_N_c_2350_n 0.0210604f $X=14.23 $Y=2.48 $X2=0
+ $Y2=0
cc_1109 N_A_2513_258#_c_1581_n N_Q_N_c_2350_n 0.00612134f $X=14.042 $Y=1.045
+ $X2=0 $Y2=0
cc_1110 N_A_2513_258#_M1020_g N_VGND_c_2412_n 0.00274214f $X=12.82 $Y=0.58 $X2=0
+ $Y2=0
cc_1111 N_A_2513_258#_c_1577_n N_VGND_c_2412_n 0.0243627f $X=13.77 $Y=1.045
+ $X2=0 $Y2=0
cc_1112 N_A_2513_258#_c_1579_n N_VGND_c_2412_n 0.0165294f $X=13.935 $Y=0.58
+ $X2=0 $Y2=0
cc_1113 N_A_2513_258#_c_1579_n N_VGND_c_2413_n 0.0280059f $X=13.935 $Y=0.58
+ $X2=0 $Y2=0
cc_1114 N_A_2513_258#_M1020_g N_VGND_c_2422_n 0.00461464f $X=12.82 $Y=0.58 $X2=0
+ $Y2=0
cc_1115 N_A_2513_258#_c_1579_n N_VGND_c_2424_n 0.0145639f $X=13.935 $Y=0.58
+ $X2=0 $Y2=0
cc_1116 N_A_2513_258#_M1020_g N_VGND_c_2439_n 0.00908738f $X=12.82 $Y=0.58 $X2=0
+ $Y2=0
cc_1117 N_A_2513_258#_c_1579_n N_VGND_c_2439_n 0.0119984f $X=13.935 $Y=0.58
+ $X2=0 $Y2=0
cc_1118 N_A_2067_74#_M1000_g N_A_3177_368#_M1047_g 0.0213843f $X=16.255 $Y=2.34
+ $X2=0 $Y2=0
cc_1119 N_A_2067_74#_M1012_g N_A_3177_368#_M1001_g 0.0139828f $X=16.27 $Y=0.79
+ $X2=0 $Y2=0
cc_1120 N_A_2067_74#_M1025_g N_A_3177_368#_c_1892_n 0.00365834f $X=15.23 $Y=0.74
+ $X2=0 $Y2=0
cc_1121 N_A_2067_74#_M1012_g N_A_3177_368#_c_1892_n 0.016091f $X=16.27 $Y=0.79
+ $X2=0 $Y2=0
cc_1122 N_A_2067_74#_M1029_g N_A_3177_368#_c_1893_n 0.00689158f $X=15.245 $Y=2.4
+ $X2=0 $Y2=0
cc_1123 N_A_2067_74#_M1000_g N_A_3177_368#_c_1893_n 0.0218825f $X=16.255 $Y=2.34
+ $X2=0 $Y2=0
cc_1124 N_A_2067_74#_M1000_g N_A_3177_368#_c_1894_n 0.00959884f $X=16.255
+ $Y=2.34 $X2=0 $Y2=0
cc_1125 N_A_2067_74#_c_1682_n N_A_3177_368#_c_1894_n 0.0090289f $X=16.255
+ $Y=1.375 $X2=0 $Y2=0
cc_1126 N_A_2067_74#_M1029_g N_A_3177_368#_c_1895_n 0.00515495f $X=15.245 $Y=2.4
+ $X2=0 $Y2=0
cc_1127 N_A_2067_74#_c_1676_n N_A_3177_368#_c_1895_n 0.0204535f $X=16.165
+ $Y=1.375 $X2=0 $Y2=0
cc_1128 N_A_2067_74#_M1000_g N_A_3177_368#_c_1895_n 0.00582757f $X=16.255
+ $Y=2.34 $X2=0 $Y2=0
cc_1129 N_A_2067_74#_c_1682_n N_A_3177_368#_c_1895_n 7.76856e-19 $X=16.255
+ $Y=1.375 $X2=0 $Y2=0
cc_1130 N_A_2067_74#_c_1682_n N_A_3177_368#_c_1896_n 0.0214984f $X=16.255
+ $Y=1.375 $X2=0 $Y2=0
cc_1131 N_A_2067_74#_c_1697_n N_VPWR_c_1963_n 0.0122262f $X=13.31 $Y=2.225 $X2=0
+ $Y2=0
cc_1132 N_A_2067_74#_c_1698_n N_VPWR_c_1963_n 0.01643f $X=13.475 $Y=2.75 $X2=0
+ $Y2=0
cc_1133 N_A_2067_74#_c_1670_n N_VPWR_c_1964_n 0.00428832f $X=14.705 $Y=1.375
+ $X2=0 $Y2=0
cc_1134 N_A_2067_74#_c_1689_n N_VPWR_c_1964_n 0.0079696f $X=14.17 $Y=2.235 $X2=0
+ $Y2=0
cc_1135 N_A_2067_74#_M1004_g N_VPWR_c_1964_n 0.00346304f $X=14.795 $Y=2.4 $X2=0
+ $Y2=0
cc_1136 N_A_2067_74#_M1004_g N_VPWR_c_1965_n 7.38193e-19 $X=14.795 $Y=2.4 $X2=0
+ $Y2=0
cc_1137 N_A_2067_74#_M1029_g N_VPWR_c_1965_n 0.0220886f $X=15.245 $Y=2.4 $X2=0
+ $Y2=0
cc_1138 N_A_2067_74#_c_1676_n N_VPWR_c_1965_n 0.00694774f $X=16.165 $Y=1.375
+ $X2=0 $Y2=0
cc_1139 N_A_2067_74#_M1000_g N_VPWR_c_1965_n 0.00476325f $X=16.255 $Y=2.34 $X2=0
+ $Y2=0
cc_1140 N_A_2067_74#_M1000_g N_VPWR_c_1966_n 0.012418f $X=16.255 $Y=2.34 $X2=0
+ $Y2=0
cc_1141 N_A_2067_74#_M1045_g N_VPWR_c_1973_n 0.00493294f $X=14.26 $Y=2.68 $X2=0
+ $Y2=0
cc_1142 N_A_2067_74#_c_1698_n N_VPWR_c_1973_n 0.0145333f $X=13.475 $Y=2.75 $X2=0
+ $Y2=0
cc_1143 N_A_2067_74#_M1004_g N_VPWR_c_1975_n 0.00515235f $X=14.795 $Y=2.4 $X2=0
+ $Y2=0
cc_1144 N_A_2067_74#_M1029_g N_VPWR_c_1975_n 0.00460063f $X=15.245 $Y=2.4 $X2=0
+ $Y2=0
cc_1145 N_A_2067_74#_M1000_g N_VPWR_c_1980_n 0.00567889f $X=16.255 $Y=2.34 $X2=0
+ $Y2=0
cc_1146 N_A_2067_74#_M1045_g N_VPWR_c_1956_n 0.00628405f $X=14.26 $Y=2.68 $X2=0
+ $Y2=0
cc_1147 N_A_2067_74#_M1004_g N_VPWR_c_1956_n 0.00969055f $X=14.795 $Y=2.4 $X2=0
+ $Y2=0
cc_1148 N_A_2067_74#_M1029_g N_VPWR_c_1956_n 0.00908554f $X=15.245 $Y=2.4 $X2=0
+ $Y2=0
cc_1149 N_A_2067_74#_M1000_g N_VPWR_c_1956_n 0.00610055f $X=16.255 $Y=2.34 $X2=0
+ $Y2=0
cc_1150 N_A_2067_74#_c_1698_n N_VPWR_c_1956_n 0.0119681f $X=13.475 $Y=2.75 $X2=0
+ $Y2=0
cc_1151 N_A_2067_74#_c_1695_n N_A_1789_424#_M1031_s 0.00237053f $X=11.82
+ $Y=2.125 $X2=0 $Y2=0
cc_1152 N_A_2067_74#_c_1720_n N_A_1789_424#_c_2269_n 0.00476347f $X=10.575
+ $Y=2.125 $X2=0 $Y2=0
cc_1153 N_A_2067_74#_M1028_d N_A_1789_424#_c_2270_n 0.00179769f $X=10.355
+ $Y=2.12 $X2=0 $Y2=0
cc_1154 N_A_2067_74#_c_1719_n N_A_1789_424#_c_2270_n 0.0118192f $X=10.49 $Y=2.46
+ $X2=0 $Y2=0
cc_1155 N_A_2067_74#_c_1695_n N_A_1789_424#_c_2272_n 0.0219539f $X=11.82
+ $Y=2.125 $X2=0 $Y2=0
cc_1156 N_A_2067_74#_c_1695_n N_A_2277_455#_c_2317_n 0.0202283f $X=11.82
+ $Y=2.125 $X2=0 $Y2=0
cc_1157 N_A_2067_74#_c_1696_n N_A_2277_455#_c_2317_n 0.0118748f $X=11.985
+ $Y=2.485 $X2=0 $Y2=0
cc_1158 N_A_2067_74#_c_1695_n N_A_2277_455#_c_2318_n 0.00513377f $X=11.82
+ $Y=2.125 $X2=0 $Y2=0
cc_1159 N_A_2067_74#_c_1696_n N_A_2277_455#_c_2318_n 0.0313337f $X=11.985
+ $Y=2.485 $X2=0 $Y2=0
cc_1160 N_A_2067_74#_c_1697_n N_A_2277_455#_c_2318_n 6.30153e-19 $X=13.31
+ $Y=2.225 $X2=0 $Y2=0
cc_1161 N_A_2067_74#_c_1701_n N_A_2277_455#_c_2318_n 0.0049692f $X=12.105
+ $Y=2.125 $X2=0 $Y2=0
cc_1162 N_A_2067_74#_c_1696_n N_A_2277_455#_c_2320_n 0.0143942f $X=11.985
+ $Y=2.485 $X2=0 $Y2=0
cc_1163 N_A_2067_74#_c_1697_n N_A_2277_455#_c_2320_n 0.0231608f $X=13.31
+ $Y=2.225 $X2=0 $Y2=0
cc_1164 N_A_2067_74#_M1004_g N_Q_N_c_2349_n 0.0264909f $X=14.795 $Y=2.4 $X2=0
+ $Y2=0
cc_1165 N_A_2067_74#_c_1673_n N_Q_N_c_2349_n 0.00477651f $X=15.155 $Y=1.375
+ $X2=0 $Y2=0
cc_1166 N_A_2067_74#_M1029_g N_Q_N_c_2349_n 0.0101354f $X=15.245 $Y=2.4 $X2=0
+ $Y2=0
cc_1167 N_A_2067_74#_c_1680_n N_Q_N_c_2349_n 0.00114549f $X=14.795 $Y=1.375
+ $X2=0 $Y2=0
cc_1168 N_A_2067_74#_M1023_g N_Q_N_c_2350_n 0.0183249f $X=14.78 $Y=0.74 $X2=0
+ $Y2=0
cc_1169 N_A_2067_74#_M1025_g N_Q_N_c_2350_n 0.0165206f $X=15.23 $Y=0.74 $X2=0
+ $Y2=0
cc_1170 N_A_2067_74#_M1023_g Q_N 0.00250547f $X=14.78 $Y=0.74 $X2=0 $Y2=0
cc_1171 N_A_2067_74#_c_1673_n Q_N 0.00824205f $X=15.155 $Y=1.375 $X2=0 $Y2=0
cc_1172 N_A_2067_74#_M1025_g Q_N 0.00308648f $X=15.23 $Y=0.74 $X2=0 $Y2=0
cc_1173 N_A_2067_74#_c_1680_n Q_N 0.0032858f $X=14.795 $Y=1.375 $X2=0 $Y2=0
cc_1174 N_A_2067_74#_c_1681_n Q_N 0.00811537f $X=15.245 $Y=1.375 $X2=0 $Y2=0
cc_1175 N_A_2067_74#_M1040_g N_VGND_c_2412_n 0.0054334f $X=13.72 $Y=0.58 $X2=0
+ $Y2=0
cc_1176 N_A_2067_74#_M1040_g N_VGND_c_2413_n 0.00358244f $X=13.72 $Y=0.58 $X2=0
+ $Y2=0
cc_1177 N_A_2067_74#_c_1670_n N_VGND_c_2413_n 0.00760021f $X=14.705 $Y=1.375
+ $X2=0 $Y2=0
cc_1178 N_A_2067_74#_M1023_g N_VGND_c_2413_n 0.00639614f $X=14.78 $Y=0.74 $X2=0
+ $Y2=0
cc_1179 N_A_2067_74#_M1025_g N_VGND_c_2414_n 0.00819758f $X=15.23 $Y=0.74 $X2=0
+ $Y2=0
cc_1180 N_A_2067_74#_c_1676_n N_VGND_c_2414_n 0.0103331f $X=16.165 $Y=1.375
+ $X2=0 $Y2=0
cc_1181 N_A_2067_74#_M1012_g N_VGND_c_2414_n 0.00377536f $X=16.27 $Y=0.79 $X2=0
+ $Y2=0
cc_1182 N_A_2067_74#_M1012_g N_VGND_c_2415_n 0.00886999f $X=16.27 $Y=0.79 $X2=0
+ $Y2=0
cc_1183 N_A_2067_74#_c_1754_n N_VGND_c_2422_n 0.0279753f $X=12.22 $Y=0.565 $X2=0
+ $Y2=0
cc_1184 N_A_2067_74#_c_1684_n N_VGND_c_2422_n 0.00610577f $X=11.55 $Y=0.565
+ $X2=0 $Y2=0
cc_1185 N_A_2067_74#_M1040_g N_VGND_c_2424_n 0.00434272f $X=13.72 $Y=0.58 $X2=0
+ $Y2=0
cc_1186 N_A_2067_74#_M1023_g N_VGND_c_2426_n 0.00456932f $X=14.78 $Y=0.74 $X2=0
+ $Y2=0
cc_1187 N_A_2067_74#_M1025_g N_VGND_c_2426_n 0.00371957f $X=15.23 $Y=0.74 $X2=0
+ $Y2=0
cc_1188 N_A_2067_74#_M1012_g N_VGND_c_2432_n 0.00485498f $X=16.27 $Y=0.79 $X2=0
+ $Y2=0
cc_1189 N_A_2067_74#_M1040_g N_VGND_c_2439_n 0.00826076f $X=13.72 $Y=0.58 $X2=0
+ $Y2=0
cc_1190 N_A_2067_74#_M1023_g N_VGND_c_2439_n 0.00894397f $X=14.78 $Y=0.74 $X2=0
+ $Y2=0
cc_1191 N_A_2067_74#_M1025_g N_VGND_c_2439_n 0.00624688f $X=15.23 $Y=0.74 $X2=0
+ $Y2=0
cc_1192 N_A_2067_74#_M1012_g N_VGND_c_2439_n 0.00514438f $X=16.27 $Y=0.79 $X2=0
+ $Y2=0
cc_1193 N_A_2067_74#_c_1683_n N_VGND_c_2439_n 0.00674927f $X=11.38 $Y=0.945
+ $X2=0 $Y2=0
cc_1194 N_A_2067_74#_c_1754_n N_VGND_c_2439_n 0.0292546f $X=12.22 $Y=0.565 $X2=0
+ $Y2=0
cc_1195 N_A_2067_74#_c_1684_n N_VGND_c_2439_n 0.00599714f $X=11.55 $Y=0.565
+ $X2=0 $Y2=0
cc_1196 N_A_2067_74#_c_1683_n N_A_1794_74#_M1039_d 0.00457257f $X=11.38 $Y=0.945
+ $X2=0 $Y2=0
cc_1197 N_A_2067_74#_c_1687_n N_A_1794_74#_c_2594_n 0.00184691f $X=10.545
+ $Y=0.81 $X2=0 $Y2=0
cc_1198 N_A_2067_74#_M1032_s N_A_1794_74#_c_2596_n 0.00250873f $X=10.335 $Y=0.37
+ $X2=0 $Y2=0
cc_1199 N_A_2067_74#_c_1683_n N_A_1794_74#_c_2596_n 0.00337267f $X=11.38
+ $Y=0.945 $X2=0 $Y2=0
cc_1200 N_A_2067_74#_c_1687_n N_A_1794_74#_c_2596_n 0.0190143f $X=10.545 $Y=0.81
+ $X2=0 $Y2=0
cc_1201 N_A_2067_74#_c_1683_n N_A_1794_74#_c_2598_n 0.02441f $X=11.38 $Y=0.945
+ $X2=0 $Y2=0
cc_1202 N_A_2067_74#_c_1684_n N_A_1794_74#_c_2598_n 0.0229927f $X=11.55 $Y=0.565
+ $X2=0 $Y2=0
cc_1203 N_A_3177_368#_c_1893_n N_VPWR_c_1965_n 0.0701151f $X=16.03 $Y=1.985
+ $X2=0 $Y2=0
cc_1204 N_A_3177_368#_M1047_g N_VPWR_c_1966_n 0.00533694f $X=16.805 $Y=2.4 $X2=0
+ $Y2=0
cc_1205 N_A_3177_368#_c_1893_n N_VPWR_c_1966_n 0.0648796f $X=16.03 $Y=1.985
+ $X2=0 $Y2=0
cc_1206 N_A_3177_368#_c_1894_n N_VPWR_c_1966_n 0.0198206f $X=16.72 $Y=1.465
+ $X2=0 $Y2=0
cc_1207 N_A_3177_368#_c_1896_n N_VPWR_c_1966_n 0.00251384f $X=17.255 $Y=1.465
+ $X2=0 $Y2=0
cc_1208 N_A_3177_368#_M1049_g N_VPWR_c_1968_n 0.00647357f $X=17.255 $Y=2.4 $X2=0
+ $Y2=0
cc_1209 N_A_3177_368#_c_1893_n N_VPWR_c_1980_n 0.00975961f $X=16.03 $Y=1.985
+ $X2=0 $Y2=0
cc_1210 N_A_3177_368#_M1047_g N_VPWR_c_1981_n 0.005209f $X=16.805 $Y=2.4 $X2=0
+ $Y2=0
cc_1211 N_A_3177_368#_M1049_g N_VPWR_c_1981_n 0.0048691f $X=17.255 $Y=2.4 $X2=0
+ $Y2=0
cc_1212 N_A_3177_368#_M1047_g N_VPWR_c_1956_n 0.00987399f $X=16.805 $Y=2.4 $X2=0
+ $Y2=0
cc_1213 N_A_3177_368#_M1049_g N_VPWR_c_1956_n 0.00875947f $X=17.255 $Y=2.4 $X2=0
+ $Y2=0
cc_1214 N_A_3177_368#_c_1893_n N_VPWR_c_1956_n 0.0111753f $X=16.03 $Y=1.985
+ $X2=0 $Y2=0
cc_1215 N_A_3177_368#_c_1892_n N_Q_N_c_2350_n 0.00502622f $X=16.055 $Y=0.615
+ $X2=0 $Y2=0
cc_1216 N_A_3177_368#_c_1895_n Q_N 0.00298092f $X=16.042 $Y=1.465 $X2=0 $Y2=0
cc_1217 N_A_3177_368#_M1047_g N_Q_c_2378_n 0.0129009f $X=16.805 $Y=2.4 $X2=0
+ $Y2=0
cc_1218 N_A_3177_368#_M1049_g N_Q_c_2378_n 0.0149161f $X=17.255 $Y=2.4 $X2=0
+ $Y2=0
cc_1219 N_A_3177_368#_M1047_g N_Q_c_2379_n 0.00320336f $X=16.805 $Y=2.4 $X2=0
+ $Y2=0
cc_1220 N_A_3177_368#_M1049_g N_Q_c_2379_n 0.00270934f $X=17.255 $Y=2.4 $X2=0
+ $Y2=0
cc_1221 N_A_3177_368#_c_1894_n N_Q_c_2379_n 0.00138666f $X=16.72 $Y=1.465 $X2=0
+ $Y2=0
cc_1222 N_A_3177_368#_c_1896_n N_Q_c_2379_n 0.00310238f $X=17.255 $Y=1.465 $X2=0
+ $Y2=0
cc_1223 N_A_3177_368#_M1047_g N_Q_c_2375_n 0.00293165f $X=16.805 $Y=2.4 $X2=0
+ $Y2=0
cc_1224 N_A_3177_368#_M1001_g N_Q_c_2375_n 0.0025553f $X=16.835 $Y=0.74 $X2=0
+ $Y2=0
cc_1225 N_A_3177_368#_M1049_g N_Q_c_2375_n 0.00994275f $X=17.255 $Y=2.4 $X2=0
+ $Y2=0
cc_1226 N_A_3177_368#_M1022_g N_Q_c_2375_n 0.00866774f $X=17.265 $Y=0.74 $X2=0
+ $Y2=0
cc_1227 N_A_3177_368#_c_1894_n N_Q_c_2375_n 0.0249855f $X=16.72 $Y=1.465 $X2=0
+ $Y2=0
cc_1228 N_A_3177_368#_c_1896_n N_Q_c_2375_n 0.0238044f $X=17.255 $Y=1.465 $X2=0
+ $Y2=0
cc_1229 N_A_3177_368#_M1001_g Q 0.00761048f $X=16.835 $Y=0.74 $X2=0 $Y2=0
cc_1230 N_A_3177_368#_M1022_g Q 0.0081896f $X=17.265 $Y=0.74 $X2=0 $Y2=0
cc_1231 N_A_3177_368#_M1001_g Q 0.00326771f $X=16.835 $Y=0.74 $X2=0 $Y2=0
cc_1232 N_A_3177_368#_M1022_g Q 0.00215589f $X=17.265 $Y=0.74 $X2=0 $Y2=0
cc_1233 N_A_3177_368#_c_1896_n Q 0.00244427f $X=17.255 $Y=1.465 $X2=0 $Y2=0
cc_1234 N_A_3177_368#_c_1892_n N_VGND_c_2414_n 0.048096f $X=16.055 $Y=0.615
+ $X2=0 $Y2=0
cc_1235 N_A_3177_368#_M1001_g N_VGND_c_2415_n 0.00501537f $X=16.835 $Y=0.74
+ $X2=0 $Y2=0
cc_1236 N_A_3177_368#_c_1892_n N_VGND_c_2415_n 0.0405787f $X=16.055 $Y=0.615
+ $X2=0 $Y2=0
cc_1237 N_A_3177_368#_c_1894_n N_VGND_c_2415_n 0.0213234f $X=16.72 $Y=1.465
+ $X2=0 $Y2=0
cc_1238 N_A_3177_368#_c_1896_n N_VGND_c_2415_n 0.00347105f $X=17.255 $Y=1.465
+ $X2=0 $Y2=0
cc_1239 N_A_3177_368#_M1022_g N_VGND_c_2417_n 0.00646793f $X=17.265 $Y=0.74
+ $X2=0 $Y2=0
cc_1240 N_A_3177_368#_c_1892_n N_VGND_c_2432_n 0.0111427f $X=16.055 $Y=0.615
+ $X2=0 $Y2=0
cc_1241 N_A_3177_368#_M1001_g N_VGND_c_2433_n 0.00434272f $X=16.835 $Y=0.74
+ $X2=0 $Y2=0
cc_1242 N_A_3177_368#_M1022_g N_VGND_c_2433_n 0.00422942f $X=17.265 $Y=0.74
+ $X2=0 $Y2=0
cc_1243 N_A_3177_368#_M1001_g N_VGND_c_2439_n 0.00825283f $X=16.835 $Y=0.74
+ $X2=0 $Y2=0
cc_1244 N_A_3177_368#_M1022_g N_VGND_c_2439_n 0.00787255f $X=17.265 $Y=0.74
+ $X2=0 $Y2=0
cc_1245 N_A_3177_368#_c_1892_n N_VGND_c_2439_n 0.0122012f $X=16.055 $Y=0.615
+ $X2=0 $Y2=0
cc_1246 N_VPWR_c_1956_n N_A_307_74#_c_2157_n 0.0155167f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1247 N_VPWR_M1041_d N_A_307_74#_c_2159_n 0.0030394f $X=2.525 $Y=2.32 $X2=0
+ $Y2=0
cc_1248 N_VPWR_M1036_d N_A_307_74#_c_2159_n 0.00307632f $X=3.555 $Y=1.84 $X2=0
+ $Y2=0
cc_1249 N_VPWR_c_1958_n N_A_307_74#_c_2159_n 0.0166684f $X=2.67 $Y=2.815 $X2=0
+ $Y2=0
cc_1250 N_VPWR_c_1985_n N_A_307_74#_c_2159_n 0.010348f $X=4.22 $Y=3.032 $X2=0
+ $Y2=0
cc_1251 N_VPWR_c_1956_n N_A_307_74#_c_2159_n 0.0234956f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1252 N_VPWR_M1036_d N_A_307_74#_c_2160_n 0.00836317f $X=3.555 $Y=1.84 $X2=0
+ $Y2=0
cc_1253 N_VPWR_c_1985_n N_A_307_74#_c_2160_n 0.0131433f $X=4.22 $Y=3.032 $X2=0
+ $Y2=0
cc_1254 N_VPWR_c_1957_n N_A_307_74#_c_2161_n 0.0201193f $X=0.8 $Y=2.475 $X2=0
+ $Y2=0
cc_1255 N_VPWR_c_1958_n N_A_307_74#_c_2161_n 0.00987247f $X=2.67 $Y=2.815 $X2=0
+ $Y2=0
cc_1256 N_VPWR_c_1978_n N_A_307_74#_c_2161_n 0.0197955f $X=2.495 $Y=3.33 $X2=0
+ $Y2=0
cc_1257 N_VPWR_c_1956_n N_A_307_74#_c_2161_n 0.016258f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1258 N_VPWR_M1041_d N_A_307_74#_c_2195_n 5.78969e-19 $X=2.525 $Y=2.32 $X2=0
+ $Y2=0
cc_1259 N_VPWR_c_1958_n N_A_307_74#_c_2195_n 0.0070234f $X=2.67 $Y=2.815 $X2=0
+ $Y2=0
cc_1260 N_VPWR_c_1956_n N_A_307_74#_c_2195_n 0.00144544f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1261 N_VPWR_M1036_d N_A_307_74#_c_2197_n 0.0116196f $X=3.555 $Y=1.84 $X2=0
+ $Y2=0
cc_1262 N_VPWR_c_1985_n N_A_307_74#_c_2197_n 0.0140504f $X=4.22 $Y=3.032 $X2=0
+ $Y2=0
cc_1263 N_VPWR_c_1956_n N_A_307_74#_c_2197_n 5.67209e-19 $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1264 N_VPWR_M1003_s N_A_1789_424#_c_2275_n 0.00357451f $X=9.455 $Y=2.12 $X2=0
+ $Y2=0
cc_1265 N_VPWR_c_1962_n N_A_1789_424#_c_2275_n 0.014901f $X=9.59 $Y=2.725 $X2=0
+ $Y2=0
cc_1266 N_VPWR_c_1971_n N_A_1789_424#_c_2270_n 0.0644458f $X=12.94 $Y=3.33 $X2=0
+ $Y2=0
cc_1267 N_VPWR_c_1956_n N_A_1789_424#_c_2270_n 0.0356291f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1268 N_VPWR_c_1962_n N_A_1789_424#_c_2271_n 0.0103534f $X=9.59 $Y=2.725 $X2=0
+ $Y2=0
cc_1269 N_VPWR_c_1971_n N_A_1789_424#_c_2271_n 0.0178163f $X=12.94 $Y=3.33 $X2=0
+ $Y2=0
cc_1270 N_VPWR_c_1956_n N_A_1789_424#_c_2271_n 0.00958215f $X=17.52 $Y=3.33
+ $X2=0 $Y2=0
cc_1271 N_VPWR_c_1961_n N_A_1789_424#_c_2273_n 0.0364847f $X=8.5 $Y=2.57 $X2=0
+ $Y2=0
cc_1272 N_VPWR_c_1962_n N_A_1789_424#_c_2273_n 0.0191298f $X=9.59 $Y=2.725 $X2=0
+ $Y2=0
cc_1273 N_VPWR_c_1969_n N_A_1789_424#_c_2273_n 0.0146357f $X=9.425 $Y=3.33 $X2=0
+ $Y2=0
cc_1274 N_VPWR_c_1956_n N_A_1789_424#_c_2273_n 0.0121141f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1275 N_VPWR_c_1963_n N_A_2277_455#_c_2318_n 0.0094484f $X=13.025 $Y=2.75
+ $X2=0 $Y2=0
cc_1276 N_VPWR_c_1971_n N_A_2277_455#_c_2318_n 0.0652834f $X=12.94 $Y=3.33 $X2=0
+ $Y2=0
cc_1277 N_VPWR_c_1956_n N_A_2277_455#_c_2318_n 0.0387639f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1278 N_VPWR_c_1971_n N_A_2277_455#_c_2319_n 0.0162012f $X=12.94 $Y=3.33 $X2=0
+ $Y2=0
cc_1279 N_VPWR_c_1956_n N_A_2277_455#_c_2319_n 0.00879606f $X=17.52 $Y=3.33
+ $X2=0 $Y2=0
cc_1280 N_VPWR_c_1963_n N_A_2277_455#_c_2320_n 0.0126297f $X=13.025 $Y=2.75
+ $X2=0 $Y2=0
cc_1281 N_VPWR_c_1964_n N_Q_N_c_2349_n 0.0387846f $X=14.57 $Y=1.985 $X2=0 $Y2=0
cc_1282 N_VPWR_c_1965_n N_Q_N_c_2349_n 0.0395727f $X=15.47 $Y=1.985 $X2=0 $Y2=0
cc_1283 N_VPWR_c_1975_n N_Q_N_c_2349_n 0.0111875f $X=15.305 $Y=3.33 $X2=0 $Y2=0
cc_1284 N_VPWR_c_1956_n N_Q_N_c_2349_n 0.00918014f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1285 N_VPWR_c_1981_n N_Q_c_2378_n 0.0157112f $X=17.395 $Y=3.33 $X2=0 $Y2=0
cc_1286 N_VPWR_c_1956_n N_Q_c_2378_n 0.0127977f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1287 N_VPWR_c_1966_n N_Q_c_2379_n 0.0400476f $X=16.58 $Y=1.985 $X2=0 $Y2=0
cc_1288 N_VPWR_c_1968_n N_Q_c_2379_n 0.0455874f $X=17.48 $Y=1.985 $X2=0 $Y2=0
cc_1289 N_A_307_74#_c_2157_n A_421_464# 0.00255471f $X=2.465 $Y=2.395 $X2=-0.19
+ $Y2=-0.245
cc_1290 N_A_307_74#_c_2154_n N_VGND_c_2407_n 0.00316404f $X=2.55 $Y=2.31 $X2=0
+ $Y2=0
cc_1291 N_A_307_74#_c_2177_n N_VGND_c_2407_n 0.0172749f $X=2.155 $Y=0.565 $X2=0
+ $Y2=0
cc_1292 N_A_307_74#_c_2177_n N_VGND_c_2418_n 0.0178113f $X=2.155 $Y=0.565 $X2=0
+ $Y2=0
cc_1293 N_A_307_74#_c_2177_n N_VGND_c_2439_n 0.0216127f $X=2.155 $Y=0.565 $X2=0
+ $Y2=0
cc_1294 N_A_307_74#_c_2154_n A_495_74# 5.40786e-19 $X=2.55 $Y=2.31 $X2=-0.19
+ $Y2=-0.245
cc_1295 N_A_307_74#_c_2177_n A_495_74# 0.00326443f $X=2.155 $Y=0.565 $X2=-0.19
+ $Y2=-0.245
cc_1296 N_A_1789_424#_c_2272_n N_A_2277_455#_c_2317_n 0.0302976f $X=10.94
+ $Y=2.465 $X2=0 $Y2=0
cc_1297 N_A_1789_424#_c_2270_n N_A_2277_455#_c_2319_n 0.0104058f $X=10.775
+ $Y=2.99 $X2=0 $Y2=0
cc_1298 N_A_1789_424#_c_2272_n N_A_2277_455#_c_2319_n 0.0012809f $X=10.94
+ $Y=2.465 $X2=0 $Y2=0
cc_1299 N_Q_N_c_2350_n N_VGND_c_2413_n 0.0176944f $X=15.015 $Y=0.515 $X2=0 $Y2=0
cc_1300 N_Q_N_c_2350_n N_VGND_c_2414_n 0.0600324f $X=15.015 $Y=0.515 $X2=0 $Y2=0
cc_1301 N_Q_N_c_2350_n N_VGND_c_2426_n 0.0168417f $X=15.015 $Y=0.515 $X2=0 $Y2=0
cc_1302 N_Q_N_c_2350_n N_VGND_c_2439_n 0.0137451f $X=15.015 $Y=0.515 $X2=0 $Y2=0
cc_1303 Q N_VGND_c_2415_n 0.0295042f $X=16.955 $Y=0.47 $X2=0 $Y2=0
cc_1304 Q N_VGND_c_2417_n 0.0308798f $X=16.955 $Y=0.47 $X2=0 $Y2=0
cc_1305 Q N_VGND_c_2433_n 0.0149085f $X=16.955 $Y=0.47 $X2=0 $Y2=0
cc_1306 Q N_VGND_c_2439_n 0.0122037f $X=16.955 $Y=0.47 $X2=0 $Y2=0
cc_1307 N_VGND_c_2410_n N_A_1794_74#_c_2593_n 0.0117303f $X=8.365 $Y=0.515 $X2=0
+ $Y2=0
cc_1308 N_VGND_c_2411_n N_A_1794_74#_c_2593_n 0.0189563f $X=9.615 $Y=0.59 $X2=0
+ $Y2=0
cc_1309 N_VGND_c_2420_n N_A_1794_74#_c_2593_n 0.011066f $X=9.45 $Y=0 $X2=0 $Y2=0
cc_1310 N_VGND_c_2439_n N_A_1794_74#_c_2593_n 0.00915947f $X=17.52 $Y=0 $X2=0
+ $Y2=0
cc_1311 N_VGND_M1005_d N_A_1794_74#_c_2594_n 0.00197722f $X=9.455 $Y=0.37 $X2=0
+ $Y2=0
cc_1312 N_VGND_c_2411_n N_A_1794_74#_c_2594_n 0.0172656f $X=9.615 $Y=0.59 $X2=0
+ $Y2=0
cc_1313 N_VGND_c_2422_n N_A_1794_74#_c_2596_n 0.0423335f $X=13.26 $Y=0 $X2=0
+ $Y2=0
cc_1314 N_VGND_c_2439_n N_A_1794_74#_c_2596_n 0.0239357f $X=17.52 $Y=0 $X2=0
+ $Y2=0
cc_1315 N_VGND_c_2411_n N_A_1794_74#_c_2597_n 0.0112234f $X=9.615 $Y=0.59 $X2=0
+ $Y2=0
cc_1316 N_VGND_c_2422_n N_A_1794_74#_c_2597_n 0.0178338f $X=13.26 $Y=0 $X2=0
+ $Y2=0
cc_1317 N_VGND_c_2439_n N_A_1794_74#_c_2597_n 0.00960503f $X=17.52 $Y=0 $X2=0
+ $Y2=0
cc_1318 N_VGND_c_2422_n N_A_1794_74#_c_2598_n 0.0227418f $X=13.26 $Y=0 $X2=0
+ $Y2=0
cc_1319 N_VGND_c_2439_n N_A_1794_74#_c_2598_n 0.0126077f $X=17.52 $Y=0 $X2=0
+ $Y2=0

* NGSPICE file created from sky130_fd_sc_ms__clkbuf_4.ext - technology: sky130A

.subckt sky130_fd_sc_ms__clkbuf_4 A VGND VNB VPB VPWR X
M1000 VGND a_83_270# X VNB nlowvt w=420000u l=150000u
+  ad=3.969e+11p pd=4.41e+06u as=2.52e+11p ps=2.88e+06u
M1001 X a_83_270# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=9.744e+11p ps=8.46e+06u
M1002 VPWR a_83_270# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_83_270# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_83_270# A VGND VNB nlowvt w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1005 a_83_270# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1006 VPWR a_83_270# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_83_270# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_83_270# VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_83_270# X VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


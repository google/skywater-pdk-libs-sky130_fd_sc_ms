# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__a21bo_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.725000 1.260000 3.235000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.450000 3.735000 1.780000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.208000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.510000 1.550000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.543200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.020000 0.840000 1.395000 1.040000 ;
        RECT 1.020000 1.040000 1.190000 1.820000 ;
        RECT 1.020000 1.820000 1.415000 2.070000 ;
        RECT 1.225000 0.350000 1.565000 0.750000 ;
        RECT 1.225000 0.750000 1.395000 0.840000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.120000  1.820000 0.450000 2.240000 ;
      RECT 0.120000  2.240000 1.810000 2.410000 ;
      RECT 0.120000  2.410000 0.450000 2.700000 ;
      RECT 0.270000  0.540000 0.600000 0.840000 ;
      RECT 0.270000  0.840000 0.850000 1.010000 ;
      RECT 0.635000  2.580000 0.965000 3.245000 ;
      RECT 0.680000  1.010000 0.850000 2.240000 ;
      RECT 0.805000  0.085000 1.055000 0.670000 ;
      RECT 1.360000  1.220000 1.735000 1.550000 ;
      RECT 1.535000  2.580000 1.865000 3.245000 ;
      RECT 1.565000  0.920000 2.810000 1.090000 ;
      RECT 1.565000  1.090000 1.735000 1.220000 ;
      RECT 1.605000  1.720000 2.075000 1.890000 ;
      RECT 1.605000  1.890000 1.810000 2.240000 ;
      RECT 1.735000  0.085000 2.310000 0.750000 ;
      RECT 1.905000  1.260000 2.215000 1.590000 ;
      RECT 1.905000  1.590000 2.075000 1.720000 ;
      RECT 2.055000  2.060000 2.415000 2.980000 ;
      RECT 2.245000  1.760000 2.555000 1.930000 ;
      RECT 2.245000  1.930000 2.415000 2.060000 ;
      RECT 2.385000  1.090000 2.555000 1.760000 ;
      RECT 2.480000  0.350000 2.810000 0.920000 ;
      RECT 2.585000  2.100000 3.735000 2.270000 ;
      RECT 2.585000  2.270000 2.755000 2.980000 ;
      RECT 2.955000  2.440000 3.205000 3.245000 ;
      RECT 3.380000  0.085000 3.710000 1.090000 ;
      RECT 3.405000  1.950000 3.735000 2.100000 ;
      RECT 3.405000  2.270000 3.735000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_ms__a21bo_2

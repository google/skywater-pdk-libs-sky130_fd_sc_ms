* File: sky130_fd_sc_ms__a21o_1.pxi.spice
* Created: Fri Aug 28 16:59:05 2020
* 
x_PM_SKY130_FD_SC_MS__A21O_1%A_81_264# N_A_81_264#_M1003_d N_A_81_264#_M1006_s
+ N_A_81_264#_M1005_g N_A_81_264#_c_63_n N_A_81_264#_c_64_n N_A_81_264#_M1000_g
+ N_A_81_264#_c_65_n N_A_81_264#_c_70_n N_A_81_264#_c_76_p N_A_81_264#_c_66_n
+ N_A_81_264#_c_67_n N_A_81_264#_c_71_n N_A_81_264#_c_72_n N_A_81_264#_c_68_n
+ PM_SKY130_FD_SC_MS__A21O_1%A_81_264#
x_PM_SKY130_FD_SC_MS__A21O_1%B1 N_B1_M1006_g N_B1_M1003_g B1 N_B1_c_129_n
+ PM_SKY130_FD_SC_MS__A21O_1%B1
x_PM_SKY130_FD_SC_MS__A21O_1%A1 N_A1_M1007_g N_A1_M1004_g A1 N_A1_c_164_n
+ PM_SKY130_FD_SC_MS__A21O_1%A1
x_PM_SKY130_FD_SC_MS__A21O_1%A2 N_A2_M1001_g N_A2_c_200_n N_A2_M1002_g
+ N_A2_c_202_n A2 N_A2_c_204_n PM_SKY130_FD_SC_MS__A21O_1%A2
x_PM_SKY130_FD_SC_MS__A21O_1%X N_X_M1000_s N_X_M1005_s N_X_c_233_n N_X_c_234_n
+ N_X_c_235_n X X X X N_X_c_236_n PM_SKY130_FD_SC_MS__A21O_1%X
x_PM_SKY130_FD_SC_MS__A21O_1%VPWR N_VPWR_M1005_d N_VPWR_M1007_d N_VPWR_c_254_n
+ N_VPWR_c_255_n N_VPWR_c_256_n N_VPWR_c_257_n VPWR N_VPWR_c_258_n
+ N_VPWR_c_259_n N_VPWR_c_253_n N_VPWR_c_261_n PM_SKY130_FD_SC_MS__A21O_1%VPWR
x_PM_SKY130_FD_SC_MS__A21O_1%A_367_392# N_A_367_392#_M1006_d
+ N_A_367_392#_M1002_d N_A_367_392#_c_290_n N_A_367_392#_c_291_n
+ N_A_367_392#_c_292_n N_A_367_392#_c_293_n N_A_367_392#_c_294_n
+ PM_SKY130_FD_SC_MS__A21O_1%A_367_392#
x_PM_SKY130_FD_SC_MS__A21O_1%VGND N_VGND_M1000_d N_VGND_M1001_d N_VGND_c_323_n
+ N_VGND_c_324_n N_VGND_c_357_n N_VGND_c_349_n N_VGND_c_325_n N_VGND_c_326_n
+ N_VGND_c_327_n N_VGND_c_328_n N_VGND_c_329_n VGND N_VGND_c_330_n
+ N_VGND_c_331_n PM_SKY130_FD_SC_MS__A21O_1%VGND
cc_1 VNB N_A_81_264#_M1005_g 6.61219e-19 $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_2 VNB N_A_81_264#_c_63_n 0.03594f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.47
cc_3 VNB N_A_81_264#_c_64_n 0.0196825f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.395
cc_4 VNB N_A_81_264#_c_65_n 0.0196318f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=1.485
cc_5 VNB N_A_81_264#_c_66_n 0.00381609f $X=-0.19 $Y=-0.245 $X2=1.97 $Y2=0.805
cc_6 VNB N_A_81_264#_c_67_n 0.00278456f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.38
cc_7 VNB N_A_81_264#_c_68_n 0.0389821f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=1.485
cc_8 VNB N_B1_M1003_g 0.0197271f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.65
cc_9 VNB B1 8.71858e-19 $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_10 VNB N_B1_c_129_n 0.0197423f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=1.47
cc_11 VNB N_A1_M1004_g 0.0191344f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.65
cc_12 VNB A1 0.0032213f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_13 VNB N_A1_c_164_n 0.0194421f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=1.47
cc_14 VNB N_A2_M1001_g 0.012615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_c_200_n 0.00850929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A2_M1002_g 0.0145107f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.65
cc_17 VNB N_A2_c_202_n 0.050643f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.395
cc_18 VNB A2 0.0277287f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.95
cc_19 VNB N_A2_c_204_n 5.28587e-19 $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.95
cc_20 VNB N_X_c_233_n 0.0282147f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_21 VNB N_X_c_234_n 0.0149129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_X_c_235_n 0.0121113f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.395
cc_23 VNB N_X_c_236_n 0.0283248f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.38
cc_24 VNB N_VPWR_c_253_n 0.143779f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.95
cc_25 VNB N_VGND_c_323_n 0.0280514f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_26 VNB N_VGND_c_324_n 0.0219582f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=1.47
cc_27 VNB N_VGND_c_325_n 0.0410501f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=1.485
cc_28 VNB N_VGND_c_326_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.485
cc_29 VNB N_VGND_c_327_n 0.0214589f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.485
cc_30 VNB N_VGND_c_328_n 0.00326658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_329_n 0.0245056f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=1.65
cc_32 VNB N_VGND_c_330_n 0.0245652f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.485
cc_33 VNB N_VGND_c_331_n 0.243932f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=1.485
cc_34 VPB N_A_81_264#_M1005_g 0.0303398f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_35 VPB N_A_81_264#_c_70_n 0.0167165f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=2.815
cc_36 VPB N_A_81_264#_c_71_n 0.00509728f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=2.115
cc_37 VPB N_A_81_264#_c_72_n 0.00738973f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.95
cc_38 VPB N_B1_M1006_g 0.0274882f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB B1 0.00206873f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_40 VPB N_B1_c_129_n 0.0129182f $X=-0.19 $Y=1.66 $X2=0.755 $Y2=1.47
cc_41 VPB N_A1_M1007_g 0.0236294f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB A1 0.00137164f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_43 VPB N_A1_c_164_n 0.0124339f $X=-0.19 $Y=1.66 $X2=0.755 $Y2=1.47
cc_44 VPB N_A2_M1002_g 0.0420646f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.65
cc_45 VPB X 0.00928864f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=0.95
cc_46 VPB X 0.0418804f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=2.815
cc_47 VPB N_X_c_236_n 0.00778611f $X=-0.19 $Y=1.66 $X2=1.33 $Y2=1.38
cc_48 VPB N_VPWR_c_254_n 0.0294637f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_49 VPB N_VPWR_c_255_n 0.00833138f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=0.95
cc_50 VPB N_VPWR_c_256_n 0.0407193f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.485
cc_51 VPB N_VPWR_c_257_n 0.00382106f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.485
cc_52 VPB N_VPWR_c_258_n 0.0196317f $X=-0.19 $Y=1.66 $X2=1.33 $Y2=1.95
cc_53 VPB N_VPWR_c_259_n 0.0258341f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=2.115
cc_54 VPB N_VPWR_c_253_n 0.0846155f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.95
cc_55 VPB N_VPWR_c_261_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.485
cc_56 VPB N_A_367_392#_c_290_n 0.00401924f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.65
cc_57 VPB N_A_367_392#_c_291_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_58 VPB N_A_367_392#_c_292_n 0.00778237f $X=-0.19 $Y=1.66 $X2=1.13 $Y2=1.47
cc_59 VPB N_A_367_392#_c_293_n 0.0131653f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=1.395
cc_60 VPB N_A_367_392#_c_294_n 0.0358769f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=0.95
cc_61 N_A_81_264#_c_71_n N_B1_M1006_g 7.1053e-19 $X=1.52 $Y=2.115 $X2=0 $Y2=0
cc_62 N_A_81_264#_c_72_n N_B1_M1006_g 0.00547941f $X=1.425 $Y=1.95 $X2=0 $Y2=0
cc_63 N_A_81_264#_c_64_n N_B1_M1003_g 0.0176258f $X=1.205 $Y=1.395 $X2=0 $Y2=0
cc_64 N_A_81_264#_c_76_p N_B1_M1003_g 0.0121724f $X=1.805 $Y=1.195 $X2=0 $Y2=0
cc_65 N_A_81_264#_c_66_n N_B1_M1003_g 0.00723827f $X=1.97 $Y=0.805 $X2=0 $Y2=0
cc_66 N_A_81_264#_c_67_n N_B1_M1003_g 0.00411569f $X=1.33 $Y=1.38 $X2=0 $Y2=0
cc_67 N_A_81_264#_c_76_p B1 0.0159378f $X=1.805 $Y=1.195 $X2=0 $Y2=0
cc_68 N_A_81_264#_c_67_n B1 0.0165507f $X=1.33 $Y=1.38 $X2=0 $Y2=0
cc_69 N_A_81_264#_c_71_n B1 0.00152541f $X=1.52 $Y=2.115 $X2=0 $Y2=0
cc_70 N_A_81_264#_c_72_n B1 0.00952856f $X=1.425 $Y=1.95 $X2=0 $Y2=0
cc_71 N_A_81_264#_c_63_n N_B1_c_129_n 0.00540357f $X=1.13 $Y=1.47 $X2=0 $Y2=0
cc_72 N_A_81_264#_c_76_p N_B1_c_129_n 0.00275021f $X=1.805 $Y=1.195 $X2=0 $Y2=0
cc_73 N_A_81_264#_c_67_n N_B1_c_129_n 0.00340356f $X=1.33 $Y=1.38 $X2=0 $Y2=0
cc_74 N_A_81_264#_c_71_n N_B1_c_129_n 0.00258674f $X=1.52 $Y=2.115 $X2=0 $Y2=0
cc_75 N_A_81_264#_c_72_n N_B1_c_129_n 0.00320156f $X=1.425 $Y=1.95 $X2=0 $Y2=0
cc_76 N_A_81_264#_c_76_p N_A1_M1004_g 0.00346932f $X=1.805 $Y=1.195 $X2=0 $Y2=0
cc_77 N_A_81_264#_c_66_n N_A1_M1004_g 0.00599966f $X=1.97 $Y=0.805 $X2=0 $Y2=0
cc_78 N_A_81_264#_c_76_p A1 0.00468798f $X=1.805 $Y=1.195 $X2=0 $Y2=0
cc_79 N_A_81_264#_c_76_p N_A1_c_164_n 3.32624e-19 $X=1.805 $Y=1.195 $X2=0 $Y2=0
cc_80 N_A_81_264#_c_76_p N_A2_M1001_g 5.14251e-19 $X=1.805 $Y=1.195 $X2=0 $Y2=0
cc_81 N_A_81_264#_c_66_n N_A2_M1001_g 4.72693e-19 $X=1.97 $Y=0.805 $X2=0 $Y2=0
cc_82 N_A_81_264#_c_63_n N_X_c_233_n 0.00199362f $X=1.13 $Y=1.47 $X2=0 $Y2=0
cc_83 N_A_81_264#_c_65_n N_X_c_233_n 0.0514037f $X=1.245 $Y=1.485 $X2=0 $Y2=0
cc_84 N_A_81_264#_c_68_n N_X_c_233_n 0.0086547f $X=0.755 $Y=1.485 $X2=0 $Y2=0
cc_85 N_A_81_264#_M1005_g X 0.00322931f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_86 N_A_81_264#_c_65_n X 7.18422e-19 $X=1.245 $Y=1.485 $X2=0 $Y2=0
cc_87 N_A_81_264#_M1005_g X 0.0140232f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_88 N_A_81_264#_c_65_n N_X_c_236_n 0.0262118f $X=1.245 $Y=1.485 $X2=0 $Y2=0
cc_89 N_A_81_264#_c_68_n N_X_c_236_n 0.014292f $X=0.755 $Y=1.485 $X2=0 $Y2=0
cc_90 N_A_81_264#_M1005_g N_VPWR_c_254_n 0.00649215f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_91 N_A_81_264#_c_63_n N_VPWR_c_254_n 7.91918e-19 $X=1.13 $Y=1.47 $X2=0 $Y2=0
cc_92 N_A_81_264#_c_65_n N_VPWR_c_254_n 0.0214461f $X=1.245 $Y=1.485 $X2=0 $Y2=0
cc_93 N_A_81_264#_c_72_n N_VPWR_c_254_n 0.056301f $X=1.425 $Y=1.95 $X2=0 $Y2=0
cc_94 N_A_81_264#_c_68_n N_VPWR_c_254_n 0.00277218f $X=0.755 $Y=1.485 $X2=0
+ $Y2=0
cc_95 N_A_81_264#_c_70_n N_VPWR_c_256_n 0.0159743f $X=1.52 $Y=2.815 $X2=0 $Y2=0
cc_96 N_A_81_264#_M1005_g N_VPWR_c_258_n 0.005209f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_97 N_A_81_264#_M1005_g N_VPWR_c_253_n 0.00991105f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_98 N_A_81_264#_c_70_n N_VPWR_c_253_n 0.0132221f $X=1.52 $Y=2.815 $X2=0 $Y2=0
cc_99 N_A_81_264#_c_76_p N_A_367_392#_c_290_n 0.00628319f $X=1.805 $Y=1.195
+ $X2=0 $Y2=0
cc_100 N_A_81_264#_c_71_n N_A_367_392#_c_290_n 0.00662256f $X=1.52 $Y=2.115
+ $X2=0 $Y2=0
cc_101 N_A_81_264#_c_70_n N_A_367_392#_c_291_n 0.0290144f $X=1.52 $Y=2.815 $X2=0
+ $Y2=0
cc_102 N_A_81_264#_c_76_p N_VGND_M1000_d 0.00682387f $X=1.805 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_103 N_A_81_264#_c_67_n N_VGND_M1000_d 0.00136247f $X=1.33 $Y=1.38 $X2=-0.19
+ $Y2=-0.245
cc_104 N_A_81_264#_c_64_n N_VGND_c_323_n 0.0157678f $X=1.205 $Y=1.395 $X2=0
+ $Y2=0
cc_105 N_A_81_264#_c_76_p N_VGND_c_323_n 0.0137131f $X=1.805 $Y=1.195 $X2=0
+ $Y2=0
cc_106 N_A_81_264#_c_66_n N_VGND_c_323_n 0.0178602f $X=1.97 $Y=0.805 $X2=0 $Y2=0
cc_107 N_A_81_264#_c_67_n N_VGND_c_323_n 0.00902191f $X=1.33 $Y=1.38 $X2=0 $Y2=0
cc_108 N_A_81_264#_c_66_n N_VGND_c_324_n 0.00746887f $X=1.97 $Y=0.805 $X2=0
+ $Y2=0
cc_109 N_A_81_264#_c_64_n N_VGND_c_325_n 0.00365567f $X=1.205 $Y=1.395 $X2=0
+ $Y2=0
cc_110 N_A_81_264#_c_66_n N_VGND_c_327_n 0.00615803f $X=1.97 $Y=0.805 $X2=0
+ $Y2=0
cc_111 N_A_81_264#_c_76_p N_VGND_c_329_n 0.00495397f $X=1.805 $Y=1.195 $X2=0
+ $Y2=0
cc_112 N_A_81_264#_c_66_n N_VGND_c_329_n 0.00276199f $X=1.97 $Y=0.805 $X2=0
+ $Y2=0
cc_113 N_A_81_264#_c_64_n N_VGND_c_331_n 0.00404919f $X=1.205 $Y=1.395 $X2=0
+ $Y2=0
cc_114 N_A_81_264#_c_66_n N_VGND_c_331_n 0.00967008f $X=1.97 $Y=0.805 $X2=0
+ $Y2=0
cc_115 N_B1_M1006_g N_A1_M1007_g 0.0155445f $X=1.745 $Y=2.46 $X2=0 $Y2=0
cc_116 N_B1_M1003_g N_A1_M1004_g 0.0117284f $X=1.755 $Y=1 $X2=0 $Y2=0
cc_117 B1 A1 0.0204777f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_118 N_B1_c_129_n A1 0.00114936f $X=1.67 $Y=1.615 $X2=0 $Y2=0
cc_119 B1 N_A1_c_164_n 0.00115083f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_120 N_B1_c_129_n N_A1_c_164_n 0.0201104f $X=1.67 $Y=1.615 $X2=0 $Y2=0
cc_121 N_B1_M1006_g N_VPWR_c_256_n 0.005209f $X=1.745 $Y=2.46 $X2=0 $Y2=0
cc_122 N_B1_M1006_g N_VPWR_c_253_n 0.00988607f $X=1.745 $Y=2.46 $X2=0 $Y2=0
cc_123 N_B1_M1006_g N_A_367_392#_c_290_n 0.00265845f $X=1.745 $Y=2.46 $X2=0
+ $Y2=0
cc_124 B1 N_A_367_392#_c_290_n 0.00232699f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_125 N_B1_M1006_g N_A_367_392#_c_291_n 0.0112601f $X=1.745 $Y=2.46 $X2=0 $Y2=0
cc_126 N_B1_M1003_g N_VGND_c_323_n 0.00552238f $X=1.755 $Y=1 $X2=0 $Y2=0
cc_127 N_B1_M1003_g N_VGND_c_327_n 0.0037378f $X=1.755 $Y=1 $X2=0 $Y2=0
cc_128 N_B1_M1003_g N_VGND_c_331_n 0.00454494f $X=1.755 $Y=1 $X2=0 $Y2=0
cc_129 A1 N_A2_c_200_n 0.00223091f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_130 N_A1_c_164_n N_A2_c_200_n 0.0214073f $X=2.21 $Y=1.615 $X2=0 $Y2=0
cc_131 N_A1_M1007_g N_A2_M1002_g 0.0250263f $X=2.195 $Y=2.46 $X2=0 $Y2=0
cc_132 N_A1_M1004_g N_A2_c_202_n 0.0301488f $X=2.185 $Y=1 $X2=0 $Y2=0
cc_133 N_A1_M1007_g N_VPWR_c_255_n 0.00291344f $X=2.195 $Y=2.46 $X2=0 $Y2=0
cc_134 N_A1_M1007_g N_VPWR_c_256_n 0.005209f $X=2.195 $Y=2.46 $X2=0 $Y2=0
cc_135 N_A1_M1007_g N_VPWR_c_253_n 0.00982765f $X=2.195 $Y=2.46 $X2=0 $Y2=0
cc_136 N_A1_M1007_g N_A_367_392#_c_290_n 0.00100081f $X=2.195 $Y=2.46 $X2=0
+ $Y2=0
cc_137 A1 N_A_367_392#_c_290_n 0.00740718f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_138 N_A1_c_164_n N_A_367_392#_c_290_n 4.66969e-19 $X=2.21 $Y=1.615 $X2=0
+ $Y2=0
cc_139 N_A1_M1007_g N_A_367_392#_c_291_n 0.0120811f $X=2.195 $Y=2.46 $X2=0 $Y2=0
cc_140 N_A1_M1007_g N_A_367_392#_c_292_n 0.0130622f $X=2.195 $Y=2.46 $X2=0 $Y2=0
cc_141 A1 N_A_367_392#_c_292_n 0.0174558f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_142 N_A1_c_164_n N_A_367_392#_c_292_n 6.27403e-19 $X=2.21 $Y=1.615 $X2=0
+ $Y2=0
cc_143 N_A1_M1007_g N_A_367_392#_c_294_n 6.43066e-19 $X=2.195 $Y=2.46 $X2=0
+ $Y2=0
cc_144 N_A1_M1004_g N_VGND_c_324_n 0.00365891f $X=2.185 $Y=1 $X2=0 $Y2=0
cc_145 A1 N_VGND_c_349_n 0.00247219f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_146 N_A1_c_164_n N_VGND_c_349_n 4.2417e-19 $X=2.21 $Y=1.615 $X2=0 $Y2=0
cc_147 N_A1_M1004_g N_VGND_c_327_n 0.0037378f $X=2.185 $Y=1 $X2=0 $Y2=0
cc_148 N_A1_M1004_g N_VGND_c_329_n 0.00110784f $X=2.185 $Y=1 $X2=0 $Y2=0
cc_149 N_A1_M1004_g N_VGND_c_331_n 0.00454494f $X=2.185 $Y=1 $X2=0 $Y2=0
cc_150 N_A2_M1002_g N_VPWR_c_255_n 0.00291344f $X=2.675 $Y=2.46 $X2=0 $Y2=0
cc_151 N_A2_M1002_g N_VPWR_c_259_n 0.005209f $X=2.675 $Y=2.46 $X2=0 $Y2=0
cc_152 N_A2_M1002_g N_VPWR_c_253_n 0.0098688f $X=2.675 $Y=2.46 $X2=0 $Y2=0
cc_153 N_A2_M1002_g N_A_367_392#_c_291_n 6.43066e-19 $X=2.675 $Y=2.46 $X2=0
+ $Y2=0
cc_154 N_A2_M1002_g N_A_367_392#_c_292_n 0.0172343f $X=2.675 $Y=2.46 $X2=0 $Y2=0
cc_155 N_A2_M1002_g N_A_367_392#_c_293_n 0.00179363f $X=2.675 $Y=2.46 $X2=0
+ $Y2=0
cc_156 N_A2_M1002_g N_A_367_392#_c_294_n 0.0122477f $X=2.675 $Y=2.46 $X2=0 $Y2=0
cc_157 N_A2_c_202_n N_VGND_c_324_n 0.0130563f $X=2.81 $Y=0.405 $X2=0 $Y2=0
cc_158 A2 N_VGND_c_324_n 0.0034499f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_159 N_A2_c_204_n N_VGND_c_324_n 0.02473f $X=3.005 $Y=0.462 $X2=0 $Y2=0
cc_160 N_A2_M1001_g N_VGND_c_357_n 0.0124199f $X=2.66 $Y=1 $X2=0 $Y2=0
cc_161 N_A2_c_204_n N_VGND_c_357_n 0.0029673f $X=3.005 $Y=0.462 $X2=0 $Y2=0
cc_162 N_A2_M1001_g N_VGND_c_329_n 0.0103623f $X=2.66 $Y=1 $X2=0 $Y2=0
cc_163 N_A2_c_200_n N_VGND_c_329_n 0.00113525f $X=2.675 $Y=1.485 $X2=0 $Y2=0
cc_164 N_A2_c_202_n N_VGND_c_329_n 0.0050123f $X=2.81 $Y=0.405 $X2=0 $Y2=0
cc_165 A2 N_VGND_c_329_n 0.00291185f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_166 N_A2_c_204_n N_VGND_c_329_n 0.0137799f $X=3.005 $Y=0.462 $X2=0 $Y2=0
cc_167 N_A2_c_202_n N_VGND_c_330_n 0.00760015f $X=2.81 $Y=0.405 $X2=0 $Y2=0
cc_168 N_A2_c_204_n N_VGND_c_330_n 0.0389306f $X=3.005 $Y=0.462 $X2=0 $Y2=0
cc_169 N_A2_c_202_n N_VGND_c_331_n 0.00934546f $X=2.81 $Y=0.405 $X2=0 $Y2=0
cc_170 N_A2_c_204_n N_VGND_c_331_n 0.0210356f $X=3.005 $Y=0.462 $X2=0 $Y2=0
cc_171 X N_VPWR_c_254_n 0.0398812f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_172 X N_VPWR_c_258_n 0.0154414f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_173 X N_VPWR_c_253_n 0.0127129f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_174 N_X_c_235_n N_VGND_c_325_n 0.00435429f $X=0.99 $Y=0.885 $X2=0 $Y2=0
cc_175 N_X_c_235_n N_VGND_c_331_n 0.00720812f $X=0.99 $Y=0.885 $X2=0 $Y2=0
cc_176 N_VPWR_c_255_n N_A_367_392#_c_291_n 0.0233858f $X=2.435 $Y=2.455 $X2=0
+ $Y2=0
cc_177 N_VPWR_c_256_n N_A_367_392#_c_291_n 0.0144623f $X=2.335 $Y=3.33 $X2=0
+ $Y2=0
cc_178 N_VPWR_c_253_n N_A_367_392#_c_291_n 0.0118344f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_179 N_VPWR_M1007_d N_A_367_392#_c_292_n 0.00197722f $X=2.285 $Y=1.96 $X2=0
+ $Y2=0
cc_180 N_VPWR_c_255_n N_A_367_392#_c_292_n 0.0151327f $X=2.435 $Y=2.455 $X2=0
+ $Y2=0
cc_181 N_VPWR_c_255_n N_A_367_392#_c_294_n 0.0233858f $X=2.435 $Y=2.455 $X2=0
+ $Y2=0
cc_182 N_VPWR_c_259_n N_A_367_392#_c_294_n 0.014549f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_183 N_VPWR_c_253_n N_A_367_392#_c_294_n 0.0119743f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_184 N_A_367_392#_c_292_n N_VGND_c_329_n 6.04679e-19 $X=2.735 $Y=2.035 $X2=0
+ $Y2=0
cc_185 N_A_367_392#_c_293_n N_VGND_c_329_n 0.0113708f $X=2.9 $Y=2.12 $X2=0 $Y2=0
cc_186 N_VGND_c_324_n A_452_136# 0.00255642f $X=2.39 $Y=0.84 $X2=-0.19
+ $Y2=-0.245
cc_187 N_VGND_c_357_n A_452_136# 0.00302954f $X=2.71 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_188 N_VGND_c_349_n A_452_136# 0.00617481f $X=2.475 $Y=0.925 $X2=-0.19
+ $Y2=-0.245

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
M1000 a_702_463# a_303_395# a_37_78# VNB nlowvt w=420000u l=150000u
+  ad=1.47e+11p pd=1.54e+06u as=2.31e+11p ps=2.78e+06u
M1001 VGND CLK a_303_395# VNB nlowvt w=740000u l=150000u
+  ad=2.086e+12p pd=1.709e+07u as=2.45475e+11p ps=2.15e+06u
M1002 a_497_395# a_303_395# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.262e+11p pd=2.14e+06u as=0p ps=0u
M1003 VGND a_2013_409# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.847e+11p ps=4.27e+06u
M1004 a_1353_392# a_497_395# a_834_355# VNB nlowvt w=740000u l=150000u
+  ad=4.58e+11p pd=3.28e+06u as=9.435e+11p ps=4.03e+06u
M1005 VGND RESET_B a_124_78# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1006 VPWR a_834_355# a_792_463# VPB pshort w=420000u l=180000u
+  ad=2.9869e+12p pd=2.378e+07u as=8.82e+10p ps=1.26e+06u
M1007 a_1630_493# a_497_395# a_1353_392# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=6.511e+11p ps=4.41e+06u
M1008 VPWR a_1353_392# a_2013_409# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.268e+11p ps=2.22e+06u
M1009 Q a_2013_409# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.552e+11p pd=5.65e+06u as=0p ps=0u
M1010 VPWR CLK a_303_395# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.32375e+11p ps=2.92e+06u
M1011 a_834_355# a_702_463# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_1678_395# a_1630_493# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_497_395# a_303_395# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1014 a_702_463# a_497_395# a_37_78# VPB pshort w=420000u l=180000u
+  ad=2.289e+11p pd=2.77e+06u as=2.289e+11p ps=2.77e+06u
M1015 a_834_355# a_702_463# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1016 a_702_463# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_124_78# D a_37_78# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_2013_409# a_1353_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1019 a_792_463# a_303_395# a_702_463# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1353_392# a_303_395# a_834_355# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_2013_409# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_1678_395# a_1647_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1023 VGND a_2013_409# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_890_138# a_834_355# a_812_138# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.008e+11p ps=1.32e+06u
M1025 a_2013_409# a_1353_392# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1678_395# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1027 VPWR a_1353_392# a_1678_395# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Q a_2013_409# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_2013_409# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1827_81# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1031 a_1678_395# a_1353_392# a_1827_81# VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1032 Q a_2013_409# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND RESET_B a_890_138# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_37_78# D VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR RESET_B a_37_78# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_812_138# a_497_395# a_702_463# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1647_81# a_303_395# a_1353_392# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 Q a_2013_409# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

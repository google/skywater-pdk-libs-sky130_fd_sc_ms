* NGSPICE file created from sky130_fd_sc_ms__einvn_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__einvn_2 A TE_B VGND VNB VPB VPWR Z
M1000 VGND a_117_74# a_231_74# VNB nlowvt w=740000u l=150000u
+  ad=3.269e+11p pd=3.45e+06u as=6.176e+11p ps=6.17e+06u
M1001 a_231_74# A Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1002 VPWR TE_B a_227_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.784e+11p pd=4.61e+06u as=9.296e+11p ps=8.38e+06u
M1003 a_227_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Z A a_227_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1005 a_227_368# A Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_117_74# TE_B VPWR VPB pshort w=640000u l=180000u
+  ad=1.76e+11p pd=1.83e+06u as=0p ps=0u
M1007 a_231_74# a_117_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Z A a_231_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_117_74# TE_B VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
.ends


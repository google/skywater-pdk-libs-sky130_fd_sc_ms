* File: sky130_fd_sc_ms__and4bb_1.pex.spice
* Created: Wed Sep  2 11:58:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__AND4BB_1%A_N 3 7 9 13 16
c30 7 0 1.61433e-19 $X=0.495 $Y=0.645
r31 15 16 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.465
+ $X2=0.505 $Y2=1.465
r32 12 15 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.27 $Y=1.465
+ $X2=0.495 $Y2=1.465
r33 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r34 9 13 7.81317 $w=2.93e-07 $l=2e-07 $layer=LI1_cond $X=0.252 $Y=1.665
+ $X2=0.252 $Y2=1.465
r35 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.465
r36 5 7 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=0.645
r37 1 16 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=1.465
r38 1 3 244.887 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_1%A_179_48# 1 2 3 12 16 19 21 22 23 25 28 30
+ 34 38 40 43 47
c107 22 0 6.72583e-20 $X=1.82 $Y=0.945
c108 21 0 1.23538e-19 $X=1.525 $Y=1.3
c109 12 0 9.12013e-20 $X=0.97 $Y=0.74
r110 37 40 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.38 $Y=1.465
+ $X2=1.525 $Y2=1.465
r111 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.38
+ $Y=1.465 $X2=1.38 $Y2=1.465
r112 32 34 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=3.46 $Y=2.2
+ $X2=3.46 $Y2=2.265
r113 31 47 2.76166 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.625 $Y=2.115
+ $X2=2.42 $Y2=2.115
r114 30 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.295 $Y=2.115
+ $X2=3.46 $Y2=2.2
r115 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.295 $Y=2.115
+ $X2=2.625 $Y2=2.115
r116 26 47 3.70735 $w=2.5e-07 $l=1.03078e-07 $layer=LI1_cond $X=2.46 $Y=2.2
+ $X2=2.42 $Y2=2.115
r117 26 28 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=2.46 $Y=2.2
+ $X2=2.46 $Y2=2.265
r118 25 47 3.70735 $w=2.5e-07 $l=1.56844e-07 $layer=LI1_cond $X=2.3 $Y=2.03
+ $X2=2.42 $Y2=2.115
r119 25 46 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=2.3 $Y=2.03 $X2=2.3
+ $Y2=1.03
r120 22 46 8.23509 $w=5.63e-07 $l=8.5e-08 $layer=LI1_cond $X=2.102 $Y=0.945
+ $X2=2.102 $Y2=1.03
r121 22 43 9.1029 $w=5.63e-07 $l=4.3e-07 $layer=LI1_cond $X=2.102 $Y=0.945
+ $X2=2.102 $Y2=0.515
r122 22 23 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.82 $Y=0.945
+ $X2=1.61 $Y2=0.945
r123 21 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.525 $Y=1.3
+ $X2=1.525 $Y2=1.465
r124 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.525 $Y=1.03
+ $X2=1.61 $Y2=0.945
r125 20 21 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.525 $Y=1.03
+ $X2=1.525 $Y2=1.3
r126 18 38 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=1.13 $Y=1.465
+ $X2=1.38 $Y2=1.465
r127 18 19 3.90195 $w=3.3e-07 $l=3.06594e-07 $layer=POLY_cond $X=1.13 $Y=1.465
+ $X2=0.895 $Y2=1.3
r128 14 19 34.7346 $w=1.65e-07 $l=3.95917e-07 $layer=POLY_cond $X=1.04 $Y=1.63
+ $X2=0.895 $Y2=1.3
r129 14 16 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.04 $Y=1.63
+ $X2=1.04 $Y2=2.4
r130 10 19 34.7346 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=0.97 $Y=1.3
+ $X2=0.895 $Y2=1.3
r131 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.97 $Y=1.3
+ $X2=0.97 $Y2=0.74
r132 3 34 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.325
+ $Y=2.12 $X2=3.46 $Y2=2.265
r133 2 28 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=2.275
+ $Y=2.12 $X2=2.46 $Y2=2.265
r134 1 43 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.37 $X2=1.985 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_1%A_27_74# 1 2 9 13 17 19 20 22 23 27 28 31
c86 28 0 2.14739e-19 $X=1.92 $Y=1.455
c87 13 0 2.32305e-19 $X=2.2 $Y=0.69
r88 31 32 6.52768 $w=5.42e-07 $l=2.9e-07 $layer=LI1_cond $X=0.427 $Y=2.115
+ $X2=0.427 $Y2=2.405
r89 28 35 76.3137 $w=5.2e-07 $l=5.05e-07 $layer=POLY_cond $X=2.015 $Y=1.455
+ $X2=2.015 $Y2=1.96
r90 28 34 47.1166 $w=5.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.015 $Y=1.455
+ $X2=2.015 $Y2=1.29
r91 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.92
+ $Y=1.455 $X2=1.92 $Y2=1.455
r92 25 27 37.6175 $w=2.63e-07 $l=8.65e-07 $layer=LI1_cond $X=1.912 $Y=2.32
+ $X2=1.912 $Y2=1.455
r93 24 32 7.66608 $w=1.7e-07 $l=3.13e-07 $layer=LI1_cond $X=0.74 $Y=2.405
+ $X2=0.427 $Y2=2.405
r94 23 25 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=1.78 $Y=2.405
+ $X2=1.912 $Y2=2.32
r95 23 24 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=1.78 $Y=2.405
+ $X2=0.74 $Y2=2.405
r96 22 31 9.97635 $w=5.42e-07 $l=2.99339e-07 $layer=LI1_cond $X=0.655 $Y=1.95
+ $X2=0.427 $Y2=2.115
r97 21 22 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.655 $Y=1.13
+ $X2=0.655 $Y2=1.95
r98 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.57 $Y=1.045
+ $X2=0.655 $Y2=1.13
r99 19 20 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.57 $Y=1.045
+ $X2=0.365 $Y2=1.045
r100 15 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.96
+ $X2=0.365 $Y2=1.045
r101 15 17 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=0.24 $Y=0.96
+ $X2=0.24 $Y2=0.645
r102 13 34 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.2 $Y=0.69 $X2=2.2
+ $Y2=1.29
r103 9 35 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=2.185 $Y=2.54
+ $X2=2.185 $Y2=1.96
r104 2 31 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r105 1 17 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_1%A_503_48# 1 2 9 12 15 16 17 20 21 24 26 27
+ 29 31 35
c89 24 0 1.65047e-19 $X=2.845 $Y=0.935
r90 34 35 5.28416 $w=1.78e-07 $l=8.5e-08 $layer=LI1_cond $X=4.145 $Y=0.94
+ $X2=4.06 $Y2=0.94
r91 31 34 23.1061 $w=1.78e-07 $l=3.75e-07 $layer=LI1_cond $X=4.52 $Y=0.94
+ $X2=4.145 $Y2=0.94
r92 31 33 4.25152 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=4.52 $Y=0.85
+ $X2=4.52 $Y2=0.735
r93 27 38 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.48 $Y=2.035
+ $X2=4.145 $Y2=2.035
r94 27 29 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=4.48 $Y=2.12
+ $X2=4.48 $Y2=2.265
r95 26 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.145 $Y=1.95
+ $X2=4.145 $Y2=2.035
r96 25 34 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=4.145 $Y=1.03 $X2=4.145
+ $Y2=0.94
r97 25 26 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.145 $Y=1.03
+ $X2=4.145 $Y2=1.95
r98 24 35 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=2.845 $Y=0.935
+ $X2=4.06 $Y2=0.935
r99 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.68
+ $Y=1.285 $X2=2.68 $Y2=1.285
r100 18 24 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=2.7 $Y=1.02
+ $X2=2.845 $Y2=0.935
r101 18 20 10.5309 $w=2.88e-07 $l=2.65e-07 $layer=LI1_cond $X=2.7 $Y=1.02
+ $X2=2.7 $Y2=1.285
r102 16 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.68 $Y=1.625
+ $X2=2.68 $Y2=1.285
r103 16 17 34.9753 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.625
+ $X2=2.68 $Y2=1.79
r104 15 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.12
+ $X2=2.68 $Y2=1.285
r105 12 17 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=2.685 $Y=2.54
+ $X2=2.685 $Y2=1.79
r106 9 15 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.59 $Y=0.69
+ $X2=2.59 $Y2=1.12
r107 2 29 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=4.345
+ $Y=2.12 $X2=4.48 $Y2=2.265
r108 1 33 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=4.38
+ $Y=0.46 $X2=4.52 $Y2=0.735
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_1%C 3 7 11 12 13 16 17
r43 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.22
+ $Y=1.355 $X2=3.22 $Y2=1.355
r44 13 17 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=3.18 $Y=1.665
+ $X2=3.18 $Y2=1.355
r45 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.22 $Y=1.695
+ $X2=3.22 $Y2=1.355
r46 11 12 35.4289 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.695
+ $X2=3.22 $Y2=1.86
r47 10 16 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.19
+ $X2=3.22 $Y2=1.355
r48 7 12 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=3.235 $Y=2.54
+ $X2=3.235 $Y2=1.86
r49 3 10 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.16 $Y=0.69 $X2=3.16
+ $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_1%D 3 7 11 12 13 16 17
r43 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.76
+ $Y=1.355 $X2=3.76 $Y2=1.355
r44 13 17 2.85631 $w=6.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.6 $Y=1.525
+ $X2=3.76 $Y2=1.525
r45 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.76 $Y=1.695
+ $X2=3.76 $Y2=1.355
r46 11 12 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.76 $Y=1.695
+ $X2=3.76 $Y2=1.86
r47 10 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.76 $Y=1.19
+ $X2=3.76 $Y2=1.355
r48 7 12 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=3.685 $Y=2.54
+ $X2=3.685 $Y2=1.86
r49 3 10 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.67 $Y=0.69 $X2=3.67
+ $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_1%B_N 3 7 9 15 16
r30 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.53
+ $Y=1.465 $X2=4.53 $Y2=1.465
r31 13 15 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=4.305 $Y=1.465
+ $X2=4.53 $Y2=1.465
r32 11 13 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=4.255 $Y=1.465
+ $X2=4.305 $Y2=1.465
r33 9 16 7.81317 $w=2.93e-07 $l=2e-07 $layer=LI1_cond $X=4.547 $Y=1.665
+ $X2=4.547 $Y2=1.465
r34 5 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.305 $Y=1.3
+ $X2=4.305 $Y2=1.465
r35 5 7 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=4.305 $Y=1.3
+ $X2=4.305 $Y2=0.735
r36 1 11 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.255 $Y=1.63
+ $X2=4.255 $Y2=1.465
r37 1 3 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=4.255 $Y=1.63
+ $X2=4.255 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_1%VPWR 1 2 3 4 17 21 25 29 32 33 35 36 38 39
+ 40 53 54 57
r65 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r66 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r67 51 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r68 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r69 48 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r70 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r71 45 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r72 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r73 42 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r74 42 44 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.98 $Y=3.33 $X2=1.68
+ $Y2=3.33
r75 40 48 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r76 40 45 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=1.68 $Y2=3.33
r77 38 50 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.815 $Y=3.33
+ $X2=3.6 $Y2=3.33
r78 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.815 $Y=3.33
+ $X2=3.98 $Y2=3.33
r79 37 53 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.145 $Y=3.33
+ $X2=4.56 $Y2=3.33
r80 37 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.145 $Y=3.33
+ $X2=3.98 $Y2=3.33
r81 35 47 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.795 $Y=3.33
+ $X2=2.64 $Y2=3.33
r82 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.795 $Y=3.33
+ $X2=2.96 $Y2=3.33
r83 34 50 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.125 $Y=3.33
+ $X2=3.6 $Y2=3.33
r84 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.125 $Y=3.33
+ $X2=2.96 $Y2=3.33
r85 32 44 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.795 $Y=3.33
+ $X2=1.68 $Y2=3.33
r86 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=3.33
+ $X2=1.96 $Y2=3.33
r87 31 47 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=2.125 $Y=3.33
+ $X2=2.64 $Y2=3.33
r88 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=3.33
+ $X2=1.96 $Y2=3.33
r89 27 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.98 $Y=3.245
+ $X2=3.98 $Y2=3.33
r90 27 29 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=3.98 $Y=3.245
+ $X2=3.98 $Y2=2.39
r91 23 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.96 $Y=3.245
+ $X2=2.96 $Y2=3.33
r92 23 25 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.96 $Y=3.245
+ $X2=2.96 $Y2=2.455
r93 19 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=3.245
+ $X2=1.96 $Y2=3.33
r94 19 21 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.96 $Y=3.245
+ $X2=1.96 $Y2=2.78
r95 15 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r96 15 17 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.78
r97 4 29 300 $w=1.7e-07 $l=3.5812e-07 $layer=licon1_PDIFF $count=2 $X=3.775
+ $Y=2.12 $X2=3.98 $Y2=2.39
r98 3 25 300 $w=1.7e-07 $l=4.17373e-07 $layer=licon1_PDIFF $count=2 $X=2.775
+ $Y=2.12 $X2=2.96 $Y2=2.455
r99 2 21 600 $w=1.7e-07 $l=7.28903e-07 $layer=licon1_PDIFF $count=1 $X=1.815
+ $Y=2.12 $X2=1.96 $Y2=2.78
r100 1 17 600 $w=1.7e-07 $l=1.04422e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.815 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_1%X 1 2 8 11 15 17 18 23
c36 17 0 1.19198e-19 $X=1.08 $Y=1.985
c37 15 0 1.61433e-19 $X=1.175 $Y=1.045
r38 18 23 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=1.2 $Y=1.985
+ $X2=1.33 $Y2=1.985
r39 17 18 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.08 $Y=1.985 $X2=1.2
+ $Y2=1.985
r40 13 15 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.995 $Y=1.045
+ $X2=1.175 $Y2=1.045
r41 9 15 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=0.96
+ $X2=1.175 $Y2=1.045
r42 9 11 25.9761 $w=1.88e-07 $l=4.45e-07 $layer=LI1_cond $X=1.175 $Y=0.96
+ $X2=1.175 $Y2=0.515
r43 8 17 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.995 $Y=1.82
+ $X2=1.08 $Y2=1.985
r44 7 13 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.995 $Y=1.13
+ $X2=0.995 $Y2=1.045
r45 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.995 $Y=1.13 $X2=0.995
+ $Y2=1.82
r46 2 23 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=1.84 $X2=1.33 $Y2=1.985
r47 1 11 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.045
+ $Y=0.37 $X2=1.185 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__AND4BB_1%VGND 1 2 9 13 16 17 18 20 33 34 37
r47 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r48 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r49 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r50 30 31 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r51 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r52 27 30 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r53 27 28 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r55 25 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r56 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r57 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r58 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r59 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r60 18 31 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.6
+ $Y2=0
r61 18 28 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.2
+ $Y2=0
r62 16 30 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.72 $Y=0 $X2=3.6
+ $Y2=0
r63 16 17 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=3.72 $Y=0 $X2=3.915
+ $Y2=0
r64 15 33 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.11 $Y=0 $X2=4.56
+ $Y2=0
r65 15 17 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.11 $Y=0 $X2=3.915
+ $Y2=0
r66 11 17 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.915 $Y=0.085
+ $X2=3.915 $Y2=0
r67 11 13 12.7064 $w=3.88e-07 $l=4.3e-07 $layer=LI1_cond $X=3.915 $Y=0.085
+ $X2=3.915 $Y2=0.515
r68 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0
r69 7 9 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0.625
r70 2 13 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=3.745
+ $Y=0.37 $X2=3.945 $Y2=0.515
r71 1 9 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.625
.ends


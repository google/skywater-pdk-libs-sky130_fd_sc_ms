* File: sky130_fd_sc_ms__mux4_4.spice
* Created: Fri Aug 28 17:41:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__mux4_4.pex.spice"
.subckt sky130_fd_sc_ms__mux4_4  VNB VPB A1 A0 S0 A2 A3 S1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* S1	S1
* A3	A3
* A2	A2
* S0	S0
* A0	A0
* A1	A1
* VPB	VPB
* VNB	VNB
MM1025 N_VGND_M1025_d N_A1_M1025_g N_A_114_126#_M1025_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1033 N_VGND_M1033_d N_A1_M1033_g N_A_114_126#_M1025_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1104 AS=0.0896 PD=0.985 PS=0.92 NRD=5.616 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1022 N_A_299_126#_M1022_d N_A0_M1022_g N_VGND_M1033_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1104 PD=0.92 PS=0.985 NRD=0 NRS=6.552 M=1 R=4.26667 SA=75001.1
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1023 N_A_299_126#_M1022_d N_A0_M1023_g N_VGND_M1023_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.3525 PD=0.92 PS=2.83 NRD=0 NRS=92.952 M=1 R=4.26667 SA=75001.6
+ SB=75000.3 A=0.096 P=1.58 MULT=1
MM1009 N_A_509_392#_M1009_d N_S0_M1009_g N_A_114_126#_M1009_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.31625 AS=0.104 PD=2.58 PS=0.965 NRD=82.332 NRS=0 M=1 R=4.26667
+ SA=75000.3 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1047 N_A_509_392#_M1047_d N_S0_M1047_g N_A_114_126#_M1009_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.104 PD=0.92 PS=0.965 NRD=0 NRS=8.436 M=1 R=4.26667
+ SA=75000.8 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1039 N_A_299_126#_M1039_d N_A_758_306#_M1039_g N_A_509_392#_M1047_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1043 N_A_299_126#_M1039_d N_A_758_306#_M1043_g N_A_509_392#_M1043_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1016 N_VGND_M1016_d N_S0_M1016_g N_A_758_306#_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_1278_121#_M1002_d N_A_758_306#_M1002_g N_A_1191_121#_M1002_s VNB
+ NLOWVT L=0.15 W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1006 N_A_1278_121#_M1002_d N_A_758_306#_M1006_g N_A_1191_121#_M1006_s VNB
+ NLOWVT L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1012 N_A_1450_121#_M1012_d N_S0_M1012_g N_A_1191_121#_M1006_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1041 N_A_1450_121#_M1012_d N_S0_M1041_g N_A_1191_121#_M1041_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.2336 PD=0.92 PS=2.01 NRD=0 NRS=14.988 M=1
+ R=4.26667 SA=75001.5 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1021 N_A_1278_121#_M1021_d N_A2_M1021_g N_VGND_M1021_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.2887 PD=0.92 PS=2.39 NRD=0 NRS=74.256 M=1 R=4.26667
+ SA=75000.3 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1040 N_A_1278_121#_M1021_d N_A2_M1040_g N_VGND_M1040_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1018 N_A_1450_121#_M1018_d N_A3_M1018_g N_VGND_M1040_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1031 N_A_1450_121#_M1018_d N_A3_M1031_g N_VGND_M1031_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1017 N_A_1191_121#_M1017_d N_S1_M1017_g N_A_2199_74#_M1017_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.166175 AS=0.1824 PD=1.255 PS=1.85 NRD=38.364 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1019 N_A_1191_121#_M1017_d N_S1_M1019_g N_A_2199_74#_M1019_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.166175 AS=0.224 PD=1.255 PS=1.34 NRD=38.364 NRS=0 M=1 R=4.26667
+ SA=75000.8 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1015 N_A_2199_74#_M1019_s N_A_2489_347#_M1015_g N_A_509_392#_M1015_s VNB
+ NLOWVT L=0.15 W=0.64 AD=0.224 AS=0.0896 PD=1.34 PS=0.92 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75001.6 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1048 N_A_2199_74#_M1048_d N_A_2489_347#_M1048_g N_A_509_392#_M1015_s VNB
+ NLOWVT L=0.15 W=0.64 AD=0.2272 AS=0.0896 PD=1.99 PS=0.92 NRD=6.552 NRS=0 M=1
+ R=4.26667 SA=75002.1 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1014 N_VGND_M1014_d N_S1_M1014_g N_A_2489_347#_M1014_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2146 AS=0.2109 PD=1.32 PS=2.05 NRD=48.648 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.2 A=0.111 P=1.78 MULT=1
MM1020 N_X_M1020_d N_A_2199_74#_M1020_g N_VGND_M1014_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2146 PD=1.02 PS=1.32 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.9
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1027 N_X_M1020_d N_A_2199_74#_M1027_g N_VGND_M1027_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.4
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1035 N_X_M1035_d N_A_2199_74#_M1035_g N_VGND_M1027_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.8
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1051 N_X_M1035_d N_A_2199_74#_M1051_g N_VGND_M1051_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_A_119_392#_M1003_d N_A1_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1004 N_A_119_392#_M1003_d N_A1_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.6
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1004_s N_A0_M1007_g N_A_299_392#_M1007_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.16 PD=1.27 PS=1.32 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90001.1
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1011_d N_A0_M1011_g N_A_299_392#_M1007_s VPB PSHORT L=0.18 W=1
+ AD=0.28 AS=0.16 PD=2.56 PS=1.32 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1000 N_A_509_392#_M1000_d N_S0_M1000_g N_A_299_392#_M1000_s VPB PSHORT L=0.18
+ W=1 AD=0.295 AS=0.1475 PD=2.59 PS=1.295 NRD=0.9653 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1042 N_A_509_392#_M1042_d N_S0_M1042_g N_A_299_392#_M1000_s VPB PSHORT L=0.18
+ W=1 AD=0.1475 AS=0.1475 PD=1.295 PS=1.295 NRD=3.9203 NRS=3.9203 M=1 R=5.55556
+ SA=90000.7 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1045 N_A_119_392#_M1045_d N_A_758_306#_M1045_g N_A_509_392#_M1042_d VPB PSHORT
+ L=0.18 W=1 AD=0.135 AS=0.1475 PD=1.27 PS=1.295 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90001.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1049 N_A_119_392#_M1045_d N_A_758_306#_M1049_g N_A_509_392#_M1049_s VPB PSHORT
+ L=0.18 W=1 AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1013_d N_S0_M1013_g N_A_758_306#_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.3136 PD=2.8 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1046 N_A_1288_377#_M1046_d N_A_758_306#_M1046_g N_A_1191_121#_M1046_s VPB
+ PSHORT L=0.18 W=1 AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1050 N_A_1288_377#_M1046_d N_A_758_306#_M1050_g N_A_1191_121#_M1050_s VPB
+ PSHORT L=0.18 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1001 N_A_1468_377#_M1001_d N_S0_M1001_g N_A_1191_121#_M1050_s VPB PSHORT
+ L=0.18 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1008 N_A_1468_377#_M1001_d N_S0_M1008_g N_A_1191_121#_M1008_s VPB PSHORT
+ L=0.18 W=1 AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90001.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1036 N_A_1468_377#_M1036_d N_A2_M1036_g N_VPWR_M1036_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.43315 PD=1.27 PS=3.2 NRD=0 NRS=74.4857 M=1 R=5.55556 SA=90000.3
+ SB=90001.7 A=0.18 P=2.36 MULT=1
MM1038 N_A_1468_377#_M1036_d N_A2_M1038_g N_VPWR_M1038_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.26025 PD=1.27 PS=1.685 NRD=0 NRS=40.4244 M=1 R=5.55556
+ SA=90000.7 SB=90001.3 A=0.18 P=2.36 MULT=1
MM1005 N_A_1288_377#_M1005_d N_A3_M1005_g N_VPWR_M1038_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.26025 PD=1.27 PS=1.685 NRD=0 NRS=40.4244 M=1 R=5.55556
+ SA=90001.4 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1024 N_A_1288_377#_M1005_d N_A3_M1024_g N_VPWR_M1024_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1032 N_A_2199_74#_M1032_d N_S1_M1032_g N_A_509_392#_M1032_s VPB PSHORT L=0.18
+ W=1 AD=0.28 AS=0.16 PD=2.56 PS=1.32 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90000.2
+ SB=90001.7 A=0.18 P=2.36 MULT=1
MM1037 N_A_2199_74#_M1037_d N_S1_M1037_g N_A_509_392#_M1032_s VPB PSHORT L=0.18
+ W=1 AD=0.16 AS=0.16 PD=1.32 PS=1.32 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90000.7
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1028 N_A_1191_121#_M1028_d N_A_2489_347#_M1028_g N_A_2199_74#_M1037_d VPB
+ PSHORT L=0.18 W=1 AD=0.16 AS=0.16 PD=1.32 PS=1.32 NRD=8.8453 NRS=0 M=1
+ R=5.55556 SA=90001.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1029 N_A_1191_121#_M1028_d N_A_2489_347#_M1029_g N_A_2199_74#_M1029_s VPB
+ PSHORT L=0.18 W=1 AD=0.16 AS=0.33 PD=1.32 PS=2.66 NRD=0 NRS=8.8453 M=1
+ R=5.55556 SA=90001.7 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1044 N_VPWR_M1044_d N_S1_M1044_g N_A_2489_347#_M1044_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1876 AS=0.3528 PD=1.455 PS=2.87 NRD=1.7533 NRS=5.2599 M=1
+ R=6.22222 SA=90000.2 SB=90002.2 A=0.2016 P=2.6 MULT=1
MM1010 N_X_M1010_d N_A_2199_74#_M1010_g N_VPWR_M1044_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1876 PD=1.39 PS=1.455 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.7
+ SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1026 N_X_M1010_d N_A_2199_74#_M1026_g N_VPWR_M1026_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.2
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1030 N_X_M1030_d N_A_2199_74#_M1030_g N_VPWR_M1026_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.7
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1034 N_X_M1030_d N_A_2199_74#_M1034_g N_VPWR_M1034_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX52_noxref VNB VPB NWDIODE A=31.9548 P=38.08
*
.include "sky130_fd_sc_ms__mux4_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__fahcin_1.spice
* Created: Wed Sep  2 12:09:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__fahcin_1.pex.spice"
.subckt sky130_fd_sc_ms__fahcin_1  VNB VPB A B CIN VPWR COUT SUM VGND
* 
* VGND	VGND
* SUM	SUM
* COUT	COUT
* VPWR	VPWR
* CIN	CIN
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_A_M1017_g N_A_28_74#_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.279859 AS=0.2109 PD=1.6087 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001 A=0.111 P=1.78 MULT=1
MM1009 N_A_259_368#_M1009_d N_A_28_74#_M1009_g N_VGND_M1017_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.242041 PD=1.85 PS=1.3913 NRD=0 NRS=76.872 M=1 R=4.26667
+ SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1014 N_A_28_74#_M1014_d N_A_492_48#_M1014_g N_A_430_418#_M1014_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1004 N_A_608_74#_M1004_d N_B_M1004_g N_A_28_74#_M1014_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.170162 AS=0.0896 PD=1.395 PS=0.92 NRD=46.872 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1025 N_A_259_368#_M1025_d N_A_492_48#_M1025_g N_A_608_74#_M1004_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1632 AS=0.170162 PD=1.15 PS=1.395 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.9 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1030 N_A_430_418#_M1030_d N_B_M1030_g N_A_259_368#_M1025_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1952 AS=0.1632 PD=1.89 PS=1.15 NRD=3.744 NRS=43.116 M=1 R=4.26667
+ SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1016 N_VGND_M1016_d N_B_M1016_g N_A_492_48#_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.212455 AS=0.222 PD=1.41565 PS=2.08 NRD=22.692 NRS=2.424 M=1 R=4.93333
+ SA=75000.2 SB=75005 A=0.111 P=1.78 MULT=1
MM1026 N_A_1200_368#_M1026_d N_A_492_48#_M1026_g N_VGND_M1016_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.183745 PD=0.92 PS=1.22435 NRD=0 NRS=29.988 M=1
+ R=4.26667 SA=75001 SB=75005.1 A=0.096 P=1.58 MULT=1
MM1001 N_COUT_M1001_d N_A_430_418#_M1001_g N_A_1200_368#_M1026_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.4528 AS=0.0896 PD=2.055 PS=0.92 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75001.4 SB=75004.6 A=0.096 P=1.58 MULT=1
MM1023 N_A_1598_400#_M1023_d N_A_608_74#_M1023_g N_COUT_M1001_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.112 AS=0.4528 PD=0.99 PS=2.055 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75002.9 SB=75003.1 A=0.096 P=1.58 MULT=1
MM1020 N_VGND_M1020_d N_CIN_M1020_g N_A_1598_400#_M1023_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.220012 AS=0.112 PD=1.53043 PS=0.99 NRD=14.052 NRS=0 M=1 R=4.26667
+ SA=75003.4 SB=75002.6 A=0.096 P=1.58 MULT=1
MM1002 N_A_1857_368#_M1002_d N_CIN_M1002_g N_VGND_M1020_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.124942 AS=0.254388 PD=1.14217 PS=1.76957 NRD=5.664 NRS=62.016 M=1
+ R=4.93333 SA=75002.8 SB=75002.6 A=0.111 P=1.78 MULT=1
MM1018 N_A_2004_136#_M1018_d N_A_608_74#_M1018_g N_A_1857_368#_M1002_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.2544 AS=0.108058 PD=1.435 PS=0.987826 NRD=14.052
+ NRS=1.872 M=1 R=4.26667 SA=75003 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1010 N_A_1967_384#_M1010_d N_A_430_418#_M1010_g N_A_2004_136#_M1018_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.1404 AS=0.2544 PD=1.145 PS=1.435 NRD=27.648 NRS=0
+ M=1 R=4.26667 SA=75004 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1000_d N_A_1857_368#_M1000_g N_A_1967_384#_M1010_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.276638 AS=0.1404 PD=1.47478 PS=1.145 NRD=78.744 NRS=0 M=1
+ R=4.26667 SA=75004.3 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1021 N_SUM_M1021_d N_A_2004_136#_M1021_g N_VGND_M1000_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.319862 PD=2.05 PS=1.70522 NRD=0 NRS=25.128 M=1 R=4.93333
+ SA=75004.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1027 N_VPWR_M1027_d N_A_M1027_g N_A_28_74#_M1027_s VPB PSHORT L=0.18 W=1.12
+ AD=0.287185 AS=0.3136 PD=1.72226 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.8 A=0.2016 P=2.6 MULT=1
MM1024 N_A_259_368#_M1024_d N_A_28_74#_M1024_g N_VPWR_M1027_d VPB PSHORT L=0.18
+ W=1 AD=0.28 AS=0.256415 PD=2.56 PS=1.53774 NRD=0 NRS=46.6102 M=1 R=5.55556
+ SA=90000.9 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1006 N_A_259_368#_M1006_d N_A_492_48#_M1006_g N_A_430_418#_M1006_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1302 AS=0.2604 PD=1.15 PS=2.3 NRD=8.1952 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90001.6 A=0.1512 P=2.04 MULT=1
MM1022 N_A_608_74#_M1022_d N_B_M1022_g N_A_259_368#_M1006_d VPB PSHORT L=0.18
+ W=0.84 AD=0.166162 AS=0.1302 PD=1.39 PS=1.15 NRD=51.5943 NRS=0 M=1 R=4.66667
+ SA=90000.7 SB=90001.2 A=0.1512 P=2.04 MULT=1
MM1007 N_A_28_74#_M1007_d N_A_492_48#_M1007_g N_A_608_74#_M1022_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2247 AS=0.166162 PD=1.375 PS=1.39 NRD=10.5395 NRS=0 M=1
+ R=4.66667 SA=90001 SB=90000.9 A=0.1512 P=2.04 MULT=1
MM1008 N_A_430_418#_M1008_d N_B_M1008_g N_A_28_74#_M1007_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2478 AS=0.2247 PD=2.27 PS=1.375 NRD=2.3443 NRS=49.2303 M=1
+ R=4.66667 SA=90001.7 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1031 N_VPWR_M1031_d N_B_M1031_g N_A_492_48#_M1031_s VPB PSHORT L=0.18 W=1.12
+ AD=0.223049 AS=0.3136 PD=1.59019 PS=2.8 NRD=1.7533 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90003.2 A=0.2016 P=2.6 MULT=1
MM1005 N_A_1200_368#_M1005_d N_A_492_48#_M1005_g N_VPWR_M1031_d VPB PSHORT
+ L=0.18 W=1 AD=0.209239 AS=0.199151 PD=1.52717 PS=1.41981 NRD=0 NRS=19.6803 M=1
+ R=5.55556 SA=90000.8 SB=90002.9 A=0.18 P=2.36 MULT=1
MM1019 N_COUT_M1019_d N_A_608_74#_M1019_g N_A_1200_368#_M1005_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.5145 AS=0.175761 PD=2.065 PS=1.28283 NRD=45.7237
+ NRS=31.6579 M=1 R=4.66667 SA=90001.3 SB=90002.9 A=0.1512 P=2.04 MULT=1
MM1013 N_A_1598_400#_M1013_d N_A_430_418#_M1013_g N_COUT_M1019_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.181696 AS=0.5145 PD=1.28739 PS=2.065 NRD=19.3454
+ NRS=39.8531 M=1 R=4.66667 SA=90002.7 SB=90001.5 A=0.1512 P=2.04 MULT=1
MM1028 N_VPWR_M1028_d N_CIN_M1028_g N_A_1598_400#_M1013_d VPB PSHORT L=0.18 W=1
+ AD=0.263491 AS=0.216304 PD=1.55189 PS=1.53261 NRD=49.7228 NRS=9.8303 M=1
+ R=5.55556 SA=90002.8 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1003 N_A_1857_368#_M1003_d N_CIN_M1003_g N_VPWR_M1028_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.295109 PD=2.8 PS=1.73811 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90003.2 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1012 N_A_2004_136#_M1012_d N_A_608_74#_M1012_g N_A_1967_384#_M1012_s VPB
+ PSHORT L=0.18 W=0.84 AD=0.1134 AS=0.2352 PD=1.11 PS=2.24 NRD=0 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1015 N_A_1857_368#_M1015_d N_A_430_418#_M1015_g N_A_2004_136#_M1012_d VPB
+ PSHORT L=0.18 W=0.84 AD=0.41895 AS=0.1134 PD=3.04 PS=1.11 NRD=104.055 NRS=0
+ M=1 R=4.66667 SA=90000.6 SB=90000.3 A=0.1512 P=2.04 MULT=1
MM1029 N_VPWR_M1029_d N_A_1857_368#_M1029_g N_A_1967_384#_M1029_s VPB PSHORT
+ L=0.18 W=1 AD=0.251698 AS=0.28 PD=1.5283 PS=2.56 NRD=44.6402 NRS=0 M=1
+ R=5.55556 SA=90000.2 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1011 N_SUM_M1011_d N_A_2004_136#_M1011_g N_VPWR_M1029_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.281902 PD=2.8 PS=1.7117 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.8 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX32_noxref VNB VPB NWDIODE A=24.8124 P=30.4
c_125 VNB 0 2.57866e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__fahcin_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__a311o_4.pxi.spice
* Created: Fri Aug 28 17:05:41 2020
* 
x_PM_SKY130_FD_SC_MS__A311O_4%C1 N_C1_M1000_g N_C1_M1017_g N_C1_M1001_g
+ N_C1_M1027_g C1 N_C1_c_141_n PM_SKY130_FD_SC_MS__A311O_4%C1
x_PM_SKY130_FD_SC_MS__A311O_4%B1 N_B1_M1005_g N_B1_M1002_g N_B1_M1012_g
+ N_B1_M1024_g B1 N_B1_c_201_n PM_SKY130_FD_SC_MS__A311O_4%B1
x_PM_SKY130_FD_SC_MS__A311O_4%A_157_392# N_A_157_392#_M1017_s
+ N_A_157_392#_M1002_s N_A_157_392#_M1007_d N_A_157_392#_M1000_d
+ N_A_157_392#_M1003_g N_A_157_392#_M1013_g N_A_157_392#_c_274_n
+ N_A_157_392#_M1019_g N_A_157_392#_M1018_g N_A_157_392#_c_275_n
+ N_A_157_392#_M1021_g N_A_157_392#_M1022_g N_A_157_392#_c_276_n
+ N_A_157_392#_M1023_g N_A_157_392#_c_262_n N_A_157_392#_c_278_n
+ N_A_157_392#_M1025_g N_A_157_392#_c_263_n N_A_157_392#_c_264_n
+ N_A_157_392#_c_265_n N_A_157_392#_c_266_n N_A_157_392#_c_267_n
+ N_A_157_392#_c_268_n N_A_157_392#_c_280_n N_A_157_392#_c_281_n
+ N_A_157_392#_c_355_p N_A_157_392#_c_269_n N_A_157_392#_c_293_n
+ N_A_157_392#_c_270_n N_A_157_392#_c_271_n N_A_157_392#_c_320_p
+ N_A_157_392#_c_272_n N_A_157_392#_c_273_n
+ PM_SKY130_FD_SC_MS__A311O_4%A_157_392#
x_PM_SKY130_FD_SC_MS__A311O_4%A3 N_A3_c_467_n N_A3_M1014_g N_A3_c_468_n
+ N_A3_c_469_n N_A3_c_470_n N_A3_M1016_g N_A3_M1004_g N_A3_M1026_g A3
+ N_A3_c_471_n N_A3_c_475_n PM_SKY130_FD_SC_MS__A311O_4%A3
x_PM_SKY130_FD_SC_MS__A311O_4%A1 N_A1_M1006_g N_A1_M1007_g N_A1_M1010_g
+ N_A1_M1009_g A1 A1 A1 N_A1_c_532_n PM_SKY130_FD_SC_MS__A311O_4%A1
x_PM_SKY130_FD_SC_MS__A311O_4%A2 N_A2_M1008_g N_A2_M1015_g N_A2_M1011_g
+ N_A2_M1020_g A2 N_A2_c_584_n PM_SKY130_FD_SC_MS__A311O_4%A2
x_PM_SKY130_FD_SC_MS__A311O_4%A_69_392# N_A_69_392#_M1000_s N_A_69_392#_M1001_s
+ N_A_69_392#_M1012_s N_A_69_392#_c_618_n N_A_69_392#_c_619_n
+ N_A_69_392#_c_620_n N_A_69_392#_c_621_n PM_SKY130_FD_SC_MS__A311O_4%A_69_392#
x_PM_SKY130_FD_SC_MS__A311O_4%A_337_392# N_A_337_392#_M1005_d
+ N_A_337_392#_M1004_s N_A_337_392#_M1006_d N_A_337_392#_M1008_d
+ N_A_337_392#_c_654_n N_A_337_392#_c_670_n N_A_337_392#_c_655_n
+ N_A_337_392#_c_656_n N_A_337_392#_c_657_n N_A_337_392#_c_658_n
+ N_A_337_392#_c_659_n N_A_337_392#_c_692_n N_A_337_392#_c_660_n
+ PM_SKY130_FD_SC_MS__A311O_4%A_337_392#
x_PM_SKY130_FD_SC_MS__A311O_4%VPWR N_VPWR_M1019_s N_VPWR_M1021_s N_VPWR_M1025_s
+ N_VPWR_M1026_d N_VPWR_M1010_s N_VPWR_M1011_s N_VPWR_c_724_n N_VPWR_c_725_n
+ N_VPWR_c_726_n N_VPWR_c_727_n N_VPWR_c_728_n N_VPWR_c_729_n N_VPWR_c_730_n
+ N_VPWR_c_731_n N_VPWR_c_732_n VPWR N_VPWR_c_733_n N_VPWR_c_734_n
+ N_VPWR_c_735_n N_VPWR_c_736_n N_VPWR_c_737_n N_VPWR_c_738_n N_VPWR_c_739_n
+ N_VPWR_c_740_n N_VPWR_c_741_n N_VPWR_c_723_n PM_SKY130_FD_SC_MS__A311O_4%VPWR
x_PM_SKY130_FD_SC_MS__A311O_4%X N_X_M1003_s N_X_M1018_s N_X_M1019_d N_X_M1023_d
+ N_X_c_832_n N_X_c_840_n N_X_c_841_n N_X_c_853_n N_X_c_854_n N_X_c_842_n
+ N_X_c_843_n N_X_c_893_n N_X_c_833_n N_X_c_834_n N_X_c_844_n N_X_c_835_n
+ N_X_c_836_n N_X_c_872_n X N_X_c_837_n N_X_c_838_n
+ PM_SKY130_FD_SC_MS__A311O_4%X
x_PM_SKY130_FD_SC_MS__A311O_4%VGND N_VGND_M1017_d N_VGND_M1027_d N_VGND_M1024_d
+ N_VGND_M1013_d N_VGND_M1022_d N_VGND_M1016_s N_VGND_c_965_n N_VGND_c_966_n
+ N_VGND_c_967_n N_VGND_c_968_n N_VGND_c_969_n N_VGND_c_970_n N_VGND_c_971_n
+ N_VGND_c_972_n N_VGND_c_973_n N_VGND_c_974_n N_VGND_c_975_n N_VGND_c_976_n
+ N_VGND_c_977_n VGND N_VGND_c_978_n N_VGND_c_979_n N_VGND_c_980_n
+ N_VGND_c_981_n N_VGND_c_982_n N_VGND_c_983_n PM_SKY130_FD_SC_MS__A311O_4%VGND
x_PM_SKY130_FD_SC_MS__A311O_4%A_888_105# N_A_888_105#_M1014_d
+ N_A_888_105#_M1015_s N_A_888_105#_c_1072_n N_A_888_105#_c_1081_n
+ N_A_888_105#_c_1073_n PM_SKY130_FD_SC_MS__A311O_4%A_888_105#
x_PM_SKY130_FD_SC_MS__A311O_4%A_1081_39# N_A_1081_39#_M1007_s
+ N_A_1081_39#_M1009_s N_A_1081_39#_M1020_d N_A_1081_39#_c_1102_n
+ N_A_1081_39#_c_1103_n N_A_1081_39#_c_1104_n N_A_1081_39#_c_1105_n
+ PM_SKY130_FD_SC_MS__A311O_4%A_1081_39#
cc_1 VNB N_C1_M1017_g 0.0351446f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.73
cc_2 VNB N_C1_M1027_g 0.0281669f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.73
cc_3 VNB C1 0.00185546f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_C1_c_141_n 0.0415109f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.62
cc_5 VNB N_B1_M1002_g 0.0302599f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.73
cc_6 VNB N_B1_M1024_g 0.0303089f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.73
cc_7 VNB B1 7.52309e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_8 VNB N_B1_c_201_n 0.0235592f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.62
cc_9 VNB N_A_157_392#_M1003_g 0.0199403f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.73
cc_10 VNB N_A_157_392#_M1013_g 0.0195521f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.62
cc_11 VNB N_A_157_392#_M1018_g 0.0188157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_157_392#_M1022_g 0.0201088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_157_392#_c_262_n 0.0135845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_157_392#_c_263_n 0.00349591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_157_392#_c_264_n 0.00131296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_157_392#_c_265_n 0.00811861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_157_392#_c_266_n 0.00336243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_157_392#_c_267_n 0.00800934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_157_392#_c_268_n 0.00741641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_157_392#_c_269_n 0.00604817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_157_392#_c_270_n 0.00443304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_157_392#_c_271_n 0.00348695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_157_392#_c_272_n 0.00364225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_157_392#_c_273_n 0.0783331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A3_c_467_n 0.0150962f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.8
cc_26 VNB N_A3_c_468_n 0.0137616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A3_c_469_n 0.00808421f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.44
cc_28 VNB N_A3_c_470_n 0.0187447f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.73
cc_29 VNB N_A3_c_471_n 0.0580992f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.62
cc_30 VNB N_A1_M1007_g 0.0264016f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.73
cc_31 VNB N_A1_M1009_g 0.0229491f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.73
cc_32 VNB A1 0.0023816f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.62
cc_33 VNB N_A1_c_532_n 0.0271611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A2_M1015_g 0.0228767f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=0.73
cc_35 VNB N_A2_M1020_g 0.0283746f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.73
cc_36 VNB A2 0.00431308f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_37 VNB N_A2_c_584_n 0.0477827f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.62
cc_38 VNB N_VPWR_c_723_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_X_c_832_n 0.0311159f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.73
cc_40 VNB N_X_c_833_n 0.00123375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_834_n 0.00225295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_X_c_835_n 0.00237374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_X_c_836_n 0.0254155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_X_c_837_n 0.0025697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_X_c_838_n 0.0105207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_965_n 0.0209749f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.635
cc_47 VNB N_VGND_c_966_n 0.00367233f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.62
cc_48 VNB N_VGND_c_967_n 0.0155164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_968_n 0.00680981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_969_n 0.0205594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_970_n 0.0101167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_971_n 0.0106292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_972_n 0.00119403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_973_n 0.0101383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_974_n 0.014713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_975_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_976_n 0.0155164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_977_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_978_n 0.0176086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_979_n 0.0884208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_980_n 0.452843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_981_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_982_n 0.00413547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_983_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_888_105#_c_1072_n 0.0030352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_888_105#_c_1073_n 0.00828173f $X=-0.19 $Y=-0.245 $X2=1.205
+ $Y2=0.73
cc_67 VNB N_A_1081_39#_c_1102_n 0.0519611f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=2.46
cc_68 VNB N_A_1081_39#_c_1103_n 0.00591587f $X=-0.19 $Y=-0.245 $X2=1.205
+ $Y2=0.73
cc_69 VNB N_A_1081_39#_c_1104_n 0.0126892f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.62
cc_70 VNB N_A_1081_39#_c_1105_n 0.024407f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.635
cc_71 VPB N_C1_M1000_g 0.0261292f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=2.46
cc_72 VPB N_C1_M1001_g 0.0204885f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=2.46
cc_73 VPB C1 0.00136459f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_74 VPB N_C1_c_141_n 0.0236142f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=1.62
cc_75 VPB N_B1_M1005_g 0.0207637f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=2.46
cc_76 VPB N_B1_M1012_g 0.0244065f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=2.46
cc_77 VPB B1 8.25483e-19 $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_78 VPB N_B1_c_201_n 0.0193069f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=1.62
cc_79 VPB N_A_157_392#_c_274_n 0.021272f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.635
cc_80 VPB N_A_157_392#_c_275_n 0.0167901f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_157_392#_c_276_n 0.0167871f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_157_392#_c_262_n 0.00815045f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_157_392#_c_278_n 0.0175672f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_157_392#_c_264_n 0.00158091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_157_392#_c_280_n 0.00305242f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_157_392#_c_281_n 0.0073332f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_157_392#_c_269_n 0.0023813f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_157_392#_c_273_n 0.0325223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A3_M1004_g 0.0250116f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=2.46
cc_90 VPB N_A3_M1026_g 0.0242211f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=0.73
cc_91 VPB N_A3_c_471_n 0.0122762f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.62
cc_92 VPB N_A3_c_475_n 0.0025127f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=1.62
cc_93 VPB N_A1_M1006_g 0.0210195f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=2.46
cc_94 VPB N_A1_M1010_g 0.022314f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=2.46
cc_95 VPB A1 0.0019514f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.62
cc_96 VPB N_A1_c_532_n 0.0162798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A2_M1008_g 0.022341f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=2.46
cc_98 VPB N_A2_M1011_g 0.0291182f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=2.46
cc_99 VPB A2 0.0037002f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_100 VPB N_A2_c_584_n 0.0314395f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.62
cc_101 VPB N_A_69_392#_c_618_n 0.00192243f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=0.73
cc_102 VPB N_A_69_392#_c_619_n 0.0169785f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_69_392#_c_620_n 0.00194885f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.62
cc_104 VPB N_A_69_392#_c_621_n 0.00656004f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.635
cc_105 VPB N_A_337_392#_c_654_n 0.00781107f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=1.44
cc_106 VPB N_A_337_392#_c_655_n 0.00135388f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.62
cc_107 VPB N_A_337_392#_c_656_n 0.00179594f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=1.62
cc_108 VPB N_A_337_392#_c_657_n 0.00337017f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=1.62
cc_109 VPB N_A_337_392#_c_658_n 0.00135978f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_337_392#_c_659_n 0.00179594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_337_392#_c_660_n 0.00231675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_724_n 0.00863475f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.635
cc_113 VPB N_VPWR_c_725_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=1.62
cc_114 VPB N_VPWR_c_726_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_727_n 0.00574883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_728_n 0.0201268f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_729_n 0.0048755f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_730_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_731_n 0.0124752f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_732_n 0.0501805f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_733_n 0.0667141f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_734_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_735_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_736_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_737_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_738_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_739_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_740_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_741_n 0.00656574f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_723_n 0.0844475f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_X_c_832_n 0.035007f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=0.73
cc_132 VPB N_X_c_840_n 0.00248381f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=0.73
cc_133 VPB N_X_c_841_n 0.0113009f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_X_c_842_n 0.0061059f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.635
cc_135 VPB N_X_c_843_n 0.00799938f $X=-0.19 $Y=1.66 $X2=1.205 $Y2=1.62
cc_136 VPB N_X_c_844_n 0.00328209f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 N_C1_M1001_g N_B1_M1005_g 0.0262313f $X=1.145 $Y=2.46 $X2=0 $Y2=0
cc_138 N_C1_M1027_g N_B1_M1002_g 0.0247525f $X=1.205 $Y=0.73 $X2=0 $Y2=0
cc_139 N_C1_c_141_n B1 0.00142809f $X=1.145 $Y=1.62 $X2=0 $Y2=0
cc_140 N_C1_c_141_n N_B1_c_201_n 0.0339424f $X=1.145 $Y=1.62 $X2=0 $Y2=0
cc_141 N_C1_M1017_g N_A_157_392#_c_263_n 0.00158318f $X=0.775 $Y=0.73 $X2=0
+ $Y2=0
cc_142 N_C1_M1027_g N_A_157_392#_c_263_n 0.00145882f $X=1.205 $Y=0.73 $X2=0
+ $Y2=0
cc_143 N_C1_M1000_g N_A_157_392#_c_264_n 0.00414972f $X=0.695 $Y=2.46 $X2=0
+ $Y2=0
cc_144 N_C1_M1017_g N_A_157_392#_c_264_n 0.00296395f $X=0.775 $Y=0.73 $X2=0
+ $Y2=0
cc_145 N_C1_M1001_g N_A_157_392#_c_264_n 0.00596014f $X=1.145 $Y=2.46 $X2=0
+ $Y2=0
cc_146 N_C1_M1027_g N_A_157_392#_c_264_n 0.00344202f $X=1.205 $Y=0.73 $X2=0
+ $Y2=0
cc_147 C1 N_A_157_392#_c_264_n 0.023546f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_148 N_C1_c_141_n N_A_157_392#_c_264_n 0.0167081f $X=1.145 $Y=1.62 $X2=0 $Y2=0
cc_149 N_C1_M1027_g N_A_157_392#_c_265_n 0.0102889f $X=1.205 $Y=0.73 $X2=0 $Y2=0
cc_150 N_C1_M1000_g N_A_157_392#_c_293_n 0.00404969f $X=0.695 $Y=2.46 $X2=0
+ $Y2=0
cc_151 N_C1_M1001_g N_A_157_392#_c_293_n 0.00460667f $X=1.145 $Y=2.46 $X2=0
+ $Y2=0
cc_152 C1 N_A_157_392#_c_293_n 0.00293704f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_153 N_C1_c_141_n N_A_157_392#_c_293_n 0.00345617f $X=1.145 $Y=1.62 $X2=0
+ $Y2=0
cc_154 N_C1_M1017_g N_A_157_392#_c_270_n 0.00266773f $X=0.775 $Y=0.73 $X2=0
+ $Y2=0
cc_155 N_C1_M1027_g N_A_157_392#_c_270_n 0.00272436f $X=1.205 $Y=0.73 $X2=0
+ $Y2=0
cc_156 N_C1_c_141_n N_A_157_392#_c_270_n 0.00265774f $X=1.145 $Y=1.62 $X2=0
+ $Y2=0
cc_157 N_C1_M1000_g N_A_69_392#_c_619_n 0.0125535f $X=0.695 $Y=2.46 $X2=0 $Y2=0
cc_158 N_C1_M1001_g N_A_69_392#_c_619_n 0.0106634f $X=1.145 $Y=2.46 $X2=0 $Y2=0
cc_159 N_C1_M1000_g N_A_69_392#_c_620_n 4.43424e-19 $X=0.695 $Y=2.46 $X2=0 $Y2=0
cc_160 N_C1_M1001_g N_A_69_392#_c_620_n 0.00455239f $X=1.145 $Y=2.46 $X2=0 $Y2=0
cc_161 N_C1_M1000_g N_VPWR_c_733_n 0.00349978f $X=0.695 $Y=2.46 $X2=0 $Y2=0
cc_162 N_C1_M1001_g N_VPWR_c_733_n 0.00347303f $X=1.145 $Y=2.46 $X2=0 $Y2=0
cc_163 N_C1_M1000_g N_VPWR_c_723_n 0.00433763f $X=0.695 $Y=2.46 $X2=0 $Y2=0
cc_164 N_C1_M1001_g N_VPWR_c_723_n 0.00428491f $X=1.145 $Y=2.46 $X2=0 $Y2=0
cc_165 N_C1_M1000_g N_X_c_832_n 0.0150035f $X=0.695 $Y=2.46 $X2=0 $Y2=0
cc_166 N_C1_M1017_g N_X_c_832_n 0.00828409f $X=0.775 $Y=0.73 $X2=0 $Y2=0
cc_167 C1 N_X_c_832_n 0.0219102f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_168 N_C1_c_141_n N_X_c_832_n 0.00345081f $X=1.145 $Y=1.62 $X2=0 $Y2=0
cc_169 N_C1_M1000_g N_X_c_840_n 0.0153579f $X=0.695 $Y=2.46 $X2=0 $Y2=0
cc_170 N_C1_M1001_g N_X_c_840_n 0.0137397f $X=1.145 $Y=2.46 $X2=0 $Y2=0
cc_171 C1 N_X_c_840_n 0.00636046f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_172 N_C1_c_141_n N_X_c_840_n 0.0016791f $X=1.145 $Y=1.62 $X2=0 $Y2=0
cc_173 N_C1_M1001_g N_X_c_853_n 0.00415377f $X=1.145 $Y=2.46 $X2=0 $Y2=0
cc_174 N_C1_M1001_g N_X_c_854_n 0.00127742f $X=1.145 $Y=2.46 $X2=0 $Y2=0
cc_175 N_C1_M1017_g N_X_c_835_n 0.0106431f $X=0.775 $Y=0.73 $X2=0 $Y2=0
cc_176 N_C1_M1027_g N_X_c_835_n 0.00641472f $X=1.205 $Y=0.73 $X2=0 $Y2=0
cc_177 C1 N_X_c_835_n 0.0103097f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_178 N_C1_c_141_n N_X_c_835_n 0.00454582f $X=1.145 $Y=1.62 $X2=0 $Y2=0
cc_179 N_C1_M1017_g N_X_c_836_n 0.001969f $X=0.775 $Y=0.73 $X2=0 $Y2=0
cc_180 N_C1_M1017_g N_X_c_838_n 0.00338785f $X=0.775 $Y=0.73 $X2=0 $Y2=0
cc_181 N_C1_M1017_g N_VGND_c_965_n 0.00806526f $X=0.775 $Y=0.73 $X2=0 $Y2=0
cc_182 N_C1_M1027_g N_VGND_c_965_n 3.98426e-19 $X=1.205 $Y=0.73 $X2=0 $Y2=0
cc_183 N_C1_M1017_g N_VGND_c_966_n 5.23778e-19 $X=0.775 $Y=0.73 $X2=0 $Y2=0
cc_184 N_C1_M1027_g N_VGND_c_966_n 0.00953485f $X=1.205 $Y=0.73 $X2=0 $Y2=0
cc_185 N_C1_M1017_g N_VGND_c_976_n 0.00455951f $X=0.775 $Y=0.73 $X2=0 $Y2=0
cc_186 N_C1_M1027_g N_VGND_c_976_n 0.00455951f $X=1.205 $Y=0.73 $X2=0 $Y2=0
cc_187 N_C1_M1017_g N_VGND_c_980_n 0.00447788f $X=0.775 $Y=0.73 $X2=0 $Y2=0
cc_188 N_C1_M1027_g N_VGND_c_980_n 0.00447788f $X=1.205 $Y=0.73 $X2=0 $Y2=0
cc_189 N_B1_M1024_g N_A_157_392#_M1003_g 0.0163992f $X=2.065 $Y=0.73 $X2=0 $Y2=0
cc_190 N_B1_M1002_g N_A_157_392#_c_264_n 8.44792e-19 $X=1.635 $Y=0.73 $X2=0
+ $Y2=0
cc_191 B1 N_A_157_392#_c_264_n 0.0126148f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_192 N_B1_c_201_n N_A_157_392#_c_264_n 0.00219292f $X=2.045 $Y=1.635 $X2=0
+ $Y2=0
cc_193 N_B1_M1002_g N_A_157_392#_c_265_n 0.0105611f $X=1.635 $Y=0.73 $X2=0 $Y2=0
cc_194 B1 N_A_157_392#_c_265_n 0.0153097f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_195 N_B1_c_201_n N_A_157_392#_c_265_n 0.00113676f $X=2.045 $Y=1.635 $X2=0
+ $Y2=0
cc_196 N_B1_M1002_g N_A_157_392#_c_266_n 0.00145882f $X=1.635 $Y=0.73 $X2=0
+ $Y2=0
cc_197 N_B1_M1024_g N_A_157_392#_c_266_n 0.00137192f $X=2.065 $Y=0.73 $X2=0
+ $Y2=0
cc_198 N_B1_M1002_g N_A_157_392#_c_267_n 9.18327e-19 $X=1.635 $Y=0.73 $X2=0
+ $Y2=0
cc_199 N_B1_M1024_g N_A_157_392#_c_267_n 0.0164591f $X=2.065 $Y=0.73 $X2=0 $Y2=0
cc_200 B1 N_A_157_392#_c_267_n 0.0220632f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_201 N_B1_c_201_n N_A_157_392#_c_267_n 0.0100451f $X=2.045 $Y=1.635 $X2=0
+ $Y2=0
cc_202 B1 N_A_157_392#_c_273_n 5.44412e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_203 N_B1_c_201_n N_A_157_392#_c_273_n 0.0224918f $X=2.045 $Y=1.635 $X2=0
+ $Y2=0
cc_204 N_B1_M1005_g N_A_69_392#_c_618_n 0.0116345f $X=1.595 $Y=2.46 $X2=0 $Y2=0
cc_205 N_B1_M1012_g N_A_69_392#_c_618_n 0.00894618f $X=2.045 $Y=2.46 $X2=0 $Y2=0
cc_206 N_B1_M1005_g N_A_69_392#_c_620_n 0.00636584f $X=1.595 $Y=2.46 $X2=0 $Y2=0
cc_207 N_B1_M1012_g N_A_69_392#_c_620_n 5.05447e-19 $X=2.045 $Y=2.46 $X2=0 $Y2=0
cc_208 N_B1_M1005_g N_A_69_392#_c_621_n 5.95939e-19 $X=1.595 $Y=2.46 $X2=0 $Y2=0
cc_209 N_B1_M1012_g N_A_69_392#_c_621_n 0.00794474f $X=2.045 $Y=2.46 $X2=0 $Y2=0
cc_210 N_B1_M1012_g N_A_337_392#_c_654_n 0.0131276f $X=2.045 $Y=2.46 $X2=0 $Y2=0
cc_211 N_B1_M1012_g N_VPWR_c_724_n 0.00127336f $X=2.045 $Y=2.46 $X2=0 $Y2=0
cc_212 N_B1_M1005_g N_VPWR_c_733_n 0.00333926f $X=1.595 $Y=2.46 $X2=0 $Y2=0
cc_213 N_B1_M1012_g N_VPWR_c_733_n 0.00335119f $X=2.045 $Y=2.46 $X2=0 $Y2=0
cc_214 N_B1_M1005_g N_VPWR_c_723_n 0.00422798f $X=1.595 $Y=2.46 $X2=0 $Y2=0
cc_215 N_B1_M1012_g N_VPWR_c_723_n 0.00426909f $X=2.045 $Y=2.46 $X2=0 $Y2=0
cc_216 N_B1_M1005_g N_X_c_840_n 0.00178373f $X=1.595 $Y=2.46 $X2=0 $Y2=0
cc_217 N_B1_M1005_g N_X_c_854_n 0.0012795f $X=1.595 $Y=2.46 $X2=0 $Y2=0
cc_218 N_B1_M1012_g N_X_c_842_n 0.00523412f $X=2.045 $Y=2.46 $X2=0 $Y2=0
cc_219 N_B1_M1024_g N_X_c_833_n 5.77553e-19 $X=2.065 $Y=0.73 $X2=0 $Y2=0
cc_220 N_B1_M1005_g N_X_c_844_n 0.0149842f $X=1.595 $Y=2.46 $X2=0 $Y2=0
cc_221 N_B1_M1012_g N_X_c_844_n 0.015785f $X=2.045 $Y=2.46 $X2=0 $Y2=0
cc_222 B1 N_X_c_844_n 0.0219009f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_223 N_B1_c_201_n N_X_c_844_n 6.2505e-19 $X=2.045 $Y=1.635 $X2=0 $Y2=0
cc_224 N_B1_M1002_g N_X_c_835_n 0.00641498f $X=1.635 $Y=0.73 $X2=0 $Y2=0
cc_225 N_B1_M1024_g N_X_c_835_n 0.00645808f $X=2.065 $Y=0.73 $X2=0 $Y2=0
cc_226 B1 N_X_c_835_n 4.24688e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_227 N_B1_M1024_g N_X_c_872_n 2.2693e-19 $X=2.065 $Y=0.73 $X2=0 $Y2=0
cc_228 N_B1_M1024_g N_X_c_837_n 3.3543e-19 $X=2.065 $Y=0.73 $X2=0 $Y2=0
cc_229 N_B1_M1002_g N_VGND_c_966_n 0.00953485f $X=1.635 $Y=0.73 $X2=0 $Y2=0
cc_230 N_B1_M1024_g N_VGND_c_966_n 5.23778e-19 $X=2.065 $Y=0.73 $X2=0 $Y2=0
cc_231 N_B1_M1002_g N_VGND_c_967_n 0.00455951f $X=1.635 $Y=0.73 $X2=0 $Y2=0
cc_232 N_B1_M1024_g N_VGND_c_967_n 0.00455951f $X=2.065 $Y=0.73 $X2=0 $Y2=0
cc_233 N_B1_M1002_g N_VGND_c_968_n 5.34522e-19 $X=1.635 $Y=0.73 $X2=0 $Y2=0
cc_234 N_B1_M1024_g N_VGND_c_968_n 0.0113902f $X=2.065 $Y=0.73 $X2=0 $Y2=0
cc_235 N_B1_M1002_g N_VGND_c_980_n 0.00447788f $X=1.635 $Y=0.73 $X2=0 $Y2=0
cc_236 N_B1_M1024_g N_VGND_c_980_n 0.00447788f $X=2.065 $Y=0.73 $X2=0 $Y2=0
cc_237 N_A_157_392#_M1022_g N_A3_c_467_n 0.0189143f $X=3.875 $Y=0.795 $X2=-0.19
+ $Y2=-0.245
cc_238 N_A_157_392#_c_268_n N_A3_c_468_n 0.00466849f $X=4.475 $Y=1.565 $X2=0
+ $Y2=0
cc_239 N_A_157_392#_c_281_n N_A3_c_468_n 0.00204554f $X=5.545 $Y=2.035 $X2=0
+ $Y2=0
cc_240 N_A_157_392#_c_262_n N_A3_c_469_n 0.0108318f $X=4.275 $Y=1.675 $X2=0
+ $Y2=0
cc_241 N_A_157_392#_c_268_n N_A3_c_469_n 0.00201387f $X=4.475 $Y=1.565 $X2=0
+ $Y2=0
cc_242 N_A_157_392#_c_320_p N_A3_c_469_n 4.05596e-19 $X=3.905 $Y=1.485 $X2=0
+ $Y2=0
cc_243 N_A_157_392#_c_273_n N_A3_c_469_n 0.00390388f $X=4.005 $Y=1.535 $X2=0
+ $Y2=0
cc_244 N_A_157_392#_c_272_n N_A3_c_470_n 0.00259763f $X=6.02 $Y=1.1 $X2=0 $Y2=0
cc_245 N_A_157_392#_c_278_n N_A3_M1004_g 0.0222201f $X=4.365 $Y=1.75 $X2=0 $Y2=0
cc_246 N_A_157_392#_c_281_n N_A3_M1004_g 0.015893f $X=5.545 $Y=2.035 $X2=0 $Y2=0
cc_247 N_A_157_392#_c_281_n N_A3_M1026_g 0.0151614f $X=5.545 $Y=2.035 $X2=0
+ $Y2=0
cc_248 N_A_157_392#_c_262_n N_A3_c_471_n 0.0222201f $X=4.275 $Y=1.675 $X2=0
+ $Y2=0
cc_249 N_A_157_392#_c_268_n N_A3_c_471_n 0.00304129f $X=4.475 $Y=1.565 $X2=0
+ $Y2=0
cc_250 N_A_157_392#_c_280_n N_A3_c_471_n 0.00491326f $X=4.56 $Y=1.95 $X2=0 $Y2=0
cc_251 N_A_157_392#_c_281_n N_A3_c_471_n 0.00290899f $X=5.545 $Y=2.035 $X2=0
+ $Y2=0
cc_252 N_A_157_392#_c_269_n N_A3_c_471_n 0.0103262f $X=5.63 $Y=1.95 $X2=0 $Y2=0
cc_253 N_A_157_392#_c_273_n N_A3_c_471_n 0.00320654f $X=4.005 $Y=1.535 $X2=0
+ $Y2=0
cc_254 N_A_157_392#_c_268_n N_A3_c_475_n 0.009987f $X=4.475 $Y=1.565 $X2=0 $Y2=0
cc_255 N_A_157_392#_c_280_n N_A3_c_475_n 0.00670292f $X=4.56 $Y=1.95 $X2=0 $Y2=0
cc_256 N_A_157_392#_c_281_n N_A3_c_475_n 0.0287463f $X=5.545 $Y=2.035 $X2=0
+ $Y2=0
cc_257 N_A_157_392#_c_269_n N_A3_c_475_n 0.020375f $X=5.63 $Y=1.95 $X2=0 $Y2=0
cc_258 N_A_157_392#_c_281_n N_A1_M1006_g 0.00425625f $X=5.545 $Y=2.035 $X2=0
+ $Y2=0
cc_259 N_A_157_392#_c_269_n N_A1_M1006_g 0.00413506f $X=5.63 $Y=1.95 $X2=0 $Y2=0
cc_260 N_A_157_392#_c_269_n N_A1_M1007_g 0.00704871f $X=5.63 $Y=1.95 $X2=0 $Y2=0
cc_261 N_A_157_392#_c_272_n N_A1_M1007_g 0.0201456f $X=6.02 $Y=1.1 $X2=0 $Y2=0
cc_262 N_A_157_392#_c_269_n N_A1_M1010_g 8.01884e-19 $X=5.63 $Y=1.95 $X2=0 $Y2=0
cc_263 N_A_157_392#_c_272_n N_A1_M1009_g 7.51231e-19 $X=6.02 $Y=1.1 $X2=0 $Y2=0
cc_264 N_A_157_392#_c_269_n A1 0.0249855f $X=5.63 $Y=1.95 $X2=0 $Y2=0
cc_265 N_A_157_392#_c_272_n A1 0.0163424f $X=6.02 $Y=1.1 $X2=0 $Y2=0
cc_266 N_A_157_392#_c_269_n N_A1_c_532_n 0.00797126f $X=5.63 $Y=1.95 $X2=0 $Y2=0
cc_267 N_A_157_392#_c_272_n N_A1_c_532_n 0.0031437f $X=6.02 $Y=1.1 $X2=0 $Y2=0
cc_268 N_A_157_392#_M1000_d N_A_69_392#_c_619_n 0.00166646f $X=0.785 $Y=1.96
+ $X2=0 $Y2=0
cc_269 N_A_157_392#_c_274_n N_A_69_392#_c_621_n 9.21806e-19 $X=3.015 $Y=1.75
+ $X2=0 $Y2=0
cc_270 N_A_157_392#_c_281_n N_A_337_392#_M1004_s 0.00165831f $X=5.545 $Y=2.035
+ $X2=0 $Y2=0
cc_271 N_A_157_392#_c_274_n N_A_337_392#_c_654_n 0.0152054f $X=3.015 $Y=1.75
+ $X2=0 $Y2=0
cc_272 N_A_157_392#_c_275_n N_A_337_392#_c_654_n 0.0130823f $X=3.465 $Y=1.75
+ $X2=0 $Y2=0
cc_273 N_A_157_392#_c_276_n N_A_337_392#_c_654_n 0.0130823f $X=3.915 $Y=1.75
+ $X2=0 $Y2=0
cc_274 N_A_157_392#_c_278_n N_A_337_392#_c_654_n 0.015687f $X=4.365 $Y=1.75
+ $X2=0 $Y2=0
cc_275 N_A_157_392#_c_268_n N_A_337_392#_c_654_n 0.00350516f $X=4.475 $Y=1.565
+ $X2=0 $Y2=0
cc_276 N_A_157_392#_c_281_n N_A_337_392#_c_654_n 0.0145314f $X=5.545 $Y=2.035
+ $X2=0 $Y2=0
cc_277 N_A_157_392#_c_355_p N_A_337_392#_c_654_n 0.00949953f $X=4.645 $Y=2.035
+ $X2=0 $Y2=0
cc_278 N_A_157_392#_c_281_n N_A_337_392#_c_670_n 0.0240577f $X=5.545 $Y=2.035
+ $X2=0 $Y2=0
cc_279 N_A_157_392#_c_281_n N_A_337_392#_c_655_n 0.00655272f $X=5.545 $Y=2.035
+ $X2=0 $Y2=0
cc_280 N_A_157_392#_c_278_n N_A_337_392#_c_660_n 7.03175e-19 $X=4.365 $Y=1.75
+ $X2=0 $Y2=0
cc_281 N_A_157_392#_c_281_n N_A_337_392#_c_660_n 0.0171986f $X=5.545 $Y=2.035
+ $X2=0 $Y2=0
cc_282 N_A_157_392#_c_280_n N_VPWR_M1025_s 0.0018358f $X=4.56 $Y=1.95 $X2=0
+ $Y2=0
cc_283 N_A_157_392#_c_281_n N_VPWR_M1025_s 0.00211299f $X=5.545 $Y=2.035 $X2=0
+ $Y2=0
cc_284 N_A_157_392#_c_355_p N_VPWR_M1025_s 0.00248996f $X=4.645 $Y=2.035 $X2=0
+ $Y2=0
cc_285 N_A_157_392#_c_281_n N_VPWR_M1026_d 0.00169018f $X=5.545 $Y=2.035 $X2=0
+ $Y2=0
cc_286 N_A_157_392#_c_274_n N_VPWR_c_724_n 0.0118211f $X=3.015 $Y=1.75 $X2=0
+ $Y2=0
cc_287 N_A_157_392#_c_275_n N_VPWR_c_724_n 0.00125818f $X=3.465 $Y=1.75 $X2=0
+ $Y2=0
cc_288 N_A_157_392#_c_274_n N_VPWR_c_725_n 0.00460063f $X=3.015 $Y=1.75 $X2=0
+ $Y2=0
cc_289 N_A_157_392#_c_275_n N_VPWR_c_725_n 0.00460063f $X=3.465 $Y=1.75 $X2=0
+ $Y2=0
cc_290 N_A_157_392#_c_274_n N_VPWR_c_726_n 0.00125818f $X=3.015 $Y=1.75 $X2=0
+ $Y2=0
cc_291 N_A_157_392#_c_275_n N_VPWR_c_726_n 0.0107196f $X=3.465 $Y=1.75 $X2=0
+ $Y2=0
cc_292 N_A_157_392#_c_276_n N_VPWR_c_726_n 0.0107196f $X=3.915 $Y=1.75 $X2=0
+ $Y2=0
cc_293 N_A_157_392#_c_278_n N_VPWR_c_726_n 0.00125818f $X=4.365 $Y=1.75 $X2=0
+ $Y2=0
cc_294 N_A_157_392#_c_276_n N_VPWR_c_727_n 0.00125818f $X=3.915 $Y=1.75 $X2=0
+ $Y2=0
cc_295 N_A_157_392#_c_278_n N_VPWR_c_727_n 0.010725f $X=4.365 $Y=1.75 $X2=0
+ $Y2=0
cc_296 N_A_157_392#_c_276_n N_VPWR_c_734_n 0.00460063f $X=3.915 $Y=1.75 $X2=0
+ $Y2=0
cc_297 N_A_157_392#_c_278_n N_VPWR_c_734_n 0.00460063f $X=4.365 $Y=1.75 $X2=0
+ $Y2=0
cc_298 N_A_157_392#_c_274_n N_VPWR_c_723_n 0.0046086f $X=3.015 $Y=1.75 $X2=0
+ $Y2=0
cc_299 N_A_157_392#_c_275_n N_VPWR_c_723_n 0.0046086f $X=3.465 $Y=1.75 $X2=0
+ $Y2=0
cc_300 N_A_157_392#_c_276_n N_VPWR_c_723_n 0.0046086f $X=3.915 $Y=1.75 $X2=0
+ $Y2=0
cc_301 N_A_157_392#_c_278_n N_VPWR_c_723_n 0.0046086f $X=4.365 $Y=1.75 $X2=0
+ $Y2=0
cc_302 N_A_157_392#_c_263_n N_X_c_832_n 0.00256949f $X=0.99 $Y=0.555 $X2=0 $Y2=0
cc_303 N_A_157_392#_c_293_n N_X_c_832_n 0.00608889f $X=1.08 $Y=2.105 $X2=0 $Y2=0
cc_304 N_A_157_392#_c_270_n N_X_c_832_n 0.00582022f $X=1.035 $Y=1.215 $X2=0
+ $Y2=0
cc_305 N_A_157_392#_M1000_d N_X_c_840_n 0.003163f $X=0.785 $Y=1.96 $X2=0 $Y2=0
cc_306 N_A_157_392#_c_293_n N_X_c_840_n 0.0205731f $X=1.08 $Y=2.105 $X2=0 $Y2=0
cc_307 N_A_157_392#_c_293_n N_X_c_853_n 0.0036619f $X=1.08 $Y=2.105 $X2=0 $Y2=0
cc_308 N_A_157_392#_c_264_n N_X_c_854_n 0.0039465f $X=1.08 $Y=2.02 $X2=0 $Y2=0
cc_309 N_A_157_392#_c_265_n N_X_c_854_n 0.00420668f $X=1.755 $Y=1.215 $X2=0
+ $Y2=0
cc_310 N_A_157_392#_c_293_n N_X_c_854_n 0.0100278f $X=1.08 $Y=2.105 $X2=0 $Y2=0
cc_311 N_A_157_392#_c_271_n N_X_c_842_n 0.0684517f $X=3.74 $Y=1.485 $X2=0 $Y2=0
cc_312 N_A_157_392#_c_273_n N_X_c_842_n 0.0117314f $X=4.005 $Y=1.535 $X2=0 $Y2=0
cc_313 N_A_157_392#_c_274_n N_X_c_843_n 0.018308f $X=3.015 $Y=1.75 $X2=0 $Y2=0
cc_314 N_A_157_392#_c_275_n N_X_c_843_n 0.0145924f $X=3.465 $Y=1.75 $X2=0 $Y2=0
cc_315 N_A_157_392#_c_276_n N_X_c_843_n 0.0145924f $X=3.915 $Y=1.75 $X2=0 $Y2=0
cc_316 N_A_157_392#_c_262_n N_X_c_843_n 0.00197799f $X=4.275 $Y=1.675 $X2=0
+ $Y2=0
cc_317 N_A_157_392#_c_278_n N_X_c_843_n 0.00502642f $X=4.365 $Y=1.75 $X2=0 $Y2=0
cc_318 N_A_157_392#_c_280_n N_X_c_843_n 0.00611406f $X=4.56 $Y=1.95 $X2=0 $Y2=0
cc_319 N_A_157_392#_c_320_p N_X_c_843_n 0.0684517f $X=3.905 $Y=1.485 $X2=0 $Y2=0
cc_320 N_A_157_392#_c_273_n N_X_c_843_n 0.00496666f $X=4.005 $Y=1.535 $X2=0
+ $Y2=0
cc_321 N_A_157_392#_M1013_g N_X_c_893_n 0.0113003f $X=2.97 $Y=0.78 $X2=0 $Y2=0
cc_322 N_A_157_392#_M1018_g N_X_c_893_n 0.0121433f $X=3.445 $Y=0.795 $X2=0 $Y2=0
cc_323 N_A_157_392#_c_271_n N_X_c_893_n 0.0554913f $X=3.74 $Y=1.485 $X2=0 $Y2=0
cc_324 N_A_157_392#_c_273_n N_X_c_893_n 0.00614392f $X=4.005 $Y=1.535 $X2=0
+ $Y2=0
cc_325 N_A_157_392#_M1003_g N_X_c_833_n 0.00454864f $X=2.54 $Y=0.78 $X2=0 $Y2=0
cc_326 N_A_157_392#_M1013_g N_X_c_833_n 7.32094e-19 $X=2.97 $Y=0.78 $X2=0 $Y2=0
cc_327 N_A_157_392#_c_266_n N_X_c_833_n 0.00293534f $X=1.85 $Y=0.555 $X2=0 $Y2=0
cc_328 N_A_157_392#_c_267_n N_X_c_833_n 0.00148317f $X=2.325 $Y=1.485 $X2=0
+ $Y2=0
cc_329 N_A_157_392#_c_271_n N_X_c_833_n 0.0249499f $X=3.74 $Y=1.485 $X2=0 $Y2=0
cc_330 N_A_157_392#_c_273_n N_X_c_833_n 0.0024556f $X=4.005 $Y=1.535 $X2=0 $Y2=0
cc_331 N_A_157_392#_M1013_g N_X_c_834_n 6.24169e-19 $X=2.97 $Y=0.78 $X2=0 $Y2=0
cc_332 N_A_157_392#_M1018_g N_X_c_834_n 0.00799917f $X=3.445 $Y=0.795 $X2=0
+ $Y2=0
cc_333 N_A_157_392#_M1022_g N_X_c_834_n 2.50179e-19 $X=3.875 $Y=0.795 $X2=0
+ $Y2=0
cc_334 N_A_157_392#_c_265_n N_X_c_844_n 7.63409e-19 $X=1.755 $Y=1.215 $X2=0
+ $Y2=0
cc_335 N_A_157_392#_c_267_n N_X_c_844_n 0.0163818f $X=2.325 $Y=1.485 $X2=0 $Y2=0
cc_336 N_A_157_392#_c_271_n N_X_c_844_n 0.00982063f $X=3.74 $Y=1.485 $X2=0 $Y2=0
cc_337 N_A_157_392#_c_273_n N_X_c_844_n 0.00158201f $X=4.005 $Y=1.535 $X2=0
+ $Y2=0
cc_338 N_A_157_392#_M1017_s N_X_c_835_n 0.00599498f $X=0.85 $Y=0.41 $X2=0 $Y2=0
cc_339 N_A_157_392#_M1002_s N_X_c_835_n 0.00438342f $X=1.71 $Y=0.41 $X2=0 $Y2=0
cc_340 N_A_157_392#_M1003_g N_X_c_835_n 0.0014982f $X=2.54 $Y=0.78 $X2=0 $Y2=0
cc_341 N_A_157_392#_c_263_n N_X_c_835_n 0.0232559f $X=0.99 $Y=0.555 $X2=0 $Y2=0
cc_342 N_A_157_392#_c_265_n N_X_c_835_n 0.0189106f $X=1.755 $Y=1.215 $X2=0 $Y2=0
cc_343 N_A_157_392#_c_266_n N_X_c_835_n 0.0197063f $X=1.85 $Y=0.555 $X2=0 $Y2=0
cc_344 N_A_157_392#_c_267_n N_X_c_835_n 0.0134082f $X=2.325 $Y=1.485 $X2=0 $Y2=0
cc_345 N_A_157_392#_c_270_n N_X_c_835_n 0.00402907f $X=1.035 $Y=1.215 $X2=0
+ $Y2=0
cc_346 N_A_157_392#_c_271_n N_X_c_835_n 0.00616549f $X=3.74 $Y=1.485 $X2=0 $Y2=0
cc_347 N_A_157_392#_c_263_n N_X_c_836_n 0.00207279f $X=0.99 $Y=0.555 $X2=0 $Y2=0
cc_348 N_A_157_392#_M1003_g N_X_c_872_n 0.00295692f $X=2.54 $Y=0.78 $X2=0 $Y2=0
cc_349 N_A_157_392#_c_266_n N_X_c_872_n 8.47036e-19 $X=1.85 $Y=0.555 $X2=0 $Y2=0
cc_350 N_A_157_392#_c_271_n N_X_c_872_n 0.00293137f $X=3.74 $Y=1.485 $X2=0 $Y2=0
cc_351 N_A_157_392#_M1003_g N_X_c_837_n 0.00926342f $X=2.54 $Y=0.78 $X2=0 $Y2=0
cc_352 N_A_157_392#_M1013_g N_X_c_837_n 0.00845441f $X=2.97 $Y=0.78 $X2=0 $Y2=0
cc_353 N_A_157_392#_M1018_g N_X_c_837_n 6.25583e-19 $X=3.445 $Y=0.795 $X2=0
+ $Y2=0
cc_354 N_A_157_392#_c_263_n N_X_c_838_n 0.00295826f $X=0.99 $Y=0.555 $X2=0 $Y2=0
cc_355 N_A_157_392#_c_267_n N_VGND_M1024_d 0.00127279f $X=2.325 $Y=1.485 $X2=0
+ $Y2=0
cc_356 N_A_157_392#_c_263_n N_VGND_c_965_n 0.00965289f $X=0.99 $Y=0.555 $X2=0
+ $Y2=0
cc_357 N_A_157_392#_c_263_n N_VGND_c_966_n 0.0234498f $X=0.99 $Y=0.555 $X2=0
+ $Y2=0
cc_358 N_A_157_392#_c_265_n N_VGND_c_966_n 0.0194236f $X=1.755 $Y=1.215 $X2=0
+ $Y2=0
cc_359 N_A_157_392#_c_266_n N_VGND_c_966_n 0.0234498f $X=1.85 $Y=0.555 $X2=0
+ $Y2=0
cc_360 N_A_157_392#_c_266_n N_VGND_c_967_n 0.00684063f $X=1.85 $Y=0.555 $X2=0
+ $Y2=0
cc_361 N_A_157_392#_M1003_g N_VGND_c_968_n 0.00516427f $X=2.54 $Y=0.78 $X2=0
+ $Y2=0
cc_362 N_A_157_392#_c_266_n N_VGND_c_968_n 0.0216242f $X=1.85 $Y=0.555 $X2=0
+ $Y2=0
cc_363 N_A_157_392#_c_267_n N_VGND_c_968_n 0.0137705f $X=2.325 $Y=1.485 $X2=0
+ $Y2=0
cc_364 N_A_157_392#_c_271_n N_VGND_c_968_n 0.00120712f $X=3.74 $Y=1.485 $X2=0
+ $Y2=0
cc_365 N_A_157_392#_M1003_g N_VGND_c_969_n 0.00467156f $X=2.54 $Y=0.78 $X2=0
+ $Y2=0
cc_366 N_A_157_392#_M1013_g N_VGND_c_969_n 0.00523933f $X=2.97 $Y=0.78 $X2=0
+ $Y2=0
cc_367 N_A_157_392#_M1013_g N_VGND_c_970_n 0.00322768f $X=2.97 $Y=0.78 $X2=0
+ $Y2=0
cc_368 N_A_157_392#_M1018_g N_VGND_c_970_n 0.00168511f $X=3.445 $Y=0.795 $X2=0
+ $Y2=0
cc_369 N_A_157_392#_M1018_g N_VGND_c_971_n 5.1451e-19 $X=3.445 $Y=0.795 $X2=0
+ $Y2=0
cc_370 N_A_157_392#_M1022_g N_VGND_c_971_n 0.0104924f $X=3.875 $Y=0.795 $X2=0
+ $Y2=0
cc_371 N_A_157_392#_M1022_g N_VGND_c_972_n 0.00356909f $X=3.875 $Y=0.795 $X2=0
+ $Y2=0
cc_372 N_A_157_392#_c_262_n N_VGND_c_972_n 0.00167287f $X=4.275 $Y=1.675 $X2=0
+ $Y2=0
cc_373 N_A_157_392#_c_268_n N_VGND_c_972_n 0.0235203f $X=4.475 $Y=1.565 $X2=0
+ $Y2=0
cc_374 N_A_157_392#_c_268_n N_VGND_c_973_n 0.0125065f $X=4.475 $Y=1.565 $X2=0
+ $Y2=0
cc_375 N_A_157_392#_c_272_n N_VGND_c_973_n 0.0128578f $X=6.02 $Y=1.1 $X2=0 $Y2=0
cc_376 N_A_157_392#_c_263_n N_VGND_c_976_n 0.00684063f $X=0.99 $Y=0.555 $X2=0
+ $Y2=0
cc_377 N_A_157_392#_M1018_g N_VGND_c_978_n 0.00514022f $X=3.445 $Y=0.795 $X2=0
+ $Y2=0
cc_378 N_A_157_392#_M1022_g N_VGND_c_978_n 0.00447026f $X=3.875 $Y=0.795 $X2=0
+ $Y2=0
cc_379 N_A_157_392#_M1003_g N_VGND_c_980_n 0.00533081f $X=2.54 $Y=0.78 $X2=0
+ $Y2=0
cc_380 N_A_157_392#_M1013_g N_VGND_c_980_n 0.00533081f $X=2.97 $Y=0.78 $X2=0
+ $Y2=0
cc_381 N_A_157_392#_M1018_g N_VGND_c_980_n 0.00528353f $X=3.445 $Y=0.795 $X2=0
+ $Y2=0
cc_382 N_A_157_392#_M1022_g N_VGND_c_980_n 0.00443817f $X=3.875 $Y=0.795 $X2=0
+ $Y2=0
cc_383 N_A_157_392#_c_263_n N_VGND_c_980_n 0.00641317f $X=0.99 $Y=0.555 $X2=0
+ $Y2=0
cc_384 N_A_157_392#_c_266_n N_VGND_c_980_n 0.00641317f $X=1.85 $Y=0.555 $X2=0
+ $Y2=0
cc_385 N_A_157_392#_M1007_d N_A_888_105#_c_1073_n 0.00338281f $X=5.88 $Y=0.585
+ $X2=0 $Y2=0
cc_386 N_A_157_392#_c_272_n N_A_888_105#_c_1073_n 0.0331424f $X=6.02 $Y=1.1
+ $X2=0 $Y2=0
cc_387 N_A_157_392#_c_272_n N_A_1081_39#_M1007_s 0.00591467f $X=6.02 $Y=1.1
+ $X2=-0.19 $Y2=-0.245
cc_388 N_A_157_392#_c_272_n N_A_1081_39#_c_1103_n 0.0112106f $X=6.02 $Y=1.1
+ $X2=0 $Y2=0
cc_389 N_A3_M1026_g N_A1_M1006_g 0.0297616f $X=5.33 $Y=2.46 $X2=0 $Y2=0
cc_390 N_A3_c_471_n N_A1_M1007_g 0.00101692f $X=5.13 $Y=1.585 $X2=0 $Y2=0
cc_391 N_A3_c_471_n N_A1_c_532_n 0.0297616f $X=5.13 $Y=1.585 $X2=0 $Y2=0
cc_392 N_A3_c_475_n N_A1_c_532_n 2.78819e-19 $X=5.13 $Y=1.585 $X2=0 $Y2=0
cc_393 N_A3_M1004_g N_A_337_392#_c_654_n 0.0102892f $X=4.88 $Y=2.46 $X2=0 $Y2=0
cc_394 N_A3_M1026_g N_A_337_392#_c_670_n 0.0126573f $X=5.33 $Y=2.46 $X2=0 $Y2=0
cc_395 N_A3_M1004_g N_A_337_392#_c_660_n 0.00914406f $X=4.88 $Y=2.46 $X2=0 $Y2=0
cc_396 N_A3_M1026_g N_A_337_392#_c_660_n 0.00897124f $X=5.33 $Y=2.46 $X2=0 $Y2=0
cc_397 N_A3_M1004_g N_VPWR_c_727_n 0.00491511f $X=4.88 $Y=2.46 $X2=0 $Y2=0
cc_398 N_A3_M1004_g N_VPWR_c_728_n 0.005209f $X=4.88 $Y=2.46 $X2=0 $Y2=0
cc_399 N_A3_M1026_g N_VPWR_c_728_n 0.005209f $X=5.33 $Y=2.46 $X2=0 $Y2=0
cc_400 N_A3_M1026_g N_VPWR_c_729_n 0.002979f $X=5.33 $Y=2.46 $X2=0 $Y2=0
cc_401 N_A3_M1004_g N_VPWR_c_723_n 0.0053328f $X=4.88 $Y=2.46 $X2=0 $Y2=0
cc_402 N_A3_M1026_g N_VPWR_c_723_n 0.00982376f $X=5.33 $Y=2.46 $X2=0 $Y2=0
cc_403 N_A3_M1004_g N_X_c_843_n 2.78366e-19 $X=4.88 $Y=2.46 $X2=0 $Y2=0
cc_404 N_A3_c_467_n N_VGND_c_971_n 0.00897916f $X=4.365 $Y=1.24 $X2=0 $Y2=0
cc_405 N_A3_c_467_n N_VGND_c_972_n 0.0136936f $X=4.365 $Y=1.24 $X2=0 $Y2=0
cc_406 N_A3_c_467_n N_VGND_c_973_n 0.0036589f $X=4.365 $Y=1.24 $X2=0 $Y2=0
cc_407 N_A3_c_468_n N_VGND_c_973_n 0.00241111f $X=4.72 $Y=1.315 $X2=0 $Y2=0
cc_408 N_A3_c_470_n N_VGND_c_973_n 0.0155579f $X=4.795 $Y=1.24 $X2=0 $Y2=0
cc_409 N_A3_c_471_n N_VGND_c_973_n 0.00822512f $X=5.13 $Y=1.585 $X2=0 $Y2=0
cc_410 N_A3_c_475_n N_VGND_c_973_n 0.0152955f $X=5.13 $Y=1.585 $X2=0 $Y2=0
cc_411 N_A3_c_467_n N_VGND_c_979_n 0.00452201f $X=4.365 $Y=1.24 $X2=0 $Y2=0
cc_412 N_A3_c_470_n N_VGND_c_979_n 0.0035868f $X=4.795 $Y=1.24 $X2=0 $Y2=0
cc_413 N_A3_c_467_n N_VGND_c_980_n 0.0049796f $X=4.365 $Y=1.24 $X2=0 $Y2=0
cc_414 N_A3_c_470_n N_VGND_c_980_n 0.0049796f $X=4.795 $Y=1.24 $X2=0 $Y2=0
cc_415 N_A3_c_467_n N_A_888_105#_c_1072_n 0.00395841f $X=4.365 $Y=1.24 $X2=0
+ $Y2=0
cc_416 N_A3_c_470_n N_A_888_105#_c_1072_n 0.00514108f $X=4.795 $Y=1.24 $X2=0
+ $Y2=0
cc_417 N_A3_c_470_n N_A_888_105#_c_1073_n 0.00989589f $X=4.795 $Y=1.24 $X2=0
+ $Y2=0
cc_418 N_A3_c_471_n N_A_888_105#_c_1073_n 0.00550459f $X=5.13 $Y=1.585 $X2=0
+ $Y2=0
cc_419 N_A3_c_475_n N_A_888_105#_c_1073_n 0.0032428f $X=5.13 $Y=1.585 $X2=0
+ $Y2=0
cc_420 N_A3_c_470_n N_A_1081_39#_c_1102_n 8.47669e-19 $X=4.795 $Y=1.24 $X2=0
+ $Y2=0
cc_421 N_A1_M1010_g N_A2_M1008_g 0.0263264f $X=6.23 $Y=2.46 $X2=0 $Y2=0
cc_422 N_A1_M1009_g N_A2_M1015_g 0.0320723f $X=6.235 $Y=0.905 $X2=0 $Y2=0
cc_423 A1 A2 0.0261825f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_424 A1 N_A2_c_584_n 0.0351268f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_425 N_A1_c_532_n N_A2_c_584_n 0.0201275f $X=6.245 $Y=1.615 $X2=0 $Y2=0
cc_426 N_A1_M1006_g N_A_337_392#_c_670_n 0.0186696f $X=5.78 $Y=2.46 $X2=0 $Y2=0
cc_427 A1 N_A_337_392#_c_655_n 0.0143383f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_428 N_A1_c_532_n N_A_337_392#_c_655_n 0.00213605f $X=6.245 $Y=1.615 $X2=0
+ $Y2=0
cc_429 N_A1_M1010_g N_A_337_392#_c_657_n 0.014478f $X=6.23 $Y=2.46 $X2=0 $Y2=0
cc_430 A1 N_A_337_392#_c_657_n 0.0565645f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_431 N_A1_c_532_n N_A_337_392#_c_657_n 0.00201785f $X=6.245 $Y=1.615 $X2=0
+ $Y2=0
cc_432 A1 N_A_337_392#_c_658_n 0.0143383f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_433 N_A1_M1006_g N_A_337_392#_c_660_n 4.97555e-19 $X=5.78 $Y=2.46 $X2=0 $Y2=0
cc_434 N_A1_M1006_g N_VPWR_c_729_n 0.00830523f $X=5.78 $Y=2.46 $X2=0 $Y2=0
cc_435 N_A1_M1010_g N_VPWR_c_729_n 4.34836e-19 $X=6.23 $Y=2.46 $X2=0 $Y2=0
cc_436 N_A1_M1006_g N_VPWR_c_730_n 4.87296e-19 $X=5.78 $Y=2.46 $X2=0 $Y2=0
cc_437 N_A1_M1010_g N_VPWR_c_730_n 0.0128666f $X=6.23 $Y=2.46 $X2=0 $Y2=0
cc_438 N_A1_M1006_g N_VPWR_c_735_n 0.00460063f $X=5.78 $Y=2.46 $X2=0 $Y2=0
cc_439 N_A1_M1010_g N_VPWR_c_735_n 0.00460063f $X=6.23 $Y=2.46 $X2=0 $Y2=0
cc_440 N_A1_M1006_g N_VPWR_c_723_n 0.00908554f $X=5.78 $Y=2.46 $X2=0 $Y2=0
cc_441 N_A1_M1010_g N_VPWR_c_723_n 0.00908554f $X=6.23 $Y=2.46 $X2=0 $Y2=0
cc_442 N_A1_M1007_g N_VGND_c_973_n 0.0012915f $X=5.805 $Y=0.905 $X2=0 $Y2=0
cc_443 N_A1_M1009_g N_A_888_105#_c_1081_n 2.33042e-19 $X=6.235 $Y=0.905 $X2=0
+ $Y2=0
cc_444 N_A1_M1007_g N_A_888_105#_c_1073_n 0.0117891f $X=5.805 $Y=0.905 $X2=0
+ $Y2=0
cc_445 N_A1_M1009_g N_A_888_105#_c_1073_n 0.0138986f $X=6.235 $Y=0.905 $X2=0
+ $Y2=0
cc_446 N_A1_M1007_g N_A_1081_39#_c_1102_n 0.00466389f $X=5.805 $Y=0.905 $X2=0
+ $Y2=0
cc_447 N_A1_M1009_g N_A_1081_39#_c_1102_n 0.00466389f $X=6.235 $Y=0.905 $X2=0
+ $Y2=0
cc_448 N_A1_M1009_g N_A_1081_39#_c_1103_n 0.00368712f $X=6.235 $Y=0.905 $X2=0
+ $Y2=0
cc_449 A1 N_A_1081_39#_c_1103_n 0.0536343f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_450 N_A1_c_532_n N_A_1081_39#_c_1103_n 0.00225398f $X=6.245 $Y=1.615 $X2=0
+ $Y2=0
cc_451 N_A2_M1008_g N_A_337_392#_c_657_n 0.014478f $X=6.71 $Y=2.46 $X2=0 $Y2=0
cc_452 N_A2_c_584_n N_A_337_392#_c_658_n 0.00209661f $X=7.16 $Y=1.615 $X2=0
+ $Y2=0
cc_453 N_A2_M1008_g N_VPWR_c_730_n 0.0128889f $X=6.71 $Y=2.46 $X2=0 $Y2=0
cc_454 N_A2_M1011_g N_VPWR_c_730_n 5.40619e-19 $X=7.16 $Y=2.46 $X2=0 $Y2=0
cc_455 N_A2_M1008_g N_VPWR_c_732_n 6.51931e-19 $X=6.71 $Y=2.46 $X2=0 $Y2=0
cc_456 N_A2_M1011_g N_VPWR_c_732_n 0.0189242f $X=7.16 $Y=2.46 $X2=0 $Y2=0
cc_457 A2 N_VPWR_c_732_n 0.0256597f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_458 N_A2_c_584_n N_VPWR_c_732_n 0.00236651f $X=7.16 $Y=1.615 $X2=0 $Y2=0
cc_459 N_A2_M1008_g N_VPWR_c_736_n 0.00460063f $X=6.71 $Y=2.46 $X2=0 $Y2=0
cc_460 N_A2_M1011_g N_VPWR_c_736_n 0.00460063f $X=7.16 $Y=2.46 $X2=0 $Y2=0
cc_461 N_A2_M1008_g N_VPWR_c_723_n 0.00908554f $X=6.71 $Y=2.46 $X2=0 $Y2=0
cc_462 N_A2_M1011_g N_VPWR_c_723_n 0.00908554f $X=7.16 $Y=2.46 $X2=0 $Y2=0
cc_463 N_A2_M1015_g N_A_888_105#_c_1081_n 0.00186627f $X=6.725 $Y=0.905 $X2=0
+ $Y2=0
cc_464 N_A2_M1020_g N_A_888_105#_c_1081_n 0.00292963f $X=7.155 $Y=0.905 $X2=0
+ $Y2=0
cc_465 N_A2_M1015_g N_A_888_105#_c_1073_n 0.00727757f $X=6.725 $Y=0.905 $X2=0
+ $Y2=0
cc_466 N_A2_M1015_g N_A_1081_39#_c_1102_n 0.00466389f $X=6.725 $Y=0.905 $X2=0
+ $Y2=0
cc_467 N_A2_M1020_g N_A_1081_39#_c_1102_n 0.0053097f $X=7.155 $Y=0.905 $X2=0
+ $Y2=0
cc_468 N_A2_M1015_g N_A_1081_39#_c_1103_n 0.014894f $X=6.725 $Y=0.905 $X2=0
+ $Y2=0
cc_469 N_A2_M1020_g N_A_1081_39#_c_1103_n 0.0173745f $X=7.155 $Y=0.905 $X2=0
+ $Y2=0
cc_470 A2 N_A_1081_39#_c_1103_n 0.00260801f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_471 N_A2_c_584_n N_A_1081_39#_c_1103_n 0.00334091f $X=7.16 $Y=1.615 $X2=0
+ $Y2=0
cc_472 A2 N_A_1081_39#_c_1104_n 0.0183965f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_473 N_A2_c_584_n N_A_1081_39#_c_1104_n 0.00193272f $X=7.16 $Y=1.615 $X2=0
+ $Y2=0
cc_474 N_A2_M1020_g N_A_1081_39#_c_1105_n 0.00526146f $X=7.155 $Y=0.905 $X2=0
+ $Y2=0
cc_475 N_A_69_392#_c_618_n N_A_337_392#_M1005_d 0.00165831f $X=2.105 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_476 N_A_69_392#_M1012_s N_A_337_392#_c_654_n 0.00508813f $X=2.135 $Y=1.96
+ $X2=0 $Y2=0
cc_477 N_A_69_392#_c_618_n N_A_337_392#_c_654_n 0.00421866f $X=2.105 $Y=2.99
+ $X2=0 $Y2=0
cc_478 N_A_69_392#_c_621_n N_A_337_392#_c_654_n 0.0206355f $X=2.27 $Y=2.78 $X2=0
+ $Y2=0
cc_479 N_A_69_392#_c_618_n N_A_337_392#_c_692_n 0.0114573f $X=2.105 $Y=2.99
+ $X2=0 $Y2=0
cc_480 N_A_69_392#_c_621_n N_VPWR_c_724_n 0.0319559f $X=2.27 $Y=2.78 $X2=0 $Y2=0
cc_481 N_A_69_392#_c_619_n N_VPWR_c_733_n 0.0366651f $X=1.205 $Y=2.887 $X2=0
+ $Y2=0
cc_482 N_A_69_392#_c_620_n N_VPWR_c_733_n 0.0581081f $X=1.535 $Y=2.887 $X2=0
+ $Y2=0
cc_483 N_A_69_392#_c_621_n N_VPWR_c_733_n 0.0225681f $X=2.27 $Y=2.78 $X2=0 $Y2=0
cc_484 N_A_69_392#_c_619_n N_VPWR_c_723_n 0.0306984f $X=1.205 $Y=2.887 $X2=0
+ $Y2=0
cc_485 N_A_69_392#_c_620_n N_VPWR_c_723_n 0.0324188f $X=1.535 $Y=2.887 $X2=0
+ $Y2=0
cc_486 N_A_69_392#_c_621_n N_VPWR_c_723_n 0.0124607f $X=2.27 $Y=2.78 $X2=0 $Y2=0
cc_487 N_A_69_392#_M1000_s N_X_c_840_n 0.00946353f $X=0.345 $Y=1.96 $X2=0 $Y2=0
cc_488 N_A_69_392#_M1001_s N_X_c_840_n 0.0035617f $X=1.235 $Y=1.96 $X2=0 $Y2=0
cc_489 N_A_69_392#_c_619_n N_X_c_840_n 0.0570304f $X=1.205 $Y=2.887 $X2=0 $Y2=0
cc_490 N_A_69_392#_c_620_n N_X_c_840_n 0.00928591f $X=1.535 $Y=2.887 $X2=0 $Y2=0
cc_491 N_A_69_392#_M1001_s N_X_c_853_n 0.0023626f $X=1.235 $Y=1.96 $X2=0 $Y2=0
cc_492 N_A_69_392#_M1001_s N_X_c_854_n 0.0039287f $X=1.235 $Y=1.96 $X2=0 $Y2=0
cc_493 N_A_69_392#_M1012_s N_X_c_844_n 0.00585802f $X=2.135 $Y=1.96 $X2=0 $Y2=0
cc_494 N_A_69_392#_c_620_n N_X_c_844_n 7.85183e-19 $X=1.535 $Y=2.887 $X2=0 $Y2=0
cc_495 N_A_337_392#_c_654_n N_VPWR_M1019_s 0.00483505f $X=4.94 $Y=2.405
+ $X2=-0.19 $Y2=1.66
cc_496 N_A_337_392#_c_654_n N_VPWR_M1021_s 0.00320919f $X=4.94 $Y=2.405 $X2=0
+ $Y2=0
cc_497 N_A_337_392#_c_654_n N_VPWR_M1025_s 0.00482714f $X=4.94 $Y=2.405 $X2=0
+ $Y2=0
cc_498 N_A_337_392#_c_670_n N_VPWR_M1026_d 0.00331838f $X=5.92 $Y=2.375 $X2=0
+ $Y2=0
cc_499 N_A_337_392#_c_657_n N_VPWR_M1010_s 0.00197722f $X=6.85 $Y=2.035 $X2=0
+ $Y2=0
cc_500 N_A_337_392#_c_654_n N_VPWR_c_724_n 0.0214945f $X=4.94 $Y=2.405 $X2=0
+ $Y2=0
cc_501 N_A_337_392#_c_654_n N_VPWR_c_726_n 0.0166513f $X=4.94 $Y=2.405 $X2=0
+ $Y2=0
cc_502 N_A_337_392#_c_654_n N_VPWR_c_727_n 0.019705f $X=4.94 $Y=2.405 $X2=0
+ $Y2=0
cc_503 N_A_337_392#_c_660_n N_VPWR_c_727_n 0.0119651f $X=5.105 $Y=2.455 $X2=0
+ $Y2=0
cc_504 N_A_337_392#_c_660_n N_VPWR_c_728_n 0.0144776f $X=5.105 $Y=2.455 $X2=0
+ $Y2=0
cc_505 N_A_337_392#_c_670_n N_VPWR_c_729_n 0.0148589f $X=5.92 $Y=2.375 $X2=0
+ $Y2=0
cc_506 N_A_337_392#_c_656_n N_VPWR_c_729_n 0.0116881f $X=6.005 $Y=2.465 $X2=0
+ $Y2=0
cc_507 N_A_337_392#_c_660_n N_VPWR_c_729_n 0.0122069f $X=5.105 $Y=2.455 $X2=0
+ $Y2=0
cc_508 N_A_337_392#_c_656_n N_VPWR_c_730_n 0.0179988f $X=6.005 $Y=2.465 $X2=0
+ $Y2=0
cc_509 N_A_337_392#_c_657_n N_VPWR_c_730_n 0.0194666f $X=6.85 $Y=2.035 $X2=0
+ $Y2=0
cc_510 N_A_337_392#_c_659_n N_VPWR_c_730_n 0.0236746f $X=6.935 $Y=2.815 $X2=0
+ $Y2=0
cc_511 N_A_337_392#_c_658_n N_VPWR_c_732_n 0.00599715f $X=6.935 $Y=2.12 $X2=0
+ $Y2=0
cc_512 N_A_337_392#_c_659_n N_VPWR_c_732_n 0.0289706f $X=6.935 $Y=2.815 $X2=0
+ $Y2=0
cc_513 N_A_337_392#_c_656_n N_VPWR_c_735_n 0.00749631f $X=6.005 $Y=2.465 $X2=0
+ $Y2=0
cc_514 N_A_337_392#_c_659_n N_VPWR_c_736_n 0.00749631f $X=6.935 $Y=2.815 $X2=0
+ $Y2=0
cc_515 N_A_337_392#_c_654_n N_VPWR_c_723_n 0.0513045f $X=4.94 $Y=2.405 $X2=0
+ $Y2=0
cc_516 N_A_337_392#_c_656_n N_VPWR_c_723_n 0.0062048f $X=6.005 $Y=2.465 $X2=0
+ $Y2=0
cc_517 N_A_337_392#_c_659_n N_VPWR_c_723_n 0.0062048f $X=6.935 $Y=2.815 $X2=0
+ $Y2=0
cc_518 N_A_337_392#_c_660_n N_VPWR_c_723_n 0.0118404f $X=5.105 $Y=2.455 $X2=0
+ $Y2=0
cc_519 N_A_337_392#_c_654_n N_X_M1019_d 0.00470972f $X=4.94 $Y=2.405 $X2=0 $Y2=0
cc_520 N_A_337_392#_c_654_n N_X_M1023_d 0.00470972f $X=4.94 $Y=2.405 $X2=0 $Y2=0
cc_521 N_A_337_392#_c_654_n N_X_c_842_n 0.102894f $X=4.94 $Y=2.405 $X2=0 $Y2=0
cc_522 N_A_337_392#_M1005_d N_X_c_844_n 0.00346931f $X=1.685 $Y=1.96 $X2=0 $Y2=0
cc_523 N_A_337_392#_c_654_n N_X_c_844_n 0.0351514f $X=4.94 $Y=2.405 $X2=0 $Y2=0
cc_524 N_A_337_392#_c_692_n N_X_c_844_n 0.0122205f $X=1.82 $Y=2.405 $X2=0 $Y2=0
cc_525 N_VPWR_c_723_n N_X_c_840_n 0.00176908f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_526 N_VPWR_c_723_n N_X_c_841_n 0.00690149f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_527 N_VPWR_M1019_s N_X_c_842_n 6.9948e-19 $X=2.665 $Y=1.84 $X2=0 $Y2=0
cc_528 N_VPWR_M1019_s N_X_c_843_n 0.00284862f $X=2.665 $Y=1.84 $X2=0 $Y2=0
cc_529 N_VPWR_M1021_s N_X_c_843_n 0.00169665f $X=3.555 $Y=1.84 $X2=0 $Y2=0
cc_530 N_X_c_835_n N_VGND_M1017_d 0.00713477f $X=2.495 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_531 N_X_c_835_n N_VGND_M1027_d 0.00212101f $X=2.495 $Y=0.925 $X2=0 $Y2=0
cc_532 N_X_c_835_n N_VGND_M1024_d 0.00654612f $X=2.495 $Y=0.925 $X2=0 $Y2=0
cc_533 N_X_c_893_n N_VGND_M1013_d 0.0041598f $X=3.495 $Y=1.065 $X2=0 $Y2=0
cc_534 N_X_c_835_n N_VGND_c_965_n 0.0162807f $X=2.495 $Y=0.925 $X2=0 $Y2=0
cc_535 N_X_c_835_n N_VGND_c_966_n 0.0241426f $X=2.495 $Y=0.925 $X2=0 $Y2=0
cc_536 N_X_c_835_n N_VGND_c_968_n 0.0189501f $X=2.495 $Y=0.925 $X2=0 $Y2=0
cc_537 N_X_c_872_n N_VGND_c_968_n 0.00118216f $X=2.64 $Y=0.925 $X2=0 $Y2=0
cc_538 N_X_c_837_n N_VGND_c_968_n 0.042245f $X=2.755 $Y=0.555 $X2=0 $Y2=0
cc_539 N_X_c_837_n N_VGND_c_969_n 0.014429f $X=2.755 $Y=0.555 $X2=0 $Y2=0
cc_540 N_X_c_893_n N_VGND_c_970_n 0.0171667f $X=3.495 $Y=1.065 $X2=0 $Y2=0
cc_541 N_X_c_834_n N_VGND_c_970_n 0.0146226f $X=3.66 $Y=0.57 $X2=0 $Y2=0
cc_542 N_X_c_837_n N_VGND_c_970_n 0.0161242f $X=2.755 $Y=0.555 $X2=0 $Y2=0
cc_543 N_X_c_834_n N_VGND_c_971_n 0.0188983f $X=3.66 $Y=0.57 $X2=0 $Y2=0
cc_544 N_X_c_834_n N_VGND_c_978_n 0.00899058f $X=3.66 $Y=0.57 $X2=0 $Y2=0
cc_545 N_X_c_834_n N_VGND_c_980_n 0.00882735f $X=3.66 $Y=0.57 $X2=0 $Y2=0
cc_546 N_X_c_837_n N_VGND_c_980_n 0.0137073f $X=2.755 $Y=0.555 $X2=0 $Y2=0
cc_547 N_X_c_838_n N_VGND_c_980_n 0.00489676f $X=0.24 $Y=0.925 $X2=0 $Y2=0
cc_548 N_VGND_c_973_n N_A_888_105#_M1014_d 0.00179007f $X=5.01 $Y=1.02 $X2=-0.19
+ $Y2=-0.245
cc_549 N_VGND_c_971_n N_A_888_105#_c_1072_n 0.0156621f $X=4.09 $Y=0.57 $X2=0
+ $Y2=0
cc_550 N_VGND_c_972_n N_A_888_105#_c_1072_n 7.25226e-19 $X=4.425 $Y=1.06 $X2=0
+ $Y2=0
cc_551 N_VGND_c_973_n N_A_888_105#_c_1072_n 0.0429099f $X=5.01 $Y=1.02 $X2=0
+ $Y2=0
cc_552 N_VGND_c_979_n N_A_888_105#_c_1072_n 0.00828248f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_553 N_VGND_c_980_n N_A_888_105#_c_1072_n 0.0105304f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_554 N_VGND_M1016_s N_A_888_105#_c_1073_n 0.00629528f $X=4.87 $Y=0.525 $X2=0
+ $Y2=0
cc_555 N_VGND_c_979_n N_A_888_105#_c_1073_n 0.0114112f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_556 N_VGND_c_980_n N_A_888_105#_c_1073_n 0.0216401f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_557 N_VGND_c_980_n N_A_1081_39#_M1007_s 0.00243084f $X=7.44 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_558 N_VGND_c_979_n N_A_1081_39#_c_1102_n 0.141318f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_559 N_VGND_c_980_n N_A_1081_39#_c_1102_n 0.0819032f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_560 N_A_888_105#_c_1073_n N_A_1081_39#_M1007_s 0.0104558f $X=6.775 $Y=0.705
+ $X2=-0.19 $Y2=-0.245
cc_561 N_A_888_105#_c_1073_n N_A_1081_39#_M1009_s 0.00495268f $X=6.775 $Y=0.705
+ $X2=0 $Y2=0
cc_562 N_A_888_105#_c_1073_n N_A_1081_39#_c_1102_n 0.107329f $X=6.775 $Y=0.705
+ $X2=0 $Y2=0
cc_563 N_A_888_105#_M1015_s N_A_1081_39#_c_1103_n 0.00179223f $X=6.8 $Y=0.585
+ $X2=0 $Y2=0
cc_564 N_A_888_105#_c_1081_n N_A_1081_39#_c_1103_n 0.016192f $X=6.94 $Y=0.73
+ $X2=0 $Y2=0
cc_565 N_A_888_105#_c_1073_n N_A_1081_39#_c_1103_n 0.0225078f $X=6.775 $Y=0.705
+ $X2=0 $Y2=0

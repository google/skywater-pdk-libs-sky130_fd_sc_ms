* File: sky130_fd_sc_ms__o21ai_2.pxi.spice
* Created: Fri Aug 28 17:54:59 2020
* 
x_PM_SKY130_FD_SC_MS__O21AI_2%A1 N_A1_M1000_g N_A1_M1009_g N_A1_M1010_g
+ N_A1_M1002_g N_A1_c_68_n N_A1_c_69_n N_A1_c_80_p N_A1_c_104_p A1 N_A1_c_70_n
+ N_A1_c_71_n PM_SKY130_FD_SC_MS__O21AI_2%A1
x_PM_SKY130_FD_SC_MS__O21AI_2%A2 N_A2_M1001_g N_A2_M1007_g N_A2_M1011_g
+ N_A2_M1003_g A2 N_A2_c_147_n N_A2_c_148_n PM_SKY130_FD_SC_MS__O21AI_2%A2
x_PM_SKY130_FD_SC_MS__O21AI_2%B1 N_B1_M1004_g N_B1_M1005_g N_B1_c_205_n
+ N_B1_c_206_n N_B1_M1006_g N_B1_c_208_n N_B1_M1008_g N_B1_c_209_n B1
+ PM_SKY130_FD_SC_MS__O21AI_2%B1
x_PM_SKY130_FD_SC_MS__O21AI_2%VPWR N_VPWR_M1000_d N_VPWR_M1002_d N_VPWR_M1006_s
+ N_VPWR_c_254_n N_VPWR_c_255_n N_VPWR_c_256_n N_VPWR_c_257_n N_VPWR_c_258_n
+ VPWR N_VPWR_c_259_n N_VPWR_c_260_n N_VPWR_c_261_n N_VPWR_c_253_n
+ PM_SKY130_FD_SC_MS__O21AI_2%VPWR
x_PM_SKY130_FD_SC_MS__O21AI_2%A_119_368# N_A_119_368#_M1000_s
+ N_A_119_368#_M1003_d N_A_119_368#_c_308_n N_A_119_368#_c_302_n
+ N_A_119_368#_c_303_n N_A_119_368#_c_304_n
+ PM_SKY130_FD_SC_MS__O21AI_2%A_119_368#
x_PM_SKY130_FD_SC_MS__O21AI_2%Y N_Y_M1005_d N_Y_M1001_s N_Y_M1004_d N_Y_c_338_n
+ N_Y_c_374_p N_Y_c_341_n N_Y_c_332_n Y Y Y Y N_Y_c_333_n
+ PM_SKY130_FD_SC_MS__O21AI_2%Y
x_PM_SKY130_FD_SC_MS__O21AI_2%A_27_74# N_A_27_74#_M1009_d N_A_27_74#_M1007_d
+ N_A_27_74#_M1010_d N_A_27_74#_M1008_s N_A_27_74#_c_375_n N_A_27_74#_c_376_n
+ N_A_27_74#_c_377_n N_A_27_74#_c_378_n N_A_27_74#_c_379_n N_A_27_74#_c_380_n
+ N_A_27_74#_c_381_n N_A_27_74#_c_382_n N_A_27_74#_c_383_n
+ PM_SKY130_FD_SC_MS__O21AI_2%A_27_74#
x_PM_SKY130_FD_SC_MS__O21AI_2%VGND N_VGND_M1009_s N_VGND_M1011_s N_VGND_c_435_n
+ N_VGND_c_436_n VGND N_VGND_c_437_n N_VGND_c_438_n N_VGND_c_439_n
+ N_VGND_c_440_n N_VGND_c_441_n N_VGND_c_442_n PM_SKY130_FD_SC_MS__O21AI_2%VGND
cc_1 VNB N_A1_M1009_g 0.0340607f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A1_M1010_g 0.0246779f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.74
cc_3 VNB N_A1_c_68_n 0.00166865f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_4 VNB N_A1_c_69_n 0.0374241f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_5 VNB N_A1_c_70_n 0.024839f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.515
cc_6 VNB N_A1_c_71_n 0.00562447f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.515
cc_7 VNB N_A2_M1007_g 0.0239739f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_8 VNB N_A2_M1011_g 0.0245225f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.74
cc_9 VNB N_A2_c_147_n 0.00175883f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.035
cc_10 VNB N_A2_c_148_n 0.0400448f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=1.95
cc_11 VNB N_B1_M1004_g 0.00232718f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_12 VNB N_B1_M1005_g 0.0262343f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_13 VNB N_B1_c_205_n 0.0134021f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=1.35
cc_14 VNB N_B1_c_206_n 0.0581295f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.74
cc_15 VNB N_B1_M1006_g 0.00368836f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.68
cc_16 VNB N_B1_c_208_n 0.0233164f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_17 VNB N_B1_c_209_n 0.0094716f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_18 VNB B1 0.00877571f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_19 VNB N_VPWR_c_253_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_332_n 0.00235393f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.035
cc_21 VNB N_Y_c_333_n 0.00472487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_375_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_23 VNB N_A_27_74#_c_376_n 0.00973995f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.95
cc_24 VNB N_A_27_74#_c_377_n 0.0143688f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_25 VNB N_A_27_74#_c_378_n 0.00220643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_74#_c_379_n 0.0124022f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.035
cc_27 VNB N_A_27_74#_c_380_n 0.00232545f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_28 VNB N_A_27_74#_c_381_n 0.00279725f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.515
cc_29 VNB N_A_27_74#_c_382_n 0.00187632f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.515
cc_30 VNB N_A_27_74#_c_383_n 0.0287634f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=1.515
cc_31 VNB N_VGND_c_435_n 0.00578139f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=1.35
cc_32 VNB N_VGND_c_436_n 0.00557884f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.68
cc_33 VNB N_VGND_c_437_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.95
cc_34 VNB N_VGND_c_438_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=1.755 $Y2=2.035
cc_35 VNB N_VGND_c_439_n 0.0399491f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.515
cc_36 VNB N_VGND_c_440_n 0.207539f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.35
cc_37 VNB N_VGND_c_441_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_442_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_A1_M1000_g 0.023717f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_40 VPB N_A1_M1002_g 0.0203785f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_41 VPB N_A1_c_68_n 0.00596297f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_42 VPB N_A1_c_69_n 0.00634597f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_43 VPB N_A1_c_70_n 0.00551453f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.515
cc_44 VPB N_A1_c_71_n 0.00263171f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.515
cc_45 VPB N_A2_M1001_g 0.0203431f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_46 VPB N_A2_M1003_g 0.0214531f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_47 VPB N_A2_c_147_n 0.00388537f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=2.035
cc_48 VPB N_A2_c_148_n 0.00674225f $X=-0.19 $Y=1.66 $X2=2.015 $Y2=1.95
cc_49 VPB N_B1_M1004_g 0.022029f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_50 VPB N_B1_M1006_g 0.0280409f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.68
cc_51 VPB N_VPWR_c_254_n 0.0106521f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=0.74
cc_52 VPB N_VPWR_c_255_n 0.0373625f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_256_n 0.00464707f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_257_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_55 VPB N_VPWR_c_258_n 0.055961f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.515
cc_56 VPB N_VPWR_c_259_n 0.0419549f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_260_n 0.0183691f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.515
cc_58 VPB N_VPWR_c_261_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_253_n 0.0605894f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_119_368#_c_302_n 0.00265439f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=0.74
cc_61 VPB N_A_119_368#_c_303_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_119_368#_c_304_n 0.00237138f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_63 VPB Y 0.0013896f $X=-0.19 $Y=1.66 $X2=2.015 $Y2=1.95
cc_64 VPB Y 0.00220527f $X=-0.19 $Y=1.66 $X2=2.075 $Y2=1.58
cc_65 VPB N_Y_c_333_n 0.00256909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 N_A1_M1000_g N_A2_M1001_g 0.0341819f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_67 N_A1_c_68_n N_A2_M1001_g 0.00121371f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_68 N_A1_c_80_p N_A2_M1001_g 0.0165241f $X=1.755 $Y=2.035 $X2=0 $Y2=0
cc_69 N_A1_M1009_g N_A2_M1007_g 0.0292811f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_70 N_A1_M1010_g N_A2_M1011_g 0.0256098f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_71 N_A1_M1002_g N_A2_M1003_g 0.0412709f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_72 N_A1_c_80_p N_A2_M1003_g 0.0130032f $X=1.755 $Y=2.035 $X2=0 $Y2=0
cc_73 N_A1_c_71_n N_A2_M1003_g 0.00496455f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_74 N_A1_M1000_g N_A2_c_147_n 6.52196e-19 $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_75 N_A1_c_68_n N_A2_c_147_n 0.0255068f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_76 N_A1_c_69_n N_A2_c_147_n 0.00123009f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_77 N_A1_c_80_p N_A2_c_147_n 0.0464043f $X=1.755 $Y=2.035 $X2=0 $Y2=0
cc_78 N_A1_c_70_n N_A2_c_147_n 0.00114794f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_79 N_A1_c_71_n N_A2_c_147_n 0.0271976f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_80 N_A1_c_68_n N_A2_c_148_n 0.00141946f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_81 N_A1_c_69_n N_A2_c_148_n 0.0171992f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_82 N_A1_c_80_p N_A2_c_148_n 7.6027e-19 $X=1.755 $Y=2.035 $X2=0 $Y2=0
cc_83 N_A1_c_70_n N_A2_c_148_n 0.0198923f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_84 N_A1_c_71_n N_A2_c_148_n 0.00136715f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_85 N_A1_M1002_g N_B1_M1004_g 0.0481146f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_86 N_A1_M1010_g N_B1_M1005_g 0.0156839f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_87 N_A1_c_70_n N_B1_M1005_g 0.00921114f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_88 N_A1_c_71_n N_B1_M1005_g 0.00173955f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_89 N_A1_c_70_n N_B1_c_209_n 0.00887611f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_90 N_A1_c_71_n N_B1_c_209_n 0.00358579f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_91 N_A1_c_68_n N_VPWR_M1000_d 0.00450592f $X=0.43 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_92 N_A1_c_104_p N_VPWR_M1000_d 0.00868688f $X=0.595 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_93 N_A1_c_80_p N_VPWR_M1002_d 0.00202466f $X=1.755 $Y=2.035 $X2=0 $Y2=0
cc_94 N_A1_M1000_g N_VPWR_c_255_n 0.00330306f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_95 N_A1_c_69_n N_VPWR_c_255_n 3.12191e-19 $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_96 N_A1_c_104_p N_VPWR_c_255_n 0.00833996f $X=0.595 $Y=2.035 $X2=0 $Y2=0
cc_97 N_A1_M1002_g N_VPWR_c_256_n 0.00126485f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_98 N_A1_M1000_g N_VPWR_c_259_n 0.00517089f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_99 N_A1_M1002_g N_VPWR_c_259_n 0.00518311f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_100 N_A1_M1000_g N_VPWR_c_253_n 0.0098133f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_101 N_A1_M1002_g N_VPWR_c_253_n 0.0098186f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_102 N_A1_c_80_p N_A_119_368#_M1000_s 0.00761058f $X=1.755 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_103 N_A1_c_80_p N_A_119_368#_M1003_d 0.00799623f $X=1.755 $Y=2.035 $X2=0
+ $Y2=0
cc_104 N_A1_c_71_n N_A_119_368#_M1003_d 0.00148857f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_105 N_A1_M1000_g N_A_119_368#_c_308_n 0.00809354f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A1_c_80_p N_A_119_368#_c_308_n 0.0148589f $X=1.755 $Y=2.035 $X2=0 $Y2=0
cc_107 N_A1_c_104_p N_A_119_368#_c_308_n 0.00237022f $X=0.595 $Y=2.035 $X2=0
+ $Y2=0
cc_108 N_A1_M1000_g N_A_119_368#_c_303_n 0.00358315f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_109 N_A1_M1002_g N_A_119_368#_c_304_n 0.00711276f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_110 N_A1_c_80_p N_Y_M1001_s 0.00410538f $X=1.755 $Y=2.035 $X2=0 $Y2=0
cc_111 N_A1_M1002_g N_Y_c_338_n 0.0162371f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_112 N_A1_c_80_p N_Y_c_338_n 0.0519142f $X=1.755 $Y=2.035 $X2=0 $Y2=0
cc_113 N_A1_c_70_n N_Y_c_338_n 2.57541e-19 $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_114 N_A1_M1002_g N_Y_c_341_n 8.26958e-19 $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_115 N_A1_c_80_p N_Y_c_341_n 0.0183291f $X=1.755 $Y=2.035 $X2=0 $Y2=0
cc_116 N_A1_c_71_n N_Y_c_333_n 0.0301737f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_117 N_A1_M1009_g N_A_27_74#_c_375_n 0.0101985f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_118 N_A1_M1009_g N_A_27_74#_c_376_n 0.0114775f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_119 N_A1_c_68_n N_A_27_74#_c_376_n 0.0114058f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_120 N_A1_M1009_g N_A_27_74#_c_377_n 0.00214612f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_121 N_A1_c_68_n N_A_27_74#_c_377_n 0.0158461f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_122 N_A1_c_69_n N_A_27_74#_c_377_n 0.0012184f $X=0.43 $Y=1.515 $X2=0 $Y2=0
cc_123 N_A1_M1010_g N_A_27_74#_c_378_n 9.34885e-19 $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_124 N_A1_M1010_g N_A_27_74#_c_379_n 0.0133221f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A1_c_70_n N_A_27_74#_c_379_n 0.0012814f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_126 N_A1_c_71_n N_A_27_74#_c_379_n 0.0436794f $X=1.92 $Y=1.515 $X2=0 $Y2=0
cc_127 N_A1_M1009_g N_VGND_c_435_n 0.00565822f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A1_M1010_g N_VGND_c_436_n 0.0106192f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_129 N_A1_M1009_g N_VGND_c_437_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A1_M1010_g N_VGND_c_439_n 0.00383152f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A1_M1009_g N_VGND_c_440_n 0.00824429f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A1_M1010_g N_VGND_c_440_n 0.00758041f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A2_M1001_g N_VPWR_c_259_n 0.00333896f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_134 N_A2_M1003_g N_VPWR_c_259_n 0.00333926f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_135 N_A2_M1001_g N_VPWR_c_253_n 0.00423284f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_136 N_A2_M1003_g N_VPWR_c_253_n 0.00423742f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A2_M1001_g N_A_119_368#_c_308_n 0.00894678f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_138 N_A2_M1003_g N_A_119_368#_c_308_n 6.52581e-19 $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A2_M1001_g N_A_119_368#_c_302_n 0.0118818f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A2_M1003_g N_A_119_368#_c_302_n 0.0103386f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_141 N_A2_M1001_g N_A_119_368#_c_303_n 0.001916f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_142 N_A2_M1003_g N_A_119_368#_c_304_n 4.1224e-19 $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_143 N_A2_M1003_g N_Y_c_338_n 0.010604f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A2_M1003_g N_Y_c_341_n 0.00697729f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_145 N_A2_M1007_g N_A_27_74#_c_375_n 9.46832e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A2_M1007_g N_A_27_74#_c_376_n 0.0134647f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A2_c_147_n N_A_27_74#_c_376_n 0.0209068f $X=1.35 $Y=1.515 $X2=0 $Y2=0
cc_148 N_A2_c_148_n N_A_27_74#_c_376_n 5.16483e-19 $X=1.44 $Y=1.515 $X2=0 $Y2=0
cc_149 N_A2_M1007_g N_A_27_74#_c_378_n 4.13268e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A2_M1011_g N_A_27_74#_c_378_n 0.00837823f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A2_M1011_g N_A_27_74#_c_379_n 0.0124938f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A2_c_147_n N_A_27_74#_c_379_n 0.0101599f $X=1.35 $Y=1.515 $X2=0 $Y2=0
cc_153 N_A2_c_148_n N_A_27_74#_c_379_n 0.0010611f $X=1.44 $Y=1.515 $X2=0 $Y2=0
cc_154 N_A2_M1011_g N_A_27_74#_c_382_n 0.00115653f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A2_c_147_n N_A_27_74#_c_382_n 0.0215332f $X=1.35 $Y=1.515 $X2=0 $Y2=0
cc_156 N_A2_c_148_n N_A_27_74#_c_382_n 9.10195e-19 $X=1.44 $Y=1.515 $X2=0 $Y2=0
cc_157 N_A2_M1007_g N_VGND_c_435_n 0.0106183f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A2_M1011_g N_VGND_c_435_n 5.10607e-19 $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A2_M1011_g N_VGND_c_436_n 0.00233634f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A2_M1007_g N_VGND_c_438_n 0.00383152f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A2_M1011_g N_VGND_c_438_n 0.00451267f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A2_M1007_g N_VGND_c_440_n 0.00757689f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A2_M1011_g N_VGND_c_440_n 0.00875489f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_164 N_B1_M1004_g N_VPWR_c_256_n 0.00834492f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_165 N_B1_M1006_g N_VPWR_c_256_n 4.43428e-19 $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_166 N_B1_c_206_n N_VPWR_c_258_n 0.00178067f $X=2.855 $Y=1.615 $X2=0 $Y2=0
cc_167 N_B1_M1006_g N_VPWR_c_258_n 0.00517389f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_168 B1 N_VPWR_c_258_n 0.0143742f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_169 N_B1_M1004_g N_VPWR_c_260_n 0.00460063f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_170 N_B1_M1006_g N_VPWR_c_260_n 0.005209f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_171 N_B1_M1004_g N_VPWR_c_253_n 0.00908554f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_172 N_B1_M1006_g N_VPWR_c_253_n 0.00986008f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_173 N_B1_M1004_g N_Y_c_338_n 0.0194478f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_174 N_B1_M1005_g N_Y_c_332_n 3.52947e-19 $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_175 N_B1_c_208_n N_Y_c_332_n 0.00177298f $X=2.865 $Y=1.22 $X2=0 $Y2=0
cc_176 N_B1_M1006_g Y 0.00337098f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_177 N_B1_M1004_g Y 2.66702e-19 $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_178 N_B1_M1006_g Y 0.00932618f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_179 N_B1_M1006_g Y 0.00440001f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_180 N_B1_M1004_g N_Y_c_333_n 0.00209013f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_181 N_B1_M1005_g N_Y_c_333_n 0.00491952f $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_182 N_B1_c_205_n N_Y_c_333_n 0.0181024f $X=2.765 $Y=1.492 $X2=0 $Y2=0
cc_183 N_B1_c_206_n N_Y_c_333_n 0.00177298f $X=2.855 $Y=1.615 $X2=0 $Y2=0
cc_184 N_B1_M1006_g N_Y_c_333_n 0.00524105f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_185 B1 N_Y_c_333_n 0.0275294f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_186 N_B1_M1005_g N_A_27_74#_c_379_n 7.03414e-19 $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_187 N_B1_M1005_g N_A_27_74#_c_381_n 0.0128435f $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_188 N_B1_c_208_n N_A_27_74#_c_381_n 0.0107617f $X=2.865 $Y=1.22 $X2=0 $Y2=0
cc_189 N_B1_M1005_g N_A_27_74#_c_383_n 6.09607e-19 $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_190 N_B1_c_206_n N_A_27_74#_c_383_n 0.00191451f $X=2.855 $Y=1.615 $X2=0 $Y2=0
cc_191 N_B1_c_208_n N_A_27_74#_c_383_n 0.00847698f $X=2.865 $Y=1.22 $X2=0 $Y2=0
cc_192 B1 N_A_27_74#_c_383_n 0.0251165f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_193 N_B1_M1005_g N_VGND_c_436_n 5.93944e-19 $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_194 N_B1_M1005_g N_VGND_c_439_n 0.00291649f $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_195 N_B1_c_208_n N_VGND_c_439_n 0.00291626f $X=2.865 $Y=1.22 $X2=0 $Y2=0
cc_196 N_B1_M1005_g N_VGND_c_440_n 0.00359962f $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_197 N_B1_c_208_n N_VGND_c_440_n 0.00363101f $X=2.865 $Y=1.22 $X2=0 $Y2=0
cc_198 N_VPWR_c_259_n N_A_119_368#_c_302_n 0.0421734f $X=2.095 $Y=3.33 $X2=0
+ $Y2=0
cc_199 N_VPWR_c_253_n N_A_119_368#_c_302_n 0.0236854f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_200 N_VPWR_c_255_n N_A_119_368#_c_303_n 0.0103534f $X=0.28 $Y=2.455 $X2=0
+ $Y2=0
cc_201 N_VPWR_c_259_n N_A_119_368#_c_303_n 0.0234131f $X=2.095 $Y=3.33 $X2=0
+ $Y2=0
cc_202 N_VPWR_c_253_n N_A_119_368#_c_303_n 0.0125504f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_203 N_VPWR_c_256_n N_A_119_368#_c_304_n 0.0187169f $X=2.18 $Y=2.805 $X2=0
+ $Y2=0
cc_204 N_VPWR_c_259_n N_A_119_368#_c_304_n 0.0226835f $X=2.095 $Y=3.33 $X2=0
+ $Y2=0
cc_205 N_VPWR_c_253_n N_A_119_368#_c_304_n 0.0124822f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_206 N_VPWR_M1002_d N_Y_c_338_n 0.00331662f $X=2.045 $Y=1.84 $X2=0 $Y2=0
cc_207 N_VPWR_c_256_n N_Y_c_338_n 0.0148589f $X=2.18 $Y=2.805 $X2=0 $Y2=0
cc_208 N_VPWR_c_258_n Y 0.0156277f $X=3.08 $Y=1.985 $X2=0 $Y2=0
cc_209 N_VPWR_c_256_n Y 0.0127584f $X=2.18 $Y=2.805 $X2=0 $Y2=0
cc_210 N_VPWR_c_258_n Y 0.017257f $X=3.08 $Y=1.985 $X2=0 $Y2=0
cc_211 N_VPWR_c_260_n Y 0.0118717f $X=2.995 $Y=3.33 $X2=0 $Y2=0
cc_212 N_VPWR_c_253_n Y 0.00975826f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_213 N_A_119_368#_c_302_n N_Y_M1001_s 0.00218982f $X=1.565 $Y=2.99 $X2=0 $Y2=0
cc_214 N_A_119_368#_M1003_d N_Y_c_338_n 0.00432698f $X=1.545 $Y=1.84 $X2=0 $Y2=0
cc_215 N_A_119_368#_c_302_n N_Y_c_338_n 0.00464895f $X=1.565 $Y=2.99 $X2=0 $Y2=0
cc_216 N_A_119_368#_c_304_n N_Y_c_338_n 0.0182896f $X=1.73 $Y=2.805 $X2=0 $Y2=0
cc_217 N_A_119_368#_c_302_n N_Y_c_341_n 0.0171805f $X=1.565 $Y=2.99 $X2=0 $Y2=0
cc_218 N_Y_c_332_n N_A_27_74#_c_379_n 0.00427071f $X=2.605 $Y=1.13 $X2=0 $Y2=0
cc_219 N_Y_c_333_n N_A_27_74#_c_379_n 0.00353683f $X=2.66 $Y=1.82 $X2=0 $Y2=0
cc_220 N_Y_M1005_d N_A_27_74#_c_381_n 0.00226551f $X=2.475 $Y=0.37 $X2=0 $Y2=0
cc_221 N_Y_c_374_p N_A_27_74#_c_381_n 0.0138835f $X=2.645 $Y=0.88 $X2=0 $Y2=0
cc_222 N_A_27_74#_c_376_n N_VGND_M1009_s 0.00256964f $X=1.125 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_223 N_A_27_74#_c_379_n N_VGND_M1011_s 0.00240632f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_224 N_A_27_74#_c_375_n N_VGND_c_435_n 0.0188012f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_225 N_A_27_74#_c_376_n N_VGND_c_435_n 0.0201026f $X=1.125 $Y=1.095 $X2=0
+ $Y2=0
cc_226 N_A_27_74#_c_378_n N_VGND_c_435_n 0.0179318f $X=1.21 $Y=0.515 $X2=0 $Y2=0
cc_227 N_A_27_74#_c_378_n N_VGND_c_436_n 0.018051f $X=1.21 $Y=0.515 $X2=0 $Y2=0
cc_228 N_A_27_74#_c_379_n N_VGND_c_436_n 0.0189333f $X=2.055 $Y=1.095 $X2=0
+ $Y2=0
cc_229 N_A_27_74#_c_380_n N_VGND_c_436_n 0.00697079f $X=2.18 $Y=0.52 $X2=0 $Y2=0
cc_230 N_A_27_74#_c_375_n N_VGND_c_437_n 0.0145639f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_231 N_A_27_74#_c_378_n N_VGND_c_438_n 0.0110391f $X=1.21 $Y=0.515 $X2=0 $Y2=0
cc_232 N_A_27_74#_c_380_n N_VGND_c_439_n 0.0111552f $X=2.18 $Y=0.52 $X2=0 $Y2=0
cc_233 N_A_27_74#_c_381_n N_VGND_c_439_n 0.0239026f $X=2.915 $Y=0.435 $X2=0
+ $Y2=0
cc_234 N_A_27_74#_c_383_n N_VGND_c_439_n 0.0146186f $X=3.08 $Y=0.515 $X2=0 $Y2=0
cc_235 N_A_27_74#_c_375_n N_VGND_c_440_n 0.0119984f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_236 N_A_27_74#_c_378_n N_VGND_c_440_n 0.00911606f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_237 N_A_27_74#_c_380_n N_VGND_c_440_n 0.00923333f $X=2.18 $Y=0.52 $X2=0 $Y2=0
cc_238 N_A_27_74#_c_381_n N_VGND_c_440_n 0.02025f $X=2.915 $Y=0.435 $X2=0 $Y2=0
cc_239 N_A_27_74#_c_383_n N_VGND_c_440_n 0.0120551f $X=3.08 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__a31oi_4.spice
* Created: Fri Aug 28 17:07:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a31oi_4.pex.spice"
.subckt sky130_fd_sc_ms__a31oi_4  VNB VPB A3 A2 A1 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1015 N_A_30_74#_M1015_d N_A3_M1015_g N_VGND_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1021 N_A_30_74#_M1021_d N_A3_M1021_g N_VGND_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1028 N_A_30_74#_M1021_d N_A3_M1028_g N_VGND_M1028_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1029 N_A_30_74#_M1029_d N_A3_M1029_g N_VGND_M1028_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.6
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1003 N_A_475_74#_M1003_d N_A2_M1003_g N_A_30_74#_M1029_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1073 AS=0.1036 PD=1.03 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333
+ SA=75002 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1012 N_A_475_74#_M1003_d N_A2_M1012_g N_A_30_74#_M1012_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1073 AS=0.1036 PD=1.03 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1022 N_A_475_74#_M1022_d N_A2_M1022_g N_A_30_74#_M1012_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75002.9 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1026 N_A_475_74#_M1022_d N_A2_M1026_g N_A_30_74#_M1026_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1554 AS=0.202325 PD=1.16 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75003.4 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A1_M1000_g N_A_475_74#_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.19805 AS=0.2109 PD=2.07 PS=1.31 NRD=0.804 NRS=23.508 M=1 R=4.93333
+ SA=75000.2 SB=75003.6 A=0.111 P=1.78 MULT=1
MM1005 N_Y_M1005_d N_A1_M1005_g N_A_475_74#_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=1.31 NRD=0 NRS=23.508 M=1 R=4.93333 SA=75000.9
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1024 N_Y_M1005_d N_A1_M1024_g N_A_475_74#_M1024_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.4
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1025 N_Y_M1025_d N_A1_M1025_g N_A_475_74#_M1024_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.8
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1023 N_Y_M1025_d N_B1_M1023_g N_VGND_M1023_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.40885 PD=1.09 PS=1.845 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1027 N_Y_M1027_d N_B1_M1027_g N_VGND_M1023_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.40885 PD=2.05 PS=1.845 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VPWR_M1008_d N_A3_M1008_g N_A_27_368#_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90007.8 A=0.2016 P=2.6 MULT=1
MM1009 N_VPWR_M1008_d N_A3_M1009_g N_A_27_368#_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90007.4 A=0.2016 P=2.6 MULT=1
MM1011 N_VPWR_M1011_d N_A3_M1011_g N_A_27_368#_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90006.9 A=0.2016 P=2.6 MULT=1
MM1013 N_VPWR_M1011_d N_A3_M1013_g N_A_27_368#_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90006.5 A=0.2016 P=2.6 MULT=1
MM1014 N_A_27_368#_M1013_s N_A2_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90006 A=0.2016 P=2.6 MULT=1
MM1016 N_A_27_368#_M1016_d N_A2_M1016_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.5
+ SB=90005.5 A=0.2016 P=2.6 MULT=1
MM1019 N_A_27_368#_M1016_d N_A2_M1019_g N_VPWR_M1019_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.9
+ SB=90005.1 A=0.2016 P=2.6 MULT=1
MM1020 N_A_27_368#_M1020_d N_A2_M1020_g N_VPWR_M1019_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90003.4
+ SB=90004.6 A=0.2016 P=2.6 MULT=1
MM1002 N_A_27_368#_M1020_d N_A1_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003.9
+ SB=90004.1 A=0.2016 P=2.6 MULT=1
MM1006 N_A_27_368#_M1006_d N_A1_M1006_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.448 AS=0.1792 PD=1.92 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.4
+ SB=90003.6 A=0.2016 P=2.6 MULT=1
MM1017 N_A_27_368#_M1006_d N_A1_M1017_g N_VPWR_M1017_s VPB PSHORT L=0.18 W=1.12
+ AD=0.448 AS=0.2072 PD=1.92 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90005.4
+ SB=90002.6 A=0.2016 P=2.6 MULT=1
MM1018 N_A_27_368#_M1018_d N_A1_M1018_g N_VPWR_M1017_s VPB PSHORT L=0.18 W=1.12
+ AD=0.168 AS=0.2072 PD=1.42 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90006
+ SB=90002 A=0.2016 P=2.6 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g N_A_27_368#_M1018_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1624 AS=0.168 PD=1.41 PS=1.42 NRD=2.6201 NRS=4.3931 M=1 R=6.22222
+ SA=90006.4 SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1001_d N_B1_M1004_g N_A_27_368#_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1624 AS=0.1512 PD=1.41 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90006.9
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1007 N_Y_M1007_d N_B1_M1007_g N_A_27_368#_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90007.4
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1010 N_Y_M1007_d N_B1_M1010_g N_A_27_368#_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90007.8
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX30_noxref VNB VPB NWDIODE A=16.7772 P=21.76
*
.include "sky130_fd_sc_ms__a31oi_4.pxi.spice"
*
.ends
*
*

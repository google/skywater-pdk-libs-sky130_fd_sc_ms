* File: sky130_fd_sc_ms__dfstp_2.pxi.spice
* Created: Fri Aug 28 17:24:11 2020
* 
x_PM_SKY130_FD_SC_MS__DFSTP_2%D N_D_c_246_n N_D_M1020_g N_D_M1031_g D D
+ N_D_c_248_n N_D_c_249_n N_D_c_253_n PM_SKY130_FD_SC_MS__DFSTP_2%D
x_PM_SKY130_FD_SC_MS__DFSTP_2%CLK N_CLK_M1033_g N_CLK_M1014_g CLK N_CLK_c_281_n
+ N_CLK_c_282_n PM_SKY130_FD_SC_MS__DFSTP_2%CLK
x_PM_SKY130_FD_SC_MS__DFSTP_2%A_398_74# N_A_398_74#_M1015_d N_A_398_74#_M1017_d
+ N_A_398_74#_c_318_n N_A_398_74#_c_337_n N_A_398_74#_M1023_g
+ N_A_398_74#_c_319_n N_A_398_74#_c_320_n N_A_398_74#_M1012_g
+ N_A_398_74#_M1001_g N_A_398_74#_M1010_g N_A_398_74#_c_342_n
+ N_A_398_74#_c_322_n N_A_398_74#_c_440_p N_A_398_74#_c_323_n
+ N_A_398_74#_c_324_n N_A_398_74#_c_343_n N_A_398_74#_c_344_n
+ N_A_398_74#_c_325_n N_A_398_74#_c_326_n N_A_398_74#_c_347_n
+ N_A_398_74#_c_348_n N_A_398_74#_c_349_n N_A_398_74#_c_350_n
+ N_A_398_74#_c_351_n N_A_398_74#_c_352_n N_A_398_74#_c_382_p
+ N_A_398_74#_c_418_p N_A_398_74#_c_327_n N_A_398_74#_c_328_n
+ N_A_398_74#_c_329_n N_A_398_74#_c_330_n N_A_398_74#_c_331_n
+ N_A_398_74#_c_332_n N_A_398_74#_c_355_n N_A_398_74#_c_333_n
+ N_A_398_74#_c_334_n N_A_398_74#_c_356_n N_A_398_74#_c_335_n
+ PM_SKY130_FD_SC_MS__DFSTP_2%A_398_74#
x_PM_SKY130_FD_SC_MS__DFSTP_2%A_767_384# N_A_767_384#_M1002_s
+ N_A_767_384#_M1009_d N_A_767_384#_M1032_g N_A_767_384#_c_588_n
+ N_A_767_384#_c_589_n N_A_767_384#_c_583_n N_A_767_384#_M1024_g
+ N_A_767_384#_c_590_n N_A_767_384#_c_591_n N_A_767_384#_c_584_n
+ N_A_767_384#_c_592_n N_A_767_384#_c_593_n N_A_767_384#_c_585_n
+ N_A_767_384#_c_586_n PM_SKY130_FD_SC_MS__DFSTP_2%A_767_384#
x_PM_SKY130_FD_SC_MS__DFSTP_2%A_612_74# N_A_612_74#_M1018_d N_A_612_74#_M1023_d
+ N_A_612_74#_M1009_g N_A_612_74#_M1002_g N_A_612_74#_M1011_g
+ N_A_612_74#_M1000_g N_A_612_74#_c_664_n N_A_612_74#_c_665_n
+ N_A_612_74#_c_666_n N_A_612_74#_c_667_n N_A_612_74#_c_668_n
+ N_A_612_74#_c_677_n N_A_612_74#_c_669_n N_A_612_74#_c_670_n
+ N_A_612_74#_c_671_n N_A_612_74#_c_679_n N_A_612_74#_c_672_n
+ N_A_612_74#_c_673_n N_A_612_74#_c_674_n PM_SKY130_FD_SC_MS__DFSTP_2%A_612_74#
x_PM_SKY130_FD_SC_MS__DFSTP_2%SET_B N_SET_B_M1016_g N_SET_B_M1022_g
+ N_SET_B_M1004_g N_SET_B_M1007_g N_SET_B_c_796_n N_SET_B_c_803_n
+ N_SET_B_c_804_n N_SET_B_c_805_n N_SET_B_c_806_n SET_B N_SET_B_c_797_n
+ N_SET_B_c_798_n N_SET_B_c_809_n PM_SKY130_FD_SC_MS__DFSTP_2%SET_B
x_PM_SKY130_FD_SC_MS__DFSTP_2%A_225_74# N_A_225_74#_M1033_s N_A_225_74#_M1014_s
+ N_A_225_74#_M1015_g N_A_225_74#_M1017_g N_A_225_74#_c_918_n
+ N_A_225_74#_c_932_n N_A_225_74#_c_919_n N_A_225_74#_c_920_n
+ N_A_225_74#_c_933_n N_A_225_74#_c_934_n N_A_225_74#_M1018_g
+ N_A_225_74#_M1021_g N_A_225_74#_c_936_n N_A_225_74#_M1003_g
+ N_A_225_74#_c_922_n N_A_225_74#_c_923_n N_A_225_74#_M1008_g
+ N_A_225_74#_c_925_n N_A_225_74#_c_926_n N_A_225_74#_c_927_n
+ N_A_225_74#_c_943_n N_A_225_74#_c_928_n N_A_225_74#_c_945_n
+ N_A_225_74#_c_946_n N_A_225_74#_c_947_n N_A_225_74#_c_929_n
+ N_A_225_74#_c_930_n N_A_225_74#_c_949_n PM_SKY130_FD_SC_MS__DFSTP_2%A_225_74#
x_PM_SKY130_FD_SC_MS__DFSTP_2%A_1566_92# N_A_1566_92#_M1027_d
+ N_A_1566_92#_M1019_d N_A_1566_92#_M1030_g N_A_1566_92#_M1028_g
+ N_A_1566_92#_c_1103_n N_A_1566_92#_c_1112_n N_A_1566_92#_c_1104_n
+ N_A_1566_92#_c_1105_n N_A_1566_92#_c_1106_n N_A_1566_92#_c_1107_n
+ N_A_1566_92#_c_1108_n N_A_1566_92#_c_1109_n N_A_1566_92#_c_1110_n
+ N_A_1566_92#_c_1115_n PM_SKY130_FD_SC_MS__DFSTP_2%A_1566_92#
x_PM_SKY130_FD_SC_MS__DFSTP_2%A_1356_74# N_A_1356_74#_M1001_d
+ N_A_1356_74#_M1003_d N_A_1356_74#_M1007_d N_A_1356_74#_M1027_g
+ N_A_1356_74#_M1019_g N_A_1356_74#_c_1182_n N_A_1356_74#_M1013_g
+ N_A_1356_74#_c_1191_n N_A_1356_74#_M1006_g N_A_1356_74#_c_1184_n
+ N_A_1356_74#_c_1193_n N_A_1356_74#_c_1185_n N_A_1356_74#_c_1195_n
+ N_A_1356_74#_c_1186_n N_A_1356_74#_c_1216_n N_A_1356_74#_c_1196_n
+ N_A_1356_74#_c_1197_n N_A_1356_74#_c_1198_n N_A_1356_74#_c_1199_n
+ N_A_1356_74#_c_1187_n N_A_1356_74#_c_1201_n N_A_1356_74#_c_1188_n
+ N_A_1356_74#_c_1202_n N_A_1356_74#_c_1227_n N_A_1356_74#_c_1203_n
+ PM_SKY130_FD_SC_MS__DFSTP_2%A_1356_74#
x_PM_SKY130_FD_SC_MS__DFSTP_2%A_2022_94# N_A_2022_94#_M1013_s
+ N_A_2022_94#_M1006_s N_A_2022_94#_M1026_g N_A_2022_94#_M1005_g
+ N_A_2022_94#_M1025_g N_A_2022_94#_M1029_g N_A_2022_94#_c_1339_n
+ N_A_2022_94#_c_1345_n N_A_2022_94#_c_1340_n N_A_2022_94#_c_1341_n
+ N_A_2022_94#_c_1342_n PM_SKY130_FD_SC_MS__DFSTP_2%A_2022_94#
x_PM_SKY130_FD_SC_MS__DFSTP_2%A_27_74# N_A_27_74#_M1031_s N_A_27_74#_M1018_s
+ N_A_27_74#_M1020_s N_A_27_74#_M1023_s N_A_27_74#_c_1405_n N_A_27_74#_c_1410_n
+ N_A_27_74#_c_1411_n N_A_27_74#_c_1412_n N_A_27_74#_c_1406_n
+ N_A_27_74#_c_1407_n N_A_27_74#_c_1414_n N_A_27_74#_c_1459_n
+ N_A_27_74#_c_1408_n PM_SKY130_FD_SC_MS__DFSTP_2%A_27_74#
x_PM_SKY130_FD_SC_MS__DFSTP_2%VPWR N_VPWR_M1020_d N_VPWR_M1014_d N_VPWR_M1032_d
+ N_VPWR_M1016_d N_VPWR_M1028_d N_VPWR_M1019_s N_VPWR_M1006_d N_VPWR_M1029_s
+ N_VPWR_c_1476_n N_VPWR_c_1477_n N_VPWR_c_1478_n N_VPWR_c_1479_n
+ N_VPWR_c_1480_n N_VPWR_c_1481_n N_VPWR_c_1482_n N_VPWR_c_1483_n
+ N_VPWR_c_1484_n N_VPWR_c_1485_n N_VPWR_c_1486_n N_VPWR_c_1487_n VPWR
+ N_VPWR_c_1488_n N_VPWR_c_1489_n N_VPWR_c_1490_n N_VPWR_c_1491_n
+ N_VPWR_c_1492_n N_VPWR_c_1493_n N_VPWR_c_1494_n N_VPWR_c_1495_n
+ N_VPWR_c_1496_n N_VPWR_c_1497_n N_VPWR_c_1498_n N_VPWR_c_1499_n
+ N_VPWR_c_1500_n N_VPWR_c_1475_n PM_SKY130_FD_SC_MS__DFSTP_2%VPWR
x_PM_SKY130_FD_SC_MS__DFSTP_2%Q N_Q_M1005_s N_Q_M1026_d N_Q_c_1629_n
+ N_Q_c_1632_n N_Q_c_1630_n N_Q_c_1631_n Q Q N_Q_c_1635_n
+ PM_SKY130_FD_SC_MS__DFSTP_2%Q
x_PM_SKY130_FD_SC_MS__DFSTP_2%VGND N_VGND_M1031_d N_VGND_M1033_d N_VGND_M1024_d
+ N_VGND_M1022_d N_VGND_M1004_d N_VGND_M1013_d N_VGND_M1025_d N_VGND_c_1668_n
+ N_VGND_c_1669_n N_VGND_c_1670_n N_VGND_c_1671_n N_VGND_c_1672_n
+ N_VGND_c_1673_n N_VGND_c_1674_n N_VGND_c_1675_n VGND N_VGND_c_1676_n
+ N_VGND_c_1677_n N_VGND_c_1678_n N_VGND_c_1679_n N_VGND_c_1680_n
+ N_VGND_c_1681_n N_VGND_c_1682_n N_VGND_c_1683_n N_VGND_c_1684_n
+ N_VGND_c_1685_n N_VGND_c_1686_n N_VGND_c_1687_n
+ PM_SKY130_FD_SC_MS__DFSTP_2%VGND
cc_1 VNB N_D_c_246_n 0.0447809f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.795
cc_2 VNB N_D_M1031_g 0.0288784f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_3 VNB N_D_c_248_n 0.025337f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_4 VNB N_D_c_249_n 0.00269121f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_5 VNB N_CLK_M1014_g 0.00385449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB CLK 0.00873773f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_7 VNB N_CLK_c_281_n 0.0322418f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_8 VNB N_CLK_c_282_n 0.019964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_398_74#_c_318_n 0.0168103f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.98
cc_10 VNB N_A_398_74#_c_319_n 0.0368422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_398_74#_c_320_n 0.0112016f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_12 VNB N_A_398_74#_M1012_g 0.0507397f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_13 VNB N_A_398_74#_c_322_n 0.00150841f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_14 VNB N_A_398_74#_c_323_n 0.0158463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_398_74#_c_324_n 0.00264685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_398_74#_c_325_n 0.00190286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_398_74#_c_326_n 0.0012865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_398_74#_c_327_n 0.00247322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_398_74#_c_328_n 0.00213614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_398_74#_c_329_n 0.0230647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_398_74#_c_330_n 0.00190332f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_398_74#_c_331_n 0.0153419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_398_74#_c_332_n 0.00680136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_398_74#_c_333_n 0.00734472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_398_74#_c_334_n 0.031744f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_398_74#_c_335_n 0.0197653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_767_384#_c_583_n 0.0195194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_767_384#_c_584_n 0.0240574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_767_384#_c_585_n 0.0224227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_767_384#_c_586_n 0.0535767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_612_74#_M1009_g 0.00366225f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_32 VNB N_A_612_74#_M1002_g 0.0241071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_612_74#_M1000_g 0.0253106f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_34 VNB N_A_612_74#_c_664_n 0.00685615f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.295
cc_35 VNB N_A_612_74#_c_665_n 0.0205132f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_36 VNB N_A_612_74#_c_666_n 0.00415803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_612_74#_c_667_n 0.00363794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_612_74#_c_668_n 0.00239084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_612_74#_c_669_n 0.00313488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_612_74#_c_670_n 0.00482349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_612_74#_c_671_n 0.00993512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_612_74#_c_672_n 0.0192723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_612_74#_c_673_n 0.0304134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_612_74#_c_674_n 0.0332086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_SET_B_M1022_g 0.0410395f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.98
cc_46 VNB N_SET_B_M1004_g 0.04772f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_47 VNB N_SET_B_c_796_n 9.90083e-19 $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.825
cc_48 VNB N_SET_B_c_797_n 0.0178127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_SET_B_c_798_n 0.00389433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_225_74#_M1015_g 0.0224523f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_51 VNB N_A_225_74#_c_918_n 0.00808021f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_52 VNB N_A_225_74#_c_919_n 0.0340583f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.825
cc_53 VNB N_A_225_74#_c_920_n 0.010226f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_54 VNB N_A_225_74#_M1018_g 0.0265626f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.295
cc_55 VNB N_A_225_74#_c_922_n 0.0106772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_225_74#_c_923_n 0.00106815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_225_74#_M1008_g 0.0502374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_225_74#_c_925_n 0.0123708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_225_74#_c_926_n 0.0195044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_225_74#_c_927_n 0.00971956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_225_74#_c_928_n 0.0104758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_225_74#_c_929_n 0.00365457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_225_74#_c_930_n 0.0133435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1566_92#_c_1103_n 0.0188877f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_65 VNB N_A_1566_92#_c_1104_n 0.0161793f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.825
cc_66 VNB N_A_1566_92#_c_1105_n 0.0283476f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.99
cc_67 VNB N_A_1566_92#_c_1106_n 0.0447681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1566_92#_c_1107_n 0.00788489f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.295
cc_69 VNB N_A_1566_92#_c_1108_n 0.00499052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1566_92#_c_1109_n 0.00759688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1566_92#_c_1110_n 0.00570228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1356_74#_M1027_g 0.0604445f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_73 VNB N_A_1356_74#_c_1182_n 0.0264413f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.98
cc_74 VNB N_A_1356_74#_M1013_g 0.0460006f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.99
cc_75 VNB N_A_1356_74#_c_1184_n 0.0107945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1356_74#_c_1185_n 0.00337811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1356_74#_c_1186_n 0.00606384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1356_74#_c_1187_n 0.00342147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1356_74#_c_1188_n 0.00446853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_2022_94#_M1026_g 0.00167809f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_81 VNB N_A_2022_94#_M1005_g 0.0229692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_2022_94#_M1025_g 0.0260335f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_83 VNB N_A_2022_94#_M1029_g 0.00231818f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_84 VNB N_A_2022_94#_c_1339_n 0.0125258f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.295
cc_85 VNB N_A_2022_94#_c_1340_n 0.0084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_2022_94#_c_1341_n 0.00309584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_2022_94#_c_1342_n 0.0647641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_27_74#_c_1405_n 0.0420755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_27_74#_c_1406_n 0.00574528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_27_74#_c_1407_n 0.0137638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_27_74#_c_1408_n 0.00619147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VPWR_c_1475_n 0.502022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_Q_c_1629_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_94 VNB N_Q_c_1630_n 0.00143777f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_95 VNB N_Q_c_1631_n 0.00457514f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_96 VNB N_VGND_c_1668_n 0.00619735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1669_n 0.0224525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1670_n 0.00559476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1671_n 0.0163103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1672_n 0.0214836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1673_n 0.0164768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1674_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1675_n 0.0505491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1676_n 0.0175546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1677_n 0.0636081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1678_n 0.0313742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1679_n 0.113496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1680_n 0.0357284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1681_n 0.0195351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1682_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1683_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1684_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1685_n 0.0112736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1686_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1687_n 0.696385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VPB N_D_c_246_n 0.0126737f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.795
cc_117 VPB N_D_M1020_g 0.0635978f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.75
cc_118 VPB N_D_c_249_n 0.00207792f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_119 VPB N_D_c_253_n 0.0244074f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_120 VPB N_CLK_M1014_g 0.0238474f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_398_74#_c_318_n 0.00525997f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.98
cc_122 VPB N_A_398_74#_c_337_n 0.0132143f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_123 VPB N_A_398_74#_M1023_g 0.0253475f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_124 VPB N_A_398_74#_c_319_n 0.0253435f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_398_74#_c_320_n 0.00803075f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.145
cc_126 VPB N_A_398_74#_M1010_g 0.0248072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_398_74#_c_342_n 0.0176902f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_398_74#_c_343_n 0.0220334f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_398_74#_c_344_n 0.00294918f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_398_74#_c_325_n 0.00207712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_398_74#_c_326_n 0.00587279f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_398_74#_c_347_n 0.0033448f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_398_74#_c_348_n 0.00842907f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_398_74#_c_349_n 0.00469668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_398_74#_c_350_n 0.015777f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_398_74#_c_351_n 0.00428736f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_398_74#_c_352_n 0.00229189f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_398_74#_c_328_n 0.00419354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_398_74#_c_331_n 0.0132977f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_398_74#_c_355_n 2.604e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_398_74#_c_356_n 0.033949f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_767_384#_M1032_g 0.0278706f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_143 VPB N_A_767_384#_c_588_n 0.0150258f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_144 VPB N_A_767_384#_c_589_n 0.0121391f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_145 VPB N_A_767_384#_c_590_n 0.0134053f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_146 VPB N_A_767_384#_c_591_n 0.0357903f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_147 VPB N_A_767_384#_c_592_n 0.00144661f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_767_384#_c_593_n 0.00167787f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_767_384#_c_585_n 0.00840486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_612_74#_M1009_g 0.0516324f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_151 VPB N_A_612_74#_M1011_g 0.0225169f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_152 VPB N_A_612_74#_c_677_n 0.00494346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_612_74#_c_669_n 0.00808184f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_612_74#_c_679_n 0.00253708f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_612_74#_c_672_n 0.00168218f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_612_74#_c_674_n 0.0106991f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_SET_B_M1016_g 0.0209795f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.99
cc_158 VPB N_SET_B_M1022_g 0.0116829f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.98
cc_159 VPB N_SET_B_M1007_g 0.0399977f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.145
cc_160 VPB N_SET_B_c_796_n 0.0229134f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.825
cc_161 VPB N_SET_B_c_803_n 0.0160157f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_162 VPB N_SET_B_c_804_n 0.0178302f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_163 VPB N_SET_B_c_805_n 4.31814e-19 $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.99
cc_164 VPB N_SET_B_c_806_n 0.0043956f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.295
cc_165 VPB SET_B 0.00404524f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_166 VPB N_SET_B_c_798_n 0.00416461f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_SET_B_c_809_n 0.0349351f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_225_74#_M1017_g 0.0197043f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_225_74#_c_932_n 0.0744311f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_170 VPB N_A_225_74#_c_933_n 0.0560671f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_171 VPB N_A_225_74#_c_934_n 0.0125859f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.99
cc_172 VPB N_A_225_74#_M1021_g 0.0379581f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_173 VPB N_A_225_74#_c_936_n 0.233439f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_225_74#_M1003_g 0.0188865f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_225_74#_c_922_n 0.0399382f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_225_74#_c_923_n 0.00891769f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_225_74#_c_925_n 0.00170265f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_225_74#_c_926_n 0.00577555f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_225_74#_c_927_n 5.35904e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_225_74#_c_943_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_225_74#_c_928_n 0.00240536f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_225_74#_c_945_n 0.0058961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_225_74#_c_946_n 0.00539283f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_225_74#_c_947_n 0.00446037f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_225_74#_c_929_n 5.33031e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_225_74#_c_949_n 7.70291e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_1566_92#_M1028_g 0.0350904f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_188 VPB N_A_1566_92#_c_1112_n 0.00129748f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_189 VPB N_A_1566_92#_c_1105_n 0.0232163f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.99
cc_190 VPB N_A_1566_92#_c_1109_n 0.0229941f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_1566_92#_c_1115_n 0.0160359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_1356_74#_M1019_g 0.0353734f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_193 VPB N_A_1356_74#_c_1182_n 0.0312876f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_194 VPB N_A_1356_74#_c_1191_n 0.0191262f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_1356_74#_c_1184_n 0.0076044f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_1356_74#_c_1193_n 0.0298932f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_1356_74#_c_1185_n 0.00469003f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_1356_74#_c_1195_n 0.00201305f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_1356_74#_c_1196_n 0.00335263f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_1356_74#_c_1197_n 0.00291284f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_1356_74#_c_1198_n 0.00680625f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_1356_74#_c_1199_n 0.0162059f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_1356_74#_c_1187_n 4.98981e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_1356_74#_c_1201_n 0.0280862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_1356_74#_c_1202_n 0.00518849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_1356_74#_c_1203_n 0.00856327f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_2022_94#_M1026_g 0.0243722f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_208 VPB N_A_2022_94#_M1029_g 0.0273866f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_209 VPB N_A_2022_94#_c_1345_n 0.0135438f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_210 VPB N_A_27_74#_c_1405_n 0.0250181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_27_74#_c_1410_n 0.0274742f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_212 VPB N_A_27_74#_c_1411_n 0.0257471f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.825
cc_213 VPB N_A_27_74#_c_1412_n 0.0158417f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_214 VPB N_A_27_74#_c_1406_n 0.00273955f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_27_74#_c_1414_n 0.0109364f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_216 VPB N_VPWR_c_1476_n 0.0169911f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_217 VPB N_VPWR_c_1477_n 0.0065563f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1478_n 0.00509177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1479_n 0.00662535f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1480_n 0.00650405f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1481_n 0.0097693f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1482_n 0.0102774f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1483_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1484_n 0.0637781f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1485_n 0.0055215f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1486_n 0.0549518f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1487_n 0.00612813f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1488_n 0.0180274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1489_n 0.0215753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1490_n 0.0523685f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1491_n 0.0384523f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1492_n 0.01948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1493_n 0.0342956f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1494_n 0.0180566f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1495_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1496_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1497_n 0.00223285f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1498_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1499_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1500_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1475_n 0.120727f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_Q_c_1632_n 0.00229073f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_Q_c_1630_n 0.0010488f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_244 VPB Q 0.00365809f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.825
cc_245 VPB N_Q_c_1635_n 0.0030239f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.99
cc_246 N_D_c_246_n N_CLK_M1014_g 0.00408937f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_247 N_D_c_246_n N_CLK_c_281_n 0.00572583f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_248 N_D_c_248_n N_CLK_c_282_n 0.00223659f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_249 N_D_c_246_n N_A_225_74#_c_928_n 0.003576f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_250 N_D_c_246_n N_A_225_74#_c_946_n 0.00298111f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_251 N_D_M1020_g N_A_225_74#_c_946_n 9.40485e-19 $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_252 N_D_c_249_n N_A_225_74#_c_946_n 0.0224944f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_253 N_D_M1031_g N_A_225_74#_c_930_n 0.00721478f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_254 N_D_c_248_n N_A_225_74#_c_930_n 0.003576f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_255 N_D_c_249_n N_A_225_74#_c_930_n 0.0556869f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_256 N_D_M1031_g N_A_27_74#_c_1405_n 0.00743437f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_257 N_D_c_248_n N_A_27_74#_c_1405_n 0.0320429f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_258 N_D_c_249_n N_A_27_74#_c_1405_n 0.0697394f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_259 N_D_M1020_g N_A_27_74#_c_1410_n 0.0083684f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_260 N_D_M1020_g N_A_27_74#_c_1411_n 0.0218367f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_261 N_D_c_249_n N_A_27_74#_c_1411_n 0.0227191f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_262 N_D_c_253_n N_A_27_74#_c_1411_n 0.00140505f $X=0.64 $Y=1.825 $X2=0 $Y2=0
cc_263 N_D_M1020_g N_VPWR_c_1476_n 0.0148304f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_264 N_D_M1020_g N_VPWR_c_1488_n 0.00460063f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_265 N_D_M1020_g N_VPWR_c_1475_n 0.00912296f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_266 N_D_M1031_g N_VGND_c_1668_n 0.0140619f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_267 N_D_c_248_n N_VGND_c_1668_n 0.00150697f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_268 N_D_c_249_n N_VGND_c_1668_n 0.0158023f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_269 N_D_M1031_g N_VGND_c_1676_n 0.00383152f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_270 N_D_M1031_g N_VGND_c_1687_n 0.00761198f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_271 CLK N_A_225_74#_M1015_g 0.00369616f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_272 N_CLK_c_281_n N_A_225_74#_M1015_g 0.0210236f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_273 N_CLK_c_282_n N_A_225_74#_M1015_g 0.0131399f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_274 N_CLK_M1014_g N_A_225_74#_M1017_g 0.0488038f $X=1.515 $Y=2.35 $X2=0 $Y2=0
cc_275 N_CLK_M1014_g N_A_225_74#_c_925_n 0.00479904f $X=1.515 $Y=2.35 $X2=0
+ $Y2=0
cc_276 N_CLK_M1014_g N_A_225_74#_c_928_n 0.00354737f $X=1.515 $Y=2.35 $X2=0
+ $Y2=0
cc_277 CLK N_A_225_74#_c_928_n 0.0286813f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_278 N_CLK_c_281_n N_A_225_74#_c_928_n 0.00297156f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_279 N_CLK_c_282_n N_A_225_74#_c_928_n 0.00321998f $X=1.465 $Y=1.22 $X2=0
+ $Y2=0
cc_280 N_CLK_c_281_n N_A_225_74#_c_945_n 0.00313913f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_281 N_CLK_M1014_g N_A_225_74#_c_947_n 0.009076f $X=1.515 $Y=2.35 $X2=0 $Y2=0
cc_282 N_CLK_c_281_n N_A_225_74#_c_947_n 5.60514e-19 $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_283 N_CLK_M1014_g N_A_225_74#_c_929_n 9.11681e-19 $X=1.515 $Y=2.35 $X2=0
+ $Y2=0
cc_284 CLK N_A_225_74#_c_929_n 0.0203335f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_285 N_CLK_c_281_n N_A_225_74#_c_929_n 2.00661e-19 $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_286 CLK N_A_225_74#_c_930_n 0.00762435f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_287 N_CLK_c_281_n N_A_225_74#_c_930_n 0.00114511f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_288 N_CLK_c_282_n N_A_225_74#_c_930_n 0.00791767f $X=1.465 $Y=1.22 $X2=0
+ $Y2=0
cc_289 N_CLK_M1014_g N_A_225_74#_c_949_n 0.00508679f $X=1.515 $Y=2.35 $X2=0
+ $Y2=0
cc_290 CLK N_A_225_74#_c_949_n 0.0352423f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_291 N_CLK_M1014_g N_A_27_74#_c_1411_n 0.0177479f $X=1.515 $Y=2.35 $X2=0 $Y2=0
cc_292 CLK N_A_27_74#_c_1406_n 0.00323107f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_293 N_CLK_M1014_g N_VPWR_c_1476_n 0.0132363f $X=1.515 $Y=2.35 $X2=0 $Y2=0
cc_294 N_CLK_M1014_g N_VPWR_c_1477_n 0.025074f $X=1.515 $Y=2.35 $X2=0 $Y2=0
cc_295 N_CLK_M1014_g N_VPWR_c_1489_n 0.00540231f $X=1.515 $Y=2.35 $X2=0 $Y2=0
cc_296 N_CLK_M1014_g N_VPWR_c_1475_n 0.00533457f $X=1.515 $Y=2.35 $X2=0 $Y2=0
cc_297 N_CLK_c_282_n N_VGND_c_1668_n 0.00295547f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_298 N_CLK_c_282_n N_VGND_c_1669_n 0.00434272f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_299 CLK N_VGND_c_1670_n 0.013855f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_300 N_CLK_c_282_n N_VGND_c_1670_n 0.00294833f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_301 N_CLK_c_282_n N_VGND_c_1687_n 0.00825381f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_302 N_A_398_74#_c_326_n N_A_767_384#_M1032_g 0.0101657f $X=3.77 $Y=1.545
+ $X2=0 $Y2=0
cc_303 N_A_398_74#_c_347_n N_A_767_384#_M1032_g 0.00222549f $X=3.71 $Y=2.89
+ $X2=0 $Y2=0
cc_304 N_A_398_74#_c_348_n N_A_767_384#_M1032_g 0.0111646f $X=4.745 $Y=2.325
+ $X2=0 $Y2=0
cc_305 N_A_398_74#_c_355_n N_A_767_384#_M1032_g 0.00445046f $X=3.77 $Y=2.325
+ $X2=0 $Y2=0
cc_306 N_A_398_74#_c_348_n N_A_767_384#_c_588_n 0.0138336f $X=4.745 $Y=2.325
+ $X2=0 $Y2=0
cc_307 N_A_398_74#_c_320_n N_A_767_384#_c_589_n 0.0067588f $X=3.83 $Y=1.38 $X2=0
+ $Y2=0
cc_308 N_A_398_74#_c_342_n N_A_767_384#_c_589_n 0.00118696f $X=2.95 $Y=2.05
+ $X2=0 $Y2=0
cc_309 N_A_398_74#_c_326_n N_A_767_384#_c_589_n 0.00714225f $X=3.77 $Y=1.545
+ $X2=0 $Y2=0
cc_310 N_A_398_74#_M1012_g N_A_767_384#_c_583_n 0.043019f $X=3.83 $Y=0.58 $X2=0
+ $Y2=0
cc_311 N_A_398_74#_c_326_n N_A_767_384#_c_590_n 0.0165446f $X=3.77 $Y=1.545
+ $X2=0 $Y2=0
cc_312 N_A_398_74#_c_348_n N_A_767_384#_c_590_n 0.0544703f $X=4.745 $Y=2.325
+ $X2=0 $Y2=0
cc_313 N_A_398_74#_c_326_n N_A_767_384#_c_591_n 0.00117498f $X=3.77 $Y=1.545
+ $X2=0 $Y2=0
cc_314 N_A_398_74#_M1012_g N_A_767_384#_c_584_n 6.56857e-19 $X=3.83 $Y=0.58
+ $X2=0 $Y2=0
cc_315 N_A_398_74#_c_349_n N_A_767_384#_c_592_n 0.0119623f $X=4.83 $Y=2.89 $X2=0
+ $Y2=0
cc_316 N_A_398_74#_c_350_n N_A_767_384#_c_592_n 0.0203683f $X=5.52 $Y=2.975
+ $X2=0 $Y2=0
cc_317 N_A_398_74#_c_352_n N_A_767_384#_c_592_n 0.00852554f $X=5.605 $Y=2.89
+ $X2=0 $Y2=0
cc_318 N_A_398_74#_c_348_n N_A_767_384#_c_593_n 0.00778909f $X=4.745 $Y=2.325
+ $X2=0 $Y2=0
cc_319 N_A_398_74#_c_320_n N_A_767_384#_c_585_n 0.00809956f $X=3.83 $Y=1.38
+ $X2=0 $Y2=0
cc_320 N_A_398_74#_c_326_n N_A_767_384#_c_585_n 0.00165073f $X=3.77 $Y=1.545
+ $X2=0 $Y2=0
cc_321 N_A_398_74#_M1012_g N_A_767_384#_c_586_n 0.00534415f $X=3.83 $Y=0.58
+ $X2=0 $Y2=0
cc_322 N_A_398_74#_c_348_n N_A_612_74#_M1009_g 0.00363124f $X=4.745 $Y=2.325
+ $X2=0 $Y2=0
cc_323 N_A_398_74#_c_349_n N_A_612_74#_M1009_g 0.00956386f $X=4.83 $Y=2.89 $X2=0
+ $Y2=0
cc_324 N_A_398_74#_c_350_n N_A_612_74#_M1009_g 0.00373127f $X=5.52 $Y=2.975
+ $X2=0 $Y2=0
cc_325 N_A_398_74#_c_352_n N_A_612_74#_M1009_g 4.25499e-19 $X=5.605 $Y=2.89
+ $X2=0 $Y2=0
cc_326 N_A_398_74#_c_352_n N_A_612_74#_M1011_g 0.00299314f $X=5.605 $Y=2.89
+ $X2=0 $Y2=0
cc_327 N_A_398_74#_c_382_p N_A_612_74#_M1011_g 0.0125554f $X=6.415 $Y=2.405
+ $X2=0 $Y2=0
cc_328 N_A_398_74#_c_328_n N_A_612_74#_M1011_g 0.0144679f $X=6.5 $Y=2.32 $X2=0
+ $Y2=0
cc_329 N_A_398_74#_c_327_n N_A_612_74#_M1000_g 0.00450375f $X=6.5 $Y=1.12 $X2=0
+ $Y2=0
cc_330 N_A_398_74#_c_330_n N_A_612_74#_M1000_g 0.0010322f $X=6.585 $Y=0.365
+ $X2=0 $Y2=0
cc_331 N_A_398_74#_c_333_n N_A_612_74#_M1000_g 0.00497904f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_332 N_A_398_74#_c_335_n N_A_612_74#_M1000_g 0.0283335f $X=6.795 $Y=1.12 $X2=0
+ $Y2=0
cc_333 N_A_398_74#_M1012_g N_A_612_74#_c_664_n 0.0143447f $X=3.83 $Y=0.58 $X2=0
+ $Y2=0
cc_334 N_A_398_74#_c_332_n N_A_612_74#_c_664_n 0.0343771f $X=2.95 $Y=1.38 $X2=0
+ $Y2=0
cc_335 N_A_398_74#_c_319_n N_A_612_74#_c_665_n 0.0013004f $X=3.755 $Y=1.545
+ $X2=0 $Y2=0
cc_336 N_A_398_74#_c_320_n N_A_612_74#_c_665_n 8.52337e-19 $X=3.83 $Y=1.38 $X2=0
+ $Y2=0
cc_337 N_A_398_74#_M1012_g N_A_612_74#_c_665_n 0.0169962f $X=3.83 $Y=0.58 $X2=0
+ $Y2=0
cc_338 N_A_398_74#_c_326_n N_A_612_74#_c_665_n 0.0224126f $X=3.77 $Y=1.545 $X2=0
+ $Y2=0
cc_339 N_A_398_74#_M1012_g N_A_612_74#_c_666_n 0.0020456f $X=3.83 $Y=0.58 $X2=0
+ $Y2=0
cc_340 N_A_398_74#_c_326_n N_A_612_74#_c_666_n 0.00145075f $X=3.77 $Y=1.545
+ $X2=0 $Y2=0
cc_341 N_A_398_74#_c_320_n N_A_612_74#_c_667_n 0.00187189f $X=3.83 $Y=1.38 $X2=0
+ $Y2=0
cc_342 N_A_398_74#_c_326_n N_A_612_74#_c_667_n 0.0142106f $X=3.77 $Y=1.545 $X2=0
+ $Y2=0
cc_343 N_A_398_74#_c_348_n N_A_612_74#_c_667_n 0.00453594f $X=4.745 $Y=2.325
+ $X2=0 $Y2=0
cc_344 N_A_398_74#_M1023_g N_A_612_74#_c_677_n 5.0381e-19 $X=3.005 $Y=2.49 $X2=0
+ $Y2=0
cc_345 N_A_398_74#_c_319_n N_A_612_74#_c_677_n 0.00478473f $X=3.755 $Y=1.545
+ $X2=0 $Y2=0
cc_346 N_A_398_74#_c_343_n N_A_612_74#_c_677_n 0.0260867f $X=3.625 $Y=2.975
+ $X2=0 $Y2=0
cc_347 N_A_398_74#_c_347_n N_A_612_74#_c_677_n 0.0124001f $X=3.71 $Y=2.89 $X2=0
+ $Y2=0
cc_348 N_A_398_74#_c_337_n N_A_612_74#_c_669_n 0.00608994f $X=2.95 $Y=1.885
+ $X2=0 $Y2=0
cc_349 N_A_398_74#_M1023_g N_A_612_74#_c_669_n 0.00355454f $X=3.005 $Y=2.49
+ $X2=0 $Y2=0
cc_350 N_A_398_74#_c_319_n N_A_612_74#_c_669_n 0.0222071f $X=3.755 $Y=1.545
+ $X2=0 $Y2=0
cc_351 N_A_398_74#_M1012_g N_A_612_74#_c_669_n 0.00339481f $X=3.83 $Y=0.58 $X2=0
+ $Y2=0
cc_352 N_A_398_74#_c_326_n N_A_612_74#_c_669_n 0.0645348f $X=3.77 $Y=1.545 $X2=0
+ $Y2=0
cc_353 N_A_398_74#_c_332_n N_A_612_74#_c_669_n 0.0617327f $X=2.95 $Y=1.38 $X2=0
+ $Y2=0
cc_354 N_A_398_74#_c_355_n N_A_612_74#_c_669_n 0.0081461f $X=3.77 $Y=2.325 $X2=0
+ $Y2=0
cc_355 N_A_398_74#_c_319_n N_A_612_74#_c_670_n 0.00711061f $X=3.755 $Y=1.545
+ $X2=0 $Y2=0
cc_356 N_A_398_74#_c_332_n N_A_612_74#_c_670_n 0.0143569f $X=2.95 $Y=1.38 $X2=0
+ $Y2=0
cc_357 N_A_398_74#_c_328_n N_A_612_74#_c_679_n 0.00946656f $X=6.5 $Y=2.32 $X2=0
+ $Y2=0
cc_358 N_A_398_74#_c_333_n N_A_612_74#_c_679_n 0.0204128f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_359 N_A_398_74#_c_328_n N_A_612_74#_c_674_n 0.00272661f $X=6.5 $Y=2.32 $X2=0
+ $Y2=0
cc_360 N_A_398_74#_c_334_n N_A_612_74#_c_674_n 0.0283335f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_361 N_A_398_74#_c_350_n N_SET_B_M1016_g 0.00296118f $X=5.52 $Y=2.975 $X2=0
+ $Y2=0
cc_362 N_A_398_74#_c_352_n N_SET_B_M1016_g 0.00987429f $X=5.605 $Y=2.89 $X2=0
+ $Y2=0
cc_363 N_A_398_74#_c_418_p N_SET_B_M1016_g 0.00640039f $X=5.69 $Y=2.405 $X2=0
+ $Y2=0
cc_364 N_A_398_74#_c_382_p N_SET_B_c_804_n 0.0103532f $X=6.415 $Y=2.405 $X2=0
+ $Y2=0
cc_365 N_A_398_74#_c_328_n N_SET_B_c_804_n 0.0176826f $X=6.5 $Y=2.32 $X2=0 $Y2=0
cc_366 N_A_398_74#_c_331_n N_SET_B_c_804_n 0.026653f $X=7.575 $Y=1.98 $X2=0
+ $Y2=0
cc_367 N_A_398_74#_c_333_n N_SET_B_c_804_n 0.00743298f $X=6.795 $Y=1.285 $X2=0
+ $Y2=0
cc_368 N_A_398_74#_c_334_n N_SET_B_c_804_n 0.0015352f $X=6.795 $Y=1.285 $X2=0
+ $Y2=0
cc_369 N_A_398_74#_c_356_n N_SET_B_c_804_n 4.9449e-19 $X=7.455 $Y=2.215 $X2=0
+ $Y2=0
cc_370 N_A_398_74#_c_382_p N_SET_B_c_805_n 0.00857725f $X=6.415 $Y=2.405 $X2=0
+ $Y2=0
cc_371 N_A_398_74#_c_328_n N_SET_B_c_805_n 0.0024765f $X=6.5 $Y=2.32 $X2=0 $Y2=0
cc_372 N_A_398_74#_c_382_p N_SET_B_c_806_n 0.029398f $X=6.415 $Y=2.405 $X2=0
+ $Y2=0
cc_373 N_A_398_74#_c_418_p N_SET_B_c_806_n 0.0118584f $X=5.69 $Y=2.405 $X2=0
+ $Y2=0
cc_374 N_A_398_74#_c_328_n N_SET_B_c_806_n 0.00959664f $X=6.5 $Y=2.32 $X2=0
+ $Y2=0
cc_375 N_A_398_74#_c_331_n SET_B 4.96175e-19 $X=7.575 $Y=1.98 $X2=0 $Y2=0
cc_376 N_A_398_74#_c_331_n N_SET_B_c_798_n 3.31672e-19 $X=7.575 $Y=1.98 $X2=0
+ $Y2=0
cc_377 N_A_398_74#_c_382_p N_SET_B_c_809_n 4.19495e-19 $X=6.415 $Y=2.405 $X2=0
+ $Y2=0
cc_378 N_A_398_74#_c_418_p N_SET_B_c_809_n 6.31522e-19 $X=5.69 $Y=2.405 $X2=0
+ $Y2=0
cc_379 N_A_398_74#_c_322_n N_A_225_74#_M1015_g 0.00164183f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_380 N_A_398_74#_c_324_n N_A_225_74#_M1015_g 0.00266901f $X=2.215 $Y=0.34
+ $X2=0 $Y2=0
cc_381 N_A_398_74#_c_344_n N_A_225_74#_M1017_g 0.00140222f $X=2.275 $Y=2.975
+ $X2=0 $Y2=0
cc_382 N_A_398_74#_c_332_n N_A_225_74#_c_918_n 8.19668e-19 $X=2.95 $Y=1.38 $X2=0
+ $Y2=0
cc_383 N_A_398_74#_c_337_n N_A_225_74#_c_932_n 0.0196818f $X=2.95 $Y=1.885 $X2=0
+ $Y2=0
cc_384 N_A_398_74#_M1023_g N_A_225_74#_c_932_n 0.0192466f $X=3.005 $Y=2.49 $X2=0
+ $Y2=0
cc_385 N_A_398_74#_c_440_p N_A_225_74#_c_932_n 0.00595179f $X=2.19 $Y=2.665
+ $X2=0 $Y2=0
cc_386 N_A_398_74#_c_343_n N_A_225_74#_c_932_n 0.0107799f $X=3.625 $Y=2.975
+ $X2=0 $Y2=0
cc_387 N_A_398_74#_c_325_n N_A_225_74#_c_932_n 3.78496e-19 $X=2.95 $Y=1.545
+ $X2=0 $Y2=0
cc_388 N_A_398_74#_c_318_n N_A_225_74#_c_919_n 0.0147005f $X=2.95 $Y=1.71 $X2=0
+ $Y2=0
cc_389 N_A_398_74#_c_323_n N_A_225_74#_c_919_n 0.00256866f $X=2.945 $Y=0.34
+ $X2=0 $Y2=0
cc_390 N_A_398_74#_c_325_n N_A_225_74#_c_919_n 0.00105733f $X=2.95 $Y=1.545
+ $X2=0 $Y2=0
cc_391 N_A_398_74#_c_332_n N_A_225_74#_c_919_n 0.0074497f $X=2.95 $Y=1.38 $X2=0
+ $Y2=0
cc_392 N_A_398_74#_c_322_n N_A_225_74#_c_920_n 0.00127231f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_393 N_A_398_74#_c_323_n N_A_225_74#_c_920_n 9.7974e-19 $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_394 N_A_398_74#_M1023_g N_A_225_74#_c_933_n 0.00859895f $X=3.005 $Y=2.49
+ $X2=0 $Y2=0
cc_395 N_A_398_74#_c_343_n N_A_225_74#_c_933_n 0.0128486f $X=3.625 $Y=2.975
+ $X2=0 $Y2=0
cc_396 N_A_398_74#_M1012_g N_A_225_74#_M1018_g 0.0087307f $X=3.83 $Y=0.58 $X2=0
+ $Y2=0
cc_397 N_A_398_74#_c_322_n N_A_225_74#_M1018_g 0.00387291f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_398 N_A_398_74#_c_323_n N_A_225_74#_M1018_g 0.0106029f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_399 N_A_398_74#_c_332_n N_A_225_74#_M1018_g 0.021296f $X=2.95 $Y=1.38 $X2=0
+ $Y2=0
cc_400 N_A_398_74#_M1023_g N_A_225_74#_M1021_g 0.0107343f $X=3.005 $Y=2.49 $X2=0
+ $Y2=0
cc_401 N_A_398_74#_c_319_n N_A_225_74#_M1021_g 0.00663151f $X=3.755 $Y=1.545
+ $X2=0 $Y2=0
cc_402 N_A_398_74#_c_343_n N_A_225_74#_M1021_g 0.0184259f $X=3.625 $Y=2.975
+ $X2=0 $Y2=0
cc_403 N_A_398_74#_c_326_n N_A_225_74#_M1021_g 6.57837e-19 $X=3.77 $Y=1.545
+ $X2=0 $Y2=0
cc_404 N_A_398_74#_c_347_n N_A_225_74#_M1021_g 0.00639544f $X=3.71 $Y=2.89 $X2=0
+ $Y2=0
cc_405 N_A_398_74#_c_355_n N_A_225_74#_M1021_g 8.45643e-19 $X=3.77 $Y=2.325
+ $X2=0 $Y2=0
cc_406 N_A_398_74#_c_343_n N_A_225_74#_c_936_n 0.00270445f $X=3.625 $Y=2.975
+ $X2=0 $Y2=0
cc_407 N_A_398_74#_c_348_n N_A_225_74#_c_936_n 0.004087f $X=4.745 $Y=2.325 $X2=0
+ $Y2=0
cc_408 N_A_398_74#_c_350_n N_A_225_74#_c_936_n 0.0125191f $X=5.52 $Y=2.975 $X2=0
+ $Y2=0
cc_409 N_A_398_74#_c_351_n N_A_225_74#_c_936_n 0.00417961f $X=4.915 $Y=2.975
+ $X2=0 $Y2=0
cc_410 N_A_398_74#_c_382_p N_A_225_74#_c_936_n 0.0104482f $X=6.415 $Y=2.405
+ $X2=0 $Y2=0
cc_411 N_A_398_74#_c_355_n N_A_225_74#_c_936_n 2.34075e-19 $X=3.77 $Y=2.325
+ $X2=0 $Y2=0
cc_412 N_A_398_74#_M1010_g N_A_225_74#_M1003_g 0.00633344f $X=7.53 $Y=2.75 $X2=0
+ $Y2=0
cc_413 N_A_398_74#_c_382_p N_A_225_74#_M1003_g 0.0016282f $X=6.415 $Y=2.405
+ $X2=0 $Y2=0
cc_414 N_A_398_74#_c_331_n N_A_225_74#_M1003_g 7.71644e-19 $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_415 N_A_398_74#_c_356_n N_A_225_74#_M1003_g 0.00420587f $X=7.455 $Y=2.215
+ $X2=0 $Y2=0
cc_416 N_A_398_74#_c_331_n N_A_225_74#_c_922_n 0.00260094f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_417 N_A_398_74#_c_356_n N_A_225_74#_c_922_n 0.00860284f $X=7.455 $Y=2.215
+ $X2=0 $Y2=0
cc_418 N_A_398_74#_c_328_n N_A_225_74#_c_923_n 0.00548401f $X=6.5 $Y=2.32 $X2=0
+ $Y2=0
cc_419 N_A_398_74#_c_333_n N_A_225_74#_c_923_n 0.00131539f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_420 N_A_398_74#_c_334_n N_A_225_74#_c_923_n 0.0197635f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_421 N_A_398_74#_c_329_n N_A_225_74#_M1008_g 0.00697755f $X=7.49 $Y=0.365
+ $X2=0 $Y2=0
cc_422 N_A_398_74#_c_331_n N_A_225_74#_M1008_g 0.0129179f $X=7.575 $Y=1.98 $X2=0
+ $Y2=0
cc_423 N_A_398_74#_c_333_n N_A_225_74#_M1008_g 3.37207e-19 $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_424 N_A_398_74#_c_334_n N_A_225_74#_M1008_g 0.0118136f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_425 N_A_398_74#_c_335_n N_A_225_74#_M1008_g 0.0128826f $X=6.795 $Y=1.12 $X2=0
+ $Y2=0
cc_426 N_A_398_74#_c_322_n N_A_225_74#_c_926_n 0.00105443f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_427 N_A_398_74#_c_318_n N_A_225_74#_c_927_n 0.0196818f $X=2.95 $Y=1.71 $X2=0
+ $Y2=0
cc_428 N_A_398_74#_c_325_n N_A_225_74#_c_927_n 3.78496e-19 $X=2.95 $Y=1.545
+ $X2=0 $Y2=0
cc_429 N_A_398_74#_M1017_d N_A_225_74#_c_947_n 0.00277287f $X=2.055 $Y=1.79
+ $X2=0 $Y2=0
cc_430 N_A_398_74#_c_322_n N_A_225_74#_c_929_n 0.0147852f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_431 N_A_398_74#_c_331_n N_A_1566_92#_M1028_g 0.00132255f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_432 N_A_398_74#_c_356_n N_A_1566_92#_M1028_g 0.0511021f $X=7.455 $Y=2.215
+ $X2=0 $Y2=0
cc_433 N_A_398_74#_c_331_n N_A_1566_92#_c_1103_n 0.013857f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_434 N_A_398_74#_c_331_n N_A_1566_92#_c_1112_n 0.0656794f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_435 N_A_398_74#_c_331_n N_A_1566_92#_c_1104_n 0.00795872f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_436 N_A_398_74#_c_331_n N_A_1566_92#_c_1107_n 0.0135436f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_437 N_A_398_74#_c_331_n N_A_1566_92#_c_1115_n 0.00154377f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_438 N_A_398_74#_c_356_n N_A_1566_92#_c_1115_n 0.00529714f $X=7.455 $Y=2.215
+ $X2=0 $Y2=0
cc_439 N_A_398_74#_c_329_n N_A_1356_74#_M1001_d 0.00227017f $X=7.49 $Y=0.365
+ $X2=-0.19 $Y2=-0.245
cc_440 N_A_398_74#_M1010_g N_A_1356_74#_c_1195_n 0.00337976f $X=7.53 $Y=2.75
+ $X2=0 $Y2=0
cc_441 N_A_398_74#_c_382_p N_A_1356_74#_c_1195_n 0.0107347f $X=6.415 $Y=2.405
+ $X2=0 $Y2=0
cc_442 N_A_398_74#_c_328_n N_A_1356_74#_c_1195_n 0.0285493f $X=6.5 $Y=2.32 $X2=0
+ $Y2=0
cc_443 N_A_398_74#_c_331_n N_A_1356_74#_c_1195_n 0.0313601f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_444 N_A_398_74#_c_356_n N_A_1356_74#_c_1195_n 0.00125052f $X=7.455 $Y=2.215
+ $X2=0 $Y2=0
cc_445 N_A_398_74#_c_327_n N_A_1356_74#_c_1186_n 0.00444057f $X=6.5 $Y=1.12
+ $X2=0 $Y2=0
cc_446 N_A_398_74#_c_328_n N_A_1356_74#_c_1186_n 0.00556347f $X=6.5 $Y=2.32
+ $X2=0 $Y2=0
cc_447 N_A_398_74#_c_331_n N_A_1356_74#_c_1186_n 0.0456192f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_448 N_A_398_74#_c_333_n N_A_1356_74#_c_1186_n 0.0236708f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_449 N_A_398_74#_c_334_n N_A_1356_74#_c_1186_n 0.00110295f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_450 N_A_398_74#_c_335_n N_A_1356_74#_c_1186_n 0.00140588f $X=6.795 $Y=1.12
+ $X2=0 $Y2=0
cc_451 N_A_398_74#_M1010_g N_A_1356_74#_c_1216_n 0.0088883f $X=7.53 $Y=2.75
+ $X2=0 $Y2=0
cc_452 N_A_398_74#_c_331_n N_A_1356_74#_c_1216_n 0.00197328f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_453 N_A_398_74#_c_331_n N_A_1356_74#_c_1197_n 0.00449885f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_454 N_A_398_74#_c_356_n N_A_1356_74#_c_1197_n 0.00397026f $X=7.455 $Y=2.215
+ $X2=0 $Y2=0
cc_455 N_A_398_74#_c_328_n N_A_1356_74#_c_1188_n 0.0103198f $X=6.5 $Y=2.32 $X2=0
+ $Y2=0
cc_456 N_A_398_74#_c_331_n N_A_1356_74#_c_1188_n 0.014742f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_457 N_A_398_74#_c_333_n N_A_1356_74#_c_1188_n 0.0101698f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_458 N_A_398_74#_c_334_n N_A_1356_74#_c_1188_n 7.38251e-19 $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_459 N_A_398_74#_M1010_g N_A_1356_74#_c_1202_n 0.00784819f $X=7.53 $Y=2.75
+ $X2=0 $Y2=0
cc_460 N_A_398_74#_c_331_n N_A_1356_74#_c_1202_n 0.020369f $X=7.575 $Y=1.98
+ $X2=0 $Y2=0
cc_461 N_A_398_74#_c_356_n N_A_1356_74#_c_1202_n 9.81303e-19 $X=7.455 $Y=2.215
+ $X2=0 $Y2=0
cc_462 N_A_398_74#_c_329_n N_A_1356_74#_c_1227_n 0.0330935f $X=7.49 $Y=0.365
+ $X2=0 $Y2=0
cc_463 N_A_398_74#_c_333_n N_A_1356_74#_c_1227_n 0.00999825f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_464 N_A_398_74#_c_334_n N_A_1356_74#_c_1227_n 0.00304494f $X=6.795 $Y=1.285
+ $X2=0 $Y2=0
cc_465 N_A_398_74#_c_323_n N_A_27_74#_M1018_s 0.00404388f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_466 N_A_398_74#_M1017_d N_A_27_74#_c_1412_n 0.00574311f $X=2.055 $Y=1.79
+ $X2=0 $Y2=0
cc_467 N_A_398_74#_M1023_g N_A_27_74#_c_1412_n 0.00907948f $X=3.005 $Y=2.49
+ $X2=0 $Y2=0
cc_468 N_A_398_74#_c_342_n N_A_27_74#_c_1412_n 9.41961e-19 $X=2.95 $Y=2.05 $X2=0
+ $Y2=0
cc_469 N_A_398_74#_c_440_p N_A_27_74#_c_1412_n 0.0376834f $X=2.19 $Y=2.665 $X2=0
+ $Y2=0
cc_470 N_A_398_74#_c_343_n N_A_27_74#_c_1412_n 0.0423044f $X=3.625 $Y=2.975
+ $X2=0 $Y2=0
cc_471 N_A_398_74#_c_325_n N_A_27_74#_c_1412_n 0.0115715f $X=2.95 $Y=1.545 $X2=0
+ $Y2=0
cc_472 N_A_398_74#_c_318_n N_A_27_74#_c_1406_n 0.0038721f $X=2.95 $Y=1.71 $X2=0
+ $Y2=0
cc_473 N_A_398_74#_c_322_n N_A_27_74#_c_1406_n 0.0116911f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_474 N_A_398_74#_c_325_n N_A_27_74#_c_1406_n 0.0502423f $X=2.95 $Y=1.545 $X2=0
+ $Y2=0
cc_475 N_A_398_74#_c_332_n N_A_27_74#_c_1406_n 0.0201904f $X=2.95 $Y=1.38 $X2=0
+ $Y2=0
cc_476 N_A_398_74#_c_322_n N_A_27_74#_c_1408_n 0.0206593f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_477 N_A_398_74#_c_323_n N_A_27_74#_c_1408_n 0.0239262f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_478 N_A_398_74#_c_332_n N_A_27_74#_c_1408_n 0.0244211f $X=2.95 $Y=1.38 $X2=0
+ $Y2=0
cc_479 N_A_398_74#_c_348_n N_VPWR_M1032_d 0.0129436f $X=4.745 $Y=2.325 $X2=0
+ $Y2=0
cc_480 N_A_398_74#_c_349_n N_VPWR_M1032_d 0.0101029f $X=4.83 $Y=2.89 $X2=0 $Y2=0
cc_481 N_A_398_74#_c_352_n N_VPWR_M1016_d 0.00292219f $X=5.605 $Y=2.89 $X2=0
+ $Y2=0
cc_482 N_A_398_74#_c_382_p N_VPWR_M1016_d 0.0099895f $X=6.415 $Y=2.405 $X2=0
+ $Y2=0
cc_483 N_A_398_74#_c_418_p N_VPWR_M1016_d 4.66606e-19 $X=5.69 $Y=2.405 $X2=0
+ $Y2=0
cc_484 N_A_398_74#_c_344_n N_VPWR_c_1477_n 0.0118993f $X=2.275 $Y=2.975 $X2=0
+ $Y2=0
cc_485 N_A_398_74#_c_343_n N_VPWR_c_1478_n 0.00905466f $X=3.625 $Y=2.975 $X2=0
+ $Y2=0
cc_486 N_A_398_74#_c_351_n N_VPWR_c_1478_n 0.0059477f $X=4.915 $Y=2.975 $X2=0
+ $Y2=0
cc_487 N_A_398_74#_c_350_n N_VPWR_c_1479_n 0.0146305f $X=5.52 $Y=2.975 $X2=0
+ $Y2=0
cc_488 N_A_398_74#_c_352_n N_VPWR_c_1479_n 0.0174179f $X=5.605 $Y=2.89 $X2=0
+ $Y2=0
cc_489 N_A_398_74#_c_382_p N_VPWR_c_1479_n 0.0189076f $X=6.415 $Y=2.405 $X2=0
+ $Y2=0
cc_490 N_A_398_74#_c_343_n N_VPWR_c_1485_n 0.00124242f $X=3.625 $Y=2.975 $X2=0
+ $Y2=0
cc_491 N_A_398_74#_c_347_n N_VPWR_c_1485_n 0.0110897f $X=3.71 $Y=2.89 $X2=0
+ $Y2=0
cc_492 N_A_398_74#_c_348_n N_VPWR_c_1485_n 0.0384402f $X=4.745 $Y=2.325 $X2=0
+ $Y2=0
cc_493 N_A_398_74#_c_349_n N_VPWR_c_1485_n 0.0250726f $X=4.83 $Y=2.89 $X2=0
+ $Y2=0
cc_494 N_A_398_74#_c_351_n N_VPWR_c_1485_n 0.00174131f $X=4.915 $Y=2.975 $X2=0
+ $Y2=0
cc_495 N_A_398_74#_M1010_g N_VPWR_c_1486_n 0.00380697f $X=7.53 $Y=2.75 $X2=0
+ $Y2=0
cc_496 N_A_398_74#_c_343_n N_VPWR_c_1490_n 0.0896403f $X=3.625 $Y=2.975 $X2=0
+ $Y2=0
cc_497 N_A_398_74#_c_344_n N_VPWR_c_1490_n 0.0111058f $X=2.275 $Y=2.975 $X2=0
+ $Y2=0
cc_498 N_A_398_74#_c_350_n N_VPWR_c_1491_n 0.0466947f $X=5.52 $Y=2.975 $X2=0
+ $Y2=0
cc_499 N_A_398_74#_c_351_n N_VPWR_c_1491_n 0.0111256f $X=4.915 $Y=2.975 $X2=0
+ $Y2=0
cc_500 N_A_398_74#_M1010_g N_VPWR_c_1475_n 0.00478f $X=7.53 $Y=2.75 $X2=0 $Y2=0
cc_501 N_A_398_74#_c_343_n N_VPWR_c_1475_n 0.051041f $X=3.625 $Y=2.975 $X2=0
+ $Y2=0
cc_502 N_A_398_74#_c_344_n N_VPWR_c_1475_n 0.0065564f $X=2.275 $Y=2.975 $X2=0
+ $Y2=0
cc_503 N_A_398_74#_c_350_n N_VPWR_c_1475_n 0.0260024f $X=5.52 $Y=2.975 $X2=0
+ $Y2=0
cc_504 N_A_398_74#_c_351_n N_VPWR_c_1475_n 0.00588338f $X=4.915 $Y=2.975 $X2=0
+ $Y2=0
cc_505 N_A_398_74#_c_382_p N_VPWR_c_1475_n 0.0208508f $X=6.415 $Y=2.405 $X2=0
+ $Y2=0
cc_506 N_A_398_74#_c_347_n A_719_456# 7.96878e-19 $X=3.71 $Y=2.89 $X2=-0.19
+ $Y2=-0.245
cc_507 N_A_398_74#_c_382_p A_1269_341# 0.00412529f $X=6.415 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_508 N_A_398_74#_c_328_n A_1269_341# 0.0159788f $X=6.5 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_509 N_A_398_74#_c_324_n N_VGND_c_1670_n 0.0109685f $X=2.215 $Y=0.34 $X2=0
+ $Y2=0
cc_510 N_A_398_74#_M1012_g N_VGND_c_1671_n 0.00175448f $X=3.83 $Y=0.58 $X2=0
+ $Y2=0
cc_511 N_A_398_74#_c_327_n N_VGND_c_1672_n 0.02453f $X=6.5 $Y=1.12 $X2=0 $Y2=0
cc_512 N_A_398_74#_c_330_n N_VGND_c_1672_n 0.0111625f $X=6.585 $Y=0.365 $X2=0
+ $Y2=0
cc_513 N_A_398_74#_c_335_n N_VGND_c_1672_n 5.00668e-19 $X=6.795 $Y=1.12 $X2=0
+ $Y2=0
cc_514 N_A_398_74#_M1012_g N_VGND_c_1677_n 0.00461464f $X=3.83 $Y=0.58 $X2=0
+ $Y2=0
cc_515 N_A_398_74#_c_323_n N_VGND_c_1677_n 0.0586507f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_516 N_A_398_74#_c_324_n N_VGND_c_1677_n 0.0121867f $X=2.215 $Y=0.34 $X2=0
+ $Y2=0
cc_517 N_A_398_74#_c_329_n N_VGND_c_1679_n 0.0604764f $X=7.49 $Y=0.365 $X2=0
+ $Y2=0
cc_518 N_A_398_74#_c_330_n N_VGND_c_1679_n 0.0105206f $X=6.585 $Y=0.365 $X2=0
+ $Y2=0
cc_519 N_A_398_74#_c_335_n N_VGND_c_1679_n 0.00281891f $X=6.795 $Y=1.12 $X2=0
+ $Y2=0
cc_520 N_A_398_74#_M1012_g N_VGND_c_1687_n 0.00911847f $X=3.83 $Y=0.58 $X2=0
+ $Y2=0
cc_521 N_A_398_74#_c_323_n N_VGND_c_1687_n 0.0333627f $X=2.945 $Y=0.34 $X2=0
+ $Y2=0
cc_522 N_A_398_74#_c_324_n N_VGND_c_1687_n 0.00660921f $X=2.215 $Y=0.34 $X2=0
+ $Y2=0
cc_523 N_A_398_74#_c_329_n N_VGND_c_1687_n 0.0393398f $X=7.49 $Y=0.365 $X2=0
+ $Y2=0
cc_524 N_A_398_74#_c_330_n N_VGND_c_1687_n 0.00652894f $X=6.585 $Y=0.365 $X2=0
+ $Y2=0
cc_525 N_A_398_74#_c_335_n N_VGND_c_1687_n 0.00358754f $X=6.795 $Y=1.12 $X2=0
+ $Y2=0
cc_526 N_A_398_74#_c_327_n A_1278_74# 0.00221695f $X=6.5 $Y=1.12 $X2=-0.19
+ $Y2=-0.245
cc_527 N_A_398_74#_c_331_n A_1489_118# 0.00846132f $X=7.575 $Y=1.98 $X2=-0.19
+ $Y2=-0.245
cc_528 N_A_767_384#_c_590_n N_A_612_74#_M1009_g 0.0217099f $X=5.085 $Y=1.905
+ $X2=0 $Y2=0
cc_529 N_A_767_384#_c_591_n N_A_612_74#_M1009_g 0.0127717f $X=4.395 $Y=1.905
+ $X2=0 $Y2=0
cc_530 N_A_767_384#_c_592_n N_A_612_74#_M1009_g 0.00564729f $X=5.265 $Y=2.52
+ $X2=0 $Y2=0
cc_531 N_A_767_384#_c_593_n N_A_612_74#_M1009_g 0.00979381f $X=5.217 $Y=2.32
+ $X2=0 $Y2=0
cc_532 N_A_767_384#_c_584_n N_A_612_74#_M1002_g 0.0137077f $X=4.575 $Y=1.065
+ $X2=0 $Y2=0
cc_533 N_A_767_384#_c_586_n N_A_612_74#_M1002_g 0.00740402f $X=4.485 $Y=1.065
+ $X2=0 $Y2=0
cc_534 N_A_767_384#_c_584_n N_A_612_74#_c_665_n 0.0144466f $X=4.575 $Y=1.065
+ $X2=0 $Y2=0
cc_535 N_A_767_384#_c_586_n N_A_612_74#_c_665_n 0.00990744f $X=4.485 $Y=1.065
+ $X2=0 $Y2=0
cc_536 N_A_767_384#_c_584_n N_A_612_74#_c_666_n 0.00147785f $X=4.575 $Y=1.065
+ $X2=0 $Y2=0
cc_537 N_A_767_384#_c_586_n N_A_612_74#_c_666_n 0.00411471f $X=4.485 $Y=1.065
+ $X2=0 $Y2=0
cc_538 N_A_767_384#_c_588_n N_A_612_74#_c_667_n 0.00298868f $X=4.23 $Y=1.995
+ $X2=0 $Y2=0
cc_539 N_A_767_384#_c_590_n N_A_612_74#_c_667_n 0.00206546f $X=5.085 $Y=1.905
+ $X2=0 $Y2=0
cc_540 N_A_767_384#_c_591_n N_A_612_74#_c_667_n 2.83197e-19 $X=4.395 $Y=1.905
+ $X2=0 $Y2=0
cc_541 N_A_767_384#_c_590_n N_A_612_74#_c_668_n 0.0146716f $X=5.085 $Y=1.905
+ $X2=0 $Y2=0
cc_542 N_A_767_384#_c_584_n N_A_612_74#_c_668_n 0.0178654f $X=4.575 $Y=1.065
+ $X2=0 $Y2=0
cc_543 N_A_767_384#_c_585_n N_A_612_74#_c_668_n 9.72701e-19 $X=4.395 $Y=1.74
+ $X2=0 $Y2=0
cc_544 N_A_767_384#_c_589_n N_A_612_74#_c_669_n 7.6011e-19 $X=4.015 $Y=1.995
+ $X2=0 $Y2=0
cc_545 N_A_767_384#_c_590_n N_A_612_74#_c_671_n 0.0633465f $X=5.085 $Y=1.905
+ $X2=0 $Y2=0
cc_546 N_A_767_384#_c_591_n N_A_612_74#_c_671_n 0.00165087f $X=4.395 $Y=1.905
+ $X2=0 $Y2=0
cc_547 N_A_767_384#_c_584_n N_A_612_74#_c_671_n 0.0347181f $X=4.575 $Y=1.065
+ $X2=0 $Y2=0
cc_548 N_A_767_384#_c_585_n N_A_612_74#_c_671_n 0.0118646f $X=4.395 $Y=1.74
+ $X2=0 $Y2=0
cc_549 N_A_767_384#_c_586_n N_A_612_74#_c_671_n 0.00436216f $X=4.485 $Y=1.065
+ $X2=0 $Y2=0
cc_550 N_A_767_384#_c_590_n N_A_612_74#_c_673_n 9.26944e-19 $X=5.085 $Y=1.905
+ $X2=0 $Y2=0
cc_551 N_A_767_384#_c_584_n N_A_612_74#_c_673_n 0.00500011f $X=4.575 $Y=1.065
+ $X2=0 $Y2=0
cc_552 N_A_767_384#_c_585_n N_A_612_74#_c_673_n 0.0127717f $X=4.395 $Y=1.74
+ $X2=0 $Y2=0
cc_553 N_A_767_384#_c_586_n N_A_612_74#_c_673_n 6.53703e-19 $X=4.485 $Y=1.065
+ $X2=0 $Y2=0
cc_554 N_A_767_384#_c_590_n N_SET_B_M1022_g 0.00127041f $X=5.085 $Y=1.905 $X2=0
+ $Y2=0
cc_555 N_A_767_384#_c_584_n N_SET_B_M1022_g 0.0013988f $X=4.575 $Y=1.065 $X2=0
+ $Y2=0
cc_556 N_A_767_384#_c_590_n N_SET_B_c_805_n 5.40656e-19 $X=5.085 $Y=1.905 $X2=0
+ $Y2=0
cc_557 N_A_767_384#_c_593_n N_SET_B_c_805_n 2.51551e-19 $X=5.217 $Y=2.32 $X2=0
+ $Y2=0
cc_558 N_A_767_384#_c_590_n N_SET_B_c_806_n 0.0245674f $X=5.085 $Y=1.905 $X2=0
+ $Y2=0
cc_559 N_A_767_384#_c_593_n N_SET_B_c_806_n 0.00609923f $X=5.217 $Y=2.32 $X2=0
+ $Y2=0
cc_560 N_A_767_384#_c_590_n N_SET_B_c_809_n 0.0020735f $X=5.085 $Y=1.905 $X2=0
+ $Y2=0
cc_561 N_A_767_384#_c_593_n N_SET_B_c_809_n 0.0041187f $X=5.217 $Y=2.32 $X2=0
+ $Y2=0
cc_562 N_A_767_384#_M1032_g N_A_225_74#_M1021_g 0.0315834f $X=3.925 $Y=2.49
+ $X2=0 $Y2=0
cc_563 N_A_767_384#_M1032_g N_A_225_74#_c_936_n 0.0102052f $X=3.925 $Y=2.49
+ $X2=0 $Y2=0
cc_564 N_A_767_384#_M1032_g N_VPWR_c_1485_n 0.00568621f $X=3.925 $Y=2.49 $X2=0
+ $Y2=0
cc_565 N_A_767_384#_M1032_g N_VPWR_c_1475_n 0.00114186f $X=3.925 $Y=2.49 $X2=0
+ $Y2=0
cc_566 N_A_767_384#_c_583_n N_VGND_c_1671_n 0.0129647f $X=4.22 $Y=0.9 $X2=0
+ $Y2=0
cc_567 N_A_767_384#_c_584_n N_VGND_c_1671_n 0.0271148f $X=4.575 $Y=1.065 $X2=0
+ $Y2=0
cc_568 N_A_767_384#_c_586_n N_VGND_c_1671_n 0.00527761f $X=4.485 $Y=1.065 $X2=0
+ $Y2=0
cc_569 N_A_767_384#_c_584_n N_VGND_c_1672_n 0.015698f $X=4.575 $Y=1.065 $X2=0
+ $Y2=0
cc_570 N_A_767_384#_c_583_n N_VGND_c_1677_n 0.00383152f $X=4.22 $Y=0.9 $X2=0
+ $Y2=0
cc_571 N_A_767_384#_c_584_n N_VGND_c_1678_n 0.00880728f $X=4.575 $Y=1.065 $X2=0
+ $Y2=0
cc_572 N_A_767_384#_c_583_n N_VGND_c_1687_n 0.0075725f $X=4.22 $Y=0.9 $X2=0
+ $Y2=0
cc_573 N_A_767_384#_c_584_n N_VGND_c_1687_n 0.012195f $X=4.575 $Y=1.065 $X2=0
+ $Y2=0
cc_574 N_A_612_74#_M1011_g N_SET_B_M1016_g 0.0120091f $X=6.255 $Y=2.205 $X2=0
+ $Y2=0
cc_575 N_A_612_74#_M1009_g N_SET_B_M1022_g 0.00824355f $X=5.04 $Y=2.49 $X2=0
+ $Y2=0
cc_576 N_A_612_74#_M1002_g N_SET_B_M1022_g 0.0572199f $X=5.21 $Y=0.8 $X2=0 $Y2=0
cc_577 N_A_612_74#_M1011_g N_SET_B_M1022_g 0.0072922f $X=6.255 $Y=2.205 $X2=0
+ $Y2=0
cc_578 N_A_612_74#_M1000_g N_SET_B_M1022_g 0.00913306f $X=6.315 $Y=0.69 $X2=0
+ $Y2=0
cc_579 N_A_612_74#_c_672_n N_SET_B_M1022_g 0.0211117f $X=5.915 $Y=1.392 $X2=0
+ $Y2=0
cc_580 N_A_612_74#_c_674_n N_SET_B_M1022_g 0.0181307f $X=6.315 $Y=1.38 $X2=0
+ $Y2=0
cc_581 N_A_612_74#_M1011_g N_SET_B_c_804_n 0.00907747f $X=6.255 $Y=2.205 $X2=0
+ $Y2=0
cc_582 N_A_612_74#_c_679_n N_SET_B_c_804_n 0.00333308f $X=6.08 $Y=1.38 $X2=0
+ $Y2=0
cc_583 N_A_612_74#_c_674_n N_SET_B_c_804_n 0.00108234f $X=6.315 $Y=1.38 $X2=0
+ $Y2=0
cc_584 N_A_612_74#_M1011_g N_SET_B_c_805_n 0.00167961f $X=6.255 $Y=2.205 $X2=0
+ $Y2=0
cc_585 N_A_612_74#_c_679_n N_SET_B_c_805_n 0.00126859f $X=6.08 $Y=1.38 $X2=0
+ $Y2=0
cc_586 N_A_612_74#_c_672_n N_SET_B_c_805_n 0.00154953f $X=5.915 $Y=1.392 $X2=0
+ $Y2=0
cc_587 N_A_612_74#_M1009_g N_SET_B_c_806_n 3.5359e-19 $X=5.04 $Y=2.49 $X2=0
+ $Y2=0
cc_588 N_A_612_74#_M1011_g N_SET_B_c_806_n 0.00267248f $X=6.255 $Y=2.205 $X2=0
+ $Y2=0
cc_589 N_A_612_74#_c_672_n N_SET_B_c_806_n 0.044128f $X=5.915 $Y=1.392 $X2=0
+ $Y2=0
cc_590 N_A_612_74#_c_674_n N_SET_B_c_806_n 0.0013286f $X=6.315 $Y=1.38 $X2=0
+ $Y2=0
cc_591 N_A_612_74#_M1009_g N_SET_B_c_809_n 0.0293725f $X=5.04 $Y=2.49 $X2=0
+ $Y2=0
cc_592 N_A_612_74#_M1011_g N_SET_B_c_809_n 0.00866216f $X=6.255 $Y=2.205 $X2=0
+ $Y2=0
cc_593 N_A_612_74#_c_672_n N_SET_B_c_809_n 0.00541653f $X=5.915 $Y=1.392 $X2=0
+ $Y2=0
cc_594 N_A_612_74#_c_670_n N_A_225_74#_c_919_n 4.37445e-19 $X=3.45 $Y=1.125
+ $X2=0 $Y2=0
cc_595 N_A_612_74#_c_664_n N_A_225_74#_M1018_g 0.00255027f $X=3.45 $Y=0.585
+ $X2=0 $Y2=0
cc_596 N_A_612_74#_c_677_n N_A_225_74#_M1021_g 0.00678965f $X=3.28 $Y=2.49 $X2=0
+ $Y2=0
cc_597 N_A_612_74#_c_669_n N_A_225_74#_M1021_g 0.00279843f $X=3.285 $Y=2.26
+ $X2=0 $Y2=0
cc_598 N_A_612_74#_M1009_g N_A_225_74#_c_936_n 0.00859895f $X=5.04 $Y=2.49 $X2=0
+ $Y2=0
cc_599 N_A_612_74#_M1011_g N_A_225_74#_c_936_n 0.0103493f $X=6.255 $Y=2.205
+ $X2=0 $Y2=0
cc_600 N_A_612_74#_M1011_g N_A_225_74#_c_923_n 0.0404199f $X=6.255 $Y=2.205
+ $X2=0 $Y2=0
cc_601 N_A_612_74#_M1011_g N_A_1356_74#_c_1195_n 6.38193e-19 $X=6.255 $Y=2.205
+ $X2=0 $Y2=0
cc_602 N_A_612_74#_M1011_g N_A_1356_74#_c_1202_n 0.00131527f $X=6.255 $Y=2.205
+ $X2=0 $Y2=0
cc_603 N_A_612_74#_c_677_n N_A_27_74#_c_1412_n 0.0200861f $X=3.28 $Y=2.49 $X2=0
+ $Y2=0
cc_604 N_A_612_74#_c_669_n N_A_27_74#_c_1412_n 0.00626792f $X=3.285 $Y=2.26
+ $X2=0 $Y2=0
cc_605 N_A_612_74#_c_669_n N_A_27_74#_c_1406_n 2.70958e-19 $X=3.285 $Y=2.26
+ $X2=0 $Y2=0
cc_606 N_A_612_74#_M1011_g N_VPWR_c_1479_n 0.00424426f $X=6.255 $Y=2.205 $X2=0
+ $Y2=0
cc_607 N_A_612_74#_M1011_g N_VPWR_c_1475_n 0.00113998f $X=6.255 $Y=2.205 $X2=0
+ $Y2=0
cc_608 N_A_612_74#_M1002_g N_VGND_c_1671_n 0.00304548f $X=5.21 $Y=0.8 $X2=0
+ $Y2=0
cc_609 N_A_612_74#_c_664_n N_VGND_c_1671_n 0.00823525f $X=3.45 $Y=0.585 $X2=0
+ $Y2=0
cc_610 N_A_612_74#_M1002_g N_VGND_c_1672_n 0.00183638f $X=5.21 $Y=0.8 $X2=0
+ $Y2=0
cc_611 N_A_612_74#_M1000_g N_VGND_c_1672_n 0.0162104f $X=6.315 $Y=0.69 $X2=0
+ $Y2=0
cc_612 N_A_612_74#_c_679_n N_VGND_c_1672_n 0.0261475f $X=6.08 $Y=1.38 $X2=0
+ $Y2=0
cc_613 N_A_612_74#_c_672_n N_VGND_c_1672_n 0.021427f $X=5.915 $Y=1.392 $X2=0
+ $Y2=0
cc_614 N_A_612_74#_c_674_n N_VGND_c_1672_n 0.00780578f $X=6.315 $Y=1.38 $X2=0
+ $Y2=0
cc_615 N_A_612_74#_c_664_n N_VGND_c_1677_n 0.0118117f $X=3.45 $Y=0.585 $X2=0
+ $Y2=0
cc_616 N_A_612_74#_M1002_g N_VGND_c_1678_n 0.00416964f $X=5.21 $Y=0.8 $X2=0
+ $Y2=0
cc_617 N_A_612_74#_M1000_g N_VGND_c_1679_n 0.00444681f $X=6.315 $Y=0.69 $X2=0
+ $Y2=0
cc_618 N_A_612_74#_M1002_g N_VGND_c_1687_n 0.00479212f $X=5.21 $Y=0.8 $X2=0
+ $Y2=0
cc_619 N_A_612_74#_M1000_g N_VGND_c_1687_n 0.00877228f $X=6.315 $Y=0.69 $X2=0
+ $Y2=0
cc_620 N_A_612_74#_c_664_n N_VGND_c_1687_n 0.011742f $X=3.45 $Y=0.585 $X2=0
+ $Y2=0
cc_621 N_SET_B_M1016_g N_A_225_74#_c_936_n 0.00861849f $X=5.49 $Y=2.49 $X2=0
+ $Y2=0
cc_622 N_SET_B_c_804_n N_A_225_74#_M1003_g 0.00924927f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_623 N_SET_B_c_804_n N_A_225_74#_c_922_n 0.00682877f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_624 N_SET_B_c_803_n N_A_1566_92#_M1028_g 0.0255676f $X=8.565 $Y=2.15 $X2=0
+ $Y2=0
cc_625 SET_B N_A_1566_92#_M1028_g 3.05387e-19 $X=8.315 $Y=1.95 $X2=0 $Y2=0
cc_626 N_SET_B_M1004_g N_A_1566_92#_c_1103_n 0.0205048f $X=8.475 $Y=0.8 $X2=0
+ $Y2=0
cc_627 N_SET_B_M1004_g N_A_1566_92#_c_1112_n 0.00149238f $X=8.475 $Y=0.8 $X2=0
+ $Y2=0
cc_628 N_SET_B_c_804_n N_A_1566_92#_c_1112_n 0.027726f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_629 SET_B N_A_1566_92#_c_1112_n 0.00213174f $X=8.315 $Y=1.95 $X2=0 $Y2=0
cc_630 N_SET_B_c_797_n N_A_1566_92#_c_1112_n 7.54692e-19 $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_631 N_SET_B_c_798_n N_A_1566_92#_c_1112_n 0.0495655f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_632 N_SET_B_M1004_g N_A_1566_92#_c_1104_n 0.0182739f $X=8.475 $Y=0.8 $X2=0
+ $Y2=0
cc_633 SET_B N_A_1566_92#_c_1105_n 7.33174e-19 $X=8.315 $Y=1.95 $X2=0 $Y2=0
cc_634 N_SET_B_c_797_n N_A_1566_92#_c_1105_n 0.0182739f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_635 N_SET_B_c_798_n N_A_1566_92#_c_1105_n 0.0038385f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_636 N_SET_B_M1004_g N_A_1566_92#_c_1106_n 0.0165527f $X=8.475 $Y=0.8 $X2=0
+ $Y2=0
cc_637 N_SET_B_c_797_n N_A_1566_92#_c_1106_n 0.00116081f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_638 N_SET_B_c_798_n N_A_1566_92#_c_1106_n 0.0252292f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_639 N_SET_B_c_796_n N_A_1566_92#_c_1115_n 0.0182739f $X=8.565 $Y=1.985 $X2=0
+ $Y2=0
cc_640 N_SET_B_c_804_n N_A_1566_92#_c_1115_n 0.00323607f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_641 SET_B N_A_1566_92#_c_1115_n 4.08782e-19 $X=8.315 $Y=1.95 $X2=0 $Y2=0
cc_642 N_SET_B_c_804_n N_A_1356_74#_M1003_d 0.00115767f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_643 N_SET_B_c_797_n N_A_1356_74#_M1027_g 0.00259971f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_644 N_SET_B_c_798_n N_A_1356_74#_M1027_g 6.32828e-19 $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_645 N_SET_B_c_797_n N_A_1356_74#_c_1184_n 0.00494777f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_646 N_SET_B_c_798_n N_A_1356_74#_c_1184_n 0.0024583f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_647 N_SET_B_M1007_g N_A_1356_74#_c_1193_n 0.00328286f $X=8.49 $Y=2.75 $X2=0
+ $Y2=0
cc_648 N_SET_B_c_803_n N_A_1356_74#_c_1193_n 0.00494777f $X=8.565 $Y=2.15 $X2=0
+ $Y2=0
cc_649 N_SET_B_c_804_n N_A_1356_74#_c_1195_n 0.0144054f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_650 N_SET_B_c_804_n N_A_1356_74#_c_1216_n 0.00350245f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_651 N_SET_B_M1007_g N_A_1356_74#_c_1196_n 0.0185963f $X=8.49 $Y=2.75 $X2=0
+ $Y2=0
cc_652 N_SET_B_c_803_n N_A_1356_74#_c_1196_n 3.53728e-19 $X=8.565 $Y=2.15 $X2=0
+ $Y2=0
cc_653 N_SET_B_c_804_n N_A_1356_74#_c_1196_n 0.00640638f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_654 SET_B N_A_1356_74#_c_1196_n 0.00471918f $X=8.315 $Y=1.95 $X2=0 $Y2=0
cc_655 N_SET_B_c_798_n N_A_1356_74#_c_1196_n 0.0215664f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_656 N_SET_B_M1007_g N_A_1356_74#_c_1197_n 6.94529e-19 $X=8.49 $Y=2.75 $X2=0
+ $Y2=0
cc_657 N_SET_B_c_804_n N_A_1356_74#_c_1197_n 0.00403539f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_658 N_SET_B_M1007_g N_A_1356_74#_c_1198_n 8.70751e-19 $X=8.49 $Y=2.75 $X2=0
+ $Y2=0
cc_659 N_SET_B_M1007_g N_A_1356_74#_c_1187_n 0.00157501f $X=8.49 $Y=2.75 $X2=0
+ $Y2=0
cc_660 SET_B N_A_1356_74#_c_1187_n 0.00107107f $X=8.315 $Y=1.95 $X2=0 $Y2=0
cc_661 N_SET_B_c_797_n N_A_1356_74#_c_1187_n 0.00225352f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_662 N_SET_B_c_798_n N_A_1356_74#_c_1187_n 0.018807f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_663 N_SET_B_c_796_n N_A_1356_74#_c_1201_n 0.00494777f $X=8.565 $Y=1.985 $X2=0
+ $Y2=0
cc_664 N_SET_B_c_804_n N_A_1356_74#_c_1188_n 0.0111047f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_665 N_SET_B_c_804_n N_A_1356_74#_c_1202_n 0.0108184f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_666 N_SET_B_c_803_n N_A_1356_74#_c_1203_n 7.69224e-19 $X=8.565 $Y=2.15 $X2=0
+ $Y2=0
cc_667 N_SET_B_c_798_n N_A_1356_74#_c_1203_n 0.00879631f $X=8.565 $Y=1.645 $X2=0
+ $Y2=0
cc_668 N_SET_B_c_804_n N_VPWR_M1016_d 3.55183e-19 $X=8.255 $Y=2.035 $X2=0 $Y2=0
cc_669 N_SET_B_c_805_n N_VPWR_M1016_d 0.00299204f $X=6.145 $Y=2.035 $X2=0 $Y2=0
cc_670 N_SET_B_c_806_n N_VPWR_M1016_d 0.00617186f $X=6 $Y=2.035 $X2=0 $Y2=0
cc_671 N_SET_B_M1016_g N_VPWR_c_1479_n 5.38053e-19 $X=5.49 $Y=2.49 $X2=0 $Y2=0
cc_672 N_SET_B_M1007_g N_VPWR_c_1480_n 0.0105772f $X=8.49 $Y=2.75 $X2=0 $Y2=0
cc_673 N_SET_B_M1007_g N_VPWR_c_1481_n 0.00336103f $X=8.49 $Y=2.75 $X2=0 $Y2=0
cc_674 N_SET_B_M1007_g N_VPWR_c_1492_n 0.00460063f $X=8.49 $Y=2.75 $X2=0 $Y2=0
cc_675 N_SET_B_M1007_g N_VPWR_c_1475_n 0.004509f $X=8.49 $Y=2.75 $X2=0 $Y2=0
cc_676 N_SET_B_c_804_n A_1269_341# 0.00663364f $X=8.255 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_677 N_SET_B_M1022_g N_VGND_c_1672_n 0.0149224f $X=5.6 $Y=0.8 $X2=0 $Y2=0
cc_678 N_SET_B_M1022_g N_VGND_c_1678_n 0.00360926f $X=5.6 $Y=0.8 $X2=0 $Y2=0
cc_679 N_SET_B_M1004_g N_VGND_c_1679_n 0.0172888f $X=8.475 $Y=0.8 $X2=0 $Y2=0
cc_680 N_SET_B_M1022_g N_VGND_c_1687_n 0.00402538f $X=5.6 $Y=0.8 $X2=0 $Y2=0
cc_681 N_SET_B_M1004_g N_VGND_c_1687_n 0.00402538f $X=8.475 $Y=0.8 $X2=0 $Y2=0
cc_682 N_A_225_74#_M1008_g N_A_1566_92#_c_1103_n 0.0158751f $X=7.37 $Y=0.8 $X2=0
+ $Y2=0
cc_683 N_A_225_74#_c_922_n N_A_1566_92#_c_1104_n 0.0158751f $X=7.295 $Y=1.735
+ $X2=0 $Y2=0
cc_684 N_A_225_74#_M1003_g N_A_1356_74#_c_1195_n 0.0125297f $X=6.76 $Y=2.46
+ $X2=0 $Y2=0
cc_685 N_A_225_74#_c_922_n N_A_1356_74#_c_1195_n 0.00672058f $X=7.295 $Y=1.735
+ $X2=0 $Y2=0
cc_686 N_A_225_74#_c_923_n N_A_1356_74#_c_1195_n 3.44404e-19 $X=6.85 $Y=1.735
+ $X2=0 $Y2=0
cc_687 N_A_225_74#_c_922_n N_A_1356_74#_c_1186_n 0.0015047f $X=7.295 $Y=1.735
+ $X2=0 $Y2=0
cc_688 N_A_225_74#_M1008_g N_A_1356_74#_c_1186_n 0.0149235f $X=7.37 $Y=0.8 $X2=0
+ $Y2=0
cc_689 N_A_225_74#_c_922_n N_A_1356_74#_c_1188_n 0.0155989f $X=7.295 $Y=1.735
+ $X2=0 $Y2=0
cc_690 N_A_225_74#_c_923_n N_A_1356_74#_c_1188_n 0.00183273f $X=6.85 $Y=1.735
+ $X2=0 $Y2=0
cc_691 N_A_225_74#_M1008_g N_A_1356_74#_c_1188_n 0.00131824f $X=7.37 $Y=0.8
+ $X2=0 $Y2=0
cc_692 N_A_225_74#_M1003_g N_A_1356_74#_c_1202_n 0.0179354f $X=6.76 $Y=2.46
+ $X2=0 $Y2=0
cc_693 N_A_225_74#_M1008_g N_A_1356_74#_c_1227_n 0.00926501f $X=7.37 $Y=0.8
+ $X2=0 $Y2=0
cc_694 N_A_225_74#_M1014_s N_A_27_74#_c_1411_n 0.0117593f $X=1.145 $Y=1.79 $X2=0
+ $Y2=0
cc_695 N_A_225_74#_c_945_n N_A_27_74#_c_1411_n 0.0189258f $X=1.305 $Y=1.87 $X2=0
+ $Y2=0
cc_696 N_A_225_74#_c_946_n N_A_27_74#_c_1411_n 0.0142272f $X=1.145 $Y=1.87 $X2=0
+ $Y2=0
cc_697 N_A_225_74#_c_947_n N_A_27_74#_c_1411_n 0.00643406f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_698 N_A_225_74#_M1017_g N_A_27_74#_c_1412_n 0.0165851f $X=1.965 $Y=2.35 $X2=0
+ $Y2=0
cc_699 N_A_225_74#_c_932_n N_A_27_74#_c_1412_n 0.0262382f $X=2.485 $Y=3.075
+ $X2=0 $Y2=0
cc_700 N_A_225_74#_c_926_n N_A_27_74#_c_1412_n 0.00180813f $X=2.41 $Y=1.465
+ $X2=0 $Y2=0
cc_701 N_A_225_74#_c_947_n N_A_27_74#_c_1412_n 0.0277303f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_702 N_A_225_74#_M1015_g N_A_27_74#_c_1406_n 7.54241e-19 $X=1.915 $Y=0.74
+ $X2=0 $Y2=0
cc_703 N_A_225_74#_M1017_g N_A_27_74#_c_1406_n 0.00119828f $X=1.965 $Y=2.35
+ $X2=0 $Y2=0
cc_704 N_A_225_74#_c_918_n N_A_27_74#_c_1406_n 0.00518646f $X=2.485 $Y=1.3 $X2=0
+ $Y2=0
cc_705 N_A_225_74#_c_932_n N_A_27_74#_c_1406_n 0.00987763f $X=2.485 $Y=3.075
+ $X2=0 $Y2=0
cc_706 N_A_225_74#_c_919_n N_A_27_74#_c_1406_n 0.00578804f $X=2.91 $Y=1.065
+ $X2=0 $Y2=0
cc_707 N_A_225_74#_c_920_n N_A_27_74#_c_1406_n 0.00450019f $X=2.56 $Y=1.065
+ $X2=0 $Y2=0
cc_708 N_A_225_74#_M1018_g N_A_27_74#_c_1406_n 0.00115087f $X=2.985 $Y=0.58
+ $X2=0 $Y2=0
cc_709 N_A_225_74#_c_927_n N_A_27_74#_c_1406_n 0.0101071f $X=2.485 $Y=1.465
+ $X2=0 $Y2=0
cc_710 N_A_225_74#_c_947_n N_A_27_74#_c_1406_n 0.0135406f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_711 N_A_225_74#_c_929_n N_A_27_74#_c_1406_n 0.0302859f $X=2.11 $Y=1.465 $X2=0
+ $Y2=0
cc_712 N_A_225_74#_M1017_g N_A_27_74#_c_1459_n 0.00187706f $X=1.965 $Y=2.35
+ $X2=0 $Y2=0
cc_713 N_A_225_74#_c_947_n N_A_27_74#_c_1459_n 0.0100622f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_714 N_A_225_74#_c_919_n N_A_27_74#_c_1408_n 0.00669646f $X=2.91 $Y=1.065
+ $X2=0 $Y2=0
cc_715 N_A_225_74#_c_920_n N_A_27_74#_c_1408_n 0.00134438f $X=2.56 $Y=1.065
+ $X2=0 $Y2=0
cc_716 N_A_225_74#_M1018_g N_A_27_74#_c_1408_n 0.0066603f $X=2.985 $Y=0.58 $X2=0
+ $Y2=0
cc_717 N_A_225_74#_c_947_n N_VPWR_M1014_d 0.00164828f $X=1.945 $Y=1.805 $X2=0
+ $Y2=0
cc_718 N_A_225_74#_M1017_g N_VPWR_c_1477_n 0.00884425f $X=1.965 $Y=2.35 $X2=0
+ $Y2=0
cc_719 N_A_225_74#_c_932_n N_VPWR_c_1477_n 0.00346637f $X=2.485 $Y=3.075 $X2=0
+ $Y2=0
cc_720 N_A_225_74#_M1021_g N_VPWR_c_1478_n 0.00103154f $X=3.505 $Y=2.49 $X2=0
+ $Y2=0
cc_721 N_A_225_74#_c_936_n N_VPWR_c_1478_n 0.0160168f $X=6.67 $Y=3.15 $X2=0
+ $Y2=0
cc_722 N_A_225_74#_c_936_n N_VPWR_c_1479_n 0.021028f $X=6.67 $Y=3.15 $X2=0 $Y2=0
cc_723 N_A_225_74#_M1003_g N_VPWR_c_1479_n 0.00617957f $X=6.76 $Y=2.46 $X2=0
+ $Y2=0
cc_724 N_A_225_74#_M1021_g N_VPWR_c_1485_n 2.53362e-19 $X=3.505 $Y=2.49 $X2=0
+ $Y2=0
cc_725 N_A_225_74#_c_936_n N_VPWR_c_1485_n 0.00817058f $X=6.67 $Y=3.15 $X2=0
+ $Y2=0
cc_726 N_A_225_74#_c_936_n N_VPWR_c_1486_n 0.0266714f $X=6.67 $Y=3.15 $X2=0
+ $Y2=0
cc_727 N_A_225_74#_M1017_g N_VPWR_c_1490_n 0.00540231f $X=1.965 $Y=2.35 $X2=0
+ $Y2=0
cc_728 N_A_225_74#_c_934_n N_VPWR_c_1490_n 0.0400301f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_729 N_A_225_74#_c_936_n N_VPWR_c_1491_n 0.0386563f $X=6.67 $Y=3.15 $X2=0
+ $Y2=0
cc_730 N_A_225_74#_M1017_g N_VPWR_c_1475_n 0.00533457f $X=1.965 $Y=2.35 $X2=0
+ $Y2=0
cc_731 N_A_225_74#_c_933_n N_VPWR_c_1475_n 0.0201442f $X=3.415 $Y=3.15 $X2=0
+ $Y2=0
cc_732 N_A_225_74#_c_934_n N_VPWR_c_1475_n 0.00604809f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_733 N_A_225_74#_c_936_n N_VPWR_c_1475_n 0.0908446f $X=6.67 $Y=3.15 $X2=0
+ $Y2=0
cc_734 N_A_225_74#_c_943_n N_VPWR_c_1475_n 0.00445365f $X=3.505 $Y=3.15 $X2=0
+ $Y2=0
cc_735 N_A_225_74#_c_930_n N_VGND_c_1668_n 0.0327823f $X=1.27 $Y=0.51 $X2=0
+ $Y2=0
cc_736 N_A_225_74#_c_930_n N_VGND_c_1669_n 0.0203368f $X=1.27 $Y=0.51 $X2=0
+ $Y2=0
cc_737 N_A_225_74#_M1015_g N_VGND_c_1670_n 0.0115598f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_738 N_A_225_74#_c_930_n N_VGND_c_1670_n 0.0256161f $X=1.27 $Y=0.51 $X2=0
+ $Y2=0
cc_739 N_A_225_74#_M1015_g N_VGND_c_1677_n 0.00383152f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_740 N_A_225_74#_M1018_g N_VGND_c_1677_n 0.00278159f $X=2.985 $Y=0.58 $X2=0
+ $Y2=0
cc_741 N_A_225_74#_M1015_g N_VGND_c_1687_n 0.00762539f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_742 N_A_225_74#_M1018_g N_VGND_c_1687_n 0.00361237f $X=2.985 $Y=0.58 $X2=0
+ $Y2=0
cc_743 N_A_225_74#_c_930_n N_VGND_c_1687_n 0.0167889f $X=1.27 $Y=0.51 $X2=0
+ $Y2=0
cc_744 N_A_1566_92#_c_1106_n N_A_1356_74#_M1027_g 0.0152849f $X=9.53 $Y=1.155
+ $X2=0 $Y2=0
cc_745 N_A_1566_92#_c_1108_n N_A_1356_74#_M1027_g 0.0121665f $X=9.695 $Y=0.8
+ $X2=0 $Y2=0
cc_746 N_A_1566_92#_c_1109_n N_A_1356_74#_M1027_g 0.0147061f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_747 N_A_1566_92#_c_1110_n N_A_1356_74#_M1027_g 0.00513932f $X=9.71 $Y=1.155
+ $X2=0 $Y2=0
cc_748 N_A_1566_92#_c_1109_n N_A_1356_74#_c_1182_n 0.0188128f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_749 N_A_1566_92#_c_1109_n N_A_1356_74#_M1013_g 0.0014319f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_750 N_A_1566_92#_c_1110_n N_A_1356_74#_M1013_g 6.25308e-19 $X=9.71 $Y=1.155
+ $X2=0 $Y2=0
cc_751 N_A_1566_92#_c_1109_n N_A_1356_74#_c_1191_n 0.00454641f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_752 N_A_1566_92#_c_1106_n N_A_1356_74#_c_1184_n 0.00155183f $X=9.53 $Y=1.155
+ $X2=0 $Y2=0
cc_753 N_A_1566_92#_M1028_g N_A_1356_74#_c_1216_n 2.21133e-19 $X=7.95 $Y=2.75
+ $X2=0 $Y2=0
cc_754 N_A_1566_92#_M1028_g N_A_1356_74#_c_1196_n 0.0103155f $X=7.95 $Y=2.75
+ $X2=0 $Y2=0
cc_755 N_A_1566_92#_c_1112_n N_A_1356_74#_c_1196_n 0.0141202f $X=7.995 $Y=1.285
+ $X2=0 $Y2=0
cc_756 N_A_1566_92#_c_1115_n N_A_1356_74#_c_1196_n 0.00139354f $X=7.995 $Y=2.13
+ $X2=0 $Y2=0
cc_757 N_A_1566_92#_M1028_g N_A_1356_74#_c_1197_n 0.0106077f $X=7.95 $Y=2.75
+ $X2=0 $Y2=0
cc_758 N_A_1566_92#_c_1112_n N_A_1356_74#_c_1197_n 0.00668502f $X=7.995 $Y=1.285
+ $X2=0 $Y2=0
cc_759 N_A_1566_92#_c_1115_n N_A_1356_74#_c_1197_n 2.12417e-19 $X=7.995 $Y=2.13
+ $X2=0 $Y2=0
cc_760 N_A_1566_92#_c_1109_n N_A_1356_74#_c_1199_n 0.0139713f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_761 N_A_1566_92#_c_1106_n N_A_1356_74#_c_1187_n 0.0142071f $X=9.53 $Y=1.155
+ $X2=0 $Y2=0
cc_762 N_A_1566_92#_c_1109_n N_A_1356_74#_c_1187_n 0.0538376f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_763 N_A_1566_92#_c_1109_n N_A_1356_74#_c_1201_n 0.0222711f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_764 N_A_1566_92#_M1028_g N_A_1356_74#_c_1202_n 7.30961e-19 $X=7.95 $Y=2.75
+ $X2=0 $Y2=0
cc_765 N_A_1566_92#_c_1108_n N_A_2022_94#_c_1339_n 0.0324928f $X=9.695 $Y=0.8
+ $X2=0 $Y2=0
cc_766 N_A_1566_92#_c_1109_n N_A_2022_94#_c_1339_n 0.00429293f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_767 N_A_1566_92#_c_1110_n N_A_2022_94#_c_1339_n 0.0134078f $X=9.71 $Y=1.155
+ $X2=0 $Y2=0
cc_768 N_A_1566_92#_c_1109_n N_A_2022_94#_c_1345_n 0.0889488f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_769 N_A_1566_92#_c_1109_n N_A_2022_94#_c_1341_n 0.0253904f $X=9.725 $Y=2.75
+ $X2=0 $Y2=0
cc_770 N_A_1566_92#_M1028_g N_VPWR_c_1480_n 0.00694744f $X=7.95 $Y=2.75 $X2=0
+ $Y2=0
cc_771 N_A_1566_92#_c_1109_n N_VPWR_c_1481_n 0.0112185f $X=9.725 $Y=2.75 $X2=0
+ $Y2=0
cc_772 N_A_1566_92#_M1028_g N_VPWR_c_1486_n 0.00489722f $X=7.95 $Y=2.75 $X2=0
+ $Y2=0
cc_773 N_A_1566_92#_c_1109_n N_VPWR_c_1493_n 0.011066f $X=9.725 $Y=2.75 $X2=0
+ $Y2=0
cc_774 N_A_1566_92#_M1028_g N_VPWR_c_1475_n 0.00515927f $X=7.95 $Y=2.75 $X2=0
+ $Y2=0
cc_775 N_A_1566_92#_c_1109_n N_VPWR_c_1475_n 0.00915947f $X=9.725 $Y=2.75 $X2=0
+ $Y2=0
cc_776 N_A_1566_92#_c_1103_n N_VGND_c_1679_n 0.00633226f $X=7.995 $Y=1.12 $X2=0
+ $Y2=0
cc_777 N_A_1566_92#_c_1106_n N_VGND_c_1679_n 0.0656301f $X=9.53 $Y=1.155 $X2=0
+ $Y2=0
cc_778 N_A_1566_92#_c_1108_n N_VGND_c_1680_n 0.00636076f $X=9.695 $Y=0.8 $X2=0
+ $Y2=0
cc_779 N_A_1566_92#_c_1103_n N_VGND_c_1687_n 0.00479212f $X=7.995 $Y=1.12 $X2=0
+ $Y2=0
cc_780 N_A_1566_92#_c_1108_n N_VGND_c_1687_n 0.010804f $X=9.695 $Y=0.8 $X2=0
+ $Y2=0
cc_781 N_A_1356_74#_c_1185_n N_A_2022_94#_M1026_g 0.0291277f $X=10.497 $Y=1.69
+ $X2=0 $Y2=0
cc_782 N_A_1356_74#_M1013_g N_A_2022_94#_M1005_g 0.0194305f $X=10.47 $Y=0.79
+ $X2=0 $Y2=0
cc_783 N_A_1356_74#_M1027_g N_A_2022_94#_c_1339_n 0.00555362f $X=9.48 $Y=0.8
+ $X2=0 $Y2=0
cc_784 N_A_1356_74#_M1013_g N_A_2022_94#_c_1339_n 0.0151436f $X=10.47 $Y=0.79
+ $X2=0 $Y2=0
cc_785 N_A_1356_74#_c_1182_n N_A_2022_94#_c_1345_n 0.0116701f $X=10.395 $Y=1.69
+ $X2=0 $Y2=0
cc_786 N_A_1356_74#_c_1191_n N_A_2022_94#_c_1345_n 0.0176844f $X=10.51 $Y=1.765
+ $X2=0 $Y2=0
cc_787 N_A_1356_74#_c_1185_n N_A_2022_94#_c_1345_n 0.00308043f $X=10.497 $Y=1.69
+ $X2=0 $Y2=0
cc_788 N_A_1356_74#_M1013_g N_A_2022_94#_c_1340_n 0.0107422f $X=10.47 $Y=0.79
+ $X2=0 $Y2=0
cc_789 N_A_1356_74#_c_1185_n N_A_2022_94#_c_1340_n 0.00855895f $X=10.497 $Y=1.69
+ $X2=0 $Y2=0
cc_790 N_A_1356_74#_c_1182_n N_A_2022_94#_c_1341_n 0.00584559f $X=10.395 $Y=1.69
+ $X2=0 $Y2=0
cc_791 N_A_1356_74#_M1013_g N_A_2022_94#_c_1341_n 0.00952755f $X=10.47 $Y=0.79
+ $X2=0 $Y2=0
cc_792 N_A_1356_74#_M1013_g N_A_2022_94#_c_1342_n 0.0153086f $X=10.47 $Y=0.79
+ $X2=0 $Y2=0
cc_793 N_A_1356_74#_c_1185_n N_A_2022_94#_c_1342_n 9.99338e-19 $X=10.497 $Y=1.69
+ $X2=0 $Y2=0
cc_794 N_A_1356_74#_c_1196_n N_VPWR_M1028_d 0.00254801f $X=8.63 $Y=2.435 $X2=0
+ $Y2=0
cc_795 N_A_1356_74#_c_1196_n N_VPWR_c_1480_n 0.0211289f $X=8.63 $Y=2.435 $X2=0
+ $Y2=0
cc_796 N_A_1356_74#_c_1197_n N_VPWR_c_1480_n 7.39923e-19 $X=7.93 $Y=2.435 $X2=0
+ $Y2=0
cc_797 N_A_1356_74#_c_1198_n N_VPWR_c_1480_n 0.00924182f $X=8.715 $Y=2.75 $X2=0
+ $Y2=0
cc_798 N_A_1356_74#_c_1202_n N_VPWR_c_1480_n 0.00722809f $X=7.47 $Y=2.765 $X2=0
+ $Y2=0
cc_799 N_A_1356_74#_M1019_g N_VPWR_c_1481_n 0.0123584f $X=9.5 $Y=2.75 $X2=0
+ $Y2=0
cc_800 N_A_1356_74#_c_1193_n N_VPWR_c_1481_n 0.00119861f $X=9.365 $Y=2.285 $X2=0
+ $Y2=0
cc_801 N_A_1356_74#_c_1198_n N_VPWR_c_1481_n 0.0211298f $X=8.715 $Y=2.75 $X2=0
+ $Y2=0
cc_802 N_A_1356_74#_c_1199_n N_VPWR_c_1481_n 0.0263373f $X=9.14 $Y=2.405 $X2=0
+ $Y2=0
cc_803 N_A_1356_74#_c_1191_n N_VPWR_c_1482_n 0.00609461f $X=10.51 $Y=1.765 $X2=0
+ $Y2=0
cc_804 N_A_1356_74#_c_1216_n N_VPWR_c_1486_n 0.00485016f $X=7.76 $Y=2.64 $X2=0
+ $Y2=0
cc_805 N_A_1356_74#_c_1197_n N_VPWR_c_1486_n 0.0027555f $X=7.93 $Y=2.435 $X2=0
+ $Y2=0
cc_806 N_A_1356_74#_c_1202_n N_VPWR_c_1486_n 0.0277579f $X=7.47 $Y=2.765 $X2=0
+ $Y2=0
cc_807 N_A_1356_74#_c_1198_n N_VPWR_c_1492_n 0.0110419f $X=8.715 $Y=2.75 $X2=0
+ $Y2=0
cc_808 N_A_1356_74#_M1019_g N_VPWR_c_1493_n 0.00460063f $X=9.5 $Y=2.75 $X2=0
+ $Y2=0
cc_809 N_A_1356_74#_c_1191_n N_VPWR_c_1493_n 0.00567889f $X=10.51 $Y=1.765 $X2=0
+ $Y2=0
cc_810 N_A_1356_74#_M1019_g N_VPWR_c_1475_n 0.00821725f $X=9.5 $Y=2.75 $X2=0
+ $Y2=0
cc_811 N_A_1356_74#_c_1191_n N_VPWR_c_1475_n 0.00610055f $X=10.51 $Y=1.765 $X2=0
+ $Y2=0
cc_812 N_A_1356_74#_c_1216_n N_VPWR_c_1475_n 0.00777687f $X=7.76 $Y=2.64 $X2=0
+ $Y2=0
cc_813 N_A_1356_74#_c_1196_n N_VPWR_c_1475_n 0.0131548f $X=8.63 $Y=2.435 $X2=0
+ $Y2=0
cc_814 N_A_1356_74#_c_1197_n N_VPWR_c_1475_n 0.0047639f $X=7.93 $Y=2.435 $X2=0
+ $Y2=0
cc_815 N_A_1356_74#_c_1198_n N_VPWR_c_1475_n 0.00915013f $X=8.715 $Y=2.75 $X2=0
+ $Y2=0
cc_816 N_A_1356_74#_c_1199_n N_VPWR_c_1475_n 0.0101037f $X=9.14 $Y=2.405 $X2=0
+ $Y2=0
cc_817 N_A_1356_74#_c_1202_n N_VPWR_c_1475_n 0.0233342f $X=7.47 $Y=2.765 $X2=0
+ $Y2=0
cc_818 N_A_1356_74#_c_1216_n A_1524_508# 0.00327035f $X=7.76 $Y=2.64 $X2=-0.19
+ $Y2=-0.245
cc_819 N_A_1356_74#_c_1197_n A_1524_508# 0.00127389f $X=7.93 $Y=2.435 $X2=-0.19
+ $Y2=-0.245
cc_820 N_A_1356_74#_c_1191_n N_Q_c_1635_n 0.00326353f $X=10.51 $Y=1.765 $X2=0
+ $Y2=0
cc_821 N_A_1356_74#_M1013_g N_VGND_c_1673_n 0.00744268f $X=10.47 $Y=0.79 $X2=0
+ $Y2=0
cc_822 N_A_1356_74#_M1027_g N_VGND_c_1679_n 0.0120948f $X=9.48 $Y=0.8 $X2=0
+ $Y2=0
cc_823 N_A_1356_74#_M1027_g N_VGND_c_1680_n 0.00418347f $X=9.48 $Y=0.8 $X2=0
+ $Y2=0
cc_824 N_A_1356_74#_M1013_g N_VGND_c_1680_n 0.00485498f $X=10.47 $Y=0.79 $X2=0
+ $Y2=0
cc_825 N_A_1356_74#_M1027_g N_VGND_c_1687_n 0.00479212f $X=9.48 $Y=0.8 $X2=0
+ $Y2=0
cc_826 N_A_1356_74#_M1013_g N_VGND_c_1687_n 0.00514438f $X=10.47 $Y=0.79 $X2=0
+ $Y2=0
cc_827 N_A_2022_94#_M1026_g N_VPWR_c_1482_n 0.0133705f $X=11.045 $Y=2.4 $X2=0
+ $Y2=0
cc_828 N_A_2022_94#_M1029_g N_VPWR_c_1482_n 5.31852e-19 $X=11.495 $Y=2.4 $X2=0
+ $Y2=0
cc_829 N_A_2022_94#_c_1345_n N_VPWR_c_1482_n 0.0183701f $X=10.285 $Y=1.985 $X2=0
+ $Y2=0
cc_830 N_A_2022_94#_M1029_g N_VPWR_c_1484_n 0.005155f $X=11.495 $Y=2.4 $X2=0
+ $Y2=0
cc_831 N_A_2022_94#_c_1345_n N_VPWR_c_1493_n 0.0106591f $X=10.285 $Y=1.985 $X2=0
+ $Y2=0
cc_832 N_A_2022_94#_M1026_g N_VPWR_c_1494_n 0.00460063f $X=11.045 $Y=2.4 $X2=0
+ $Y2=0
cc_833 N_A_2022_94#_M1029_g N_VPWR_c_1494_n 0.0048691f $X=11.495 $Y=2.4 $X2=0
+ $Y2=0
cc_834 N_A_2022_94#_M1026_g N_VPWR_c_1475_n 0.00908554f $X=11.045 $Y=2.4 $X2=0
+ $Y2=0
cc_835 N_A_2022_94#_M1029_g N_VPWR_c_1475_n 0.00875947f $X=11.495 $Y=2.4 $X2=0
+ $Y2=0
cc_836 N_A_2022_94#_c_1345_n N_VPWR_c_1475_n 0.0122002f $X=10.285 $Y=1.985 $X2=0
+ $Y2=0
cc_837 N_A_2022_94#_M1005_g N_Q_c_1629_n 0.00735215f $X=11.05 $Y=0.74 $X2=0
+ $Y2=0
cc_838 N_A_2022_94#_M1025_g N_Q_c_1629_n 0.00930275f $X=11.48 $Y=0.74 $X2=0
+ $Y2=0
cc_839 N_A_2022_94#_M1026_g N_Q_c_1632_n 3.85373e-19 $X=11.045 $Y=2.4 $X2=0
+ $Y2=0
cc_840 N_A_2022_94#_M1029_g N_Q_c_1632_n 0.0126857f $X=11.495 $Y=2.4 $X2=0 $Y2=0
cc_841 N_A_2022_94#_M1026_g N_Q_c_1630_n 0.00293165f $X=11.045 $Y=2.4 $X2=0
+ $Y2=0
cc_842 N_A_2022_94#_M1005_g N_Q_c_1630_n 0.00247818f $X=11.05 $Y=0.74 $X2=0
+ $Y2=0
cc_843 N_A_2022_94#_M1025_g N_Q_c_1630_n 0.00892862f $X=11.48 $Y=0.74 $X2=0
+ $Y2=0
cc_844 N_A_2022_94#_M1029_g N_Q_c_1630_n 0.00994275f $X=11.495 $Y=2.4 $X2=0
+ $Y2=0
cc_845 N_A_2022_94#_c_1340_n N_Q_c_1630_n 0.0249855f $X=10.975 $Y=1.465 $X2=0
+ $Y2=0
cc_846 N_A_2022_94#_c_1342_n N_Q_c_1630_n 0.0231811f $X=11.495 $Y=1.465 $X2=0
+ $Y2=0
cc_847 N_A_2022_94#_M1005_g N_Q_c_1631_n 0.00245603f $X=11.05 $Y=0.74 $X2=0
+ $Y2=0
cc_848 N_A_2022_94#_M1025_g N_Q_c_1631_n 0.00259764f $X=11.48 $Y=0.74 $X2=0
+ $Y2=0
cc_849 N_A_2022_94#_c_1340_n N_Q_c_1631_n 0.00191579f $X=10.975 $Y=1.465 $X2=0
+ $Y2=0
cc_850 N_A_2022_94#_c_1342_n N_Q_c_1631_n 0.00359474f $X=11.495 $Y=1.465 $X2=0
+ $Y2=0
cc_851 N_A_2022_94#_M1029_g Q 0.00478479f $X=11.495 $Y=2.4 $X2=0 $Y2=0
cc_852 N_A_2022_94#_c_1342_n Q 0.00304448f $X=11.495 $Y=1.465 $X2=0 $Y2=0
cc_853 N_A_2022_94#_M1026_g N_Q_c_1635_n 0.0201096f $X=11.045 $Y=2.4 $X2=0 $Y2=0
cc_854 N_A_2022_94#_c_1345_n N_Q_c_1635_n 0.0212714f $X=10.285 $Y=1.985 $X2=0
+ $Y2=0
cc_855 N_A_2022_94#_c_1340_n N_Q_c_1635_n 0.0318525f $X=10.975 $Y=1.465 $X2=0
+ $Y2=0
cc_856 N_A_2022_94#_c_1342_n N_Q_c_1635_n 0.00326486f $X=11.495 $Y=1.465 $X2=0
+ $Y2=0
cc_857 N_A_2022_94#_M1005_g N_VGND_c_1673_n 0.00946427f $X=11.05 $Y=0.74 $X2=0
+ $Y2=0
cc_858 N_A_2022_94#_c_1339_n N_VGND_c_1673_n 0.0258905f $X=10.255 $Y=0.615 $X2=0
+ $Y2=0
cc_859 N_A_2022_94#_c_1340_n N_VGND_c_1673_n 0.0285241f $X=10.975 $Y=1.465 $X2=0
+ $Y2=0
cc_860 N_A_2022_94#_c_1342_n N_VGND_c_1673_n 0.00277218f $X=11.495 $Y=1.465
+ $X2=0 $Y2=0
cc_861 N_A_2022_94#_M1025_g N_VGND_c_1675_n 0.00842499f $X=11.48 $Y=0.74 $X2=0
+ $Y2=0
cc_862 N_A_2022_94#_c_1339_n N_VGND_c_1680_n 0.0103491f $X=10.255 $Y=0.615 $X2=0
+ $Y2=0
cc_863 N_A_2022_94#_M1005_g N_VGND_c_1681_n 0.00434272f $X=11.05 $Y=0.74 $X2=0
+ $Y2=0
cc_864 N_A_2022_94#_M1025_g N_VGND_c_1681_n 0.00394617f $X=11.48 $Y=0.74 $X2=0
+ $Y2=0
cc_865 N_A_2022_94#_M1005_g N_VGND_c_1687_n 0.00825059f $X=11.05 $Y=0.74 $X2=0
+ $Y2=0
cc_866 N_A_2022_94#_M1025_g N_VGND_c_1687_n 0.00696181f $X=11.48 $Y=0.74 $X2=0
+ $Y2=0
cc_867 N_A_2022_94#_c_1339_n N_VGND_c_1687_n 0.0113354f $X=10.255 $Y=0.615 $X2=0
+ $Y2=0
cc_868 N_A_27_74#_c_1412_n N_VPWR_M1014_d 9.71305e-19 $X=2.445 $Y=2.145 $X2=0
+ $Y2=0
cc_869 N_A_27_74#_c_1459_n N_VPWR_M1014_d 0.00499461f $X=1.71 $Y=2.145 $X2=0
+ $Y2=0
cc_870 N_A_27_74#_c_1410_n N_VPWR_c_1476_n 0.0158217f $X=0.28 $Y=2.75 $X2=0
+ $Y2=0
cc_871 N_A_27_74#_c_1411_n N_VPWR_c_1476_n 0.0274627f $X=1.625 $Y=2.275 $X2=0
+ $Y2=0
cc_872 N_A_27_74#_c_1411_n N_VPWR_c_1477_n 0.00220908f $X=1.625 $Y=2.275 $X2=0
+ $Y2=0
cc_873 N_A_27_74#_c_1412_n N_VPWR_c_1477_n 0.00262985f $X=2.445 $Y=2.145 $X2=0
+ $Y2=0
cc_874 N_A_27_74#_c_1459_n N_VPWR_c_1477_n 0.0112212f $X=1.71 $Y=2.145 $X2=0
+ $Y2=0
cc_875 N_A_27_74#_c_1410_n N_VPWR_c_1488_n 0.011066f $X=0.28 $Y=2.75 $X2=0 $Y2=0
cc_876 N_A_27_74#_c_1410_n N_VPWR_c_1475_n 0.00915947f $X=0.28 $Y=2.75 $X2=0
+ $Y2=0
cc_877 N_A_27_74#_c_1407_n N_VGND_c_1676_n 0.00897649f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_878 N_A_27_74#_c_1407_n N_VGND_c_1687_n 0.00884022f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_879 N_VPWR_c_1482_n N_Q_c_1632_n 0.0255478f $X=10.82 $Y=2.405 $X2=0 $Y2=0
cc_880 N_VPWR_c_1484_n N_Q_c_1632_n 0.0315676f $X=11.72 $Y=1.985 $X2=0 $Y2=0
cc_881 N_VPWR_c_1494_n N_Q_c_1632_n 0.0135669f $X=11.635 $Y=3.33 $X2=0 $Y2=0
cc_882 N_VPWR_c_1475_n N_Q_c_1632_n 0.0110909f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_883 N_VPWR_c_1484_n Q 0.0146621f $X=11.72 $Y=1.985 $X2=0 $Y2=0
cc_884 N_VPWR_M1006_d N_Q_c_1635_n 0.00684067f $X=10.6 $Y=1.84 $X2=0 $Y2=0
cc_885 N_VPWR_c_1482_n N_Q_c_1635_n 0.0204127f $X=10.82 $Y=2.405 $X2=0 $Y2=0
cc_886 N_Q_c_1629_n N_VGND_c_1673_n 0.0312654f $X=11.265 $Y=0.515 $X2=0 $Y2=0
cc_887 N_Q_c_1629_n N_VGND_c_1675_n 0.0597505f $X=11.265 $Y=0.515 $X2=0 $Y2=0
cc_888 N_Q_c_1629_n N_VGND_c_1681_n 0.0159493f $X=11.265 $Y=0.515 $X2=0 $Y2=0
cc_889 N_Q_c_1629_n N_VGND_c_1687_n 0.0130065f $X=11.265 $Y=0.515 $X2=0 $Y2=0

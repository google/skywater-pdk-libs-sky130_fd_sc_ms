* File: sky130_fd_sc_ms__a31o_4.pex.spice
* Created: Fri Aug 28 17:06:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A31O_4%A_83_274# 1 2 3 4 15 17 19 22 24 26 27 29 32
+ 34 36 39 41 51 53 54 59 61 65 72 73 75 85
c141 85 0 9.90067e-20 $X=1.955 $Y=1.385
c142 75 0 2.72384e-19 $X=3.405 $Y=1.13
c143 73 0 1.68626e-19 $X=3.35 $Y=1.97
c144 65 0 9.60428e-20 $X=4.585 $Y=0.76
c145 61 0 1.54719e-19 $X=4.42 $Y=1.195
c146 15 0 7.10079e-20 $X=0.505 $Y=2.4
r147 84 85 11.055 $w=3.27e-07 $l=7.5e-08 $layer=POLY_cond $X=1.88 $Y=1.385
+ $X2=1.955 $Y2=1.385
r148 81 82 11.792 $w=3.27e-07 $l=8e-08 $layer=POLY_cond $X=1.425 $Y=1.385
+ $X2=1.505 $Y2=1.385
r149 78 79 5.89602 $w=3.27e-07 $l=4e-08 $layer=POLY_cond $X=0.955 $Y=1.385
+ $X2=0.995 $Y2=1.385
r150 77 78 64.1193 $w=3.27e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=1.385
+ $X2=0.955 $Y2=1.385
r151 76 77 2.21101 $w=3.27e-07 $l=1.5e-08 $layer=POLY_cond $X=0.505 $Y=1.385
+ $X2=0.52 $Y2=1.385
r152 72 73 7.89515 $w=4.48e-07 $l=1.15e-07 $layer=LI1_cond $X=3.35 $Y=2.085
+ $X2=3.35 $Y2=1.97
r153 69 85 31.6911 $w=3.27e-07 $l=2.15e-07 $layer=POLY_cond $X=2.17 $Y=1.385
+ $X2=1.955 $Y2=1.385
r154 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.17
+ $Y=1.385 $X2=2.17 $Y2=1.385
r155 63 65 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=4.585 $Y=1.11
+ $X2=4.585 $Y2=0.76
r156 62 75 4.30018 $w=1.7e-07 $l=3.76098e-07 $layer=LI1_cond $X=3.75 $Y=1.195
+ $X2=3.405 $Y2=1.13
r157 61 63 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.42 $Y=1.195
+ $X2=4.585 $Y2=1.11
r158 61 62 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.42 $Y=1.195
+ $X2=3.75 $Y2=1.195
r159 57 75 1.96316 $w=3.3e-07 $l=1.89737e-07 $layer=LI1_cond $X=3.585 $Y=1.11
+ $X2=3.405 $Y2=1.13
r160 57 59 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=3.585 $Y=1.11
+ $X2=3.585 $Y2=0.515
r161 55 75 1.96316 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.49 $Y=1.3
+ $X2=3.405 $Y2=1.13
r162 55 73 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.49 $Y=1.3
+ $X2=3.49 $Y2=1.97
r163 53 75 4.30018 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.405 $Y=1.215
+ $X2=3.405 $Y2=1.13
r164 53 54 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.405 $Y=1.215
+ $X2=2.74 $Y2=1.215
r165 49 54 7.35534 $w=3e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.615 $Y=1.13
+ $X2=2.74 $Y2=1.215
r166 49 68 18.0967 $w=3e-07 $l=5.39884e-07 $layer=LI1_cond $X=2.615 $Y=1.13
+ $X2=2.17 $Y2=1.34
r167 49 51 28.3501 $w=2.48e-07 $l=6.15e-07 $layer=LI1_cond $X=2.615 $Y=1.13
+ $X2=2.615 $Y2=0.515
r168 48 84 7.37003 $w=3.27e-07 $l=5e-08 $layer=POLY_cond $X=1.83 $Y=1.385
+ $X2=1.88 $Y2=1.385
r169 48 82 47.9052 $w=3.27e-07 $l=3.25e-07 $layer=POLY_cond $X=1.83 $Y=1.385
+ $X2=1.505 $Y2=1.385
r170 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.83
+ $Y=1.385 $X2=1.83 $Y2=1.385
r171 44 81 40.5352 $w=3.27e-07 $l=2.75e-07 $layer=POLY_cond $X=1.15 $Y=1.385
+ $X2=1.425 $Y2=1.385
r172 44 79 22.8471 $w=3.27e-07 $l=1.55e-07 $layer=POLY_cond $X=1.15 $Y=1.385
+ $X2=0.995 $Y2=1.385
r173 43 47 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.15 $Y=1.385
+ $X2=1.83 $Y2=1.385
r174 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.385 $X2=1.15 $Y2=1.385
r175 41 68 10.2918 $w=3.3e-07 $l=2.96648e-07 $layer=LI1_cond $X=1.895 $Y=1.385
+ $X2=2.17 $Y2=1.34
r176 41 47 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=1.895 $Y=1.385
+ $X2=1.83 $Y2=1.385
r177 37 85 16.7191 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.955 $Y=1.55
+ $X2=1.955 $Y2=1.385
r178 37 39 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.955 $Y=1.55
+ $X2=1.955 $Y2=2.4
r179 34 84 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.88 $Y=1.22
+ $X2=1.88 $Y2=1.385
r180 34 36 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.88 $Y=1.22
+ $X2=1.88 $Y2=0.74
r181 30 82 16.7191 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.505 $Y=1.55
+ $X2=1.505 $Y2=1.385
r182 30 32 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.505 $Y=1.55
+ $X2=1.505 $Y2=2.4
r183 27 81 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.22
+ $X2=1.425 $Y2=1.385
r184 27 29 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.425 $Y=1.22
+ $X2=1.425 $Y2=0.74
r185 24 79 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.22
+ $X2=0.995 $Y2=1.385
r186 24 26 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.995 $Y=1.22
+ $X2=0.995 $Y2=0.74
r187 20 78 16.7191 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.55
+ $X2=0.955 $Y2=1.385
r188 20 22 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.955 $Y=1.55
+ $X2=0.955 $Y2=2.4
r189 17 77 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=1.22
+ $X2=0.52 $Y2=1.385
r190 17 19 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.52 $Y=1.22
+ $X2=0.52 $Y2=0.74
r191 13 76 16.7191 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.55
+ $X2=0.505 $Y2=1.385
r192 13 15 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.505 $Y=1.55
+ $X2=0.505 $Y2=2.4
r193 4 72 300 $w=1.7e-07 $l=2.498e-07 $layer=licon1_PDIFF $count=2 $X=3.105
+ $Y=1.96 $X2=3.3 $Y2=2.085
r194 3 65 182 $w=1.7e-07 $l=4.83735e-07 $layer=licon1_NDIFF $count=1 $X=4.375
+ $Y=0.37 $X2=4.585 $Y2=0.76
r195 2 59 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.445
+ $Y=0.37 $X2=3.585 $Y2=0.515
r196 1 51 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=2.51
+ $Y=0.37 $X2=2.655 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A31O_4%B1 3 7 11 15 17 24
c61 24 0 7.22101e-20 $X=3.37 $Y=1.635
c62 17 0 9.90067e-20 $X=3.12 $Y=1.665
c63 3 0 9.37482e-20 $X=2.87 $Y=0.69
r64 22 24 48.3612 $w=2.99e-07 $l=3e-07 $layer=POLY_cond $X=3.07 $Y=1.635
+ $X2=3.37 $Y2=1.635
r65 20 22 8.86622 $w=2.99e-07 $l=5.5e-08 $layer=POLY_cond $X=3.015 $Y=1.635
+ $X2=3.07 $Y2=1.635
r66 19 20 23.3746 $w=2.99e-07 $l=1.45e-07 $layer=POLY_cond $X=2.87 $Y=1.635
+ $X2=3.015 $Y2=1.635
r67 17 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.07
+ $Y=1.635 $X2=3.07 $Y2=1.635
r68 13 24 26.5987 $w=2.99e-07 $l=2.33345e-07 $layer=POLY_cond $X=3.535 $Y=1.8
+ $X2=3.37 $Y2=1.635
r69 13 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.535 $Y=1.8
+ $X2=3.535 $Y2=2.46
r70 9 24 18.89 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.37 $Y=1.47 $X2=3.37
+ $Y2=1.635
r71 9 11 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=3.37 $Y=1.47 $X2=3.37
+ $Y2=0.69
r72 5 20 14.6425 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.015 $Y=1.8
+ $X2=3.015 $Y2=1.635
r73 5 7 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.015 $Y=1.8 $X2=3.015
+ $Y2=2.46
r74 1 19 18.89 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.87 $Y=1.47 $X2=2.87
+ $Y2=1.635
r75 1 3 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.87 $Y=1.47 $X2=2.87
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__A31O_4%A1 1 3 4 5 7 10 12 14 17 19 20 21 30
c67 10 0 1.68626e-19 $X=4.135 $Y=2.46
r68 28 30 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=4.55 $Y=1.615
+ $X2=4.685 $Y2=1.615
r69 26 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.21 $Y=1.615
+ $X2=4.55 $Y2=1.615
r70 24 26 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.135 $Y=1.615
+ $X2=4.21 $Y2=1.615
r71 21 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.55
+ $Y=1.615 $X2=4.55 $Y2=1.615
r72 20 21 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=4.08 $Y=1.615
+ $X2=4.55 $Y2=1.615
r73 15 30 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.685 $Y=1.78
+ $X2=4.685 $Y2=1.615
r74 15 17 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=4.685 $Y=1.78
+ $X2=4.685 $Y2=2.46
r75 12 19 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.3 $Y=1.085
+ $X2=4.21 $Y2=1.16
r76 12 14 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.3 $Y=1.085
+ $X2=4.3 $Y2=0.69
r77 8 24 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.135 $Y=1.78
+ $X2=4.135 $Y2=1.615
r78 8 10 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=4.135 $Y=1.78
+ $X2=4.135 $Y2=2.46
r79 7 26 2.83073 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.21 $Y=1.45
+ $X2=4.21 $Y2=1.615
r80 6 19 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=4.21 $Y=1.235
+ $X2=4.21 $Y2=1.16
r81 6 7 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=4.21 $Y=1.235
+ $X2=4.21 $Y2=1.45
r82 4 19 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.045 $Y=1.16
+ $X2=4.21 $Y2=1.16
r83 4 5 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.045 $Y=1.16
+ $X2=3.875 $Y2=1.16
r84 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.8 $Y=1.085
+ $X2=3.875 $Y2=1.16
r85 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.8 $Y=1.085 $X2=3.8
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__A31O_4%A2 3 6 7 9 11 14 18 20 23 25 26 30 31
c68 23 0 9.60428e-20 $X=5.36 $Y=1.16
c69 20 0 1.63311e-19 $X=5.045 $Y=1.6
c70 18 0 1.03588e-19 $X=5.79 $Y=0.69
r71 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.7
+ $Y=1.615 $X2=5.7 $Y2=1.615
r72 26 31 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=5.52 $Y=1.615
+ $X2=5.7 $Y2=1.615
r73 25 26 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.615
+ $X2=5.52 $Y2=1.615
r74 21 23 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.15 $Y=1.16
+ $X2=5.36 $Y2=1.16
r75 16 30 34.7346 $w=1.65e-07 $l=1.90526e-07 $layer=POLY_cond $X=5.79 $Y=1.45
+ $X2=5.735 $Y2=1.615
r76 16 18 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=5.79 $Y=1.45
+ $X2=5.79 $Y2=0.69
r77 12 30 34.7346 $w=1.65e-07 $l=1.83916e-07 $layer=POLY_cond $X=5.695 $Y=1.78
+ $X2=5.735 $Y2=1.615
r78 12 14 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=5.695 $Y=1.78
+ $X2=5.695 $Y2=2.46
r79 9 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.36 $Y=1.085
+ $X2=5.36 $Y2=1.16
r80 9 11 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.36 $Y=1.085
+ $X2=5.36 $Y2=0.69
r81 8 20 3.90195 $w=3.3e-07 $l=1.8735e-07 $layer=POLY_cond $X=5.225 $Y=1.615
+ $X2=5.045 $Y2=1.6
r82 7 30 3.90195 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=5.605 $Y=1.615
+ $X2=5.735 $Y2=1.615
r83 7 8 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=5.605 $Y=1.615
+ $X2=5.225 $Y2=1.615
r84 6 20 34.7346 $w=1.65e-07 $l=1.95576e-07 $layer=POLY_cond $X=5.15 $Y=1.45
+ $X2=5.045 $Y2=1.6
r85 5 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.15 $Y=1.235
+ $X2=5.15 $Y2=1.16
r86 5 6 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=5.15 $Y=1.235
+ $X2=5.15 $Y2=1.45
r87 1 20 34.7346 $w=1.65e-07 $l=2.20454e-07 $layer=POLY_cond $X=5.135 $Y=1.78
+ $X2=5.045 $Y2=1.6
r88 1 3 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=5.135 $Y=1.78
+ $X2=5.135 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A31O_4%A3 3 7 11 15 17 18 28
c41 3 0 1.72297e-19 $X=6.195 $Y=2.46
r42 27 28 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=6.65 $Y=1.615
+ $X2=6.695 $Y2=1.615
r43 25 27 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=6.62 $Y=1.615 $X2=6.65
+ $Y2=1.615
r44 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.62
+ $Y=1.615 $X2=6.62 $Y2=1.615
r45 23 25 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=6.22 $Y=1.615 $X2=6.62
+ $Y2=1.615
r46 21 23 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=6.195 $Y=1.615
+ $X2=6.22 $Y2=1.615
r47 18 26 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=6.96 $Y=1.615
+ $X2=6.62 $Y2=1.615
r48 17 26 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=6.48 $Y=1.615
+ $X2=6.62 $Y2=1.615
r49 13 28 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.695 $Y=1.78
+ $X2=6.695 $Y2=1.615
r50 13 15 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=6.695 $Y=1.78
+ $X2=6.695 $Y2=2.46
r51 9 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.65 $Y=1.45
+ $X2=6.65 $Y2=1.615
r52 9 11 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=6.65 $Y=1.45 $X2=6.65
+ $Y2=0.69
r53 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.22 $Y=1.45
+ $X2=6.22 $Y2=1.615
r54 5 7 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=6.22 $Y=1.45 $X2=6.22
+ $Y2=0.69
r55 1 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.195 $Y=1.78
+ $X2=6.195 $Y2=1.615
r56 1 3 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=6.195 $Y=1.78
+ $X2=6.195 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A31O_4%VPWR 1 2 3 4 5 6 19 21 27 33 39 43 47 50 51
+ 53 54 55 57 62 77 83 84 90 93 96
r95 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r96 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r97 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r98 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r99 84 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r100 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r101 81 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.585 $Y=3.33
+ $X2=6.42 $Y2=3.33
r102 81 83 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.585 $Y=3.33
+ $X2=6.96 $Y2=3.33
r103 80 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r104 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r105 77 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.255 $Y=3.33
+ $X2=6.42 $Y2=3.33
r106 77 79 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.255 $Y=3.33
+ $X2=6 $Y2=3.33
r107 76 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r108 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r109 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r110 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r111 70 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r112 69 72 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r113 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r114 67 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.23 $Y2=3.33
r115 67 69 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.64 $Y2=3.33
r116 66 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r117 66 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r118 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r119 63 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.23 $Y2=3.33
r120 63 65 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.68 $Y2=3.33
r121 62 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=2.23 $Y2=3.33
r122 62 65 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=1.68 $Y2=3.33
r123 61 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r124 61 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r125 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r126 58 87 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r127 58 60 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r128 57 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.23 $Y2=3.33
r129 57 60 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.72 $Y2=3.33
r130 55 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r131 55 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r132 53 75 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.245 $Y=3.33
+ $X2=5.04 $Y2=3.33
r133 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.245 $Y=3.33
+ $X2=5.41 $Y2=3.33
r134 52 79 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=5.575 $Y=3.33
+ $X2=6 $Y2=3.33
r135 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.575 $Y=3.33
+ $X2=5.41 $Y2=3.33
r136 50 72 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.245 $Y=3.33
+ $X2=4.08 $Y2=3.33
r137 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.245 $Y=3.33
+ $X2=4.41 $Y2=3.33
r138 49 75 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=4.575 $Y=3.33
+ $X2=5.04 $Y2=3.33
r139 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.575 $Y=3.33
+ $X2=4.41 $Y2=3.33
r140 45 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=3.245
+ $X2=6.42 $Y2=3.33
r141 45 47 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=6.42 $Y=3.245
+ $X2=6.42 $Y2=2.425
r142 41 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.41 $Y=3.245
+ $X2=5.41 $Y2=3.33
r143 41 43 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=5.41 $Y=3.245
+ $X2=5.41 $Y2=2.425
r144 37 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.41 $Y=3.245
+ $X2=4.41 $Y2=3.33
r145 37 39 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=4.41 $Y=3.245
+ $X2=4.41 $Y2=2.425
r146 33 36 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.23 $Y=1.985
+ $X2=2.23 $Y2=2.815
r147 31 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=3.245
+ $X2=2.23 $Y2=3.33
r148 31 36 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.23 $Y=3.245
+ $X2=2.23 $Y2=2.815
r149 27 30 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.23 $Y=2.145
+ $X2=1.23 $Y2=2.825
r150 25 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=3.33
r151 25 30 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=2.825
r152 21 24 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r153 19 87 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r154 19 24 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r155 6 47 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=6.285
+ $Y=1.96 $X2=6.42 $Y2=2.425
r156 5 43 300 $w=1.7e-07 $l=5.49773e-07 $layer=licon1_PDIFF $count=2 $X=5.225
+ $Y=1.96 $X2=5.41 $Y2=2.425
r157 4 39 300 $w=1.7e-07 $l=5.49773e-07 $layer=licon1_PDIFF $count=2 $X=4.225
+ $Y=1.96 $X2=4.41 $Y2=2.425
r158 3 36 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.84 $X2=2.23 $Y2=2.815
r159 3 33 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.84 $X2=2.23 $Y2=1.985
r160 2 30 400 $w=1.7e-07 $l=1.07352e-06 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.23 $Y2=2.825
r161 2 27 400 $w=1.7e-07 $l=3.86588e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.23 $Y2=2.145
r162 1 24 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r163 1 21 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__A31O_4%X 1 2 3 4 15 19 21 25 29 35 36 37 38 54
c57 21 0 1.43218e-19 $X=1.565 $Y=1.805
r58 43 56 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.89
+ $X2=0.73 $Y2=1.805
r59 37 38 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.73 $Y=2.405
+ $X2=0.73 $Y2=2.775
r60 36 37 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=0.73 $Y=1.985
+ $X2=0.73 $Y2=2.405
r61 36 43 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.73 $Y=1.985
+ $X2=0.73 $Y2=1.89
r62 35 56 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=1.805
r63 35 54 4.72076 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=1.55
r64 29 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.73 $Y=1.985
+ $X2=1.73 $Y2=2.815
r65 27 29 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.73 $Y=1.89
+ $X2=1.73 $Y2=1.985
r66 23 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.64 $Y=0.83
+ $X2=1.64 $Y2=0.495
r67 22 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=1.805
+ $X2=0.73 $Y2=1.805
r68 21 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.565 $Y=1.805
+ $X2=1.73 $Y2=1.89
r69 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.565 $Y=1.805
+ $X2=0.895 $Y2=1.805
r70 20 34 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.865 $Y=0.915
+ $X2=0.74 $Y2=0.915
r71 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.555 $Y=0.915
+ $X2=1.64 $Y2=0.83
r72 19 20 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.555 $Y=0.915
+ $X2=0.865 $Y2=0.915
r73 17 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=1 $X2=0.74
+ $Y2=0.915
r74 17 54 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=0.74 $Y=1 $X2=0.74
+ $Y2=1.55
r75 13 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0.83 $X2=0.74
+ $Y2=0.915
r76 13 15 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=0.74 $Y=0.83
+ $X2=0.74 $Y2=0.515
r77 4 31 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.84 $X2=1.73 $Y2=2.815
r78 4 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.84 $X2=1.73 $Y2=1.985
r79 3 38 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.815
r80 3 36 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=1.985
r81 2 25 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.5
+ $Y=0.37 $X2=1.64 $Y2=0.495
r82 1 34 182 $w=1.7e-07 $l=6.81249e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.37 $X2=0.78 $Y2=0.965
r83 1 15 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A31O_4%A_529_392# 1 2 3 4 5 16 18 20 22 23 24 28 30
+ 34 36 38 40 49 51
c90 49 0 1.54719e-19 $X=4.91 $Y=2.115
c91 36 0 1.47061e-19 $X=6.755 $Y=2.035
c92 34 0 1.72297e-19 $X=5.92 $Y=2.815
c93 22 0 1.78636e-19 $X=3.91 $Y=2.12
r94 38 53 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.92 $Y=2.12 $X2=6.92
+ $Y2=2.035
r95 38 40 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=6.92 $Y=2.12
+ $X2=6.92 $Y2=2.815
r96 37 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.085 $Y=2.035
+ $X2=5.92 $Y2=2.035
r97 36 53 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.755 $Y=2.035
+ $X2=6.92 $Y2=2.035
r98 36 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.755 $Y=2.035
+ $X2=6.085 $Y2=2.035
r99 32 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=2.12 $X2=5.92
+ $Y2=2.035
r100 32 34 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.92 $Y=2.12
+ $X2=5.92 $Y2=2.815
r101 31 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.075 $Y=2.035
+ $X2=4.91 $Y2=2.035
r102 30 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.755 $Y=2.035
+ $X2=5.92 $Y2=2.035
r103 30 31 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.755 $Y=2.035
+ $X2=5.075 $Y2=2.035
r104 26 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.91 $Y=2.12
+ $X2=4.91 $Y2=2.035
r105 26 28 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.91 $Y=2.12
+ $X2=4.91 $Y2=2.815
r106 25 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.075 $Y=2.035
+ $X2=3.91 $Y2=2.035
r107 24 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.745 $Y=2.035
+ $X2=4.91 $Y2=2.035
r108 24 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.745 $Y=2.035
+ $X2=4.075 $Y2=2.035
r109 23 47 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.91 $Y=2.81 $X2=3.91
+ $Y2=2.895
r110 22 45 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.91 $Y=2.12 $X2=3.91
+ $Y2=2.035
r111 22 23 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=3.91 $Y=2.12
+ $X2=3.91 $Y2=2.81
r112 21 43 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.955 $Y=2.895
+ $X2=2.79 $Y2=2.895
r113 20 47 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.745 $Y=2.895
+ $X2=3.91 $Y2=2.895
r114 20 21 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=3.745 $Y=2.895
+ $X2=2.955 $Y2=2.895
r115 16 43 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.79 $Y=2.81 $X2=2.79
+ $Y2=2.895
r116 16 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.79 $Y=2.81
+ $X2=2.79 $Y2=2.135
r117 5 53 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=6.785
+ $Y=1.96 $X2=6.92 $Y2=2.115
r118 5 40 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.785
+ $Y=1.96 $X2=6.92 $Y2=2.815
r119 4 51 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=5.785
+ $Y=1.96 $X2=5.92 $Y2=2.115
r120 4 34 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.785
+ $Y=1.96 $X2=5.92 $Y2=2.815
r121 3 49 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=4.775
+ $Y=1.96 $X2=4.91 $Y2=2.115
r122 3 28 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.775
+ $Y=1.96 $X2=4.91 $Y2=2.815
r123 2 47 400 $w=1.7e-07 $l=9.87269e-07 $layer=licon1_PDIFF $count=1 $X=3.625
+ $Y=1.96 $X2=3.91 $Y2=2.815
r124 2 45 400 $w=1.7e-07 $l=3.54119e-07 $layer=licon1_PDIFF $count=1 $X=3.625
+ $Y=1.96 $X2=3.91 $Y2=2.115
r125 1 43 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.645
+ $Y=1.96 $X2=2.79 $Y2=2.815
r126 1 18 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.645
+ $Y=1.96 $X2=2.79 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_MS__A31O_4%VGND 1 2 3 4 5 16 18 22 26 30 34 36 38 43 48
+ 53 63 64 70 73 76 79
r90 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r91 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r92 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r93 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r94 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r95 64 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r96 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r97 61 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.6 $Y=0 $X2=6.435
+ $Y2=0
r98 61 63 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.6 $Y=0 $X2=6.96
+ $Y2=0
r99 60 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r100 59 60 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=0 $X2=6 $Y2=0
r101 56 59 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=6
+ $Y2=0
r102 54 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.25 $Y=0 $X2=3.085
+ $Y2=0
r103 54 56 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.25 $Y=0 $X2=3.6
+ $Y2=0
r104 53 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.27 $Y=0 $X2=6.435
+ $Y2=0
r105 53 59 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.27 $Y=0 $X2=6
+ $Y2=0
r106 52 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r107 52 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r108 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r109 49 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=0 $X2=2.095
+ $Y2=0
r110 49 51 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.26 $Y=0 $X2=2.64
+ $Y2=0
r111 48 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.92 $Y=0 $X2=3.085
+ $Y2=0
r112 48 51 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.92 $Y=0 $X2=2.64
+ $Y2=0
r113 47 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r114 47 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r115 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r116 44 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.21
+ $Y2=0
r117 44 46 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.375 $Y=0
+ $X2=1.68 $Y2=0
r118 43 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.93 $Y=0 $X2=2.095
+ $Y2=0
r119 43 46 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.93 $Y=0 $X2=1.68
+ $Y2=0
r120 42 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r121 42 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r122 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r123 39 67 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r124 39 41 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r125 38 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.21
+ $Y2=0
r126 38 41 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=0
+ $X2=0.72 $Y2=0
r127 36 60 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=6
+ $Y2=0
r128 36 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r129 36 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r130 32 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.435 $Y=0.085
+ $X2=6.435 $Y2=0
r131 32 34 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.435 $Y=0.085
+ $X2=6.435 $Y2=0.495
r132 28 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=0.085
+ $X2=3.085 $Y2=0
r133 28 30 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.085 $Y=0.085
+ $X2=3.085 $Y2=0.495
r134 24 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.095 $Y=0.085
+ $X2=2.095 $Y2=0
r135 24 26 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.095 $Y=0.085
+ $X2=2.095 $Y2=0.515
r136 20 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0
r137 20 22 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0.565
r138 16 67 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r139 16 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.515
r140 5 34 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=6.295
+ $Y=0.37 $X2=6.435 $Y2=0.495
r141 4 30 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.945
+ $Y=0.37 $X2=3.085 $Y2=0.495
r142 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.955
+ $Y=0.37 $X2=2.095 $Y2=0.515
r143 2 22 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.21 $Y2=0.565
r144 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A31O_4%A_775_74# 1 2 9 11 12 15
r27 13 15 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=5.575 $Y=0.425
+ $X2=5.575 $Y2=0.495
r28 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.41 $Y=0.34
+ $X2=5.575 $Y2=0.425
r29 11 12 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=5.41 $Y=0.34
+ $X2=4.25 $Y2=0.34
r30 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.085 $Y=0.425
+ $X2=4.25 $Y2=0.34
r31 7 9 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=4.085 $Y=0.425 $X2=4.085
+ $Y2=0.495
r32 2 15 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=5.435
+ $Y=0.37 $X2=5.575 $Y2=0.495
r33 1 9 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=3.875
+ $Y=0.37 $X2=4.085 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_MS__A31O_4%A_1000_74# 1 2 3 12 14 15 18 20 24 26
c40 26 0 1.47061e-19 $X=6.005 $Y=1.195
c41 15 0 1.63311e-19 $X=5.23 $Y=1.195
c42 12 0 1.03588e-19 $X=5.145 $Y=0.76
r43 22 24 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=6.905 $Y=1.11
+ $X2=6.905 $Y2=0.515
r44 21 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.09 $Y=1.195
+ $X2=6.005 $Y2=1.195
r45 20 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.78 $Y=1.195
+ $X2=6.905 $Y2=1.11
r46 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.78 $Y=1.195
+ $X2=6.09 $Y2=1.195
r47 16 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=1.11
+ $X2=6.005 $Y2=1.195
r48 16 18 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=6.005 $Y=1.11
+ $X2=6.005 $Y2=0.515
r49 14 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=1.195
+ $X2=6.005 $Y2=1.195
r50 14 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.92 $Y=1.195
+ $X2=5.23 $Y2=1.195
r51 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.105 $Y=1.11
+ $X2=5.23 $Y2=1.195
r52 10 12 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=5.105 $Y=1.11
+ $X2=5.105 $Y2=0.76
r53 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.725
+ $Y=0.37 $X2=6.865 $Y2=0.515
r54 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.865
+ $Y=0.37 $X2=6.005 $Y2=0.515
r55 1 12 182 $w=1.7e-07 $l=4.56782e-07 $layer=licon1_NDIFF $count=1 $X=5 $Y=0.37
+ $X2=5.145 $Y2=0.76
.ends


* File: sky130_fd_sc_ms__or3b_2.spice
* Created: Fri Aug 28 18:08:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__or3b_2.pex.spice"
.subckt sky130_fd_sc_ms__or3b_2  VNB VPB C_N A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_C_N_M1005_g N_A_27_368#_M1005_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.107506 AS=0.15675 PD=0.937984 PS=1.67 NRD=18.54 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75002.9 A=0.0825 P=1.4 MULT=1
MM1004 N_X_M1004_d N_A_190_260#_M1004_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.144644 PD=1.02 PS=1.26202 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1008 N_X_M1004_d N_A_190_260#_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.210739 PD=1.02 PS=1.41029 NRD=0 NRS=29.184 M=1 R=4.93333
+ SA=75001 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1007 N_A_190_260#_M1007_d N_A_M1007_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.182261 PD=0.99 PS=1.21971 NRD=13.116 NRS=21.552 M=1 R=4.26667
+ SA=75001.8 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1006_d N_B_M1006_g N_A_190_260#_M1007_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1344 AS=0.112 PD=1.06 PS=0.99 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75002.3
+ SB=75000.8 A=0.096 P=1.58 MULT=1
MM1000 N_A_190_260#_M1000_d N_A_27_368#_M1000_g N_VGND_M1006_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.1344 PD=1.85 PS=1.06 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75002.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1002 N_VPWR_M1002_d N_C_N_M1002_g N_A_27_368#_M1002_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1614 AS=0.2352 PD=1.26429 PS=2.24 NRD=32.1504 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90002.9 A=0.1512 P=2.04 MULT=1
MM1010 N_X_M1010_d N_A_190_260#_M1010_g N_VPWR_M1002_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2152 PD=1.39 PS=1.68571 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90002.2 A=0.2016 P=2.6 MULT=1
MM1011 N_X_M1010_d N_A_190_260#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.319808 PD=1.39 PS=1.76981 NRD=0 NRS=22.852 M=1 R=6.22222
+ SA=90001 SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1001 A_461_368# N_A_M1001_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.285542 PD=1.24 PS=1.58019 NRD=12.7853 NRS=27.5603 M=1 R=5.55556
+ SA=90001.8 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1003 A_545_368# N_B_M1003_g A_461_368# VPB PSHORT L=0.18 W=1 AD=0.18 AS=0.12
+ PD=1.36 PS=1.24 NRD=24.6053 NRS=12.7853 M=1 R=5.55556 SA=90002.2 SB=90000.7
+ A=0.18 P=2.36 MULT=1
MM1009 N_A_190_260#_M1009_d N_A_27_368#_M1009_g A_545_368# VPB PSHORT L=0.18 W=1
+ AD=0.28 AS=0.18 PD=2.56 PS=1.36 NRD=0 NRS=24.6053 M=1 R=5.55556 SA=90002.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ms__or3b_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__a22oi_1.pex.spice
* Created: Fri Aug 28 17:03:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A22OI_1%B2 3 5 7 8 9 10 11
r32 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r33 11 16 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=0.27 $Y=1.665
+ $X2=0.27 $Y2=1.385
r34 10 16 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.385
r35 8 15 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=0.615 $Y=1.385
+ $X2=0.27 $Y2=1.385
r36 8 9 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.615 $Y=1.385 $X2=0.705
+ $Y2=1.385
r37 5 9 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=0.72 $Y=1.22
+ $X2=0.705 $Y2=1.385
r38 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.72 $Y=1.22 $X2=0.72
+ $Y2=0.74
r39 1 9 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.705 $Y=1.55
+ $X2=0.705 $Y2=1.385
r40 1 3 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.705 $Y=1.55
+ $X2=0.705 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_1%B1 3 7 9 12 13
c38 12 0 3.57792e-20 $X=1.17 $Y=1.515
c39 7 0 1.10616e-19 $X=1.155 $Y=2.4
r40 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.515
+ $X2=1.17 $Y2=1.68
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.515
+ $X2=1.17 $Y2=1.35
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.515 $X2=1.17 $Y2=1.515
r43 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.17 $Y=1.665
+ $X2=1.17 $Y2=1.515
r44 7 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.155 $Y=2.4
+ $X2=1.155 $Y2=1.68
r45 3 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.08 $Y=0.74 $X2=1.08
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_1%A1 3 7 9 12 13
c35 13 0 1.10616e-19 $X=1.71 $Y=1.515
r36 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.71 $Y=1.515
+ $X2=1.71 $Y2=1.68
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.71 $Y=1.515
+ $X2=1.71 $Y2=1.35
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.515 $X2=1.71 $Y2=1.515
r39 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.71 $Y=1.665
+ $X2=1.71 $Y2=1.515
r40 7 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.635 $Y=2.4
+ $X2=1.635 $Y2=1.68
r41 3 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.62 $Y=0.74 $X2=1.62
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_1%A2 3 7 9 10 14
r30 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.515
+ $X2=2.25 $Y2=1.68
r31 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.515
+ $X2=2.25 $Y2=1.35
r32 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.515 $X2=2.25 $Y2=1.515
r33 10 15 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.25 $Y2=1.565
r34 9 15 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=2.16 $Y=1.565 $X2=2.25
+ $Y2=1.565
r35 7 17 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.175 $Y=2.4
+ $X2=2.175 $Y2=1.68
r36 3 16 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.16 $Y=0.74 $X2=2.16
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_1%A_71_368# 1 2 3 12 14 15 16 19 20 22 24
r41 22 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.4 $Y=2.12 $X2=2.4
+ $Y2=2.035
r42 22 24 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.4 $Y=2.12 $X2=2.4
+ $Y2=2.815
r43 21 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=2.035
+ $X2=1.38 $Y2=2.035
r44 20 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=2.035
+ $X2=2.4 $Y2=2.035
r45 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.235 $Y=2.035
+ $X2=1.545 $Y2=2.035
r46 17 19 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.38 $Y=2.905 $X2=1.38
+ $Y2=2.815
r47 16 27 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.38 $Y=2.12 $X2=1.38
+ $Y2=2.035
r48 16 19 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.38 $Y=2.12
+ $X2=1.38 $Y2=2.815
r49 14 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.215 $Y=2.99
+ $X2=1.38 $Y2=2.905
r50 14 15 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.215 $Y=2.99
+ $X2=0.645 $Y2=2.99
r51 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.48 $Y=2.905
+ $X2=0.645 $Y2=2.99
r52 10 12 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.48 $Y=2.905
+ $X2=0.48 $Y2=2.455
r53 3 29 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.265
+ $Y=1.84 $X2=2.4 $Y2=2.115
r54 3 24 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.265
+ $Y=1.84 $X2=2.4 $Y2=2.815
r55 2 27 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.245
+ $Y=1.84 $X2=1.38 $Y2=2.115
r56 2 19 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.245
+ $Y=1.84 $X2=1.38 $Y2=2.815
r57 1 12 300 $w=1.7e-07 $l=6.74611e-07 $layer=licon1_PDIFF $count=2 $X=0.355
+ $Y=1.84 $X2=0.48 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_1%Y 1 2 7 8 13 20 22 23
c36 20 0 3.57792e-20 $X=0.93 $Y=2.115
r37 22 23 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=1.295
+ $X2=0.72 $Y2=1.665
r38 17 23 14.2803 $w=2.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.72 $Y=1.95
+ $X2=0.72 $Y2=1.665
r39 17 20 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.72 $Y=2.035
+ $X2=0.93 $Y2=2.035
r40 15 22 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.72 $Y=1.18
+ $X2=0.72 $Y2=1.295
r41 11 13 12.965 $w=4.38e-07 $l=4.95e-07 $layer=LI1_cond $X=1.35 $Y=1.01
+ $X2=1.35 $Y2=0.515
r42 8 15 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.835 $Y=1.095
+ $X2=0.72 $Y2=1.18
r43 7 11 8.71846 $w=1.7e-07 $l=2.59037e-07 $layer=LI1_cond $X=1.13 $Y=1.095
+ $X2=1.35 $Y2=1.01
r44 7 8 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.13 $Y=1.095
+ $X2=0.835 $Y2=1.095
r45 2 20 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=0.795
+ $Y=1.84 $X2=0.93 $Y2=2.115
r46 1 13 91 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=2 $X=1.155
+ $Y=0.37 $X2=1.35 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_1%VPWR 1 6 9 10 11 21 22
r28 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r29 19 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r30 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r31 14 18 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r32 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 11 19 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r34 11 15 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.24 $Y2=3.33
r35 9 18 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=1.68 $Y2=3.33
r36 9 10 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.715 $Y=3.33 $X2=1.89
+ $Y2=3.33
r37 8 21 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.065 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 8 10 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.065 $Y=3.33 $X2=1.89
+ $Y2=3.33
r39 4 10 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.89 $Y=3.245 $X2=1.89
+ $Y2=3.33
r40 4 6 26.0123 $w=3.48e-07 $l=7.9e-07 $layer=LI1_cond $X=1.89 $Y=3.245 $X2=1.89
+ $Y2=2.455
r41 1 6 300 $w=1.7e-07 $l=6.92604e-07 $layer=licon1_PDIFF $count=2 $X=1.725
+ $Y=1.84 $X2=1.89 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__A22OI_1%VGND 1 2 9 13 16 17 19 20 21 34 35
r30 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r31 32 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r32 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r33 28 31 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r34 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r35 25 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r36 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r37 21 32 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r38 21 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r39 19 31 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.16
+ $Y2=0
r40 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.375
+ $Y2=0
r41 18 34 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.54 $Y=0 $X2=2.64
+ $Y2=0
r42 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.54 $Y=0 $X2=2.375
+ $Y2=0
r43 16 24 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.34 $Y=0 $X2=0.24
+ $Y2=0
r44 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.34 $Y=0 $X2=0.505
+ $Y2=0
r45 15 28 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=0.67 $Y=0 $X2=0.72
+ $Y2=0
r46 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.67 $Y=0 $X2=0.505
+ $Y2=0
r47 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=0.085
+ $X2=2.375 $Y2=0
r48 11 13 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.375 $Y=0.085
+ $X2=2.375 $Y2=0.515
r49 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.505 $Y=0.085
+ $X2=0.505 $Y2=0
r50 7 9 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.505 $Y=0.085
+ $X2=0.505 $Y2=0.675
r51 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.235
+ $Y=0.37 $X2=2.375 $Y2=0.515
r52 1 9 182 $w=1.7e-07 $l=3.62146e-07 $layer=licon1_NDIFF $count=1 $X=0.38
+ $Y=0.37 $X2=0.505 $Y2=0.675
.ends


* File: sky130_fd_sc_ms__and3b_2.pxi.spice
* Created: Wed Sep  2 11:58:03 2020
* 
x_PM_SKY130_FD_SC_MS__AND3B_2%A_N N_A_N_c_79_n N_A_N_c_84_n N_A_N_M1005_g
+ N_A_N_M1009_g A_N N_A_N_c_81_n N_A_N_c_82_n PM_SKY130_FD_SC_MS__AND3B_2%A_N
x_PM_SKY130_FD_SC_MS__AND3B_2%A_27_88# N_A_27_88#_M1009_s N_A_27_88#_M1005_s
+ N_A_27_88#_c_110_n N_A_27_88#_M1002_g N_A_27_88#_c_112_n N_A_27_88#_M1008_g
+ N_A_27_88#_c_113_n N_A_27_88#_c_114_n N_A_27_88#_c_115_n N_A_27_88#_c_116_n
+ N_A_27_88#_c_120_n N_A_27_88#_c_117_n N_A_27_88#_c_118_n N_A_27_88#_c_122_n
+ N_A_27_88#_c_123_n N_A_27_88#_c_124_n PM_SKY130_FD_SC_MS__AND3B_2%A_27_88#
x_PM_SKY130_FD_SC_MS__AND3B_2%B N_B_M1006_g N_B_M1001_g B B B B N_B_c_179_n
+ N_B_c_180_n PM_SKY130_FD_SC_MS__AND3B_2%B
x_PM_SKY130_FD_SC_MS__AND3B_2%C N_C_M1000_g N_C_M1003_g C N_C_c_219_n
+ PM_SKY130_FD_SC_MS__AND3B_2%C
x_PM_SKY130_FD_SC_MS__AND3B_2%A_284_368# N_A_284_368#_M1008_s
+ N_A_284_368#_M1002_s N_A_284_368#_M1001_d N_A_284_368#_M1004_g
+ N_A_284_368#_M1007_g N_A_284_368#_M1010_g N_A_284_368#_M1011_g
+ N_A_284_368#_c_259_n N_A_284_368#_c_266_n N_A_284_368#_c_281_n
+ N_A_284_368#_c_267_n N_A_284_368#_c_268_n N_A_284_368#_c_260_n
+ N_A_284_368#_c_270_n N_A_284_368#_c_285_n N_A_284_368#_c_261_n
+ N_A_284_368#_c_262_n PM_SKY130_FD_SC_MS__AND3B_2%A_284_368#
x_PM_SKY130_FD_SC_MS__AND3B_2%VPWR N_VPWR_M1005_d N_VPWR_M1002_d N_VPWR_M1003_d
+ N_VPWR_M1011_s N_VPWR_c_358_n N_VPWR_c_359_n N_VPWR_c_360_n N_VPWR_c_361_n
+ N_VPWR_c_362_n N_VPWR_c_363_n N_VPWR_c_364_n VPWR N_VPWR_c_365_n
+ N_VPWR_c_366_n N_VPWR_c_367_n N_VPWR_c_368_n N_VPWR_c_369_n N_VPWR_c_357_n
+ PM_SKY130_FD_SC_MS__AND3B_2%VPWR
x_PM_SKY130_FD_SC_MS__AND3B_2%X N_X_M1004_d N_X_M1007_d N_X_c_413_n X X X X X
+ PM_SKY130_FD_SC_MS__AND3B_2%X
x_PM_SKY130_FD_SC_MS__AND3B_2%VGND N_VGND_M1009_d N_VGND_M1000_d N_VGND_M1010_s
+ N_VGND_c_441_n N_VGND_c_442_n N_VGND_c_443_n N_VGND_c_444_n N_VGND_c_445_n
+ N_VGND_c_446_n VGND N_VGND_c_447_n N_VGND_c_448_n N_VGND_c_449_n
+ N_VGND_c_450_n PM_SKY130_FD_SC_MS__AND3B_2%VGND
cc_1 VNB N_A_N_c_79_n 0.0195074f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.755
cc_2 VNB N_A_N_M1009_g 0.0372275f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.715
cc_3 VNB N_A_N_c_81_n 0.0204063f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.425
cc_4 VNB N_A_N_c_82_n 0.0162384f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.425
cc_5 VNB N_A_27_88#_c_110_n 0.048996f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.715
cc_6 VNB N_A_27_88#_M1002_g 0.00300324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_88#_c_112_n 0.0196408f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.425
cc_8 VNB N_A_27_88#_c_113_n 0.0170325f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.595
cc_9 VNB N_A_27_88#_c_114_n 0.0211815f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.595
cc_10 VNB N_A_27_88#_c_115_n 0.0283998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_88#_c_116_n 0.00959922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_88#_c_117_n 0.00179898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_88#_c_118_n 0.0375386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B_M1001_g 0.00587774f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.26
cc_15 VNB B 0.00518004f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.715
cc_16 VNB N_B_c_179_n 0.0306834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B_c_180_n 0.0174585f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.595
cc_18 VNB N_C_M1000_g 0.0266942f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.02
cc_19 VNB C 0.00914442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_C_c_219_n 0.0226331f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.425
cc_21 VNB N_A_284_368#_M1004_g 0.0230215f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.425
cc_22 VNB N_A_284_368#_M1007_g 0.00145058f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.595
cc_23 VNB N_A_284_368#_M1010_g 0.0260225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_284_368#_M1011_g 0.00170504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_284_368#_c_259_n 0.0191617f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_284_368#_c_260_n 0.00121168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_284_368#_c_261_n 0.00753363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_284_368#_c_262_n 0.0846127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_357_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB X 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.425
cc_31 VNB X 0.00185591f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.425
cc_32 VNB N_VGND_c_441_n 0.0185992f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.425
cc_33 VNB N_VGND_c_442_n 0.00925448f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.595
cc_34 VNB N_VGND_c_443_n 0.0125919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_444_n 0.0419252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_445_n 0.0561173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_446_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_447_n 0.0177296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_448_n 0.0212406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_449_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_450_n 0.289569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VPB N_A_N_c_79_n 0.0385545f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.755
cc_43 VPB N_A_N_c_84_n 0.0264756f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.02
cc_44 VPB N_A_N_c_82_n 0.0112383f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.425
cc_45 VPB N_A_27_88#_M1002_g 0.027318f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_27_88#_c_120_n 0.0204899f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_27_88#_c_118_n 0.0249392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_27_88#_c_122_n 0.00515744f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_27_88#_c_123_n 0.0386655f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_27_88#_c_124_n 0.00647567f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_B_M1001_g 0.0230306f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.26
cc_52 VPB B 0.00305328f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.715
cc_53 VPB N_C_M1003_g 0.0210646f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.715
cc_54 VPB C 0.00671662f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_C_c_219_n 0.00545122f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.425
cc_56 VPB N_A_284_368#_M1007_g 0.0239413f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.595
cc_57 VPB N_A_284_368#_M1011_g 0.0248625f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_284_368#_c_259_n 0.00257159f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_284_368#_c_266_n 0.0180257f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_284_368#_c_267_n 0.0028233f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_284_368#_c_268_n 0.00769764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_284_368#_c_260_n 0.0218353f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_284_368#_c_270_n 0.00217379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_358_n 0.0202931f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=1.26
cc_65 VPB N_VPWR_c_359_n 0.0198884f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.595
cc_66 VPB N_VPWR_c_360_n 0.0102062f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_361_n 0.0119967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_362_n 0.0238914f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_363_n 0.0297343f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_364_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_365_n 0.017913f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_366_n 0.0211424f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_367_n 0.0182362f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_368_n 0.00613202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_369_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_357_n 0.0993241f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_X_c_413_n 3.60567e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB X 0.0011589f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.425
cc_79 N_A_N_M1009_g N_A_27_88#_c_114_n 0.00218986f $X=0.495 $Y=0.715 $X2=0 $Y2=0
cc_80 N_A_N_M1009_g N_A_27_88#_c_115_n 0.0180286f $X=0.495 $Y=0.715 $X2=0 $Y2=0
cc_81 N_A_N_c_81_n N_A_27_88#_c_115_n 0.00116829f $X=0.385 $Y=1.425 $X2=0 $Y2=0
cc_82 N_A_N_c_82_n N_A_27_88#_c_115_n 0.0133787f $X=0.385 $Y=1.425 $X2=0 $Y2=0
cc_83 N_A_N_c_81_n N_A_27_88#_c_116_n 0.00415347f $X=0.385 $Y=1.425 $X2=0 $Y2=0
cc_84 N_A_N_c_82_n N_A_27_88#_c_116_n 0.022566f $X=0.385 $Y=1.425 $X2=0 $Y2=0
cc_85 N_A_N_c_79_n N_A_27_88#_c_120_n 3.8731e-19 $X=0.395 $Y=1.755 $X2=0 $Y2=0
cc_86 N_A_N_c_84_n N_A_27_88#_c_120_n 0.0178226f $X=0.505 $Y=2.02 $X2=0 $Y2=0
cc_87 N_A_N_c_82_n N_A_27_88#_c_120_n 0.0113738f $X=0.385 $Y=1.425 $X2=0 $Y2=0
cc_88 N_A_N_M1009_g N_A_27_88#_c_117_n 0.00441126f $X=0.495 $Y=0.715 $X2=0 $Y2=0
cc_89 N_A_N_c_82_n N_A_27_88#_c_117_n 0.0287652f $X=0.385 $Y=1.425 $X2=0 $Y2=0
cc_90 N_A_N_M1009_g N_A_27_88#_c_118_n 0.0250202f $X=0.495 $Y=0.715 $X2=0 $Y2=0
cc_91 N_A_N_c_82_n N_A_27_88#_c_118_n 0.00256857f $X=0.385 $Y=1.425 $X2=0 $Y2=0
cc_92 N_A_N_c_79_n N_A_27_88#_c_122_n 0.00665196f $X=0.395 $Y=1.755 $X2=0 $Y2=0
cc_93 N_A_N_c_79_n N_A_27_88#_c_123_n 0.00483226f $X=0.395 $Y=1.755 $X2=0 $Y2=0
cc_94 N_A_N_c_84_n N_A_27_88#_c_123_n 0.00382138f $X=0.505 $Y=2.02 $X2=0 $Y2=0
cc_95 N_A_N_c_82_n N_A_27_88#_c_123_n 0.0248079f $X=0.385 $Y=1.425 $X2=0 $Y2=0
cc_96 N_A_N_c_81_n N_A_27_88#_c_124_n 0.00145659f $X=0.385 $Y=1.425 $X2=0 $Y2=0
cc_97 N_A_N_c_84_n N_VPWR_c_358_n 0.0175594f $X=0.505 $Y=2.02 $X2=0 $Y2=0
cc_98 N_A_N_c_84_n N_VPWR_c_365_n 0.00475445f $X=0.505 $Y=2.02 $X2=0 $Y2=0
cc_99 N_A_N_c_84_n N_VPWR_c_357_n 0.00942403f $X=0.505 $Y=2.02 $X2=0 $Y2=0
cc_100 N_A_N_M1009_g N_VGND_c_441_n 0.0117471f $X=0.495 $Y=0.715 $X2=0 $Y2=0
cc_101 N_A_N_M1009_g N_VGND_c_447_n 0.00438299f $X=0.495 $Y=0.715 $X2=0 $Y2=0
cc_102 N_A_N_M1009_g N_VGND_c_450_n 0.00439883f $X=0.495 $Y=0.715 $X2=0 $Y2=0
cc_103 N_A_27_88#_c_113_n N_B_M1001_g 0.0287775f $X=1.79 $Y=1.397 $X2=0 $Y2=0
cc_104 N_A_27_88#_c_112_n B 0.0107746f $X=1.805 $Y=1.185 $X2=0 $Y2=0
cc_105 N_A_27_88#_c_113_n N_B_c_179_n 0.0342483f $X=1.79 $Y=1.397 $X2=0 $Y2=0
cc_106 N_A_27_88#_c_112_n N_B_c_180_n 0.0342483f $X=1.805 $Y=1.185 $X2=0 $Y2=0
cc_107 N_A_27_88#_c_110_n N_A_284_368#_c_259_n 0.0305284f $X=1.7 $Y=1.397 $X2=0
+ $Y2=0
cc_108 N_A_27_88#_M1002_g N_A_284_368#_c_259_n 0.00978545f $X=1.79 $Y=2.34 $X2=0
+ $Y2=0
cc_109 N_A_27_88#_c_112_n N_A_284_368#_c_259_n 0.0144396f $X=1.805 $Y=1.185
+ $X2=0 $Y2=0
cc_110 N_A_27_88#_c_113_n N_A_284_368#_c_259_n 0.00742094f $X=1.79 $Y=1.397
+ $X2=0 $Y2=0
cc_111 N_A_27_88#_c_115_n N_A_284_368#_c_259_n 0.0151173f $X=0.9 $Y=1.005 $X2=0
+ $Y2=0
cc_112 N_A_27_88#_c_117_n N_A_284_368#_c_259_n 0.059451f $X=1.065 $Y=1.35 $X2=0
+ $Y2=0
cc_113 N_A_27_88#_c_118_n N_A_284_368#_c_259_n 0.00216806f $X=1.065 $Y=1.35
+ $X2=0 $Y2=0
cc_114 N_A_27_88#_c_122_n N_A_284_368#_c_259_n 0.00473672f $X=0.985 $Y=2.1 $X2=0
+ $Y2=0
cc_115 N_A_27_88#_M1002_g N_A_284_368#_c_266_n 0.0107668f $X=1.79 $Y=2.34 $X2=0
+ $Y2=0
cc_116 N_A_27_88#_c_120_n N_A_284_368#_c_266_n 0.0083406f $X=0.9 $Y=2.185 $X2=0
+ $Y2=0
cc_117 N_A_27_88#_M1002_g N_A_284_368#_c_281_n 0.0154646f $X=1.79 $Y=2.34 $X2=0
+ $Y2=0
cc_118 N_A_27_88#_M1002_g N_A_284_368#_c_270_n 0.0021104f $X=1.79 $Y=2.34 $X2=0
+ $Y2=0
cc_119 N_A_27_88#_c_120_n N_A_284_368#_c_270_n 0.00117914f $X=0.9 $Y=2.185 $X2=0
+ $Y2=0
cc_120 N_A_27_88#_c_122_n N_A_284_368#_c_270_n 0.00796471f $X=0.985 $Y=2.1 $X2=0
+ $Y2=0
cc_121 N_A_27_88#_M1002_g N_A_284_368#_c_285_n 7.11668e-19 $X=1.79 $Y=2.34 $X2=0
+ $Y2=0
cc_122 N_A_27_88#_c_120_n N_VPWR_M1005_d 0.00338403f $X=0.9 $Y=2.185 $X2=-0.19
+ $Y2=-0.245
cc_123 N_A_27_88#_c_120_n N_VPWR_c_358_n 0.0219251f $X=0.9 $Y=2.185 $X2=0 $Y2=0
cc_124 N_A_27_88#_c_123_n N_VPWR_c_358_n 0.0210352f $X=0.28 $Y=2.265 $X2=0 $Y2=0
cc_125 N_A_27_88#_M1002_g N_VPWR_c_359_n 0.00349882f $X=1.79 $Y=2.34 $X2=0 $Y2=0
cc_126 N_A_27_88#_M1002_g N_VPWR_c_363_n 0.00567889f $X=1.79 $Y=2.34 $X2=0 $Y2=0
cc_127 N_A_27_88#_c_123_n N_VPWR_c_365_n 0.0126277f $X=0.28 $Y=2.265 $X2=0 $Y2=0
cc_128 N_A_27_88#_M1002_g N_VPWR_c_357_n 0.00610055f $X=1.79 $Y=2.34 $X2=0 $Y2=0
cc_129 N_A_27_88#_c_123_n N_VPWR_c_357_n 0.0104521f $X=0.28 $Y=2.265 $X2=0 $Y2=0
cc_130 N_A_27_88#_c_115_n N_VGND_M1009_d 0.00296919f $X=0.9 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_131 N_A_27_88#_c_114_n N_VGND_c_441_n 0.0131449f $X=0.28 $Y=0.715 $X2=0 $Y2=0
cc_132 N_A_27_88#_c_115_n N_VGND_c_441_n 0.0219096f $X=0.9 $Y=1.005 $X2=0 $Y2=0
cc_133 N_A_27_88#_c_112_n N_VGND_c_445_n 0.00434272f $X=1.805 $Y=1.185 $X2=0
+ $Y2=0
cc_134 N_A_27_88#_c_114_n N_VGND_c_447_n 0.0089644f $X=0.28 $Y=0.715 $X2=0 $Y2=0
cc_135 N_A_27_88#_c_112_n N_VGND_c_450_n 0.00825979f $X=1.805 $Y=1.185 $X2=0
+ $Y2=0
cc_136 N_A_27_88#_c_114_n N_VGND_c_450_n 0.00911107f $X=0.28 $Y=0.715 $X2=0
+ $Y2=0
cc_137 B N_C_M1000_g 0.00907035f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_138 N_B_c_179_n N_C_M1000_g 0.012271f $X=2.285 $Y=1.385 $X2=0 $Y2=0
cc_139 N_B_c_180_n N_C_M1000_g 0.0240719f $X=2.285 $Y=1.22 $X2=0 $Y2=0
cc_140 N_B_M1001_g N_C_M1003_g 0.0135368f $X=2.36 $Y=2.34 $X2=0 $Y2=0
cc_141 N_B_M1001_g C 6.31308e-19 $X=2.36 $Y=2.34 $X2=0 $Y2=0
cc_142 B C 0.0262562f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_143 N_B_c_179_n C 0.00115663f $X=2.285 $Y=1.385 $X2=0 $Y2=0
cc_144 N_B_M1001_g N_C_c_219_n 0.012271f $X=2.36 $Y=2.34 $X2=0 $Y2=0
cc_145 B N_C_c_219_n 4.19042e-19 $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_146 N_B_M1001_g N_A_284_368#_c_259_n 9.88241e-19 $X=2.36 $Y=2.34 $X2=0 $Y2=0
cc_147 B N_A_284_368#_c_259_n 0.071653f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_148 N_B_c_180_n N_A_284_368#_c_259_n 0.00150231f $X=2.285 $Y=1.22 $X2=0 $Y2=0
cc_149 N_B_M1001_g N_A_284_368#_c_266_n 8.84754e-19 $X=2.36 $Y=2.34 $X2=0 $Y2=0
cc_150 N_B_M1001_g N_A_284_368#_c_281_n 0.0140859f $X=2.36 $Y=2.34 $X2=0 $Y2=0
cc_151 B N_A_284_368#_c_281_n 0.0279681f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_152 N_B_c_179_n N_A_284_368#_c_281_n 5.34801e-19 $X=2.285 $Y=1.385 $X2=0
+ $Y2=0
cc_153 N_B_M1001_g N_A_284_368#_c_267_n 0.00589514f $X=2.36 $Y=2.34 $X2=0 $Y2=0
cc_154 N_B_M1001_g N_A_284_368#_c_285_n 0.00636139f $X=2.36 $Y=2.34 $X2=0 $Y2=0
cc_155 B N_A_284_368#_c_285_n 0.00237022f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_156 N_B_M1001_g N_VPWR_c_359_n 0.00672099f $X=2.36 $Y=2.34 $X2=0 $Y2=0
cc_157 N_B_M1001_g N_VPWR_c_366_n 0.00567889f $X=2.36 $Y=2.34 $X2=0 $Y2=0
cc_158 N_B_M1001_g N_VPWR_c_357_n 0.00610055f $X=2.36 $Y=2.34 $X2=0 $Y2=0
cc_159 B N_VGND_c_442_n 0.030309f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_160 N_B_c_180_n N_VGND_c_442_n 0.0015178f $X=2.285 $Y=1.22 $X2=0 $Y2=0
cc_161 B N_VGND_c_445_n 0.0108342f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_162 N_B_c_180_n N_VGND_c_445_n 0.00303293f $X=2.285 $Y=1.22 $X2=0 $Y2=0
cc_163 B N_VGND_c_450_n 0.0133038f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_164 N_B_c_180_n N_VGND_c_450_n 0.00372643f $X=2.285 $Y=1.22 $X2=0 $Y2=0
cc_165 B A_376_74# 0.00738039f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_166 B A_454_74# 0.00983395f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_167 N_C_M1000_g N_A_284_368#_M1004_g 0.0181973f $X=2.765 $Y=0.74 $X2=0 $Y2=0
cc_168 N_C_M1003_g N_A_284_368#_M1007_g 0.0355577f $X=2.81 $Y=2.34 $X2=0 $Y2=0
cc_169 N_C_M1003_g N_A_284_368#_c_267_n 0.00747868f $X=2.81 $Y=2.34 $X2=0 $Y2=0
cc_170 N_C_M1003_g N_A_284_368#_c_268_n 0.0151438f $X=2.81 $Y=2.34 $X2=0 $Y2=0
cc_171 C N_A_284_368#_c_268_n 0.0164611f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_172 N_C_c_219_n N_A_284_368#_c_268_n 4.15225e-19 $X=2.855 $Y=1.515 $X2=0
+ $Y2=0
cc_173 N_C_M1003_g N_A_284_368#_c_285_n 0.00738163f $X=2.81 $Y=2.34 $X2=0 $Y2=0
cc_174 C N_A_284_368#_c_285_n 0.00362344f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_175 C N_A_284_368#_c_262_n 0.00403615f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_176 N_C_c_219_n N_A_284_368#_c_262_n 0.0178587f $X=2.855 $Y=1.515 $X2=0 $Y2=0
cc_177 N_C_M1003_g N_VPWR_c_360_n 0.00569686f $X=2.81 $Y=2.34 $X2=0 $Y2=0
cc_178 N_C_M1003_g N_VPWR_c_366_n 0.00567889f $X=2.81 $Y=2.34 $X2=0 $Y2=0
cc_179 N_C_M1003_g N_VPWR_c_357_n 0.00610055f $X=2.81 $Y=2.34 $X2=0 $Y2=0
cc_180 N_C_M1000_g X 2.59942e-19 $X=2.765 $Y=0.74 $X2=0 $Y2=0
cc_181 N_C_M1000_g X 2.16826e-19 $X=2.765 $Y=0.74 $X2=0 $Y2=0
cc_182 N_C_M1003_g X 0.0012194f $X=2.81 $Y=2.34 $X2=0 $Y2=0
cc_183 C X 0.034443f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_184 N_C_c_219_n X 2.31392e-19 $X=2.855 $Y=1.515 $X2=0 $Y2=0
cc_185 N_C_M1000_g N_VGND_c_442_n 0.0179953f $X=2.765 $Y=0.74 $X2=0 $Y2=0
cc_186 C N_VGND_c_442_n 0.0236581f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_187 N_C_c_219_n N_VGND_c_442_n 0.00430878f $X=2.855 $Y=1.515 $X2=0 $Y2=0
cc_188 N_C_M1000_g N_VGND_c_445_n 0.00383152f $X=2.765 $Y=0.74 $X2=0 $Y2=0
cc_189 N_C_M1000_g N_VGND_c_450_n 0.00758792f $X=2.765 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A_284_368#_c_281_n N_VPWR_M1002_d 0.00900736f $X=2.42 $Y=2.035 $X2=0
+ $Y2=0
cc_191 N_A_284_368#_c_268_n N_VPWR_M1003_d 0.00667869f $X=4.045 $Y=2.325 $X2=0
+ $Y2=0
cc_192 N_A_284_368#_c_268_n N_VPWR_M1011_s 0.00468907f $X=4.045 $Y=2.325 $X2=0
+ $Y2=0
cc_193 N_A_284_368#_c_260_n N_VPWR_M1011_s 0.00697509f $X=4.13 $Y=2.24 $X2=0
+ $Y2=0
cc_194 N_A_284_368#_c_266_n N_VPWR_c_358_n 0.0165803f $X=1.565 $Y=2.695 $X2=0
+ $Y2=0
cc_195 N_A_284_368#_c_266_n N_VPWR_c_359_n 0.0221782f $X=1.565 $Y=2.695 $X2=0
+ $Y2=0
cc_196 N_A_284_368#_c_281_n N_VPWR_c_359_n 0.022455f $X=2.42 $Y=2.035 $X2=0
+ $Y2=0
cc_197 N_A_284_368#_c_285_n N_VPWR_c_359_n 0.020261f $X=2.585 $Y=2.035 $X2=0
+ $Y2=0
cc_198 N_A_284_368#_M1007_g N_VPWR_c_360_n 0.0140648f $X=3.35 $Y=2.4 $X2=0 $Y2=0
cc_199 N_A_284_368#_M1011_g N_VPWR_c_360_n 0.0015105f $X=3.815 $Y=2.4 $X2=0
+ $Y2=0
cc_200 N_A_284_368#_c_267_n N_VPWR_c_360_n 0.018506f $X=2.585 $Y=2.715 $X2=0
+ $Y2=0
cc_201 N_A_284_368#_c_268_n N_VPWR_c_360_n 0.0218557f $X=4.045 $Y=2.325 $X2=0
+ $Y2=0
cc_202 N_A_284_368#_M1007_g N_VPWR_c_362_n 0.0015105f $X=3.35 $Y=2.4 $X2=0 $Y2=0
cc_203 N_A_284_368#_M1011_g N_VPWR_c_362_n 0.014544f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_204 N_A_284_368#_c_268_n N_VPWR_c_362_n 0.0232411f $X=4.045 $Y=2.325 $X2=0
+ $Y2=0
cc_205 N_A_284_368#_c_266_n N_VPWR_c_363_n 0.00975961f $X=1.565 $Y=2.695 $X2=0
+ $Y2=0
cc_206 N_A_284_368#_c_267_n N_VPWR_c_366_n 0.00967309f $X=2.585 $Y=2.715 $X2=0
+ $Y2=0
cc_207 N_A_284_368#_M1007_g N_VPWR_c_367_n 0.00460063f $X=3.35 $Y=2.4 $X2=0
+ $Y2=0
cc_208 N_A_284_368#_M1011_g N_VPWR_c_367_n 0.00460063f $X=3.815 $Y=2.4 $X2=0
+ $Y2=0
cc_209 N_A_284_368#_M1007_g N_VPWR_c_357_n 0.00908706f $X=3.35 $Y=2.4 $X2=0
+ $Y2=0
cc_210 N_A_284_368#_M1011_g N_VPWR_c_357_n 0.00908706f $X=3.815 $Y=2.4 $X2=0
+ $Y2=0
cc_211 N_A_284_368#_c_266_n N_VPWR_c_357_n 0.0111753f $X=1.565 $Y=2.695 $X2=0
+ $Y2=0
cc_212 N_A_284_368#_c_267_n N_VPWR_c_357_n 0.0111395f $X=2.585 $Y=2.715 $X2=0
+ $Y2=0
cc_213 N_A_284_368#_c_268_n N_X_M1007_d 0.00824948f $X=4.045 $Y=2.325 $X2=0
+ $Y2=0
cc_214 N_A_284_368#_M1007_g N_X_c_413_n 0.00582782f $X=3.35 $Y=2.4 $X2=0 $Y2=0
cc_215 N_A_284_368#_M1011_g N_X_c_413_n 0.00567836f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_216 N_A_284_368#_c_268_n N_X_c_413_n 0.0180796f $X=4.045 $Y=2.325 $X2=0 $Y2=0
cc_217 N_A_284_368#_c_260_n N_X_c_413_n 0.0123186f $X=4.13 $Y=2.24 $X2=0 $Y2=0
cc_218 N_A_284_368#_c_285_n N_X_c_413_n 0.00291109f $X=2.585 $Y=2.035 $X2=0
+ $Y2=0
cc_219 N_A_284_368#_M1004_g X 0.00855013f $X=3.335 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A_284_368#_M1010_g X 0.00788704f $X=3.765 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A_284_368#_M1004_g X 0.00345332f $X=3.335 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A_284_368#_M1010_g X 0.00202916f $X=3.765 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A_284_368#_M1004_g X 0.00483694f $X=3.335 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A_284_368#_M1007_g X 0.00440628f $X=3.35 $Y=2.4 $X2=0 $Y2=0
cc_225 N_A_284_368#_M1010_g X 0.00892301f $X=3.765 $Y=0.74 $X2=0 $Y2=0
cc_226 N_A_284_368#_M1011_g X 0.00211441f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_227 N_A_284_368#_c_260_n X 0.00937947f $X=4.13 $Y=2.24 $X2=0 $Y2=0
cc_228 N_A_284_368#_c_261_n X 0.0246163f $X=4.05 $Y=1.465 $X2=0 $Y2=0
cc_229 N_A_284_368#_c_262_n X 0.0221511f $X=4.05 $Y=1.465 $X2=0 $Y2=0
cc_230 N_A_284_368#_c_259_n N_VGND_c_441_n 0.0153399f $X=1.59 $Y=0.515 $X2=0
+ $Y2=0
cc_231 N_A_284_368#_M1004_g N_VGND_c_442_n 0.0100794f $X=3.335 $Y=0.74 $X2=0
+ $Y2=0
cc_232 N_A_284_368#_M1010_g N_VGND_c_444_n 0.00647412f $X=3.765 $Y=0.74 $X2=0
+ $Y2=0
cc_233 N_A_284_368#_c_261_n N_VGND_c_444_n 0.0214533f $X=4.05 $Y=1.465 $X2=0
+ $Y2=0
cc_234 N_A_284_368#_c_262_n N_VGND_c_444_n 0.001962f $X=4.05 $Y=1.465 $X2=0
+ $Y2=0
cc_235 N_A_284_368#_c_259_n N_VGND_c_445_n 0.0156794f $X=1.59 $Y=0.515 $X2=0
+ $Y2=0
cc_236 N_A_284_368#_M1004_g N_VGND_c_448_n 0.00434272f $X=3.335 $Y=0.74 $X2=0
+ $Y2=0
cc_237 N_A_284_368#_M1010_g N_VGND_c_448_n 0.00434272f $X=3.765 $Y=0.74 $X2=0
+ $Y2=0
cc_238 N_A_284_368#_M1004_g N_VGND_c_450_n 0.00822522f $X=3.335 $Y=0.74 $X2=0
+ $Y2=0
cc_239 N_A_284_368#_M1010_g N_VGND_c_450_n 0.0082413f $X=3.765 $Y=0.74 $X2=0
+ $Y2=0
cc_240 N_A_284_368#_c_259_n N_VGND_c_450_n 0.0129217f $X=1.59 $Y=0.515 $X2=0
+ $Y2=0
cc_241 X N_VGND_c_442_n 0.0465051f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_242 X N_VGND_c_444_n 0.0293763f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_243 X N_VGND_c_448_n 0.0144922f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_244 X N_VGND_c_450_n 0.0118826f $X=3.515 $Y=0.47 $X2=0 $Y2=0

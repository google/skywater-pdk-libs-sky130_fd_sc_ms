* File: sky130_fd_sc_ms__a21oi_1.pex.spice
* Created: Wed Sep  2 11:51:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A21OI_1%A2 3 5 7 8 15
c25 8 0 1.40395e-19 $X=0.24 $Y=1.295
r26 14 15 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.385
+ $X2=0.51 $Y2=1.385
r27 11 14 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.27 $Y=1.385
+ $X2=0.495 $Y2=1.385
r28 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r29 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.385
r30 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.22
+ $X2=0.51 $Y2=1.385
r31 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.51 $Y=1.22 $X2=0.51
+ $Y2=0.74
r32 1 14 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.55
+ $X2=0.495 $Y2=1.385
r33 1 3 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.495 $Y=1.55
+ $X2=0.495 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A21OI_1%A1 3 7 9 12 13
c37 12 0 3.37569e-19 $X=0.96 $Y=1.515
r38 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.515
+ $X2=0.96 $Y2=1.68
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.515
+ $X2=0.96 $Y2=1.35
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.96
+ $Y=1.515 $X2=0.96 $Y2=1.515
r41 9 13 6.43224 $w=4.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.96 $Y2=1.565
r42 7 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.975 $Y=2.4
+ $X2=0.975 $Y2=1.68
r43 3 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.87 $Y=0.74 $X2=0.87
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__A21OI_1%B1 1 3 6 8 14
r29 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.385 $X2=1.65 $Y2=1.385
r30 12 14 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=1.425 $Y=1.385
+ $X2=1.65 $Y2=1.385
r31 10 12 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.41 $Y=1.385
+ $X2=1.425 $Y2=1.385
r32 8 15 4.06745 $w=2.53e-07 $l=9e-08 $layer=LI1_cond $X=1.687 $Y=1.295
+ $X2=1.687 $Y2=1.385
r33 4 12 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.55
+ $X2=1.425 $Y2=1.385
r34 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.425 $Y=1.55
+ $X2=1.425 $Y2=2.4
r35 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.22
+ $X2=1.41 $Y2=1.385
r36 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.41 $Y=1.22 $X2=1.41
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A21OI_1%A_29_368# 1 2 7 9 11 18
c25 11 0 1.97174e-19 $X=0.833 $Y=2.107
r26 12 16 3.62238 $w=2.45e-07 $l=2.01879e-07 $layer=LI1_cond $X=0.435 $Y=2.107
+ $X2=0.27 $Y2=2.025
r27 11 18 18.9889 $w=2.45e-07 $l=3.67e-07 $layer=LI1_cond $X=0.833 $Y=2.107
+ $X2=1.2 $Y2=2.107
r28 11 12 18.7213 $w=2.43e-07 $l=3.98e-07 $layer=LI1_cond $X=0.833 $Y=2.107
+ $X2=0.435 $Y2=2.107
r29 7 16 3.2704 $w=2.95e-07 $l=2.13811e-07 $layer=LI1_cond $X=0.252 $Y=2.23
+ $X2=0.27 $Y2=2.025
r30 7 9 6.6412 $w=2.93e-07 $l=1.7e-07 $layer=LI1_cond $X=0.252 $Y=2.23 $X2=0.252
+ $Y2=2.4
r31 2 18 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=1.065
+ $Y=1.84 $X2=1.2 $Y2=2.225
r32 1 16 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=1.985
r33 1 9 300 $w=1.7e-07 $l=6.19354e-07 $layer=licon1_PDIFF $count=2 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A21OI_1%VPWR 1 6 8 10 17 18 21
r25 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r26 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r27 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.9 $Y=3.33
+ $X2=0.735 $Y2=3.33
r28 15 17 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=0.9 $Y=3.33 $X2=1.68
+ $Y2=3.33
r29 13 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r30 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r31 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.735 $Y2=3.33
r32 10 12 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 8 18 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r34 8 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r35 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=3.33
r36 4 6 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=2.485
r37 1 6 300 $w=1.7e-07 $l=7.16083e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=0.735 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_MS__A21OI_1%Y 1 2 9 12 13 14 16 18 19 20
r39 19 20 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.69 $Y=2.405
+ $X2=1.69 $Y2=2.775
r40 18 19 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=1.69 $Y=1.985
+ $X2=1.69 $Y2=2.405
r41 17 18 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=1.69 $Y=1.89
+ $X2=1.69 $Y2=1.985
r42 15 16 8.69455 $w=3.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.155 $Y=1.01
+ $X2=1.155 $Y2=1.18
r43 13 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.565 $Y=1.805
+ $X2=1.69 $Y2=1.89
r44 13 14 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.565 $Y=1.805
+ $X2=1.39 $Y2=1.805
r45 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.305 $Y=1.72
+ $X2=1.39 $Y2=1.805
r46 12 16 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=1.305 $Y=1.72
+ $X2=1.305 $Y2=1.18
r47 9 15 15.4178 $w=3.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.105 $Y=0.515
+ $X2=1.105 $Y2=1.01
r48 2 20 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.515
+ $Y=1.84 $X2=1.65 $Y2=2.815
r49 2 18 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.515
+ $Y=1.84 $X2=1.65 $Y2=1.985
r50 1 9 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=0.945
+ $Y=0.37 $X2=1.105 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A21OI_1%VGND 1 2 7 9 11 13 15 17 27
r24 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r25 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r26 21 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r27 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r28 18 23 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.46 $Y=0 $X2=0.23
+ $Y2=0
r29 18 20 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.46 $Y=0 $X2=1.2
+ $Y2=0
r30 17 26 3.82794 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.74
+ $Y2=0
r31 17 20 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.2
+ $Y2=0
r32 15 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r33 15 24 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.24
+ $Y2=0
r34 11 26 3.18995 $w=2.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=1.675 $Y=0.085
+ $X2=1.74 $Y2=0
r35 11 13 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.675 $Y=0.085
+ $X2=1.675 $Y2=0.515
r36 7 23 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.295 $Y=0.085
+ $X2=0.23 $Y2=0
r37 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.295 $Y=0.085
+ $X2=0.295 $Y2=0.515
r38 2 13 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=1.485
+ $Y=0.37 $X2=1.645 $Y2=0.515
r39 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.17
+ $Y=0.37 $X2=0.295 $Y2=0.515
.ends


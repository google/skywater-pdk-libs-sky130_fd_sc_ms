* File: sky130_fd_sc_ms__nor2_8.pxi.spice
* Created: Fri Aug 28 17:47:10 2020
* 
x_PM_SKY130_FD_SC_MS__NOR2_8%A N_A_c_134_n N_A_M1001_g N_A_c_122_n N_A_c_123_n
+ N_A_c_137_n N_A_M1003_g N_A_c_124_n N_A_c_139_n N_A_M1004_g N_A_c_125_n
+ N_A_M1002_g N_A_c_141_n N_A_M1006_g N_A_M1005_g N_A_c_142_n N_A_M1007_g
+ N_A_c_143_n N_A_M1010_g N_A_M1014_g N_A_c_144_n N_A_M1011_g N_A_M1016_g
+ N_A_c_145_n N_A_M1015_g N_A_c_130_n N_A_c_131_n A A A A A N_A_c_133_n
+ PM_SKY130_FD_SC_MS__NOR2_8%A
x_PM_SKY130_FD_SC_MS__NOR2_8%B N_B_c_251_n N_B_M1000_g N_B_M1012_g N_B_c_253_n
+ N_B_M1013_g N_B_c_255_n N_B_M1017_g N_B_c_257_n N_B_M1008_g N_B_c_258_n
+ N_B_M1018_g N_B_c_260_n N_B_M1009_g N_B_M1019_g N_B_c_262_n N_B_M1023_g
+ N_B_c_263_n N_B_c_264_n N_B_M1020_g N_B_c_266_n N_B_M1021_g N_B_M1022_g
+ N_B_c_269_n N_B_c_270_n N_B_c_271_n N_B_c_272_n N_B_c_273_n B B N_B_c_274_n
+ N_B_c_275_n PM_SKY130_FD_SC_MS__NOR2_8%B
x_PM_SKY130_FD_SC_MS__NOR2_8%A_27_368# N_A_27_368#_M1001_d N_A_27_368#_M1003_d
+ N_A_27_368#_M1006_d N_A_27_368#_M1010_d N_A_27_368#_M1015_d
+ N_A_27_368#_M1013_s N_A_27_368#_M1018_s N_A_27_368#_M1020_s
+ N_A_27_368#_M1022_s N_A_27_368#_c_385_n N_A_27_368#_c_386_n
+ N_A_27_368#_c_387_n N_A_27_368#_c_388_n N_A_27_368#_c_409_n
+ N_A_27_368#_c_389_n N_A_27_368#_c_415_n N_A_27_368#_c_390_n
+ N_A_27_368#_c_421_n N_A_27_368#_c_425_n N_A_27_368#_c_426_n
+ N_A_27_368#_c_391_n N_A_27_368#_c_392_n N_A_27_368#_c_444_n
+ N_A_27_368#_c_393_n N_A_27_368#_c_394_n N_A_27_368#_c_395_n
+ N_A_27_368#_c_396_n N_A_27_368#_c_397_n N_A_27_368#_c_398_n
+ N_A_27_368#_c_399_n N_A_27_368#_c_431_n N_A_27_368#_c_434_n
+ N_A_27_368#_c_400_n N_A_27_368#_c_401_n N_A_27_368#_c_402_n
+ PM_SKY130_FD_SC_MS__NOR2_8%A_27_368#
x_PM_SKY130_FD_SC_MS__NOR2_8%VPWR N_VPWR_M1001_s N_VPWR_M1004_s N_VPWR_M1007_s
+ N_VPWR_M1011_s N_VPWR_c_516_n N_VPWR_c_517_n N_VPWR_c_518_n N_VPWR_c_519_n
+ VPWR N_VPWR_c_520_n N_VPWR_c_521_n N_VPWR_c_522_n N_VPWR_c_523_n
+ N_VPWR_c_524_n N_VPWR_c_515_n N_VPWR_c_526_n N_VPWR_c_527_n N_VPWR_c_528_n
+ N_VPWR_c_529_n PM_SKY130_FD_SC_MS__NOR2_8%VPWR
x_PM_SKY130_FD_SC_MS__NOR2_8%Y N_Y_M1002_s N_Y_M1014_s N_Y_M1000_s N_Y_M1009_s
+ N_Y_M1012_d N_Y_M1017_d N_Y_M1019_d N_Y_M1021_d N_Y_c_614_n N_Y_c_615_n
+ N_Y_c_616_n N_Y_c_617_n N_Y_c_618_n N_Y_c_623_n N_Y_c_647_n N_Y_c_619_n
+ N_Y_c_654_n N_Y_c_620_n N_Y_c_621_n N_Y_c_681_n N_Y_c_622_n Y Y
+ PM_SKY130_FD_SC_MS__NOR2_8%Y
x_PM_SKY130_FD_SC_MS__NOR2_8%VGND N_VGND_M1002_d N_VGND_M1005_d N_VGND_M1016_d
+ N_VGND_M1008_d N_VGND_M1023_d N_VGND_c_723_n N_VGND_c_724_n N_VGND_c_725_n
+ N_VGND_c_726_n N_VGND_c_727_n N_VGND_c_728_n N_VGND_c_729_n VGND
+ N_VGND_c_730_n N_VGND_c_731_n N_VGND_c_732_n N_VGND_c_733_n N_VGND_c_734_n
+ N_VGND_c_735_n N_VGND_c_736_n N_VGND_c_737_n N_VGND_c_738_n
+ PM_SKY130_FD_SC_MS__NOR2_8%VGND
cc_1 VNB N_A_c_122_n 0.0136212f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.65
cc_2 VNB N_A_c_123_n 0.0162708f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.65
cc_3 VNB N_A_c_124_n 0.0105251f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=1.65
cc_4 VNB N_A_c_125_n 0.00713292f $X=-0.19 $Y=-0.245 $X2=1.735 $Y2=1.65
cc_5 VNB N_A_M1002_g 0.0315514f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=0.74
cc_6 VNB N_A_M1005_g 0.0315587f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=0.74
cc_7 VNB N_A_M1014_g 0.0307539f $X=-0.19 $Y=-0.245 $X2=3.21 $Y2=0.74
cc_8 VNB N_A_M1016_g 0.0247574f $X=-0.19 $Y=-0.245 $X2=3.71 $Y2=0.74
cc_9 VNB N_A_c_130_n 0.00735408f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.65
cc_10 VNB N_A_c_131_n 0.00735408f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=1.65
cc_11 VNB A 0.012161f $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=1.58
cc_12 VNB N_A_c_133_n 0.110949f $X=-0.19 $Y=-0.245 $X2=3.71 $Y2=1.537
cc_13 VNB N_B_c_251_n 0.0200058f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.725
cc_14 VNB N_B_M1012_g 0.0196625f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.725
cc_15 VNB N_B_c_253_n 0.0181613f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_16 VNB N_B_M1013_g 0.0158298f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=2.4
cc_17 VNB N_B_c_255_n 0.0166202f $X=-0.19 $Y=-0.245 $X2=1.735 $Y2=1.65
cc_18 VNB N_B_M1017_g 0.015177f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=0.74
cc_19 VNB N_B_c_257_n 0.020416f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.725
cc_20 VNB N_B_c_258_n 0.0117381f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=1.35
cc_21 VNB N_B_M1018_g 0.0145655f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=1.725
cc_22 VNB N_B_c_260_n 0.0157738f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=2.4
cc_23 VNB N_B_M1019_g 0.015156f $X=-0.19 $Y=-0.245 $X2=3.21 $Y2=0.74
cc_24 VNB N_B_c_262_n 0.0169231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B_c_263_n 0.00635223f $X=-0.19 $Y=-0.245 $X2=3.305 $Y2=2.4
cc_26 VNB N_B_c_264_n 0.0193653f $X=-0.19 $Y=-0.245 $X2=3.71 $Y2=1.35
cc_27 VNB N_B_M1020_g 0.0163843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B_c_266_n 0.0188047f $X=-0.19 $Y=-0.245 $X2=3.855 $Y2=2.4
cc_29 VNB N_B_M1021_g 0.0164034f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_30 VNB N_B_M1022_g 0.0264902f $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=1.58
cc_31 VNB N_B_c_269_n 0.0109817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_B_c_270_n 0.00800249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_B_c_271_n 0.00294508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_B_c_272_n 0.0073596f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=1.515
cc_35 VNB N_B_c_273_n 0.0206427f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=1.537
cc_36 VNB N_B_c_274_n 0.150322f $X=-0.19 $Y=-0.245 $X2=3.42 $Y2=1.515
cc_37 VNB N_B_c_275_n 0.00258269f $X=-0.19 $Y=-0.245 $X2=3.71 $Y2=1.537
cc_38 VNB N_VPWR_c_515_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_Y_c_614_n 0.00280455f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=1.725
cc_40 VNB N_Y_c_615_n 0.00636217f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=2.4
cc_41 VNB N_Y_c_616_n 0.00231148f $X=-0.19 $Y=-0.245 $X2=2.855 $Y2=1.725
cc_42 VNB N_Y_c_617_n 0.00280455f $X=-0.19 $Y=-0.245 $X2=3.21 $Y2=1.35
cc_43 VNB N_Y_c_618_n 0.00879444f $X=-0.19 $Y=-0.245 $X2=3.21 $Y2=0.74
cc_44 VNB N_Y_c_619_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.58
cc_45 VNB N_Y_c_620_n 0.0135921f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.537
cc_46 VNB N_Y_c_621_n 0.0298908f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.537
cc_47 VNB N_Y_c_622_n 0.00231148f $X=-0.19 $Y=-0.245 $X2=3.21 $Y2=1.537
cc_48 VNB N_VGND_c_723_n 0.065313f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.725
cc_49 VNB N_VGND_c_724_n 0.00936836f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=0.74
cc_50 VNB N_VGND_c_725_n 0.00585698f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=2.4
cc_51 VNB N_VGND_c_726_n 0.0351261f $X=-0.19 $Y=-0.245 $X2=2.855 $Y2=2.4
cc_52 VNB N_VGND_c_727_n 0.00899973f $X=-0.19 $Y=-0.245 $X2=3.21 $Y2=0.74
cc_53 VNB N_VGND_c_728_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=3.305 $Y2=1.725
cc_54 VNB N_VGND_c_729_n 0.0211799f $X=-0.19 $Y=-0.245 $X2=3.71 $Y2=0.74
cc_55 VNB N_VGND_c_730_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=3.855 $Y2=2.4
cc_56 VNB N_VGND_c_731_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_57 VNB N_VGND_c_732_n 0.0433909f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.537
cc_58 VNB N_VGND_c_733_n 0.474712f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=1.537
cc_59 VNB N_VGND_c_734_n 0.0428317f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=1.537
cc_60 VNB N_VGND_c_735_n 0.0138518f $X=-0.19 $Y=-0.245 $X2=3.42 $Y2=1.537
cc_61 VNB N_VGND_c_736_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=3.71 $Y2=1.537
cc_62 VNB N_VGND_c_737_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_738_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.565
cc_64 VPB N_A_c_134_n 0.0251108f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.725
cc_65 VPB N_A_c_122_n 0.00517211f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=1.65
cc_66 VPB N_A_c_123_n 0.00483437f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.65
cc_67 VPB N_A_c_137_n 0.0182323f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.725
cc_68 VPB N_A_c_124_n 0.00376305f $X=-0.19 $Y=1.66 $X2=1.365 $Y2=1.65
cc_69 VPB N_A_c_139_n 0.0182691f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.725
cc_70 VPB N_A_c_125_n 0.00387443f $X=-0.19 $Y=1.66 $X2=1.735 $Y2=1.65
cc_71 VPB N_A_c_141_n 0.0178412f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.725
cc_72 VPB N_A_c_142_n 0.0189558f $X=-0.19 $Y=1.66 $X2=2.355 $Y2=1.725
cc_73 VPB N_A_c_143_n 0.0183678f $X=-0.19 $Y=1.66 $X2=2.855 $Y2=1.725
cc_74 VPB N_A_c_144_n 0.0193923f $X=-0.19 $Y=1.66 $X2=3.305 $Y2=1.725
cc_75 VPB N_A_c_145_n 0.019655f $X=-0.19 $Y=1.66 $X2=3.855 $Y2=1.725
cc_76 VPB N_A_c_130_n 0.00124171f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.65
cc_77 VPB N_A_c_131_n 0.00124171f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=1.65
cc_78 VPB A 0.014499f $X=-0.19 $Y=1.66 $X2=3.515 $Y2=1.58
cc_79 VPB N_A_c_133_n 0.0310853f $X=-0.19 $Y=1.66 $X2=3.71 $Y2=1.537
cc_80 VPB N_B_M1012_g 0.0224743f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.725
cc_81 VPB N_B_M1013_g 0.0215292f $X=-0.19 $Y=1.66 $X2=1.455 $Y2=2.4
cc_82 VPB N_B_M1017_g 0.0209105f $X=-0.19 $Y=1.66 $X2=1.81 $Y2=0.74
cc_83 VPB N_B_M1018_g 0.0207781f $X=-0.19 $Y=1.66 $X2=2.355 $Y2=1.725
cc_84 VPB N_B_M1019_g 0.020791f $X=-0.19 $Y=1.66 $X2=3.21 $Y2=0.74
cc_85 VPB N_B_M1020_g 0.0214124f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_B_M1021_g 0.0214124f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_87 VPB N_B_M1022_g 0.0280697f $X=-0.19 $Y=1.66 $X2=3.515 $Y2=1.58
cc_88 VPB N_A_27_368#_c_385_n 0.0417114f $X=-0.19 $Y=1.66 $X2=2.855 $Y2=1.725
cc_89 VPB N_A_27_368#_c_386_n 0.006229f $X=-0.19 $Y=1.66 $X2=3.21 $Y2=0.74
cc_90 VPB N_A_27_368#_c_387_n 0.0194896f $X=-0.19 $Y=1.66 $X2=3.21 $Y2=0.74
cc_91 VPB N_A_27_368#_c_388_n 0.00179594f $X=-0.19 $Y=1.66 $X2=3.305 $Y2=2.4
cc_92 VPB N_A_27_368#_c_389_n 0.00202354f $X=-0.19 $Y=1.66 $X2=3.855 $Y2=1.725
cc_93 VPB N_A_27_368#_c_390_n 0.00202354f $X=-0.19 $Y=1.66 $X2=2.075 $Y2=1.58
cc_94 VPB N_A_27_368#_c_391_n 0.00248492f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_27_368#_c_392_n 0.00196551f $X=-0.19 $Y=1.66 $X2=1.81 $Y2=1.537
cc_96 VPB N_A_27_368#_c_393_n 0.00233539f $X=-0.19 $Y=1.66 $X2=2.855 $Y2=1.537
cc_97 VPB N_A_27_368#_c_394_n 0.00201002f $X=-0.19 $Y=1.66 $X2=3.42 $Y2=1.515
cc_98 VPB N_A_27_368#_c_395_n 0.00237099f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.565
cc_99 VPB N_A_27_368#_c_396_n 0.0024533f $X=-0.19 $Y=1.66 $X2=2.16 $Y2=1.565
cc_100 VPB N_A_27_368#_c_397_n 0.0123539f $X=-0.19 $Y=1.66 $X2=3.12 $Y2=1.565
cc_101 VPB N_A_27_368#_c_398_n 0.0548516f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_27_368#_c_399_n 0.00284703f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_27_368#_c_400_n 0.00189272f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_27_368#_c_401_n 0.00149233f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_27_368#_c_402_n 0.00189272f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_516_n 0.00568435f $X=-0.19 $Y=1.66 $X2=1.545 $Y2=1.65
cc_107 VPB N_VPWR_c_517_n 0.0026822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_518_n 0.0049562f $X=-0.19 $Y=1.66 $X2=2.31 $Y2=1.35
cc_109 VPB N_VPWR_c_519_n 0.0084909f $X=-0.19 $Y=1.66 $X2=2.355 $Y2=1.725
cc_110 VPB N_VPWR_c_520_n 0.0191515f $X=-0.19 $Y=1.66 $X2=2.855 $Y2=2.4
cc_111 VPB N_VPWR_c_521_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_522_n 0.0175706f $X=-0.19 $Y=1.66 $X2=3.71 $Y2=0.74
cc_113 VPB N_VPWR_c_523_n 0.0175706f $X=-0.19 $Y=1.66 $X2=3.855 $Y2=2.4
cc_114 VPB N_VPWR_c_524_n 0.102584f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_515_n 0.0833148f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_526_n 0.0061274f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.537
cc_117 VPB N_VPWR_c_527_n 0.00601644f $X=-0.19 $Y=1.66 $X2=2.06 $Y2=1.515
cc_118 VPB N_VPWR_c_528_n 0.0061274f $X=-0.19 $Y=1.66 $X2=2.855 $Y2=1.537
cc_119 VPB N_VPWR_c_529_n 0.00631788f $X=-0.19 $Y=1.66 $X2=3.42 $Y2=1.537
cc_120 VPB N_Y_c_623_n 8.06968e-19 $X=-0.19 $Y=1.66 $X2=3.305 $Y2=2.4
cc_121 VPB N_Y_c_621_n 0.00675591f $X=-0.19 $Y=1.66 $X2=1.905 $Y2=1.537
cc_122 N_A_M1016_g N_B_c_251_n 0.0286926f $X=3.71 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_123 N_A_M1016_g N_B_M1012_g 0.00677313f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_124 A N_B_M1012_g 0.001746f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_125 N_A_c_133_n N_B_M1012_g 0.0196342f $X=3.71 $Y=1.537 $X2=0 $Y2=0
cc_126 N_A_c_134_n N_A_27_368#_c_385_n 0.0147224f $X=0.505 $Y=1.725 $X2=0 $Y2=0
cc_127 N_A_c_137_n N_A_27_368#_c_385_n 9.98799e-19 $X=1.005 $Y=1.725 $X2=0 $Y2=0
cc_128 N_A_c_134_n N_A_27_368#_c_386_n 0.0169566f $X=0.505 $Y=1.725 $X2=0 $Y2=0
cc_129 N_A_c_122_n N_A_27_368#_c_386_n 0.00388793f $X=0.915 $Y=1.65 $X2=0 $Y2=0
cc_130 N_A_c_137_n N_A_27_368#_c_386_n 0.0162266f $X=1.005 $Y=1.725 $X2=0 $Y2=0
cc_131 N_A_c_134_n N_A_27_368#_c_387_n 0.00303312f $X=0.505 $Y=1.725 $X2=0 $Y2=0
cc_132 N_A_c_139_n N_A_27_368#_c_409_n 0.0191004f $X=1.455 $Y=1.725 $X2=0 $Y2=0
cc_133 N_A_c_125_n N_A_27_368#_c_409_n 5.54179e-19 $X=1.735 $Y=1.65 $X2=0 $Y2=0
cc_134 N_A_c_141_n N_A_27_368#_c_409_n 0.0142175f $X=1.905 $Y=1.725 $X2=0 $Y2=0
cc_135 A N_A_27_368#_c_409_n 0.0317652f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_136 N_A_c_142_n N_A_27_368#_c_389_n 0.0115755f $X=2.355 $Y=1.725 $X2=0 $Y2=0
cc_137 N_A_c_143_n N_A_27_368#_c_389_n 9.01797e-19 $X=2.855 $Y=1.725 $X2=0 $Y2=0
cc_138 N_A_c_142_n N_A_27_368#_c_415_n 0.0132272f $X=2.355 $Y=1.725 $X2=0 $Y2=0
cc_139 N_A_c_143_n N_A_27_368#_c_415_n 0.0145524f $X=2.855 $Y=1.725 $X2=0 $Y2=0
cc_140 A N_A_27_368#_c_415_n 0.047525f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_141 N_A_c_133_n N_A_27_368#_c_415_n 8.48758e-19 $X=3.71 $Y=1.537 $X2=0 $Y2=0
cc_142 N_A_c_144_n N_A_27_368#_c_390_n 0.0119537f $X=3.305 $Y=1.725 $X2=0 $Y2=0
cc_143 N_A_c_145_n N_A_27_368#_c_390_n 6.01945e-19 $X=3.855 $Y=1.725 $X2=0 $Y2=0
cc_144 N_A_c_144_n N_A_27_368#_c_421_n 0.0134861f $X=3.305 $Y=1.725 $X2=0 $Y2=0
cc_145 N_A_c_145_n N_A_27_368#_c_421_n 0.017588f $X=3.855 $Y=1.725 $X2=0 $Y2=0
cc_146 A N_A_27_368#_c_421_n 0.0340746f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_147 N_A_c_133_n N_A_27_368#_c_421_n 0.00114327f $X=3.71 $Y=1.537 $X2=0 $Y2=0
cc_148 N_A_c_145_n N_A_27_368#_c_425_n 0.00184802f $X=3.855 $Y=1.725 $X2=0 $Y2=0
cc_149 N_A_c_144_n N_A_27_368#_c_426_n 5.84028e-19 $X=3.305 $Y=1.725 $X2=0 $Y2=0
cc_150 N_A_c_145_n N_A_27_368#_c_426_n 0.0106645f $X=3.855 $Y=1.725 $X2=0 $Y2=0
cc_151 N_A_c_145_n N_A_27_368#_c_392_n 0.00338824f $X=3.855 $Y=1.725 $X2=0 $Y2=0
cc_152 N_A_c_124_n N_A_27_368#_c_399_n 0.00280743f $X=1.365 $Y=1.65 $X2=0 $Y2=0
cc_153 N_A_c_139_n N_A_27_368#_c_399_n 0.00142373f $X=1.455 $Y=1.725 $X2=0 $Y2=0
cc_154 N_A_c_142_n N_A_27_368#_c_431_n 8.84614e-19 $X=2.355 $Y=1.725 $X2=0 $Y2=0
cc_155 A N_A_27_368#_c_431_n 0.0189743f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_156 N_A_c_133_n N_A_27_368#_c_431_n 6.13576e-19 $X=3.71 $Y=1.537 $X2=0 $Y2=0
cc_157 N_A_c_144_n N_A_27_368#_c_434_n 8.84614e-19 $X=3.305 $Y=1.725 $X2=0 $Y2=0
cc_158 A N_A_27_368#_c_434_n 0.0189743f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_159 N_A_c_133_n N_A_27_368#_c_434_n 6.10251e-19 $X=3.71 $Y=1.537 $X2=0 $Y2=0
cc_160 N_A_c_134_n N_VPWR_c_516_n 0.00408927f $X=0.505 $Y=1.725 $X2=0 $Y2=0
cc_161 N_A_c_137_n N_VPWR_c_516_n 0.0163605f $X=1.005 $Y=1.725 $X2=0 $Y2=0
cc_162 N_A_c_139_n N_VPWR_c_516_n 5.9496e-19 $X=1.455 $Y=1.725 $X2=0 $Y2=0
cc_163 N_A_c_137_n N_VPWR_c_517_n 5.41206e-19 $X=1.005 $Y=1.725 $X2=0 $Y2=0
cc_164 N_A_c_139_n N_VPWR_c_517_n 0.0127835f $X=1.455 $Y=1.725 $X2=0 $Y2=0
cc_165 N_A_c_141_n N_VPWR_c_517_n 0.0128656f $X=1.905 $Y=1.725 $X2=0 $Y2=0
cc_166 N_A_c_142_n N_VPWR_c_517_n 5.56271e-19 $X=2.355 $Y=1.725 $X2=0 $Y2=0
cc_167 N_A_c_142_n N_VPWR_c_518_n 0.00188411f $X=2.355 $Y=1.725 $X2=0 $Y2=0
cc_168 N_A_c_143_n N_VPWR_c_518_n 0.0128297f $X=2.855 $Y=1.725 $X2=0 $Y2=0
cc_169 N_A_c_144_n N_VPWR_c_518_n 5.56271e-19 $X=3.305 $Y=1.725 $X2=0 $Y2=0
cc_170 N_A_c_144_n N_VPWR_c_519_n 0.00197411f $X=3.305 $Y=1.725 $X2=0 $Y2=0
cc_171 N_A_c_145_n N_VPWR_c_519_n 0.00150551f $X=3.855 $Y=1.725 $X2=0 $Y2=0
cc_172 N_A_c_134_n N_VPWR_c_520_n 0.005209f $X=0.505 $Y=1.725 $X2=0 $Y2=0
cc_173 N_A_c_137_n N_VPWR_c_521_n 0.00460063f $X=1.005 $Y=1.725 $X2=0 $Y2=0
cc_174 N_A_c_139_n N_VPWR_c_521_n 0.00460063f $X=1.455 $Y=1.725 $X2=0 $Y2=0
cc_175 N_A_c_141_n N_VPWR_c_522_n 0.00460063f $X=1.905 $Y=1.725 $X2=0 $Y2=0
cc_176 N_A_c_142_n N_VPWR_c_522_n 0.005209f $X=2.355 $Y=1.725 $X2=0 $Y2=0
cc_177 N_A_c_143_n N_VPWR_c_523_n 0.00460063f $X=2.855 $Y=1.725 $X2=0 $Y2=0
cc_178 N_A_c_144_n N_VPWR_c_523_n 0.005209f $X=3.305 $Y=1.725 $X2=0 $Y2=0
cc_179 N_A_c_145_n N_VPWR_c_524_n 0.00517089f $X=3.855 $Y=1.725 $X2=0 $Y2=0
cc_180 N_A_c_134_n N_VPWR_c_515_n 0.00985824f $X=0.505 $Y=1.725 $X2=0 $Y2=0
cc_181 N_A_c_137_n N_VPWR_c_515_n 0.00908554f $X=1.005 $Y=1.725 $X2=0 $Y2=0
cc_182 N_A_c_139_n N_VPWR_c_515_n 0.00908554f $X=1.455 $Y=1.725 $X2=0 $Y2=0
cc_183 N_A_c_141_n N_VPWR_c_515_n 0.00908554f $X=1.905 $Y=1.725 $X2=0 $Y2=0
cc_184 N_A_c_142_n N_VPWR_c_515_n 0.00982082f $X=2.355 $Y=1.725 $X2=0 $Y2=0
cc_185 N_A_c_143_n N_VPWR_c_515_n 0.00908554f $X=2.855 $Y=1.725 $X2=0 $Y2=0
cc_186 N_A_c_144_n N_VPWR_c_515_n 0.00982526f $X=3.305 $Y=1.725 $X2=0 $Y2=0
cc_187 N_A_c_145_n N_VPWR_c_515_n 0.00977848f $X=3.855 $Y=1.725 $X2=0 $Y2=0
cc_188 N_A_M1002_g N_Y_c_614_n 0.00821243f $X=1.81 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A_M1005_g N_Y_c_614_n 0.00350341f $X=2.31 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A_M1005_g N_Y_c_615_n 0.0167736f $X=2.31 $Y=0.74 $X2=0 $Y2=0
cc_191 N_A_M1014_g N_Y_c_615_n 0.0131906f $X=3.21 $Y=0.74 $X2=0 $Y2=0
cc_192 A N_Y_c_615_n 0.0809793f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_193 N_A_c_133_n N_Y_c_615_n 0.0145243f $X=3.71 $Y=1.537 $X2=0 $Y2=0
cc_194 N_A_M1002_g N_Y_c_616_n 0.00499186f $X=1.81 $Y=0.74 $X2=0 $Y2=0
cc_195 A N_Y_c_616_n 0.0282341f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_196 N_A_c_133_n N_Y_c_616_n 0.00443007f $X=3.71 $Y=1.537 $X2=0 $Y2=0
cc_197 N_A_M1014_g N_Y_c_617_n 0.0137366f $X=3.21 $Y=0.74 $X2=0 $Y2=0
cc_198 N_A_M1016_g N_Y_c_617_n 0.00350341f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A_M1016_g N_Y_c_618_n 0.0172035f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_200 A N_Y_c_618_n 0.00925196f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_201 N_A_c_133_n N_Y_c_618_n 0.0052328f $X=3.71 $Y=1.537 $X2=0 $Y2=0
cc_202 N_A_M1016_g N_Y_c_621_n 0.00133266f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A_M1014_g N_Y_c_622_n 0.00173883f $X=3.21 $Y=0.74 $X2=0 $Y2=0
cc_204 A N_Y_c_622_n 0.0282341f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_205 N_A_c_133_n N_Y_c_622_n 0.00443007f $X=3.71 $Y=1.537 $X2=0 $Y2=0
cc_206 N_A_c_122_n N_VGND_c_723_n 0.0237644f $X=0.915 $Y=1.65 $X2=0 $Y2=0
cc_207 N_A_c_125_n N_VGND_c_723_n 5.99493e-19 $X=1.735 $Y=1.65 $X2=0 $Y2=0
cc_208 N_A_M1002_g N_VGND_c_723_n 0.00556557f $X=1.81 $Y=0.74 $X2=0 $Y2=0
cc_209 A N_VGND_c_723_n 0.00932589f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_210 N_A_M1002_g N_VGND_c_724_n 4.95933e-19 $X=1.81 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A_M1005_g N_VGND_c_724_n 0.0137423f $X=2.31 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A_M1014_g N_VGND_c_724_n 0.00607183f $X=3.21 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A_M1014_g N_VGND_c_725_n 4.99121e-19 $X=3.21 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A_M1016_g N_VGND_c_725_n 0.0109084f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A_M1002_g N_VGND_c_730_n 0.00434272f $X=1.81 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A_M1005_g N_VGND_c_730_n 0.00383152f $X=2.31 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A_M1014_g N_VGND_c_731_n 0.00434272f $X=3.21 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A_M1016_g N_VGND_c_731_n 0.00383152f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A_M1002_g N_VGND_c_733_n 0.00825717f $X=1.81 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A_M1005_g N_VGND_c_733_n 0.00758198f $X=2.31 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A_M1014_g N_VGND_c_733_n 0.00825717f $X=3.21 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A_M1016_g N_VGND_c_733_n 0.00758198f $X=3.71 $Y=0.74 $X2=0 $Y2=0
cc_223 N_B_M1012_g N_A_27_368#_c_425_n 0.00342914f $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_224 N_B_c_269_n N_A_27_368#_c_425_n 0.00157102f $X=4.265 $Y=1.26 $X2=0 $Y2=0
cc_225 N_B_M1012_g N_A_27_368#_c_426_n 0.0103846f $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_226 N_B_M1013_g N_A_27_368#_c_426_n 5.42618e-19 $X=4.805 $Y=2.4 $X2=0 $Y2=0
cc_227 N_B_M1012_g N_A_27_368#_c_391_n 0.0119307f $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_228 N_B_M1013_g N_A_27_368#_c_391_n 0.0145175f $X=4.805 $Y=2.4 $X2=0 $Y2=0
cc_229 N_B_M1012_g N_A_27_368#_c_392_n 0.001916f $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_230 N_B_c_255_n N_A_27_368#_c_444_n 4.59311e-19 $X=5.215 $Y=1.26 $X2=0 $Y2=0
cc_231 N_B_M1017_g N_A_27_368#_c_393_n 0.0142213f $X=5.305 $Y=2.4 $X2=0 $Y2=0
cc_232 N_B_M1018_g N_A_27_368#_c_393_n 0.0140221f $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_233 N_B_M1018_g N_A_27_368#_c_394_n 3.74607e-19 $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_234 N_B_M1019_g N_A_27_368#_c_394_n 3.72209e-19 $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_235 N_B_c_264_n N_A_27_368#_c_394_n 3.5899e-19 $X=6.4 $Y=1.26 $X2=0 $Y2=0
cc_236 N_B_M1019_g N_A_27_368#_c_395_n 0.0140221f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_237 N_B_M1020_g N_A_27_368#_c_395_n 0.0142213f $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_238 N_B_M1020_g N_A_27_368#_c_396_n 4.28085e-19 $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_239 N_B_M1021_g N_A_27_368#_c_396_n 4.28085e-19 $X=7.155 $Y=2.4 $X2=0 $Y2=0
cc_240 N_B_M1021_g N_A_27_368#_c_397_n 0.0142213f $X=7.155 $Y=2.4 $X2=0 $Y2=0
cc_241 N_B_M1022_g N_A_27_368#_c_397_n 0.0150709f $X=7.605 $Y=2.4 $X2=0 $Y2=0
cc_242 N_B_M1022_g N_A_27_368#_c_398_n 0.00151912f $X=7.605 $Y=2.4 $X2=0 $Y2=0
cc_243 N_B_M1012_g N_VPWR_c_524_n 0.00333896f $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_244 N_B_M1013_g N_VPWR_c_524_n 0.00333926f $X=4.805 $Y=2.4 $X2=0 $Y2=0
cc_245 N_B_M1017_g N_VPWR_c_524_n 0.00333926f $X=5.305 $Y=2.4 $X2=0 $Y2=0
cc_246 N_B_M1018_g N_VPWR_c_524_n 0.00333926f $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_247 N_B_M1019_g N_VPWR_c_524_n 0.00333926f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_248 N_B_M1020_g N_VPWR_c_524_n 0.00333926f $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_249 N_B_M1021_g N_VPWR_c_524_n 0.00333926f $X=7.155 $Y=2.4 $X2=0 $Y2=0
cc_250 N_B_M1022_g N_VPWR_c_524_n 0.00333926f $X=7.605 $Y=2.4 $X2=0 $Y2=0
cc_251 N_B_M1012_g N_VPWR_c_515_n 0.00423284f $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_252 N_B_M1013_g N_VPWR_c_515_n 0.00423664f $X=4.805 $Y=2.4 $X2=0 $Y2=0
cc_253 N_B_M1017_g N_VPWR_c_515_n 0.00423176f $X=5.305 $Y=2.4 $X2=0 $Y2=0
cc_254 N_B_M1018_g N_VPWR_c_515_n 0.00422687f $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_255 N_B_M1019_g N_VPWR_c_515_n 0.00422687f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_256 N_B_M1020_g N_VPWR_c_515_n 0.00423176f $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_257 N_B_M1021_g N_VPWR_c_515_n 0.00423176f $X=7.155 $Y=2.4 $X2=0 $Y2=0
cc_258 N_B_M1022_g N_VPWR_c_515_n 0.00426591f $X=7.605 $Y=2.4 $X2=0 $Y2=0
cc_259 N_B_c_251_n N_Y_c_618_n 0.0148088f $X=4.21 $Y=1.185 $X2=0 $Y2=0
cc_260 N_B_M1012_g N_Y_c_623_n 0.00169841f $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_261 N_B_M1013_g N_Y_c_623_n 0.0135032f $X=4.805 $Y=2.4 $X2=0 $Y2=0
cc_262 N_B_M1017_g N_Y_c_623_n 6.43827e-19 $X=5.305 $Y=2.4 $X2=0 $Y2=0
cc_263 N_B_M1013_g N_Y_c_647_n 6.43827e-19 $X=4.805 $Y=2.4 $X2=0 $Y2=0
cc_264 N_B_M1017_g N_Y_c_647_n 0.0135194f $X=5.305 $Y=2.4 $X2=0 $Y2=0
cc_265 N_B_M1018_g N_Y_c_647_n 0.0122666f $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_266 N_B_M1019_g N_Y_c_647_n 3.7839e-19 $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_267 N_B_c_257_n N_Y_c_619_n 6.54586e-19 $X=5.325 $Y=1.185 $X2=0 $Y2=0
cc_268 N_B_c_260_n N_Y_c_619_n 0.0113581f $X=5.895 $Y=1.185 $X2=0 $Y2=0
cc_269 N_B_c_262_n N_Y_c_619_n 0.0102239f $X=6.325 $Y=1.185 $X2=0 $Y2=0
cc_270 N_B_M1018_g N_Y_c_654_n 7.64932e-19 $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_271 N_B_M1019_g N_Y_c_654_n 0.0163769f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_272 N_B_M1020_g N_Y_c_654_n 0.0165314f $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_273 N_B_M1021_g N_Y_c_654_n 7.44743e-19 $X=7.155 $Y=2.4 $X2=0 $Y2=0
cc_274 N_B_M1020_g N_Y_c_620_n 0.0136621f $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_275 N_B_c_266_n N_Y_c_620_n 0.00492465f $X=7.065 $Y=1.26 $X2=0 $Y2=0
cc_276 N_B_M1021_g N_Y_c_620_n 0.021071f $X=7.155 $Y=2.4 $X2=0 $Y2=0
cc_277 N_B_M1022_g N_Y_c_620_n 0.0105573f $X=7.605 $Y=2.4 $X2=0 $Y2=0
cc_278 N_B_c_273_n N_Y_c_620_n 0.00252388f $X=7.38 $Y=1.26 $X2=0 $Y2=0
cc_279 N_B_c_275_n N_Y_c_620_n 0.0282229f $X=7.39 $Y=0.465 $X2=0 $Y2=0
cc_280 N_B_c_251_n N_Y_c_621_n 0.0127495f $X=4.21 $Y=1.185 $X2=0 $Y2=0
cc_281 N_B_M1012_g N_Y_c_621_n 0.0150437f $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_282 N_B_c_253_n N_Y_c_621_n 0.0172053f $X=4.715 $Y=1.26 $X2=0 $Y2=0
cc_283 N_B_M1013_g N_Y_c_621_n 0.0237113f $X=4.805 $Y=2.4 $X2=0 $Y2=0
cc_284 N_B_c_255_n N_Y_c_621_n 0.0140604f $X=5.215 $Y=1.26 $X2=0 $Y2=0
cc_285 N_B_M1017_g N_Y_c_621_n 0.023828f $X=5.305 $Y=2.4 $X2=0 $Y2=0
cc_286 N_B_c_257_n N_Y_c_621_n 0.0190402f $X=5.325 $Y=1.185 $X2=0 $Y2=0
cc_287 N_B_c_258_n N_Y_c_621_n 0.00848084f $X=5.665 $Y=1.26 $X2=0 $Y2=0
cc_288 N_B_M1018_g N_Y_c_621_n 0.0216264f $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_289 N_B_c_260_n N_Y_c_621_n 0.00632967f $X=5.895 $Y=1.185 $X2=0 $Y2=0
cc_290 N_B_M1019_g N_Y_c_621_n 0.0195098f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_291 N_B_c_262_n N_Y_c_621_n 0.00260099f $X=6.325 $Y=1.185 $X2=0 $Y2=0
cc_292 N_B_c_264_n N_Y_c_621_n 0.0256234f $X=6.4 $Y=1.26 $X2=0 $Y2=0
cc_293 N_B_M1020_g N_Y_c_621_n 0.00382311f $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_294 N_B_c_269_n N_Y_c_621_n 0.0114296f $X=4.265 $Y=1.26 $X2=0 $Y2=0
cc_295 N_B_c_270_n N_Y_c_621_n 0.00706721f $X=4.805 $Y=1.26 $X2=0 $Y2=0
cc_296 N_B_c_271_n N_Y_c_621_n 0.00261306f $X=5.307 $Y=1.26 $X2=0 $Y2=0
cc_297 N_B_M1020_g N_Y_c_681_n 7.44743e-19 $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_298 N_B_M1021_g N_Y_c_681_n 0.0165314f $X=7.155 $Y=2.4 $X2=0 $Y2=0
cc_299 N_B_M1022_g N_Y_c_681_n 0.0207961f $X=7.605 $Y=2.4 $X2=0 $Y2=0
cc_300 N_B_c_251_n N_VGND_c_725_n 0.00571001f $X=4.21 $Y=1.185 $X2=0 $Y2=0
cc_301 N_B_c_251_n N_VGND_c_726_n 0.00433139f $X=4.21 $Y=1.185 $X2=0 $Y2=0
cc_302 N_B_c_257_n N_VGND_c_726_n 0.00433139f $X=5.325 $Y=1.185 $X2=0 $Y2=0
cc_303 N_B_c_257_n N_VGND_c_727_n 0.00701523f $X=5.325 $Y=1.185 $X2=0 $Y2=0
cc_304 N_B_c_258_n N_VGND_c_727_n 0.00167292f $X=5.665 $Y=1.26 $X2=0 $Y2=0
cc_305 N_B_c_260_n N_VGND_c_727_n 0.00563364f $X=5.895 $Y=1.185 $X2=0 $Y2=0
cc_306 N_B_c_260_n N_VGND_c_728_n 0.00434272f $X=5.895 $Y=1.185 $X2=0 $Y2=0
cc_307 N_B_c_262_n N_VGND_c_728_n 0.00434272f $X=6.325 $Y=1.185 $X2=0 $Y2=0
cc_308 N_B_c_262_n N_VGND_c_729_n 0.00963146f $X=6.325 $Y=1.185 $X2=0 $Y2=0
cc_309 N_B_c_263_n N_VGND_c_729_n 0.00981619f $X=6.565 $Y=1.26 $X2=0 $Y2=0
cc_310 N_B_c_274_n N_VGND_c_729_n 0.0104159f $X=7.39 $Y=0.465 $X2=0 $Y2=0
cc_311 N_B_c_275_n N_VGND_c_729_n 0.0317365f $X=7.39 $Y=0.465 $X2=0 $Y2=0
cc_312 N_B_c_274_n N_VGND_c_732_n 0.0127398f $X=7.39 $Y=0.465 $X2=0 $Y2=0
cc_313 N_B_c_275_n N_VGND_c_732_n 0.0172176f $X=7.39 $Y=0.465 $X2=0 $Y2=0
cc_314 N_B_c_251_n N_VGND_c_733_n 0.00822102f $X=4.21 $Y=1.185 $X2=0 $Y2=0
cc_315 N_B_c_257_n N_VGND_c_733_n 0.00822624f $X=5.325 $Y=1.185 $X2=0 $Y2=0
cc_316 N_B_c_260_n N_VGND_c_733_n 0.00821294f $X=5.895 $Y=1.185 $X2=0 $Y2=0
cc_317 N_B_c_262_n N_VGND_c_733_n 0.00825059f $X=6.325 $Y=1.185 $X2=0 $Y2=0
cc_318 N_B_c_274_n N_VGND_c_733_n 0.010606f $X=7.39 $Y=0.465 $X2=0 $Y2=0
cc_319 N_B_c_275_n N_VGND_c_733_n 0.0122345f $X=7.39 $Y=0.465 $X2=0 $Y2=0
cc_320 N_A_27_368#_c_386_n N_VPWR_M1001_s 0.00218982f $X=1.145 $Y=1.865
+ $X2=-0.19 $Y2=1.66
cc_321 N_A_27_368#_c_409_n N_VPWR_M1004_s 0.00313001f $X=2.045 $Y=2.035 $X2=0
+ $Y2=0
cc_322 N_A_27_368#_c_415_n N_VPWR_M1007_s 0.00408841f $X=2.995 $Y=2.035 $X2=0
+ $Y2=0
cc_323 N_A_27_368#_c_421_n N_VPWR_M1011_s 0.00513979f $X=3.915 $Y=2.035 $X2=0
+ $Y2=0
cc_324 N_A_27_368#_c_385_n N_VPWR_c_516_n 0.0330597f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_325 N_A_27_368#_c_386_n N_VPWR_c_516_n 0.0189268f $X=1.145 $Y=1.865 $X2=0
+ $Y2=0
cc_326 N_A_27_368#_c_388_n N_VPWR_c_516_n 0.0289706f $X=1.23 $Y=2.435 $X2=0
+ $Y2=0
cc_327 N_A_27_368#_c_388_n N_VPWR_c_517_n 0.0233699f $X=1.23 $Y=2.435 $X2=0
+ $Y2=0
cc_328 N_A_27_368#_c_409_n N_VPWR_c_517_n 0.0170259f $X=2.045 $Y=2.035 $X2=0
+ $Y2=0
cc_329 N_A_27_368#_c_389_n N_VPWR_c_517_n 0.0234083f $X=2.13 $Y=2.435 $X2=0
+ $Y2=0
cc_330 N_A_27_368#_c_389_n N_VPWR_c_518_n 0.0256025f $X=2.13 $Y=2.435 $X2=0
+ $Y2=0
cc_331 N_A_27_368#_c_415_n N_VPWR_c_518_n 0.0189268f $X=2.995 $Y=2.035 $X2=0
+ $Y2=0
cc_332 N_A_27_368#_c_390_n N_VPWR_c_518_n 0.0234083f $X=3.08 $Y=2.435 $X2=0
+ $Y2=0
cc_333 N_A_27_368#_c_390_n N_VPWR_c_519_n 0.0256025f $X=3.08 $Y=2.435 $X2=0
+ $Y2=0
cc_334 N_A_27_368#_c_421_n N_VPWR_c_519_n 0.0208278f $X=3.915 $Y=2.035 $X2=0
+ $Y2=0
cc_335 N_A_27_368#_c_392_n N_VPWR_c_519_n 0.0119238f $X=4.245 $Y=2.99 $X2=0
+ $Y2=0
cc_336 N_A_27_368#_c_385_n N_VPWR_c_520_n 0.014549f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_337 N_A_27_368#_c_388_n N_VPWR_c_521_n 0.00749631f $X=1.23 $Y=2.435 $X2=0
+ $Y2=0
cc_338 N_A_27_368#_c_389_n N_VPWR_c_522_n 0.0109793f $X=2.13 $Y=2.435 $X2=0
+ $Y2=0
cc_339 N_A_27_368#_c_390_n N_VPWR_c_523_n 0.0109793f $X=3.08 $Y=2.435 $X2=0
+ $Y2=0
cc_340 N_A_27_368#_c_391_n N_VPWR_c_524_n 0.0427884f $X=4.925 $Y=2.99 $X2=0
+ $Y2=0
cc_341 N_A_27_368#_c_392_n N_VPWR_c_524_n 0.0234458f $X=4.245 $Y=2.99 $X2=0
+ $Y2=0
cc_342 N_A_27_368#_c_393_n N_VPWR_c_524_n 0.0433424f $X=5.875 $Y=2.99 $X2=0
+ $Y2=0
cc_343 N_A_27_368#_c_395_n N_VPWR_c_524_n 0.0436645f $X=6.775 $Y=2.99 $X2=0
+ $Y2=0
cc_344 N_A_27_368#_c_397_n N_VPWR_c_524_n 0.0663548f $X=7.715 $Y=2.99 $X2=0
+ $Y2=0
cc_345 N_A_27_368#_c_400_n N_VPWR_c_524_n 0.0186386f $X=5.055 $Y=2.99 $X2=0
+ $Y2=0
cc_346 N_A_27_368#_c_401_n N_VPWR_c_524_n 0.0146958f $X=5.977 $Y=2.99 $X2=0
+ $Y2=0
cc_347 N_A_27_368#_c_402_n N_VPWR_c_524_n 0.0186386f $X=6.905 $Y=2.99 $X2=0
+ $Y2=0
cc_348 N_A_27_368#_c_385_n N_VPWR_c_515_n 0.0119743f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_349 N_A_27_368#_c_388_n N_VPWR_c_515_n 0.0062048f $X=1.23 $Y=2.435 $X2=0
+ $Y2=0
cc_350 N_A_27_368#_c_389_n N_VPWR_c_515_n 0.00901959f $X=2.13 $Y=2.435 $X2=0
+ $Y2=0
cc_351 N_A_27_368#_c_390_n N_VPWR_c_515_n 0.00901959f $X=3.08 $Y=2.435 $X2=0
+ $Y2=0
cc_352 N_A_27_368#_c_391_n N_VPWR_c_515_n 0.0240573f $X=4.925 $Y=2.99 $X2=0
+ $Y2=0
cc_353 N_A_27_368#_c_392_n N_VPWR_c_515_n 0.0125551f $X=4.245 $Y=2.99 $X2=0
+ $Y2=0
cc_354 N_A_27_368#_c_393_n N_VPWR_c_515_n 0.0242962f $X=5.875 $Y=2.99 $X2=0
+ $Y2=0
cc_355 N_A_27_368#_c_395_n N_VPWR_c_515_n 0.0244842f $X=6.775 $Y=2.99 $X2=0
+ $Y2=0
cc_356 N_A_27_368#_c_397_n N_VPWR_c_515_n 0.0367499f $X=7.715 $Y=2.99 $X2=0
+ $Y2=0
cc_357 N_A_27_368#_c_400_n N_VPWR_c_515_n 0.0101082f $X=5.055 $Y=2.99 $X2=0
+ $Y2=0
cc_358 N_A_27_368#_c_401_n N_VPWR_c_515_n 0.00796993f $X=5.977 $Y=2.99 $X2=0
+ $Y2=0
cc_359 N_A_27_368#_c_402_n N_VPWR_c_515_n 0.0101082f $X=6.905 $Y=2.99 $X2=0
+ $Y2=0
cc_360 N_A_27_368#_c_391_n N_Y_M1012_d 0.00218982f $X=4.925 $Y=2.99 $X2=0 $Y2=0
cc_361 N_A_27_368#_c_393_n N_Y_M1017_d 0.00165831f $X=5.875 $Y=2.99 $X2=0 $Y2=0
cc_362 N_A_27_368#_c_395_n N_Y_M1019_d 0.00165831f $X=6.775 $Y=2.99 $X2=0 $Y2=0
cc_363 N_A_27_368#_c_397_n N_Y_M1021_d 0.00165831f $X=7.715 $Y=2.99 $X2=0 $Y2=0
cc_364 N_A_27_368#_c_391_n N_Y_c_623_n 0.0177084f $X=4.925 $Y=2.99 $X2=0 $Y2=0
cc_365 N_A_27_368#_c_393_n N_Y_c_647_n 0.0159318f $X=5.875 $Y=2.99 $X2=0 $Y2=0
cc_366 N_A_27_368#_c_394_n N_Y_c_647_n 0.0335012f $X=5.98 $Y=1.985 $X2=0 $Y2=0
cc_367 N_A_27_368#_c_394_n N_Y_c_654_n 0.0327761f $X=5.98 $Y=1.985 $X2=0 $Y2=0
cc_368 N_A_27_368#_c_395_n N_Y_c_654_n 0.0159318f $X=6.775 $Y=2.99 $X2=0 $Y2=0
cc_369 N_A_27_368#_c_396_n N_Y_c_654_n 0.0335271f $X=6.93 $Y=1.985 $X2=0 $Y2=0
cc_370 N_A_27_368#_c_396_n N_Y_c_620_n 0.0217907f $X=6.93 $Y=1.985 $X2=0 $Y2=0
cc_371 N_A_27_368#_c_444_n N_Y_c_621_n 0.0213737f $X=5.08 $Y=2.115 $X2=0 $Y2=0
cc_372 N_A_27_368#_c_394_n N_Y_c_621_n 0.0189809f $X=5.98 $Y=1.985 $X2=0 $Y2=0
cc_373 N_A_27_368#_c_396_n N_Y_c_681_n 0.0335271f $X=6.93 $Y=1.985 $X2=0 $Y2=0
cc_374 N_A_27_368#_c_397_n N_Y_c_681_n 0.0159318f $X=7.715 $Y=2.99 $X2=0 $Y2=0
cc_375 N_A_27_368#_c_398_n N_Y_c_681_n 0.0351234f $X=7.88 $Y=1.985 $X2=0 $Y2=0
cc_376 N_A_27_368#_c_386_n N_VGND_c_723_n 0.0155831f $X=1.145 $Y=1.865 $X2=0
+ $Y2=0
cc_377 N_A_27_368#_c_399_n N_VGND_c_723_n 0.00609516f $X=1.23 $Y=1.865 $X2=0
+ $Y2=0
cc_378 N_Y_c_615_n N_VGND_M1005_d 0.00889788f $X=3.26 $Y=1.095 $X2=0 $Y2=0
cc_379 N_Y_c_618_n N_VGND_M1016_d 0.00250873f $X=4.26 $Y=1.095 $X2=0 $Y2=0
cc_380 N_Y_c_614_n N_VGND_c_723_n 0.0256093f $X=2.025 $Y=0.515 $X2=0 $Y2=0
cc_381 N_Y_c_616_n N_VGND_c_723_n 0.00594067f $X=2.19 $Y=1.095 $X2=0 $Y2=0
cc_382 N_Y_c_614_n N_VGND_c_724_n 0.0213338f $X=2.025 $Y=0.515 $X2=0 $Y2=0
cc_383 N_Y_c_615_n N_VGND_c_724_n 0.0535301f $X=3.26 $Y=1.095 $X2=0 $Y2=0
cc_384 N_Y_c_617_n N_VGND_c_724_n 0.019268f $X=3.425 $Y=0.515 $X2=0 $Y2=0
cc_385 N_Y_c_617_n N_VGND_c_725_n 0.0191765f $X=3.425 $Y=0.515 $X2=0 $Y2=0
cc_386 N_Y_c_618_n N_VGND_c_725_n 0.0209867f $X=4.26 $Y=1.095 $X2=0 $Y2=0
cc_387 N_Y_c_621_n N_VGND_c_725_n 0.0214346f $X=6.595 $Y=1.565 $X2=0 $Y2=0
cc_388 N_Y_c_621_n N_VGND_c_726_n 0.0451408f $X=6.595 $Y=1.565 $X2=0 $Y2=0
cc_389 N_Y_c_619_n N_VGND_c_727_n 0.0240544f $X=6.11 $Y=0.515 $X2=0 $Y2=0
cc_390 N_Y_c_621_n N_VGND_c_727_n 0.0560141f $X=6.595 $Y=1.565 $X2=0 $Y2=0
cc_391 N_Y_c_619_n N_VGND_c_728_n 0.0144922f $X=6.11 $Y=0.515 $X2=0 $Y2=0
cc_392 N_Y_c_619_n N_VGND_c_729_n 0.0308485f $X=6.11 $Y=0.515 $X2=0 $Y2=0
cc_393 N_Y_c_620_n N_VGND_c_729_n 0.0085367f $X=7.215 $Y=1.565 $X2=0 $Y2=0
cc_394 N_Y_c_621_n N_VGND_c_729_n 0.00828005f $X=6.595 $Y=1.565 $X2=0 $Y2=0
cc_395 N_Y_c_614_n N_VGND_c_730_n 0.0145639f $X=2.025 $Y=0.515 $X2=0 $Y2=0
cc_396 N_Y_c_617_n N_VGND_c_731_n 0.0145639f $X=3.425 $Y=0.515 $X2=0 $Y2=0
cc_397 N_Y_c_614_n N_VGND_c_733_n 0.0119984f $X=2.025 $Y=0.515 $X2=0 $Y2=0
cc_398 N_Y_c_617_n N_VGND_c_733_n 0.0119984f $X=3.425 $Y=0.515 $X2=0 $Y2=0
cc_399 N_Y_c_619_n N_VGND_c_733_n 0.0118826f $X=6.11 $Y=0.515 $X2=0 $Y2=0
cc_400 N_Y_c_621_n N_VGND_c_733_n 0.0372462f $X=6.595 $Y=1.565 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__a311o_1.pxi.spice
* Created: Fri Aug 28 17:05:23 2020
* 
x_PM_SKY130_FD_SC_MS__A311O_1%A_89_270# N_A_89_270#_M1007_d N_A_89_270#_M1003_d
+ N_A_89_270#_M1005_d N_A_89_270#_M1010_g N_A_89_270#_c_75_n N_A_89_270#_M1006_g
+ N_A_89_270#_c_76_n N_A_89_270#_c_77_n N_A_89_270#_c_78_n N_A_89_270#_c_86_n
+ N_A_89_270#_c_79_n N_A_89_270#_c_80_n N_A_89_270#_c_87_n N_A_89_270#_c_81_n
+ N_A_89_270#_c_82_n N_A_89_270#_c_83_n PM_SKY130_FD_SC_MS__A311O_1%A_89_270#
x_PM_SKY130_FD_SC_MS__A311O_1%A3 N_A3_M1000_g N_A3_M1004_g A3 N_A3_c_176_n
+ PM_SKY130_FD_SC_MS__A311O_1%A3
x_PM_SKY130_FD_SC_MS__A311O_1%A2 N_A2_M1002_g N_A2_M1011_g A2 N_A2_c_212_n
+ PM_SKY130_FD_SC_MS__A311O_1%A2
x_PM_SKY130_FD_SC_MS__A311O_1%A1 N_A1_M1007_g N_A1_c_245_n N_A1_M1008_g A1 A1
+ N_A1_c_247_n N_A1_c_248_n N_A1_c_249_n PM_SKY130_FD_SC_MS__A311O_1%A1
x_PM_SKY130_FD_SC_MS__A311O_1%B1 N_B1_M1001_g N_B1_M1009_g N_B1_c_296_n B1
+ N_B1_c_298_n PM_SKY130_FD_SC_MS__A311O_1%B1
x_PM_SKY130_FD_SC_MS__A311O_1%C1 N_C1_M1005_g N_C1_M1003_g N_C1_c_337_n
+ N_C1_c_338_n C1 N_C1_c_339_n N_C1_c_340_n PM_SKY130_FD_SC_MS__A311O_1%C1
x_PM_SKY130_FD_SC_MS__A311O_1%X N_X_M1006_s N_X_M1010_s N_X_c_375_n N_X_c_376_n
+ X X X X N_X_c_377_n PM_SKY130_FD_SC_MS__A311O_1%X
x_PM_SKY130_FD_SC_MS__A311O_1%VPWR N_VPWR_M1010_d N_VPWR_M1002_d N_VPWR_c_397_n
+ N_VPWR_c_398_n N_VPWR_c_399_n N_VPWR_c_400_n VPWR N_VPWR_c_401_n
+ N_VPWR_c_396_n N_VPWR_c_403_n PM_SKY130_FD_SC_MS__A311O_1%VPWR
x_PM_SKY130_FD_SC_MS__A311O_1%A_261_392# N_A_261_392#_M1000_d
+ N_A_261_392#_M1008_d N_A_261_392#_c_439_n N_A_261_392#_c_440_n
+ N_A_261_392#_c_441_n N_A_261_392#_c_442_n N_A_261_392#_c_443_n
+ PM_SKY130_FD_SC_MS__A311O_1%A_261_392#
x_PM_SKY130_FD_SC_MS__A311O_1%VGND N_VGND_M1006_d N_VGND_M1001_d N_VGND_c_480_n
+ N_VGND_c_481_n N_VGND_c_482_n N_VGND_c_483_n VGND N_VGND_c_484_n
+ N_VGND_c_485_n N_VGND_c_486_n N_VGND_c_487_n PM_SKY130_FD_SC_MS__A311O_1%VGND
cc_1 VNB N_A_89_270#_c_75_n 0.0215076f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.35
cc_2 VNB N_A_89_270#_c_76_n 0.0109532f $X=-0.19 $Y=-0.245 $X2=2.24 $Y2=1.195
cc_3 VNB N_A_89_270#_c_77_n 0.00627074f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.195
cc_4 VNB N_A_89_270#_c_78_n 0.0106288f $X=-0.19 $Y=-0.245 $X2=3.245 $Y2=1.53
cc_5 VNB N_A_89_270#_c_79_n 0.0175711f $X=-0.19 $Y=-0.245 $X2=3.41 $Y2=1.105
cc_6 VNB N_A_89_270#_c_80_n 0.003271f $X=-0.19 $Y=-0.245 $X2=2.405 $Y2=1.005
cc_7 VNB N_A_89_270#_c_81_n 0.00228403f $X=-0.19 $Y=-0.245 $X2=3.34 $Y2=1.94
cc_8 VNB N_A_89_270#_c_82_n 0.00770964f $X=-0.19 $Y=-0.245 $X2=3.41 $Y2=1.53
cc_9 VNB N_A_89_270#_c_83_n 0.0294391f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.515
cc_10 VNB N_A3_M1004_g 0.0239645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB A3 9.08959e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A3_c_176_n 0.0191325f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_13 VNB N_A2_M1011_g 0.0208933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB A2 0.00320338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_c_212_n 0.016088f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_16 VNB N_A1_M1007_g 0.00828724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_c_245_n 0.005531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_M1008_g 0.011874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_247_n 0.0466861f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.87
cc_20 VNB N_A1_c_248_n 9.2097e-19 $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.87
cc_21 VNB N_A1_c_249_n 0.00608405f $X=-0.19 $Y=-0.245 $X2=3.245 $Y2=1.53
cc_22 VNB N_B1_M1001_g 0.00907604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B1_M1009_g 0.00809716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B1_c_296_n 0.0100012f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.68
cc_25 VNB B1 0.00737349f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_26 VNB N_B1_c_298_n 0.0353796f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.35
cc_27 VNB N_C1_M1005_g 0.0103317f $X=-0.19 $Y=-0.245 $X2=3.135 $Y2=1.96
cc_28 VNB N_C1_M1003_g 0.0111186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_C1_c_337_n 0.0199494f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_30 VNB N_C1_c_338_n 0.0137028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_C1_c_339_n 0.0599949f $X=-0.19 $Y=-0.245 $X2=2.24 $Y2=1.195
cc_32 VNB N_C1_c_340_n 0.0126535f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.195
cc_33 VNB N_X_c_375_n 0.0182499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_376_n 0.0228556f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_35 VNB N_X_c_377_n 0.0234973f $X=-0.19 $Y=-0.245 $X2=2.405 $Y2=1.005
cc_36 VNB N_VPWR_c_396_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.515
cc_37 VNB N_VGND_c_480_n 0.0203545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_481_n 0.00567404f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_39 VNB N_VGND_c_482_n 0.0256231f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.35
cc_40 VNB N_VGND_c_483_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.87
cc_41 VNB N_VGND_c_484_n 0.0507439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_485_n 0.0181991f $X=-0.19 $Y=-0.245 $X2=3.41 $Y2=1.94
cc_43 VNB N_VGND_c_486_n 0.249518f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.195
cc_44 VNB N_VGND_c_487_n 0.00270401f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.515
cc_45 VPB N_A_89_270#_M1010_g 0.0282035f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.4
cc_46 VPB N_A_89_270#_c_77_n 0.00421697f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.195
cc_47 VPB N_A_89_270#_c_86_n 0.0404369f $X=-0.19 $Y=1.66 $X2=3.27 $Y2=2.815
cc_48 VPB N_A_89_270#_c_87_n 0.0115428f $X=-0.19 $Y=1.66 $X2=3.27 $Y2=2.105
cc_49 VPB N_A_89_270#_c_81_n 0.0158759f $X=-0.19 $Y=1.66 $X2=3.34 $Y2=1.94
cc_50 VPB N_A_89_270#_c_83_n 0.00675718f $X=-0.19 $Y=1.66 $X2=0.735 $Y2=1.515
cc_51 VPB N_A3_M1000_g 0.0256571f $X=-0.19 $Y=1.66 $X2=3.135 $Y2=1.96
cc_52 VPB A3 8.81819e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A3_c_176_n 0.0131733f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.4
cc_54 VPB N_A2_M1002_g 0.0242687f $X=-0.19 $Y=1.66 $X2=3.135 $Y2=1.96
cc_55 VPB A2 0.00214309f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A2_c_212_n 0.0103295f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.4
cc_57 VPB N_A1_M1008_g 0.0307961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_B1_M1009_g 0.0291714f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_C1_M1005_g 0.0338431f $X=-0.19 $Y=1.66 $X2=3.135 $Y2=1.96
cc_60 VPB X 0.00695105f $X=-0.19 $Y=1.66 $X2=2.24 $Y2=1.195
cc_61 VPB X 0.0406888f $X=-0.19 $Y=1.66 $X2=3.41 $Y2=1.105
cc_62 VPB N_X_c_377_n 0.0090928f $X=-0.19 $Y=1.66 $X2=2.405 $Y2=1.005
cc_63 VPB N_VPWR_c_397_n 0.0142832f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.4
cc_64 VPB N_VPWR_c_398_n 0.00931005f $X=-0.19 $Y=1.66 $X2=2.24 $Y2=1.195
cc_65 VPB N_VPWR_c_399_n 0.0196495f $X=-0.19 $Y=1.66 $X2=2.57 $Y2=1.53
cc_66 VPB N_VPWR_c_400_n 0.00555219f $X=-0.19 $Y=1.66 $X2=3.34 $Y2=2.175
cc_67 VPB N_VPWR_c_401_n 0.0514544f $X=-0.19 $Y=1.66 $X2=0.712 $Y2=1.515
cc_68 VPB N_VPWR_c_396_n 0.0752344f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.515
cc_69 VPB N_VPWR_c_403_n 0.028772f $X=-0.19 $Y=1.66 $X2=2.405 $Y2=1.005
cc_70 VPB N_A_261_392#_c_439_n 0.00394251f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_261_392#_c_440_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_261_392#_c_441_n 0.00442833f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.4
cc_73 VPB N_A_261_392#_c_442_n 0.00320906f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_261_392#_c_443_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.735 $Y2=0.87
cc_75 N_A_89_270#_M1010_g N_A3_M1000_g 0.0215268f $X=0.535 $Y=2.4 $X2=0 $Y2=0
cc_76 N_A_89_270#_c_75_n N_A3_M1004_g 0.0233429f $X=0.735 $Y=1.35 $X2=0 $Y2=0
cc_77 N_A_89_270#_c_76_n N_A3_M1004_g 0.0154265f $X=2.24 $Y=1.195 $X2=0 $Y2=0
cc_78 N_A_89_270#_c_77_n N_A3_M1004_g 0.00384761f $X=0.945 $Y=1.195 $X2=0 $Y2=0
cc_79 N_A_89_270#_M1010_g A3 5.05051e-19 $X=0.535 $Y=2.4 $X2=0 $Y2=0
cc_80 N_A_89_270#_c_76_n A3 0.0181696f $X=2.24 $Y=1.195 $X2=0 $Y2=0
cc_81 N_A_89_270#_c_77_n A3 0.0184377f $X=0.945 $Y=1.195 $X2=0 $Y2=0
cc_82 N_A_89_270#_M1010_g N_A3_c_176_n 0.003303f $X=0.535 $Y=2.4 $X2=0 $Y2=0
cc_83 N_A_89_270#_c_76_n N_A3_c_176_n 0.00302365f $X=2.24 $Y=1.195 $X2=0 $Y2=0
cc_84 N_A_89_270#_c_77_n N_A3_c_176_n 0.00163481f $X=0.945 $Y=1.195 $X2=0 $Y2=0
cc_85 N_A_89_270#_c_83_n N_A3_c_176_n 0.0130342f $X=0.735 $Y=1.515 $X2=0 $Y2=0
cc_86 N_A_89_270#_c_76_n N_A2_M1011_g 0.0122853f $X=2.24 $Y=1.195 $X2=0 $Y2=0
cc_87 N_A_89_270#_c_80_n N_A2_M1011_g 0.00218849f $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_88 N_A_89_270#_c_76_n A2 0.0250329f $X=2.24 $Y=1.195 $X2=0 $Y2=0
cc_89 N_A_89_270#_c_80_n A2 0.00718333f $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_90 N_A_89_270#_c_76_n N_A2_c_212_n 0.00431149f $X=2.24 $Y=1.195 $X2=0 $Y2=0
cc_91 N_A_89_270#_c_76_n N_A1_M1007_g 0.011152f $X=2.24 $Y=1.195 $X2=0 $Y2=0
cc_92 N_A_89_270#_c_80_n N_A1_M1007_g 0.00877504f $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_93 N_A_89_270#_c_80_n N_A1_c_245_n 0.00358622f $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_94 N_A_89_270#_c_80_n N_A1_M1008_g 0.00660486f $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_95 N_A_89_270#_c_76_n N_A1_c_247_n 3.32499e-19 $X=2.24 $Y=1.195 $X2=0 $Y2=0
cc_96 N_A_89_270#_c_80_n N_A1_c_247_n 2.43363e-19 $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_97 N_A_89_270#_M1007_d N_A1_c_248_n 6.27105e-19 $X=2.265 $Y=0.615 $X2=0 $Y2=0
cc_98 N_A_89_270#_c_76_n N_A1_c_248_n 0.00623312f $X=2.24 $Y=1.195 $X2=0 $Y2=0
cc_99 N_A_89_270#_c_80_n N_A1_c_248_n 0.00288651f $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_100 N_A_89_270#_c_76_n N_A1_c_249_n 0.0113079f $X=2.24 $Y=1.195 $X2=0 $Y2=0
cc_101 N_A_89_270#_c_79_n N_B1_M1001_g 4.84241e-19 $X=3.41 $Y=1.105 $X2=0 $Y2=0
cc_102 N_A_89_270#_c_80_n N_B1_M1001_g 0.00848117f $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_103 N_A_89_270#_c_78_n N_B1_M1009_g 0.0108987f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_104 N_A_89_270#_c_80_n N_B1_M1009_g 0.00197044f $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_105 N_A_89_270#_c_87_n N_B1_M1009_g 0.00282815f $X=3.27 $Y=2.105 $X2=0 $Y2=0
cc_106 N_A_89_270#_c_78_n N_B1_c_296_n 0.00839397f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_107 N_A_89_270#_c_79_n N_B1_c_296_n 2.58467e-19 $X=3.41 $Y=1.105 $X2=0 $Y2=0
cc_108 N_A_89_270#_c_80_n N_B1_c_296_n 0.00446272f $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_109 N_A_89_270#_c_80_n B1 0.00186884f $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_110 N_A_89_270#_c_78_n N_C1_M1005_g 0.0135718f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_111 N_A_89_270#_c_86_n N_C1_M1005_g 0.0150763f $X=3.27 $Y=2.815 $X2=0 $Y2=0
cc_112 N_A_89_270#_c_87_n N_C1_M1005_g 0.00517796f $X=3.27 $Y=2.105 $X2=0 $Y2=0
cc_113 N_A_89_270#_c_81_n N_C1_M1005_g 0.0130735f $X=3.34 $Y=1.94 $X2=0 $Y2=0
cc_114 N_A_89_270#_c_79_n N_C1_M1003_g 0.00737166f $X=3.41 $Y=1.105 $X2=0 $Y2=0
cc_115 N_A_89_270#_c_80_n N_C1_M1003_g 5.26759e-19 $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_116 N_A_89_270#_c_78_n N_C1_c_337_n 0.00906085f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_117 N_A_89_270#_c_79_n N_C1_c_337_n 0.00493627f $X=3.41 $Y=1.105 $X2=0 $Y2=0
cc_118 N_A_89_270#_c_80_n N_C1_c_337_n 4.1554e-19 $X=2.405 $Y=1.005 $X2=0 $Y2=0
cc_119 N_A_89_270#_c_87_n N_C1_c_337_n 6.35295e-19 $X=3.27 $Y=2.105 $X2=0 $Y2=0
cc_120 N_A_89_270#_c_82_n N_C1_c_337_n 0.00141795f $X=3.41 $Y=1.53 $X2=0 $Y2=0
cc_121 N_A_89_270#_c_79_n N_C1_c_339_n 0.00363944f $X=3.41 $Y=1.105 $X2=0 $Y2=0
cc_122 N_A_89_270#_M1003_d N_C1_c_340_n 0.00273424f $X=3.27 $Y=0.615 $X2=0 $Y2=0
cc_123 N_A_89_270#_c_79_n N_C1_c_340_n 0.00981852f $X=3.41 $Y=1.105 $X2=0 $Y2=0
cc_124 N_A_89_270#_c_77_n N_X_c_375_n 0.00920337f $X=0.945 $Y=1.195 $X2=0 $Y2=0
cc_125 N_A_89_270#_c_83_n N_X_c_375_n 0.00202112f $X=0.735 $Y=1.515 $X2=0 $Y2=0
cc_126 N_A_89_270#_c_75_n N_X_c_376_n 4.43891e-19 $X=0.735 $Y=1.35 $X2=0 $Y2=0
cc_127 N_A_89_270#_M1010_g X 0.00385747f $X=0.535 $Y=2.4 $X2=0 $Y2=0
cc_128 N_A_89_270#_M1010_g X 0.0120548f $X=0.535 $Y=2.4 $X2=0 $Y2=0
cc_129 N_A_89_270#_c_75_n N_X_c_377_n 0.00256161f $X=0.735 $Y=1.35 $X2=0 $Y2=0
cc_130 N_A_89_270#_c_77_n N_X_c_377_n 0.0299346f $X=0.945 $Y=1.195 $X2=0 $Y2=0
cc_131 N_A_89_270#_c_83_n N_X_c_377_n 0.0136465f $X=0.735 $Y=1.515 $X2=0 $Y2=0
cc_132 N_A_89_270#_M1010_g N_VPWR_c_397_n 0.0115992f $X=0.535 $Y=2.4 $X2=0 $Y2=0
cc_133 N_A_89_270#_c_76_n N_VPWR_c_397_n 0.00508495f $X=2.24 $Y=1.195 $X2=0
+ $Y2=0
cc_134 N_A_89_270#_c_77_n N_VPWR_c_397_n 0.0173496f $X=0.945 $Y=1.195 $X2=0
+ $Y2=0
cc_135 N_A_89_270#_c_83_n N_VPWR_c_397_n 0.00107868f $X=0.735 $Y=1.515 $X2=0
+ $Y2=0
cc_136 N_A_89_270#_c_86_n N_VPWR_c_401_n 0.0207959f $X=3.27 $Y=2.815 $X2=0 $Y2=0
cc_137 N_A_89_270#_M1010_g N_VPWR_c_396_n 0.00987339f $X=0.535 $Y=2.4 $X2=0
+ $Y2=0
cc_138 N_A_89_270#_c_86_n N_VPWR_c_396_n 0.0171449f $X=3.27 $Y=2.815 $X2=0 $Y2=0
cc_139 N_A_89_270#_M1010_g N_VPWR_c_403_n 0.005209f $X=0.535 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A_89_270#_c_76_n N_A_261_392#_c_439_n 0.00649318f $X=2.24 $Y=1.195
+ $X2=0 $Y2=0
cc_141 N_A_89_270#_c_76_n N_A_261_392#_c_441_n 0.00875899f $X=2.24 $Y=1.195
+ $X2=0 $Y2=0
cc_142 N_A_89_270#_c_80_n N_A_261_392#_c_441_n 0.00103949f $X=2.405 $Y=1.005
+ $X2=0 $Y2=0
cc_143 N_A_89_270#_c_78_n N_A_261_392#_c_442_n 0.00113092f $X=3.245 $Y=1.53
+ $X2=0 $Y2=0
cc_144 N_A_89_270#_c_80_n N_A_261_392#_c_442_n 0.0177922f $X=2.405 $Y=1.005
+ $X2=0 $Y2=0
cc_145 N_A_89_270#_c_87_n N_A_261_392#_c_442_n 0.00597448f $X=3.27 $Y=2.105
+ $X2=0 $Y2=0
cc_146 N_A_89_270#_c_87_n N_A_261_392#_c_443_n 0.0270058f $X=3.27 $Y=2.105 $X2=0
+ $Y2=0
cc_147 N_A_89_270#_c_76_n N_VGND_M1006_d 0.00177524f $X=2.24 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_148 N_A_89_270#_c_77_n N_VGND_M1006_d 8.58534e-19 $X=0.945 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_149 N_A_89_270#_c_75_n N_VGND_c_480_n 0.0140304f $X=0.735 $Y=1.35 $X2=0 $Y2=0
cc_150 N_A_89_270#_c_76_n N_VGND_c_480_n 0.0136318f $X=2.24 $Y=1.195 $X2=0 $Y2=0
cc_151 N_A_89_270#_c_77_n N_VGND_c_480_n 0.00890417f $X=0.945 $Y=1.195 $X2=0
+ $Y2=0
cc_152 N_A_89_270#_c_78_n N_VGND_c_481_n 0.0212375f $X=3.245 $Y=1.53 $X2=0 $Y2=0
cc_153 N_A_89_270#_c_80_n N_VGND_c_481_n 6.88425e-19 $X=2.405 $Y=1.005 $X2=0
+ $Y2=0
cc_154 N_A_89_270#_c_75_n N_VGND_c_482_n 0.00405273f $X=0.735 $Y=1.35 $X2=0
+ $Y2=0
cc_155 N_A_89_270#_c_75_n N_VGND_c_486_n 0.00424518f $X=0.735 $Y=1.35 $X2=0
+ $Y2=0
cc_156 N_A_89_270#_c_80_n N_VGND_c_486_n 0.00775516f $X=2.405 $Y=1.005 $X2=0
+ $Y2=0
cc_157 N_A_89_270#_c_76_n A_264_120# 0.00756132f $X=2.24 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_158 N_A_89_270#_c_76_n A_359_123# 0.00335572f $X=2.24 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_159 N_A3_M1000_g N_A2_M1002_g 0.0155375f $X=1.215 $Y=2.46 $X2=0 $Y2=0
cc_160 N_A3_M1004_g N_A2_M1011_g 0.0378038f $X=1.245 $Y=0.92 $X2=0 $Y2=0
cc_161 A3 A2 0.0226838f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_162 N_A3_c_176_n A2 0.00187659f $X=1.2 $Y=1.615 $X2=0 $Y2=0
cc_163 A3 N_A2_c_212_n 4.06578e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_164 N_A3_c_176_n N_A2_c_212_n 0.0207467f $X=1.2 $Y=1.615 $X2=0 $Y2=0
cc_165 N_A3_M1004_g N_A1_c_249_n 0.00181953f $X=1.245 $Y=0.92 $X2=0 $Y2=0
cc_166 N_A3_M1000_g X 5.91015e-19 $X=1.215 $Y=2.46 $X2=0 $Y2=0
cc_167 N_A3_M1000_g N_VPWR_c_397_n 0.0116329f $X=1.215 $Y=2.46 $X2=0 $Y2=0
cc_168 N_A3_c_176_n N_VPWR_c_397_n 0.00208216f $X=1.2 $Y=1.615 $X2=0 $Y2=0
cc_169 N_A3_M1000_g N_VPWR_c_399_n 0.005209f $X=1.215 $Y=2.46 $X2=0 $Y2=0
cc_170 N_A3_M1000_g N_VPWR_c_396_n 0.00983608f $X=1.215 $Y=2.46 $X2=0 $Y2=0
cc_171 N_A3_M1000_g N_A_261_392#_c_439_n 0.00249896f $X=1.215 $Y=2.46 $X2=0
+ $Y2=0
cc_172 A3 N_A_261_392#_c_439_n 0.00740718f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_173 N_A3_c_176_n N_A_261_392#_c_439_n 4.65552e-19 $X=1.2 $Y=1.615 $X2=0 $Y2=0
cc_174 N_A3_M1000_g N_A_261_392#_c_440_n 0.0103799f $X=1.215 $Y=2.46 $X2=0 $Y2=0
cc_175 N_A3_M1004_g N_VGND_c_480_n 0.00343181f $X=1.245 $Y=0.92 $X2=0 $Y2=0
cc_176 N_A3_M1004_g N_VGND_c_484_n 0.00428744f $X=1.245 $Y=0.92 $X2=0 $Y2=0
cc_177 N_A3_M1004_g N_VGND_c_486_n 0.00476395f $X=1.245 $Y=0.92 $X2=0 $Y2=0
cc_178 N_A2_M1011_g N_A1_M1007_g 0.0378467f $X=1.72 $Y=0.935 $X2=0 $Y2=0
cc_179 N_A2_M1002_g N_A1_M1008_g 0.0289122f $X=1.665 $Y=2.46 $X2=0 $Y2=0
cc_180 A2 N_A1_M1008_g 0.00167797f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_181 N_A2_c_212_n N_A1_M1008_g 0.0198993f $X=1.74 $Y=1.615 $X2=0 $Y2=0
cc_182 N_A2_M1011_g N_A1_c_247_n 0.00129249f $X=1.72 $Y=0.935 $X2=0 $Y2=0
cc_183 N_A2_M1011_g N_A1_c_249_n 0.0113054f $X=1.72 $Y=0.935 $X2=0 $Y2=0
cc_184 N_A2_M1002_g N_VPWR_c_398_n 0.00321888f $X=1.665 $Y=2.46 $X2=0 $Y2=0
cc_185 N_A2_M1002_g N_VPWR_c_399_n 0.005209f $X=1.665 $Y=2.46 $X2=0 $Y2=0
cc_186 N_A2_M1002_g N_VPWR_c_396_n 0.00983279f $X=1.665 $Y=2.46 $X2=0 $Y2=0
cc_187 N_A2_M1002_g N_A_261_392#_c_439_n 0.00100213f $X=1.665 $Y=2.46 $X2=0
+ $Y2=0
cc_188 A2 N_A_261_392#_c_439_n 0.00327936f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_189 N_A2_M1002_g N_A_261_392#_c_440_n 0.0123627f $X=1.665 $Y=2.46 $X2=0 $Y2=0
cc_190 N_A2_M1002_g N_A_261_392#_c_441_n 0.0133817f $X=1.665 $Y=2.46 $X2=0 $Y2=0
cc_191 A2 N_A_261_392#_c_441_n 0.0219515f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_192 N_A2_c_212_n N_A_261_392#_c_441_n 0.00352068f $X=1.74 $Y=1.615 $X2=0
+ $Y2=0
cc_193 N_A2_M1002_g N_A_261_392#_c_443_n 6.0235e-19 $X=1.665 $Y=2.46 $X2=0 $Y2=0
cc_194 N_A2_M1011_g N_VGND_c_484_n 6.8294e-19 $X=1.72 $Y=0.935 $X2=0 $Y2=0
cc_195 N_A1_M1007_g N_B1_M1001_g 0.0198607f $X=2.19 $Y=0.935 $X2=0 $Y2=0
cc_196 N_A1_c_248_n N_B1_M1001_g 5.66657e-19 $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_197 N_A1_M1008_g N_B1_M1009_g 0.0307367f $X=2.205 $Y=2.46 $X2=0 $Y2=0
cc_198 N_A1_c_245_n N_B1_c_296_n 0.00777372f $X=2.205 $Y=1.42 $X2=0 $Y2=0
cc_199 N_A1_M1007_g B1 3.45758e-19 $X=2.19 $Y=0.935 $X2=0 $Y2=0
cc_200 N_A1_c_247_n B1 0.00143004f $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_201 N_A1_c_248_n B1 0.0285655f $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_202 N_A1_c_247_n N_B1_c_298_n 0.0213815f $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_203 N_A1_c_248_n N_B1_c_298_n 3.01834e-19 $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_204 N_A1_M1008_g N_VPWR_c_398_n 0.00726917f $X=2.205 $Y=2.46 $X2=0 $Y2=0
cc_205 N_A1_M1008_g N_VPWR_c_401_n 0.005209f $X=2.205 $Y=2.46 $X2=0 $Y2=0
cc_206 N_A1_M1008_g N_VPWR_c_396_n 0.00982607f $X=2.205 $Y=2.46 $X2=0 $Y2=0
cc_207 N_A1_M1008_g N_A_261_392#_c_440_n 6.97719e-19 $X=2.205 $Y=2.46 $X2=0
+ $Y2=0
cc_208 N_A1_M1008_g N_A_261_392#_c_441_n 0.0154068f $X=2.205 $Y=2.46 $X2=0 $Y2=0
cc_209 N_A1_M1008_g N_A_261_392#_c_442_n 0.00150612f $X=2.205 $Y=2.46 $X2=0
+ $Y2=0
cc_210 N_A1_M1008_g N_A_261_392#_c_443_n 0.0118717f $X=2.205 $Y=2.46 $X2=0 $Y2=0
cc_211 N_A1_c_249_n N_VGND_c_480_n 0.00827599f $X=2.005 $Y=0.555 $X2=0 $Y2=0
cc_212 N_A1_c_247_n N_VGND_c_484_n 0.0066215f $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_213 N_A1_c_248_n N_VGND_c_484_n 0.0215843f $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_214 N_A1_c_249_n N_VGND_c_484_n 0.0132973f $X=2.005 $Y=0.555 $X2=0 $Y2=0
cc_215 N_A1_c_247_n N_VGND_c_486_n 0.00960263f $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_216 N_A1_c_248_n N_VGND_c_486_n 0.0110944f $X=2.17 $Y=0.34 $X2=0 $Y2=0
cc_217 N_A1_c_249_n N_VGND_c_486_n 0.0147336f $X=2.005 $Y=0.555 $X2=0 $Y2=0
cc_218 N_A1_c_249_n A_264_120# 0.00131491f $X=2.005 $Y=0.555 $X2=-0.19
+ $Y2=-0.245
cc_219 N_A1_c_248_n A_359_123# 0.00103536f $X=2.17 $Y=0.34 $X2=-0.19 $Y2=-0.245
cc_220 N_A1_c_249_n A_359_123# 0.00273639f $X=2.005 $Y=0.555 $X2=-0.19
+ $Y2=-0.245
cc_221 N_B1_M1009_g N_C1_M1005_g 0.0538715f $X=2.655 $Y=2.46 $X2=0 $Y2=0
cc_222 N_B1_M1001_g N_C1_M1003_g 0.0179711f $X=2.62 $Y=0.935 $X2=0 $Y2=0
cc_223 B1 N_C1_M1003_g 4.01526e-19 $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_224 N_B1_c_296_n N_C1_c_337_n 0.0538715f $X=2.645 $Y=1.48 $X2=0 $Y2=0
cc_225 B1 N_C1_c_338_n 2.72693e-19 $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_226 N_B1_c_298_n N_C1_c_338_n 0.0179383f $X=2.71 $Y=0.34 $X2=0 $Y2=0
cc_227 N_B1_M1009_g N_VPWR_c_401_n 0.005209f $X=2.655 $Y=2.46 $X2=0 $Y2=0
cc_228 N_B1_M1009_g N_VPWR_c_396_n 0.0098298f $X=2.655 $Y=2.46 $X2=0 $Y2=0
cc_229 N_B1_M1009_g N_A_261_392#_c_442_n 0.00396143f $X=2.655 $Y=2.46 $X2=0
+ $Y2=0
cc_230 N_B1_M1009_g N_A_261_392#_c_443_n 0.015809f $X=2.655 $Y=2.46 $X2=0 $Y2=0
cc_231 N_B1_M1001_g N_VGND_c_481_n 0.00474594f $X=2.62 $Y=0.935 $X2=0 $Y2=0
cc_232 B1 N_VGND_c_481_n 0.0304236f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_233 N_B1_c_298_n N_VGND_c_481_n 0.00291452f $X=2.71 $Y=0.34 $X2=0 $Y2=0
cc_234 B1 N_VGND_c_484_n 0.0227602f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_235 N_B1_c_298_n N_VGND_c_484_n 0.00659434f $X=2.71 $Y=0.34 $X2=0 $Y2=0
cc_236 B1 N_VGND_c_486_n 0.011864f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_237 N_B1_c_298_n N_VGND_c_486_n 0.00886835f $X=2.71 $Y=0.34 $X2=0 $Y2=0
cc_238 N_C1_M1005_g N_VPWR_c_401_n 0.005209f $X=3.045 $Y=2.46 $X2=0 $Y2=0
cc_239 N_C1_M1005_g N_VPWR_c_396_n 0.00987283f $X=3.045 $Y=2.46 $X2=0 $Y2=0
cc_240 N_C1_M1005_g N_A_261_392#_c_442_n 4.88988e-19 $X=3.045 $Y=2.46 $X2=0
+ $Y2=0
cc_241 N_C1_M1005_g N_A_261_392#_c_443_n 0.00234524f $X=3.045 $Y=2.46 $X2=0
+ $Y2=0
cc_242 N_C1_M1003_g N_VGND_c_481_n 0.0170264f $X=3.195 $Y=0.935 $X2=0 $Y2=0
cc_243 N_C1_c_337_n N_VGND_c_481_n 0.0034605f $X=3.195 $Y=1.405 $X2=0 $Y2=0
cc_244 N_C1_c_338_n N_VGND_c_481_n 0.0116775f $X=3.27 $Y=0.34 $X2=0 $Y2=0
cc_245 N_C1_c_340_n N_VGND_c_481_n 0.030194f $X=3.55 $Y=0.34 $X2=0 $Y2=0
cc_246 N_C1_c_338_n N_VGND_c_485_n 0.011998f $X=3.27 $Y=0.34 $X2=0 $Y2=0
cc_247 N_C1_c_340_n N_VGND_c_485_n 0.0215843f $X=3.55 $Y=0.34 $X2=0 $Y2=0
cc_248 N_C1_c_338_n N_VGND_c_486_n 0.00332328f $X=3.27 $Y=0.34 $X2=0 $Y2=0
cc_249 N_C1_c_339_n N_VGND_c_486_n 0.0149884f $X=3.55 $Y=0.34 $X2=0 $Y2=0
cc_250 N_C1_c_340_n N_VGND_c_486_n 0.0110944f $X=3.55 $Y=0.34 $X2=0 $Y2=0
cc_251 X N_VPWR_c_397_n 0.039791f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_252 X N_VPWR_c_396_n 0.0127129f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_253 X N_VPWR_c_403_n 0.0154414f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_254 N_X_c_376_n N_VGND_c_480_n 0.017215f $X=0.52 $Y=0.645 $X2=0 $Y2=0
cc_255 N_X_c_376_n N_VGND_c_482_n 0.00710472f $X=0.52 $Y=0.645 $X2=0 $Y2=0
cc_256 N_X_c_376_n N_VGND_c_486_n 0.00832885f $X=0.52 $Y=0.645 $X2=0 $Y2=0
cc_257 N_VPWR_c_397_n N_A_261_392#_c_439_n 0.00755647f $X=0.875 $Y=2.115 $X2=0
+ $Y2=0
cc_258 N_VPWR_c_397_n N_A_261_392#_c_440_n 0.0330629f $X=0.875 $Y=2.115 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_398_n N_A_261_392#_c_440_n 0.0234237f $X=1.91 $Y=2.455 $X2=0
+ $Y2=0
cc_260 N_VPWR_c_399_n N_A_261_392#_c_440_n 0.0144623f $X=1.805 $Y=3.33 $X2=0
+ $Y2=0
cc_261 N_VPWR_c_396_n N_A_261_392#_c_440_n 0.0118344f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_262 N_VPWR_M1002_d N_A_261_392#_c_441_n 0.00261503f $X=1.755 $Y=1.96 $X2=0
+ $Y2=0
cc_263 N_VPWR_c_398_n N_A_261_392#_c_441_n 0.0200142f $X=1.91 $Y=2.455 $X2=0
+ $Y2=0
cc_264 N_VPWR_c_398_n N_A_261_392#_c_443_n 0.0266656f $X=1.91 $Y=2.455 $X2=0
+ $Y2=0
cc_265 N_VPWR_c_401_n N_A_261_392#_c_443_n 0.0144436f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_266 N_VPWR_c_396_n N_A_261_392#_c_443_n 0.0118287f $X=3.6 $Y=3.33 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__mux2i_1.spice
* Created: Wed Sep  2 12:11:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__mux2i_1.pex.spice"
.subckt sky130_fd_sc_ms__mux2i_1  VNB VPB S A0 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A0	A0
* S	S
* VPB	VPB
* VNB	VNB
MM1007 N_A_114_74#_M1007_d N_S_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.15675 AS=0.15675 PD=1.67 PS=1.67 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1008 N_VGND_M1008_d N_S_M1008_g N_A_225_74#_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.2109 PD=1.16 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1001 A_426_74# N_A_114_74#_M1001_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.0888 AS=0.1554 PD=0.98 PS=1.16 NRD=10.536 NRS=11.34 M=1 R=4.93333
+ SA=75000.8 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A0_M1000_g A_426_74# VNB NLOWVT L=0.15 W=0.74 AD=0.26085
+ AS=0.0888 PD=1.445 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75001.2
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1004 N_A_225_74#_M1004_d N_A1_M1004_g N_Y_M1000_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.26085 PD=2.05 PS=1.445 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_A_114_74#_M1009_d N_S_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=0.84
+ AD=0.2184 AS=0.2268 PD=2.2 PS=2.22 NRD=0 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1002 N_VPWR_M1002_d N_S_M1002_g N_A_223_368#_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2968 PD=1.39 PS=2.77 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1003 N_A_402_368#_M1003_d N_A_114_74#_M1003_g N_VPWR_M1002_d VPB PSHORT L=0.18
+ W=1.12 AD=0.2912 AS=0.1512 PD=2.76 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1005 N_Y_M1005_d N_A0_M1005_g N_A_223_368#_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2968 PD=1.39 PS=2.77 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1006 N_A_402_368#_M1006_d N_A1_M1006_g N_Y_M1005_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3024 AS=0.1512 PD=2.78 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ms__mux2i_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__nor4bb_2.spice
* Created: Fri Aug 28 17:50:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nor4bb_2.pex.spice"
.subckt sky130_fd_sc_ms__nor4bb_2  VNB VPB C_N D_N B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* D_N	D_N
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1019 N_VGND_M1019_d N_C_N_M1019_g N_A_27_392#_M1019_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.180725 AS=0.1824 PD=1.42 PS=1.85 NRD=15.936 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1013 N_A_311_124#_M1013_d N_D_N_M1013_g N_VGND_M1019_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.2496 AS=0.180725 PD=2.06 PS=1.42 NRD=17.808 NRS=42.624 M=1
+ R=4.26667 SA=75000.6 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1009 N_Y_M1009_d N_A_311_124#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.4735 PD=1.02 PS=2.86 NRD=0 NRS=29.184 M=1 R=4.93333 SA=75000.5
+ SB=75004.1 A=0.111 P=1.78 MULT=1
MM1017 N_Y_M1009_d N_A_311_124#_M1017_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2096 PD=1.02 PS=1.405 NRD=0 NRS=37.008 M=1 R=4.93333 SA=75000.9
+ SB=75003.6 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1017_s N_A_27_392#_M1011_g N_Y_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2096 AS=0.1036 PD=1.405 PS=1.02 NRD=37.008 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1018_d N_A_27_392#_M1018_g N_Y_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_B_M1002_g N_VGND_M1018_d VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.5 SB=75002.1
+ A=0.111 P=1.78 MULT=1
MM1016 N_Y_M1002_d N_B_M1016_g N_VGND_M1016_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.30155 PD=1.02 PS=1.555 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.9 SB=75001.6
+ A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1016_s N_A_M1000_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.30155 AS=0.12025 PD=1.555 PS=1.065 NRD=0 NRS=7.296 M=1 R=4.93333
+ SA=75003.9 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_A_M1015_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.12025 PD=2.05 PS=1.065 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.3 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1003 N_VPWR_M1003_d N_C_N_M1003_g N_A_27_392#_M1003_s VPB PSHORT L=0.18 W=1
+ AD=0.57 AS=0.28 PD=2.14 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.5 A=0.18 P=2.36 MULT=1
MM1014 N_A_311_124#_M1014_d N_D_N_M1014_g N_VPWR_M1003_d VPB PSHORT L=0.18 W=1
+ AD=0.28 AS=0.57 PD=2.56 PS=2.14 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.5
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1001 N_Y_M1001_d N_A_311_124#_M1001_g N_A_493_368#_M1001_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1007 N_Y_M1001_d N_A_311_124#_M1007_g N_A_493_368#_M1007_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90000.6 SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1004 N_A_775_368#_M1004_d N_A_27_392#_M1004_g N_A_493_368#_M1007_s VPB PSHORT
+ L=0.18 W=1.12 AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=7.8997 NRS=0 M=1
+ R=6.22222 SA=90001.1 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1005 N_A_775_368#_M1004_d N_A_27_392#_M1005_g N_A_493_368#_M1005_s VPB PSHORT
+ L=0.18 W=1.12 AD=0.1792 AS=0.3136 PD=1.44 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1006 N_A_775_368#_M1006_d N_B_M1006_g N_A_985_368#_M1006_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1010 N_A_775_368#_M1006_d N_B_M1010_g N_A_985_368#_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90000.6 SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1008 N_VPWR_M1008_d N_A_M1008_g N_A_985_368#_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1012 N_VPWR_M1008_d N_A_M1012_g N_A_985_368#_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX20_noxref VNB VPB NWDIODE A=14.0988 P=18.88
*
.include "sky130_fd_sc_ms__nor4bb_2.pxi.spice"
*
.ends
*
*

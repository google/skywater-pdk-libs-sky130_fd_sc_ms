* File: sky130_fd_sc_ms__fa_4.spice
* Created: Wed Sep  2 12:09:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__fa_4.pex.spice"
.subckt sky130_fd_sc_ms__fa_4  VNB VPB B CIN A VPWR SUM COUT VGND
* 
* VGND	VGND
* COUT	COUT
* SUM	SUM
* VPWR	VPWR
* A	A
* CIN	CIN
* B	B
* VPB	VPB
* VNB	VNB
MM1034 N_VGND_M1034_d N_A_M1034_g N_A_27_74#_M1034_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.39435 AS=0.2109 PD=1.87 PS=2.05 NRD=77.496 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75010.1 A=0.111 P=1.78 MULT=1
MM1030 N_A_27_74#_M1030_d N_B_M1030_g N_VGND_M1034_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.39435 PD=1.02 PS=1.87 NRD=0 NRS=77.496 M=1 R=4.93333 SA=75001.3
+ SB=75009 A=0.111 P=1.78 MULT=1
MM1001 N_A_418_74#_M1001_d N_CIN_M1001_g N_A_27_74#_M1030_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75001.7 SB=75008.5 A=0.111 P=1.78 MULT=1
MM1026 A_532_74# N_B_M1026_g N_A_418_74#_M1001_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.1554 PD=1.13 PS=1.16 NRD=22.692 NRS=11.34 M=1 R=4.93333
+ SA=75002.3 SB=75008 A=0.111 P=1.78 MULT=1
MM1035 N_VGND_M1035_d N_A_M1035_g A_532_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1184
+ AS=0.1443 PD=1.06 PS=1.13 NRD=0 NRS=22.692 M=1 R=4.93333 SA=75002.8 SB=75007.4
+ A=0.111 P=1.78 MULT=1
MM1032 N_A_734_74#_M1032_d N_CIN_M1032_g N_VGND_M1035_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1184 PD=1.02 PS=1.06 NRD=0 NRS=6.48 M=1 R=4.93333 SA=75003.3
+ SB=75007 A=0.111 P=1.78 MULT=1
MM1033 N_VGND_M1033_d N_B_M1033_g N_A_734_74#_M1032_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.19035 AS=0.1036 PD=1.37 PS=1.02 NRD=32.784 NRS=0 M=1 R=4.93333 SA=75003.7
+ SB=75006.5 A=0.111 P=1.78 MULT=1
MM1015 N_A_734_74#_M1015_d N_A_M1015_g N_VGND_M1033_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.19035 PD=1.02 PS=1.37 NRD=0 NRS=32.784 M=1 R=4.93333 SA=75004.3
+ SB=75005.9 A=0.111 P=1.78 MULT=1
MM1016 N_A_1024_74#_M1016_d N_A_418_74#_M1016_g N_A_734_74#_M1015_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1961 AS=0.1036 PD=1.27 PS=1.02 NRD=40.536 NRS=0 M=1
+ R=4.93333 SA=75004.8 SB=75005.5 A=0.111 P=1.78 MULT=1
MM1028 A_1160_74# N_CIN_M1028_g N_A_1024_74#_M1016_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.0888 AS=0.1961 PD=0.98 PS=1.27 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75005.4
+ SB=75004.8 A=0.111 P=1.78 MULT=1
MM1039 A_1238_74# N_B_M1039_g A_1160_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1332
+ AS=0.0888 PD=1.1 PS=0.98 NRD=20.268 NRS=10.536 M=1 R=4.93333 SA=75005.8
+ SB=75004.4 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_A_M1002_g A_1238_74# VNB NLOWVT L=0.15 W=0.74 AD=0.19385
+ AS=0.1332 PD=1.41 PS=1.1 NRD=13.776 NRS=20.268 M=1 R=4.93333 SA=75006.3
+ SB=75003.9 A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1002_d N_A_1024_74#_M1022_g N_SUM_M1022_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.19385 AS=0.1036 PD=1.41 PS=1.02 NRD=33.552 NRS=0 M=1 R=4.93333
+ SA=75006.6 SB=75003.5 A=0.111 P=1.78 MULT=1
MM1024 N_VGND_M1024_d N_A_1024_74#_M1024_g N_SUM_M1022_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.19615 AS=0.1036 PD=1.41 PS=1.02 NRD=34.056 NRS=0 M=1 R=4.93333
+ SA=75007 SB=75003.1 A=0.111 P=1.78 MULT=1
MM1036 N_VGND_M1024_d N_A_1024_74#_M1036_g N_SUM_M1036_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.19615 AS=0.1036 PD=1.41 PS=1.02 NRD=34.056 NRS=0 M=1 R=4.93333
+ SA=75007.6 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1038 N_VGND_M1038_d N_A_1024_74#_M1038_g N_SUM_M1036_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.19615 AS=0.1036 PD=1.41 PS=1.02 NRD=34.056 NRS=0 M=1 R=4.93333
+ SA=75008 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1011 N_COUT_M1011_d N_A_418_74#_M1011_g N_VGND_M1038_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.19615 PD=1.02 PS=1.41 NRD=0 NRS=34.056 M=1 R=4.93333
+ SA=75008.6 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1014 N_COUT_M1011_d N_A_418_74#_M1014_g N_VGND_M1014_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75009
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1025 N_COUT_M1025_d N_A_418_74#_M1025_g N_VGND_M1014_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75009.5 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1037 N_COUT_M1025_d N_A_418_74#_M1037_g N_VGND_M1037_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75009.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_A_27_392#_M1003_s VPB PSHORT L=0.18 W=1
+ AD=0.238375 AS=0.28 PD=1.695 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90007.9 A=0.18 P=2.36 MULT=1
MM1017 N_A_27_392#_M1017_d N_B_M1017_g N_VPWR_M1003_d VPB PSHORT L=0.18 W=1
+ AD=0.475662 AS=0.238375 PD=2.02 PS=1.695 NRD=82.8582 NRS=13.7703 M=1 R=5.55556
+ SA=90000.7 SB=90009.1 A=0.18 P=2.36 MULT=1
MM1027 N_A_418_74#_M1027_d N_CIN_M1027_g N_A_27_392#_M1017_d VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.475662 PD=1.27 PS=2.02 NRD=0 NRS=82.8582 M=1 R=5.55556
+ SA=90001.7 SB=90008.1 A=0.18 P=2.36 MULT=1
MM1029 A_538_347# N_B_M1029_g N_A_418_74#_M1027_d VPB PSHORT L=0.18 W=1 AD=0.165
+ AS=0.135 PD=1.33 PS=1.27 NRD=21.6503 NRS=0 M=1 R=5.55556 SA=90002.1 SB=90007.6
+ A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g A_538_347# VPB PSHORT L=0.18 W=1 AD=0.16
+ AS=0.165 PD=1.32 PS=1.33 NRD=0 NRS=21.6503 M=1 R=5.55556 SA=90002.6 SB=90007.1
+ A=0.18 P=2.36 MULT=1
MM1006 N_A_740_347#_M1006_d N_CIN_M1006_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.16 PD=1.27 PS=1.32 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90003.1
+ SB=90006.6 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_B_M1012_g N_A_740_347#_M1006_d VPB PSHORT L=0.18 W=1
+ AD=0.195 AS=0.135 PD=1.39 PS=1.27 NRD=15.7403 NRS=0 M=1 R=5.55556 SA=90003.6
+ SB=90006.2 A=0.18 P=2.36 MULT=1
MM1004 N_A_740_347#_M1004_d N_A_M1004_g N_VPWR_M1012_d VPB PSHORT L=0.18 W=1
+ AD=0.16 AS=0.195 PD=1.32 PS=1.39 NRD=8.8453 NRS=5.8903 M=1 R=5.55556
+ SA=90004.2 SB=90005.6 A=0.18 P=2.36 MULT=1
MM1013 N_A_1024_74#_M1013_d N_A_418_74#_M1013_g N_A_740_347#_M1004_d VPB PSHORT
+ L=0.18 W=1 AD=0.16 AS=0.16 PD=1.32 PS=1.32 NRD=8.8453 NRS=0 M=1 R=5.55556
+ SA=90004.7 SB=90005.1 A=0.18 P=2.36 MULT=1
MM1009 A_1144_347# N_CIN_M1009_g N_A_1024_74#_M1013_d VPB PSHORT L=0.18 W=1
+ AD=0.145 AS=0.16 PD=1.29 PS=1.32 NRD=17.7103 NRS=0 M=1 R=5.55556 SA=90005.2
+ SB=90004.6 A=0.18 P=2.36 MULT=1
MM1031 A_1238_347# N_B_M1031_g A_1144_347# VPB PSHORT L=0.18 W=1 AD=0.18735
+ AS=0.145 PD=1.465 PS=1.29 NRD=26.0631 NRS=17.7103 M=1 R=5.55556 SA=90005.6
+ SB=90004.1 A=0.18 P=2.36 MULT=1
MM1018 N_VPWR_M1018_d N_A_M1018_g A_1238_347# VPB PSHORT L=0.18 W=1 AD=0.188019
+ AS=0.18735 PD=1.40094 PS=1.465 NRD=18.2028 NRS=26.0631 M=1 R=5.55556
+ SA=90005.6 SB=90004 A=0.18 P=2.36 MULT=1
MM1007 N_SUM_M1007_d N_A_1024_74#_M1007_g N_VPWR_M1018_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.210581 PD=1.39 PS=1.56906 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90005.5 SB=90003.5 A=0.2016 P=2.6 MULT=1
MM1008 N_SUM_M1007_d N_A_1024_74#_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90006
+ SB=90003 A=0.2016 P=2.6 MULT=1
MM1010 N_SUM_M1010_d N_A_1024_74#_M1010_g N_VPWR_M1008_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90006.5 SB=90002.5 A=0.2016 P=2.6 MULT=1
MM1020 N_SUM_M1010_d N_A_1024_74#_M1020_g N_VPWR_M1020_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90006.9 SB=90002.1 A=0.2016 P=2.6 MULT=1
MM1000 N_VPWR_M1020_s N_A_418_74#_M1000_g N_COUT_M1000_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90007.4 SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1019 N_VPWR_M1019_d N_A_418_74#_M1019_g N_COUT_M1000_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90007.9 SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1021 N_VPWR_M1019_d N_A_418_74#_M1021_g N_COUT_M1021_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90008.4 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1023 N_VPWR_M1023_d N_A_418_74#_M1023_g N_COUT_M1021_s VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90008.8
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX40_noxref VNB VPB NWDIODE A=21.8696 P=26.77
c_98 VNB 0 3.2512e-19 $X=0 $Y=0
c_188 VPB 0 1.94609e-19 $X=0 $Y=3.085
c_1385 A_538_347# 0 1.16364e-19 $X=2.69 $Y=1.735
*
.include "sky130_fd_sc_ms__fa_4.pxi.spice"
*
.ends
*
*

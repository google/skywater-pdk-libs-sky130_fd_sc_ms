* File: sky130_fd_sc_ms__sdlclkp_2.pex.spice
* Created: Fri Aug 28 18:15:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SDLCLKP_2%SCE 2 5 9 11 12 15 16
r32 15 17 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.455
+ $X2=0.402 $Y2=1.29
r33 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.455 $X2=0.385 $Y2=1.455
r34 12 16 2.58853 $w=6.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.625
+ $X2=0.385 $Y2=1.625
r35 9 17 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.495 $Y=0.835
+ $X2=0.495 $Y2=1.29
r36 5 11 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=0.495 $Y=2.54
+ $X2=0.495 $Y2=1.96
r37 2 11 43.6083 $w=3.65e-07 $l=1.82e-07 $layer=POLY_cond $X=0.402 $Y=1.778
+ $X2=0.402 $Y2=1.96
r38 1 15 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=0.402 $Y=1.472
+ $X2=0.402 $Y2=1.455
r39 1 2 48.3767 $w=3.65e-07 $l=3.06e-07 $layer=POLY_cond $X=0.402 $Y=1.472
+ $X2=0.402 $Y2=1.778
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_2%GATE 3 7 9 12 13
r41 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.795
+ $X2=0.96 $Y2=1.96
r42 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.795
+ $X2=0.96 $Y2=1.63
r43 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.96
+ $Y=1.795 $X2=0.96 $Y2=1.795
r44 9 13 5.68433 $w=5.03e-07 $l=2.4e-07 $layer=LI1_cond $X=1.047 $Y=2.035
+ $X2=1.047 $Y2=1.795
r45 7 14 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=0.925 $Y=0.835
+ $X2=0.925 $Y2=1.63
r46 3 15 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=0.885 $Y=2.54
+ $X2=0.885 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_2%A_318_74# 1 2 9 13 16 17 22 28 30 36
c80 36 0 1.42669e-19 $X=2.94 $Y=1.455
c81 30 0 4.32489e-20 $X=2.855 $Y=1.55
c82 13 0 3.10502e-20 $X=3.35 $Y=0.615
r83 31 36 12.2299 $w=3.35e-07 $l=8.5e-08 $layer=POLY_cond $X=2.855 $Y=1.455
+ $X2=2.94 $Y2=1.455
r84 30 33 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.855 $Y=1.55 $X2=2.855
+ $Y2=1.63
r85 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.855
+ $Y=1.55 $X2=2.855 $Y2=1.55
r86 27 28 10.1887 $w=6.03e-07 $l=1.65e-07 $layer=LI1_cond $X=2.175 $Y=1.847
+ $X2=2.34 $Y2=1.847
r87 20 22 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.73 $Y=0.965
+ $X2=1.895 $Y2=0.965
r88 17 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=1.63
+ $X2=2.855 $Y2=1.63
r89 17 28 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.69 $Y=1.63
+ $X2=2.34 $Y2=1.63
r90 16 27 5.53557 $w=6.03e-07 $l=2.8e-07 $layer=LI1_cond $X=1.895 $Y=1.847
+ $X2=2.175 $Y2=1.847
r91 15 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=1.05
+ $X2=1.895 $Y2=0.965
r92 15 16 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.895 $Y=1.05
+ $X2=1.895 $Y2=1.545
r93 11 36 58.991 $w=3.35e-07 $l=5.24118e-07 $layer=POLY_cond $X=3.35 $Y=1.195
+ $X2=2.94 $Y2=1.455
r94 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.35 $Y=1.195
+ $X2=3.35 $Y2=0.615
r95 7 36 17.2825 $w=1.8e-07 $l=2.6e-07 $layer=POLY_cond $X=2.94 $Y=1.715
+ $X2=2.94 $Y2=1.455
r96 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=2.94 $Y=1.715 $X2=2.94
+ $Y2=2.315
r97 2 27 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.04
+ $Y=1.84 $X2=2.175 $Y2=1.985
r98 1 20 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.59
+ $Y=0.37 $X2=1.73 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_2%A_288_48# 1 2 7 9 10 11 15 16 17 18 19 20
+ 22 25 28 29 30 32 33 34 36 37 38 42 46 49 51 52
c155 42 0 1.44698e-19 $X=5.195 $Y=0.515
c156 38 0 1.9008e-19 $X=4.38 $Y=0.34
c157 37 0 9.22391e-20 $X=4.995 $Y=0.34
c158 28 0 3.10502e-20 $X=2.63 $Y=1.03
r159 51 52 8.46257 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=5.152 $Y=1.885
+ $X2=5.152 $Y2=1.72
r160 49 52 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=5.08 $Y=1.01
+ $X2=5.08 $Y2=1.72
r161 46 48 14.6122 $w=2.63e-07 $l=3.15e-07 $layer=LI1_cond $X=2.315 $Y=1.195
+ $X2=2.63 $Y2=1.195
r162 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.315
+ $Y=1.195 $X2=2.315 $Y2=1.195
r163 40 49 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=5.177 $Y=0.828
+ $X2=5.177 $Y2=1.01
r164 40 42 9.88259 $w=3.63e-07 $l=3.13e-07 $layer=LI1_cond $X=5.177 $Y=0.828
+ $X2=5.177 $Y2=0.515
r165 39 42 2.84164 $w=3.63e-07 $l=9e-08 $layer=LI1_cond $X=5.177 $Y=0.425
+ $X2=5.177 $Y2=0.515
r166 37 39 8.06639 $w=1.7e-07 $l=2.2044e-07 $layer=LI1_cond $X=4.995 $Y=0.34
+ $X2=5.177 $Y2=0.425
r167 37 38 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.995 $Y=0.34
+ $X2=4.38 $Y2=0.34
r168 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.295 $Y=0.425
+ $X2=4.38 $Y2=0.34
r169 35 36 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.295 $Y=0.425
+ $X2=4.295 $Y2=0.905
r170 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.21 $Y=0.99
+ $X2=4.295 $Y2=0.905
r171 33 34 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.21 $Y=0.99
+ $X2=3.7 $Y2=0.99
r172 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.615 $Y=0.905
+ $X2=3.7 $Y2=0.99
r173 31 32 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.615 $Y=0.425
+ $X2=3.615 $Y2=0.905
r174 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.53 $Y=0.34
+ $X2=3.615 $Y2=0.425
r175 29 30 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=3.53 $Y=0.34
+ $X2=2.715 $Y2=0.34
r176 28 48 3.29066 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.63 $Y=1.03
+ $X2=2.63 $Y2=1.195
r177 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.63 $Y=0.425
+ $X2=2.715 $Y2=0.34
r178 27 28 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.63 $Y=0.425
+ $X2=2.63 $Y2=1.03
r179 23 25 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=3.465 $Y=3.075
+ $X2=3.465 $Y2=2.465
r180 20 22 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.825 $Y=0.995
+ $X2=2.825 $Y2=0.645
r181 19 47 39.0383 $w=2.64e-07 $l=2.11849e-07 $layer=POLY_cond $X=2.48 $Y=1.07
+ $X2=2.315 $Y2=1.177
r182 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.75 $Y=1.07
+ $X2=2.825 $Y2=0.995
r183 18 19 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.75 $Y=1.07
+ $X2=2.48 $Y2=1.07
r184 16 23 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.375 $Y=3.15
+ $X2=3.465 $Y2=3.075
r185 16 17 684.543 $w=1.5e-07 $l=1.335e-06 $layer=POLY_cond $X=3.375 $Y=3.15
+ $X2=2.04 $Y2=3.15
r186 13 17 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.95 $Y=3.075
+ $X2=2.04 $Y2=3.15
r187 13 15 316.798 $w=1.8e-07 $l=8.15e-07 $layer=POLY_cond $X=1.95 $Y=3.075
+ $X2=1.95 $Y2=2.26
r188 12 47 66.6402 $w=2.64e-07 $l=4.47236e-07 $layer=POLY_cond $X=1.95 $Y=1.36
+ $X2=2.315 $Y2=1.177
r189 12 15 349.839 $w=1.8e-07 $l=9e-07 $layer=POLY_cond $X=1.95 $Y=1.36 $X2=1.95
+ $Y2=2.26
r190 10 12 25.3451 $w=2.64e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.86 $Y=1.285
+ $X2=1.95 $Y2=1.36
r191 10 11 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.86 $Y=1.285
+ $X2=1.59 $Y2=1.285
r192 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.515 $Y=1.21
+ $X2=1.59 $Y2=1.285
r193 7 9 151.027 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.515 $Y=1.21
+ $X2=1.515 $Y2=0.74
r194 2 51 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.01
+ $Y=1.74 $X2=5.145 $Y2=1.885
r195 1 42 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.05
+ $Y=0.37 $X2=5.195 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_2%A_706_317# 1 2 9 13 17 21 23 26 31 35 38
+ 39 42 43 45 49 54 55 56 60 65
c134 65 0 1.1118e-19 $X=6.565 $Y=1.465
c135 49 0 1.42669e-19 $X=3.695 $Y=1.75
c136 9 0 4.32489e-20 $X=3.74 $Y=0.615
r137 59 60 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=3.74 $Y=1.75
+ $X2=3.855 $Y2=1.75
r138 50 59 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=3.695 $Y=1.75
+ $X2=3.74 $Y2=1.75
r139 49 52 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.695 $Y=1.75
+ $X2=3.695 $Y2=1.84
r140 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.695
+ $Y=1.75 $X2=3.695 $Y2=1.75
r141 46 65 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=6.365 $Y=1.465
+ $X2=6.565 $Y2=1.465
r142 46 62 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.365 $Y=1.465
+ $X2=6.275 $Y2=1.465
r143 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.365
+ $Y=1.465 $X2=6.365 $Y2=1.465
r144 43 45 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=6.005 $Y=1.465
+ $X2=6.365 $Y2=1.465
r145 41 43 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.92 $Y=1.63
+ $X2=6.005 $Y2=1.465
r146 41 42 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.92 $Y=1.63
+ $X2=5.92 $Y2=2.22
r147 40 55 4.39717 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=4.825 $Y=2.305
+ $X2=4.632 $Y2=2.305
r148 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.835 $Y=2.305
+ $X2=5.92 $Y2=2.22
r149 39 40 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=5.835 $Y=2.305
+ $X2=4.825 $Y2=2.305
r150 38 54 3.37808 $w=2.77e-07 $l=1.44375e-07 $layer=LI1_cond $X=4.74 $Y=1.755
+ $X2=4.632 $Y2=1.84
r151 38 56 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.74 $Y=1.755
+ $X2=4.74 $Y2=1.075
r152 33 56 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=4.687 $Y=0.938
+ $X2=4.687 $Y2=1.075
r153 33 35 4.31642 $w=2.73e-07 $l=1.03e-07 $layer=LI1_cond $X=4.687 $Y=0.938
+ $X2=4.687 $Y2=0.835
r154 29 55 2.50573 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.632 $Y=2.39
+ $X2=4.632 $Y2=2.305
r155 29 31 10.9258 $w=3.83e-07 $l=3.65e-07 $layer=LI1_cond $X=4.632 $Y=2.39
+ $X2=4.632 $Y2=2.755
r156 28 54 3.37808 $w=2.77e-07 $l=8.5e-08 $layer=LI1_cond $X=4.632 $Y=1.925
+ $X2=4.632 $Y2=1.84
r157 26 55 2.50573 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.632 $Y=2.22
+ $X2=4.632 $Y2=2.305
r158 26 28 8.83041 $w=3.83e-07 $l=2.95e-07 $layer=LI1_cond $X=4.632 $Y=2.22
+ $X2=4.632 $Y2=1.925
r159 24 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.86 $Y=1.84
+ $X2=3.695 $Y2=1.84
r160 23 54 3.15366 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=4.44 $Y=1.84
+ $X2=4.632 $Y2=1.84
r161 23 24 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.44 $Y=1.84
+ $X2=3.86 $Y2=1.84
r162 19 65 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.565 $Y=1.63
+ $X2=6.565 $Y2=1.465
r163 19 21 287.645 $w=1.8e-07 $l=7.4e-07 $layer=POLY_cond $X=6.565 $Y=1.63
+ $X2=6.565 $Y2=2.37
r164 15 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.275 $Y=1.3
+ $X2=6.275 $Y2=1.465
r165 15 17 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.275 $Y=1.3
+ $X2=6.275 $Y2=0.74
r166 11 60 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.855 $Y=1.915
+ $X2=3.855 $Y2=1.75
r167 11 13 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=3.855 $Y=1.915
+ $X2=3.855 $Y2=2.465
r168 7 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.74 $Y=1.585
+ $X2=3.74 $Y2=1.75
r169 7 9 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=3.74 $Y=1.585
+ $X2=3.74 $Y2=0.615
r170 2 31 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.47
+ $Y=1.78 $X2=4.605 $Y2=2.755
r171 2 28 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.47
+ $Y=1.78 $X2=4.605 $Y2=1.925
r172 1 35 182 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_NDIFF $count=1 $X=4.495
+ $Y=0.405 $X2=4.635 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_2%A_580_74# 1 2 9 13 14 19 22 25 26 28 29 33
+ 36
r84 33 37 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=4.325 $Y=1.42
+ $X2=4.325 $Y2=1.585
r85 33 36 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=4.325 $Y=1.42
+ $X2=4.325 $Y2=1.255
r86 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.32
+ $Y=1.42 $X2=4.32 $Y2=1.42
r87 29 32 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.32 $Y=1.33 $X2=4.32
+ $Y2=1.42
r88 25 26 10.5918 $w=3.58e-07 $l=2.3e-07 $layer=LI1_cond $X=3.18 $Y=2.465
+ $X2=3.18 $Y2=2.235
r89 23 28 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.36 $Y=1.33
+ $X2=3.275 $Y2=1.33
r90 22 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.155 $Y=1.33
+ $X2=4.32 $Y2=1.33
r91 22 23 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=4.155 $Y=1.33
+ $X2=3.36 $Y2=1.33
r92 20 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=1.415
+ $X2=3.275 $Y2=1.33
r93 20 26 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=3.275 $Y=1.415
+ $X2=3.275 $Y2=2.235
r94 19 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.275 $Y=1.245
+ $X2=3.275 $Y2=1.33
r95 18 19 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.275 $Y=0.845
+ $X2=3.275 $Y2=1.245
r96 14 18 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.19 $Y=0.72
+ $X2=3.275 $Y2=0.845
r97 14 16 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=3.19 $Y=0.72
+ $X2=3.05 $Y2=0.72
r98 13 36 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.42 $Y=0.775
+ $X2=4.42 $Y2=1.255
r99 9 37 293.476 $w=1.8e-07 $l=7.55e-07 $layer=POLY_cond $X=4.38 $Y=2.34
+ $X2=4.38 $Y2=1.585
r100 2 25 600 $w=1.7e-07 $l=6.33916e-07 $layer=licon1_PDIFF $count=1 $X=3.03
+ $Y=1.895 $X2=3.165 $Y2=2.465
r101 1 16 182 $w=1.7e-07 $l=3.77624e-07 $layer=licon1_NDIFF $count=1 $X=2.9
+ $Y=0.37 $X2=3.05 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_2%CLK 3 5 7 10 12 14 15 24
c53 15 0 1.1118e-19 $X=5.52 $Y=1.295
c54 12 0 2.36937e-19 $X=5.915 $Y=1.22
r55 23 24 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.9 $Y=1.385
+ $X2=5.915 $Y2=1.385
r56 21 23 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=5.5 $Y=1.385 $X2=5.9
+ $Y2=1.385
r57 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.5
+ $Y=1.385 $X2=5.5 $Y2=1.385
r58 19 21 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.41 $Y=1.385 $X2=5.5
+ $Y2=1.385
r59 17 19 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=5.37 $Y=1.385 $X2=5.41
+ $Y2=1.385
r60 15 22 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.5 $Y=1.295 $X2=5.5
+ $Y2=1.385
r61 12 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.915 $Y=1.22
+ $X2=5.915 $Y2=1.385
r62 12 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.915 $Y=1.22
+ $X2=5.915 $Y2=0.74
r63 8 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.9 $Y=1.55 $X2=5.9
+ $Y2=1.385
r64 8 10 318.742 $w=1.8e-07 $l=8.2e-07 $layer=POLY_cond $X=5.9 $Y=1.55 $X2=5.9
+ $Y2=2.37
r65 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.41 $Y=1.22
+ $X2=5.41 $Y2=1.385
r66 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.41 $Y=1.22 $X2=5.41
+ $Y2=0.74
r67 1 17 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.37 $Y=1.55
+ $X2=5.37 $Y2=1.385
r68 1 3 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=5.37 $Y=1.55 $X2=5.37
+ $Y2=2.16
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_2%A_1198_374# 1 2 9 13 17 21 25 31 33 34 35
+ 36 40 42 44 49
r90 49 50 11.4038 $w=3.17e-07 $l=7.5e-08 $layer=POLY_cond $X=7.6 $Y=1.465
+ $X2=7.675 $Y2=1.465
r91 48 49 53.9779 $w=3.17e-07 $l=3.55e-07 $layer=POLY_cond $X=7.245 $Y=1.465
+ $X2=7.6 $Y2=1.465
r92 47 48 14.4448 $w=3.17e-07 $l=9.5e-08 $layer=POLY_cond $X=7.15 $Y=1.465
+ $X2=7.245 $Y2=1.465
r93 43 47 13.6845 $w=3.17e-07 $l=9e-08 $layer=POLY_cond $X=7.06 $Y=1.465
+ $X2=7.15 $Y2=1.465
r94 42 45 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=7.047 $Y=1.465
+ $X2=7.047 $Y2=1.63
r95 42 44 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=7.047 $Y=1.465
+ $X2=7.047 $Y2=1.3
r96 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.06
+ $Y=1.465 $X2=7.06 $Y2=1.465
r97 40 45 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.955 $Y=1.8
+ $X2=6.955 $Y2=1.63
r98 37 44 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.955 $Y=1.13
+ $X2=6.955 $Y2=1.3
r99 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.87 $Y=1.045
+ $X2=6.955 $Y2=1.13
r100 35 36 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.87 $Y=1.045
+ $X2=6.655 $Y2=1.045
r101 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.87 $Y=1.885
+ $X2=6.955 $Y2=1.8
r102 33 34 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.87 $Y=1.885
+ $X2=6.505 $Y2=1.885
r103 29 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.49 $Y=0.96
+ $X2=6.655 $Y2=1.045
r104 29 31 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=6.49 $Y=0.96
+ $X2=6.49 $Y2=0.515
r105 25 27 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=6.34 $Y=2.015
+ $X2=6.34 $Y2=2.725
r106 23 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.34 $Y=1.97
+ $X2=6.505 $Y2=1.885
r107 23 25 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=6.34 $Y=1.97
+ $X2=6.34 $Y2=2.015
r108 19 50 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.675 $Y=1.3
+ $X2=7.675 $Y2=1.465
r109 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.675 $Y=1.3
+ $X2=7.675 $Y2=0.74
r110 15 49 15.9969 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.6 $Y=1.63
+ $X2=7.6 $Y2=1.465
r111 15 17 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=7.6 $Y=1.63 $X2=7.6
+ $Y2=2.4
r112 11 48 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.245 $Y=1.3
+ $X2=7.245 $Y2=1.465
r113 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.245 $Y=1.3
+ $X2=7.245 $Y2=0.74
r114 7 47 15.9969 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.15 $Y=1.63
+ $X2=7.15 $Y2=1.465
r115 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=7.15 $Y=1.63 $X2=7.15
+ $Y2=2.4
r116 2 27 400 $w=1.7e-07 $l=1.01502e-06 $layer=licon1_PDIFF $count=1 $X=5.99
+ $Y=1.87 $X2=6.34 $Y2=2.725
r117 2 25 400 $w=1.7e-07 $l=4.16233e-07 $layer=licon1_PDIFF $count=1 $X=5.99
+ $Y=1.87 $X2=6.34 $Y2=2.015
r118 1 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.35
+ $Y=0.37 $X2=6.49 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_2%VPWR 1 2 3 4 5 6 19 21 25 29 35 39 43 45
+ 50 51 52 54 59 67 76 84 87 90 94
r92 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r93 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r94 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r95 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r96 79 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r97 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r98 76 93 3.94754 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=7.74 $Y=3.33 $X2=7.95
+ $Y2=3.33
r99 76 78 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=7.74 $Y=3.33 $X2=7.44
+ $Y2=3.33
r100 75 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r101 75 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=5.52 $Y2=3.33
r102 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r103 72 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.84 $Y=3.33
+ $X2=5.675 $Y2=3.33
r104 72 74 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.84 $Y=3.33
+ $X2=6.48 $Y2=3.33
r105 71 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r106 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r107 68 87 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.24 $Y=3.33
+ $X2=4.115 $Y2=3.33
r108 68 70 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.24 $Y=3.33
+ $X2=4.56 $Y2=3.33
r109 67 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.51 $Y=3.33
+ $X2=5.675 $Y2=3.33
r110 67 70 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=5.51 $Y=3.33
+ $X2=4.56 $Y2=3.33
r111 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r112 63 66 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r113 63 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r114 62 65 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r115 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r116 60 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=1.65 $Y2=3.33
r117 60 62 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=2.16 $Y2=3.33
r118 59 87 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.99 $Y=3.33
+ $X2=4.115 $Y2=3.33
r119 59 65 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.99 $Y=3.33
+ $X2=3.6 $Y2=3.33
r120 58 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r121 58 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r122 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r123 55 81 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.217 $Y2=3.33
r124 55 57 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=1.2 $Y2=3.33
r125 54 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.65 $Y2=3.33
r126 54 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.2 $Y2=3.33
r127 52 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r128 52 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r129 52 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r130 50 74 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.71 $Y=3.33
+ $X2=6.48 $Y2=3.33
r131 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.71 $Y=3.33
+ $X2=6.875 $Y2=3.33
r132 49 78 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=7.04 $Y=3.33 $X2=7.44
+ $Y2=3.33
r133 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.04 $Y=3.33
+ $X2=6.875 $Y2=3.33
r134 45 48 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=7.865 $Y=1.985
+ $X2=7.865 $Y2=2.815
r135 43 93 3.19563 $w=2.5e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.865 $Y=3.245
+ $X2=7.95 $Y2=3.33
r136 43 48 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.865 $Y=3.245
+ $X2=7.865 $Y2=2.815
r137 39 42 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=6.875 $Y=2.305
+ $X2=6.875 $Y2=2.815
r138 37 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.875 $Y=3.245
+ $X2=6.875 $Y2=3.33
r139 37 42 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.875 $Y=3.245
+ $X2=6.875 $Y2=2.815
r140 33 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.675 $Y=3.245
+ $X2=5.675 $Y2=3.33
r141 33 35 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=5.675 $Y=3.245
+ $X2=5.675 $Y2=2.725
r142 29 32 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=4.115 $Y=2.26
+ $X2=4.115 $Y2=2.755
r143 27 87 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.115 $Y=3.245
+ $X2=4.115 $Y2=3.33
r144 27 32 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=4.115 $Y=3.245
+ $X2=4.115 $Y2=2.755
r145 23 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.65 $Y=3.245
+ $X2=1.65 $Y2=3.33
r146 23 25 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.65 $Y=3.245
+ $X2=1.65 $Y2=2.825
r147 19 81 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.217 $Y2=3.33
r148 19 21 33.1764 $w=3.28e-07 $l=9.5e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.27 $Y2=2.295
r149 6 48 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.69
+ $Y=1.84 $X2=7.825 $Y2=2.815
r150 6 45 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.69
+ $Y=1.84 $X2=7.825 $Y2=1.985
r151 5 42 600 $w=1.7e-07 $l=1.04925e-06 $layer=licon1_PDIFF $count=1 $X=6.655
+ $Y=1.87 $X2=6.875 $Y2=2.815
r152 5 39 600 $w=1.7e-07 $l=5.33784e-07 $layer=licon1_PDIFF $count=1 $X=6.655
+ $Y=1.87 $X2=6.875 $Y2=2.305
r153 4 35 600 $w=1.7e-07 $l=1.0872e-06 $layer=licon1_PDIFF $count=1 $X=5.46
+ $Y=1.74 $X2=5.675 $Y2=2.725
r154 3 32 600 $w=1.7e-07 $l=5.95819e-07 $layer=licon1_PDIFF $count=1 $X=3.945
+ $Y=2.255 $X2=4.155 $Y2=2.755
r155 3 29 600 $w=1.7e-07 $l=2.12485e-07 $layer=licon1_PDIFF $count=1 $X=3.945
+ $Y=2.255 $X2=4.155 $Y2=2.26
r156 2 25 600 $w=1.7e-07 $l=1.05033e-06 $layer=licon1_PDIFF $count=1 $X=1.515
+ $Y=1.84 $X2=1.65 $Y2=2.825
r157 1 21 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.27 $Y2=2.295
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_2%A_114_112# 1 2 3 4 14 16 17 18 19 23 26 27
+ 31 35 36 38
r98 38 40 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=2.25 $Y=0.53
+ $X2=2.25 $Y2=0.625
r99 29 31 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=2.675 $Y=2.32
+ $X2=2.675 $Y2=2.05
r100 28 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=2.405
+ $X2=1.555 $Y2=2.405
r101 27 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.55 $Y=2.405
+ $X2=2.675 $Y2=2.32
r102 27 28 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=2.55 $Y=2.405
+ $X2=1.64 $Y2=2.405
r103 26 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.555 $Y=2.32
+ $X2=1.555 $Y2=2.405
r104 25 26 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=1.555 $Y=1.39
+ $X2=1.555 $Y2=2.32
r105 24 35 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.275 $Y=2.405
+ $X2=1.11 $Y2=2.405
r106 23 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.47 $Y=2.405
+ $X2=1.555 $Y2=2.405
r107 23 24 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.47 $Y=2.405
+ $X2=1.275 $Y2=2.405
r108 20 33 2.70854 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.89 $Y=1.305
+ $X2=0.72 $Y2=1.305
r109 19 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.47 $Y=1.305
+ $X2=1.555 $Y2=1.39
r110 19 20 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=1.47 $Y=1.305
+ $X2=0.89 $Y2=1.305
r111 17 40 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.125 $Y=0.625
+ $X2=2.25 $Y2=0.625
r112 17 18 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=2.125 $Y=0.625
+ $X2=0.89 $Y2=0.625
r113 14 33 13.8085 $w=3.45e-07 $l=3.58497e-07 $layer=LI1_cond $X=0.717 $Y=0.948
+ $X2=0.72 $Y2=1.305
r114 14 16 3.94169 $w=3.43e-07 $l=1.18e-07 $layer=LI1_cond $X=0.717 $Y=0.948
+ $X2=0.717 $Y2=0.83
r115 13 18 7.89393 $w=1.7e-07 $l=2.11268e-07 $layer=LI1_cond $X=0.717 $Y=0.71
+ $X2=0.89 $Y2=0.625
r116 13 16 4.0085 $w=3.43e-07 $l=1.2e-07 $layer=LI1_cond $X=0.717 $Y=0.71
+ $X2=0.717 $Y2=0.83
r117 4 31 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=2.58
+ $Y=1.895 $X2=2.715 $Y2=2.05
r118 3 35 300 $w=1.7e-07 $l=3.45977e-07 $layer=licon1_PDIFF $count=2 $X=0.975
+ $Y=2.12 $X2=1.11 $Y2=2.405
r119 2 38 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=2.145
+ $Y=0.37 $X2=2.29 $Y2=0.53
r120 1 16 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.56 $X2=0.71 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_2%GCLK 1 2 9 13 14 15 16 23 32
r37 21 23 1.2336 $w=3.53e-07 $l=3.8e-08 $layer=LI1_cond $X=7.387 $Y=1.997
+ $X2=7.387 $Y2=2.035
r38 15 16 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=7.387 $Y=2.405
+ $X2=7.387 $Y2=2.775
r39 14 21 0.779116 $w=3.53e-07 $l=2.4e-08 $layer=LI1_cond $X=7.387 $Y=1.973
+ $X2=7.387 $Y2=1.997
r40 14 32 8.1095 $w=3.53e-07 $l=1.53e-07 $layer=LI1_cond $X=7.387 $Y=1.973
+ $X2=7.387 $Y2=1.82
r41 14 15 11.2647 $w=3.53e-07 $l=3.47e-07 $layer=LI1_cond $X=7.387 $Y=2.058
+ $X2=7.387 $Y2=2.405
r42 14 23 0.746653 $w=3.53e-07 $l=2.3e-08 $layer=LI1_cond $X=7.387 $Y=2.058
+ $X2=7.387 $Y2=2.035
r43 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.48 $Y=1.13 $X2=7.48
+ $Y2=1.82
r44 7 13 7.30505 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.46 $Y=0.965
+ $X2=7.46 $Y2=1.13
r45 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=7.46 $Y=0.965 $X2=7.46
+ $Y2=0.515
r46 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.24
+ $Y=1.84 $X2=7.375 $Y2=1.985
r47 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.24
+ $Y=1.84 $X2=7.375 $Y2=2.815
r48 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.32
+ $Y=0.37 $X2=7.46 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDLCLKP_2%VGND 1 2 3 4 5 6 19 21 25 29 33 35 37 40
+ 41 43 44 45 47 65 69 79 85 89
c93 3 0 1.9008e-19 $X=3.815 $Y=0.405
r94 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r95 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r96 79 82 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.22 $Y=0 $X2=1.22
+ $Y2=0.285
r97 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r98 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r99 73 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r100 73 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r101 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r102 70 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.115 $Y=0 $X2=6.99
+ $Y2=0
r103 70 72 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.115 $Y=0
+ $X2=7.44 $Y2=0
r104 69 88 4.02656 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=7.805 $Y=0
+ $X2=7.982 $Y2=0
r105 69 72 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.805 $Y=0
+ $X2=7.44 $Y2=0
r106 68 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r107 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r108 65 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.865 $Y=0 $X2=6.99
+ $Y2=0
r109 65 67 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.865 $Y=0
+ $X2=6.48 $Y2=0
r110 64 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r111 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r112 60 63 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.52
+ $Y2=0
r113 57 58 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r114 55 58 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=3.6
+ $Y2=0
r115 55 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r116 54 57 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.6
+ $Y2=0
r117 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r118 52 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.22
+ $Y2=0
r119 52 54 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.68
+ $Y2=0
r120 51 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r121 51 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r122 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r123 48 75 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r124 48 50 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.72 $Y2=0
r125 47 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.22
+ $Y2=0
r126 47 50 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=0.72 $Y2=0
r127 45 64 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=5.52 $Y2=0
r128 45 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r129 45 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r130 43 63 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=5.53 $Y=0 $X2=5.52
+ $Y2=0
r131 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.53 $Y=0 $X2=5.695
+ $Y2=0
r132 42 67 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=5.86 $Y=0 $X2=6.48
+ $Y2=0
r133 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.86 $Y=0 $X2=5.695
+ $Y2=0
r134 40 57 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.87 $Y=0 $X2=3.6
+ $Y2=0
r135 40 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.87 $Y=0 $X2=3.955
+ $Y2=0
r136 39 60 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=4.04 $Y=0 $X2=4.08
+ $Y2=0
r137 39 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=0 $X2=3.955
+ $Y2=0
r138 35 88 3.1166 $w=2.5e-07 $l=1.07912e-07 $layer=LI1_cond $X=7.93 $Y=0.085
+ $X2=7.982 $Y2=0
r139 35 37 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.93 $Y=0.085
+ $X2=7.93 $Y2=0.515
r140 31 85 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.99 $Y=0.085
+ $X2=6.99 $Y2=0
r141 31 33 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=6.99 $Y=0.085
+ $X2=6.99 $Y2=0.57
r142 27 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.695 $Y=0.085
+ $X2=5.695 $Y2=0
r143 27 29 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.695 $Y=0.085
+ $X2=5.695 $Y2=0.515
r144 23 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.955 $Y=0.085
+ $X2=3.955 $Y2=0
r145 23 25 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.955 $Y=0.085
+ $X2=3.955 $Y2=0.56
r146 19 75 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r147 19 21 34.3428 $w=2.48e-07 $l=7.45e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.83
r148 6 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.75
+ $Y=0.37 $X2=7.89 $Y2=0.515
r149 5 33 182 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_NDIFF $count=1 $X=6.895
+ $Y=0.37 $X2=7.03 $Y2=0.57
r150 4 29 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=5.485
+ $Y=0.37 $X2=5.695 $Y2=0.515
r151 3 25 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=3.815
+ $Y=0.405 $X2=3.955 $Y2=0.56
r152 2 82 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.56 $X2=1.22 $Y2=0.285
r153 1 21 182 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.28 $Y2=0.83
.ends


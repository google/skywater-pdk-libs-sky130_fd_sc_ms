* File: sky130_fd_sc_ms__nand3b_1.spice
* Created: Fri Aug 28 17:43:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nand3b_1.pex.spice"
.subckt sky130_fd_sc_ms__nand3b_1  VNB VPB A_N C B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* C	C
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_N_M1004_g N_A_27_116#_M1004_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.191114 AS=0.15675 PD=1.16395 PS=1.67 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75002.1 A=0.0825 P=1.4 MULT=1
MM1006 A_269_78# N_C_M1006_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.257136 PD=0.98 PS=1.56605 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.9
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1007 A_347_78# N_B_M1007_g A_269_78# VNB NLOWVT L=0.15 W=0.74 AD=0.1443
+ AS=0.0888 PD=1.13 PS=0.98 NRD=22.692 NRS=10.536 M=1 R=4.93333 SA=75001.2
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_A_27_116#_M1002_g A_347_78# VNB NLOWVT L=0.15 W=0.74
+ AD=0.3404 AS=0.1443 PD=2.4 PS=1.13 NRD=14.184 NRS=22.692 M=1 R=4.93333
+ SA=75001.8 SB=75000.4 A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_A_N_M1005_g N_A_27_116#_M1005_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1854 AS=0.2352 PD=1.30714 PS=2.24 NRD=18.7544 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90001.8 A=0.1512 P=2.04 MULT=1
MM1001 N_Y_M1001_d N_C_M1001_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.2472 PD=1.39 PS=1.74286 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.6
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1003 N_VPWR_M1003_d N_B_M1003_g N_Y_M1001_d VPB PSHORT L=0.18 W=1.12 AD=0.2072
+ AS=0.1512 PD=1.49 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90001.1 SB=90000.7
+ A=0.2016 P=2.6 MULT=1
MM1000 N_Y_M1000_d N_A_27_116#_M1000_g N_VPWR_M1003_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.2072 PD=2.8 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ms__nand3b_1.pxi.spice"
*
.ends
*
*

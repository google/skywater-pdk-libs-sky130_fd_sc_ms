* File: sky130_fd_sc_ms__mux2i_4.spice
* Created: Fri Aug 28 17:40:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__mux2i_4.pex.spice"
.subckt sky130_fd_sc_ms__mux2i_4  VNB VPB A1 A0 S Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* S	S
* A0	A0
* A1	A1
* VPB	VPB
* VNB	VNB
MM1000 N_Y_M1000_d N_A1_M1000_g N_A_114_85#_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1005 N_Y_M1005_d N_A1_M1005_g N_A_114_85#_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1022 N_Y_M1005_d N_A1_M1022_g N_A_114_85#_M1022_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.13505 PD=1.02 PS=1.105 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1023 N_Y_M1023_d N_A1_M1023_g N_A_114_85#_M1022_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.13505 PD=1.02 PS=1.105 NRD=0 NRS=13.776 M=1 R=4.93333
+ SA=75001.6 SB=75002 A=0.111 P=1.78 MULT=1
MM1007 N_A_475_85#_M1007_d N_A0_M1007_g N_Y_M1023_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1030 N_A_475_85#_M1007_d N_A0_M1030_g N_Y_M1030_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.12025 PD=1.09 PS=1.065 NRD=0 NRS=3.24 M=1 R=4.93333 SA=75002.5
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1031 N_A_475_85#_M1031_d N_A0_M1031_g N_Y_M1030_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.12025 PD=1.02 PS=1.065 NRD=0 NRS=4.044 M=1 R=4.93333 SA=75003
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1034 N_A_475_85#_M1031_d N_A0_M1034_g N_Y_M1034_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.4
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1013 N_A_475_85#_M1013_d N_A_1030_268#_M1013_g N_VGND_M1013_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1036 AS=0.36 PD=1.02 PS=2.83 NRD=0 NRS=69.96 M=1 R=4.93333
+ SA=75000.3 SB=75003.9 A=0.111 P=1.78 MULT=1
MM1014 N_A_475_85#_M1013_d N_A_1030_268#_M1014_g N_VGND_M1014_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1036 AS=0.20315 PD=1.02 PS=1.49 NRD=0 NRS=35.592 M=1
+ R=4.93333 SA=75000.7 SB=75003.5 A=0.111 P=1.78 MULT=1
MM1026 N_A_475_85#_M1026_d N_A_1030_268#_M1026_g N_VGND_M1014_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1036 AS=0.20315 PD=1.02 PS=1.49 NRD=0 NRS=35.592 M=1
+ R=4.93333 SA=75001.2 SB=75003.3 A=0.111 P=1.78 MULT=1
MM1029 N_A_475_85#_M1026_d N_A_1030_268#_M1029_g N_VGND_M1029_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1036 AS=0.19615 PD=1.02 PS=1.41 NRD=0 NRS=34.056 M=1
+ R=4.93333 SA=75001.6 SB=75002.9 A=0.111 P=1.78 MULT=1
MM1010 N_A_114_85#_M1010_d N_S_M1010_g N_VGND_M1029_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.19615 PD=1.02 PS=1.41 NRD=0 NRS=34.056 M=1 R=4.93333 SA=75002.2
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1017 N_A_114_85#_M1010_d N_S_M1017_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1887 PD=1.02 PS=1.25 NRD=0 NRS=18.648 M=1 R=4.93333 SA=75002.6
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1025 N_A_114_85#_M1025_d N_S_M1025_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1887 PD=1.02 PS=1.25 NRD=0 NRS=18.648 M=1 R=4.93333 SA=75003.3
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1028 N_A_114_85#_M1025_d N_S_M1028_g N_VGND_M1028_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003.7
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1024 N_A_1030_268#_M1024_d N_S_M1024_g N_VGND_M1028_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.1295 PD=2.19 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75004.2
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1008 N_A_119_368#_M1008_d N_A1_M1008_g N_Y_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003.5 A=0.2016 P=2.6 MULT=1
MM1009 N_A_119_368#_M1008_d N_A1_M1009_g N_Y_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90003.1 A=0.2016 P=2.6 MULT=1
MM1011 N_A_119_368#_M1011_d N_A1_M1011_g N_Y_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90002.6 A=0.2016 P=2.6 MULT=1
MM1015 N_A_119_368#_M1011_d N_A1_M1015_g N_Y_M1015_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1568 PD=1.39 PS=1.4 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90002.2 A=0.2016 P=2.6 MULT=1
MM1001 N_A_481_368#_M1001_d N_A0_M1001_g N_Y_M1015_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1736 AS=0.1568 PD=1.43 PS=1.4 NRD=6.1464 NRS=0.8668 M=1 R=6.22222
+ SA=90002 SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1016 N_A_481_368#_M1001_d N_A0_M1016_g N_Y_M1016_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1736 AS=0.1792 PD=1.43 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.5
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1018 N_A_481_368#_M1018_d N_A0_M1018_g N_Y_M1016_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90003
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1019 N_A_481_368#_M1018_d N_A0_M1019_g N_Y_M1019_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.3696 PD=1.44 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1002 N_VPWR_M1002_d N_A_1030_268#_M1002_g N_A_119_368#_M1002_s VPB PSHORT
+ L=0.18 W=1.12 AD=0.7336 AS=0.1512 PD=3.55 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90004.3 A=0.2016 P=2.6 MULT=1
MM1012 N_VPWR_M1012_d N_A_1030_268#_M1012_g N_A_119_368#_M1002_s VPB PSHORT
+ L=0.18 W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001 SB=90003.8 A=0.2016 P=2.6 MULT=1
MM1020 N_VPWR_M1012_d N_A_1030_268#_M1020_g N_A_119_368#_M1020_s VPB PSHORT
+ L=0.18 W=1.12 AD=0.1512 AS=0.196 PD=1.39 PS=1.47 NRD=0 NRS=1.7533 M=1
+ R=6.22222 SA=90001.5 SB=90003.4 A=0.2016 P=2.6 MULT=1
MM1021 N_VPWR_M1021_d N_A_1030_268#_M1021_g N_A_119_368#_M1020_s VPB PSHORT
+ L=0.18 W=1.12 AD=0.1792 AS=0.196 PD=1.44 PS=1.47 NRD=0 NRS=10.5395 M=1
+ R=6.22222 SA=90002 SB=90002.8 A=0.2016 P=2.6 MULT=1
MM1003 N_A_481_368#_M1003_d N_S_M1003_g N_VPWR_M1021_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.5
+ SB=90002.3 A=0.2016 P=2.6 MULT=1
MM1004 N_A_481_368#_M1003_d N_S_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.9
+ SB=90001.9 A=0.2016 P=2.6 MULT=1
MM1006 N_A_481_368#_M1006_d N_S_M1006_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003.5
+ SB=90001.3 A=0.2016 P=2.6 MULT=1
MM1032 N_A_481_368#_M1006_d N_S_M1032_g N_VPWR_M1032_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.196 PD=1.39 PS=1.65143 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.9
+ SB=90000.9 A=0.2016 P=2.6 MULT=1
MM1027 N_A_1030_268#_M1027_d N_S_M1027_g N_VPWR_M1032_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.147 PD=1.11 PS=1.23857 NRD=0 NRS=11.7215 M=1 R=4.66667
+ SA=90004.4 SB=90000.6 A=0.1512 P=2.04 MULT=1
MM1033 N_A_1030_268#_M1027_d N_S_M1033_g N_VPWR_M1033_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.2352 PD=1.11 PS=2.24 NRD=0 NRS=0 M=1 R=4.66667 SA=90004.9
+ SB=90000.2 A=0.1512 P=2.04 MULT=1
DX35_noxref VNB VPB NWDIODE A=19.4556 P=24.64
*
.include "sky130_fd_sc_ms__mux2i_4.pxi.spice"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_245_94# B1 a_456_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X1 a_245_94# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 a_465_392# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X3 X a_83_264# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VPWR A1 a_267_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X5 VPWR C1 a_83_264# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X6 VGND A1 a_245_94# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X7 a_267_392# A2 a_83_264# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X8 X a_83_264# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X9 a_83_264# B2 a_465_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X10 a_456_74# B2 a_245_94# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X11 a_456_74# C1 a_83_264# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends

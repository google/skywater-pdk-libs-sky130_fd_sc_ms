* File: sky130_fd_sc_ms__a2111o_1.spice
* Created: Fri Aug 28 16:55:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a2111o_1.pex.spice"
.subckt sky130_fd_sc_ms__a2111o_1  VNB VPB A1 A2 B1 C1 D1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D1	D1
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1002 A_168_136# N_A1_M1002_g N_A_85_136#_M1002_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1696 PD=0.85 PS=1.81 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g A_168_136# VNB NLOWVT L=0.15 W=0.64 AD=0.1248
+ AS=0.0672 PD=1.03 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667 SA=75000.6 SB=75001.8
+ A=0.096 P=1.58 MULT=1
MM1006 N_A_85_136#_M1006_d N_B1_M1006_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1248 PD=0.92 PS=1.03 NRD=0 NRS=20.616 M=1 R=4.26667 SA=75001.1
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1007 N_VGND_M1007_d N_C1_M1007_g N_A_85_136#_M1006_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1504 AS=0.0896 PD=1.11 PS=0.92 NRD=35.616 NRS=0 M=1 R=4.26667 SA=75001.5
+ SB=75000.8 A=0.096 P=1.58 MULT=1
MM1003 N_A_85_136#_M1003_d N_D1_M1003_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1696 AS=0.1504 PD=1.81 PS=1.11 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.1
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 N_X_M1008_d N_A_85_136#_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1961 PD=2.01 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_VPWR_M1010_d N_A1_M1010_g N_A_80_392#_M1010_s VPB PSHORT L=0.18 W=1
+ AD=0.155 AS=0.26 PD=1.31 PS=2.52 NRD=2.9353 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.9 A=0.18 P=2.36 MULT=1
MM1000 N_A_80_392#_M1000_d N_A2_M1000_g N_VPWR_M1010_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.155 PD=1.27 PS=1.31 NRD=0 NRS=2.9353 M=1 R=5.55556 SA=90000.7
+ SB=90001.4 A=0.18 P=2.36 MULT=1
MM1001 A_356_392# N_B1_M1001_g N_A_80_392#_M1000_d VPB PSHORT L=0.18 W=1
+ AD=0.105 AS=0.135 PD=1.21 PS=1.27 NRD=9.8303 NRS=0 M=1 R=5.55556 SA=90001.1
+ SB=90000.9 A=0.18 P=2.36 MULT=1
MM1009 A_434_392# N_C1_M1009_g A_356_392# VPB PSHORT L=0.18 W=1 AD=0.105
+ AS=0.105 PD=1.21 PS=1.21 NRD=9.8303 NRS=9.8303 M=1 R=5.55556 SA=90001.5
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1004 N_A_85_136#_M1004_d N_D1_M1004_g A_434_392# VPB PSHORT L=0.18 W=1 AD=0.26
+ AS=0.105 PD=2.52 PS=1.21 NRD=0 NRS=9.8303 M=1 R=5.55556 SA=90001.9 SB=90000.2
+ A=0.18 P=2.36 MULT=1
MM1011 N_X_M1011_d N_A_85_136#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2912 AS=0.2912 PD=2.76 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__a2111o_1.pxi.spice"
*
.ends
*
*

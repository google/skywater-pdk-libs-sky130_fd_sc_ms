* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
X0 VGND B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_345_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X2 a_159_368# C1 a_237_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 Y C1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 Y A1 a_461_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 VPWR A2 a_345_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X6 a_461_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_237_368# B1 a_345_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 Y D1 a_159_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X9 VGND D1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

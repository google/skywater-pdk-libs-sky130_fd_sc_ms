* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
X0 a_2022_94# a_1356_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X1 Q a_2022_94# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X2 a_1489_118# a_1566_92# a_1596_118# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 a_719_456# a_767_384# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X4 VGND a_2022_94# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 VPWR SET_B a_1356_74# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X6 a_27_74# a_225_74# a_612_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X7 VPWR a_1356_74# a_1566_92# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X8 a_1356_74# a_225_74# a_1489_118# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X9 a_1356_74# a_398_74# a_1524_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X10 a_781_74# a_767_384# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X11 Q a_2022_94# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 a_1057_118# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X13 VPWR a_2022_94# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X14 a_1596_118# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X15 VPWR a_225_74# a_398_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X16 VPWR a_612_74# a_1269_341# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X17 a_27_74# D VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X18 a_612_74# a_398_74# a_781_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X19 VGND a_225_74# a_398_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 a_27_74# a_398_74# a_612_74# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X21 a_1269_341# a_225_74# a_1356_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X22 VPWR a_612_74# a_767_384# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X23 a_225_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 a_767_384# a_612_74# a_1057_118# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X25 a_1524_508# a_1566_92# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X26 a_767_384# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X27 a_1278_74# a_398_74# a_1356_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X28 a_612_74# a_225_74# a_719_456# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X29 a_27_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X30 VGND a_612_74# a_1278_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X31 a_225_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X32 VGND a_1356_74# a_1566_92# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X33 a_2022_94# a_1356_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends

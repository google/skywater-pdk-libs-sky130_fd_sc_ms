* File: sky130_fd_sc_ms__bufinv_16.pxi.spice
* Created: Fri Aug 28 17:16:35 2020
* 
x_PM_SKY130_FD_SC_MS__BUFINV_16%A N_A_M1000_g N_A_M1001_g N_A_M1002_g
+ N_A_M1035_g N_A_M1005_g N_A_M1047_g A A A N_A_c_234_n N_A_c_235_n
+ PM_SKY130_FD_SC_MS__BUFINV_16%A
x_PM_SKY130_FD_SC_MS__BUFINV_16%A_27_74# N_A_27_74#_M1000_d N_A_27_74#_M1035_d
+ N_A_27_74#_M1001_s N_A_27_74#_M1002_s N_A_27_74#_M1011_g N_A_27_74#_M1009_g
+ N_A_27_74#_M1015_g N_A_27_74#_M1016_g N_A_27_74#_M1018_g N_A_27_74#_M1019_g
+ N_A_27_74#_M1026_g N_A_27_74#_M1025_g N_A_27_74#_M1048_g N_A_27_74#_M1029_g
+ N_A_27_74#_c_308_n N_A_27_74#_M1049_g N_A_27_74#_M1033_g N_A_27_74#_c_311_n
+ N_A_27_74#_c_312_n N_A_27_74#_c_328_n N_A_27_74#_c_329_n N_A_27_74#_c_313_n
+ N_A_27_74#_c_314_n N_A_27_74#_c_344_n N_A_27_74#_c_330_n N_A_27_74#_c_315_n
+ N_A_27_74#_c_316_n N_A_27_74#_c_356_n N_A_27_74#_c_317_n N_A_27_74#_c_318_n
+ N_A_27_74#_c_359_n N_A_27_74#_c_319_n N_A_27_74#_c_320_n N_A_27_74#_c_321_n
+ PM_SKY130_FD_SC_MS__BUFINV_16%A_27_74#
x_PM_SKY130_FD_SC_MS__BUFINV_16%A_384_74# N_A_384_74#_M1011_d
+ N_A_384_74#_M1018_d N_A_384_74#_M1048_d N_A_384_74#_M1009_d
+ N_A_384_74#_M1019_d N_A_384_74#_M1029_d N_A_384_74#_M1003_g
+ N_A_384_74#_M1004_g N_A_384_74#_M1007_g N_A_384_74#_M1006_g
+ N_A_384_74#_M1013_g N_A_384_74#_M1008_g N_A_384_74#_M1021_g
+ N_A_384_74#_M1010_g N_A_384_74#_M1022_g N_A_384_74#_M1012_g
+ N_A_384_74#_M1023_g N_A_384_74#_M1014_g N_A_384_74#_M1017_g
+ N_A_384_74#_M1027_g N_A_384_74#_M1028_g N_A_384_74#_M1020_g
+ N_A_384_74#_M1024_g N_A_384_74#_M1032_g N_A_384_74#_M1030_g
+ N_A_384_74#_M1036_g N_A_384_74#_M1031_g N_A_384_74#_M1038_g
+ N_A_384_74#_M1034_g N_A_384_74#_M1039_g N_A_384_74#_M1037_g
+ N_A_384_74#_M1041_g N_A_384_74#_M1042_g N_A_384_74#_M1040_g
+ N_A_384_74#_M1043_g N_A_384_74#_M1044_g N_A_384_74#_M1046_g
+ N_A_384_74#_M1045_g N_A_384_74#_c_570_n N_A_384_74#_c_537_n
+ N_A_384_74#_c_538_n N_A_384_74#_c_539_n N_A_384_74#_c_571_n
+ N_A_384_74#_c_572_n N_A_384_74#_c_540_n N_A_384_74#_c_573_n
+ N_A_384_74#_c_541_n N_A_384_74#_c_574_n N_A_384_74#_c_542_n
+ N_A_384_74#_c_543_n N_A_384_74#_c_576_n N_A_384_74#_c_544_n
+ N_A_384_74#_c_577_n N_A_384_74#_c_545_n N_A_384_74#_c_546_n
+ N_A_384_74#_c_547_n N_A_384_74#_c_548_n N_A_384_74#_c_549_n
+ N_A_384_74#_c_550_n N_A_384_74#_c_551_n N_A_384_74#_c_552_n
+ N_A_384_74#_c_553_n PM_SKY130_FD_SC_MS__BUFINV_16%A_384_74#
x_PM_SKY130_FD_SC_MS__BUFINV_16%VPWR N_VPWR_M1001_d N_VPWR_M1005_d
+ N_VPWR_M1016_s N_VPWR_M1025_s N_VPWR_M1033_s N_VPWR_M1006_s N_VPWR_M1010_s
+ N_VPWR_M1014_s N_VPWR_M1020_s N_VPWR_M1030_s N_VPWR_M1034_s N_VPWR_M1040_s
+ N_VPWR_M1045_s N_VPWR_c_974_n N_VPWR_c_975_n N_VPWR_c_976_n N_VPWR_c_977_n
+ N_VPWR_c_978_n N_VPWR_c_979_n N_VPWR_c_980_n N_VPWR_c_981_n N_VPWR_c_982_n
+ N_VPWR_c_983_n N_VPWR_c_984_n N_VPWR_c_985_n N_VPWR_c_986_n N_VPWR_c_987_n
+ N_VPWR_c_988_n N_VPWR_c_989_n N_VPWR_c_990_n N_VPWR_c_991_n N_VPWR_c_992_n
+ N_VPWR_c_993_n N_VPWR_c_994_n N_VPWR_c_995_n N_VPWR_c_996_n N_VPWR_c_997_n
+ N_VPWR_c_998_n N_VPWR_c_999_n N_VPWR_c_1000_n N_VPWR_c_1001_n N_VPWR_c_1002_n
+ VPWR N_VPWR_c_1003_n N_VPWR_c_1004_n N_VPWR_c_1005_n N_VPWR_c_1006_n
+ N_VPWR_c_1007_n N_VPWR_c_1008_n N_VPWR_c_1009_n N_VPWR_c_1010_n
+ N_VPWR_c_1011_n N_VPWR_c_973_n PM_SKY130_FD_SC_MS__BUFINV_16%VPWR
x_PM_SKY130_FD_SC_MS__BUFINV_16%Y N_Y_M1003_s N_Y_M1013_s N_Y_M1022_s
+ N_Y_M1027_s N_Y_M1032_s N_Y_M1038_s N_Y_M1041_s N_Y_M1044_s N_Y_M1004_d
+ N_Y_M1008_d N_Y_M1012_d N_Y_M1017_d N_Y_M1024_d N_Y_M1031_d N_Y_M1037_d
+ N_Y_M1043_d N_Y_c_1195_n N_Y_c_1196_n N_Y_c_1197_n N_Y_c_1198_n N_Y_c_1207_n
+ N_Y_c_1262_n N_Y_c_1208_n N_Y_c_1199_n N_Y_c_1277_n N_Y_c_1210_n N_Y_c_1200_n
+ N_Y_c_1201_n N_Y_c_1202_n N_Y_c_1311_n N_Y_c_1314_n N_Y_c_1318_n N_Y_c_1321_n
+ N_Y_c_1214_n Y N_Y_c_1215_n N_Y_c_1216_n N_Y_c_1217_n N_Y_c_1218_n
+ N_Y_c_1219_n N_Y_c_1336_n N_Y_c_1358_n PM_SKY130_FD_SC_MS__BUFINV_16%Y
x_PM_SKY130_FD_SC_MS__BUFINV_16%VGND N_VGND_M1000_s N_VGND_M1047_s
+ N_VGND_M1015_s N_VGND_M1026_s N_VGND_M1049_s N_VGND_M1007_d N_VGND_M1021_d
+ N_VGND_M1023_d N_VGND_M1028_d N_VGND_M1036_d N_VGND_M1039_d N_VGND_M1042_d
+ N_VGND_M1046_d N_VGND_c_1449_n N_VGND_c_1450_n N_VGND_c_1451_n N_VGND_c_1452_n
+ N_VGND_c_1453_n N_VGND_c_1454_n N_VGND_c_1455_n N_VGND_c_1456_n
+ N_VGND_c_1457_n N_VGND_c_1458_n N_VGND_c_1459_n N_VGND_c_1460_n
+ N_VGND_c_1461_n N_VGND_c_1462_n N_VGND_c_1463_n N_VGND_c_1464_n
+ N_VGND_c_1465_n N_VGND_c_1466_n N_VGND_c_1467_n N_VGND_c_1468_n
+ N_VGND_c_1469_n N_VGND_c_1470_n VGND N_VGND_c_1471_n N_VGND_c_1472_n
+ N_VGND_c_1473_n N_VGND_c_1474_n N_VGND_c_1475_n N_VGND_c_1476_n
+ N_VGND_c_1477_n N_VGND_c_1478_n N_VGND_c_1479_n N_VGND_c_1480_n
+ N_VGND_c_1481_n N_VGND_c_1482_n N_VGND_c_1483_n N_VGND_c_1484_n
+ N_VGND_c_1485_n N_VGND_c_1486_n N_VGND_c_1487_n N_VGND_c_1488_n
+ PM_SKY130_FD_SC_MS__BUFINV_16%VGND
cc_1 VNB N_A_M1000_g 0.0327337f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_M1035_g 0.0240034f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.74
cc_3 VNB N_A_M1047_g 0.0227235f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=0.74
cc_4 VNB N_A_c_234_n 0.0166485f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_5 VNB N_A_c_235_n 0.0570679f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.515
cc_6 VNB N_A_27_74#_M1011_g 0.0208043f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.74
cc_7 VNB N_A_27_74#_M1009_g 0.00161032f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=2.4
cc_8 VNB N_A_27_74#_M1015_g 0.0203546f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=0.74
cc_9 VNB N_A_27_74#_M1016_g 0.00156549f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_10 VNB N_A_27_74#_M1018_g 0.0209331f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_11 VNB N_A_27_74#_M1019_g 0.00154301f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_12 VNB N_A_27_74#_M1026_g 0.0211968f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_13 VNB N_A_27_74#_M1025_g 0.00154124f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.515
cc_14 VNB N_A_27_74#_M1048_g 0.0210803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_74#_M1029_g 0.00142151f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_16 VNB N_A_27_74#_c_308_n 0.00890084f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.565
cc_17 VNB N_A_27_74#_M1049_g 0.0215143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_74#_M1033_g 0.00937171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_311_n 0.0078775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_74#_c_312_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_74#_c_313_n 0.00360698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_314_n 0.00998227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_74#_c_315_n 0.00179995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_74#_c_316_n 0.00415915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_74#_c_317_n 4.30857e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_74#_c_318_n 6.65696e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_74#_c_319_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_74#_c_320_n 0.00563641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_74#_c_321_n 0.0981532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_384_74#_M1003_g 0.0216367f $X=-0.19 $Y=-0.245 $X2=1.415 $Y2=1.35
cc_31 VNB N_A_384_74#_M1004_g 0.00131629f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_32 VNB N_A_384_74#_M1007_g 0.0204987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_384_74#_M1006_g 0.00130405f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.515
cc_34 VNB N_A_384_74#_M1013_g 0.021162f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.515
cc_35 VNB N_A_384_74#_M1008_g 0.00130405f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_36 VNB N_A_384_74#_M1021_g 0.021363f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_37 VNB N_A_384_74#_M1010_g 0.00130405f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_38 VNB N_A_384_74#_M1022_g 0.0211843f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.565
cc_39 VNB N_A_384_74#_M1012_g 0.00130405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_384_74#_M1023_g 0.0213617f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_384_74#_M1014_g 0.00130405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_384_74#_M1017_g 0.00130405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_384_74#_M1027_g 0.0211822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_384_74#_M1028_g 0.0213612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_384_74#_M1020_g 0.00130405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_384_74#_M1024_g 0.00130405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_384_74#_M1032_g 0.0211812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_384_74#_M1030_g 0.00136248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_384_74#_M1036_g 0.0213612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_384_74#_M1031_g 0.00136264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_384_74#_M1038_g 0.0211812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_384_74#_M1034_g 0.00136248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_384_74#_M1039_g 0.0213612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_384_74#_M1037_g 0.00136264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_384_74#_M1041_g 0.0211812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_384_74#_M1042_g 0.0213612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_384_74#_M1040_g 0.00131638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_384_74#_M1043_g 0.00147155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_384_74#_M1044_g 0.021184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_384_74#_M1046_g 0.0260277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_384_74#_M1045_g 0.00247541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_384_74#_c_537_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_384_74#_c_538_n 0.00275044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_384_74#_c_539_n 0.00140873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_384_74#_c_540_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_384_74#_c_541_n 0.00374208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_384_74#_c_542_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_384_74#_c_543_n 0.00686392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_384_74#_c_544_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_384_74#_c_545_n 0.00180003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_384_74#_c_546_n 0.00109754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_384_74#_c_547_n 0.00177315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_384_74#_c_548_n 0.00176232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_384_74#_c_549_n 0.00176506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_384_74#_c_550_n 0.00176778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_384_74#_c_551_n 0.00176778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_384_74#_c_552_n 0.00183757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_384_74#_c_553_n 0.372846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VPWR_c_973_n 0.502022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_Y_c_1195_n 0.00378061f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_81 VNB N_Y_c_1196_n 0.00574953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_Y_c_1197_n 0.00397969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_Y_c_1198_n 0.00398355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_Y_c_1199_n 0.00398531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_Y_c_1200_n 0.00398531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_Y_c_1201_n 0.00398531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_Y_c_1202_n 0.00269539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1449_n 0.00563075f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.515
cc_89 VNB N_VGND_c_1450_n 0.00258815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1451_n 0.0040939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1452_n 0.00495983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1453_n 0.00754943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1454_n 0.00419598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1455_n 0.00502158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1456_n 0.00498499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1457_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1458_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1459_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1460_n 0.00508214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1461_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1462_n 0.0547214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1463_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1464_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1465_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1466_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1467_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1468_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1469_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1470_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1471_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1472_n 0.0172409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1473_n 0.0175258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1474_n 0.0170514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1475_n 0.0169733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1476_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1477_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1478_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1479_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1480_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1481_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1482_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1483_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1484_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1485_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1486_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1487_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1488_n 0.623946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VPB N_A_M1001_g 0.027583f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_129 VPB N_A_M1002_g 0.0204965f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_130 VPB N_A_M1005_g 0.0213785f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=2.4
cc_131 VPB N_A_c_234_n 0.0131369f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_132 VPB N_A_c_235_n 0.00839531f $X=-0.19 $Y=1.66 $X2=1.415 $Y2=1.515
cc_133 VPB N_A_27_74#_M1009_g 0.0229895f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=2.4
cc_134 VPB N_A_27_74#_M1016_g 0.0223087f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_135 VPB N_A_27_74#_M1019_g 0.0220607f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_136 VPB N_A_27_74#_M1025_g 0.0220351f $X=-0.19 $Y=1.66 $X2=1.415 $Y2=1.515
cc_137 VPB N_A_27_74#_M1029_g 0.0214742f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_138 VPB N_A_27_74#_M1033_g 0.021519f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_27_74#_c_328_n 0.00739392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_27_74#_c_329_n 0.0352219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_27_74#_c_330_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_27_74#_c_317_n 0.00283436f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_384_74#_M1004_g 0.0215608f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_144 VPB N_A_384_74#_M1006_g 0.0214304f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.515
cc_145 VPB N_A_384_74#_M1008_g 0.0211752f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_146 VPB N_A_384_74#_M1010_g 0.021432f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_147 VPB N_A_384_74#_M1012_g 0.0211768f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_384_74#_M1014_g 0.0214314f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_384_74#_M1017_g 0.0211786f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_384_74#_M1020_g 0.0214312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_384_74#_M1024_g 0.0211808f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_384_74#_M1030_g 0.0220418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_384_74#_M1031_g 0.0217901f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_384_74#_M1034_g 0.0220414f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_384_74#_M1037_g 0.0217879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_384_74#_M1040_g 0.0215577f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_384_74#_M1043_g 0.0223417f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_384_74#_M1045_g 0.0284154f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_384_74#_c_570_n 0.00248769f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_384_74#_c_571_n 0.00219429f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_384_74#_c_572_n 0.00236567f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_384_74#_c_573_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_384_74#_c_574_n 0.002854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_384_74#_c_543_n 0.00165499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_384_74#_c_576_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_384_74#_c_577_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_384_74#_c_545_n 0.0160836f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_384_74#_c_546_n 0.00147325f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_384_74#_c_547_n 0.00153481f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_384_74#_c_548_n 0.00192338f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_384_74#_c_549_n 0.00218971f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_384_74#_c_550_n 0.0019973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_384_74#_c_551_n 0.00173921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_384_74#_c_552_n 0.00195978f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_974_n 0.00797179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_975_n 0.00797541f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.565
cc_177 VPB N_VPWR_c_976_n 0.00797179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_977_n 0.00797179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_978_n 0.00797179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_979_n 0.00797179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_980_n 0.00797179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_981_n 0.00797179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_982_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_983_n 0.00797179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_984_n 0.00862436f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_985_n 0.00873731f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_986_n 0.00850289f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_987_n 0.0111306f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_988_n 0.0645583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_989_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_990_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_991_n 0.0212277f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_992_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_993_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_994_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_995_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_996_n 0.00319223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_997_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_998_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_999_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1000_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1001_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1002_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1003_n 0.0205913f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1004_n 0.020445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1005_n 0.0201268f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1006_n 0.0207632f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1007_n 0.0234893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1008_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1009_n 0.00430193f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1010_n 0.00449427f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1011_n 0.00410958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_973_n 0.122986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_Y_c_1195_n 0.0010898f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_215 VPB N_Y_c_1196_n 0.00127452f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_Y_c_1197_n 0.00128982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_Y_c_1198_n 0.00126175f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_Y_c_1207_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_Y_c_1208_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_Y_c_1199_n 0.00125184f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_Y_c_1210_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_Y_c_1200_n 0.00125369f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_Y_c_1201_n 0.0012661f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_Y_c_1202_n 0.00126196f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_Y_c_1214_n 2.03637e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_Y_c_1215_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_Y_c_1216_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_Y_c_1217_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_Y_c_1218_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_Y_c_1219_n 0.00276853f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 N_A_M1047_g N_A_27_74#_M1011_g 0.0296537f $X=1.415 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A_M1005_g N_A_27_74#_M1009_g 0.0224044f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_233 N_A_M1000_g N_A_27_74#_c_312_n 0.00159319f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A_M1001_g N_A_27_74#_c_328_n 8.84614e-19 $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_235 N_A_c_234_n N_A_27_74#_c_328_n 0.0259449f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_236 N_A_M1001_g N_A_27_74#_c_329_n 0.0121004f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_237 N_A_M1002_g N_A_27_74#_c_329_n 6.50516e-19 $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_238 N_A_M1000_g N_A_27_74#_c_313_n 0.013995f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_239 N_A_M1035_g N_A_27_74#_c_313_n 0.0141485f $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A_c_234_n N_A_27_74#_c_313_n 0.056571f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_241 N_A_c_235_n N_A_27_74#_c_313_n 0.00386308f $X=1.415 $Y=1.515 $X2=0 $Y2=0
cc_242 N_A_c_234_n N_A_27_74#_c_314_n 0.0216404f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_243 N_A_M1001_g N_A_27_74#_c_344_n 0.012931f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_244 N_A_M1002_g N_A_27_74#_c_344_n 0.012931f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_245 N_A_c_234_n N_A_27_74#_c_344_n 0.0391869f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_246 N_A_c_235_n N_A_27_74#_c_344_n 4.90767e-19 $X=1.415 $Y=1.515 $X2=0 $Y2=0
cc_247 N_A_M1001_g N_A_27_74#_c_330_n 6.50516e-19 $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_248 N_A_M1002_g N_A_27_74#_c_330_n 0.0119382f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_249 N_A_M1005_g N_A_27_74#_c_330_n 0.01199f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_250 N_A_M1035_g N_A_27_74#_c_315_n 4.0877e-19 $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_251 N_A_M1047_g N_A_27_74#_c_315_n 3.92313e-19 $X=1.415 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A_M1047_g N_A_27_74#_c_316_n 0.0139897f $X=1.415 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A_c_234_n N_A_27_74#_c_316_n 0.0107488f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_254 N_A_c_235_n N_A_27_74#_c_316_n 4.15062e-19 $X=1.415 $Y=1.515 $X2=0 $Y2=0
cc_255 N_A_M1005_g N_A_27_74#_c_356_n 0.0150125f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_256 N_A_c_234_n N_A_27_74#_c_356_n 0.00580317f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_257 N_A_M1005_g N_A_27_74#_c_317_n 0.00353478f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_258 N_A_M1002_g N_A_27_74#_c_359_n 8.84614e-19 $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_259 N_A_M1005_g N_A_27_74#_c_359_n 8.84614e-19 $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_260 N_A_c_234_n N_A_27_74#_c_359_n 0.0235495f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_261 N_A_c_235_n N_A_27_74#_c_359_n 5.5407e-19 $X=1.415 $Y=1.515 $X2=0 $Y2=0
cc_262 N_A_c_234_n N_A_27_74#_c_319_n 0.0146029f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_263 N_A_c_235_n N_A_27_74#_c_319_n 0.00240845f $X=1.415 $Y=1.515 $X2=0 $Y2=0
cc_264 N_A_M1047_g N_A_27_74#_c_320_n 0.0040282f $X=1.415 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A_c_234_n N_A_27_74#_c_320_n 0.0341212f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_266 N_A_c_235_n N_A_27_74#_c_320_n 0.00353478f $X=1.415 $Y=1.515 $X2=0 $Y2=0
cc_267 N_A_c_235_n N_A_27_74#_c_321_n 0.0224044f $X=1.415 $Y=1.515 $X2=0 $Y2=0
cc_268 N_A_M1005_g N_A_384_74#_c_570_n 7.45782e-19 $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_269 N_A_M1001_g N_VPWR_c_974_n 0.0027763f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_270 N_A_M1002_g N_VPWR_c_974_n 0.0027763f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_271 N_A_M1005_g N_VPWR_c_975_n 0.0027763f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_272 N_A_M1002_g N_VPWR_c_989_n 0.005209f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_273 N_A_M1005_g N_VPWR_c_989_n 0.005209f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_274 N_A_M1001_g N_VPWR_c_1007_n 0.005209f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_275 N_A_M1001_g N_VPWR_c_973_n 0.00986025f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_276 N_A_M1002_g N_VPWR_c_973_n 0.00982266f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_277 N_A_M1005_g N_VPWR_c_973_n 0.00982376f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_278 N_A_M1000_g N_VGND_c_1449_n 0.0136841f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_279 N_A_M1035_g N_VGND_c_1449_n 0.00425844f $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_280 N_A_M1035_g N_VGND_c_1450_n 4.80113e-19 $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_281 N_A_M1047_g N_VGND_c_1450_n 0.0107133f $X=1.415 $Y=0.74 $X2=0 $Y2=0
cc_282 N_A_M1000_g N_VGND_c_1471_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_283 N_A_M1035_g N_VGND_c_1472_n 0.00461464f $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_284 N_A_M1047_g N_VGND_c_1472_n 0.00383152f $X=1.415 $Y=0.74 $X2=0 $Y2=0
cc_285 N_A_M1000_g N_VGND_c_1488_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_286 N_A_M1035_g N_VGND_c_1488_n 0.00908454f $X=0.985 $Y=0.74 $X2=0 $Y2=0
cc_287 N_A_M1047_g N_VGND_c_1488_n 0.0075754f $X=1.415 $Y=0.74 $X2=0 $Y2=0
cc_288 N_A_27_74#_M1049_g N_A_384_74#_M1003_g 0.020096f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_289 N_A_27_74#_M1033_g N_A_384_74#_M1004_g 0.0165919f $X=4.13 $Y=2.4 $X2=0
+ $Y2=0
cc_290 N_A_27_74#_M1009_g N_A_384_74#_c_570_n 0.0136341f $X=1.86 $Y=2.4 $X2=0
+ $Y2=0
cc_291 N_A_27_74#_M1016_g N_A_384_74#_c_570_n 0.0143533f $X=2.33 $Y=2.4 $X2=0
+ $Y2=0
cc_292 N_A_27_74#_M1019_g N_A_384_74#_c_570_n 6.97946e-19 $X=2.78 $Y=2.4 $X2=0
+ $Y2=0
cc_293 N_A_27_74#_c_330_n N_A_384_74#_c_570_n 0.00454938f $X=1.185 $Y=2.815
+ $X2=0 $Y2=0
cc_294 N_A_27_74#_c_356_n N_A_384_74#_c_570_n 0.011936f $X=1.6 $Y=2.035 $X2=0
+ $Y2=0
cc_295 N_A_27_74#_M1011_g N_A_384_74#_c_537_n 3.92313e-19 $X=1.845 $Y=0.74 $X2=0
+ $Y2=0
cc_296 N_A_27_74#_M1015_g N_A_384_74#_c_537_n 3.92313e-19 $X=2.275 $Y=0.74 $X2=0
+ $Y2=0
cc_297 N_A_27_74#_M1015_g N_A_384_74#_c_538_n 0.0124383f $X=2.275 $Y=0.74 $X2=0
+ $Y2=0
cc_298 N_A_27_74#_M1018_g N_A_384_74#_c_538_n 0.0111034f $X=2.705 $Y=0.74 $X2=0
+ $Y2=0
cc_299 N_A_27_74#_c_318_n N_A_384_74#_c_538_n 0.0447482f $X=3.295 $Y=1.465 $X2=0
+ $Y2=0
cc_300 N_A_27_74#_c_321_n N_A_384_74#_c_538_n 0.00251785f $X=3.77 $Y=1.465 $X2=0
+ $Y2=0
cc_301 N_A_27_74#_c_318_n N_A_384_74#_c_539_n 0.0143381f $X=3.295 $Y=1.465 $X2=0
+ $Y2=0
cc_302 N_A_27_74#_c_320_n N_A_384_74#_c_539_n 0.00140469f $X=1.685 $Y=1.095
+ $X2=0 $Y2=0
cc_303 N_A_27_74#_c_321_n N_A_384_74#_c_539_n 0.00244789f $X=3.77 $Y=1.465 $X2=0
+ $Y2=0
cc_304 N_A_27_74#_M1016_g N_A_384_74#_c_571_n 0.012931f $X=2.33 $Y=2.4 $X2=0
+ $Y2=0
cc_305 N_A_27_74#_M1019_g N_A_384_74#_c_571_n 0.012931f $X=2.78 $Y=2.4 $X2=0
+ $Y2=0
cc_306 N_A_27_74#_c_318_n N_A_384_74#_c_571_n 0.0416512f $X=3.295 $Y=1.465 $X2=0
+ $Y2=0
cc_307 N_A_27_74#_c_321_n N_A_384_74#_c_571_n 0.00225424f $X=3.77 $Y=1.465 $X2=0
+ $Y2=0
cc_308 N_A_27_74#_M1009_g N_A_384_74#_c_572_n 0.0023781f $X=1.86 $Y=2.4 $X2=0
+ $Y2=0
cc_309 N_A_27_74#_M1016_g N_A_384_74#_c_572_n 0.00138281f $X=2.33 $Y=2.4 $X2=0
+ $Y2=0
cc_310 N_A_27_74#_c_356_n N_A_384_74#_c_572_n 0.00169302f $X=1.6 $Y=2.035 $X2=0
+ $Y2=0
cc_311 N_A_27_74#_c_317_n N_A_384_74#_c_572_n 0.00779204f $X=1.685 $Y=1.95 $X2=0
+ $Y2=0
cc_312 N_A_27_74#_c_318_n N_A_384_74#_c_572_n 0.0276532f $X=3.295 $Y=1.465 $X2=0
+ $Y2=0
cc_313 N_A_27_74#_c_321_n N_A_384_74#_c_572_n 0.00272029f $X=3.77 $Y=1.465 $X2=0
+ $Y2=0
cc_314 N_A_27_74#_M1015_g N_A_384_74#_c_540_n 6.20738e-19 $X=2.275 $Y=0.74 $X2=0
+ $Y2=0
cc_315 N_A_27_74#_M1018_g N_A_384_74#_c_540_n 0.00866629f $X=2.705 $Y=0.74 $X2=0
+ $Y2=0
cc_316 N_A_27_74#_M1026_g N_A_384_74#_c_540_n 3.97481e-19 $X=3.135 $Y=0.74 $X2=0
+ $Y2=0
cc_317 N_A_27_74#_M1016_g N_A_384_74#_c_573_n 6.97946e-19 $X=2.33 $Y=2.4 $X2=0
+ $Y2=0
cc_318 N_A_27_74#_M1019_g N_A_384_74#_c_573_n 0.0143027f $X=2.78 $Y=2.4 $X2=0
+ $Y2=0
cc_319 N_A_27_74#_M1025_g N_A_384_74#_c_573_n 0.0143027f $X=3.23 $Y=2.4 $X2=0
+ $Y2=0
cc_320 N_A_27_74#_M1029_g N_A_384_74#_c_573_n 6.97946e-19 $X=3.68 $Y=2.4 $X2=0
+ $Y2=0
cc_321 N_A_27_74#_M1026_g N_A_384_74#_c_541_n 0.0128832f $X=3.135 $Y=0.74 $X2=0
+ $Y2=0
cc_322 N_A_27_74#_M1048_g N_A_384_74#_c_541_n 0.0133712f $X=3.635 $Y=0.74 $X2=0
+ $Y2=0
cc_323 N_A_27_74#_c_318_n N_A_384_74#_c_541_n 0.0335994f $X=3.295 $Y=1.465 $X2=0
+ $Y2=0
cc_324 N_A_27_74#_c_321_n N_A_384_74#_c_541_n 0.00429413f $X=3.77 $Y=1.465 $X2=0
+ $Y2=0
cc_325 N_A_27_74#_M1025_g N_A_384_74#_c_574_n 0.012931f $X=3.23 $Y=2.4 $X2=0
+ $Y2=0
cc_326 N_A_27_74#_M1029_g N_A_384_74#_c_574_n 0.0148841f $X=3.68 $Y=2.4 $X2=0
+ $Y2=0
cc_327 N_A_27_74#_c_318_n N_A_384_74#_c_574_n 0.0212014f $X=3.295 $Y=1.465 $X2=0
+ $Y2=0
cc_328 N_A_27_74#_c_321_n N_A_384_74#_c_574_n 0.00233302f $X=3.77 $Y=1.465 $X2=0
+ $Y2=0
cc_329 N_A_27_74#_M1026_g N_A_384_74#_c_542_n 8.7513e-19 $X=3.135 $Y=0.74 $X2=0
+ $Y2=0
cc_330 N_A_27_74#_M1048_g N_A_384_74#_c_542_n 0.00862472f $X=3.635 $Y=0.74 $X2=0
+ $Y2=0
cc_331 N_A_27_74#_M1049_g N_A_384_74#_c_542_n 3.97481e-19 $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_332 N_A_27_74#_M1026_g N_A_384_74#_c_543_n 8.02787e-19 $X=3.135 $Y=0.74 $X2=0
+ $Y2=0
cc_333 N_A_27_74#_M1025_g N_A_384_74#_c_543_n 8.00048e-19 $X=3.23 $Y=2.4 $X2=0
+ $Y2=0
cc_334 N_A_27_74#_M1048_g N_A_384_74#_c_543_n 0.00529244f $X=3.635 $Y=0.74 $X2=0
+ $Y2=0
cc_335 N_A_27_74#_M1029_g N_A_384_74#_c_543_n 0.00628049f $X=3.68 $Y=2.4 $X2=0
+ $Y2=0
cc_336 N_A_27_74#_c_308_n N_A_384_74#_c_543_n 0.0105749f $X=3.99 $Y=1.375 $X2=0
+ $Y2=0
cc_337 N_A_27_74#_M1049_g N_A_384_74#_c_543_n 0.00453721f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_338 N_A_27_74#_M1033_g N_A_384_74#_c_543_n 0.0216336f $X=4.13 $Y=2.4 $X2=0
+ $Y2=0
cc_339 N_A_27_74#_c_311_n N_A_384_74#_c_543_n 0.0113158f $X=4.105 $Y=1.375 $X2=0
+ $Y2=0
cc_340 N_A_27_74#_c_318_n N_A_384_74#_c_543_n 0.0185957f $X=3.295 $Y=1.465 $X2=0
+ $Y2=0
cc_341 N_A_27_74#_c_321_n N_A_384_74#_c_543_n 0.010562f $X=3.77 $Y=1.465 $X2=0
+ $Y2=0
cc_342 N_A_27_74#_M1025_g N_A_384_74#_c_576_n 6.97946e-19 $X=3.23 $Y=2.4 $X2=0
+ $Y2=0
cc_343 N_A_27_74#_M1029_g N_A_384_74#_c_576_n 0.0143027f $X=3.68 $Y=2.4 $X2=0
+ $Y2=0
cc_344 N_A_27_74#_M1033_g N_A_384_74#_c_576_n 0.0130665f $X=4.13 $Y=2.4 $X2=0
+ $Y2=0
cc_345 N_A_27_74#_M1018_g N_A_384_74#_c_544_n 9.7541e-19 $X=2.705 $Y=0.74 $X2=0
+ $Y2=0
cc_346 N_A_27_74#_c_318_n N_A_384_74#_c_544_n 0.0209731f $X=3.295 $Y=1.465 $X2=0
+ $Y2=0
cc_347 N_A_27_74#_c_321_n N_A_384_74#_c_544_n 0.00268454f $X=3.77 $Y=1.465 $X2=0
+ $Y2=0
cc_348 N_A_27_74#_M1019_g N_A_384_74#_c_577_n 0.00135419f $X=2.78 $Y=2.4 $X2=0
+ $Y2=0
cc_349 N_A_27_74#_M1025_g N_A_384_74#_c_577_n 0.00135419f $X=3.23 $Y=2.4 $X2=0
+ $Y2=0
cc_350 N_A_27_74#_c_318_n N_A_384_74#_c_577_n 0.0275631f $X=3.295 $Y=1.465 $X2=0
+ $Y2=0
cc_351 N_A_27_74#_c_321_n N_A_384_74#_c_577_n 0.00241214f $X=3.77 $Y=1.465 $X2=0
+ $Y2=0
cc_352 N_A_27_74#_M1033_g N_A_384_74#_c_545_n 0.00322271f $X=4.13 $Y=2.4 $X2=0
+ $Y2=0
cc_353 N_A_27_74#_c_311_n N_A_384_74#_c_553_n 0.0165919f $X=4.105 $Y=1.375 $X2=0
+ $Y2=0
cc_354 N_A_27_74#_c_344_n N_VPWR_M1001_d 0.00314376f $X=1.02 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_355 N_A_27_74#_c_356_n N_VPWR_M1005_d 0.00359894f $X=1.6 $Y=2.035 $X2=0 $Y2=0
cc_356 N_A_27_74#_c_317_n N_VPWR_M1005_d 0.00141518f $X=1.685 $Y=1.95 $X2=0
+ $Y2=0
cc_357 N_A_27_74#_c_329_n N_VPWR_c_974_n 0.0233699f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_358 N_A_27_74#_c_344_n N_VPWR_c_974_n 0.0126919f $X=1.02 $Y=2.035 $X2=0 $Y2=0
cc_359 N_A_27_74#_c_330_n N_VPWR_c_974_n 0.0233699f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_360 N_A_27_74#_M1009_g N_VPWR_c_975_n 0.00278184f $X=1.86 $Y=2.4 $X2=0 $Y2=0
cc_361 N_A_27_74#_c_330_n N_VPWR_c_975_n 0.0233699f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_362 N_A_27_74#_c_356_n N_VPWR_c_975_n 0.0136051f $X=1.6 $Y=2.035 $X2=0 $Y2=0
cc_363 N_A_27_74#_M1016_g N_VPWR_c_976_n 0.00329146f $X=2.33 $Y=2.4 $X2=0 $Y2=0
cc_364 N_A_27_74#_M1019_g N_VPWR_c_976_n 0.00329146f $X=2.78 $Y=2.4 $X2=0 $Y2=0
cc_365 N_A_27_74#_M1025_g N_VPWR_c_977_n 0.00329146f $X=3.23 $Y=2.4 $X2=0 $Y2=0
cc_366 N_A_27_74#_M1029_g N_VPWR_c_977_n 0.00329146f $X=3.68 $Y=2.4 $X2=0 $Y2=0
cc_367 N_A_27_74#_M1033_g N_VPWR_c_978_n 0.0027763f $X=4.13 $Y=2.4 $X2=0 $Y2=0
cc_368 N_A_27_74#_c_330_n N_VPWR_c_989_n 0.0144623f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_369 N_A_27_74#_M1009_g N_VPWR_c_991_n 0.0054356f $X=1.86 $Y=2.4 $X2=0 $Y2=0
cc_370 N_A_27_74#_M1016_g N_VPWR_c_991_n 0.005209f $X=2.33 $Y=2.4 $X2=0 $Y2=0
cc_371 N_A_27_74#_M1019_g N_VPWR_c_993_n 0.005209f $X=2.78 $Y=2.4 $X2=0 $Y2=0
cc_372 N_A_27_74#_M1025_g N_VPWR_c_993_n 0.005209f $X=3.23 $Y=2.4 $X2=0 $Y2=0
cc_373 N_A_27_74#_M1029_g N_VPWR_c_995_n 0.005209f $X=3.68 $Y=2.4 $X2=0 $Y2=0
cc_374 N_A_27_74#_M1033_g N_VPWR_c_995_n 0.005209f $X=4.13 $Y=2.4 $X2=0 $Y2=0
cc_375 N_A_27_74#_c_329_n N_VPWR_c_1007_n 0.014549f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_376 N_A_27_74#_M1009_g N_VPWR_c_973_n 0.0105595f $X=1.86 $Y=2.4 $X2=0 $Y2=0
cc_377 N_A_27_74#_M1016_g N_VPWR_c_973_n 0.00982467f $X=2.33 $Y=2.4 $X2=0 $Y2=0
cc_378 N_A_27_74#_M1019_g N_VPWR_c_973_n 0.00982266f $X=2.78 $Y=2.4 $X2=0 $Y2=0
cc_379 N_A_27_74#_M1025_g N_VPWR_c_973_n 0.00982266f $X=3.23 $Y=2.4 $X2=0 $Y2=0
cc_380 N_A_27_74#_M1029_g N_VPWR_c_973_n 0.00982266f $X=3.68 $Y=2.4 $X2=0 $Y2=0
cc_381 N_A_27_74#_M1033_g N_VPWR_c_973_n 0.00982376f $X=4.13 $Y=2.4 $X2=0 $Y2=0
cc_382 N_A_27_74#_c_329_n N_VPWR_c_973_n 0.0119743f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_383 N_A_27_74#_c_330_n N_VPWR_c_973_n 0.0118344f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_384 N_A_27_74#_M1049_g N_Y_c_1195_n 0.0010331f $X=4.065 $Y=0.74 $X2=0 $Y2=0
cc_385 N_A_27_74#_M1033_g N_Y_c_1195_n 4.88414e-19 $X=4.13 $Y=2.4 $X2=0 $Y2=0
cc_386 N_A_27_74#_c_311_n N_Y_c_1195_n 4.13338e-19 $X=4.105 $Y=1.375 $X2=0 $Y2=0
cc_387 N_A_27_74#_c_313_n N_VGND_M1000_s 0.00240242f $X=1.115 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_388 N_A_27_74#_c_316_n N_VGND_M1047_s 8.02634e-19 $X=1.6 $Y=1.095 $X2=0 $Y2=0
cc_389 N_A_27_74#_c_320_n N_VGND_M1047_s 0.00168914f $X=1.685 $Y=1.095 $X2=0
+ $Y2=0
cc_390 N_A_27_74#_c_312_n N_VGND_c_1449_n 0.0182902f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_391 N_A_27_74#_c_313_n N_VGND_c_1449_n 0.0201731f $X=1.115 $Y=1.095 $X2=0
+ $Y2=0
cc_392 N_A_27_74#_c_315_n N_VGND_c_1449_n 0.00118247f $X=1.2 $Y=0.515 $X2=0
+ $Y2=0
cc_393 N_A_27_74#_M1011_g N_VGND_c_1450_n 0.0108544f $X=1.845 $Y=0.74 $X2=0
+ $Y2=0
cc_394 N_A_27_74#_M1015_g N_VGND_c_1450_n 4.71636e-19 $X=2.275 $Y=0.74 $X2=0
+ $Y2=0
cc_395 N_A_27_74#_c_315_n N_VGND_c_1450_n 0.0182488f $X=1.2 $Y=0.515 $X2=0 $Y2=0
cc_396 N_A_27_74#_c_316_n N_VGND_c_1450_n 0.00609809f $X=1.6 $Y=1.095 $X2=0
+ $Y2=0
cc_397 N_A_27_74#_c_318_n N_VGND_c_1450_n 8.33225e-19 $X=3.295 $Y=1.465 $X2=0
+ $Y2=0
cc_398 N_A_27_74#_c_320_n N_VGND_c_1450_n 0.0100981f $X=1.685 $Y=1.095 $X2=0
+ $Y2=0
cc_399 N_A_27_74#_M1011_g N_VGND_c_1451_n 4.57991e-19 $X=1.845 $Y=0.74 $X2=0
+ $Y2=0
cc_400 N_A_27_74#_M1015_g N_VGND_c_1451_n 0.00900784f $X=2.275 $Y=0.74 $X2=0
+ $Y2=0
cc_401 N_A_27_74#_M1018_g N_VGND_c_1451_n 0.00183835f $X=2.705 $Y=0.74 $X2=0
+ $Y2=0
cc_402 N_A_27_74#_M1018_g N_VGND_c_1452_n 5.04273e-19 $X=2.705 $Y=0.74 $X2=0
+ $Y2=0
cc_403 N_A_27_74#_M1026_g N_VGND_c_1452_n 0.0097054f $X=3.135 $Y=0.74 $X2=0
+ $Y2=0
cc_404 N_A_27_74#_M1048_g N_VGND_c_1452_n 0.00397833f $X=3.635 $Y=0.74 $X2=0
+ $Y2=0
cc_405 N_A_27_74#_M1048_g N_VGND_c_1453_n 6.13182e-19 $X=3.635 $Y=0.74 $X2=0
+ $Y2=0
cc_406 N_A_27_74#_M1049_g N_VGND_c_1453_n 0.0134222f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_407 N_A_27_74#_c_311_n N_VGND_c_1453_n 6.25621e-19 $X=4.105 $Y=1.375 $X2=0
+ $Y2=0
cc_408 N_A_27_74#_M1011_g N_VGND_c_1463_n 0.00383152f $X=1.845 $Y=0.74 $X2=0
+ $Y2=0
cc_409 N_A_27_74#_M1015_g N_VGND_c_1463_n 0.00383152f $X=2.275 $Y=0.74 $X2=0
+ $Y2=0
cc_410 N_A_27_74#_M1018_g N_VGND_c_1465_n 0.00434272f $X=2.705 $Y=0.74 $X2=0
+ $Y2=0
cc_411 N_A_27_74#_M1026_g N_VGND_c_1465_n 0.00383152f $X=3.135 $Y=0.74 $X2=0
+ $Y2=0
cc_412 N_A_27_74#_M1048_g N_VGND_c_1467_n 0.00434272f $X=3.635 $Y=0.74 $X2=0
+ $Y2=0
cc_413 N_A_27_74#_M1049_g N_VGND_c_1467_n 0.00383152f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_414 N_A_27_74#_c_312_n N_VGND_c_1471_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_415 N_A_27_74#_c_315_n N_VGND_c_1472_n 0.00749631f $X=1.2 $Y=0.515 $X2=0
+ $Y2=0
cc_416 N_A_27_74#_M1011_g N_VGND_c_1488_n 0.0075754f $X=1.845 $Y=0.74 $X2=0
+ $Y2=0
cc_417 N_A_27_74#_M1015_g N_VGND_c_1488_n 0.0075754f $X=2.275 $Y=0.74 $X2=0
+ $Y2=0
cc_418 N_A_27_74#_M1018_g N_VGND_c_1488_n 0.00820284f $X=2.705 $Y=0.74 $X2=0
+ $Y2=0
cc_419 N_A_27_74#_M1026_g N_VGND_c_1488_n 0.0075754f $X=3.135 $Y=0.74 $X2=0
+ $Y2=0
cc_420 N_A_27_74#_M1048_g N_VGND_c_1488_n 0.00820718f $X=3.635 $Y=0.74 $X2=0
+ $Y2=0
cc_421 N_A_27_74#_M1049_g N_VGND_c_1488_n 0.0075754f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_422 N_A_27_74#_c_312_n N_VGND_c_1488_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_423 N_A_27_74#_c_315_n N_VGND_c_1488_n 0.0062048f $X=1.2 $Y=0.515 $X2=0 $Y2=0
cc_424 N_A_384_74#_c_571_n N_VPWR_M1016_s 0.00165831f $X=2.84 $Y=1.885 $X2=0
+ $Y2=0
cc_425 N_A_384_74#_c_574_n N_VPWR_M1025_s 0.00165831f $X=3.74 $Y=1.885 $X2=0
+ $Y2=0
cc_426 N_A_384_74#_c_570_n N_VPWR_c_975_n 0.0216642f $X=2.105 $Y=1.985 $X2=0
+ $Y2=0
cc_427 N_A_384_74#_c_570_n N_VPWR_c_976_n 0.0283117f $X=2.105 $Y=1.985 $X2=0
+ $Y2=0
cc_428 N_A_384_74#_c_571_n N_VPWR_c_976_n 0.0126919f $X=2.84 $Y=1.885 $X2=0
+ $Y2=0
cc_429 N_A_384_74#_c_573_n N_VPWR_c_976_n 0.0283117f $X=3.005 $Y=1.985 $X2=0
+ $Y2=0
cc_430 N_A_384_74#_c_573_n N_VPWR_c_977_n 0.0283117f $X=3.005 $Y=1.985 $X2=0
+ $Y2=0
cc_431 N_A_384_74#_c_574_n N_VPWR_c_977_n 0.0126919f $X=3.74 $Y=1.885 $X2=0
+ $Y2=0
cc_432 N_A_384_74#_c_576_n N_VPWR_c_977_n 0.0283117f $X=3.905 $Y=1.985 $X2=0
+ $Y2=0
cc_433 N_A_384_74#_M1004_g N_VPWR_c_978_n 0.0027763f $X=4.58 $Y=2.4 $X2=0 $Y2=0
cc_434 N_A_384_74#_c_543_n N_VPWR_c_978_n 0.0116873f $X=3.905 $Y=1.97 $X2=0
+ $Y2=0
cc_435 N_A_384_74#_c_576_n N_VPWR_c_978_n 0.033414f $X=3.905 $Y=1.985 $X2=0
+ $Y2=0
cc_436 N_A_384_74#_c_545_n N_VPWR_c_978_n 0.00504465f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_437 N_A_384_74#_M1006_g N_VPWR_c_979_n 0.0030956f $X=5.03 $Y=2.4 $X2=0 $Y2=0
cc_438 N_A_384_74#_M1008_g N_VPWR_c_979_n 0.00307652f $X=5.48 $Y=2.4 $X2=0 $Y2=0
cc_439 N_A_384_74#_c_545_n N_VPWR_c_979_n 7.18372e-19 $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_440 N_A_384_74#_c_546_n N_VPWR_c_979_n 0.00954925f $X=5.175 $Y=1.465 $X2=0
+ $Y2=0
cc_441 N_A_384_74#_c_553_n N_VPWR_c_979_n 4.45097e-19 $X=11.48 $Y=1.465 $X2=0
+ $Y2=0
cc_442 N_A_384_74#_M1010_g N_VPWR_c_980_n 0.0030956f $X=5.93 $Y=2.4 $X2=0 $Y2=0
cc_443 N_A_384_74#_M1012_g N_VPWR_c_980_n 0.00308294f $X=6.38 $Y=2.4 $X2=0 $Y2=0
cc_444 N_A_384_74#_c_545_n N_VPWR_c_980_n 6.09205e-19 $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_445 N_A_384_74#_c_547_n N_VPWR_c_980_n 0.0113635f $X=6.065 $Y=1.465 $X2=0
+ $Y2=0
cc_446 N_A_384_74#_c_553_n N_VPWR_c_980_n 4.47117e-19 $X=11.48 $Y=1.465 $X2=0
+ $Y2=0
cc_447 N_A_384_74#_M1014_g N_VPWR_c_981_n 0.0030956f $X=6.83 $Y=2.4 $X2=0 $Y2=0
cc_448 N_A_384_74#_M1017_g N_VPWR_c_981_n 0.0030956f $X=7.28 $Y=2.4 $X2=0 $Y2=0
cc_449 N_A_384_74#_c_545_n N_VPWR_c_981_n 5.65539e-19 $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_450 N_A_384_74#_c_548_n N_VPWR_c_981_n 0.0119865f $X=7.005 $Y=1.465 $X2=0
+ $Y2=0
cc_451 N_A_384_74#_c_553_n N_VPWR_c_981_n 4.47791e-19 $X=11.48 $Y=1.465 $X2=0
+ $Y2=0
cc_452 N_A_384_74#_M1017_g N_VPWR_c_982_n 0.005209f $X=7.28 $Y=2.4 $X2=0 $Y2=0
cc_453 N_A_384_74#_M1020_g N_VPWR_c_982_n 0.005209f $X=7.73 $Y=2.4 $X2=0 $Y2=0
cc_454 N_A_384_74#_M1020_g N_VPWR_c_983_n 0.0030956f $X=7.73 $Y=2.4 $X2=0 $Y2=0
cc_455 N_A_384_74#_M1024_g N_VPWR_c_983_n 0.00310967f $X=8.18 $Y=2.4 $X2=0 $Y2=0
cc_456 N_A_384_74#_c_545_n N_VPWR_c_983_n 5.65539e-19 $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_457 N_A_384_74#_c_549_n N_VPWR_c_983_n 0.0119865f $X=7.925 $Y=1.465 $X2=0
+ $Y2=0
cc_458 N_A_384_74#_c_553_n N_VPWR_c_983_n 4.47791e-19 $X=11.48 $Y=1.465 $X2=0
+ $Y2=0
cc_459 N_A_384_74#_M1030_g N_VPWR_c_984_n 0.00333991f $X=8.63 $Y=2.4 $X2=0 $Y2=0
cc_460 N_A_384_74#_M1031_g N_VPWR_c_984_n 0.00335915f $X=9.13 $Y=2.4 $X2=0 $Y2=0
cc_461 N_A_384_74#_c_545_n N_VPWR_c_984_n 7.50685e-19 $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_462 N_A_384_74#_c_550_n N_VPWR_c_984_n 0.0158923f $X=8.85 $Y=1.465 $X2=0
+ $Y2=0
cc_463 N_A_384_74#_c_553_n N_VPWR_c_984_n 6.96563e-19 $X=11.48 $Y=1.465 $X2=0
+ $Y2=0
cc_464 N_A_384_74#_M1034_g N_VPWR_c_985_n 0.00336509f $X=9.58 $Y=2.4 $X2=0 $Y2=0
cc_465 N_A_384_74#_M1037_g N_VPWR_c_985_n 0.00340432f $X=10.08 $Y=2.4 $X2=0
+ $Y2=0
cc_466 N_A_384_74#_c_545_n N_VPWR_c_985_n 8.28015e-19 $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_467 N_A_384_74#_c_551_n N_VPWR_c_985_n 0.0158923f $X=9.78 $Y=1.465 $X2=0
+ $Y2=0
cc_468 N_A_384_74#_c_553_n N_VPWR_c_985_n 6.96563e-19 $X=11.48 $Y=1.465 $X2=0
+ $Y2=0
cc_469 N_A_384_74#_M1040_g N_VPWR_c_986_n 0.00324453f $X=10.53 $Y=2.4 $X2=0
+ $Y2=0
cc_470 N_A_384_74#_M1043_g N_VPWR_c_986_n 0.00340385f $X=10.99 $Y=2.4 $X2=0
+ $Y2=0
cc_471 N_A_384_74#_c_545_n N_VPWR_c_986_n 6.194e-19 $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_472 N_A_384_74#_c_552_n N_VPWR_c_986_n 0.0140801f $X=10.71 $Y=1.465 $X2=0
+ $Y2=0
cc_473 N_A_384_74#_c_553_n N_VPWR_c_986_n 4.97545e-19 $X=11.48 $Y=1.465 $X2=0
+ $Y2=0
cc_474 N_A_384_74#_M1045_g N_VPWR_c_988_n 0.00649215f $X=11.48 $Y=2.4 $X2=0
+ $Y2=0
cc_475 N_A_384_74#_c_570_n N_VPWR_c_991_n 0.0145221f $X=2.105 $Y=1.985 $X2=0
+ $Y2=0
cc_476 N_A_384_74#_c_573_n N_VPWR_c_993_n 0.0144623f $X=3.005 $Y=1.985 $X2=0
+ $Y2=0
cc_477 N_A_384_74#_c_576_n N_VPWR_c_995_n 0.0144623f $X=3.905 $Y=1.985 $X2=0
+ $Y2=0
cc_478 N_A_384_74#_M1004_g N_VPWR_c_997_n 0.005209f $X=4.58 $Y=2.4 $X2=0 $Y2=0
cc_479 N_A_384_74#_M1006_g N_VPWR_c_997_n 0.005209f $X=5.03 $Y=2.4 $X2=0 $Y2=0
cc_480 N_A_384_74#_M1008_g N_VPWR_c_999_n 0.005209f $X=5.48 $Y=2.4 $X2=0 $Y2=0
cc_481 N_A_384_74#_M1010_g N_VPWR_c_999_n 0.005209f $X=5.93 $Y=2.4 $X2=0 $Y2=0
cc_482 N_A_384_74#_M1012_g N_VPWR_c_1001_n 0.005209f $X=6.38 $Y=2.4 $X2=0 $Y2=0
cc_483 N_A_384_74#_M1014_g N_VPWR_c_1001_n 0.005209f $X=6.83 $Y=2.4 $X2=0 $Y2=0
cc_484 N_A_384_74#_M1024_g N_VPWR_c_1003_n 0.005209f $X=8.18 $Y=2.4 $X2=0 $Y2=0
cc_485 N_A_384_74#_M1030_g N_VPWR_c_1003_n 0.005209f $X=8.63 $Y=2.4 $X2=0 $Y2=0
cc_486 N_A_384_74#_M1031_g N_VPWR_c_1004_n 0.005209f $X=9.13 $Y=2.4 $X2=0 $Y2=0
cc_487 N_A_384_74#_M1034_g N_VPWR_c_1004_n 0.005209f $X=9.58 $Y=2.4 $X2=0 $Y2=0
cc_488 N_A_384_74#_M1037_g N_VPWR_c_1005_n 0.005209f $X=10.08 $Y=2.4 $X2=0 $Y2=0
cc_489 N_A_384_74#_M1040_g N_VPWR_c_1005_n 0.005209f $X=10.53 $Y=2.4 $X2=0 $Y2=0
cc_490 N_A_384_74#_M1043_g N_VPWR_c_1006_n 0.00553757f $X=10.99 $Y=2.4 $X2=0
+ $Y2=0
cc_491 N_A_384_74#_M1045_g N_VPWR_c_1006_n 0.005209f $X=11.48 $Y=2.4 $X2=0 $Y2=0
cc_492 N_A_384_74#_M1004_g N_VPWR_c_973_n 0.00982376f $X=4.58 $Y=2.4 $X2=0 $Y2=0
cc_493 N_A_384_74#_M1006_g N_VPWR_c_973_n 0.00982266f $X=5.03 $Y=2.4 $X2=0 $Y2=0
cc_494 N_A_384_74#_M1008_g N_VPWR_c_973_n 0.00982266f $X=5.48 $Y=2.4 $X2=0 $Y2=0
cc_495 N_A_384_74#_M1010_g N_VPWR_c_973_n 0.00982266f $X=5.93 $Y=2.4 $X2=0 $Y2=0
cc_496 N_A_384_74#_M1012_g N_VPWR_c_973_n 0.00982266f $X=6.38 $Y=2.4 $X2=0 $Y2=0
cc_497 N_A_384_74#_M1014_g N_VPWR_c_973_n 0.00982266f $X=6.83 $Y=2.4 $X2=0 $Y2=0
cc_498 N_A_384_74#_M1017_g N_VPWR_c_973_n 0.00982266f $X=7.28 $Y=2.4 $X2=0 $Y2=0
cc_499 N_A_384_74#_M1020_g N_VPWR_c_973_n 0.00982266f $X=7.73 $Y=2.4 $X2=0 $Y2=0
cc_500 N_A_384_74#_M1024_g N_VPWR_c_973_n 0.00982266f $X=8.18 $Y=2.4 $X2=0 $Y2=0
cc_501 N_A_384_74#_M1030_g N_VPWR_c_973_n 0.00982754f $X=8.63 $Y=2.4 $X2=0 $Y2=0
cc_502 N_A_384_74#_M1031_g N_VPWR_c_973_n 0.00982642f $X=9.13 $Y=2.4 $X2=0 $Y2=0
cc_503 N_A_384_74#_M1034_g N_VPWR_c_973_n 0.00982754f $X=9.58 $Y=2.4 $X2=0 $Y2=0
cc_504 N_A_384_74#_M1037_g N_VPWR_c_973_n 0.00982418f $X=10.08 $Y=2.4 $X2=0
+ $Y2=0
cc_505 N_A_384_74#_M1040_g N_VPWR_c_973_n 0.00982367f $X=10.53 $Y=2.4 $X2=0
+ $Y2=0
cc_506 N_A_384_74#_M1043_g N_VPWR_c_973_n 0.0108837f $X=10.99 $Y=2.4 $X2=0 $Y2=0
cc_507 N_A_384_74#_M1045_g N_VPWR_c_973_n 0.00986453f $X=11.48 $Y=2.4 $X2=0
+ $Y2=0
cc_508 N_A_384_74#_c_570_n N_VPWR_c_973_n 0.0119308f $X=2.105 $Y=1.985 $X2=0
+ $Y2=0
cc_509 N_A_384_74#_c_573_n N_VPWR_c_973_n 0.0118344f $X=3.005 $Y=1.985 $X2=0
+ $Y2=0
cc_510 N_A_384_74#_c_576_n N_VPWR_c_973_n 0.0118344f $X=3.905 $Y=1.985 $X2=0
+ $Y2=0
cc_511 N_A_384_74#_M1003_g N_Y_c_1195_n 0.0138189f $X=4.565 $Y=0.74 $X2=0 $Y2=0
cc_512 N_A_384_74#_M1004_g N_Y_c_1195_n 0.00621993f $X=4.58 $Y=2.4 $X2=0 $Y2=0
cc_513 N_A_384_74#_M1007_g N_Y_c_1195_n 0.00296452f $X=4.995 $Y=0.74 $X2=0 $Y2=0
cc_514 N_A_384_74#_M1006_g N_Y_c_1195_n 0.00250389f $X=5.03 $Y=2.4 $X2=0 $Y2=0
cc_515 N_A_384_74#_c_543_n N_Y_c_1195_n 0.0375214f $X=3.905 $Y=1.97 $X2=0 $Y2=0
cc_516 N_A_384_74#_c_545_n N_Y_c_1195_n 0.0304042f $X=10.71 $Y=1.665 $X2=0 $Y2=0
cc_517 N_A_384_74#_c_546_n N_Y_c_1195_n 0.0314924f $X=5.175 $Y=1.465 $X2=0 $Y2=0
cc_518 N_A_384_74#_c_553_n N_Y_c_1195_n 0.0189128f $X=11.48 $Y=1.465 $X2=0 $Y2=0
cc_519 N_A_384_74#_M1006_g N_Y_c_1196_n 7.04819e-19 $X=5.03 $Y=2.4 $X2=0 $Y2=0
cc_520 N_A_384_74#_M1013_g N_Y_c_1196_n 0.00318673f $X=5.425 $Y=0.74 $X2=0 $Y2=0
cc_521 N_A_384_74#_M1008_g N_Y_c_1196_n 0.0064289f $X=5.48 $Y=2.4 $X2=0 $Y2=0
cc_522 N_A_384_74#_M1021_g N_Y_c_1196_n 0.00511263f $X=5.855 $Y=0.74 $X2=0 $Y2=0
cc_523 N_A_384_74#_M1010_g N_Y_c_1196_n 0.00409885f $X=5.93 $Y=2.4 $X2=0 $Y2=0
cc_524 N_A_384_74#_c_545_n N_Y_c_1196_n 0.0260544f $X=10.71 $Y=1.665 $X2=0 $Y2=0
cc_525 N_A_384_74#_c_546_n N_Y_c_1196_n 0.0263665f $X=5.175 $Y=1.465 $X2=0 $Y2=0
cc_526 N_A_384_74#_c_547_n N_Y_c_1196_n 0.0307287f $X=6.065 $Y=1.465 $X2=0 $Y2=0
cc_527 N_A_384_74#_c_553_n N_Y_c_1196_n 0.0193844f $X=11.48 $Y=1.465 $X2=0 $Y2=0
cc_528 N_A_384_74#_M1021_g N_Y_c_1197_n 0.00109749f $X=5.855 $Y=0.74 $X2=0 $Y2=0
cc_529 N_A_384_74#_M1010_g N_Y_c_1197_n 0.00106191f $X=5.93 $Y=2.4 $X2=0 $Y2=0
cc_530 N_A_384_74#_M1022_g N_Y_c_1197_n 0.0131322f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_531 N_A_384_74#_M1012_g N_Y_c_1197_n 0.00632482f $X=6.38 $Y=2.4 $X2=0 $Y2=0
cc_532 N_A_384_74#_M1023_g N_Y_c_1197_n 0.00519497f $X=6.785 $Y=0.74 $X2=0 $Y2=0
cc_533 N_A_384_74#_M1014_g N_Y_c_1197_n 0.00436893f $X=6.83 $Y=2.4 $X2=0 $Y2=0
cc_534 N_A_384_74#_c_545_n N_Y_c_1197_n 0.0280183f $X=10.71 $Y=1.665 $X2=0 $Y2=0
cc_535 N_A_384_74#_c_547_n N_Y_c_1197_n 0.0286581f $X=6.065 $Y=1.465 $X2=0 $Y2=0
cc_536 N_A_384_74#_c_548_n N_Y_c_1197_n 0.0293313f $X=7.005 $Y=1.465 $X2=0 $Y2=0
cc_537 N_A_384_74#_c_553_n N_Y_c_1197_n 0.0205921f $X=11.48 $Y=1.465 $X2=0 $Y2=0
cc_538 N_A_384_74#_M1023_g N_Y_c_1198_n 0.00110789f $X=6.785 $Y=0.74 $X2=0 $Y2=0
cc_539 N_A_384_74#_M1014_g N_Y_c_1198_n 0.00137539f $X=6.83 $Y=2.4 $X2=0 $Y2=0
cc_540 N_A_384_74#_M1017_g N_Y_c_1198_n 0.00602666f $X=7.28 $Y=2.4 $X2=0 $Y2=0
cc_541 N_A_384_74#_M1027_g N_Y_c_1198_n 0.0137331f $X=7.285 $Y=0.74 $X2=0 $Y2=0
cc_542 N_A_384_74#_M1028_g N_Y_c_1198_n 0.0052341f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_543 N_A_384_74#_M1020_g N_Y_c_1198_n 0.00287989f $X=7.73 $Y=2.4 $X2=0 $Y2=0
cc_544 N_A_384_74#_c_545_n N_Y_c_1198_n 0.0286676f $X=10.71 $Y=1.665 $X2=0 $Y2=0
cc_545 N_A_384_74#_c_548_n N_Y_c_1198_n 0.0317868f $X=7.005 $Y=1.465 $X2=0 $Y2=0
cc_546 N_A_384_74#_c_549_n N_Y_c_1198_n 0.0309223f $X=7.925 $Y=1.465 $X2=0 $Y2=0
cc_547 N_A_384_74#_c_553_n N_Y_c_1198_n 0.0204645f $X=11.48 $Y=1.465 $X2=0 $Y2=0
cc_548 N_A_384_74#_M1017_g N_Y_c_1207_n 0.0112654f $X=7.28 $Y=2.4 $X2=0 $Y2=0
cc_549 N_A_384_74#_M1020_g N_Y_c_1207_n 0.0112654f $X=7.73 $Y=2.4 $X2=0 $Y2=0
cc_550 N_A_384_74#_M1024_g N_Y_c_1262_n 0.00294766f $X=8.18 $Y=2.4 $X2=0 $Y2=0
cc_551 N_A_384_74#_M1030_g N_Y_c_1262_n 0.00316431f $X=8.63 $Y=2.4 $X2=0 $Y2=0
cc_552 N_A_384_74#_c_545_n N_Y_c_1262_n 0.0011287f $X=10.71 $Y=1.665 $X2=0 $Y2=0
cc_553 N_A_384_74#_M1024_g N_Y_c_1208_n 0.0104099f $X=8.18 $Y=2.4 $X2=0 $Y2=0
cc_554 N_A_384_74#_M1030_g N_Y_c_1208_n 0.0105267f $X=8.63 $Y=2.4 $X2=0 $Y2=0
cc_555 N_A_384_74#_M1028_g N_Y_c_1199_n 0.00111312f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_556 N_A_384_74#_M1020_g N_Y_c_1199_n 9.03138e-19 $X=7.73 $Y=2.4 $X2=0 $Y2=0
cc_557 N_A_384_74#_M1024_g N_Y_c_1199_n 0.00565525f $X=8.18 $Y=2.4 $X2=0 $Y2=0
cc_558 N_A_384_74#_M1032_g N_Y_c_1199_n 0.0140323f $X=8.215 $Y=0.74 $X2=0 $Y2=0
cc_559 N_A_384_74#_M1030_g N_Y_c_1199_n 0.00303955f $X=8.63 $Y=2.4 $X2=0 $Y2=0
cc_560 N_A_384_74#_M1036_g N_Y_c_1199_n 0.0052532f $X=8.645 $Y=0.74 $X2=0 $Y2=0
cc_561 N_A_384_74#_c_545_n N_Y_c_1199_n 0.029145f $X=10.71 $Y=1.665 $X2=0 $Y2=0
cc_562 N_A_384_74#_c_549_n N_Y_c_1199_n 0.0309801f $X=7.925 $Y=1.465 $X2=0 $Y2=0
cc_563 N_A_384_74#_c_550_n N_Y_c_1199_n 0.0317874f $X=8.85 $Y=1.465 $X2=0 $Y2=0
cc_564 N_A_384_74#_c_553_n N_Y_c_1199_n 0.020647f $X=11.48 $Y=1.465 $X2=0 $Y2=0
cc_565 N_A_384_74#_M1031_g N_Y_c_1277_n 0.00254641f $X=9.13 $Y=2.4 $X2=0 $Y2=0
cc_566 N_A_384_74#_M1034_g N_Y_c_1277_n 0.00316431f $X=9.58 $Y=2.4 $X2=0 $Y2=0
cc_567 N_A_384_74#_c_545_n N_Y_c_1277_n 9.68436e-19 $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_568 N_A_384_74#_M1031_g N_Y_c_1210_n 0.0104335f $X=9.13 $Y=2.4 $X2=0 $Y2=0
cc_569 N_A_384_74#_M1034_g N_Y_c_1210_n 0.0105267f $X=9.58 $Y=2.4 $X2=0 $Y2=0
cc_570 N_A_384_74#_M1030_g N_Y_c_1200_n 9.03726e-19 $X=8.63 $Y=2.4 $X2=0 $Y2=0
cc_571 N_A_384_74#_M1036_g N_Y_c_1200_n 0.00111312f $X=8.645 $Y=0.74 $X2=0 $Y2=0
cc_572 N_A_384_74#_M1031_g N_Y_c_1200_n 0.00609125f $X=9.13 $Y=2.4 $X2=0 $Y2=0
cc_573 N_A_384_74#_M1038_g N_Y_c_1200_n 0.0140323f $X=9.145 $Y=0.74 $X2=0 $Y2=0
cc_574 N_A_384_74#_M1034_g N_Y_c_1200_n 0.00293186f $X=9.58 $Y=2.4 $X2=0 $Y2=0
cc_575 N_A_384_74#_M1039_g N_Y_c_1200_n 0.0052532f $X=9.575 $Y=0.74 $X2=0 $Y2=0
cc_576 N_A_384_74#_c_545_n N_Y_c_1200_n 0.0291963f $X=10.71 $Y=1.665 $X2=0 $Y2=0
cc_577 N_A_384_74#_c_550_n N_Y_c_1200_n 0.0301915f $X=8.85 $Y=1.465 $X2=0 $Y2=0
cc_578 N_A_384_74#_c_551_n N_Y_c_1200_n 0.0317874f $X=9.78 $Y=1.465 $X2=0 $Y2=0
cc_579 N_A_384_74#_c_553_n N_Y_c_1200_n 0.0206962f $X=11.48 $Y=1.465 $X2=0 $Y2=0
cc_580 N_A_384_74#_M1034_g N_Y_c_1201_n 9.96342e-19 $X=9.58 $Y=2.4 $X2=0 $Y2=0
cc_581 N_A_384_74#_M1039_g N_Y_c_1201_n 0.00111312f $X=9.575 $Y=0.74 $X2=0 $Y2=0
cc_582 N_A_384_74#_M1037_g N_Y_c_1201_n 0.00640933f $X=10.08 $Y=2.4 $X2=0 $Y2=0
cc_583 N_A_384_74#_M1041_g N_Y_c_1201_n 0.0140323f $X=10.075 $Y=0.74 $X2=0 $Y2=0
cc_584 N_A_384_74#_M1042_g N_Y_c_1201_n 0.0052532f $X=10.505 $Y=0.74 $X2=0 $Y2=0
cc_585 N_A_384_74#_M1040_g N_Y_c_1201_n 0.0045289f $X=10.53 $Y=2.4 $X2=0 $Y2=0
cc_586 N_A_384_74#_c_545_n N_Y_c_1201_n 0.0291468f $X=10.71 $Y=1.665 $X2=0 $Y2=0
cc_587 N_A_384_74#_c_551_n N_Y_c_1201_n 0.0301915f $X=9.78 $Y=1.465 $X2=0 $Y2=0
cc_588 N_A_384_74#_c_552_n N_Y_c_1201_n 0.0317874f $X=10.71 $Y=1.465 $X2=0 $Y2=0
cc_589 N_A_384_74#_c_553_n N_Y_c_1201_n 0.0207067f $X=11.48 $Y=1.465 $X2=0 $Y2=0
cc_590 N_A_384_74#_M1042_g N_Y_c_1202_n 0.00110862f $X=10.505 $Y=0.74 $X2=0
+ $Y2=0
cc_591 N_A_384_74#_M1040_g N_Y_c_1202_n 8.52524e-19 $X=10.53 $Y=2.4 $X2=0 $Y2=0
cc_592 N_A_384_74#_M1043_g N_Y_c_1202_n 0.0034752f $X=10.99 $Y=2.4 $X2=0 $Y2=0
cc_593 N_A_384_74#_M1044_g N_Y_c_1202_n 0.01491f $X=11.005 $Y=0.74 $X2=0 $Y2=0
cc_594 N_A_384_74#_M1046_g N_Y_c_1202_n 0.0190845f $X=11.435 $Y=0.74 $X2=0 $Y2=0
cc_595 N_A_384_74#_M1045_g N_Y_c_1202_n 0.00469386f $X=11.48 $Y=2.4 $X2=0 $Y2=0
cc_596 N_A_384_74#_c_545_n N_Y_c_1202_n 0.0028814f $X=10.71 $Y=1.665 $X2=0 $Y2=0
cc_597 N_A_384_74#_c_552_n N_Y_c_1202_n 0.0313214f $X=10.71 $Y=1.465 $X2=0 $Y2=0
cc_598 N_A_384_74#_c_553_n N_Y_c_1202_n 0.0344515f $X=11.48 $Y=1.465 $X2=0 $Y2=0
cc_599 N_A_384_74#_M1004_g N_Y_c_1311_n 0.00254862f $X=4.58 $Y=2.4 $X2=0 $Y2=0
cc_600 N_A_384_74#_M1006_g N_Y_c_1311_n 0.00152964f $X=5.03 $Y=2.4 $X2=0 $Y2=0
cc_601 N_A_384_74#_c_545_n N_Y_c_1311_n 0.00110327f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_602 N_A_384_74#_M1008_g N_Y_c_1314_n 0.00169254f $X=5.48 $Y=2.4 $X2=0 $Y2=0
cc_603 N_A_384_74#_M1010_g N_Y_c_1314_n 0.00152964f $X=5.93 $Y=2.4 $X2=0 $Y2=0
cc_604 N_A_384_74#_c_545_n N_Y_c_1314_n 0.00141259f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_605 N_A_384_74#_c_553_n N_Y_c_1314_n 6.6154e-19 $X=11.48 $Y=1.465 $X2=0 $Y2=0
cc_606 N_A_384_74#_M1012_g N_Y_c_1318_n 0.00140803f $X=6.38 $Y=2.4 $X2=0 $Y2=0
cc_607 N_A_384_74#_M1014_g N_Y_c_1318_n 0.00152964f $X=6.83 $Y=2.4 $X2=0 $Y2=0
cc_608 N_A_384_74#_c_545_n N_Y_c_1318_n 0.0011806f $X=10.71 $Y=1.665 $X2=0 $Y2=0
cc_609 N_A_384_74#_M1037_g N_Y_c_1321_n 0.00124236f $X=10.08 $Y=2.4 $X2=0 $Y2=0
cc_610 N_A_384_74#_M1040_g N_Y_c_1321_n 0.00152964f $X=10.53 $Y=2.4 $X2=0 $Y2=0
cc_611 N_A_384_74#_c_545_n N_Y_c_1321_n 0.00102594f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_612 N_A_384_74#_M1043_g N_Y_c_1214_n 0.0044513f $X=10.99 $Y=2.4 $X2=0 $Y2=0
cc_613 N_A_384_74#_M1045_g N_Y_c_1214_n 0.00599049f $X=11.48 $Y=2.4 $X2=0 $Y2=0
cc_614 N_A_384_74#_M1004_g N_Y_c_1215_n 0.0122453f $X=4.58 $Y=2.4 $X2=0 $Y2=0
cc_615 N_A_384_74#_M1006_g N_Y_c_1215_n 0.0118259f $X=5.03 $Y=2.4 $X2=0 $Y2=0
cc_616 N_A_384_74#_M1008_g N_Y_c_1216_n 0.0118259f $X=5.48 $Y=2.4 $X2=0 $Y2=0
cc_617 N_A_384_74#_M1010_g N_Y_c_1216_n 0.0118259f $X=5.93 $Y=2.4 $X2=0 $Y2=0
cc_618 N_A_384_74#_M1012_g N_Y_c_1217_n 0.0118259f $X=6.38 $Y=2.4 $X2=0 $Y2=0
cc_619 N_A_384_74#_M1014_g N_Y_c_1217_n 0.0118259f $X=6.83 $Y=2.4 $X2=0 $Y2=0
cc_620 N_A_384_74#_M1037_g N_Y_c_1218_n 0.0115839f $X=10.08 $Y=2.4 $X2=0 $Y2=0
cc_621 N_A_384_74#_M1040_g N_Y_c_1218_n 0.0118428f $X=10.53 $Y=2.4 $X2=0 $Y2=0
cc_622 N_A_384_74#_M1043_g N_Y_c_1219_n 6.71238e-19 $X=10.99 $Y=2.4 $X2=0 $Y2=0
cc_623 N_A_384_74#_M1045_g N_Y_c_1219_n 0.0130656f $X=11.48 $Y=2.4 $X2=0 $Y2=0
cc_624 N_A_384_74#_M1006_g N_Y_c_1336_n 0.00775616f $X=5.03 $Y=2.4 $X2=0 $Y2=0
cc_625 N_A_384_74#_M1008_g N_Y_c_1336_n 0.00750888f $X=5.48 $Y=2.4 $X2=0 $Y2=0
cc_626 N_A_384_74#_M1010_g N_Y_c_1336_n 0.00763665f $X=5.93 $Y=2.4 $X2=0 $Y2=0
cc_627 N_A_384_74#_M1012_g N_Y_c_1336_n 0.00759682f $X=6.38 $Y=2.4 $X2=0 $Y2=0
cc_628 N_A_384_74#_M1014_g N_Y_c_1336_n 0.00777323f $X=6.83 $Y=2.4 $X2=0 $Y2=0
cc_629 N_A_384_74#_M1017_g N_Y_c_1336_n 0.00779332f $X=7.28 $Y=2.4 $X2=0 $Y2=0
cc_630 N_A_384_74#_M1020_g N_Y_c_1336_n 0.00784152f $X=7.73 $Y=2.4 $X2=0 $Y2=0
cc_631 N_A_384_74#_M1024_g N_Y_c_1336_n 0.00794076f $X=8.18 $Y=2.4 $X2=0 $Y2=0
cc_632 N_A_384_74#_M1030_g N_Y_c_1336_n 0.00786325f $X=8.63 $Y=2.4 $X2=0 $Y2=0
cc_633 N_A_384_74#_M1031_g N_Y_c_1336_n 0.00776487f $X=9.13 $Y=2.4 $X2=0 $Y2=0
cc_634 N_A_384_74#_M1034_g N_Y_c_1336_n 0.00779496f $X=9.58 $Y=2.4 $X2=0 $Y2=0
cc_635 N_A_384_74#_M1037_g N_Y_c_1336_n 0.00764079f $X=10.08 $Y=2.4 $X2=0 $Y2=0
cc_636 N_A_384_74#_M1040_g N_Y_c_1336_n 0.0077903f $X=10.53 $Y=2.4 $X2=0 $Y2=0
cc_637 N_A_384_74#_M1043_g N_Y_c_1336_n 0.0143268f $X=10.99 $Y=2.4 $X2=0 $Y2=0
cc_638 N_A_384_74#_c_545_n N_Y_c_1336_n 0.60514f $X=10.71 $Y=1.665 $X2=0 $Y2=0
cc_639 N_A_384_74#_c_546_n N_Y_c_1336_n 0.00187712f $X=5.175 $Y=1.465 $X2=0
+ $Y2=0
cc_640 N_A_384_74#_c_547_n N_Y_c_1336_n 0.00247972f $X=6.065 $Y=1.465 $X2=0
+ $Y2=0
cc_641 N_A_384_74#_c_548_n N_Y_c_1336_n 0.0020405f $X=7.005 $Y=1.465 $X2=0 $Y2=0
cc_642 N_A_384_74#_c_549_n N_Y_c_1336_n 0.00185369f $X=7.925 $Y=1.465 $X2=0
+ $Y2=0
cc_643 N_A_384_74#_c_550_n N_Y_c_1336_n 0.00128761f $X=8.85 $Y=1.465 $X2=0 $Y2=0
cc_644 N_A_384_74#_c_551_n N_Y_c_1336_n 0.00147955f $X=9.78 $Y=1.465 $X2=0 $Y2=0
cc_645 N_A_384_74#_c_552_n N_Y_c_1336_n 0.0019243f $X=10.71 $Y=1.465 $X2=0 $Y2=0
cc_646 N_A_384_74#_M1017_g N_Y_c_1358_n 0.00142298f $X=7.28 $Y=2.4 $X2=0 $Y2=0
cc_647 N_A_384_74#_M1020_g N_Y_c_1358_n 0.00209021f $X=7.73 $Y=2.4 $X2=0 $Y2=0
cc_648 N_A_384_74#_c_545_n N_Y_c_1358_n 9.48608e-19 $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_649 N_A_384_74#_c_538_n N_VGND_M1015_s 0.00176461f $X=2.755 $Y=1.045 $X2=0
+ $Y2=0
cc_650 N_A_384_74#_c_541_n N_VGND_M1026_s 0.00250873f $X=3.685 $Y=1.045 $X2=0
+ $Y2=0
cc_651 N_A_384_74#_c_537_n N_VGND_c_1450_n 0.0182488f $X=2.06 $Y=0.515 $X2=0
+ $Y2=0
cc_652 N_A_384_74#_c_537_n N_VGND_c_1451_n 0.0157999f $X=2.06 $Y=0.515 $X2=0
+ $Y2=0
cc_653 N_A_384_74#_c_538_n N_VGND_c_1451_n 0.0152916f $X=2.755 $Y=1.045 $X2=0
+ $Y2=0
cc_654 N_A_384_74#_c_540_n N_VGND_c_1451_n 0.0158413f $X=2.92 $Y=0.515 $X2=0
+ $Y2=0
cc_655 N_A_384_74#_c_540_n N_VGND_c_1452_n 0.0164981f $X=2.92 $Y=0.515 $X2=0
+ $Y2=0
cc_656 N_A_384_74#_c_541_n N_VGND_c_1452_n 0.0209867f $X=3.685 $Y=1.045 $X2=0
+ $Y2=0
cc_657 N_A_384_74#_c_542_n N_VGND_c_1452_n 0.0166127f $X=3.85 $Y=0.515 $X2=0
+ $Y2=0
cc_658 N_A_384_74#_M1003_g N_VGND_c_1453_n 0.00581358f $X=4.565 $Y=0.74 $X2=0
+ $Y2=0
cc_659 N_A_384_74#_c_542_n N_VGND_c_1453_n 0.0225912f $X=3.85 $Y=0.515 $X2=0
+ $Y2=0
cc_660 N_A_384_74#_c_543_n N_VGND_c_1453_n 0.0342051f $X=3.905 $Y=1.97 $X2=0
+ $Y2=0
cc_661 N_A_384_74#_c_545_n N_VGND_c_1453_n 0.00177399f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_662 N_A_384_74#_M1003_g N_VGND_c_1454_n 5.98876e-19 $X=4.565 $Y=0.74 $X2=0
+ $Y2=0
cc_663 N_A_384_74#_M1007_g N_VGND_c_1454_n 0.0121668f $X=4.995 $Y=0.74 $X2=0
+ $Y2=0
cc_664 N_A_384_74#_M1013_g N_VGND_c_1454_n 0.00174374f $X=5.425 $Y=0.74 $X2=0
+ $Y2=0
cc_665 N_A_384_74#_c_545_n N_VGND_c_1454_n 0.00123706f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_666 N_A_384_74#_c_546_n N_VGND_c_1454_n 0.0155643f $X=5.175 $Y=1.465 $X2=0
+ $Y2=0
cc_667 N_A_384_74#_c_553_n N_VGND_c_1454_n 7.7342e-19 $X=11.48 $Y=1.465 $X2=0
+ $Y2=0
cc_668 N_A_384_74#_M1013_g N_VGND_c_1455_n 5.61948e-19 $X=5.425 $Y=0.74 $X2=0
+ $Y2=0
cc_669 N_A_384_74#_M1021_g N_VGND_c_1455_n 0.0126669f $X=5.855 $Y=0.74 $X2=0
+ $Y2=0
cc_670 N_A_384_74#_M1022_g N_VGND_c_1455_n 0.00562547f $X=6.355 $Y=0.74 $X2=0
+ $Y2=0
cc_671 N_A_384_74#_c_545_n N_VGND_c_1455_n 0.00181192f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_672 N_A_384_74#_c_547_n N_VGND_c_1455_n 0.0207506f $X=6.065 $Y=1.465 $X2=0
+ $Y2=0
cc_673 N_A_384_74#_c_553_n N_VGND_c_1455_n 0.00131438f $X=11.48 $Y=1.465 $X2=0
+ $Y2=0
cc_674 N_A_384_74#_M1022_g N_VGND_c_1456_n 5.96902e-19 $X=6.355 $Y=0.74 $X2=0
+ $Y2=0
cc_675 N_A_384_74#_M1023_g N_VGND_c_1456_n 0.0126964f $X=6.785 $Y=0.74 $X2=0
+ $Y2=0
cc_676 N_A_384_74#_M1027_g N_VGND_c_1456_n 0.00562212f $X=7.285 $Y=0.74 $X2=0
+ $Y2=0
cc_677 N_A_384_74#_c_545_n N_VGND_c_1456_n 0.00179414f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_678 N_A_384_74#_c_548_n N_VGND_c_1456_n 0.020583f $X=7.005 $Y=1.465 $X2=0
+ $Y2=0
cc_679 N_A_384_74#_c_553_n N_VGND_c_1456_n 0.00131525f $X=11.48 $Y=1.465 $X2=0
+ $Y2=0
cc_680 N_A_384_74#_M1027_g N_VGND_c_1457_n 5.96902e-19 $X=7.285 $Y=0.74 $X2=0
+ $Y2=0
cc_681 N_A_384_74#_M1028_g N_VGND_c_1457_n 0.0126506f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_682 N_A_384_74#_M1032_g N_VGND_c_1457_n 0.00562044f $X=8.215 $Y=0.74 $X2=0
+ $Y2=0
cc_683 N_A_384_74#_c_545_n N_VGND_c_1457_n 0.00181192f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_684 N_A_384_74#_c_549_n N_VGND_c_1457_n 0.0207506f $X=7.925 $Y=1.465 $X2=0
+ $Y2=0
cc_685 N_A_384_74#_c_553_n N_VGND_c_1457_n 0.00131525f $X=11.48 $Y=1.465 $X2=0
+ $Y2=0
cc_686 N_A_384_74#_M1032_g N_VGND_c_1458_n 5.96902e-19 $X=8.215 $Y=0.74 $X2=0
+ $Y2=0
cc_687 N_A_384_74#_M1036_g N_VGND_c_1458_n 0.0126506f $X=8.645 $Y=0.74 $X2=0
+ $Y2=0
cc_688 N_A_384_74#_M1038_g N_VGND_c_1458_n 0.00562044f $X=9.145 $Y=0.74 $X2=0
+ $Y2=0
cc_689 N_A_384_74#_c_545_n N_VGND_c_1458_n 0.00197911f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_690 N_A_384_74#_c_550_n N_VGND_c_1458_n 0.0205727f $X=8.85 $Y=1.465 $X2=0
+ $Y2=0
cc_691 N_A_384_74#_c_553_n N_VGND_c_1458_n 0.0013196f $X=11.48 $Y=1.465 $X2=0
+ $Y2=0
cc_692 N_A_384_74#_M1038_g N_VGND_c_1459_n 5.96902e-19 $X=9.145 $Y=0.74 $X2=0
+ $Y2=0
cc_693 N_A_384_74#_M1039_g N_VGND_c_1459_n 0.0126506f $X=9.575 $Y=0.74 $X2=0
+ $Y2=0
cc_694 N_A_384_74#_M1041_g N_VGND_c_1459_n 0.00562044f $X=10.075 $Y=0.74 $X2=0
+ $Y2=0
cc_695 N_A_384_74#_c_545_n N_VGND_c_1459_n 0.00197911f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_696 N_A_384_74#_c_551_n N_VGND_c_1459_n 0.0205727f $X=9.78 $Y=1.465 $X2=0
+ $Y2=0
cc_697 N_A_384_74#_c_553_n N_VGND_c_1459_n 0.0013196f $X=11.48 $Y=1.465 $X2=0
+ $Y2=0
cc_698 N_A_384_74#_M1041_g N_VGND_c_1460_n 5.96902e-19 $X=10.075 $Y=0.74 $X2=0
+ $Y2=0
cc_699 N_A_384_74#_M1042_g N_VGND_c_1460_n 0.0126506f $X=10.505 $Y=0.74 $X2=0
+ $Y2=0
cc_700 N_A_384_74#_M1044_g N_VGND_c_1460_n 0.00570988f $X=11.005 $Y=0.74 $X2=0
+ $Y2=0
cc_701 N_A_384_74#_c_545_n N_VGND_c_1460_n 0.00149791f $X=10.71 $Y=1.665 $X2=0
+ $Y2=0
cc_702 N_A_384_74#_c_552_n N_VGND_c_1460_n 0.0206571f $X=10.71 $Y=1.465 $X2=0
+ $Y2=0
cc_703 N_A_384_74#_c_553_n N_VGND_c_1460_n 0.00131612f $X=11.48 $Y=1.465 $X2=0
+ $Y2=0
cc_704 N_A_384_74#_M1046_g N_VGND_c_1462_n 0.0184907f $X=11.435 $Y=0.74 $X2=0
+ $Y2=0
cc_705 N_A_384_74#_c_553_n N_VGND_c_1462_n 6.77396e-19 $X=11.48 $Y=1.465 $X2=0
+ $Y2=0
cc_706 N_A_384_74#_c_537_n N_VGND_c_1463_n 0.00749631f $X=2.06 $Y=0.515 $X2=0
+ $Y2=0
cc_707 N_A_384_74#_c_540_n N_VGND_c_1465_n 0.0109942f $X=2.92 $Y=0.515 $X2=0
+ $Y2=0
cc_708 N_A_384_74#_c_542_n N_VGND_c_1467_n 0.0109942f $X=3.85 $Y=0.515 $X2=0
+ $Y2=0
cc_709 N_A_384_74#_M1003_g N_VGND_c_1469_n 0.00434272f $X=4.565 $Y=0.74 $X2=0
+ $Y2=0
cc_710 N_A_384_74#_M1007_g N_VGND_c_1469_n 0.00383152f $X=4.995 $Y=0.74 $X2=0
+ $Y2=0
cc_711 N_A_384_74#_M1013_g N_VGND_c_1473_n 0.00461464f $X=5.425 $Y=0.74 $X2=0
+ $Y2=0
cc_712 N_A_384_74#_M1021_g N_VGND_c_1473_n 0.00383152f $X=5.855 $Y=0.74 $X2=0
+ $Y2=0
cc_713 N_A_384_74#_M1022_g N_VGND_c_1474_n 0.00451267f $X=6.355 $Y=0.74 $X2=0
+ $Y2=0
cc_714 N_A_384_74#_M1023_g N_VGND_c_1474_n 0.00383152f $X=6.785 $Y=0.74 $X2=0
+ $Y2=0
cc_715 N_A_384_74#_M1027_g N_VGND_c_1475_n 0.00439937f $X=7.285 $Y=0.74 $X2=0
+ $Y2=0
cc_716 N_A_384_74#_M1028_g N_VGND_c_1475_n 0.00383152f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_717 N_A_384_74#_M1032_g N_VGND_c_1476_n 0.00434272f $X=8.215 $Y=0.74 $X2=0
+ $Y2=0
cc_718 N_A_384_74#_M1036_g N_VGND_c_1476_n 0.00383152f $X=8.645 $Y=0.74 $X2=0
+ $Y2=0
cc_719 N_A_384_74#_M1038_g N_VGND_c_1477_n 0.00434272f $X=9.145 $Y=0.74 $X2=0
+ $Y2=0
cc_720 N_A_384_74#_M1039_g N_VGND_c_1477_n 0.00383152f $X=9.575 $Y=0.74 $X2=0
+ $Y2=0
cc_721 N_A_384_74#_M1041_g N_VGND_c_1478_n 0.00434272f $X=10.075 $Y=0.74 $X2=0
+ $Y2=0
cc_722 N_A_384_74#_M1042_g N_VGND_c_1478_n 0.00383152f $X=10.505 $Y=0.74 $X2=0
+ $Y2=0
cc_723 N_A_384_74#_M1044_g N_VGND_c_1479_n 0.00434272f $X=11.005 $Y=0.74 $X2=0
+ $Y2=0
cc_724 N_A_384_74#_M1046_g N_VGND_c_1479_n 0.00434272f $X=11.435 $Y=0.74 $X2=0
+ $Y2=0
cc_725 N_A_384_74#_M1003_g N_VGND_c_1488_n 0.00820772f $X=4.565 $Y=0.74 $X2=0
+ $Y2=0
cc_726 N_A_384_74#_M1007_g N_VGND_c_1488_n 0.0075754f $X=4.995 $Y=0.74 $X2=0
+ $Y2=0
cc_727 N_A_384_74#_M1013_g N_VGND_c_1488_n 0.00908333f $X=5.425 $Y=0.74 $X2=0
+ $Y2=0
cc_728 N_A_384_74#_M1021_g N_VGND_c_1488_n 0.0075754f $X=5.855 $Y=0.74 $X2=0
+ $Y2=0
cc_729 N_A_384_74#_M1022_g N_VGND_c_1488_n 0.00875749f $X=6.355 $Y=0.74 $X2=0
+ $Y2=0
cc_730 N_A_384_74#_M1023_g N_VGND_c_1488_n 0.0075754f $X=6.785 $Y=0.74 $X2=0
+ $Y2=0
cc_731 N_A_384_74#_M1027_g N_VGND_c_1488_n 0.00839062f $X=7.285 $Y=0.74 $X2=0
+ $Y2=0
cc_732 N_A_384_74#_M1028_g N_VGND_c_1488_n 0.0075754f $X=7.715 $Y=0.74 $X2=0
+ $Y2=0
cc_733 N_A_384_74#_M1032_g N_VGND_c_1488_n 0.00820718f $X=8.215 $Y=0.74 $X2=0
+ $Y2=0
cc_734 N_A_384_74#_M1036_g N_VGND_c_1488_n 0.0075754f $X=8.645 $Y=0.74 $X2=0
+ $Y2=0
cc_735 N_A_384_74#_M1038_g N_VGND_c_1488_n 0.00820718f $X=9.145 $Y=0.74 $X2=0
+ $Y2=0
cc_736 N_A_384_74#_M1039_g N_VGND_c_1488_n 0.0075754f $X=9.575 $Y=0.74 $X2=0
+ $Y2=0
cc_737 N_A_384_74#_M1041_g N_VGND_c_1488_n 0.00820718f $X=10.075 $Y=0.74 $X2=0
+ $Y2=0
cc_738 N_A_384_74#_M1042_g N_VGND_c_1488_n 0.0075754f $X=10.505 $Y=0.74 $X2=0
+ $Y2=0
cc_739 N_A_384_74#_M1044_g N_VGND_c_1488_n 0.00820718f $X=11.005 $Y=0.74 $X2=0
+ $Y2=0
cc_740 N_A_384_74#_M1046_g N_VGND_c_1488_n 0.00823934f $X=11.435 $Y=0.74 $X2=0
+ $Y2=0
cc_741 N_A_384_74#_c_537_n N_VGND_c_1488_n 0.0062048f $X=2.06 $Y=0.515 $X2=0
+ $Y2=0
cc_742 N_A_384_74#_c_540_n N_VGND_c_1488_n 0.00904371f $X=2.92 $Y=0.515 $X2=0
+ $Y2=0
cc_743 N_A_384_74#_c_542_n N_VGND_c_1488_n 0.00904371f $X=3.85 $Y=0.515 $X2=0
+ $Y2=0
cc_744 N_VPWR_c_982_n N_Y_c_1207_n 0.0144623f $X=7.87 $Y=3.33 $X2=0 $Y2=0
cc_745 N_VPWR_c_973_n N_Y_c_1207_n 0.0118344f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_746 N_VPWR_c_983_n N_Y_c_1262_n 0.0104268f $X=7.955 $Y=2.085 $X2=0 $Y2=0
cc_747 N_VPWR_c_984_n N_Y_c_1262_n 0.0109606f $X=8.855 $Y=2.085 $X2=0 $Y2=0
cc_748 N_VPWR_c_983_n N_Y_c_1208_n 0.0267962f $X=7.955 $Y=2.085 $X2=0 $Y2=0
cc_749 N_VPWR_c_984_n N_Y_c_1208_n 0.0268239f $X=8.855 $Y=2.085 $X2=0 $Y2=0
cc_750 N_VPWR_c_1003_n N_Y_c_1208_n 0.0144623f $X=8.77 $Y=3.33 $X2=0 $Y2=0
cc_751 N_VPWR_c_973_n N_Y_c_1208_n 0.0118344f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_752 N_VPWR_c_984_n N_Y_c_1277_n 0.0111375f $X=8.855 $Y=2.085 $X2=0 $Y2=0
cc_753 N_VPWR_c_985_n N_Y_c_1277_n 0.0109668f $X=9.805 $Y=2.085 $X2=0 $Y2=0
cc_754 N_VPWR_c_984_n N_Y_c_1210_n 0.0273702f $X=8.855 $Y=2.085 $X2=0 $Y2=0
cc_755 N_VPWR_c_985_n N_Y_c_1210_n 0.0268283f $X=9.805 $Y=2.085 $X2=0 $Y2=0
cc_756 N_VPWR_c_1004_n N_Y_c_1210_n 0.0144623f $X=9.72 $Y=3.33 $X2=0 $Y2=0
cc_757 N_VPWR_c_973_n N_Y_c_1210_n 0.0118344f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_758 N_VPWR_c_979_n N_Y_c_1311_n 0.0376772f $X=5.255 $Y=2.085 $X2=0 $Y2=0
cc_759 N_VPWR_c_979_n N_Y_c_1314_n 0.00502852f $X=5.255 $Y=2.085 $X2=0 $Y2=0
cc_760 N_VPWR_c_980_n N_Y_c_1314_n 0.0376775f $X=6.155 $Y=2.085 $X2=0 $Y2=0
cc_761 N_VPWR_c_980_n N_Y_c_1318_n 0.00472896f $X=6.155 $Y=2.085 $X2=0 $Y2=0
cc_762 N_VPWR_c_981_n N_Y_c_1318_n 0.0376769f $X=7.055 $Y=2.085 $X2=0 $Y2=0
cc_763 N_VPWR_c_985_n N_Y_c_1321_n 0.00504547f $X=9.805 $Y=2.085 $X2=0 $Y2=0
cc_764 N_VPWR_c_986_n N_Y_c_1321_n 0.0377254f $X=10.755 $Y=2.085 $X2=0 $Y2=0
cc_765 N_VPWR_c_986_n N_Y_c_1214_n 0.005042f $X=10.755 $Y=2.085 $X2=0 $Y2=0
cc_766 N_VPWR_c_988_n N_Y_c_1214_n 0.0396382f $X=11.705 $Y=1.985 $X2=0 $Y2=0
cc_767 N_VPWR_c_978_n N_Y_c_1215_n 0.0322322f $X=4.355 $Y=2.085 $X2=0 $Y2=0
cc_768 N_VPWR_c_997_n N_Y_c_1215_n 0.0144623f $X=5.17 $Y=3.33 $X2=0 $Y2=0
cc_769 N_VPWR_c_973_n N_Y_c_1215_n 0.0118344f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_770 N_VPWR_c_979_n N_Y_c_1216_n 0.0334492f $X=5.255 $Y=2.085 $X2=0 $Y2=0
cc_771 N_VPWR_c_999_n N_Y_c_1216_n 0.0144623f $X=6.07 $Y=3.33 $X2=0 $Y2=0
cc_772 N_VPWR_c_973_n N_Y_c_1216_n 0.0118344f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_773 N_VPWR_c_980_n N_Y_c_1217_n 0.0334492f $X=6.155 $Y=2.085 $X2=0 $Y2=0
cc_774 N_VPWR_c_1001_n N_Y_c_1217_n 0.0144623f $X=6.97 $Y=3.33 $X2=0 $Y2=0
cc_775 N_VPWR_c_973_n N_Y_c_1217_n 0.0118344f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_776 N_VPWR_c_985_n N_Y_c_1218_n 0.0357709f $X=9.805 $Y=2.085 $X2=0 $Y2=0
cc_777 N_VPWR_c_1005_n N_Y_c_1218_n 0.0144623f $X=10.67 $Y=3.33 $X2=0 $Y2=0
cc_778 N_VPWR_c_973_n N_Y_c_1218_n 0.0118344f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_779 N_VPWR_c_986_n N_Y_c_1219_n 0.00519412f $X=10.755 $Y=2.085 $X2=0 $Y2=0
cc_780 N_VPWR_c_1006_n N_Y_c_1219_n 0.014549f $X=11.62 $Y=3.33 $X2=0 $Y2=0
cc_781 N_VPWR_c_973_n N_Y_c_1219_n 0.0119743f $X=11.76 $Y=3.33 $X2=0 $Y2=0
cc_782 N_VPWR_M1006_s N_Y_c_1336_n 0.00519671f $X=5.12 $Y=1.84 $X2=0 $Y2=0
cc_783 N_VPWR_M1010_s N_Y_c_1336_n 0.00508955f $X=6.02 $Y=1.84 $X2=0 $Y2=0
cc_784 N_VPWR_M1014_s N_Y_c_1336_n 0.00500358f $X=6.92 $Y=1.84 $X2=0 $Y2=0
cc_785 N_VPWR_M1020_s N_Y_c_1336_n 0.00492968f $X=7.82 $Y=1.84 $X2=0 $Y2=0
cc_786 N_VPWR_M1030_s N_Y_c_1336_n 0.00501959f $X=8.72 $Y=1.84 $X2=0 $Y2=0
cc_787 N_VPWR_M1034_s N_Y_c_1336_n 0.00460673f $X=9.67 $Y=1.84 $X2=0 $Y2=0
cc_788 N_VPWR_M1040_s N_Y_c_1336_n 0.00388636f $X=10.62 $Y=1.84 $X2=0 $Y2=0
cc_789 N_VPWR_c_978_n N_Y_c_1336_n 0.00152375f $X=4.355 $Y=2.085 $X2=0 $Y2=0
cc_790 N_VPWR_c_979_n N_Y_c_1336_n 0.0188549f $X=5.255 $Y=2.085 $X2=0 $Y2=0
cc_791 N_VPWR_c_980_n N_Y_c_1336_n 0.0189031f $X=6.155 $Y=2.085 $X2=0 $Y2=0
cc_792 N_VPWR_c_981_n N_Y_c_1336_n 0.0189983f $X=7.055 $Y=2.085 $X2=0 $Y2=0
cc_793 N_VPWR_c_983_n N_Y_c_1336_n 0.0191011f $X=7.955 $Y=2.085 $X2=0 $Y2=0
cc_794 N_VPWR_c_984_n N_Y_c_1336_n 0.0234703f $X=8.855 $Y=2.085 $X2=0 $Y2=0
cc_795 N_VPWR_c_985_n N_Y_c_1336_n 0.0240975f $X=9.805 $Y=2.085 $X2=0 $Y2=0
cc_796 N_VPWR_c_986_n N_Y_c_1336_n 0.0228683f $X=10.755 $Y=2.085 $X2=0 $Y2=0
cc_797 N_VPWR_c_988_n N_Y_c_1336_n 0.00161542f $X=11.705 $Y=1.985 $X2=0 $Y2=0
cc_798 N_VPWR_c_981_n N_Y_c_1358_n 0.0376755f $X=7.055 $Y=2.085 $X2=0 $Y2=0
cc_799 N_VPWR_c_983_n N_Y_c_1358_n 0.0376755f $X=7.955 $Y=2.085 $X2=0 $Y2=0
cc_800 N_Y_c_1195_n N_VGND_c_1453_n 0.0296294f $X=4.78 $Y=0.515 $X2=0 $Y2=0
cc_801 N_Y_c_1195_n N_VGND_c_1454_n 0.026661f $X=4.78 $Y=0.515 $X2=0 $Y2=0
cc_802 N_Y_c_1196_n N_VGND_c_1454_n 0.00127089f $X=5.64 $Y=0.515 $X2=0 $Y2=0
cc_803 N_Y_c_1196_n N_VGND_c_1455_n 0.0277717f $X=5.64 $Y=0.515 $X2=0 $Y2=0
cc_804 N_Y_c_1197_n N_VGND_c_1455_n 0.0258753f $X=6.57 $Y=0.515 $X2=0 $Y2=0
cc_805 N_Y_c_1197_n N_VGND_c_1456_n 0.0277814f $X=6.57 $Y=0.515 $X2=0 $Y2=0
cc_806 N_Y_c_1198_n N_VGND_c_1456_n 0.0272176f $X=7.5 $Y=0.515 $X2=0 $Y2=0
cc_807 N_Y_c_1198_n N_VGND_c_1457_n 0.0277859f $X=7.5 $Y=0.515 $X2=0 $Y2=0
cc_808 N_Y_c_1199_n N_VGND_c_1457_n 0.0279399f $X=8.43 $Y=0.515 $X2=0 $Y2=0
cc_809 N_Y_c_1199_n N_VGND_c_1458_n 0.0277882f $X=8.43 $Y=0.515 $X2=0 $Y2=0
cc_810 N_Y_c_1200_n N_VGND_c_1458_n 0.0279399f $X=9.36 $Y=0.515 $X2=0 $Y2=0
cc_811 N_Y_c_1200_n N_VGND_c_1459_n 0.0277882f $X=9.36 $Y=0.515 $X2=0 $Y2=0
cc_812 N_Y_c_1201_n N_VGND_c_1459_n 0.0279399f $X=10.29 $Y=0.515 $X2=0 $Y2=0
cc_813 N_Y_c_1201_n N_VGND_c_1460_n 0.0277882f $X=10.29 $Y=0.515 $X2=0 $Y2=0
cc_814 N_Y_c_1202_n N_VGND_c_1460_n 0.0291199f $X=11.22 $Y=0.515 $X2=0 $Y2=0
cc_815 N_Y_c_1202_n N_VGND_c_1462_n 0.0308485f $X=11.22 $Y=0.515 $X2=0 $Y2=0
cc_816 N_Y_c_1195_n N_VGND_c_1469_n 0.0109942f $X=4.78 $Y=0.515 $X2=0 $Y2=0
cc_817 N_Y_c_1196_n N_VGND_c_1473_n 0.00950426f $X=5.64 $Y=0.515 $X2=0 $Y2=0
cc_818 N_Y_c_1197_n N_VGND_c_1474_n 0.0103698f $X=6.57 $Y=0.515 $X2=0 $Y2=0
cc_819 N_Y_c_1198_n N_VGND_c_1475_n 0.0107861f $X=7.5 $Y=0.515 $X2=0 $Y2=0
cc_820 N_Y_c_1199_n N_VGND_c_1476_n 0.0109942f $X=8.43 $Y=0.515 $X2=0 $Y2=0
cc_821 N_Y_c_1200_n N_VGND_c_1477_n 0.0109942f $X=9.36 $Y=0.515 $X2=0 $Y2=0
cc_822 N_Y_c_1201_n N_VGND_c_1478_n 0.0109942f $X=10.29 $Y=0.515 $X2=0 $Y2=0
cc_823 N_Y_c_1202_n N_VGND_c_1479_n 0.0144922f $X=11.22 $Y=0.515 $X2=0 $Y2=0
cc_824 N_Y_c_1195_n N_VGND_c_1488_n 0.00904371f $X=4.78 $Y=0.515 $X2=0 $Y2=0
cc_825 N_Y_c_1196_n N_VGND_c_1488_n 0.0078668f $X=5.64 $Y=0.515 $X2=0 $Y2=0
cc_826 N_Y_c_1197_n N_VGND_c_1488_n 0.00856206f $X=6.57 $Y=0.515 $X2=0 $Y2=0
cc_827 N_Y_c_1198_n N_VGND_c_1488_n 0.00888316f $X=7.5 $Y=0.515 $X2=0 $Y2=0
cc_828 N_Y_c_1199_n N_VGND_c_1488_n 0.00904371f $X=8.43 $Y=0.515 $X2=0 $Y2=0
cc_829 N_Y_c_1200_n N_VGND_c_1488_n 0.00904371f $X=9.36 $Y=0.515 $X2=0 $Y2=0
cc_830 N_Y_c_1201_n N_VGND_c_1488_n 0.00904371f $X=10.29 $Y=0.515 $X2=0 $Y2=0
cc_831 N_Y_c_1202_n N_VGND_c_1488_n 0.0118826f $X=11.22 $Y=0.515 $X2=0 $Y2=0

* NGSPICE file created from sky130_fd_sc_ms__xnor2_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__xnor2_1 A B VGND VNB VPB VPWR Y
M1000 VGND A a_293_74# VNB nlowvt w=740000u l=150000u
+  ad=5.4e+11p pd=4.52e+06u as=4.107e+11p ps=4.07e+06u
M1001 VPWR B a_141_385# VPB pshort w=840000u l=180000u
+  ad=1.13705e+12p pd=8.5e+06u as=2.268e+11p ps=2.22e+06u
M1002 a_141_385# B a_112_119# VNB nlowvt w=640000u l=150000u
+  ad=1.76e+11p pd=1.83e+06u as=1.344e+11p ps=1.7e+06u
M1003 a_379_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=0p ps=0u
M1004 Y a_141_385# a_293_74# VNB nlowvt w=740000u l=150000u
+  ad=2.294e+11p pd=2.1e+06u as=0p ps=0u
M1005 Y B a_379_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.368e+11p pd=3.02e+06u as=0p ps=0u
M1006 a_112_119# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_141_385# A VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_293_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_141_385# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__buf_4.pxi.spice
* Created: Wed Sep  2 11:59:35 2020
* 
x_PM_SKY130_FD_SC_MS__BUF_4%A_86_260# N_A_86_260#_M1007_d N_A_86_260#_M1001_d
+ N_A_86_260#_M1005_g N_A_86_260#_M1000_g N_A_86_260#_M1006_g
+ N_A_86_260#_M1003_g N_A_86_260#_M1008_g N_A_86_260#_M1004_g
+ N_A_86_260#_M1009_g N_A_86_260#_M1010_g N_A_86_260#_c_72_n N_A_86_260#_c_73_n
+ N_A_86_260#_c_74_n N_A_86_260#_c_75_n N_A_86_260#_c_153_p N_A_86_260#_c_85_n
+ N_A_86_260#_c_76_n N_A_86_260#_c_77_n N_A_86_260#_c_78_n N_A_86_260#_c_79_n
+ N_A_86_260#_c_80_n PM_SKY130_FD_SC_MS__BUF_4%A_86_260#
x_PM_SKY130_FD_SC_MS__BUF_4%A N_A_M1001_g N_A_M1002_g N_A_M1007_g A N_A_c_182_n
+ N_A_c_183_n PM_SKY130_FD_SC_MS__BUF_4%A
x_PM_SKY130_FD_SC_MS__BUF_4%VPWR N_VPWR_M1005_d N_VPWR_M1006_d N_VPWR_M1009_d
+ N_VPWR_M1002_s N_VPWR_c_221_n N_VPWR_c_222_n N_VPWR_c_223_n N_VPWR_c_224_n
+ N_VPWR_c_225_n N_VPWR_c_226_n VPWR N_VPWR_c_227_n N_VPWR_c_228_n
+ N_VPWR_c_229_n N_VPWR_c_230_n N_VPWR_c_231_n N_VPWR_c_220_n
+ PM_SKY130_FD_SC_MS__BUF_4%VPWR
x_PM_SKY130_FD_SC_MS__BUF_4%X N_X_M1000_s N_X_M1004_s N_X_M1005_s N_X_M1008_s
+ N_X_c_273_n N_X_c_274_n N_X_c_275_n N_X_c_279_n N_X_c_280_n N_X_c_276_n
+ N_X_c_281_n N_X_c_277_n N_X_c_282_n X PM_SKY130_FD_SC_MS__BUF_4%X
x_PM_SKY130_FD_SC_MS__BUF_4%VGND N_VGND_M1000_d N_VGND_M1003_d N_VGND_M1010_d
+ N_VGND_c_336_n N_VGND_c_337_n N_VGND_c_338_n N_VGND_c_339_n VGND
+ N_VGND_c_340_n N_VGND_c_341_n N_VGND_c_342_n N_VGND_c_343_n N_VGND_c_344_n
+ PM_SKY130_FD_SC_MS__BUF_4%VGND
cc_1 VNB N_A_86_260#_M1005_g 0.0175041f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.4
cc_2 VNB N_A_86_260#_M1000_g 0.0265448f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_3 VNB N_A_86_260#_M1006_g 0.0015344f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.4
cc_4 VNB N_A_86_260#_M1003_g 0.022504f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_5 VNB N_A_86_260#_M1008_g 0.00154196f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=2.4
cc_6 VNB N_A_86_260#_M1004_g 0.0225168f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=0.74
cc_7 VNB N_A_86_260#_M1009_g 0.00168554f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=2.4
cc_8 VNB N_A_86_260#_M1010_g 0.0249635f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=0.74
cc_9 VNB N_A_86_260#_c_72_n 0.0145731f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.375
cc_10 VNB N_A_86_260#_c_73_n 0.00768954f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=1.465
cc_11 VNB N_A_86_260#_c_74_n 0.00389847f $X=-0.19 $Y=-0.245 $X2=2.2 $Y2=1.3
cc_12 VNB N_A_86_260#_c_75_n 0.00548705f $X=-0.19 $Y=-0.245 $X2=2.915 $Y2=1.045
cc_13 VNB N_A_86_260#_c_76_n 0.02581f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=0.515
cc_14 VNB N_A_86_260#_c_77_n 0.0249538f $X=-0.19 $Y=-0.245 $X2=3.16 $Y2=1.95
cc_15 VNB N_A_86_260#_c_78_n 0.0124806f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=1.045
cc_16 VNB N_A_86_260#_c_79_n 0.00922324f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=1.465
cc_17 VNB N_A_86_260#_c_80_n 0.0668824f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=1.465
cc_18 VNB N_A_M1007_g 0.0330952f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.3
cc_19 VNB N_A_c_182_n 0.00412911f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.4
cc_20 VNB N_A_c_183_n 0.0436966f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.4
cc_21 VNB N_VPWR_c_220_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_X_c_273_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=1.375
cc_23 VNB N_X_c_274_n 0.00290742f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.63
cc_24 VNB N_X_c_275_n 0.00335622f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.4
cc_25 VNB N_X_c_276_n 0.00542414f $X=-0.19 $Y=-0.245 $X2=1.42 $Y2=2.4
cc_26 VNB N_X_c_277_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=1.3
cc_27 VNB N_VGND_c_336_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_337_n 0.0376574f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_29 VNB N_VGND_c_338_n 0.00830803f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.375
cc_30 VNB N_VGND_c_339_n 0.0187266f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.4
cc_31 VNB N_VGND_c_340_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_32 VNB N_VGND_c_341_n 0.0191816f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.3
cc_33 VNB N_VGND_c_342_n 0.204744f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=0.74
cc_34 VNB N_VGND_c_343_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_344_n 0.0243944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_A_86_260#_M1005_g 0.0289586f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=2.4
cc_37 VPB N_A_86_260#_M1006_g 0.021401f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=2.4
cc_38 VPB N_A_86_260#_M1008_g 0.0214376f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=2.4
cc_39 VPB N_A_86_260#_M1009_g 0.0246042f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=2.4
cc_40 VPB N_A_86_260#_c_85_n 0.0105449f $X=-0.19 $Y=1.66 $X2=3.075 $Y2=2.075
cc_41 VPB N_A_86_260#_c_77_n 0.0122364f $X=-0.19 $Y=1.66 $X2=3.16 $Y2=1.95
cc_42 VPB N_A_M1001_g 0.0223819f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A_M1002_g 0.0228274f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.45
cc_44 VPB N_A_c_182_n 0.00322424f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=2.4
cc_45 VPB N_A_c_183_n 0.00487278f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=2.4
cc_46 VPB N_VPWR_c_221_n 0.0124752f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_47 VPB N_VPWR_c_222_n 0.064803f $X=-0.19 $Y=1.66 $X2=0.88 $Y2=1.375
cc_48 VPB N_VPWR_c_223_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.3
cc_49 VPB N_VPWR_c_224_n 0.0122571f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=1.63
cc_50 VPB N_VPWR_c_225_n 0.0121909f $X=-0.19 $Y=1.66 $X2=1.565 $Y2=1.3
cc_51 VPB N_VPWR_c_226_n 0.0391172f $X=-0.19 $Y=1.66 $X2=1.565 $Y2=0.74
cc_52 VPB N_VPWR_c_227_n 0.0164074f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=2.4
cc_53 VPB N_VPWR_c_228_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_229_n 0.0207798f $X=-0.19 $Y=1.66 $X2=1.225 $Y2=1.465
cc_55 VPB N_VPWR_c_230_n 0.00601644f $X=-0.19 $Y=1.66 $X2=3.075 $Y2=2.075
cc_56 VPB N_VPWR_c_231_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_220_n 0.0752858f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_X_c_275_n 0.00272979f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=2.4
cc_59 VPB N_X_c_279_n 0.00184146f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.3
cc_60 VPB N_X_c_280_n 0.00499535f $X=-0.19 $Y=1.66 $X2=1.42 $Y2=1.63
cc_61 VPB N_X_c_281_n 0.00179594f $X=-0.19 $Y=1.66 $X2=1.565 $Y2=0.74
cc_62 VPB N_X_c_282_n 3.92079e-19 $X=-0.19 $Y=1.66 $X2=1.995 $Y2=0.74
cc_63 N_A_86_260#_c_85_n N_A_M1001_g 0.005558f $X=3.075 $Y=2.075 $X2=0 $Y2=0
cc_64 N_A_86_260#_c_85_n N_A_M1002_g 0.0200318f $X=3.075 $Y=2.075 $X2=0 $Y2=0
cc_65 N_A_86_260#_M1010_g N_A_M1007_g 0.0127822f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_66 N_A_86_260#_c_73_n N_A_M1007_g 0.00105416f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_67 N_A_86_260#_c_74_n N_A_M1007_g 0.00275276f $X=2.2 $Y=1.3 $X2=0 $Y2=0
cc_68 N_A_86_260#_c_75_n N_A_M1007_g 0.0131472f $X=2.915 $Y=1.045 $X2=0 $Y2=0
cc_69 N_A_86_260#_c_76_n N_A_M1007_g 0.0174462f $X=3.08 $Y=0.515 $X2=0 $Y2=0
cc_70 N_A_86_260#_c_77_n N_A_M1007_g 0.00778767f $X=3.16 $Y=1.95 $X2=0 $Y2=0
cc_71 N_A_86_260#_c_78_n N_A_M1007_g 0.00206782f $X=3.08 $Y=1.045 $X2=0 $Y2=0
cc_72 N_A_86_260#_M1009_g N_A_c_182_n 2.06048e-19 $X=1.87 $Y=2.4 $X2=0 $Y2=0
cc_73 N_A_86_260#_c_73_n N_A_c_182_n 0.0192045f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_74 N_A_86_260#_c_75_n N_A_c_182_n 0.0237625f $X=2.915 $Y=1.045 $X2=0 $Y2=0
cc_75 N_A_86_260#_c_85_n N_A_c_182_n 0.026883f $X=3.075 $Y=2.075 $X2=0 $Y2=0
cc_76 N_A_86_260#_c_77_n N_A_c_182_n 0.0326294f $X=3.16 $Y=1.95 $X2=0 $Y2=0
cc_77 N_A_86_260#_c_80_n N_A_c_182_n 5.66834e-19 $X=1.995 $Y=1.465 $X2=0 $Y2=0
cc_78 N_A_86_260#_M1009_g N_A_c_183_n 0.0210853f $X=1.87 $Y=2.4 $X2=0 $Y2=0
cc_79 N_A_86_260#_c_73_n N_A_c_183_n 0.00188928f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_80 N_A_86_260#_c_75_n N_A_c_183_n 0.00850991f $X=2.915 $Y=1.045 $X2=0 $Y2=0
cc_81 N_A_86_260#_c_85_n N_A_c_183_n 5.04899e-19 $X=3.075 $Y=2.075 $X2=0 $Y2=0
cc_82 N_A_86_260#_c_77_n N_A_c_183_n 0.0166059f $X=3.16 $Y=1.95 $X2=0 $Y2=0
cc_83 N_A_86_260#_c_78_n N_A_c_183_n 2.29254e-19 $X=3.08 $Y=1.045 $X2=0 $Y2=0
cc_84 N_A_86_260#_c_80_n N_A_c_183_n 0.00876655f $X=1.995 $Y=1.465 $X2=0 $Y2=0
cc_85 N_A_86_260#_c_85_n N_VPWR_M1002_s 0.00668552f $X=3.075 $Y=2.075 $X2=0
+ $Y2=0
cc_86 N_A_86_260#_c_77_n N_VPWR_M1002_s 0.00183735f $X=3.16 $Y=1.95 $X2=0 $Y2=0
cc_87 N_A_86_260#_M1005_g N_VPWR_c_222_n 0.0218617f $X=0.52 $Y=2.4 $X2=0 $Y2=0
cc_88 N_A_86_260#_M1006_g N_VPWR_c_222_n 6.98003e-19 $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_89 N_A_86_260#_M1005_g N_VPWR_c_223_n 5.82463e-19 $X=0.52 $Y=2.4 $X2=0 $Y2=0
cc_90 N_A_86_260#_M1006_g N_VPWR_c_223_n 0.0168011f $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_91 N_A_86_260#_M1008_g N_VPWR_c_223_n 0.0168979f $X=1.42 $Y=2.4 $X2=0 $Y2=0
cc_92 N_A_86_260#_M1009_g N_VPWR_c_223_n 5.88636e-19 $X=1.87 $Y=2.4 $X2=0 $Y2=0
cc_93 N_A_86_260#_M1008_g N_VPWR_c_224_n 6.98003e-19 $X=1.42 $Y=2.4 $X2=0 $Y2=0
cc_94 N_A_86_260#_M1009_g N_VPWR_c_224_n 0.0203293f $X=1.87 $Y=2.4 $X2=0 $Y2=0
cc_95 N_A_86_260#_c_73_n N_VPWR_c_224_n 0.0267415f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_96 N_A_86_260#_c_80_n N_VPWR_c_224_n 0.00296151f $X=1.995 $Y=1.465 $X2=0
+ $Y2=0
cc_97 N_A_86_260#_c_85_n N_VPWR_c_226_n 0.0235456f $X=3.075 $Y=2.075 $X2=0 $Y2=0
cc_98 N_A_86_260#_M1005_g N_VPWR_c_227_n 0.00460063f $X=0.52 $Y=2.4 $X2=0 $Y2=0
cc_99 N_A_86_260#_M1006_g N_VPWR_c_227_n 0.00460063f $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_100 N_A_86_260#_M1008_g N_VPWR_c_228_n 0.00460063f $X=1.42 $Y=2.4 $X2=0 $Y2=0
cc_101 N_A_86_260#_M1009_g N_VPWR_c_228_n 0.00460063f $X=1.87 $Y=2.4 $X2=0 $Y2=0
cc_102 N_A_86_260#_M1005_g N_VPWR_c_220_n 0.00908554f $X=0.52 $Y=2.4 $X2=0 $Y2=0
cc_103 N_A_86_260#_M1006_g N_VPWR_c_220_n 0.00908554f $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_104 N_A_86_260#_M1008_g N_VPWR_c_220_n 0.00908554f $X=1.42 $Y=2.4 $X2=0 $Y2=0
cc_105 N_A_86_260#_M1009_g N_VPWR_c_220_n 0.00908554f $X=1.87 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A_86_260#_M1000_g N_X_c_273_n 0.00767507f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_107 N_A_86_260#_M1003_g N_X_c_273_n 0.00916694f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_108 N_A_86_260#_M1004_g N_X_c_273_n 6.18925e-19 $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_109 N_A_86_260#_M1000_g N_X_c_274_n 0.0154604f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_110 N_A_86_260#_M1003_g N_X_c_274_n 0.00546031f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_111 N_A_86_260#_c_72_n N_X_c_274_n 0.00653153f $X=0.535 $Y=1.375 $X2=0 $Y2=0
cc_112 N_A_86_260#_c_73_n N_X_c_274_n 0.00679785f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_113 N_A_86_260#_c_79_n N_X_c_274_n 0.00719234f $X=0.88 $Y=1.465 $X2=0 $Y2=0
cc_114 N_A_86_260#_M1005_g N_X_c_275_n 0.00844264f $X=0.52 $Y=2.4 $X2=0 $Y2=0
cc_115 N_A_86_260#_c_73_n N_X_c_275_n 0.014004f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_116 N_A_86_260#_c_79_n N_X_c_275_n 0.00499189f $X=0.88 $Y=1.465 $X2=0 $Y2=0
cc_117 N_A_86_260#_c_80_n N_X_c_275_n 0.00586219f $X=1.995 $Y=1.465 $X2=0 $Y2=0
cc_118 N_A_86_260#_M1005_g N_X_c_279_n 3.62784e-19 $X=0.52 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A_86_260#_M1006_g N_X_c_279_n 3.65169e-19 $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A_86_260#_M1006_g N_X_c_280_n 0.0172188f $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_121 N_A_86_260#_M1008_g N_X_c_280_n 0.0145668f $X=1.42 $Y=2.4 $X2=0 $Y2=0
cc_122 N_A_86_260#_M1009_g N_X_c_280_n 8.09632e-19 $X=1.87 $Y=2.4 $X2=0 $Y2=0
cc_123 N_A_86_260#_c_73_n N_X_c_280_n 0.0512087f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_124 N_A_86_260#_c_80_n N_X_c_280_n 0.00450883f $X=1.995 $Y=1.465 $X2=0 $Y2=0
cc_125 N_A_86_260#_M1003_g N_X_c_276_n 0.0135497f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A_86_260#_M1004_g N_X_c_276_n 0.0128445f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A_86_260#_M1010_g N_X_c_276_n 0.00240508f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A_86_260#_c_73_n N_X_c_276_n 0.0687837f $X=2.115 $Y=1.465 $X2=0 $Y2=0
cc_129 N_A_86_260#_c_153_p N_X_c_276_n 0.00808483f $X=2.285 $Y=1.045 $X2=0 $Y2=0
cc_130 N_A_86_260#_c_80_n N_X_c_276_n 0.0087353f $X=1.995 $Y=1.465 $X2=0 $Y2=0
cc_131 N_A_86_260#_M1008_g N_X_c_281_n 3.62369e-19 $X=1.42 $Y=2.4 $X2=0 $Y2=0
cc_132 N_A_86_260#_M1009_g N_X_c_281_n 3.62369e-19 $X=1.87 $Y=2.4 $X2=0 $Y2=0
cc_133 N_A_86_260#_M1003_g N_X_c_277_n 6.18925e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A_86_260#_M1004_g N_X_c_277_n 0.00916694f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A_86_260#_M1010_g N_X_c_277_n 0.0167949f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A_86_260#_M1005_g N_X_c_282_n 8.09632e-19 $X=0.52 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A_86_260#_c_75_n N_VGND_M1010_d 0.00863822f $X=2.915 $Y=1.045 $X2=0
+ $Y2=0
cc_138 N_A_86_260#_c_153_p N_VGND_M1010_d 0.00351113f $X=2.285 $Y=1.045 $X2=0
+ $Y2=0
cc_139 N_A_86_260#_M1000_g N_VGND_c_337_n 0.0161039f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_140 N_A_86_260#_c_72_n N_VGND_c_337_n 3.61737e-19 $X=0.535 $Y=1.375 $X2=0
+ $Y2=0
cc_141 N_A_86_260#_M1003_g N_VGND_c_338_n 0.00454042f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_142 N_A_86_260#_M1004_g N_VGND_c_338_n 0.00454042f $X=1.565 $Y=0.74 $X2=0
+ $Y2=0
cc_143 N_A_86_260#_M1004_g N_VGND_c_339_n 0.00434272f $X=1.565 $Y=0.74 $X2=0
+ $Y2=0
cc_144 N_A_86_260#_M1010_g N_VGND_c_339_n 0.00434272f $X=1.995 $Y=0.74 $X2=0
+ $Y2=0
cc_145 N_A_86_260#_M1000_g N_VGND_c_340_n 0.00434272f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_146 N_A_86_260#_M1003_g N_VGND_c_340_n 0.00434272f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_147 N_A_86_260#_c_76_n N_VGND_c_341_n 0.0145639f $X=3.08 $Y=0.515 $X2=0 $Y2=0
cc_148 N_A_86_260#_M1000_g N_VGND_c_342_n 0.00823934f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_149 N_A_86_260#_M1003_g N_VGND_c_342_n 0.00821294f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_150 N_A_86_260#_M1004_g N_VGND_c_342_n 0.00821294f $X=1.565 $Y=0.74 $X2=0
+ $Y2=0
cc_151 N_A_86_260#_M1010_g N_VGND_c_342_n 0.00822986f $X=1.995 $Y=0.74 $X2=0
+ $Y2=0
cc_152 N_A_86_260#_c_76_n N_VGND_c_342_n 0.0119984f $X=3.08 $Y=0.515 $X2=0 $Y2=0
cc_153 N_A_86_260#_M1010_g N_VGND_c_344_n 0.00543794f $X=1.995 $Y=0.74 $X2=0
+ $Y2=0
cc_154 N_A_86_260#_c_75_n N_VGND_c_344_n 0.0251789f $X=2.915 $Y=1.045 $X2=0
+ $Y2=0
cc_155 N_A_86_260#_c_153_p N_VGND_c_344_n 0.00982229f $X=2.285 $Y=1.045 $X2=0
+ $Y2=0
cc_156 N_A_86_260#_c_76_n N_VGND_c_344_n 0.013254f $X=3.08 $Y=0.515 $X2=0 $Y2=0
cc_157 N_A_M1001_g N_VPWR_c_224_n 0.00707382f $X=2.405 $Y=2.26 $X2=0 $Y2=0
cc_158 N_A_M1001_g N_VPWR_c_226_n 0.00132812f $X=2.405 $Y=2.26 $X2=0 $Y2=0
cc_159 N_A_M1002_g N_VPWR_c_226_n 0.0126632f $X=2.855 $Y=2.26 $X2=0 $Y2=0
cc_160 N_A_M1001_g N_VPWR_c_229_n 0.00482866f $X=2.405 $Y=2.26 $X2=0 $Y2=0
cc_161 N_A_M1002_g N_VPWR_c_229_n 0.00401533f $X=2.855 $Y=2.26 $X2=0 $Y2=0
cc_162 N_A_M1001_g N_VPWR_c_220_n 0.00555093f $X=2.405 $Y=2.26 $X2=0 $Y2=0
cc_163 N_A_M1002_g N_VPWR_c_220_n 0.00465661f $X=2.855 $Y=2.26 $X2=0 $Y2=0
cc_164 N_A_M1007_g N_VGND_c_341_n 0.00434272f $X=2.865 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A_M1007_g N_VGND_c_342_n 0.00826644f $X=2.865 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A_M1007_g N_VGND_c_344_n 0.00703669f $X=2.865 $Y=0.74 $X2=0 $Y2=0
cc_167 N_VPWR_c_222_n N_X_c_279_n 0.0339152f $X=0.295 $Y=1.985 $X2=0 $Y2=0
cc_168 N_VPWR_c_223_n N_X_c_279_n 0.0288913f $X=1.195 $Y=2.225 $X2=0 $Y2=0
cc_169 N_VPWR_c_227_n N_X_c_279_n 0.00771942f $X=1.03 $Y=3.33 $X2=0 $Y2=0
cc_170 N_VPWR_c_220_n N_X_c_279_n 0.00638947f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_171 N_VPWR_M1006_d N_X_c_280_n 0.00165831f $X=1.06 $Y=1.84 $X2=0 $Y2=0
cc_172 N_VPWR_c_223_n N_X_c_280_n 0.0170259f $X=1.195 $Y=2.225 $X2=0 $Y2=0
cc_173 N_VPWR_c_224_n N_X_c_280_n 0.00575112f $X=2.095 $Y=1.985 $X2=0 $Y2=0
cc_174 N_VPWR_c_223_n N_X_c_281_n 0.0283117f $X=1.195 $Y=2.225 $X2=0 $Y2=0
cc_175 N_VPWR_c_224_n N_X_c_281_n 0.0339124f $X=2.095 $Y=1.985 $X2=0 $Y2=0
cc_176 N_VPWR_c_228_n N_X_c_281_n 0.00749631f $X=1.93 $Y=3.33 $X2=0 $Y2=0
cc_177 N_VPWR_c_220_n N_X_c_281_n 0.0062048f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_178 N_VPWR_c_222_n N_X_c_282_n 0.00575112f $X=0.295 $Y=1.985 $X2=0 $Y2=0
cc_179 N_X_c_276_n N_VGND_M1003_d 0.00374767f $X=1.615 $Y=1.045 $X2=0 $Y2=0
cc_180 N_X_c_273_n N_VGND_c_337_n 0.0236416f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_181 N_X_c_273_n N_VGND_c_338_n 0.0173003f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_182 N_X_c_276_n N_VGND_c_338_n 0.0248957f $X=1.615 $Y=1.045 $X2=0 $Y2=0
cc_183 N_X_c_277_n N_VGND_c_338_n 0.0173003f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_184 N_X_c_277_n N_VGND_c_339_n 0.0144922f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_185 N_X_c_273_n N_VGND_c_340_n 0.0144922f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_186 N_X_c_273_n N_VGND_c_342_n 0.0118826f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_187 N_X_c_277_n N_VGND_c_342_n 0.0118826f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_188 N_X_c_277_n N_VGND_c_344_n 0.013254f $X=1.78 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__nor3b_1.spice
* Created: Wed Sep  2 12:16:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nor3b_1.pex.spice"
.subckt sky130_fd_sc_ms__nor3b_1  VNB VPB C_N A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_C_N_M1004_g N_A_27_112#_M1004_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.116971 AS=0.2695 PD=0.963566 PS=2.08 NRD=18 NRS=0 M=1 R=3.66667
+ SA=75000.4 SB=75001.8 A=0.0825 P=1.4 MULT=1
MM1007 N_Y_M1007_d N_A_M1007_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.74 AD=0.1184
+ AS=0.157379 PD=1.06 PS=1.29643 NRD=6.48 NRS=4.86 M=1 R=4.93333 SA=75000.8
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_B_M1005_g N_Y_M1007_d VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.1184 PD=1.16 PS=1.06 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.2 SB=75000.8
+ A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A_27_112#_M1000_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.8
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_VPWR_M1006_d N_C_N_M1006_g N_A_27_112#_M1006_s VPB PSHORT L=0.18 W=0.84
+ AD=0.174 AS=0.2352 PD=1.29429 PS=2.24 NRD=26.9693 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90001.7 A=0.1512 P=2.04 MULT=1
MM1003 A_263_368# N_A_M1003_g N_VPWR_M1006_d VPB PSHORT L=0.18 W=1.12 AD=0.1344
+ AS=0.232 PD=1.36 PS=1.72571 NRD=11.426 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1002 A_347_368# N_B_M1002_g A_263_368# VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.1344 PD=1.51 PS=1.36 NRD=24.6053 NRS=11.426 M=1 R=6.22222 SA=90001
+ SB=90000.8 A=0.2016 P=2.6 MULT=1
MM1001 N_Y_M1001_d N_A_27_112#_M1001_g A_347_368# VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.2184 PD=2.8 PS=1.51 NRD=0 NRS=24.6053 M=1 R=6.22222 SA=90001.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ms__nor3b_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__nand3_2.pxi.spice
* Created: Wed Sep  2 12:13:36 2020
* 
x_PM_SKY130_FD_SC_MS__NAND3_2%C N_C_c_61_n N_C_M1000_g N_C_M1004_g N_C_c_63_n
+ N_C_M1010_g N_C_M1005_g C N_C_c_65_n N_C_c_66_n PM_SKY130_FD_SC_MS__NAND3_2%C
x_PM_SKY130_FD_SC_MS__NAND3_2%B N_B_M1007_g N_B_M1003_g N_B_M1008_g N_B_M1009_g
+ N_B_c_134_p N_B_c_164_p N_B_c_115_n N_B_c_116_n N_B_c_117_n B N_B_c_118_n
+ N_B_c_119_n B PM_SKY130_FD_SC_MS__NAND3_2%B
x_PM_SKY130_FD_SC_MS__NAND3_2%A N_A_M1002_g N_A_M1001_g N_A_M1011_g N_A_M1006_g
+ A N_A_c_209_n N_A_c_206_n PM_SKY130_FD_SC_MS__NAND3_2%A
x_PM_SKY130_FD_SC_MS__NAND3_2%VPWR N_VPWR_M1004_s N_VPWR_M1005_s N_VPWR_M1001_d
+ N_VPWR_M1008_s N_VPWR_c_259_n N_VPWR_c_260_n N_VPWR_c_261_n N_VPWR_c_262_n
+ N_VPWR_c_263_n N_VPWR_c_264_n VPWR N_VPWR_c_265_n N_VPWR_c_266_n
+ N_VPWR_c_267_n N_VPWR_c_268_n N_VPWR_c_269_n N_VPWR_c_258_n
+ PM_SKY130_FD_SC_MS__NAND3_2%VPWR
x_PM_SKY130_FD_SC_MS__NAND3_2%Y N_Y_M1002_s N_Y_M1004_d N_Y_M1003_d N_Y_M1006_s
+ N_Y_c_315_n N_Y_c_312_n N_Y_c_322_n N_Y_c_342_n N_Y_c_346_n N_Y_c_347_n
+ N_Y_c_316_n N_Y_c_317_n N_Y_c_313_n N_Y_c_314_n Y Y
+ PM_SKY130_FD_SC_MS__NAND3_2%Y
x_PM_SKY130_FD_SC_MS__NAND3_2%A_27_74# N_A_27_74#_M1000_d N_A_27_74#_M1010_d
+ N_A_27_74#_M1009_s N_A_27_74#_c_396_n N_A_27_74#_c_401_n N_A_27_74#_c_409_n
+ N_A_27_74#_c_397_n N_A_27_74#_c_398_n N_A_27_74#_c_399_n
+ PM_SKY130_FD_SC_MS__NAND3_2%A_27_74#
x_PM_SKY130_FD_SC_MS__NAND3_2%VGND N_VGND_M1000_s N_VGND_c_455_n VGND
+ N_VGND_c_456_n N_VGND_c_457_n N_VGND_c_458_n N_VGND_c_459_n
+ PM_SKY130_FD_SC_MS__NAND3_2%VGND
x_PM_SKY130_FD_SC_MS__NAND3_2%A_283_74# N_A_283_74#_M1007_d N_A_283_74#_M1011_d
+ N_A_283_74#_c_495_n PM_SKY130_FD_SC_MS__NAND3_2%A_283_74#
cc_1 VNB N_C_c_61_n 0.0221619f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.22
cc_2 VNB N_C_M1004_g 0.00915832f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_3 VNB N_C_c_63_n 0.0162301f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.22
cc_4 VNB N_C_M1005_g 8.89891e-19 $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_5 VNB N_C_c_65_n 0.0251517f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.385
cc_6 VNB N_C_c_66_n 0.0464143f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.43
cc_7 VNB N_B_M1007_g 0.0248915f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.74
cc_8 VNB N_B_M1008_g 7.20106e-19 $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.64
cc_9 VNB N_B_M1009_g 0.0280879f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB N_B_c_115_n 3.02997e-19 $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.385
cc_11 VNB N_B_c_116_n 0.01693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B_c_117_n 0.0350063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B_c_118_n 0.0232586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B_c_119_n 0.0054119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_M1002_g 0.0198416f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.74
cc_16 VNB N_A_M1011_g 0.0203106f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.64
cc_17 VNB N_A_c_206_n 0.0389992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_258_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_312_n 0.010102f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.43
cc_20 VNB N_Y_c_313_n 0.00300143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_314_n 0.00225359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_396_n 0.0172715f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_23 VNB N_A_27_74#_c_397_n 0.0110846f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.385
cc_24 VNB N_A_27_74#_c_398_n 0.00213939f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.365
cc_25 VNB N_A_27_74#_c_399_n 0.0331002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_455_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_27 VNB N_VGND_c_456_n 0.0162587f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.74
cc_28 VNB N_VGND_c_457_n 0.0629719f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.385
cc_29 VNB N_VGND_c_458_n 0.205212f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.385
cc_30 VNB N_VGND_c_459_n 0.00601569f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_31 VNB N_A_283_74#_c_495_n 0.0141546f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.64
cc_32 VPB N_C_M1004_g 0.028074f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_33 VPB N_C_M1005_g 0.0222768f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_34 VPB N_B_M1003_g 0.0219022f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_B_M1008_g 0.0276238f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.64
cc_36 VPB N_B_c_115_n 0.00150135f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.385
cc_37 VPB B 0.00120134f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_B_c_118_n 0.00541504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_B_c_119_n 0.00185734f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A_M1001_g 0.0219052f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_A_M1006_g 0.0216796f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_42 VPB N_A_c_209_n 0.00348454f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.365
cc_43 VPB N_A_c_206_n 0.00602543f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_259_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_45 VPB N_VPWR_c_260_n 0.0574987f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_46 VPB N_VPWR_c_261_n 0.00884785f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.385
cc_47 VPB N_VPWR_c_262_n 0.00578359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_263_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.365
cc_49 VPB N_VPWR_c_264_n 0.0571953f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_265_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_266_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_267_n 0.0183691f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_268_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_269_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_258_n 0.0596689f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_Y_c_315_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_57 VPB N_Y_c_316_n 0.00220582f $X=-0.19 $Y=1.66 $X2=0.57 $Y2=1.365
cc_58 VPB N_Y_c_317_n 0.00569592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_Y_c_313_n 0.0012232f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB Y 0.00235965f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 N_C_c_63_n N_B_M1007_g 0.0140681f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_62 N_C_c_66_n N_B_M1007_g 0.0166541f $X=0.91 $Y=1.43 $X2=0 $Y2=0
cc_63 N_C_M1005_g N_B_M1003_g 0.0367895f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_64 N_C_M1005_g B 2.98095e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_65 N_C_c_66_n N_B_c_118_n 0.00790688f $X=0.91 $Y=1.43 $X2=0 $Y2=0
cc_66 N_C_c_66_n N_B_c_119_n 2.77958e-19 $X=0.91 $Y=1.43 $X2=0 $Y2=0
cc_67 N_C_M1004_g N_VPWR_c_260_n 0.00649215f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_68 N_C_c_65_n N_VPWR_c_260_n 0.0154298f $X=0.57 $Y=1.385 $X2=0 $Y2=0
cc_69 N_C_M1005_g N_VPWR_c_261_n 0.00318542f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_70 N_C_M1004_g N_VPWR_c_265_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_71 N_C_M1005_g N_VPWR_c_265_n 0.005209f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_72 N_C_M1004_g N_VPWR_c_258_n 0.00986008f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_73 N_C_M1005_g N_VPWR_c_258_n 0.0098216f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_74 N_C_M1004_g N_Y_c_315_n 0.00729841f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_75 N_C_M1005_g N_Y_c_315_n 0.00815638f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_76 N_C_c_61_n N_Y_c_322_n 5.01846e-19 $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_77 N_C_c_63_n N_Y_c_322_n 0.0049118f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_78 N_C_c_65_n N_Y_c_322_n 0.0061979f $X=0.57 $Y=1.385 $X2=0 $Y2=0
cc_79 N_C_c_66_n N_Y_c_322_n 0.00189162f $X=0.91 $Y=1.43 $X2=0 $Y2=0
cc_80 N_C_M1004_g N_Y_c_317_n 0.00905778f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_81 N_C_M1005_g N_Y_c_317_n 0.0252789f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_82 N_C_c_65_n N_Y_c_317_n 0.0100415f $X=0.57 $Y=1.385 $X2=0 $Y2=0
cc_83 N_C_c_66_n N_Y_c_317_n 0.00280483f $X=0.91 $Y=1.43 $X2=0 $Y2=0
cc_84 N_C_M1004_g N_Y_c_313_n 0.00153449f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_85 N_C_M1005_g N_Y_c_313_n 0.0052949f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_86 N_C_c_65_n N_Y_c_313_n 0.0199139f $X=0.57 $Y=1.385 $X2=0 $Y2=0
cc_87 N_C_c_66_n N_Y_c_313_n 0.0111382f $X=0.91 $Y=1.43 $X2=0 $Y2=0
cc_88 N_C_M1005_g Y 5.43358e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_89 N_C_c_61_n N_A_27_74#_c_396_n 4.43891e-19 $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_90 N_C_c_61_n N_A_27_74#_c_401_n 0.00948928f $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_91 N_C_c_63_n N_A_27_74#_c_401_n 0.0125772f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_92 N_C_c_65_n N_A_27_74#_c_401_n 0.0153562f $X=0.57 $Y=1.385 $X2=0 $Y2=0
cc_93 N_C_c_66_n N_A_27_74#_c_401_n 8.56627e-19 $X=0.91 $Y=1.43 $X2=0 $Y2=0
cc_94 N_C_c_61_n N_A_27_74#_c_397_n 0.00343023f $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_95 N_C_c_63_n N_A_27_74#_c_397_n 5.20319e-19 $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_96 N_C_c_65_n N_A_27_74#_c_397_n 0.0236506f $X=0.57 $Y=1.385 $X2=0 $Y2=0
cc_97 N_C_c_63_n N_A_27_74#_c_398_n 2.82836e-19 $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_98 N_C_c_61_n N_VGND_c_455_n 0.0095457f $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_99 N_C_c_63_n N_VGND_c_455_n 0.00663018f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_100 N_C_c_61_n N_VGND_c_456_n 0.00281948f $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_101 N_C_c_63_n N_VGND_c_457_n 0.00281141f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_102 N_C_c_61_n N_VGND_c_458_n 0.00367131f $X=0.48 $Y=1.22 $X2=0 $Y2=0
cc_103 N_C_c_63_n N_VGND_c_458_n 0.00365164f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_104 N_B_M1007_g N_A_M1002_g 0.0311226f $X=1.34 $Y=0.74 $X2=0 $Y2=0
cc_105 N_B_M1003_g N_A_M1001_g 0.0305505f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_106 N_B_c_134_p N_A_M1001_g 0.0163801f $X=2.655 $Y=2.035 $X2=0 $Y2=0
cc_107 B N_A_M1001_g 0.00302106f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_108 N_B_M1009_g N_A_M1011_g 0.0295756f $X=2.88 $Y=0.795 $X2=0 $Y2=0
cc_109 N_B_c_116_n N_A_M1011_g 6.56671e-19 $X=2.9 $Y=1.485 $X2=0 $Y2=0
cc_110 N_B_c_117_n N_A_M1011_g 9.74524e-19 $X=2.9 $Y=1.485 $X2=0 $Y2=0
cc_111 N_B_c_134_p N_A_M1006_g 0.0172229f $X=2.655 $Y=2.035 $X2=0 $Y2=0
cc_112 N_B_c_134_p N_A_c_209_n 0.0221964f $X=2.655 $Y=2.035 $X2=0 $Y2=0
cc_113 N_B_c_115_n N_A_c_209_n 0.00598812f $X=2.74 $Y=1.95 $X2=0 $Y2=0
cc_114 N_B_c_116_n N_A_c_209_n 0.0101158f $X=2.9 $Y=1.485 $X2=0 $Y2=0
cc_115 B N_A_c_209_n 0.00790543f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_116 N_B_c_118_n N_A_c_209_n 2.16173e-19 $X=1.43 $Y=1.515 $X2=0 $Y2=0
cc_117 N_B_c_119_n N_A_c_209_n 0.015572f $X=1.61 $Y=1.68 $X2=0 $Y2=0
cc_118 N_B_M1008_g N_A_c_206_n 0.0319432f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_119 N_B_c_134_p N_A_c_206_n 7.30233e-19 $X=2.655 $Y=2.035 $X2=0 $Y2=0
cc_120 N_B_c_115_n N_A_c_206_n 0.00459551f $X=2.74 $Y=1.95 $X2=0 $Y2=0
cc_121 N_B_c_116_n N_A_c_206_n 0.00414741f $X=2.9 $Y=1.485 $X2=0 $Y2=0
cc_122 N_B_c_117_n N_A_c_206_n 0.0166521f $X=2.9 $Y=1.485 $X2=0 $Y2=0
cc_123 N_B_c_118_n N_A_c_206_n 0.0209478f $X=1.43 $Y=1.515 $X2=0 $Y2=0
cc_124 N_B_c_119_n N_A_c_206_n 0.00171302f $X=1.61 $Y=1.68 $X2=0 $Y2=0
cc_125 N_B_c_134_p N_VPWR_M1001_d 0.00401408f $X=2.655 $Y=2.035 $X2=0 $Y2=0
cc_126 N_B_M1003_g N_VPWR_c_261_n 0.00306788f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_127 N_B_M1008_g N_VPWR_c_262_n 4.42323e-19 $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_128 N_B_M1008_g N_VPWR_c_264_n 0.00516461f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_129 N_B_c_115_n N_VPWR_c_264_n 0.0051298f $X=2.74 $Y=1.95 $X2=0 $Y2=0
cc_130 N_B_c_116_n N_VPWR_c_264_n 0.005819f $X=2.9 $Y=1.485 $X2=0 $Y2=0
cc_131 N_B_c_117_n N_VPWR_c_264_n 0.0016074f $X=2.9 $Y=1.485 $X2=0 $Y2=0
cc_132 N_B_M1003_g N_VPWR_c_266_n 0.005209f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_133 N_B_M1008_g N_VPWR_c_267_n 0.005209f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_134 N_B_M1003_g N_VPWR_c_258_n 0.0098299f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_135 N_B_M1008_g N_VPWR_c_258_n 0.00986118f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_136 N_B_c_164_p N_Y_M1003_d 0.0017721f $X=1.795 $Y=2.035 $X2=0 $Y2=0
cc_137 N_B_c_134_p N_Y_M1006_s 0.00554514f $X=2.655 $Y=2.035 $X2=0 $Y2=0
cc_138 N_B_c_115_n N_Y_M1006_s 0.00125604f $X=2.74 $Y=1.95 $X2=0 $Y2=0
cc_139 N_B_M1003_g N_Y_c_315_n 5.29656e-19 $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_140 N_B_M1007_g N_Y_c_312_n 0.0112384f $X=1.34 $Y=0.74 $X2=0 $Y2=0
cc_141 N_B_c_118_n N_Y_c_312_n 0.00499274f $X=1.43 $Y=1.515 $X2=0 $Y2=0
cc_142 N_B_c_119_n N_Y_c_312_n 0.0363457f $X=1.61 $Y=1.68 $X2=0 $Y2=0
cc_143 N_B_M1003_g N_Y_c_342_n 0.0133934f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_144 N_B_c_164_p N_Y_c_342_n 0.00683016f $X=1.795 $Y=2.035 $X2=0 $Y2=0
cc_145 N_B_c_118_n N_Y_c_342_n 3.20903e-19 $X=1.43 $Y=1.515 $X2=0 $Y2=0
cc_146 N_B_c_119_n N_Y_c_342_n 0.00330994f $X=1.61 $Y=1.68 $X2=0 $Y2=0
cc_147 N_B_c_134_p N_Y_c_346_n 0.0372379f $X=2.655 $Y=2.035 $X2=0 $Y2=0
cc_148 N_B_M1008_g N_Y_c_347_n 0.00254123f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_149 N_B_c_134_p N_Y_c_347_n 0.0153976f $X=2.655 $Y=2.035 $X2=0 $Y2=0
cc_150 N_B_M1008_g N_Y_c_316_n 0.00741984f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_151 N_B_M1007_g N_Y_c_313_n 0.00348765f $X=1.34 $Y=0.74 $X2=0 $Y2=0
cc_152 N_B_M1003_g N_Y_c_313_n 0.00251758f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_153 B N_Y_c_313_n 0.00985453f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_154 N_B_c_118_n N_Y_c_313_n 7.50286e-19 $X=1.43 $Y=1.515 $X2=0 $Y2=0
cc_155 N_B_c_119_n N_Y_c_313_n 0.0192485f $X=1.61 $Y=1.68 $X2=0 $Y2=0
cc_156 N_B_M1007_g N_Y_c_314_n 7.95487e-19 $X=1.34 $Y=0.74 $X2=0 $Y2=0
cc_157 N_B_M1009_g N_Y_c_314_n 0.00117715f $X=2.88 $Y=0.795 $X2=0 $Y2=0
cc_158 N_B_M1003_g Y 0.00915327f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_159 N_B_c_134_p Y 0.00186441f $X=2.655 $Y=2.035 $X2=0 $Y2=0
cc_160 N_B_c_164_p Y 0.016847f $X=1.795 $Y=2.035 $X2=0 $Y2=0
cc_161 N_B_M1007_g N_A_27_74#_c_409_n 0.00503198f $X=1.34 $Y=0.74 $X2=0 $Y2=0
cc_162 N_B_M1009_g N_A_27_74#_c_409_n 0.010205f $X=2.88 $Y=0.795 $X2=0 $Y2=0
cc_163 N_B_c_116_n N_A_27_74#_c_409_n 0.00722399f $X=2.9 $Y=1.485 $X2=0 $Y2=0
cc_164 N_B_c_117_n N_A_27_74#_c_409_n 0.00109429f $X=2.9 $Y=1.485 $X2=0 $Y2=0
cc_165 N_B_M1007_g N_A_27_74#_c_398_n 0.00980692f $X=1.34 $Y=0.74 $X2=0 $Y2=0
cc_166 N_B_M1009_g N_A_27_74#_c_399_n 0.0138289f $X=2.88 $Y=0.795 $X2=0 $Y2=0
cc_167 N_B_c_116_n N_A_27_74#_c_399_n 0.00838142f $X=2.9 $Y=1.485 $X2=0 $Y2=0
cc_168 N_B_c_117_n N_A_27_74#_c_399_n 0.00238884f $X=2.9 $Y=1.485 $X2=0 $Y2=0
cc_169 N_B_M1007_g N_VGND_c_455_n 3.89995e-19 $X=1.34 $Y=0.74 $X2=0 $Y2=0
cc_170 N_B_M1007_g N_VGND_c_457_n 0.00321733f $X=1.34 $Y=0.74 $X2=0 $Y2=0
cc_171 N_B_M1009_g N_VGND_c_457_n 0.00407143f $X=2.88 $Y=0.795 $X2=0 $Y2=0
cc_172 N_B_M1007_g N_VGND_c_458_n 0.00409122f $X=1.34 $Y=0.74 $X2=0 $Y2=0
cc_173 N_B_M1009_g N_VGND_c_458_n 0.00528353f $X=2.88 $Y=0.795 $X2=0 $Y2=0
cc_174 N_B_M1007_g N_A_283_74#_c_495_n 0.00260352f $X=1.34 $Y=0.74 $X2=0 $Y2=0
cc_175 N_B_M1009_g N_A_283_74#_c_495_n 0.00391613f $X=2.88 $Y=0.795 $X2=0 $Y2=0
cc_176 N_A_M1001_g N_VPWR_c_262_n 0.00336059f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_177 N_A_M1006_g N_VPWR_c_262_n 0.00866323f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_178 N_A_M1001_g N_VPWR_c_266_n 0.00526565f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_179 N_A_M1006_g N_VPWR_c_267_n 0.00460063f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_180 N_A_M1001_g N_VPWR_c_258_n 0.0100042f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A_M1006_g N_VPWR_c_258_n 0.00908665f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_182 N_A_M1002_g N_Y_c_312_n 0.013508f $X=1.895 $Y=0.795 $X2=0 $Y2=0
cc_183 N_A_M1001_g N_Y_c_346_n 0.0133251f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_184 N_A_M1006_g N_Y_c_346_n 0.0142879f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_185 N_A_M1006_g N_Y_c_316_n 3.78614e-19 $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_186 N_A_M1002_g N_Y_c_314_n 0.00643082f $X=1.895 $Y=0.795 $X2=0 $Y2=0
cc_187 N_A_M1011_g N_Y_c_314_n 0.00830615f $X=2.325 $Y=0.795 $X2=0 $Y2=0
cc_188 N_A_c_209_n N_Y_c_314_n 0.0245791f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_189 N_A_c_206_n N_Y_c_314_n 0.00263554f $X=2.405 $Y=1.515 $X2=0 $Y2=0
cc_190 N_A_M1001_g Y 0.0084443f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_191 N_A_M1006_g Y 8.11972e-19 $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_192 N_A_M1002_g N_A_27_74#_c_409_n 0.0117007f $X=1.895 $Y=0.795 $X2=0 $Y2=0
cc_193 N_A_M1011_g N_A_27_74#_c_409_n 0.0145843f $X=2.325 $Y=0.795 $X2=0 $Y2=0
cc_194 N_A_c_209_n N_A_27_74#_c_409_n 4.60142e-19 $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_195 N_A_c_206_n N_A_27_74#_c_409_n 0.0019193f $X=2.405 $Y=1.515 $X2=0 $Y2=0
cc_196 N_A_M1002_g N_A_27_74#_c_398_n 8.11839e-19 $X=1.895 $Y=0.795 $X2=0 $Y2=0
cc_197 N_A_M1011_g N_A_27_74#_c_399_n 0.00223206f $X=2.325 $Y=0.795 $X2=0 $Y2=0
cc_198 N_A_M1002_g N_VGND_c_457_n 8.63546e-19 $X=1.895 $Y=0.795 $X2=0 $Y2=0
cc_199 N_A_M1011_g N_VGND_c_457_n 8.63546e-19 $X=2.325 $Y=0.795 $X2=0 $Y2=0
cc_200 N_A_M1002_g N_A_283_74#_c_495_n 0.00941316f $X=1.895 $Y=0.795 $X2=0 $Y2=0
cc_201 N_A_M1011_g N_A_283_74#_c_495_n 0.00942684f $X=2.325 $Y=0.795 $X2=0 $Y2=0
cc_202 N_VPWR_c_261_n N_Y_c_315_n 0.0138908f $X=1.23 $Y=2.795 $X2=0 $Y2=0
cc_203 N_VPWR_c_265_n N_Y_c_315_n 0.0144623f $X=1.065 $Y=3.33 $X2=0 $Y2=0
cc_204 N_VPWR_c_258_n N_Y_c_315_n 0.0118344f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_205 N_VPWR_M1005_s N_Y_c_342_n 0.00915485f $X=1.045 $Y=1.84 $X2=0 $Y2=0
cc_206 N_VPWR_c_261_n N_Y_c_342_n 0.0167599f $X=1.23 $Y=2.795 $X2=0 $Y2=0
cc_207 N_VPWR_M1001_d N_Y_c_346_n 0.00415867f $X=2 $Y=1.84 $X2=0 $Y2=0
cc_208 N_VPWR_c_262_n N_Y_c_346_n 0.01852f $X=2.18 $Y=2.795 $X2=0 $Y2=0
cc_209 N_VPWR_c_262_n N_Y_c_316_n 0.0132809f $X=2.18 $Y=2.795 $X2=0 $Y2=0
cc_210 N_VPWR_c_264_n N_Y_c_316_n 0.017257f $X=3.08 $Y=1.985 $X2=0 $Y2=0
cc_211 N_VPWR_c_267_n N_Y_c_316_n 0.0118843f $X=2.995 $Y=3.33 $X2=0 $Y2=0
cc_212 N_VPWR_c_258_n N_Y_c_316_n 0.0097632f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_213 N_VPWR_c_260_n N_Y_c_317_n 0.04112f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_214 N_VPWR_c_261_n Y 0.0122069f $X=1.23 $Y=2.795 $X2=0 $Y2=0
cc_215 N_VPWR_c_262_n Y 0.0139233f $X=2.18 $Y=2.795 $X2=0 $Y2=0
cc_216 N_VPWR_c_266_n Y 0.0144926f $X=2.015 $Y=3.33 $X2=0 $Y2=0
cc_217 N_VPWR_c_258_n Y 0.0118645f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_218 N_VPWR_c_264_n N_A_27_74#_c_399_n 0.00608804f $X=3.08 $Y=1.985 $X2=0
+ $Y2=0
cc_219 N_Y_c_312_n N_A_27_74#_M1010_d 0.00119058f $X=1.945 $Y=1.175 $X2=0 $Y2=0
cc_220 N_Y_c_322_n N_A_27_74#_M1010_d 5.86511e-19 $X=1.095 $Y=1.175 $X2=0 $Y2=0
cc_221 N_Y_c_322_n N_A_27_74#_c_401_n 0.00453647f $X=1.095 $Y=1.175 $X2=0 $Y2=0
cc_222 N_Y_M1002_s N_A_27_74#_c_409_n 0.003356f $X=1.97 $Y=0.425 $X2=0 $Y2=0
cc_223 N_Y_c_312_n N_A_27_74#_c_409_n 0.0199657f $X=1.945 $Y=1.175 $X2=0 $Y2=0
cc_224 N_Y_c_314_n N_A_27_74#_c_409_n 0.0160991f $X=2.11 $Y=1.02 $X2=0 $Y2=0
cc_225 N_Y_c_312_n N_A_27_74#_c_398_n 0.0165421f $X=1.945 $Y=1.175 $X2=0 $Y2=0
cc_226 N_Y_c_322_n N_A_27_74#_c_398_n 0.00472879f $X=1.095 $Y=1.175 $X2=0 $Y2=0
cc_227 N_Y_c_314_n N_A_27_74#_c_399_n 0.00523618f $X=2.11 $Y=1.02 $X2=0 $Y2=0
cc_228 N_Y_c_312_n N_A_283_74#_M1007_d 0.00437664f $X=1.945 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_229 N_A_27_74#_c_401_n N_VGND_M1000_s 0.00447978f $X=1.04 $Y=0.835 $X2=-0.19
+ $Y2=-0.245
cc_230 N_A_27_74#_c_396_n N_VGND_c_455_n 0.00897147f $X=0.265 $Y=0.515 $X2=0
+ $Y2=0
cc_231 N_A_27_74#_c_401_n N_VGND_c_455_n 0.0165203f $X=1.04 $Y=0.835 $X2=0 $Y2=0
cc_232 N_A_27_74#_c_398_n N_VGND_c_455_n 0.0104177f $X=1.205 $Y=0.68 $X2=0 $Y2=0
cc_233 N_A_27_74#_c_396_n N_VGND_c_456_n 0.0110419f $X=0.265 $Y=0.515 $X2=0
+ $Y2=0
cc_234 N_A_27_74#_c_401_n N_VGND_c_456_n 0.00125985f $X=1.04 $Y=0.835 $X2=0
+ $Y2=0
cc_235 N_A_27_74#_c_397_n N_VGND_c_456_n 7.09218e-19 $X=0.265 $Y=0.835 $X2=0
+ $Y2=0
cc_236 N_A_27_74#_c_401_n N_VGND_c_457_n 0.00197156f $X=1.04 $Y=0.835 $X2=0
+ $Y2=0
cc_237 N_A_27_74#_c_409_n N_VGND_c_457_n 0.00390932f $X=2.93 $Y=0.68 $X2=0 $Y2=0
cc_238 N_A_27_74#_c_398_n N_VGND_c_457_n 0.0107219f $X=1.205 $Y=0.68 $X2=0 $Y2=0
cc_239 N_A_27_74#_c_399_n N_VGND_c_457_n 0.0117675f $X=3.095 $Y=0.57 $X2=0 $Y2=0
cc_240 N_A_27_74#_c_396_n N_VGND_c_458_n 0.00915013f $X=0.265 $Y=0.515 $X2=0
+ $Y2=0
cc_241 N_A_27_74#_c_401_n N_VGND_c_458_n 0.00743138f $X=1.04 $Y=0.835 $X2=0
+ $Y2=0
cc_242 N_A_27_74#_c_409_n N_VGND_c_458_n 0.00964348f $X=2.93 $Y=0.68 $X2=0 $Y2=0
cc_243 N_A_27_74#_c_397_n N_VGND_c_458_n 0.00196697f $X=0.265 $Y=0.835 $X2=0
+ $Y2=0
cc_244 N_A_27_74#_c_398_n N_VGND_c_458_n 0.0106167f $X=1.205 $Y=0.68 $X2=0 $Y2=0
cc_245 N_A_27_74#_c_399_n N_VGND_c_458_n 0.0116783f $X=3.095 $Y=0.57 $X2=0 $Y2=0
cc_246 N_A_27_74#_c_409_n N_A_283_74#_M1007_d 0.00737496f $X=2.93 $Y=0.68
+ $X2=-0.19 $Y2=-0.245
cc_247 N_A_27_74#_c_409_n N_A_283_74#_M1011_d 0.0118482f $X=2.93 $Y=0.68 $X2=0
+ $Y2=0
cc_248 N_A_27_74#_c_409_n N_A_283_74#_c_495_n 0.0797775f $X=2.93 $Y=0.68 $X2=0
+ $Y2=0
cc_249 N_A_27_74#_c_398_n N_A_283_74#_c_495_n 0.0025548f $X=1.205 $Y=0.68 $X2=0
+ $Y2=0
cc_250 N_A_27_74#_c_399_n N_A_283_74#_c_495_n 0.00153676f $X=3.095 $Y=0.57 $X2=0
+ $Y2=0
cc_251 N_VGND_c_458_n N_A_283_74#_M1007_d 0.00230295f $X=3.12 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_252 N_VGND_c_458_n N_A_283_74#_M1011_d 0.00247946f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_253 N_VGND_c_455_n N_A_283_74#_c_495_n 0.00240443f $X=0.695 $Y=0.495 $X2=0
+ $Y2=0
cc_254 N_VGND_c_457_n N_A_283_74#_c_495_n 0.0838614f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_255 N_VGND_c_458_n N_A_283_74#_c_495_n 0.0492532f $X=3.12 $Y=0 $X2=0 $Y2=0

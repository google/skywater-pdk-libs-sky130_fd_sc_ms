* File: sky130_fd_sc_ms__clkdlyinv5sd1_1.spice
* Created: Wed Sep  2 12:01:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__clkdlyinv5sd1_1.pex.spice"
.subckt sky130_fd_sc_ms__clkdlyinv5sd1_1  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_A_M1007_g N_A_28_74#_M1007_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.15435 AS=0.1113 PD=1.155 PS=1.37 NRD=15.708 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1009 N_A_288_74#_M1009_d N_A_28_74#_M1009_g N_VGND_M1007_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.1113 AS=0.15435 PD=1.37 PS=1.155 NRD=0 NRS=114.276 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_A_549_74#_M1001_d N_A_288_74#_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.1113 AS=0.2604 PD=1.37 PS=2.08 NRD=0 NRS=99.996 M=1 R=2.8
+ SA=75000.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_549_74#_M1004_g N_A_682_74#_M1004_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0966 AS=0.2583 PD=0.88 PS=2.07 NRD=51.42 NRS=99.996 M=1 R=2.8
+ SA=75000.5 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_A_682_74#_M1002_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0966 PD=1.37 PS=0.88 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_A_28_74#_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.390943 AS=0.2968 PD=1.93358 PS=2.77 NRD=2.6201 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90000.9 A=0.2016 P=2.6 MULT=1
MM1005 N_A_288_74#_M1005_d N_A_28_74#_M1005_g N_VPWR_M1006_d VPB PSHORT L=0.15
+ W=1 AD=0.26 AS=0.349057 PD=2.52 PS=1.72642 NRD=0 NRS=81.7353 M=1 R=6.66667
+ SA=75001.1 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1000 N_A_549_74#_M1000_d N_A_288_74#_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.15
+ W=1 AD=0.265 AS=0.62 PD=2.53 PS=3.24 NRD=0 NRS=69.9153 M=1 R=6.66667
+ SA=75000.5 SB=75000.2 A=0.15 P=2.3 MULT=1
MM1003 N_VPWR_M1003_d N_A_549_74#_M1003_g N_A_682_74#_M1003_s VPB PSHORT L=0.15
+ W=1 AD=0.231698 AS=0.61 PD=1.49057 PS=3.22 NRD=36.7602 NRS=67.9453 M=1
+ R=6.66667 SA=75000.5 SB=75000.8 A=0.15 P=2.3 MULT=1
MM1008 N_Y_M1008_d N_A_682_74#_M1008_g N_VPWR_M1003_d VPB PSHORT L=0.18 W=1.12
+ AD=0.2968 AS=0.259502 PD=2.77 PS=1.66943 NRD=0 NRS=0 M=1 R=6.22222 SA=90001
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=10.5276 P=15.04
*
.include "sky130_fd_sc_ms__clkdlyinv5sd1_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__ebufn_4.pxi.spice
* Created: Fri Aug 28 17:32:03 2020
* 
x_PM_SKY130_FD_SC_MS__EBUFN_4%A N_A_M1006_g N_A_M1004_g A N_A_c_131_n
+ PM_SKY130_FD_SC_MS__EBUFN_4%A
x_PM_SKY130_FD_SC_MS__EBUFN_4%TE_B N_TE_B_M1011_g N_TE_B_c_163_n N_TE_B_c_175_n
+ N_TE_B_M1001_g N_TE_B_c_164_n N_TE_B_c_177_n N_TE_B_M1013_g N_TE_B_c_165_n
+ N_TE_B_c_179_n N_TE_B_M1016_g N_TE_B_c_166_n N_TE_B_c_181_n N_TE_B_M1017_g
+ N_TE_B_c_167_n N_TE_B_c_183_n N_TE_B_M1019_g N_TE_B_c_168_n N_TE_B_c_169_n
+ N_TE_B_c_170_n N_TE_B_c_171_n TE_B N_TE_B_c_173_n N_TE_B_c_174_n
+ PM_SKY130_FD_SC_MS__EBUFN_4%TE_B
x_PM_SKY130_FD_SC_MS__EBUFN_4%A_208_74# N_A_208_74#_M1011_d N_A_208_74#_M1001_d
+ N_A_208_74#_c_282_n N_A_208_74#_c_283_n N_A_208_74#_c_284_n
+ N_A_208_74#_M1007_g N_A_208_74#_c_285_n N_A_208_74#_c_286_n
+ N_A_208_74#_M1008_g N_A_208_74#_c_287_n N_A_208_74#_c_288_n
+ N_A_208_74#_M1009_g N_A_208_74#_c_289_n N_A_208_74#_c_290_n
+ N_A_208_74#_M1015_g N_A_208_74#_c_291_n N_A_208_74#_c_292_n
+ N_A_208_74#_c_293_n N_A_208_74#_c_298_n N_A_208_74#_c_297_n
+ N_A_208_74#_c_294_n N_A_208_74#_c_295_n N_A_208_74#_c_296_n
+ PM_SKY130_FD_SC_MS__EBUFN_4%A_208_74#
x_PM_SKY130_FD_SC_MS__EBUFN_4%A_27_368# N_A_27_368#_M1004_s N_A_27_368#_M1006_s
+ N_A_27_368#_M1000_g N_A_27_368#_M1005_g N_A_27_368#_M1002_g
+ N_A_27_368#_M1012_g N_A_27_368#_M1003_g N_A_27_368#_M1014_g
+ N_A_27_368#_M1010_g N_A_27_368#_M1018_g N_A_27_368#_c_397_n
+ N_A_27_368#_c_408_n N_A_27_368#_c_409_n N_A_27_368#_c_410_n
+ N_A_27_368#_c_411_n N_A_27_368#_c_412_n N_A_27_368#_c_413_n
+ N_A_27_368#_c_414_n N_A_27_368#_c_415_n N_A_27_368#_c_398_n
+ N_A_27_368#_c_399_n N_A_27_368#_c_505_p N_A_27_368#_c_400_n
+ N_A_27_368#_c_401_n N_A_27_368#_c_417_n N_A_27_368#_c_402_n
+ N_A_27_368#_c_403_n PM_SKY130_FD_SC_MS__EBUFN_4%A_27_368#
x_PM_SKY130_FD_SC_MS__EBUFN_4%VPWR N_VPWR_M1006_d N_VPWR_M1013_d N_VPWR_M1017_d
+ N_VPWR_c_557_n N_VPWR_c_558_n N_VPWR_c_559_n N_VPWR_c_560_n N_VPWR_c_561_n
+ N_VPWR_c_562_n VPWR N_VPWR_c_563_n N_VPWR_c_564_n N_VPWR_c_556_n
+ N_VPWR_c_566_n N_VPWR_c_567_n PM_SKY130_FD_SC_MS__EBUFN_4%VPWR
x_PM_SKY130_FD_SC_MS__EBUFN_4%A_348_368# N_A_348_368#_M1013_s
+ N_A_348_368#_M1016_s N_A_348_368#_M1019_s N_A_348_368#_M1002_s
+ N_A_348_368#_M1010_s N_A_348_368#_c_635_n N_A_348_368#_c_626_n
+ N_A_348_368#_c_627_n N_A_348_368#_c_628_n N_A_348_368#_c_629_n
+ N_A_348_368#_c_644_n N_A_348_368#_c_630_n N_A_348_368#_c_631_n
+ N_A_348_368#_c_688_p N_A_348_368#_c_632_n N_A_348_368#_c_633_n
+ N_A_348_368#_c_659_n N_A_348_368#_c_634_n
+ PM_SKY130_FD_SC_MS__EBUFN_4%A_348_368#
x_PM_SKY130_FD_SC_MS__EBUFN_4%Z N_Z_M1005_s N_Z_M1014_s N_Z_M1000_d N_Z_M1003_d
+ N_Z_c_695_n N_Z_c_699_n N_Z_c_707_n N_Z_c_696_n N_Z_c_691_n N_Z_c_692_n
+ N_Z_c_722_n N_Z_c_693_n N_Z_c_694_n Z Z Z PM_SKY130_FD_SC_MS__EBUFN_4%Z
x_PM_SKY130_FD_SC_MS__EBUFN_4%VGND N_VGND_M1004_d N_VGND_M1007_d N_VGND_M1009_d
+ N_VGND_c_758_n N_VGND_c_759_n N_VGND_c_760_n N_VGND_c_761_n N_VGND_c_762_n
+ N_VGND_c_763_n N_VGND_c_764_n VGND N_VGND_c_765_n N_VGND_c_766_n
+ N_VGND_c_767_n N_VGND_c_768_n PM_SKY130_FD_SC_MS__EBUFN_4%VGND
x_PM_SKY130_FD_SC_MS__EBUFN_4%A_378_74# N_A_378_74#_M1007_s N_A_378_74#_M1008_s
+ N_A_378_74#_M1015_s N_A_378_74#_M1012_d N_A_378_74#_M1018_d
+ N_A_378_74#_c_830_n N_A_378_74#_c_831_n N_A_378_74#_c_832_n
+ N_A_378_74#_c_833_n N_A_378_74#_c_834_n N_A_378_74#_c_865_n
+ N_A_378_74#_c_835_n N_A_378_74#_c_836_n N_A_378_74#_c_887_n
+ N_A_378_74#_c_837_n N_A_378_74#_c_838_n N_A_378_74#_c_839_n
+ N_A_378_74#_c_840_n PM_SKY130_FD_SC_MS__EBUFN_4%A_378_74#
cc_1 VNB N_A_M1006_g 0.00161385f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A_M1004_g 0.0263754f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.74
cc_3 VNB A 0.00396202f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_A_c_131_n 0.0341949f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.465
cc_5 VNB N_TE_B_c_163_n 0.014558f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.3
cc_6 VNB N_TE_B_c_164_n 0.0209946f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_7 VNB N_TE_B_c_165_n 0.00652849f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.3
cc_8 VNB N_TE_B_c_166_n 0.00551218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_TE_B_c_167_n 0.0103807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_TE_B_c_168_n 0.00469483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_TE_B_c_169_n 0.00491136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_TE_B_c_170_n 0.00369526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_TE_B_c_171_n 0.00369526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB TE_B 0.00702428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_TE_B_c_173_n 0.0182217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_TE_B_c_174_n 0.0192479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_208_74#_c_282_n 0.0205453f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.74
cc_18 VNB N_A_208_74#_c_283_n 0.011951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_208_74#_c_284_n 0.0166173f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_20 VNB N_A_208_74#_c_285_n 0.0122721f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.465
cc_21 VNB N_A_208_74#_c_286_n 0.01433f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.3
cc_22 VNB N_A_208_74#_c_287_n 0.0122636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_208_74#_c_288_n 0.0143385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_208_74#_c_289_n 0.0200371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_208_74#_c_290_n 0.0146143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_208_74#_c_291_n 0.00514785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_208_74#_c_292_n 0.00511446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_208_74#_c_293_n 0.00511446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_208_74#_c_294_n 0.00848374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_208_74#_c_295_n 0.00568136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_208_74#_c_296_n 0.0754207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_368#_M1000_g 4.95336e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_33 VNB N_A_27_368#_M1005_g 0.0214935f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.465
cc_34 VNB N_A_27_368#_M1002_g 4.78697e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_368#_M1012_g 0.0209312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_27_368#_M1003_g 4.7662e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_368#_M1014_g 0.0211723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_368#_M1010_g 7.19436e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_368#_M1018_g 0.0285164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_27_368#_c_397_n 0.0280304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_368#_c_398_n 0.0025686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_27_368#_c_399_n 0.00606935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_27_368#_c_400_n 0.0112533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_27_368#_c_401_n 0.0248753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_27_368#_c_402_n 0.0135381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_27_368#_c_403_n 0.0982087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VPWR_c_556_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_Z_c_691_n 0.00225436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_Z_c_692_n 0.00229628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_Z_c_693_n 0.00122079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_Z_c_694_n 0.00176823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_758_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.465
cc_53 VNB N_VGND_c_759_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.54
cc_54 VNB N_VGND_c_760_n 0.00452091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_761_n 0.0363752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_762_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_763_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_764_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_765_n 0.018117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_766_n 0.0569796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_767_n 0.328933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_768_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_378_74#_c_830_n 0.00221841f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.54
cc_64 VNB N_A_378_74#_c_831_n 0.0063992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_378_74#_c_832_n 2.51175e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_378_74#_c_833_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_378_74#_c_834_n 0.00578259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_378_74#_c_835_n 0.0027626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_378_74#_c_836_n 0.00163793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_378_74#_c_837_n 0.0122413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_378_74#_c_838_n 0.0364928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_378_74#_c_839_n 7.52762e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_378_74#_c_840_n 0.00121874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VPB N_A_M1006_g 0.0262218f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_75 VPB A 0.00440147f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_76 VPB N_TE_B_c_175_n 0.0240272f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=0.74
cc_77 VPB N_TE_B_c_164_n 0.0245338f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_78 VPB N_TE_B_c_177_n 0.0230458f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.465
cc_79 VPB N_TE_B_c_165_n 0.00414223f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.3
cc_80 VPB N_TE_B_c_179_n 0.0178168f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.54
cc_81 VPB N_TE_B_c_166_n 0.00378507f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_TE_B_c_181_n 0.0181086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_TE_B_c_167_n 0.0063045f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_TE_B_c_183_n 0.0185246f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_TE_B_c_168_n 0.00601664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_TE_B_c_169_n 0.00124171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_TE_B_c_170_n 0.00124171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_TE_B_c_171_n 0.00124171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_208_74#_c_297_n 0.00532438f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_27_368#_M1000_g 0.0218302f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_91 VPB N_A_27_368#_M1002_g 0.0213667f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_27_368#_M1003_g 0.0213413f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_27_368#_M1010_g 0.0280581f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_27_368#_c_408_n 0.00536733f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_27_368#_c_409_n 0.0114247f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_27_368#_c_410_n 0.0187341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_27_368#_c_411_n 0.00914426f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_27_368#_c_412_n 0.00464413f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_27_368#_c_413_n 0.00513674f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_27_368#_c_414_n 0.0034454f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_27_368#_c_415_n 0.00107523f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_27_368#_c_401_n 0.0127888f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_27_368#_c_417_n 0.00723806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_557_n 0.00396699f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.465
cc_105 VPB N_VPWR_c_558_n 0.00329129f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.54
cc_106 VPB N_VPWR_c_559_n 0.0157448f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.54
cc_107 VPB N_VPWR_c_560_n 0.00454608f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_561_n 0.0377381f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_562_n 0.00601619f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_563_n 0.017793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_564_n 0.0591139f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_556_n 0.0794015f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_566_n 0.00647446f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_567_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_348_368#_c_626_n 0.00123781f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.54
cc_116 VPB N_A_348_368#_c_627_n 0.00179594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_348_368#_c_628_n 0.0021546f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_348_368#_c_629_n 0.00207253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_348_368#_c_630_n 0.00240659f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_348_368#_c_631_n 0.00160153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_348_368#_c_632_n 0.0117115f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_348_368#_c_633_n 0.0503906f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_348_368#_c_634_n 0.00167433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_Z_c_695_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.465
cc_125 VPB N_Z_c_696_n 0.00219429f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_Z_c_693_n 0.00103298f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB Z 0.00176823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 N_A_M1006_g N_TE_B_c_168_n 0.0471889f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_129 N_A_M1004_g TE_B 6.22691e-19 $X=0.535 $Y=0.74 $X2=0 $Y2=0
cc_130 A TE_B 0.0199149f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_131 N_A_c_131_n TE_B 2.12581e-19 $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_132 A N_TE_B_c_173_n 0.00476272f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_133 N_A_c_131_n N_TE_B_c_173_n 0.0206413f $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_134 N_A_M1004_g N_TE_B_c_174_n 0.0159419f $X=0.535 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A_M1006_g N_A_208_74#_c_298_n 0.00111355f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_136 N_A_M1006_g N_A_208_74#_c_297_n 5.5862e-19 $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_137 A N_A_208_74#_c_297_n 0.00383597f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_138 A N_A_208_74#_c_294_n 0.0049962f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_139 N_A_M1004_g N_A_27_368#_c_397_n 0.00241184f $X=0.535 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A_c_131_n N_A_27_368#_c_408_n 4.06489e-19 $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_141 N_A_M1006_g N_A_27_368#_c_410_n 4.7096e-19 $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_142 N_A_M1006_g N_A_27_368#_c_411_n 0.0135793f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_143 A N_A_27_368#_c_411_n 0.010284f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_144 N_A_c_131_n N_A_27_368#_c_400_n 0.00239983f $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_145 N_A_M1006_g N_A_27_368#_c_401_n 0.00724244f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_146 N_A_M1004_g N_A_27_368#_c_401_n 0.0039401f $X=0.535 $Y=0.74 $X2=0 $Y2=0
cc_147 A N_A_27_368#_c_401_n 0.0364523f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_148 N_A_c_131_n N_A_27_368#_c_401_n 0.00809677f $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_149 N_A_M1006_g N_VPWR_c_557_n 0.0105027f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_150 N_A_M1006_g N_VPWR_c_563_n 0.00460063f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_151 N_A_M1006_g N_VPWR_c_556_n 0.00446988f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_152 N_A_M1004_g N_VGND_c_758_n 0.0144322f $X=0.535 $Y=0.74 $X2=0 $Y2=0
cc_153 A N_VGND_c_758_n 0.01106f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_154 N_A_c_131_n N_VGND_c_758_n 0.00129795f $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_155 N_A_M1004_g N_VGND_c_765_n 0.00383152f $X=0.535 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A_M1004_g N_VGND_c_767_n 0.00761327f $X=0.535 $Y=0.74 $X2=0 $Y2=0
cc_157 N_TE_B_c_169_n N_A_208_74#_c_282_n 0.0169843f $X=2.11 $Y=1.65 $X2=0 $Y2=0
cc_158 N_TE_B_c_164_n N_A_208_74#_c_283_n 0.0169843f $X=2.02 $Y=1.65 $X2=0 $Y2=0
cc_159 N_TE_B_c_173_n N_A_208_74#_c_283_n 0.00761709f $X=1.075 $Y=1.385 $X2=0
+ $Y2=0
cc_160 N_TE_B_c_170_n N_A_208_74#_c_285_n 0.0169843f $X=2.56 $Y=1.65 $X2=0 $Y2=0
cc_161 N_TE_B_c_171_n N_A_208_74#_c_287_n 0.0169843f $X=3.01 $Y=1.65 $X2=0 $Y2=0
cc_162 N_TE_B_c_165_n N_A_208_74#_c_291_n 0.0169843f $X=2.47 $Y=1.65 $X2=0 $Y2=0
cc_163 N_TE_B_c_166_n N_A_208_74#_c_292_n 0.0169843f $X=2.92 $Y=1.65 $X2=0 $Y2=0
cc_164 N_TE_B_c_167_n N_A_208_74#_c_293_n 0.0169843f $X=3.37 $Y=1.65 $X2=0 $Y2=0
cc_165 N_TE_B_c_175_n N_A_208_74#_c_298_n 0.00734906f $X=0.98 $Y=1.725 $X2=0
+ $Y2=0
cc_166 N_TE_B_c_168_n N_A_208_74#_c_298_n 6.38792e-19 $X=1.065 $Y=1.65 $X2=0
+ $Y2=0
cc_167 N_TE_B_c_175_n N_A_208_74#_c_297_n 0.0057782f $X=0.98 $Y=1.725 $X2=0
+ $Y2=0
cc_168 N_TE_B_c_164_n N_A_208_74#_c_297_n 0.0173987f $X=2.02 $Y=1.65 $X2=0 $Y2=0
cc_169 N_TE_B_c_177_n N_A_208_74#_c_297_n 0.00393075f $X=2.11 $Y=1.725 $X2=0
+ $Y2=0
cc_170 N_TE_B_c_168_n N_A_208_74#_c_297_n 0.00422564f $X=1.065 $Y=1.65 $X2=0
+ $Y2=0
cc_171 TE_B N_A_208_74#_c_297_n 0.0178111f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_172 N_TE_B_c_163_n N_A_208_74#_c_294_n 6.8085e-19 $X=1.065 $Y=1.575 $X2=0
+ $Y2=0
cc_173 N_TE_B_c_164_n N_A_208_74#_c_294_n 0.0163685f $X=2.02 $Y=1.65 $X2=0 $Y2=0
cc_174 TE_B N_A_208_74#_c_294_n 0.0298967f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_175 N_TE_B_c_173_n N_A_208_74#_c_294_n 0.00152275f $X=1.075 $Y=1.385 $X2=0
+ $Y2=0
cc_176 N_TE_B_c_174_n N_A_208_74#_c_294_n 9.11108e-19 $X=1.065 $Y=1.22 $X2=0
+ $Y2=0
cc_177 N_TE_B_c_164_n N_A_208_74#_c_295_n 0.0046517f $X=2.02 $Y=1.65 $X2=0 $Y2=0
cc_178 TE_B N_A_208_74#_c_295_n 0.0164997f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_179 N_TE_B_c_173_n N_A_208_74#_c_295_n 0.0010152f $X=1.075 $Y=1.385 $X2=0
+ $Y2=0
cc_180 N_TE_B_c_174_n N_A_208_74#_c_295_n 6.76457e-19 $X=1.065 $Y=1.22 $X2=0
+ $Y2=0
cc_181 TE_B N_A_208_74#_c_296_n 0.00107199f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_182 N_TE_B_c_174_n N_A_208_74#_c_296_n 0.016396f $X=1.065 $Y=1.22 $X2=0 $Y2=0
cc_183 N_TE_B_c_183_n N_A_27_368#_M1000_g 0.0111843f $X=3.46 $Y=1.725 $X2=0
+ $Y2=0
cc_184 N_TE_B_c_175_n N_A_27_368#_c_411_n 0.019433f $X=0.98 $Y=1.725 $X2=0 $Y2=0
cc_185 N_TE_B_c_164_n N_A_27_368#_c_411_n 8.33427e-19 $X=2.02 $Y=1.65 $X2=0
+ $Y2=0
cc_186 N_TE_B_c_175_n N_A_27_368#_c_412_n 0.00440223f $X=0.98 $Y=1.725 $X2=0
+ $Y2=0
cc_187 N_TE_B_c_177_n N_A_27_368#_c_412_n 0.0041232f $X=2.11 $Y=1.725 $X2=0
+ $Y2=0
cc_188 N_TE_B_c_164_n N_A_27_368#_c_413_n 0.00514557f $X=2.02 $Y=1.65 $X2=0
+ $Y2=0
cc_189 N_TE_B_c_177_n N_A_27_368#_c_413_n 0.0186182f $X=2.11 $Y=1.725 $X2=0
+ $Y2=0
cc_190 N_TE_B_c_165_n N_A_27_368#_c_413_n 0.00199579f $X=2.47 $Y=1.65 $X2=0
+ $Y2=0
cc_191 N_TE_B_c_179_n N_A_27_368#_c_413_n 0.0050995f $X=2.56 $Y=1.725 $X2=0
+ $Y2=0
cc_192 N_TE_B_c_175_n N_A_27_368#_c_414_n 6.66989e-19 $X=0.98 $Y=1.725 $X2=0
+ $Y2=0
cc_193 N_TE_B_c_164_n N_A_27_368#_c_414_n 8.92373e-19 $X=2.02 $Y=1.65 $X2=0
+ $Y2=0
cc_194 N_TE_B_c_177_n N_A_27_368#_c_415_n 0.0051974f $X=2.11 $Y=1.725 $X2=0
+ $Y2=0
cc_195 N_TE_B_c_165_n N_A_27_368#_c_415_n 0.00303973f $X=2.47 $Y=1.65 $X2=0
+ $Y2=0
cc_196 N_TE_B_c_179_n N_A_27_368#_c_415_n 0.00711f $X=2.56 $Y=1.725 $X2=0 $Y2=0
cc_197 N_TE_B_c_181_n N_A_27_368#_c_415_n 5.38945e-19 $X=3.01 $Y=1.725 $X2=0
+ $Y2=0
cc_198 N_TE_B_c_170_n N_A_27_368#_c_415_n 0.0036841f $X=2.56 $Y=1.65 $X2=0 $Y2=0
cc_199 N_TE_B_c_165_n N_A_27_368#_c_398_n 0.00346529f $X=2.47 $Y=1.65 $X2=0
+ $Y2=0
cc_200 N_TE_B_c_170_n N_A_27_368#_c_398_n 7.22911e-19 $X=2.56 $Y=1.65 $X2=0
+ $Y2=0
cc_201 N_TE_B_c_166_n N_A_27_368#_c_402_n 0.00776016f $X=2.92 $Y=1.65 $X2=0
+ $Y2=0
cc_202 N_TE_B_c_167_n N_A_27_368#_c_402_n 0.0117412f $X=3.37 $Y=1.65 $X2=0 $Y2=0
cc_203 N_TE_B_c_170_n N_A_27_368#_c_402_n 0.00668245f $X=2.56 $Y=1.65 $X2=0
+ $Y2=0
cc_204 N_TE_B_c_171_n N_A_27_368#_c_402_n 0.0046055f $X=3.01 $Y=1.65 $X2=0 $Y2=0
cc_205 N_TE_B_c_167_n N_A_27_368#_c_403_n 0.0111843f $X=3.37 $Y=1.65 $X2=0 $Y2=0
cc_206 N_TE_B_c_175_n N_VPWR_c_557_n 0.0184935f $X=0.98 $Y=1.725 $X2=0 $Y2=0
cc_207 N_TE_B_c_177_n N_VPWR_c_558_n 0.0153136f $X=2.11 $Y=1.725 $X2=0 $Y2=0
cc_208 N_TE_B_c_179_n N_VPWR_c_558_n 0.00743975f $X=2.56 $Y=1.725 $X2=0 $Y2=0
cc_209 N_TE_B_c_181_n N_VPWR_c_558_n 3.98916e-19 $X=3.01 $Y=1.725 $X2=0 $Y2=0
cc_210 N_TE_B_c_179_n N_VPWR_c_559_n 0.00338459f $X=2.56 $Y=1.725 $X2=0 $Y2=0
cc_211 N_TE_B_c_181_n N_VPWR_c_559_n 0.00460063f $X=3.01 $Y=1.725 $X2=0 $Y2=0
cc_212 N_TE_B_c_179_n N_VPWR_c_560_n 4.54258e-19 $X=2.56 $Y=1.725 $X2=0 $Y2=0
cc_213 N_TE_B_c_181_n N_VPWR_c_560_n 0.0148175f $X=3.01 $Y=1.725 $X2=0 $Y2=0
cc_214 N_TE_B_c_183_n N_VPWR_c_560_n 0.00169232f $X=3.46 $Y=1.725 $X2=0 $Y2=0
cc_215 N_TE_B_c_175_n N_VPWR_c_561_n 0.00460063f $X=0.98 $Y=1.725 $X2=0 $Y2=0
cc_216 N_TE_B_c_177_n N_VPWR_c_561_n 0.00338459f $X=2.11 $Y=1.725 $X2=0 $Y2=0
cc_217 N_TE_B_c_183_n N_VPWR_c_564_n 0.00517089f $X=3.46 $Y=1.725 $X2=0 $Y2=0
cc_218 N_TE_B_c_175_n N_VPWR_c_556_n 0.0044838f $X=0.98 $Y=1.725 $X2=0 $Y2=0
cc_219 N_TE_B_c_177_n N_VPWR_c_556_n 0.0044586f $X=2.11 $Y=1.725 $X2=0 $Y2=0
cc_220 N_TE_B_c_179_n N_VPWR_c_556_n 0.00440727f $X=2.56 $Y=1.725 $X2=0 $Y2=0
cc_221 N_TE_B_c_181_n N_VPWR_c_556_n 0.00908554f $X=3.01 $Y=1.725 $X2=0 $Y2=0
cc_222 N_TE_B_c_183_n N_VPWR_c_556_n 0.00977588f $X=3.46 $Y=1.725 $X2=0 $Y2=0
cc_223 N_TE_B_c_177_n N_A_348_368#_c_635_n 0.011349f $X=2.11 $Y=1.725 $X2=0
+ $Y2=0
cc_224 N_TE_B_c_179_n N_A_348_368#_c_635_n 0.0149673f $X=2.56 $Y=1.725 $X2=0
+ $Y2=0
cc_225 N_TE_B_c_166_n N_A_348_368#_c_626_n 0.00197117f $X=2.92 $Y=1.65 $X2=0
+ $Y2=0
cc_226 N_TE_B_c_179_n N_A_348_368#_c_627_n 2.55042e-19 $X=2.56 $Y=1.725 $X2=0
+ $Y2=0
cc_227 N_TE_B_c_181_n N_A_348_368#_c_627_n 2.55042e-19 $X=3.01 $Y=1.725 $X2=0
+ $Y2=0
cc_228 N_TE_B_c_181_n N_A_348_368#_c_628_n 0.0142554f $X=3.01 $Y=1.725 $X2=0
+ $Y2=0
cc_229 N_TE_B_c_167_n N_A_348_368#_c_628_n 0.00187989f $X=3.37 $Y=1.65 $X2=0
+ $Y2=0
cc_230 N_TE_B_c_183_n N_A_348_368#_c_628_n 0.0127914f $X=3.46 $Y=1.725 $X2=0
+ $Y2=0
cc_231 N_TE_B_c_183_n N_A_348_368#_c_629_n 0.00104546f $X=3.46 $Y=1.725 $X2=0
+ $Y2=0
cc_232 N_TE_B_c_181_n N_A_348_368#_c_644_n 7.27629e-19 $X=3.01 $Y=1.725 $X2=0
+ $Y2=0
cc_233 N_TE_B_c_183_n N_A_348_368#_c_644_n 0.0127108f $X=3.46 $Y=1.725 $X2=0
+ $Y2=0
cc_234 N_TE_B_c_183_n N_A_348_368#_c_631_n 0.00347836f $X=3.46 $Y=1.725 $X2=0
+ $Y2=0
cc_235 N_TE_B_c_183_n N_Z_c_699_n 2.5626e-19 $X=3.46 $Y=1.725 $X2=0 $Y2=0
cc_236 N_TE_B_c_174_n N_VGND_c_758_n 0.0133028f $X=1.065 $Y=1.22 $X2=0 $Y2=0
cc_237 N_TE_B_c_174_n N_VGND_c_761_n 0.00383152f $X=1.065 $Y=1.22 $X2=0 $Y2=0
cc_238 N_TE_B_c_174_n N_VGND_c_767_n 0.00762539f $X=1.065 $Y=1.22 $X2=0 $Y2=0
cc_239 N_TE_B_c_165_n N_A_378_74#_c_831_n 4.52625e-19 $X=2.47 $Y=1.65 $X2=0
+ $Y2=0
cc_240 N_TE_B_c_169_n N_A_378_74#_c_831_n 0.0016808f $X=2.11 $Y=1.65 $X2=0 $Y2=0
cc_241 N_TE_B_c_164_n N_A_378_74#_c_832_n 0.00120343f $X=2.02 $Y=1.65 $X2=0
+ $Y2=0
cc_242 N_TE_B_c_167_n N_A_378_74#_c_834_n 6.28703e-19 $X=3.37 $Y=1.65 $X2=0
+ $Y2=0
cc_243 N_TE_B_c_171_n N_A_378_74#_c_834_n 2.85891e-19 $X=3.01 $Y=1.65 $X2=0
+ $Y2=0
cc_244 N_A_208_74#_c_290_n N_A_27_368#_M1005_g 0.0193926f $X=3.535 $Y=1.185
+ $X2=0 $Y2=0
cc_245 N_A_208_74#_M1001_d N_A_27_368#_c_411_n 0.0077488f $X=1.07 $Y=1.84 $X2=0
+ $Y2=0
cc_246 N_A_208_74#_c_298_n N_A_27_368#_c_411_n 0.0145226f $X=1.205 $Y=2.02 $X2=0
+ $Y2=0
cc_247 N_A_208_74#_c_297_n N_A_27_368#_c_411_n 0.00592951f $X=1.615 $Y=1.72
+ $X2=0 $Y2=0
cc_248 N_A_208_74#_c_297_n N_A_27_368#_c_413_n 0.0107872f $X=1.615 $Y=1.72 $X2=0
+ $Y2=0
cc_249 N_A_208_74#_c_298_n N_A_27_368#_c_414_n 0.0136473f $X=1.205 $Y=2.02 $X2=0
+ $Y2=0
cc_250 N_A_208_74#_c_297_n N_A_27_368#_c_414_n 0.0139991f $X=1.615 $Y=1.72 $X2=0
+ $Y2=0
cc_251 N_A_208_74#_c_297_n N_A_27_368#_c_415_n 0.00574523f $X=1.615 $Y=1.72
+ $X2=0 $Y2=0
cc_252 N_A_208_74#_c_294_n N_A_27_368#_c_415_n 0.00178624f $X=1.615 $Y=1.145
+ $X2=0 $Y2=0
cc_253 N_A_208_74#_c_285_n N_A_27_368#_c_398_n 0.00115704f $X=2.6 $Y=1.26 $X2=0
+ $Y2=0
cc_254 N_A_208_74#_c_294_n N_A_27_368#_c_398_n 0.00569129f $X=1.615 $Y=1.145
+ $X2=0 $Y2=0
cc_255 N_A_208_74#_c_285_n N_A_27_368#_c_402_n 0.00936976f $X=2.6 $Y=1.26 $X2=0
+ $Y2=0
cc_256 N_A_208_74#_c_289_n N_A_27_368#_c_403_n 0.0010213f $X=3.46 $Y=1.26 $X2=0
+ $Y2=0
cc_257 N_A_208_74#_c_297_n N_A_348_368#_M1013_s 0.00111748f $X=1.615 $Y=1.72
+ $X2=-0.19 $Y2=-0.245
cc_258 N_A_208_74#_c_295_n N_VGND_c_758_n 0.0285331f $X=1.615 $Y=0.465 $X2=0
+ $Y2=0
cc_259 N_A_208_74#_c_296_n N_VGND_c_758_n 4.72719e-19 $X=1.615 $Y=0.465 $X2=0
+ $Y2=0
cc_260 N_A_208_74#_c_284_n N_VGND_c_759_n 0.0122493f $X=2.245 $Y=1.185 $X2=0
+ $Y2=0
cc_261 N_A_208_74#_c_285_n N_VGND_c_759_n 7.11061e-19 $X=2.6 $Y=1.26 $X2=0 $Y2=0
cc_262 N_A_208_74#_c_286_n N_VGND_c_759_n 0.0106722f $X=2.675 $Y=1.185 $X2=0
+ $Y2=0
cc_263 N_A_208_74#_c_288_n N_VGND_c_759_n 5.10431e-19 $X=3.105 $Y=1.185 $X2=0
+ $Y2=0
cc_264 N_A_208_74#_c_295_n N_VGND_c_759_n 0.00156286f $X=1.615 $Y=0.465 $X2=0
+ $Y2=0
cc_265 N_A_208_74#_c_296_n N_VGND_c_759_n 3.15165e-19 $X=1.615 $Y=0.465 $X2=0
+ $Y2=0
cc_266 N_A_208_74#_c_286_n N_VGND_c_760_n 4.64001e-19 $X=2.675 $Y=1.185 $X2=0
+ $Y2=0
cc_267 N_A_208_74#_c_288_n N_VGND_c_760_n 0.0093975f $X=3.105 $Y=1.185 $X2=0
+ $Y2=0
cc_268 N_A_208_74#_c_290_n N_VGND_c_760_n 0.00154624f $X=3.535 $Y=1.185 $X2=0
+ $Y2=0
cc_269 N_A_208_74#_c_284_n N_VGND_c_761_n 0.00383152f $X=2.245 $Y=1.185 $X2=0
+ $Y2=0
cc_270 N_A_208_74#_c_295_n N_VGND_c_761_n 0.0367749f $X=1.615 $Y=0.465 $X2=0
+ $Y2=0
cc_271 N_A_208_74#_c_296_n N_VGND_c_761_n 0.00827872f $X=1.615 $Y=0.465 $X2=0
+ $Y2=0
cc_272 N_A_208_74#_c_286_n N_VGND_c_763_n 0.00383152f $X=2.675 $Y=1.185 $X2=0
+ $Y2=0
cc_273 N_A_208_74#_c_288_n N_VGND_c_763_n 0.00383152f $X=3.105 $Y=1.185 $X2=0
+ $Y2=0
cc_274 N_A_208_74#_c_290_n N_VGND_c_766_n 0.00430908f $X=3.535 $Y=1.185 $X2=0
+ $Y2=0
cc_275 N_A_208_74#_c_284_n N_VGND_c_767_n 0.00762539f $X=2.245 $Y=1.185 $X2=0
+ $Y2=0
cc_276 N_A_208_74#_c_286_n N_VGND_c_767_n 0.0075754f $X=2.675 $Y=1.185 $X2=0
+ $Y2=0
cc_277 N_A_208_74#_c_288_n N_VGND_c_767_n 0.0075754f $X=3.105 $Y=1.185 $X2=0
+ $Y2=0
cc_278 N_A_208_74#_c_290_n N_VGND_c_767_n 0.0081578f $X=3.535 $Y=1.185 $X2=0
+ $Y2=0
cc_279 N_A_208_74#_c_295_n N_VGND_c_767_n 0.0256312f $X=1.615 $Y=0.465 $X2=0
+ $Y2=0
cc_280 N_A_208_74#_c_296_n N_VGND_c_767_n 0.0115893f $X=1.615 $Y=0.465 $X2=0
+ $Y2=0
cc_281 N_A_208_74#_c_284_n N_A_378_74#_c_830_n 0.00122164f $X=2.245 $Y=1.185
+ $X2=0 $Y2=0
cc_282 N_A_208_74#_c_294_n N_A_378_74#_c_830_n 0.00957786f $X=1.615 $Y=1.145
+ $X2=0 $Y2=0
cc_283 N_A_208_74#_c_295_n N_A_378_74#_c_830_n 0.0518232f $X=1.615 $Y=0.465
+ $X2=0 $Y2=0
cc_284 N_A_208_74#_c_296_n N_A_378_74#_c_830_n 0.00601712f $X=1.615 $Y=0.465
+ $X2=0 $Y2=0
cc_285 N_A_208_74#_c_282_n N_A_378_74#_c_831_n 0.00129279f $X=2.17 $Y=1.26 $X2=0
+ $Y2=0
cc_286 N_A_208_74#_c_284_n N_A_378_74#_c_831_n 0.00749872f $X=2.245 $Y=1.185
+ $X2=0 $Y2=0
cc_287 N_A_208_74#_c_285_n N_A_378_74#_c_831_n 0.00643581f $X=2.6 $Y=1.26 $X2=0
+ $Y2=0
cc_288 N_A_208_74#_c_286_n N_A_378_74#_c_831_n 0.00721311f $X=2.675 $Y=1.185
+ $X2=0 $Y2=0
cc_289 N_A_208_74#_c_287_n N_A_378_74#_c_831_n 0.00129486f $X=3.03 $Y=1.26 $X2=0
+ $Y2=0
cc_290 N_A_208_74#_c_291_n N_A_378_74#_c_831_n 0.00365884f $X=2.245 $Y=1.26
+ $X2=0 $Y2=0
cc_291 N_A_208_74#_c_292_n N_A_378_74#_c_831_n 0.00251095f $X=2.675 $Y=1.26
+ $X2=0 $Y2=0
cc_292 N_A_208_74#_c_282_n N_A_378_74#_c_832_n 0.0096098f $X=2.17 $Y=1.26 $X2=0
+ $Y2=0
cc_293 N_A_208_74#_c_294_n N_A_378_74#_c_832_n 0.0137054f $X=1.615 $Y=1.145
+ $X2=0 $Y2=0
cc_294 N_A_208_74#_c_296_n N_A_378_74#_c_832_n 3.76302e-19 $X=1.615 $Y=0.465
+ $X2=0 $Y2=0
cc_295 N_A_208_74#_c_286_n N_A_378_74#_c_833_n 0.00111248f $X=2.675 $Y=1.185
+ $X2=0 $Y2=0
cc_296 N_A_208_74#_c_288_n N_A_378_74#_c_833_n 3.92313e-19 $X=3.105 $Y=1.185
+ $X2=0 $Y2=0
cc_297 N_A_208_74#_c_288_n N_A_378_74#_c_834_n 0.0122885f $X=3.105 $Y=1.185
+ $X2=0 $Y2=0
cc_298 N_A_208_74#_c_289_n N_A_378_74#_c_834_n 0.0024802f $X=3.46 $Y=1.26 $X2=0
+ $Y2=0
cc_299 N_A_208_74#_c_290_n N_A_378_74#_c_834_n 0.0121337f $X=3.535 $Y=1.185
+ $X2=0 $Y2=0
cc_300 N_A_208_74#_c_288_n N_A_378_74#_c_865_n 5.78934e-19 $X=3.105 $Y=1.185
+ $X2=0 $Y2=0
cc_301 N_A_208_74#_c_290_n N_A_378_74#_c_865_n 0.00767715f $X=3.535 $Y=1.185
+ $X2=0 $Y2=0
cc_302 N_A_208_74#_c_290_n N_A_378_74#_c_836_n 0.00322875f $X=3.535 $Y=1.185
+ $X2=0 $Y2=0
cc_303 N_A_208_74#_c_287_n N_A_378_74#_c_839_n 0.0109545f $X=3.03 $Y=1.26 $X2=0
+ $Y2=0
cc_304 N_A_208_74#_c_288_n N_A_378_74#_c_839_n 9.32193e-19 $X=3.105 $Y=1.185
+ $X2=0 $Y2=0
cc_305 N_A_27_368#_c_411_n N_VPWR_M1006_d 0.00602724f $X=1.46 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_306 N_A_27_368#_c_413_n N_VPWR_M1013_d 0.00383849f $X=2.36 $Y=2.145 $X2=0
+ $Y2=0
cc_307 N_A_27_368#_c_415_n N_VPWR_M1013_d 0.00264247f $X=2.445 $Y=2.06 $X2=0
+ $Y2=0
cc_308 N_A_27_368#_c_410_n N_VPWR_c_557_n 0.00901665f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_309 N_A_27_368#_c_411_n N_VPWR_c_557_n 0.0185259f $X=1.46 $Y=2.475 $X2=0
+ $Y2=0
cc_310 N_A_27_368#_c_410_n N_VPWR_c_563_n 0.0124046f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_311 N_A_27_368#_M1000_g N_VPWR_c_564_n 0.00333926f $X=3.91 $Y=2.4 $X2=0 $Y2=0
cc_312 N_A_27_368#_M1002_g N_VPWR_c_564_n 0.00333926f $X=4.36 $Y=2.4 $X2=0 $Y2=0
cc_313 N_A_27_368#_M1003_g N_VPWR_c_564_n 0.00333926f $X=4.81 $Y=2.4 $X2=0 $Y2=0
cc_314 N_A_27_368#_M1010_g N_VPWR_c_564_n 0.00333926f $X=5.26 $Y=2.4 $X2=0 $Y2=0
cc_315 N_A_27_368#_M1000_g N_VPWR_c_556_n 0.00422798f $X=3.91 $Y=2.4 $X2=0 $Y2=0
cc_316 N_A_27_368#_M1002_g N_VPWR_c_556_n 0.00422687f $X=4.36 $Y=2.4 $X2=0 $Y2=0
cc_317 N_A_27_368#_M1003_g N_VPWR_c_556_n 0.00422687f $X=4.81 $Y=2.4 $X2=0 $Y2=0
cc_318 N_A_27_368#_M1010_g N_VPWR_c_556_n 0.00426412f $X=5.26 $Y=2.4 $X2=0 $Y2=0
cc_319 N_A_27_368#_c_410_n N_VPWR_c_556_n 0.0102675f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_320 N_A_27_368#_c_411_n N_VPWR_c_556_n 0.0331756f $X=1.46 $Y=2.475 $X2=0
+ $Y2=0
cc_321 N_A_27_368#_c_413_n N_A_348_368#_M1013_s 0.00859863f $X=2.36 $Y=2.145
+ $X2=-0.19 $Y2=-0.245
cc_322 N_A_27_368#_c_413_n N_A_348_368#_c_635_n 0.028407f $X=2.36 $Y=2.145 $X2=0
+ $Y2=0
cc_323 N_A_27_368#_c_415_n N_A_348_368#_c_626_n 0.00667447f $X=2.445 $Y=2.06
+ $X2=0 $Y2=0
cc_324 N_A_27_368#_c_402_n N_A_348_368#_c_626_n 0.013717f $X=3.82 $Y=1.485 $X2=0
+ $Y2=0
cc_325 N_A_27_368#_c_402_n N_A_348_368#_c_628_n 0.045085f $X=3.82 $Y=1.485 $X2=0
+ $Y2=0
cc_326 N_A_27_368#_c_402_n N_A_348_368#_c_629_n 0.0208665f $X=3.82 $Y=1.485
+ $X2=0 $Y2=0
cc_327 N_A_27_368#_M1000_g N_A_348_368#_c_630_n 0.0139961f $X=3.91 $Y=2.4 $X2=0
+ $Y2=0
cc_328 N_A_27_368#_M1002_g N_A_348_368#_c_630_n 0.0140221f $X=4.36 $Y=2.4 $X2=0
+ $Y2=0
cc_329 N_A_27_368#_M1003_g N_A_348_368#_c_632_n 0.0140221f $X=4.81 $Y=2.4 $X2=0
+ $Y2=0
cc_330 N_A_27_368#_M1010_g N_A_348_368#_c_632_n 0.0148358f $X=5.26 $Y=2.4 $X2=0
+ $Y2=0
cc_331 N_A_27_368#_M1010_g N_A_348_368#_c_633_n 0.00147128f $X=5.26 $Y=2.4 $X2=0
+ $Y2=0
cc_332 N_A_27_368#_c_411_n N_A_348_368#_c_659_n 0.0133002f $X=1.46 $Y=2.475
+ $X2=0 $Y2=0
cc_333 N_A_27_368#_c_413_n N_A_348_368#_c_659_n 0.0126786f $X=2.36 $Y=2.145
+ $X2=0 $Y2=0
cc_334 N_A_27_368#_M1000_g N_Z_c_695_n 0.00267931f $X=3.91 $Y=2.4 $X2=0 $Y2=0
cc_335 N_A_27_368#_M1002_g N_Z_c_695_n 0.00112087f $X=4.36 $Y=2.4 $X2=0 $Y2=0
cc_336 N_A_27_368#_c_399_n N_Z_c_695_n 0.0275254f $X=3.985 $Y=1.485 $X2=0 $Y2=0
cc_337 N_A_27_368#_c_403_n N_Z_c_695_n 0.00225438f $X=5.275 $Y=1.485 $X2=0 $Y2=0
cc_338 N_A_27_368#_M1000_g N_Z_c_699_n 0.0092344f $X=3.91 $Y=2.4 $X2=0 $Y2=0
cc_339 N_A_27_368#_M1002_g N_Z_c_699_n 0.010067f $X=4.36 $Y=2.4 $X2=0 $Y2=0
cc_340 N_A_27_368#_M1003_g N_Z_c_699_n 5.88596e-19 $X=4.81 $Y=2.4 $X2=0 $Y2=0
cc_341 N_A_27_368#_M1005_g N_Z_c_707_n 0.00466922f $X=3.965 $Y=0.74 $X2=0 $Y2=0
cc_342 N_A_27_368#_M1012_g N_Z_c_707_n 0.00587139f $X=4.395 $Y=0.74 $X2=0 $Y2=0
cc_343 N_A_27_368#_M1014_g N_Z_c_707_n 5.63827e-19 $X=4.825 $Y=0.74 $X2=0 $Y2=0
cc_344 N_A_27_368#_M1002_g N_Z_c_696_n 0.012931f $X=4.36 $Y=2.4 $X2=0 $Y2=0
cc_345 N_A_27_368#_M1003_g N_Z_c_696_n 0.0135059f $X=4.81 $Y=2.4 $X2=0 $Y2=0
cc_346 N_A_27_368#_c_505_p N_Z_c_696_n 0.0388286f $X=4.665 $Y=1.485 $X2=0 $Y2=0
cc_347 N_A_27_368#_c_403_n N_Z_c_696_n 0.00209665f $X=5.275 $Y=1.485 $X2=0 $Y2=0
cc_348 N_A_27_368#_M1012_g N_Z_c_691_n 0.00891372f $X=4.395 $Y=0.74 $X2=0 $Y2=0
cc_349 N_A_27_368#_M1014_g N_Z_c_691_n 0.00944863f $X=4.825 $Y=0.74 $X2=0 $Y2=0
cc_350 N_A_27_368#_c_505_p N_Z_c_691_n 0.0356525f $X=4.665 $Y=1.485 $X2=0 $Y2=0
cc_351 N_A_27_368#_c_403_n N_Z_c_691_n 0.00236025f $X=5.275 $Y=1.485 $X2=0 $Y2=0
cc_352 N_A_27_368#_M1005_g N_Z_c_692_n 0.00373071f $X=3.965 $Y=0.74 $X2=0 $Y2=0
cc_353 N_A_27_368#_M1012_g N_Z_c_692_n 0.00235421f $X=4.395 $Y=0.74 $X2=0 $Y2=0
cc_354 N_A_27_368#_c_505_p N_Z_c_692_n 0.0271537f $X=4.665 $Y=1.485 $X2=0 $Y2=0
cc_355 N_A_27_368#_c_403_n N_Z_c_692_n 0.00250921f $X=5.275 $Y=1.485 $X2=0 $Y2=0
cc_356 N_A_27_368#_M1012_g N_Z_c_722_n 5.63827e-19 $X=4.395 $Y=0.74 $X2=0 $Y2=0
cc_357 N_A_27_368#_M1014_g N_Z_c_722_n 0.00640291f $X=4.825 $Y=0.74 $X2=0 $Y2=0
cc_358 N_A_27_368#_M1018_g N_Z_c_722_n 0.0047509f $X=5.275 $Y=0.74 $X2=0 $Y2=0
cc_359 N_A_27_368#_M1003_g N_Z_c_693_n 0.00259091f $X=4.81 $Y=2.4 $X2=0 $Y2=0
cc_360 N_A_27_368#_M1014_g N_Z_c_693_n 0.00261386f $X=4.825 $Y=0.74 $X2=0 $Y2=0
cc_361 N_A_27_368#_M1010_g N_Z_c_693_n 0.00868548f $X=5.26 $Y=2.4 $X2=0 $Y2=0
cc_362 N_A_27_368#_M1018_g N_Z_c_693_n 0.00843462f $X=5.275 $Y=0.74 $X2=0 $Y2=0
cc_363 N_A_27_368#_c_505_p N_Z_c_693_n 0.0214916f $X=4.665 $Y=1.485 $X2=0 $Y2=0
cc_364 N_A_27_368#_c_403_n N_Z_c_693_n 0.0257339f $X=5.275 $Y=1.485 $X2=0 $Y2=0
cc_365 N_A_27_368#_M1014_g N_Z_c_694_n 0.00227685f $X=4.825 $Y=0.74 $X2=0 $Y2=0
cc_366 N_A_27_368#_M1018_g N_Z_c_694_n 0.00363443f $X=5.275 $Y=0.74 $X2=0 $Y2=0
cc_367 N_A_27_368#_c_403_n N_Z_c_694_n 0.0013317f $X=5.275 $Y=1.485 $X2=0 $Y2=0
cc_368 N_A_27_368#_M1003_g Z 0.00153758f $X=4.81 $Y=2.4 $X2=0 $Y2=0
cc_369 N_A_27_368#_M1010_g Z 0.00239532f $X=5.26 $Y=2.4 $X2=0 $Y2=0
cc_370 N_A_27_368#_c_403_n Z 0.00135743f $X=5.275 $Y=1.485 $X2=0 $Y2=0
cc_371 N_A_27_368#_M1002_g Z 5.88486e-19 $X=4.36 $Y=2.4 $X2=0 $Y2=0
cc_372 N_A_27_368#_M1003_g Z 0.010067f $X=4.81 $Y=2.4 $X2=0 $Y2=0
cc_373 N_A_27_368#_M1010_g Z 0.00995107f $X=5.26 $Y=2.4 $X2=0 $Y2=0
cc_374 N_A_27_368#_c_397_n N_VGND_c_758_n 0.024411f $X=0.32 $Y=0.515 $X2=0 $Y2=0
cc_375 N_A_27_368#_c_397_n N_VGND_c_765_n 0.0141895f $X=0.32 $Y=0.515 $X2=0
+ $Y2=0
cc_376 N_A_27_368#_M1005_g N_VGND_c_766_n 0.00278271f $X=3.965 $Y=0.74 $X2=0
+ $Y2=0
cc_377 N_A_27_368#_M1012_g N_VGND_c_766_n 0.00278271f $X=4.395 $Y=0.74 $X2=0
+ $Y2=0
cc_378 N_A_27_368#_M1014_g N_VGND_c_766_n 0.00278271f $X=4.825 $Y=0.74 $X2=0
+ $Y2=0
cc_379 N_A_27_368#_M1018_g N_VGND_c_766_n 0.00278271f $X=5.275 $Y=0.74 $X2=0
+ $Y2=0
cc_380 N_A_27_368#_M1005_g N_VGND_c_767_n 0.00353526f $X=3.965 $Y=0.74 $X2=0
+ $Y2=0
cc_381 N_A_27_368#_M1012_g N_VGND_c_767_n 0.00353428f $X=4.395 $Y=0.74 $X2=0
+ $Y2=0
cc_382 N_A_27_368#_M1014_g N_VGND_c_767_n 0.00353626f $X=4.825 $Y=0.74 $X2=0
+ $Y2=0
cc_383 N_A_27_368#_M1018_g N_VGND_c_767_n 0.00353613f $X=5.275 $Y=0.74 $X2=0
+ $Y2=0
cc_384 N_A_27_368#_c_397_n N_VGND_c_767_n 0.0117448f $X=0.32 $Y=0.515 $X2=0
+ $Y2=0
cc_385 N_A_27_368#_c_398_n N_A_378_74#_c_831_n 0.0137157f $X=2.53 $Y=1.565 $X2=0
+ $Y2=0
cc_386 N_A_27_368#_c_402_n N_A_378_74#_c_831_n 0.0195631f $X=3.82 $Y=1.485 $X2=0
+ $Y2=0
cc_387 N_A_27_368#_M1005_g N_A_378_74#_c_834_n 3.2654e-19 $X=3.965 $Y=0.74 $X2=0
+ $Y2=0
cc_388 N_A_27_368#_c_399_n N_A_378_74#_c_834_n 0.001265f $X=3.985 $Y=1.485 $X2=0
+ $Y2=0
cc_389 N_A_27_368#_c_402_n N_A_378_74#_c_834_n 0.0402638f $X=3.82 $Y=1.485 $X2=0
+ $Y2=0
cc_390 N_A_27_368#_c_403_n N_A_378_74#_c_834_n 4.08598e-19 $X=5.275 $Y=1.485
+ $X2=0 $Y2=0
cc_391 N_A_27_368#_M1005_g N_A_378_74#_c_835_n 0.0122971f $X=3.965 $Y=0.74 $X2=0
+ $Y2=0
cc_392 N_A_27_368#_M1012_g N_A_378_74#_c_835_n 0.0102404f $X=4.395 $Y=0.74 $X2=0
+ $Y2=0
cc_393 N_A_27_368#_M1014_g N_A_378_74#_c_837_n 0.0103604f $X=4.825 $Y=0.74 $X2=0
+ $Y2=0
cc_394 N_A_27_368#_M1018_g N_A_378_74#_c_837_n 0.0139388f $X=5.275 $Y=0.74 $X2=0
+ $Y2=0
cc_395 N_A_27_368#_M1018_g N_A_378_74#_c_838_n 0.00159899f $X=5.275 $Y=0.74
+ $X2=0 $Y2=0
cc_396 N_A_27_368#_c_402_n N_A_378_74#_c_839_n 0.0134254f $X=3.82 $Y=1.485 $X2=0
+ $Y2=0
cc_397 N_VPWR_M1013_d N_A_348_368#_c_635_n 0.00320822f $X=2.2 $Y=1.84 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_558_n N_A_348_368#_c_635_n 0.0165098f $X=2.335 $Y=2.825 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_559_n N_A_348_368#_c_635_n 0.00220374f $X=3.07 $Y=3.33 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_561_n N_A_348_368#_c_635_n 0.00220374f $X=2.17 $Y=3.33 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_556_n N_A_348_368#_c_635_n 0.0100815f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_558_n N_A_348_368#_c_627_n 0.00854446f $X=2.335 $Y=2.825 $X2=0
+ $Y2=0
cc_403 N_VPWR_c_559_n N_A_348_368#_c_627_n 0.00749631f $X=3.07 $Y=3.33 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_560_n N_A_348_368#_c_627_n 0.0135825f $X=3.235 $Y=2.325 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_556_n N_A_348_368#_c_627_n 0.0062048f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_406 N_VPWR_M1017_d N_A_348_368#_c_628_n 0.00165831f $X=3.1 $Y=1.84 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_560_n N_A_348_368#_c_628_n 0.0148589f $X=3.235 $Y=2.325 $X2=0
+ $Y2=0
cc_408 N_VPWR_c_564_n N_A_348_368#_c_630_n 0.0439866f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_409 N_VPWR_c_556_n N_A_348_368#_c_630_n 0.0246722f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_560_n N_A_348_368#_c_631_n 0.0103534f $X=3.235 $Y=2.325 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_564_n N_A_348_368#_c_631_n 0.0178163f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_412 N_VPWR_c_556_n N_A_348_368#_c_631_n 0.00958215f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_413 N_VPWR_c_564_n N_A_348_368#_c_632_n 0.0619083f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_414 N_VPWR_c_556_n N_A_348_368#_c_632_n 0.0343916f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_415 N_VPWR_c_561_n N_A_348_368#_c_659_n 0.00414725f $X=2.17 $Y=3.33 $X2=0
+ $Y2=0
cc_416 N_VPWR_c_556_n N_A_348_368#_c_659_n 0.00547139f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_417 N_VPWR_c_564_n N_A_348_368#_c_634_n 0.016488f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_418 N_VPWR_c_556_n N_A_348_368#_c_634_n 0.00894187f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_419 N_A_348_368#_c_630_n N_Z_M1000_d 0.00165831f $X=4.47 $Y=2.99 $X2=0 $Y2=0
cc_420 N_A_348_368#_c_632_n N_Z_M1003_d 0.00165831f $X=5.4 $Y=2.99 $X2=0 $Y2=0
cc_421 N_A_348_368#_c_629_n N_Z_c_695_n 0.00710059f $X=3.645 $Y=1.99 $X2=0 $Y2=0
cc_422 N_A_348_368#_c_630_n N_Z_c_699_n 0.0159318f $X=4.47 $Y=2.99 $X2=0 $Y2=0
cc_423 N_A_348_368#_M1002_s N_Z_c_696_n 0.00165831f $X=4.45 $Y=1.84 $X2=0 $Y2=0
cc_424 N_A_348_368#_c_688_p N_Z_c_696_n 0.0126919f $X=4.585 $Y=2.325 $X2=0 $Y2=0
cc_425 N_A_348_368#_c_633_n Z 0.00710261f $X=5.485 $Y=1.985 $X2=0 $Y2=0
cc_426 N_A_348_368#_c_632_n Z 0.0162881f $X=5.4 $Y=2.99 $X2=0 $Y2=0
cc_427 N_Z_c_691_n N_A_378_74#_M1012_d 0.00176461f $X=4.875 $Y=1.065 $X2=0 $Y2=0
cc_428 N_Z_c_692_n N_A_378_74#_c_834_n 0.00862188f $X=4.345 $Y=1.065 $X2=0 $Y2=0
cc_429 N_Z_M1005_s N_A_378_74#_c_835_n 0.00176461f $X=4.04 $Y=0.37 $X2=0 $Y2=0
cc_430 N_Z_c_707_n N_A_378_74#_c_835_n 0.0158052f $X=4.18 $Y=0.82 $X2=0 $Y2=0
cc_431 N_Z_c_691_n N_A_378_74#_c_835_n 0.0031794f $X=4.875 $Y=1.065 $X2=0 $Y2=0
cc_432 N_Z_c_691_n N_A_378_74#_c_887_n 0.0132844f $X=4.875 $Y=1.065 $X2=0 $Y2=0
cc_433 N_Z_M1014_s N_A_378_74#_c_837_n 0.00197722f $X=4.9 $Y=0.37 $X2=0 $Y2=0
cc_434 N_Z_c_691_n N_A_378_74#_c_837_n 0.0031794f $X=4.875 $Y=1.065 $X2=0 $Y2=0
cc_435 N_Z_c_722_n N_A_378_74#_c_837_n 0.0160331f $X=5.04 $Y=0.86 $X2=0 $Y2=0
cc_436 N_Z_c_694_n N_A_378_74#_c_838_n 0.00622221f $X=5.04 $Y=1.065 $X2=0 $Y2=0
cc_437 N_VGND_c_759_n N_A_378_74#_c_830_n 0.0229082f $X=2.46 $Y=0.515 $X2=0
+ $Y2=0
cc_438 N_VGND_c_761_n N_A_378_74#_c_830_n 0.00749631f $X=2.295 $Y=0 $X2=0 $Y2=0
cc_439 N_VGND_c_767_n N_A_378_74#_c_830_n 0.0062048f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_440 N_VGND_c_759_n N_A_378_74#_c_831_n 0.0216086f $X=2.46 $Y=0.515 $X2=0
+ $Y2=0
cc_441 N_VGND_c_759_n N_A_378_74#_c_833_n 0.0229082f $X=2.46 $Y=0.515 $X2=0
+ $Y2=0
cc_442 N_VGND_c_760_n N_A_378_74#_c_833_n 0.0164868f $X=3.32 $Y=0.645 $X2=0
+ $Y2=0
cc_443 N_VGND_c_763_n N_A_378_74#_c_833_n 0.00749631f $X=3.155 $Y=0 $X2=0 $Y2=0
cc_444 N_VGND_c_767_n N_A_378_74#_c_833_n 0.0062048f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_445 N_VGND_M1009_d N_A_378_74#_c_834_n 0.00176461f $X=3.18 $Y=0.37 $X2=0
+ $Y2=0
cc_446 N_VGND_c_760_n N_A_378_74#_c_834_n 0.0152916f $X=3.32 $Y=0.645 $X2=0
+ $Y2=0
cc_447 N_VGND_c_766_n N_A_378_74#_c_835_n 0.043517f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_448 N_VGND_c_767_n N_A_378_74#_c_835_n 0.0245693f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_449 N_VGND_c_760_n N_A_378_74#_c_836_n 0.0112234f $X=3.32 $Y=0.645 $X2=0
+ $Y2=0
cc_450 N_VGND_c_766_n N_A_378_74#_c_836_n 0.0178338f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_451 N_VGND_c_767_n N_A_378_74#_c_836_n 0.00960503f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_452 N_VGND_c_766_n N_A_378_74#_c_837_n 0.0627271f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_453 N_VGND_c_767_n N_A_378_74#_c_837_n 0.0350406f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_454 N_VGND_c_766_n N_A_378_74#_c_840_n 0.0120038f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_455 N_VGND_c_767_n N_A_378_74#_c_840_n 0.00657483f $X=5.52 $Y=0 $X2=0 $Y2=0

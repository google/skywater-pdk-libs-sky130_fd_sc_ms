* File: sky130_fd_sc_ms__nor4_1.pxi.spice
* Created: Wed Sep  2 12:16:37 2020
* 
x_PM_SKY130_FD_SC_MS__NOR4_1%A N_A_M1001_g N_A_c_50_n N_A_M1000_g N_A_c_51_n
+ N_A_c_52_n A N_A_c_53_n PM_SKY130_FD_SC_MS__NOR4_1%A
x_PM_SKY130_FD_SC_MS__NOR4_1%B N_B_M1005_g N_B_M1003_g B B B B N_B_c_75_n
+ N_B_c_76_n PM_SKY130_FD_SC_MS__NOR4_1%B
x_PM_SKY130_FD_SC_MS__NOR4_1%C N_C_M1002_g N_C_M1004_g C C N_C_c_114_n
+ N_C_c_115_n PM_SKY130_FD_SC_MS__NOR4_1%C
x_PM_SKY130_FD_SC_MS__NOR4_1%D N_D_M1007_g N_D_M1006_g D N_D_c_151_n N_D_c_152_n
+ PM_SKY130_FD_SC_MS__NOR4_1%D
x_PM_SKY130_FD_SC_MS__NOR4_1%VPWR N_VPWR_M1001_s N_VPWR_c_184_n N_VPWR_c_185_n
+ VPWR N_VPWR_c_186_n N_VPWR_c_183_n PM_SKY130_FD_SC_MS__NOR4_1%VPWR
x_PM_SKY130_FD_SC_MS__NOR4_1%Y N_Y_M1000_d N_Y_M1004_d N_Y_M1006_d N_Y_c_207_n
+ N_Y_c_208_n N_Y_c_209_n N_Y_c_210_n N_Y_c_211_n N_Y_c_212_n N_Y_c_214_n
+ N_Y_c_213_n Y PM_SKY130_FD_SC_MS__NOR4_1%Y
x_PM_SKY130_FD_SC_MS__NOR4_1%VGND N_VGND_M1000_s N_VGND_M1003_d N_VGND_M1007_d
+ N_VGND_c_265_n N_VGND_c_266_n N_VGND_c_267_n N_VGND_c_268_n N_VGND_c_269_n
+ N_VGND_c_270_n N_VGND_c_271_n VGND N_VGND_c_272_n N_VGND_c_273_n
+ PM_SKY130_FD_SC_MS__NOR4_1%VGND
cc_1 VNB N_A_M1001_g 0.00922335f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.4
cc_2 VNB N_A_c_50_n 0.0211013f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.22
cc_3 VNB N_A_c_51_n 0.0412296f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.385
cc_4 VNB N_A_c_52_n 0.0133082f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.385
cc_5 VNB N_A_c_53_n 0.0240277f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.385
cc_6 VNB N_B_M1003_g 0.0267613f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=0.74
cc_7 VNB N_B_c_75_n 0.0251376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B_c_76_n 0.00390329f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.365
cc_9 VNB N_C_M1004_g 0.026814f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=0.74
cc_10 VNB N_C_c_114_n 0.0269862f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.385
cc_11 VNB N_C_c_115_n 0.00167078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_D_M1007_g 0.0264948f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.4
cc_13 VNB N_D_c_151_n 0.0270602f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.385
cc_14 VNB N_D_c_152_n 0.00419952f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.385
cc_15 VNB N_VPWR_c_183_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_Y_c_207_n 0.00215184f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.385
cc_17 VNB N_Y_c_208_n 0.0100809f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.385
cc_18 VNB N_Y_c_209_n 0.00906721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_210_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_211_n 0.0227193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_212_n 0.00789082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_213_n 0.0230393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_265_n 0.016404f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_24 VNB N_VGND_c_266_n 0.0351944f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.385
cc_25 VNB N_VGND_c_267_n 0.00900448f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_26 VNB N_VGND_c_268_n 0.0162041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_269_n 0.0323694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_270_n 0.0168561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_271_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_272_n 0.021877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_273_n 0.193176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VPB N_A_M1001_g 0.029188f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=2.4
cc_33 VPB N_B_M1005_g 0.0224038f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=2.4
cc_34 VPB N_B_c_75_n 0.00558018f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_B_c_76_n 0.00124177f $X=-0.19 $Y=1.66 $X2=0.375 $Y2=1.365
cc_36 VPB N_C_M1002_g 0.0239347f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=2.4
cc_37 VPB N_C_c_114_n 0.00566743f $X=-0.19 $Y=1.66 $X2=0.375 $Y2=1.385
cc_38 VPB N_C_c_115_n 0.00128802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_D_M1006_g 0.0278048f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=0.74
cc_40 VPB N_D_c_151_n 0.00567549f $X=-0.19 $Y=1.66 $X2=0.375 $Y2=1.385
cc_41 VPB N_D_c_152_n 0.00575749f $X=-0.19 $Y=1.66 $X2=0.375 $Y2=1.385
cc_42 VPB N_VPWR_c_184_n 0.0164625f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_185_n 0.0556262f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=0.74
cc_44 VPB N_VPWR_c_186_n 0.0687447f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_183_n 0.0900975f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_Y_c_214_n 0.0138831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_Y_c_213_n 0.0142705f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB Y 0.0405122f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 N_A_M1001_g N_B_M1005_g 0.0446155f $X=0.645 $Y=2.4 $X2=0 $Y2=0
cc_50 N_A_c_50_n N_B_M1003_g 0.0190702f $X=0.66 $Y=1.22 $X2=0 $Y2=0
cc_51 N_A_c_53_n N_B_M1003_g 5.55714e-19 $X=0.375 $Y=1.385 $X2=0 $Y2=0
cc_52 N_A_c_52_n N_B_c_75_n 0.0446155f $X=0.645 $Y=1.385 $X2=0 $Y2=0
cc_53 N_A_c_53_n N_B_c_75_n 5.45707e-19 $X=0.375 $Y=1.385 $X2=0 $Y2=0
cc_54 N_A_c_52_n N_B_c_76_n 0.00655339f $X=0.645 $Y=1.385 $X2=0 $Y2=0
cc_55 N_A_c_53_n N_B_c_76_n 0.00713992f $X=0.375 $Y=1.385 $X2=0 $Y2=0
cc_56 N_A_M1001_g N_VPWR_c_185_n 0.0267629f $X=0.645 $Y=2.4 $X2=0 $Y2=0
cc_57 N_A_c_51_n N_VPWR_c_185_n 0.00683719f $X=0.555 $Y=1.385 $X2=0 $Y2=0
cc_58 N_A_c_53_n N_VPWR_c_185_n 0.0170992f $X=0.375 $Y=1.385 $X2=0 $Y2=0
cc_59 N_A_M1001_g N_VPWR_c_186_n 0.00460063f $X=0.645 $Y=2.4 $X2=0 $Y2=0
cc_60 N_A_M1001_g N_VPWR_c_183_n 0.00908371f $X=0.645 $Y=2.4 $X2=0 $Y2=0
cc_61 N_A_c_50_n N_Y_c_207_n 4.03226e-19 $X=0.66 $Y=1.22 $X2=0 $Y2=0
cc_62 N_A_c_50_n N_Y_c_209_n 0.00221478f $X=0.66 $Y=1.22 $X2=0 $Y2=0
cc_63 N_A_c_50_n N_VGND_c_266_n 0.0131164f $X=0.66 $Y=1.22 $X2=0 $Y2=0
cc_64 N_A_c_51_n N_VGND_c_266_n 0.00230739f $X=0.555 $Y=1.385 $X2=0 $Y2=0
cc_65 N_A_c_53_n N_VGND_c_266_n 0.0282557f $X=0.375 $Y=1.385 $X2=0 $Y2=0
cc_66 N_A_c_50_n N_VGND_c_270_n 0.00383152f $X=0.66 $Y=1.22 $X2=0 $Y2=0
cc_67 N_A_c_50_n N_VGND_c_273_n 0.00757637f $X=0.66 $Y=1.22 $X2=0 $Y2=0
cc_68 N_B_M1005_g N_C_M1002_g 0.0393786f $X=1.065 $Y=2.4 $X2=0 $Y2=0
cc_69 N_B_M1003_g N_C_M1004_g 0.0195058f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_70 N_B_c_75_n N_C_c_114_n 0.0175819f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_71 N_B_c_76_n N_C_c_114_n 0.0225688f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_72 N_B_M1005_g N_C_c_115_n 4.80069e-19 $X=1.065 $Y=2.4 $X2=0 $Y2=0
cc_73 N_B_c_75_n N_C_c_115_n 4.14802e-19 $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_74 N_B_c_76_n N_C_c_115_n 0.0501177f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_75 N_B_M1005_g N_VPWR_c_185_n 0.00379458f $X=1.065 $Y=2.4 $X2=0 $Y2=0
cc_76 N_B_c_76_n N_VPWR_c_185_n 0.0412437f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_77 N_B_M1005_g N_VPWR_c_186_n 0.00365007f $X=1.065 $Y=2.4 $X2=0 $Y2=0
cc_78 N_B_c_76_n N_VPWR_c_186_n 0.00957002f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_79 N_B_M1005_g N_VPWR_c_183_n 0.00444515f $X=1.065 $Y=2.4 $X2=0 $Y2=0
cc_80 N_B_c_76_n N_VPWR_c_183_n 0.010893f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_81 N_B_c_76_n A_231_368# 0.0142235f $X=1.14 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_82 N_B_M1003_g N_Y_c_207_n 0.00968448f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_83 N_B_M1003_g N_Y_c_208_n 0.012155f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_84 N_B_c_75_n N_Y_c_208_n 9.86927e-19 $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_85 N_B_c_76_n N_Y_c_208_n 0.0214362f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_86 N_B_M1003_g N_Y_c_209_n 0.00139157f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_87 N_B_c_75_n N_Y_c_209_n 3.0499e-19 $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_88 N_B_c_76_n N_Y_c_209_n 0.0055933f $X=1.14 $Y=1.515 $X2=0 $Y2=0
cc_89 N_B_M1003_g N_Y_c_210_n 8.51666e-19 $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_90 N_B_M1003_g N_VGND_c_266_n 5.57151e-19 $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_91 N_B_M1003_g N_VGND_c_267_n 0.00543742f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_92 N_B_M1003_g N_VGND_c_270_n 0.00434272f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_93 N_B_M1003_g N_VGND_c_273_n 0.00822072f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_94 N_C_M1004_g N_D_M1007_g 0.0200614f $X=1.76 $Y=0.74 $X2=0 $Y2=0
cc_95 N_C_M1002_g N_D_M1006_g 0.0446788f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_96 N_C_c_115_n N_D_M1006_g 0.00595463f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_97 N_C_c_114_n N_D_c_151_n 0.0173872f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_98 N_C_c_115_n N_D_c_151_n 3.65288e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_99 N_C_M1002_g N_D_c_152_n 2.76671e-19 $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_100 N_C_c_114_n N_D_c_152_n 0.00202953f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_101 N_C_c_115_n N_D_c_152_n 0.0349695f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_102 N_C_M1002_g N_VPWR_c_186_n 0.00553757f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_103 N_C_M1002_g N_VPWR_c_183_n 0.0109203f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_104 N_C_c_115_n A_345_368# 0.00809156f $X=1.71 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_105 N_C_M1004_g N_Y_c_207_n 8.12002e-19 $X=1.76 $Y=0.74 $X2=0 $Y2=0
cc_106 N_C_M1004_g N_Y_c_208_n 0.012155f $X=1.76 $Y=0.74 $X2=0 $Y2=0
cc_107 N_C_c_114_n N_Y_c_208_n 9.6679e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_108 N_C_c_115_n N_Y_c_208_n 0.0205962f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_109 N_C_M1004_g N_Y_c_210_n 0.0111642f $X=1.76 $Y=0.74 $X2=0 $Y2=0
cc_110 N_C_M1004_g N_Y_c_212_n 0.0015571f $X=1.76 $Y=0.74 $X2=0 $Y2=0
cc_111 N_C_c_114_n N_Y_c_212_n 3.08675e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_112 N_C_c_115_n N_Y_c_212_n 0.0055933f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_113 N_C_M1002_g N_Y_c_214_n 0.00392019f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_114 N_C_c_115_n N_Y_c_214_n 0.00847408f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_115 N_C_M1004_g N_VGND_c_267_n 0.00782003f $X=1.76 $Y=0.74 $X2=0 $Y2=0
cc_116 N_C_M1004_g N_VGND_c_272_n 0.00434272f $X=1.76 $Y=0.74 $X2=0 $Y2=0
cc_117 N_C_M1004_g N_VGND_c_273_n 0.00823282f $X=1.76 $Y=0.74 $X2=0 $Y2=0
cc_118 N_D_M1006_g N_VPWR_c_186_n 0.005209f $X=2.205 $Y=2.4 $X2=0 $Y2=0
cc_119 N_D_M1006_g N_VPWR_c_183_n 0.00988707f $X=2.205 $Y=2.4 $X2=0 $Y2=0
cc_120 N_D_M1007_g N_Y_c_210_n 0.01371f $X=2.19 $Y=0.74 $X2=0 $Y2=0
cc_121 N_D_M1007_g N_Y_c_211_n 0.0129505f $X=2.19 $Y=0.74 $X2=0 $Y2=0
cc_122 N_D_c_151_n N_Y_c_211_n 0.00125903f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_123 N_D_c_152_n N_Y_c_211_n 0.0229301f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_124 N_D_M1007_g N_Y_c_212_n 0.0015571f $X=2.19 $Y=0.74 $X2=0 $Y2=0
cc_125 N_D_c_152_n N_Y_c_212_n 0.00829487f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_126 N_D_M1006_g N_Y_c_214_n 0.00499632f $X=2.205 $Y=2.4 $X2=0 $Y2=0
cc_127 N_D_c_151_n N_Y_c_214_n 7.74224e-19 $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_128 N_D_c_152_n N_Y_c_214_n 0.0129929f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_129 N_D_M1007_g N_Y_c_213_n 0.00477786f $X=2.19 $Y=0.74 $X2=0 $Y2=0
cc_130 N_D_M1006_g N_Y_c_213_n 0.00508892f $X=2.205 $Y=2.4 $X2=0 $Y2=0
cc_131 N_D_c_151_n N_Y_c_213_n 0.00739878f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_132 N_D_c_152_n N_Y_c_213_n 0.0332226f $X=2.28 $Y=1.515 $X2=0 $Y2=0
cc_133 N_D_M1006_g Y 0.0175455f $X=2.205 $Y=2.4 $X2=0 $Y2=0
cc_134 N_D_M1007_g N_VGND_c_269_n 0.00722118f $X=2.19 $Y=0.74 $X2=0 $Y2=0
cc_135 N_D_M1007_g N_VGND_c_272_n 0.00434272f $X=2.19 $Y=0.74 $X2=0 $Y2=0
cc_136 N_D_M1007_g N_VGND_c_273_n 0.0082432f $X=2.19 $Y=0.74 $X2=0 $Y2=0
cc_137 N_VPWR_c_186_n Y 0.0230269f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_138 N_VPWR_c_183_n Y 0.0189916f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_139 N_Y_c_208_n N_VGND_M1003_d 0.00764236f $X=1.81 $Y=1.095 $X2=0 $Y2=0
cc_140 N_Y_c_211_n N_VGND_M1007_d 0.0024352f $X=2.615 $Y=1.095 $X2=0 $Y2=0
cc_141 N_Y_c_207_n N_VGND_c_266_n 0.0262671f $X=0.875 $Y=0.515 $X2=0 $Y2=0
cc_142 N_Y_c_207_n N_VGND_c_267_n 0.0185169f $X=0.875 $Y=0.515 $X2=0 $Y2=0
cc_143 N_Y_c_208_n N_VGND_c_267_n 0.0257907f $X=1.81 $Y=1.095 $X2=0 $Y2=0
cc_144 N_Y_c_210_n N_VGND_c_267_n 0.0267123f $X=1.975 $Y=0.515 $X2=0 $Y2=0
cc_145 N_Y_c_210_n N_VGND_c_269_n 0.0191765f $X=1.975 $Y=0.515 $X2=0 $Y2=0
cc_146 N_Y_c_211_n N_VGND_c_269_n 0.0263592f $X=2.615 $Y=1.095 $X2=0 $Y2=0
cc_147 N_Y_c_207_n N_VGND_c_270_n 0.0114405f $X=0.875 $Y=0.515 $X2=0 $Y2=0
cc_148 N_Y_c_210_n N_VGND_c_272_n 0.0144922f $X=1.975 $Y=0.515 $X2=0 $Y2=0
cc_149 N_Y_c_207_n N_VGND_c_273_n 0.00941304f $X=0.875 $Y=0.515 $X2=0 $Y2=0
cc_150 N_Y_c_210_n N_VGND_c_273_n 0.0118826f $X=1.975 $Y=0.515 $X2=0 $Y2=0

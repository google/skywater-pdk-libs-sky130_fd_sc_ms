* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 X a_114_125# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=7.504e+11p pd=5.82e+06u as=2.281e+12p ps=1.709e+07u
M1001 a_27_125# B1 a_300_125# VNB nlowvt w=640000u l=150000u
+  ad=7.904e+11p pd=7.59e+06u as=7.456e+11p ps=7.45e+06u
M1002 VGND a_114_125# X VNB nlowvt w=740000u l=150000u
+  ad=1.2421e+12p pd=1.053e+07u as=4.181e+11p ps=4.09e+06u
M1003 X a_114_125# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_300_125# B2 a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_114_125# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A1 a_300_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_114_125# A2 a_766_387# VPB pshort w=1e+06u l=180000u
+  ad=8.35e+11p pd=7.67e+06u as=6.15e+11p ps=5.23e+06u
M1008 a_300_387# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.85e+11p pd=5.17e+06u as=0p ps=0u
M1009 VGND A2 a_300_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_300_125# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_300_125# B1 a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_125# C1 a_114_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1013 a_766_387# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_114_125# C1 a_27_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_114_125# C1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR C1 a_114_125# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_766_387# A2 a_114_125# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_300_125# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_114_125# B2 a_300_387# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_114_125# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_300_387# B2 a_114_125# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 X a_114_125# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR B1 a_300_387# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR A1 a_766_387# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_27_125# B2 a_300_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_114_125# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_114_125# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

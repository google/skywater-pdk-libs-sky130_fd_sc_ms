* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__mux2i_2 A0 A1 S VGND VNB VPB VPWR Y
M1000 VPWR a_922_72# a_343_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.58023e+12p pd=1.017e+07u as=1.0304e+12p ps=6.32e+06u
M1001 VGND a_922_72# a_115_74# VNB nlowvt w=740000u l=150000u
+  ad=1.10195e+12p pd=8.18e+06u as=5.18e+11p ps=4.36e+06u
M1002 Y A0 a_121_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.1312e+12p pd=8.74e+06u as=6.496e+11p ps=5.64e+06u
M1003 Y A1 a_343_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_922_72# S VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1005 a_337_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=7.8555e+11p pd=5.15e+06u as=8.4255e+11p ps=6.93e+06u
M1006 a_121_368# S VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR S a_121_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_115_74# A0 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_922_72# S VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1010 a_337_74# S VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_121_368# A0 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_343_368# a_922_72# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND S a_337_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_343_368# A1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A1 a_337_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A0 a_115_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_115_74# a_922_72# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__and2b_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__and2b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.450000 0.805000 1.780000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.494400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.975000 1.435000 1.305000 1.620000 ;
        RECT 0.975000 1.620000 2.585000 1.790000 ;
        RECT 2.045000 1.180000 2.585000 1.620000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.026600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.095000 0.350000 3.265000 0.980000 ;
        RECT 3.095000 0.980000 4.675000 1.150000 ;
        RECT 3.095000 1.820000 4.165000 1.990000 ;
        RECT 3.095000 1.990000 3.265000 2.980000 ;
        RECT 3.910000 0.350000 4.160000 0.980000 ;
        RECT 3.995000 1.480000 4.675000 1.650000 ;
        RECT 3.995000 1.650000 4.165000 1.820000 ;
        RECT 3.995000 1.990000 4.165000 2.980000 ;
        RECT 4.445000 1.150000 4.675000 1.480000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.085000  0.350000 0.540000 1.095000 ;
      RECT 0.085000  1.095000 1.845000 1.265000 ;
      RECT 0.085000  1.265000 0.255000 1.950000 ;
      RECT 0.085000  1.950000 0.355000 2.980000 ;
      RECT 0.555000  2.100000 0.885000 3.245000 ;
      RECT 0.710000  0.085000 1.040000 0.925000 ;
      RECT 1.075000  1.960000 2.925000 2.130000 ;
      RECT 1.075000  2.130000 1.405000 2.980000 ;
      RECT 1.210000  0.335000 2.400000 0.585000 ;
      RECT 1.210000  0.585000 1.470000 0.925000 ;
      RECT 1.515000  1.265000 1.845000 1.450000 ;
      RECT 1.605000  2.300000 1.855000 3.245000 ;
      RECT 1.640000  0.755000 2.925000 0.925000 ;
      RECT 2.045000  2.130000 2.375000 2.980000 ;
      RECT 2.565000  2.300000 2.895000 3.245000 ;
      RECT 2.570000  0.085000 2.900000 0.585000 ;
      RECT 2.755000  0.925000 2.925000 1.320000 ;
      RECT 2.755000  1.320000 3.825000 1.650000 ;
      RECT 2.755000  1.650000 2.925000 1.960000 ;
      RECT 3.445000  0.085000 3.695000 0.810000 ;
      RECT 3.465000  2.160000 3.795000 3.245000 ;
      RECT 4.340000  0.085000 4.670000 0.810000 ;
      RECT 4.365000  1.820000 4.695000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_ms__and2b_4

* File: sky130_fd_sc_ms__o31a_2.pex.spice
* Created: Fri Aug 28 18:02:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O31A_2%A_55_264# 1 2 9 13 15 19 23 25 27 28 29 34 36
+ 41 45 46 49 54
c107 34 0 5.17841e-20 $X=3.56 $Y=0.96
r108 54 55 32.4387 $w=3.65e-07 $l=7.5e-08 $layer=POLY_cond $X=0.457 $Y=1.395
+ $X2=0.457 $Y2=1.32
r109 47 49 1.43009 $w=4.58e-07 $l=5.5e-08 $layer=LI1_cond $X=2.995 $Y=2.405
+ $X2=2.995 $Y2=2.46
r110 45 47 7.80051 $w=4.58e-07 $l=3e-07 $layer=LI1_cond $X=2.995 $Y=2.105
+ $X2=2.995 $Y2=2.405
r111 45 46 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.995 $Y=2.105
+ $X2=2.995 $Y2=1.94
r112 42 57 40.9207 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.457 $Y=1.485
+ $X2=0.457 $Y2=1.65
r113 42 54 14.2284 $w=3.65e-07 $l=9e-08 $layer=POLY_cond $X=0.457 $Y=1.485
+ $X2=0.457 $Y2=1.395
r114 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.44
+ $Y=1.485 $X2=0.44 $Y2=1.485
r115 38 41 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.31 $Y=1.485
+ $X2=0.44 $Y2=1.485
r116 34 50 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.56 $Y=1.045
+ $X2=3.14 $Y2=1.045
r117 34 36 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.56 $Y=0.96
+ $X2=3.56 $Y2=0.515
r118 32 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=1.13
+ $X2=3.14 $Y2=1.045
r119 32 46 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=3.14 $Y=1.13
+ $X2=3.14 $Y2=1.94
r120 28 47 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=2.765 $Y=2.405
+ $X2=2.995 $Y2=2.405
r121 28 29 154.62 $w=1.68e-07 $l=2.37e-06 $layer=LI1_cond $X=2.765 $Y=2.405
+ $X2=0.395 $Y2=2.405
r122 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.31 $Y=2.32
+ $X2=0.395 $Y2=2.405
r123 26 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.31 $Y=1.65
+ $X2=0.31 $Y2=1.485
r124 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.31 $Y=1.65
+ $X2=0.31 $Y2=2.32
r125 21 25 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=1.01 $Y=1.47
+ $X2=1.01 $Y2=1.395
r126 21 23 361.5 $w=1.8e-07 $l=9.3e-07 $layer=POLY_cond $X=1.01 $Y=1.47 $X2=1.01
+ $Y2=2.4
r127 17 25 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=0.995 $Y=1.32
+ $X2=1.01 $Y2=1.395
r128 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.995 $Y=1.32
+ $X2=0.995 $Y2=0.74
r129 16 54 23.6381 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=0.64 $Y=1.395
+ $X2=0.457 $Y2=1.395
r130 15 25 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.92 $Y=1.395
+ $X2=1.01 $Y2=1.395
r131 15 16 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.92 $Y=1.395
+ $X2=0.64 $Y2=1.395
r132 13 55 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.565 $Y=0.74
+ $X2=0.565 $Y2=1.32
r133 9 57 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=0.505 $Y=2.4
+ $X2=0.505 $Y2=1.65
r134 2 49 300 $w=1.7e-07 $l=5.89491e-07 $layer=licon1_PDIFF $count=2 $X=2.735
+ $Y=1.96 $X2=2.93 $Y2=2.46
r135 2 45 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=2.735
+ $Y=1.96 $X2=2.93 $Y2=2.105
r136 1 36 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=3.35
+ $Y=0.37 $X2=3.56 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_2%A1 3 7 9 10 14 15
c40 7 0 1.1955e-19 $X=1.655 $Y=2.46
r41 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.58 $Y=1.515
+ $X2=1.58 $Y2=1.68
r42 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.58 $Y=1.515
+ $X2=1.58 $Y2=1.35
r43 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.58
+ $Y=1.515 $X2=1.58 $Y2=1.515
r44 9 10 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.605 $Y=1.665
+ $X2=1.605 $Y2=2.035
r45 9 15 4.54912 $w=3.78e-07 $l=1.5e-07 $layer=LI1_cond $X=1.605 $Y=1.665
+ $X2=1.605 $Y2=1.515
r46 7 17 303.194 $w=1.8e-07 $l=7.8e-07 $layer=POLY_cond $X=1.655 $Y=2.46
+ $X2=1.655 $Y2=1.68
r47 3 16 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.565 $Y=0.74
+ $X2=1.565 $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_2%A2 3 7 9 10 14
c36 9 0 9.66157e-20 $X=2.16 $Y=1.665
r37 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.635
+ $X2=2.15 $Y2=1.8
r38 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.635
+ $X2=2.15 $Y2=1.47
r39 9 10 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=2.15 $Y=1.635 $X2=2.15
+ $Y2=2.035
r40 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.15
+ $Y=1.635 $X2=2.15 $Y2=1.635
r41 7 17 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.075 $Y=2.46
+ $X2=2.075 $Y2=1.8
r42 3 16 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.06 $Y=0.74 $X2=2.06
+ $Y2=1.47
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_2%A3 3 6 8 11 13
c38 11 0 9.66157e-20 $X=2.72 $Y=1.385
c39 8 0 1.98306e-19 $X=2.64 $Y=1.295
r40 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.72 $Y=1.385
+ $X2=2.72 $Y2=1.55
r41 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.72 $Y=1.385
+ $X2=2.72 $Y2=1.22
r42 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.72
+ $Y=1.385 $X2=2.72 $Y2=1.385
r43 8 12 2.88111 $w=3.58e-07 $l=9e-08 $layer=LI1_cond $X=2.705 $Y=1.295
+ $X2=2.705 $Y2=1.385
r44 6 14 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=2.645 $Y=2.46
+ $X2=2.645 $Y2=1.55
r45 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.63 $Y=0.74 $X2=2.63
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_2%B1 1 3 8 10 11 17 18
c32 8 0 1.98306e-19 $X=3.275 $Y=0.74
c33 1 0 5.17841e-20 $X=3.185 $Y=1.88
r34 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.56
+ $Y=1.465 $X2=3.56 $Y2=1.465
r35 15 17 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=3.275 $Y=1.465
+ $X2=3.56 $Y2=1.465
r36 13 15 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.2 $Y=1.465
+ $X2=3.275 $Y2=1.465
r37 11 18 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.56 $Y=1.665 $X2=3.56
+ $Y2=1.465
r38 6 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.275 $Y=1.3
+ $X2=3.275 $Y2=1.465
r39 6 8 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.275 $Y=1.3 $X2=3.275
+ $Y2=0.74
r40 4 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.2 $Y=1.63 $X2=3.2
+ $Y2=1.465
r41 4 10 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=3.2 $Y=1.63 $X2=3.2
+ $Y2=1.79
r42 1 10 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.185 $Y=1.88 $X2=3.185
+ $Y2=1.79
r43 1 3 155.311 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=3.185 $Y=1.88
+ $X2=3.185 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_2%VPWR 1 2 3 10 12 16 18 20 24 26 31 43 47
r43 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r44 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r45 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r46 38 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r47 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 35 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r49 34 37 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r50 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 32 43 11.6267 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=1.595 $Y=3.33
+ $X2=1.332 $Y2=3.33
r52 32 34 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.595 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 31 46 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=3.395 $Y=3.33
+ $X2=3.617 $Y2=3.33
r54 31 37 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.395 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 30 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 30 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r57 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 27 40 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r59 27 29 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 26 43 11.6267 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=1.07 $Y=3.33
+ $X2=1.332 $Y2=3.33
r61 26 29 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.07 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 24 38 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=3.12 $Y2=3.33
r63 24 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r64 20 23 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=3.56 $Y=2.115 $X2=3.56
+ $Y2=2.815
r65 18 46 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.56 $Y=3.245
+ $X2=3.617 $Y2=3.33
r66 18 23 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.56 $Y=3.245
+ $X2=3.56 $Y2=2.815
r67 14 43 2.19831 $w=5.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.332 $Y=3.245
+ $X2=1.332 $Y2=3.33
r68 14 16 9.79645 $w=5.23e-07 $l=4.3e-07 $layer=LI1_cond $X=1.332 $Y=3.245
+ $X2=1.332 $Y2=2.815
r69 10 40 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r70 10 12 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.78
r71 3 23 400 $w=1.7e-07 $l=9.87269e-07 $layer=licon1_PDIFF $count=1 $X=3.275
+ $Y=1.96 $X2=3.56 $Y2=2.815
r72 3 20 400 $w=1.7e-07 $l=3.54119e-07 $layer=licon1_PDIFF $count=1 $X=3.275
+ $Y=1.96 $X2=3.56 $Y2=2.115
r73 2 16 600 $w=1.7e-07 $l=1.08392e-06 $layer=licon1_PDIFF $count=1 $X=1.1
+ $Y=1.84 $X2=1.33 $Y2=2.815
r74 1 12 600 $w=1.7e-07 $l=1.0099e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_2%X 1 2 9 12 13 14 20
c36 12 0 1.1955e-19 $X=0.86 $Y=1.82
r37 14 20 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=0.72 $Y=1.985
+ $X2=0.86 $Y2=1.985
r38 12 20 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.86 $Y=1.82
+ $X2=0.86 $Y2=1.985
r39 12 13 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.86 $Y=1.82 $X2=0.86
+ $Y2=1.13
r40 7 13 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.78 $Y=0.965
+ $X2=0.78 $Y2=1.13
r41 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.78 $Y=0.965 $X2=0.78
+ $Y2=0.515
r42 2 14 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.755 $Y2=1.985
r43 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.64
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_2%VGND 1 2 3 10 12 16 18 22 24 26 36 37 43 46
r48 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r49 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r50 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r51 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r52 34 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r53 34 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r54 33 36 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r55 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r56 31 46 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=2.51 $Y=0 $X2=2.312
+ $Y2=0
r57 31 33 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.51 $Y=0 $X2=2.64
+ $Y2=0
r58 30 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r59 30 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r60 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r61 27 40 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r62 27 29 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r63 26 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.28
+ $Y2=0
r64 26 29 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=0.72
+ $Y2=0
r65 24 47 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r66 24 44 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r67 20 46 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.312 $Y=0.085
+ $X2=2.312 $Y2=0
r68 20 22 12.5456 $w=3.93e-07 $l=4.3e-07 $layer=LI1_cond $X=2.312 $Y=0.085
+ $X2=2.312 $Y2=0.515
r69 19 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.28
+ $Y2=0
r70 18 46 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=2.312
+ $Y2=0
r71 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=1.445
+ $Y2=0
r72 14 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0
r73 14 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0.515
r74 10 40 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r75 10 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.515
r76 3 22 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=2.135
+ $Y=0.37 $X2=2.31 $Y2=0.515
r77 2 16 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.28 $Y2=0.515
r78 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_2%A_328_74# 1 2 7 9 11 16
r30 12 14 4.5891 $w=1.7e-07 $l=2.07123e-07 $layer=LI1_cond $X=1.945 $Y=0.855
+ $X2=1.78 $Y2=0.95
r31 11 16 6.57143 $w=4.27e-07 $l=3.69519e-07 $layer=LI1_cond $X=2.68 $Y=0.855
+ $X2=2.952 $Y2=0.625
r32 11 12 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.68 $Y=0.855
+ $X2=1.945 $Y2=0.855
r33 7 14 3.17707 $w=3.3e-07 $l=1.8e-07 $layer=LI1_cond $X=1.78 $Y=0.77 $X2=1.78
+ $Y2=0.95
r34 7 9 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.78 $Y=0.77 $X2=1.78
+ $Y2=0.515
r35 2 16 182 $w=1.7e-07 $l=3.57071e-07 $layer=licon1_NDIFF $count=1 $X=2.705
+ $Y=0.37 $X2=2.95 $Y2=0.625
r36 1 14 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.64
+ $Y=0.37 $X2=1.78 $Y2=0.965
r37 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.64
+ $Y=0.37 $X2=1.78 $Y2=0.515
.ends


* File: sky130_fd_sc_ms__mux2i_2.pxi.spice
* Created: Wed Sep  2 12:12:06 2020
* 
x_PM_SKY130_FD_SC_MS__MUX2I_2%A0 N_A0_c_92_n N_A0_M1008_g N_A0_M1002_g
+ N_A0_M1011_g N_A0_c_95_n N_A0_M1016_g A0 A0 N_A0_c_97_n
+ PM_SKY130_FD_SC_MS__MUX2I_2%A0
x_PM_SKY130_FD_SC_MS__MUX2I_2%A1 N_A1_M1005_g N_A1_M1003_g N_A1_c_145_n
+ N_A1_M1014_g N_A1_M1015_g A1 A1 A1 A1 N_A1_c_148_n N_A1_c_149_n
+ PM_SKY130_FD_SC_MS__MUX2I_2%A1
x_PM_SKY130_FD_SC_MS__MUX2I_2%S N_S_c_207_n N_S_M1010_g N_S_M1006_g N_S_M1007_g
+ N_S_c_208_n N_S_M1013_g N_S_M1004_g N_S_M1009_g N_S_c_227_p N_S_c_209_n
+ N_S_c_210_n S S S N_S_c_211_n N_S_c_212_n N_S_c_213_n N_S_c_214_n
+ PM_SKY130_FD_SC_MS__MUX2I_2%S
x_PM_SKY130_FD_SC_MS__MUX2I_2%A_922_72# N_A_922_72#_M1009_d N_A_922_72#_M1004_d
+ N_A_922_72#_c_303_n N_A_922_72#_M1001_g N_A_922_72#_M1000_g
+ N_A_922_72#_M1012_g N_A_922_72#_c_304_n N_A_922_72#_M1017_g
+ N_A_922_72#_c_305_n N_A_922_72#_c_330_n N_A_922_72#_c_362_p
+ N_A_922_72#_c_306_n N_A_922_72#_c_307_n N_A_922_72#_c_313_n
+ N_A_922_72#_c_308_n N_A_922_72#_c_309_n PM_SKY130_FD_SC_MS__MUX2I_2%A_922_72#
x_PM_SKY130_FD_SC_MS__MUX2I_2%Y N_Y_M1008_s N_Y_M1016_s N_Y_M1015_s N_Y_M1002_d
+ N_Y_M1011_d N_Y_M1014_d N_Y_c_380_n N_Y_c_386_n N_Y_c_381_n N_Y_c_382_n
+ N_Y_c_383_n N_Y_c_384_n Y Y Y N_Y_c_388_n N_Y_c_385_n Y
+ PM_SKY130_FD_SC_MS__MUX2I_2%Y
x_PM_SKY130_FD_SC_MS__MUX2I_2%A_121_368# N_A_121_368#_M1002_s
+ N_A_121_368#_M1006_d N_A_121_368#_c_459_n N_A_121_368#_c_447_n
+ N_A_121_368#_c_448_n N_A_121_368#_c_449_n
+ PM_SKY130_FD_SC_MS__MUX2I_2%A_121_368#
x_PM_SKY130_FD_SC_MS__MUX2I_2%A_343_368# N_A_343_368#_M1003_s
+ N_A_343_368#_M1000_s N_A_343_368#_c_483_n N_A_343_368#_c_490_n
+ N_A_343_368#_c_485_n N_A_343_368#_c_488_n N_A_343_368#_c_507_n
+ N_A_343_368#_c_484_n PM_SKY130_FD_SC_MS__MUX2I_2%A_343_368#
x_PM_SKY130_FD_SC_MS__MUX2I_2%VPWR N_VPWR_M1006_s N_VPWR_M1007_s N_VPWR_M1012_d
+ N_VPWR_c_527_n N_VPWR_c_528_n N_VPWR_c_529_n N_VPWR_c_530_n N_VPWR_c_531_n
+ N_VPWR_c_532_n VPWR N_VPWR_c_533_n N_VPWR_c_534_n N_VPWR_c_526_n
+ N_VPWR_c_536_n PM_SKY130_FD_SC_MS__MUX2I_2%VPWR
x_PM_SKY130_FD_SC_MS__MUX2I_2%A_115_74# N_A_115_74#_M1008_d N_A_115_74#_M1001_s
+ N_A_115_74#_c_594_n N_A_115_74#_c_592_n N_A_115_74#_c_596_n
+ N_A_115_74#_c_606_n N_A_115_74#_c_593_n N_A_115_74#_c_610_n
+ N_A_115_74#_c_611_n PM_SKY130_FD_SC_MS__MUX2I_2%A_115_74#
x_PM_SKY130_FD_SC_MS__MUX2I_2%A_337_74# N_A_337_74#_M1005_d N_A_337_74#_M1010_d
+ N_A_337_74#_c_655_n N_A_337_74#_c_656_n N_A_337_74#_c_657_n
+ PM_SKY130_FD_SC_MS__MUX2I_2%A_337_74#
x_PM_SKY130_FD_SC_MS__MUX2I_2%VGND N_VGND_M1010_s N_VGND_M1013_s N_VGND_M1017_d
+ N_VGND_c_685_n N_VGND_c_686_n N_VGND_c_687_n N_VGND_c_688_n N_VGND_c_689_n
+ N_VGND_c_690_n N_VGND_c_691_n VGND N_VGND_c_692_n N_VGND_c_693_n
+ N_VGND_c_694_n N_VGND_c_695_n PM_SKY130_FD_SC_MS__MUX2I_2%VGND
cc_1 VNB N_A0_c_92_n 0.019784f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.22
cc_2 VNB N_A0_M1002_g 0.00659492f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.4
cc_3 VNB N_A0_M1011_g 0.00680068f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_4 VNB N_A0_c_95_n 0.0181514f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=1.22
cc_5 VNB A0 0.0186724f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_6 VNB N_A0_c_97_n 0.0481091f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=1.385
cc_7 VNB N_A1_M1005_g 0.0294747f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.74
cc_8 VNB N_A1_c_145_n 0.0337283f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_9 VNB N_A1_M1015_g 0.03266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB A1 0.0149308f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.385
cc_11 VNB N_A1_c_148_n 0.0122419f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.365
cc_12 VNB N_A1_c_149_n 0.0169344f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.365
cc_13 VNB N_S_c_207_n 0.0206654f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.22
cc_14 VNB N_S_c_208_n 0.019018f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=1.22
cc_15 VNB N_S_c_209_n 0.0017739f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=1.385
cc_16 VNB N_S_c_210_n 0.0298867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_S_c_211_n 0.0440126f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_S_c_212_n 0.0227992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_S_c_213_n 0.00534662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_S_c_214_n 0.00471257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_922_72#_c_303_n 0.0185099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_922_72#_c_304_n 0.0176316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_922_72#_c_305_n 0.00113063f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.385
cc_24 VNB N_A_922_72#_c_306_n 0.0212892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_922_72#_c_307_n 0.00720662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_922_72#_c_308_n 0.0223385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_922_72#_c_309_n 0.038183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_380_n 0.0159312f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.385
cc_29 VNB N_Y_c_381_n 0.0108475f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.365
cc_30 VNB N_Y_c_382_n 0.0101912f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.365
cc_31 VNB N_Y_c_383_n 0.00723062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_384_n 0.00724446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_385_n 0.0299842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_526_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_115_74#_c_592_n 0.0059686f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_36 VNB N_A_115_74#_c_593_n 0.00384221f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.385
cc_37 VNB N_A_337_74#_c_655_n 0.00480724f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_38 VNB N_A_337_74#_c_656_n 0.00254729f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_39 VNB N_A_337_74#_c_657_n 0.023826f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_40 VNB N_VGND_c_685_n 0.0135172f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=1.22
cc_41 VNB N_VGND_c_686_n 0.0169046f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_42 VNB N_VGND_c_687_n 0.023772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_688_n 0.0740423f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.385
cc_44 VNB N_VGND_c_689_n 0.00631593f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.385
cc_45 VNB N_VGND_c_690_n 0.0203649f $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=1.385
cc_46 VNB N_VGND_c_691_n 0.00660419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_692_n 0.0202039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_693_n 0.0202442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_694_n 0.350853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_695_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VPB N_A0_M1002_g 0.0289963f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_52 VPB N_A0_M1011_g 0.0253584f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_53 VPB N_A1_M1003_g 0.0261349f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A1_c_145_n 0.0148122f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_55 VPB N_A1_M1014_g 0.0293186f $X=-0.19 $Y=1.66 $X2=1.02 $Y2=0.74
cc_56 VPB A1 0.0182834f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.385
cc_57 VPB N_A1_c_148_n 7.55233e-19 $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.365
cc_58 VPB N_A1_c_149_n 9.52843e-19 $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.365
cc_59 VPB N_S_M1006_g 0.0234017f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=2.4
cc_60 VPB N_S_M1007_g 0.0220348f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_61 VPB N_S_M1004_g 0.025742f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_S_c_209_n 0.00174584f $X=-0.19 $Y=1.66 $X2=1.02 $Y2=1.385
cc_63 VPB N_S_c_210_n 0.00626128f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_S_c_211_n 0.00606885f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_S_c_213_n 0.0100906f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_S_c_214_n 3.66167e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_922_72#_M1000_g 0.0231187f $X=-0.19 $Y=1.66 $X2=1.02 $Y2=1.22
cc_68 VPB N_A_922_72#_M1012_g 0.0234954f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.21
cc_69 VPB N_A_922_72#_c_305_n 5.53756e-19 $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.385
cc_70 VPB N_A_922_72#_c_313_n 0.0300891f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_922_72#_c_308_n 0.0208264f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_922_72#_c_309_n 0.00346598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_Y_c_386_n 0.00245455f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB Y 0.0371002f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_Y_c_388_n 0.0186517f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_Y_c_385_n 0.00776535f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_121_368#_c_447_n 0.00275735f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.21
cc_78 VPB N_A_121_368#_c_448_n 0.00556798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_121_368#_c_449_n 0.00616889f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_343_368#_c_483_n 0.00711562f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_81 VPB N_A_343_368#_c_484_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.385
cc_82 VPB N_VPWR_c_527_n 0.00782802f $X=-0.19 $Y=1.66 $X2=1.02 $Y2=1.22
cc_83 VPB N_VPWR_c_528_n 0.0141893f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.21
cc_84 VPB N_VPWR_c_529_n 0.0202609f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.385
cc_85 VPB N_VPWR_c_530_n 0.00660357f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.385
cc_86 VPB N_VPWR_c_531_n 0.018916f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.385
cc_87 VPB N_VPWR_c_532_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.385
cc_88 VPB N_VPWR_c_533_n 0.0857144f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.365
cc_89 VPB N_VPWR_c_534_n 0.0206493f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_526_n 0.0925982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_536_n 0.0160597f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 N_A0_c_95_n N_A1_M1005_g 0.0258129f $X=1.02 $Y=1.22 $X2=0 $Y2=0
cc_93 A0 N_A1_M1005_g 0.0056955f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_94 N_A0_M1011_g N_A1_M1003_g 0.0258129f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_95 A0 A1 0.00865884f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_96 N_A0_c_97_n A1 0.00138054f $X=1.02 $Y=1.385 $X2=0 $Y2=0
cc_97 A0 N_A1_c_148_n 5.47694e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_98 N_A0_c_97_n N_A1_c_148_n 0.0258129f $X=1.02 $Y=1.385 $X2=0 $Y2=0
cc_99 N_A0_c_92_n N_Y_c_380_n 0.00624207f $X=0.5 $Y=1.22 $X2=0 $Y2=0
cc_100 N_A0_c_95_n N_Y_c_380_n 9.06811e-19 $X=1.02 $Y=1.22 $X2=0 $Y2=0
cc_101 N_A0_M1002_g N_Y_c_386_n 0.0157991f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_102 N_A0_M1011_g N_Y_c_386_n 0.0141495f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_103 A0 N_Y_c_386_n 0.0306472f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_104 N_A0_c_97_n N_Y_c_386_n 0.002473f $X=1.02 $Y=1.385 $X2=0 $Y2=0
cc_105 N_A0_c_92_n N_Y_c_381_n 0.0105638f $X=0.5 $Y=1.22 $X2=0 $Y2=0
cc_106 N_A0_c_95_n N_Y_c_381_n 0.0103939f $X=1.02 $Y=1.22 $X2=0 $Y2=0
cc_107 N_A0_c_92_n N_Y_c_382_n 0.00287994f $X=0.5 $Y=1.22 $X2=0 $Y2=0
cc_108 N_A0_c_92_n N_Y_c_383_n 0.00228454f $X=0.5 $Y=1.22 $X2=0 $Y2=0
cc_109 A0 N_Y_c_383_n 0.00188965f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_110 N_A0_M1002_g Y 0.0121649f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_111 N_A0_M1002_g N_Y_c_388_n 0.0039561f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_112 N_A0_M1011_g N_Y_c_388_n 0.00119358f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_113 A0 N_Y_c_388_n 0.00105488f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_114 N_A0_c_92_n N_Y_c_385_n 0.00586267f $X=0.5 $Y=1.22 $X2=0 $Y2=0
cc_115 A0 N_Y_c_385_n 0.0293669f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_116 N_A0_c_97_n N_Y_c_385_n 0.00771343f $X=1.02 $Y=1.385 $X2=0 $Y2=0
cc_117 N_A0_M1002_g N_A_121_368#_c_447_n 4.62771e-19 $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A0_M1011_g N_A_121_368#_c_447_n 0.0133304f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A0_M1011_g N_A_121_368#_c_448_n 0.0134995f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A0_M1011_g N_A_343_368#_c_485_n 0.00144509f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_121 N_A0_M1002_g N_VPWR_c_533_n 0.0053223f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_122 N_A0_M1011_g N_VPWR_c_533_n 0.005209f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_123 N_A0_M1002_g N_VPWR_c_526_n 0.0102422f $X=0.515 $Y=2.4 $X2=0 $Y2=0
cc_124 N_A0_M1011_g N_VPWR_c_526_n 0.00985263f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_125 N_A0_c_95_n N_A_115_74#_c_594_n 0.00969651f $X=1.02 $Y=1.22 $X2=0 $Y2=0
cc_126 A0 N_A_115_74#_c_594_n 0.0124833f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_127 N_A0_c_92_n N_A_115_74#_c_596_n 0.00363306f $X=0.5 $Y=1.22 $X2=0 $Y2=0
cc_128 N_A0_c_95_n N_A_115_74#_c_596_n 0.00695442f $X=1.02 $Y=1.22 $X2=0 $Y2=0
cc_129 A0 N_A_115_74#_c_596_n 0.025093f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_130 N_A0_c_97_n N_A_115_74#_c_596_n 0.00128387f $X=1.02 $Y=1.385 $X2=0 $Y2=0
cc_131 A0 N_A_337_74#_c_655_n 0.00368238f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_132 N_A0_c_92_n N_VGND_c_688_n 0.00278247f $X=0.5 $Y=1.22 $X2=0 $Y2=0
cc_133 N_A0_c_95_n N_VGND_c_688_n 0.00278271f $X=1.02 $Y=1.22 $X2=0 $Y2=0
cc_134 N_A0_c_92_n N_VGND_c_694_n 0.00357932f $X=0.5 $Y=1.22 $X2=0 $Y2=0
cc_135 N_A0_c_95_n N_VGND_c_694_n 0.00354744f $X=1.02 $Y=1.22 $X2=0 $Y2=0
cc_136 A1 N_S_c_211_n 0.00235925f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_137 A1 N_S_c_213_n 0.024491f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_138 N_A1_M1003_g N_Y_c_386_n 0.0139701f $X=1.625 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A1_c_145_n N_Y_c_386_n 0.00259259f $X=2.365 $Y=1.515 $X2=0 $Y2=0
cc_140 N_A1_M1014_g N_Y_c_386_n 0.0111838f $X=2.455 $Y=2.4 $X2=0 $Y2=0
cc_141 A1 N_Y_c_386_n 0.093904f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_142 N_A1_M1005_g N_Y_c_381_n 0.0114875f $X=1.61 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A1_M1015_g N_Y_c_381_n 0.0119796f $X=2.47 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A1_M1015_g N_Y_c_384_n 0.00185541f $X=2.47 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A1_M1003_g N_A_121_368#_c_447_n 0.00232723f $X=1.625 $Y=2.4 $X2=0 $Y2=0
cc_146 N_A1_M1003_g N_A_121_368#_c_448_n 0.0183193f $X=1.625 $Y=2.4 $X2=0 $Y2=0
cc_147 N_A1_M1014_g N_A_121_368#_c_448_n 0.0152137f $X=2.455 $Y=2.4 $X2=0 $Y2=0
cc_148 A1 N_A_121_368#_c_448_n 0.006306f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_149 N_A1_M1014_g N_A_121_368#_c_449_n 0.00378916f $X=2.455 $Y=2.4 $X2=0 $Y2=0
cc_150 A1 N_A_121_368#_c_449_n 0.0146554f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_151 N_A1_M1014_g N_A_343_368#_c_483_n 0.0111379f $X=2.455 $Y=2.4 $X2=0 $Y2=0
cc_152 N_A1_M1003_g N_A_343_368#_c_485_n 0.00842594f $X=1.625 $Y=2.4 $X2=0 $Y2=0
cc_153 N_A1_M1014_g N_A_343_368#_c_488_n 0.00884202f $X=2.455 $Y=2.4 $X2=0 $Y2=0
cc_154 N_A1_M1003_g N_VPWR_c_533_n 0.00520465f $X=1.625 $Y=2.4 $X2=0 $Y2=0
cc_155 N_A1_M1014_g N_VPWR_c_533_n 0.00373961f $X=2.455 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A1_M1003_g N_VPWR_c_526_n 0.00984566f $X=1.625 $Y=2.4 $X2=0 $Y2=0
cc_157 N_A1_M1014_g N_VPWR_c_526_n 0.00469483f $X=2.455 $Y=2.4 $X2=0 $Y2=0
cc_158 N_A1_M1014_g N_VPWR_c_536_n 0.00326111f $X=2.455 $Y=2.4 $X2=0 $Y2=0
cc_159 N_A1_M1005_g N_A_115_74#_c_594_n 0.0147737f $X=1.61 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A1_c_145_n N_A_115_74#_c_594_n 6.3897e-19 $X=2.365 $Y=1.515 $X2=0 $Y2=0
cc_161 N_A1_M1015_g N_A_115_74#_c_594_n 3.85527e-19 $X=2.47 $Y=0.74 $X2=0 $Y2=0
cc_162 A1 N_A_115_74#_c_594_n 0.00413062f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_163 N_A1_M1015_g N_A_115_74#_c_592_n 0.010944f $X=2.47 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A1_M1005_g N_A_115_74#_c_596_n 0.00118817f $X=1.61 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A1_M1005_g N_A_115_74#_c_606_n 0.00251864f $X=1.61 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A1_M1015_g N_A_115_74#_c_606_n 0.0102998f $X=2.47 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A1_M1015_g N_A_115_74#_c_593_n 0.00176656f $X=2.47 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A1_M1005_g N_A_337_74#_c_655_n 0.00507838f $X=1.61 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A1_c_145_n N_A_337_74#_c_655_n 0.00750284f $X=2.365 $Y=1.515 $X2=0
+ $Y2=0
cc_170 N_A1_M1015_g N_A_337_74#_c_655_n 0.00374276f $X=2.47 $Y=0.74 $X2=0 $Y2=0
cc_171 A1 N_A_337_74#_c_655_n 0.0261369f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_172 N_A1_c_145_n N_A_337_74#_c_657_n 0.00592104f $X=2.365 $Y=1.515 $X2=0
+ $Y2=0
cc_173 N_A1_M1015_g N_A_337_74#_c_657_n 0.01343f $X=2.47 $Y=0.74 $X2=0 $Y2=0
cc_174 A1 N_A_337_74#_c_657_n 0.0901221f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_175 N_A1_M1015_g N_VGND_c_685_n 3.17863e-19 $X=2.47 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A1_M1005_g N_VGND_c_688_n 0.00278271f $X=1.61 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A1_M1015_g N_VGND_c_688_n 0.00278271f $X=2.47 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A1_M1005_g N_VGND_c_694_n 0.00357764f $X=1.61 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A1_M1015_g N_VGND_c_694_n 0.00360459f $X=2.47 $Y=0.74 $X2=0 $Y2=0
cc_180 N_S_c_208_n N_A_922_72#_c_303_n 0.0265275f $X=4.08 $Y=1.35 $X2=0 $Y2=0
cc_181 N_S_M1007_g N_A_922_72#_M1000_g 0.0335762f $X=4.065 $Y=2.4 $X2=0 $Y2=0
cc_182 N_S_c_227_p N_A_922_72#_M1000_g 0.0112656f $X=5.48 $Y=1.925 $X2=0 $Y2=0
cc_183 N_S_c_214_n N_A_922_72#_M1000_g 0.0116856f $X=4.675 $Y=1.72 $X2=0 $Y2=0
cc_184 N_S_M1004_g N_A_922_72#_M1012_g 0.0228079f $X=5.735 $Y=2.34 $X2=0 $Y2=0
cc_185 N_S_c_227_p N_A_922_72#_M1012_g 0.0168698f $X=5.48 $Y=1.925 $X2=0 $Y2=0
cc_186 N_S_c_209_n N_A_922_72#_M1012_g 0.00365291f $X=5.645 $Y=1.515 $X2=0 $Y2=0
cc_187 N_S_c_214_n N_A_922_72#_M1012_g 8.5127e-19 $X=4.675 $Y=1.72 $X2=0 $Y2=0
cc_188 N_S_c_212_n N_A_922_72#_c_304_n 0.021018f $X=5.652 $Y=1.35 $X2=0 $Y2=0
cc_189 N_S_c_227_p N_A_922_72#_c_305_n 0.023205f $X=5.48 $Y=1.925 $X2=0 $Y2=0
cc_190 N_S_c_209_n N_A_922_72#_c_305_n 0.0182306f $X=5.645 $Y=1.515 $X2=0 $Y2=0
cc_191 N_S_c_210_n N_A_922_72#_c_305_n 0.00118798f $X=5.645 $Y=1.515 $X2=0 $Y2=0
cc_192 N_S_c_212_n N_A_922_72#_c_305_n 9.47796e-19 $X=5.652 $Y=1.35 $X2=0 $Y2=0
cc_193 N_S_c_214_n N_A_922_72#_c_305_n 0.0147091f $X=4.675 $Y=1.72 $X2=0 $Y2=0
cc_194 N_S_c_227_p N_A_922_72#_c_330_n 0.00477724f $X=5.48 $Y=1.925 $X2=0 $Y2=0
cc_195 N_S_c_209_n N_A_922_72#_c_330_n 0.0222041f $X=5.645 $Y=1.515 $X2=0 $Y2=0
cc_196 N_S_c_210_n N_A_922_72#_c_330_n 0.00120563f $X=5.645 $Y=1.515 $X2=0 $Y2=0
cc_197 N_S_c_212_n N_A_922_72#_c_330_n 0.0115736f $X=5.652 $Y=1.35 $X2=0 $Y2=0
cc_198 N_S_c_212_n N_A_922_72#_c_306_n 0.00710009f $X=5.652 $Y=1.35 $X2=0 $Y2=0
cc_199 N_S_c_209_n N_A_922_72#_c_307_n 0.00117341f $X=5.645 $Y=1.515 $X2=0 $Y2=0
cc_200 N_S_c_212_n N_A_922_72#_c_307_n 0.00108392f $X=5.652 $Y=1.35 $X2=0 $Y2=0
cc_201 N_S_M1004_g N_A_922_72#_c_313_n 0.0108047f $X=5.735 $Y=2.34 $X2=0 $Y2=0
cc_202 N_S_c_227_p N_A_922_72#_c_313_n 0.00114029f $X=5.48 $Y=1.925 $X2=0 $Y2=0
cc_203 N_S_c_227_p N_A_922_72#_c_308_n 0.0133618f $X=5.48 $Y=1.925 $X2=0 $Y2=0
cc_204 N_S_c_209_n N_A_922_72#_c_308_n 0.036751f $X=5.645 $Y=1.515 $X2=0 $Y2=0
cc_205 N_S_c_210_n N_A_922_72#_c_308_n 0.0174221f $X=5.645 $Y=1.515 $X2=0 $Y2=0
cc_206 N_S_c_212_n N_A_922_72#_c_308_n 0.00413599f $X=5.652 $Y=1.35 $X2=0 $Y2=0
cc_207 N_S_c_227_p N_A_922_72#_c_309_n 0.00158047f $X=5.48 $Y=1.925 $X2=0 $Y2=0
cc_208 N_S_c_209_n N_A_922_72#_c_309_n 0.00139584f $X=5.645 $Y=1.515 $X2=0 $Y2=0
cc_209 N_S_c_210_n N_A_922_72#_c_309_n 0.0180157f $X=5.645 $Y=1.515 $X2=0 $Y2=0
cc_210 N_S_c_211_n N_A_922_72#_c_309_n 0.010191f $X=4.08 $Y=1.515 $X2=0 $Y2=0
cc_211 N_S_c_214_n N_A_922_72#_c_309_n 0.011295f $X=4.675 $Y=1.72 $X2=0 $Y2=0
cc_212 N_S_M1006_g N_Y_c_386_n 0.00191227f $X=3.615 $Y=2.4 $X2=0 $Y2=0
cc_213 N_S_c_207_n N_Y_c_384_n 0.00230277f $X=3.6 $Y=1.35 $X2=0 $Y2=0
cc_214 N_S_M1006_g N_A_121_368#_c_459_n 0.0180744f $X=3.615 $Y=2.4 $X2=0 $Y2=0
cc_215 N_S_M1007_g N_A_121_368#_c_459_n 0.00857755f $X=4.065 $Y=2.4 $X2=0 $Y2=0
cc_216 N_S_c_211_n N_A_121_368#_c_459_n 4.54581e-19 $X=4.08 $Y=1.515 $X2=0 $Y2=0
cc_217 N_S_c_213_n N_A_121_368#_c_459_n 0.0355443f $X=4.35 $Y=1.72 $X2=0 $Y2=0
cc_218 N_S_M1006_g N_A_121_368#_c_449_n 0.00397873f $X=3.615 $Y=2.4 $X2=0 $Y2=0
cc_219 N_S_c_227_p N_A_343_368#_M1000_s 0.00412048f $X=5.48 $Y=1.925 $X2=0 $Y2=0
cc_220 N_S_M1006_g N_A_343_368#_c_490_n 0.0112192f $X=3.615 $Y=2.4 $X2=0 $Y2=0
cc_221 N_S_M1007_g N_A_343_368#_c_490_n 0.0162985f $X=4.065 $Y=2.4 $X2=0 $Y2=0
cc_222 N_S_c_213_n N_A_343_368#_c_490_n 0.0084502f $X=4.35 $Y=1.72 $X2=0 $Y2=0
cc_223 N_S_c_214_n N_A_343_368#_c_490_n 0.0116927f $X=4.675 $Y=1.72 $X2=0 $Y2=0
cc_224 N_S_M1007_g N_A_343_368#_c_484_n 0.00231007f $X=4.065 $Y=2.4 $X2=0 $Y2=0
cc_225 N_S_c_227_p N_A_343_368#_c_484_n 0.0170259f $X=5.48 $Y=1.925 $X2=0 $Y2=0
cc_226 N_S_c_214_n N_VPWR_M1007_s 0.00690078f $X=4.675 $Y=1.72 $X2=0 $Y2=0
cc_227 N_S_c_227_p N_VPWR_M1012_d 0.00729957f $X=5.48 $Y=1.925 $X2=0 $Y2=0
cc_228 N_S_M1007_g N_VPWR_c_527_n 0.00454457f $X=4.065 $Y=2.4 $X2=0 $Y2=0
cc_229 N_S_M1004_g N_VPWR_c_528_n 0.00734822f $X=5.735 $Y=2.34 $X2=0 $Y2=0
cc_230 N_S_c_227_p N_VPWR_c_528_n 0.0245683f $X=5.48 $Y=1.925 $X2=0 $Y2=0
cc_231 N_S_c_210_n N_VPWR_c_528_n 4.22769e-19 $X=5.645 $Y=1.515 $X2=0 $Y2=0
cc_232 N_S_M1006_g N_VPWR_c_529_n 0.00393371f $X=3.615 $Y=2.4 $X2=0 $Y2=0
cc_233 N_S_M1007_g N_VPWR_c_529_n 0.00393371f $X=4.065 $Y=2.4 $X2=0 $Y2=0
cc_234 N_S_M1004_g N_VPWR_c_534_n 0.00567889f $X=5.735 $Y=2.34 $X2=0 $Y2=0
cc_235 N_S_M1006_g N_VPWR_c_526_n 0.00503521f $X=3.615 $Y=2.4 $X2=0 $Y2=0
cc_236 N_S_M1007_g N_VPWR_c_526_n 0.00499997f $X=4.065 $Y=2.4 $X2=0 $Y2=0
cc_237 N_S_M1004_g N_VPWR_c_526_n 0.00610055f $X=5.735 $Y=2.34 $X2=0 $Y2=0
cc_238 N_S_M1006_g N_VPWR_c_536_n 0.00543666f $X=3.615 $Y=2.4 $X2=0 $Y2=0
cc_239 N_S_c_207_n N_A_115_74#_c_593_n 0.00340328f $X=3.6 $Y=1.35 $X2=0 $Y2=0
cc_240 N_S_c_208_n N_A_115_74#_c_610_n 7.12069e-19 $X=4.08 $Y=1.35 $X2=0 $Y2=0
cc_241 N_S_c_207_n N_A_115_74#_c_611_n 0.0135909f $X=3.6 $Y=1.35 $X2=0 $Y2=0
cc_242 N_S_c_208_n N_A_115_74#_c_611_n 0.0143324f $X=4.08 $Y=1.35 $X2=0 $Y2=0
cc_243 N_S_c_213_n N_A_115_74#_c_611_n 0.0179481f $X=4.35 $Y=1.72 $X2=0 $Y2=0
cc_244 N_S_c_207_n N_A_337_74#_c_656_n 0.00537817f $X=3.6 $Y=1.35 $X2=0 $Y2=0
cc_245 N_S_c_208_n N_A_337_74#_c_656_n 0.00678548f $X=4.08 $Y=1.35 $X2=0 $Y2=0
cc_246 N_S_c_211_n N_A_337_74#_c_656_n 0.00399478f $X=4.08 $Y=1.515 $X2=0 $Y2=0
cc_247 N_S_c_207_n N_A_337_74#_c_657_n 0.00983725f $X=3.6 $Y=1.35 $X2=0 $Y2=0
cc_248 N_S_c_213_n N_A_337_74#_c_657_n 0.0420755f $X=4.35 $Y=1.72 $X2=0 $Y2=0
cc_249 N_S_c_207_n N_VGND_c_685_n 0.00546687f $X=3.6 $Y=1.35 $X2=0 $Y2=0
cc_250 N_S_c_208_n N_VGND_c_686_n 0.00383345f $X=4.08 $Y=1.35 $X2=0 $Y2=0
cc_251 N_S_c_212_n N_VGND_c_687_n 0.00488969f $X=5.652 $Y=1.35 $X2=0 $Y2=0
cc_252 N_S_c_207_n N_VGND_c_690_n 0.0038134f $X=3.6 $Y=1.35 $X2=0 $Y2=0
cc_253 N_S_c_208_n N_VGND_c_690_n 0.0038134f $X=4.08 $Y=1.35 $X2=0 $Y2=0
cc_254 N_S_c_212_n N_VGND_c_693_n 0.00417655f $X=5.652 $Y=1.35 $X2=0 $Y2=0
cc_255 N_S_c_207_n N_VGND_c_694_n 0.00508379f $X=3.6 $Y=1.35 $X2=0 $Y2=0
cc_256 N_S_c_208_n N_VGND_c_694_n 0.00508379f $X=4.08 $Y=1.35 $X2=0 $Y2=0
cc_257 N_S_c_212_n N_VGND_c_694_n 0.00479212f $X=5.652 $Y=1.35 $X2=0 $Y2=0
cc_258 N_A_922_72#_M1000_g N_A_121_368#_c_459_n 0.00143444f $X=4.7 $Y=2.4 $X2=0
+ $Y2=0
cc_259 N_A_922_72#_M1000_g N_A_343_368#_c_490_n 0.0131658f $X=4.7 $Y=2.4 $X2=0
+ $Y2=0
cc_260 N_A_922_72#_M1000_g N_A_343_368#_c_484_n 0.0163279f $X=4.7 $Y=2.4 $X2=0
+ $Y2=0
cc_261 N_A_922_72#_M1012_g N_A_343_368#_c_484_n 0.0118975f $X=5.15 $Y=2.4 $X2=0
+ $Y2=0
cc_262 N_A_922_72#_M1000_g N_VPWR_c_527_n 0.0041787f $X=4.7 $Y=2.4 $X2=0 $Y2=0
cc_263 N_A_922_72#_M1012_g N_VPWR_c_528_n 0.00623718f $X=5.15 $Y=2.4 $X2=0 $Y2=0
cc_264 N_A_922_72#_c_313_n N_VPWR_c_528_n 0.0228728f $X=5.96 $Y=2.265 $X2=0
+ $Y2=0
cc_265 N_A_922_72#_M1000_g N_VPWR_c_531_n 0.00387245f $X=4.7 $Y=2.4 $X2=0 $Y2=0
cc_266 N_A_922_72#_M1012_g N_VPWR_c_531_n 0.005209f $X=5.15 $Y=2.4 $X2=0 $Y2=0
cc_267 N_A_922_72#_c_313_n N_VPWR_c_534_n 0.0105092f $X=5.96 $Y=2.265 $X2=0
+ $Y2=0
cc_268 N_A_922_72#_M1000_g N_VPWR_c_526_n 0.00487387f $X=4.7 $Y=2.4 $X2=0 $Y2=0
cc_269 N_A_922_72#_M1012_g N_VPWR_c_526_n 0.00986727f $X=5.15 $Y=2.4 $X2=0 $Y2=0
cc_270 N_A_922_72#_c_313_n N_VPWR_c_526_n 0.0120294f $X=5.96 $Y=2.265 $X2=0
+ $Y2=0
cc_271 N_A_922_72#_c_305_n N_A_115_74#_M1001_s 6.07965e-19 $X=5.075 $Y=1.505
+ $X2=0 $Y2=0
cc_272 N_A_922_72#_c_362_p N_A_115_74#_M1001_s 0.00368553f $X=5.24 $Y=1.095
+ $X2=0 $Y2=0
cc_273 N_A_922_72#_c_303_n N_A_115_74#_c_610_n 0.00525305f $X=4.685 $Y=1.34
+ $X2=0 $Y2=0
cc_274 N_A_922_72#_c_304_n N_A_115_74#_c_610_n 0.00408973f $X=5.165 $Y=1.34
+ $X2=0 $Y2=0
cc_275 N_A_922_72#_c_362_p N_A_115_74#_c_610_n 0.0118787f $X=5.24 $Y=1.095 $X2=0
+ $Y2=0
cc_276 N_A_922_72#_c_309_n N_A_115_74#_c_610_n 0.00212274f $X=5.165 $Y=1.505
+ $X2=0 $Y2=0
cc_277 N_A_922_72#_c_303_n N_A_115_74#_c_611_n 0.0117154f $X=4.685 $Y=1.34 $X2=0
+ $Y2=0
cc_278 N_A_922_72#_c_303_n N_A_337_74#_c_656_n 0.0011501f $X=4.685 $Y=1.34 $X2=0
+ $Y2=0
cc_279 N_A_922_72#_c_330_n N_VGND_M1017_d 0.00890916f $X=5.795 $Y=1.095 $X2=0
+ $Y2=0
cc_280 N_A_922_72#_c_303_n N_VGND_c_686_n 0.00383345f $X=4.685 $Y=1.34 $X2=0
+ $Y2=0
cc_281 N_A_922_72#_c_304_n N_VGND_c_687_n 0.0072762f $X=5.165 $Y=1.34 $X2=0
+ $Y2=0
cc_282 N_A_922_72#_c_330_n N_VGND_c_687_n 0.0257093f $X=5.795 $Y=1.095 $X2=0
+ $Y2=0
cc_283 N_A_922_72#_c_306_n N_VGND_c_687_n 0.0105452f $X=5.96 $Y=0.735 $X2=0
+ $Y2=0
cc_284 N_A_922_72#_c_303_n N_VGND_c_692_n 0.00379069f $X=4.685 $Y=1.34 $X2=0
+ $Y2=0
cc_285 N_A_922_72#_c_304_n N_VGND_c_692_n 0.00472994f $X=5.165 $Y=1.34 $X2=0
+ $Y2=0
cc_286 N_A_922_72#_c_306_n N_VGND_c_693_n 0.00814182f $X=5.96 $Y=0.735 $X2=0
+ $Y2=0
cc_287 N_A_922_72#_c_303_n N_VGND_c_694_n 0.00508379f $X=4.685 $Y=1.34 $X2=0
+ $Y2=0
cc_288 N_A_922_72#_c_304_n N_VGND_c_694_n 0.00508379f $X=5.165 $Y=1.34 $X2=0
+ $Y2=0
cc_289 N_A_922_72#_c_306_n N_VGND_c_694_n 0.011178f $X=5.96 $Y=0.735 $X2=0 $Y2=0
cc_290 N_Y_c_386_n N_A_121_368#_M1002_s 0.00483913f $X=2.68 $Y=2.03 $X2=-0.19
+ $Y2=-0.245
cc_291 N_Y_c_386_n N_A_121_368#_c_447_n 0.0182218f $X=2.68 $Y=2.03 $X2=0 $Y2=0
cc_292 Y N_A_121_368#_c_447_n 0.0207538f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_293 N_Y_M1011_d N_A_121_368#_c_448_n 0.0166565f $X=1.095 $Y=1.84 $X2=0 $Y2=0
cc_294 N_Y_M1014_d N_A_121_368#_c_448_n 0.00568251f $X=2.545 $Y=1.84 $X2=0 $Y2=0
cc_295 N_Y_c_386_n N_A_121_368#_c_448_n 0.114813f $X=2.68 $Y=2.03 $X2=0 $Y2=0
cc_296 N_Y_c_386_n N_A_121_368#_c_449_n 0.00965074f $X=2.68 $Y=2.03 $X2=0 $Y2=0
cc_297 N_Y_c_386_n N_A_343_368#_M1003_s 0.013188f $X=2.68 $Y=2.03 $X2=-0.19
+ $Y2=-0.245
cc_298 N_Y_M1014_d N_A_343_368#_c_483_n 0.00672569f $X=2.545 $Y=1.84 $X2=0 $Y2=0
cc_299 Y N_VPWR_c_533_n 0.0159175f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_300 Y N_VPWR_c_526_n 0.0131305f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_301 N_Y_c_381_n N_A_115_74#_M1008_d 0.00299895f $X=2.58 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_302 N_Y_M1016_s N_A_115_74#_c_594_n 0.0129407f $X=1.095 $Y=0.37 $X2=0 $Y2=0
cc_303 N_Y_c_381_n N_A_115_74#_c_594_n 0.0738597f $X=2.58 $Y=0.34 $X2=0 $Y2=0
cc_304 N_Y_M1015_s N_A_115_74#_c_592_n 0.00759772f $X=2.545 $Y=0.37 $X2=0 $Y2=0
cc_305 N_Y_c_381_n N_A_115_74#_c_592_n 0.00477629f $X=2.58 $Y=0.34 $X2=0 $Y2=0
cc_306 N_Y_c_384_n N_A_115_74#_c_592_n 0.0228342f $X=2.745 $Y=0.34 $X2=0 $Y2=0
cc_307 N_Y_c_380_n N_A_115_74#_c_596_n 0.0297541f $X=0.285 $Y=0.515 $X2=0 $Y2=0
cc_308 N_Y_c_381_n N_A_115_74#_c_596_n 0.0197539f $X=2.58 $Y=0.34 $X2=0 $Y2=0
cc_309 N_Y_c_381_n N_A_115_74#_c_606_n 0.00792639f $X=2.58 $Y=0.34 $X2=0 $Y2=0
cc_310 N_Y_c_381_n N_A_337_74#_M1005_d 0.00737333f $X=2.58 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_311 N_Y_M1015_s N_A_337_74#_c_657_n 0.00324248f $X=2.545 $Y=0.37 $X2=0 $Y2=0
cc_312 N_Y_c_384_n N_VGND_c_685_n 0.0158437f $X=2.745 $Y=0.34 $X2=0 $Y2=0
cc_313 N_Y_c_381_n N_VGND_c_688_n 0.135211f $X=2.58 $Y=0.34 $X2=0 $Y2=0
cc_314 N_Y_c_382_n N_VGND_c_688_n 0.0260778f $X=0.45 $Y=0.34 $X2=0 $Y2=0
cc_315 N_Y_c_384_n N_VGND_c_688_n 0.0222656f $X=2.745 $Y=0.34 $X2=0 $Y2=0
cc_316 N_Y_M1016_s N_VGND_c_694_n 0.00246676f $X=1.095 $Y=0.37 $X2=0 $Y2=0
cc_317 N_Y_c_381_n N_VGND_c_694_n 0.0774633f $X=2.58 $Y=0.34 $X2=0 $Y2=0
cc_318 N_Y_c_382_n N_VGND_c_694_n 0.014076f $X=0.45 $Y=0.34 $X2=0 $Y2=0
cc_319 N_Y_c_384_n N_VGND_c_694_n 0.0125202f $X=2.745 $Y=0.34 $X2=0 $Y2=0
cc_320 N_A_121_368#_c_448_n N_A_343_368#_M1003_s 0.013697f $X=3.015 $Y=2.232
+ $X2=-0.19 $Y2=1.66
cc_321 N_A_121_368#_c_459_n N_A_343_368#_c_483_n 0.00885658f $X=3.84 $Y=2.175
+ $X2=0 $Y2=0
cc_322 N_A_121_368#_M1006_d N_A_343_368#_c_490_n 0.00442572f $X=3.705 $Y=1.84
+ $X2=0 $Y2=0
cc_323 N_A_121_368#_c_459_n N_A_343_368#_c_490_n 0.0268434f $X=3.84 $Y=2.175
+ $X2=0 $Y2=0
cc_324 N_A_121_368#_c_448_n N_A_343_368#_c_485_n 0.0496355f $X=3.015 $Y=2.232
+ $X2=0 $Y2=0
cc_325 N_A_121_368#_c_449_n N_A_343_368#_c_488_n 0.0496355f $X=3.185 $Y=2.232
+ $X2=0 $Y2=0
cc_326 N_A_121_368#_c_459_n N_A_343_368#_c_507_n 0.00893008f $X=3.84 $Y=2.175
+ $X2=0 $Y2=0
cc_327 N_A_121_368#_c_459_n N_VPWR_M1006_s 0.016677f $X=3.84 $Y=2.175 $X2=-0.19
+ $Y2=1.66
cc_328 N_A_121_368#_c_449_n N_VPWR_M1006_s 0.00612985f $X=3.185 $Y=2.232
+ $X2=-0.19 $Y2=1.66
cc_329 N_A_121_368#_c_447_n N_VPWR_c_533_n 0.0145721f $X=0.78 $Y=2.37 $X2=0
+ $Y2=0
cc_330 N_A_121_368#_c_447_n N_VPWR_c_526_n 0.0119833f $X=0.78 $Y=2.37 $X2=0
+ $Y2=0
cc_331 N_A_343_368#_c_483_n N_VPWR_M1006_s 0.00857931f $X=3.355 $Y=2.71
+ $X2=-0.19 $Y2=1.66
cc_332 N_A_343_368#_c_507_n N_VPWR_M1006_s 0.00726657f $X=3.44 $Y=2.595
+ $X2=-0.19 $Y2=1.66
cc_333 N_A_343_368#_c_490_n N_VPWR_M1007_s 0.0109562f $X=4.76 $Y=2.595 $X2=0
+ $Y2=0
cc_334 N_A_343_368#_c_490_n N_VPWR_c_527_n 0.0261179f $X=4.76 $Y=2.595 $X2=0
+ $Y2=0
cc_335 N_A_343_368#_c_484_n N_VPWR_c_527_n 0.00489696f $X=4.925 $Y=2.265 $X2=0
+ $Y2=0
cc_336 N_A_343_368#_c_484_n N_VPWR_c_528_n 0.0308084f $X=4.925 $Y=2.265 $X2=0
+ $Y2=0
cc_337 N_A_343_368#_c_490_n N_VPWR_c_529_n 0.00989602f $X=4.76 $Y=2.595 $X2=0
+ $Y2=0
cc_338 N_A_343_368#_c_490_n N_VPWR_c_531_n 0.0028743f $X=4.76 $Y=2.595 $X2=0
+ $Y2=0
cc_339 N_A_343_368#_c_484_n N_VPWR_c_531_n 0.0144623f $X=4.925 $Y=2.265 $X2=0
+ $Y2=0
cc_340 N_A_343_368#_c_483_n N_VPWR_c_533_n 0.0145144f $X=3.355 $Y=2.71 $X2=0
+ $Y2=0
cc_341 N_A_343_368#_c_485_n N_VPWR_c_533_n 0.0245025f $X=2.23 $Y=2.79 $X2=0
+ $Y2=0
cc_342 N_A_343_368#_c_483_n N_VPWR_c_526_n 0.0218064f $X=3.355 $Y=2.71 $X2=0
+ $Y2=0
cc_343 N_A_343_368#_c_490_n N_VPWR_c_526_n 0.0241598f $X=4.76 $Y=2.595 $X2=0
+ $Y2=0
cc_344 N_A_343_368#_c_485_n N_VPWR_c_526_n 0.0248593f $X=2.23 $Y=2.79 $X2=0
+ $Y2=0
cc_345 N_A_343_368#_c_507_n N_VPWR_c_526_n 0.00239403f $X=3.44 $Y=2.595 $X2=0
+ $Y2=0
cc_346 N_A_343_368#_c_484_n N_VPWR_c_526_n 0.0118344f $X=4.925 $Y=2.265 $X2=0
+ $Y2=0
cc_347 N_A_343_368#_c_483_n N_VPWR_c_536_n 0.0205871f $X=3.355 $Y=2.71 $X2=0
+ $Y2=0
cc_348 N_A_343_368#_c_507_n N_VPWR_c_536_n 0.00864628f $X=3.44 $Y=2.595 $X2=0
+ $Y2=0
cc_349 N_A_115_74#_c_594_n N_A_337_74#_M1005_d 0.0140992f $X=2.24 $Y=0.68
+ $X2=-0.19 $Y2=-0.245
cc_350 N_A_115_74#_c_606_n N_A_337_74#_M1005_d 0.00494202f $X=2.325 $Y=0.68
+ $X2=-0.19 $Y2=-0.245
cc_351 N_A_115_74#_c_611_n N_A_337_74#_M1010_d 0.00600194f $X=4.735 $Y=0.665
+ $X2=0 $Y2=0
cc_352 N_A_115_74#_c_594_n N_A_337_74#_c_655_n 0.0250821f $X=2.24 $Y=0.68 $X2=0
+ $Y2=0
cc_353 N_A_115_74#_c_611_n N_A_337_74#_c_656_n 0.0196351f $X=4.735 $Y=0.665
+ $X2=0 $Y2=0
cc_354 N_A_115_74#_c_594_n N_A_337_74#_c_657_n 0.00766912f $X=2.24 $Y=0.68 $X2=0
+ $Y2=0
cc_355 N_A_115_74#_c_592_n N_A_337_74#_c_657_n 0.0443759f $X=3.08 $Y=0.835 $X2=0
+ $Y2=0
cc_356 N_A_115_74#_c_606_n N_A_337_74#_c_657_n 0.00844404f $X=2.325 $Y=0.68
+ $X2=0 $Y2=0
cc_357 N_A_115_74#_c_593_n N_A_337_74#_c_657_n 0.0128864f $X=3.165 $Y=0.745
+ $X2=0 $Y2=0
cc_358 N_A_115_74#_c_611_n N_A_337_74#_c_657_n 0.0175892f $X=4.735 $Y=0.665
+ $X2=0 $Y2=0
cc_359 N_A_115_74#_c_593_n N_VGND_M1010_s 0.00472881f $X=3.165 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_360 N_A_115_74#_c_611_n N_VGND_M1010_s 0.00642911f $X=4.735 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_361 N_A_115_74#_c_611_n N_VGND_M1013_s 0.0111719f $X=4.735 $Y=0.665 $X2=0
+ $Y2=0
cc_362 N_A_115_74#_c_593_n N_VGND_c_685_n 0.0086353f $X=3.165 $Y=0.745 $X2=0
+ $Y2=0
cc_363 N_A_115_74#_c_611_n N_VGND_c_685_n 0.0167914f $X=4.735 $Y=0.665 $X2=0
+ $Y2=0
cc_364 N_A_115_74#_c_611_n N_VGND_c_686_n 0.0262846f $X=4.735 $Y=0.665 $X2=0
+ $Y2=0
cc_365 N_A_115_74#_c_592_n N_VGND_c_688_n 0.00248688f $X=3.08 $Y=0.835 $X2=0
+ $Y2=0
cc_366 N_A_115_74#_c_593_n N_VGND_c_688_n 0.00104648f $X=3.165 $Y=0.745 $X2=0
+ $Y2=0
cc_367 N_A_115_74#_c_611_n N_VGND_c_690_n 0.0102331f $X=4.735 $Y=0.665 $X2=0
+ $Y2=0
cc_368 N_A_115_74#_c_610_n N_VGND_c_692_n 0.00824986f $X=4.925 $Y=0.665 $X2=0
+ $Y2=0
cc_369 N_A_115_74#_c_611_n N_VGND_c_692_n 0.00241616f $X=4.735 $Y=0.665 $X2=0
+ $Y2=0
cc_370 N_A_115_74#_c_592_n N_VGND_c_694_n 0.00544547f $X=3.08 $Y=0.835 $X2=0
+ $Y2=0
cc_371 N_A_115_74#_c_593_n N_VGND_c_694_n 0.00220611f $X=3.165 $Y=0.745 $X2=0
+ $Y2=0
cc_372 N_A_115_74#_c_610_n N_VGND_c_694_n 0.0122645f $X=4.925 $Y=0.665 $X2=0
+ $Y2=0
cc_373 N_A_115_74#_c_611_n N_VGND_c_694_n 0.0278432f $X=4.735 $Y=0.665 $X2=0
+ $Y2=0
cc_374 N_A_337_74#_c_657_n N_VGND_M1010_s 0.00518087f $X=3.65 $Y=1.13 $X2=-0.19
+ $Y2=-0.245

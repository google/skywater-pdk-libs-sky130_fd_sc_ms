* File: sky130_fd_sc_ms__buf_16.pex.spice
* Created: Wed Sep  2 11:59:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__BUF_16%A_83_260# 1 2 3 4 5 6 21 25 29 33 37 41 45 49
+ 53 57 61 65 69 73 77 81 85 89 93 97 101 105 109 113 117 121 125 129 133 137
+ 141 145 147 148 149 150 153 157 159 161 165 169 171 173 175 177 181 186 187
+ 189 190 216 217 226 233 240 247 254 261 268 272
c469 272 0 8.31019e-20 $X=7.38 $Y=1.465
c470 216 0 8.59108e-19 $X=7.505 $Y=1.665
r471 271 272 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.305 $Y=1.465
+ $X2=7.38 $Y2=1.465
r472 270 271 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=6.95 $Y=1.465
+ $X2=7.305 $Y2=1.465
r473 269 270 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=6.855 $Y=1.465
+ $X2=6.95 $Y2=1.465
r474 267 269 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=6.665 $Y=1.465
+ $X2=6.855 $Y2=1.465
r475 267 268 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.665
+ $Y=1.465 $X2=6.665 $Y2=1.465
r476 265 267 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=6.405 $Y=1.465
+ $X2=6.665 $Y2=1.465
r477 264 265 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=6.38 $Y=1.465
+ $X2=6.405 $Y2=1.465
r478 263 264 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=5.955 $Y=1.465
+ $X2=6.38 $Y2=1.465
r479 262 263 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=5.95 $Y=1.465
+ $X2=5.955 $Y2=1.465
r480 260 262 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.74 $Y=1.465
+ $X2=5.95 $Y2=1.465
r481 260 261 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.74
+ $Y=1.465 $X2=5.74 $Y2=1.465
r482 258 260 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=5.505 $Y=1.465
+ $X2=5.74 $Y2=1.465
r483 257 258 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.38 $Y=1.465
+ $X2=5.505 $Y2=1.465
r484 256 257 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=5.055 $Y=1.465
+ $X2=5.38 $Y2=1.465
r485 255 256 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=4.95 $Y=1.465
+ $X2=5.055 $Y2=1.465
r486 253 255 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=4.72 $Y=1.465
+ $X2=4.95 $Y2=1.465
r487 253 254 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.72
+ $Y=1.465 $X2=4.72 $Y2=1.465
r488 251 253 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=4.605 $Y=1.465
+ $X2=4.72 $Y2=1.465
r489 250 251 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=4.38 $Y=1.465
+ $X2=4.605 $Y2=1.465
r490 249 250 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=4.155 $Y=1.465
+ $X2=4.38 $Y2=1.465
r491 248 249 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=3.95 $Y=1.465
+ $X2=4.155 $Y2=1.465
r492 246 248 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.86 $Y=1.465
+ $X2=3.95 $Y2=1.465
r493 246 247 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.86
+ $Y=1.465 $X2=3.86 $Y2=1.465
r494 244 246 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=3.705 $Y=1.465
+ $X2=3.86 $Y2=1.465
r495 243 244 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=3.52 $Y=1.465
+ $X2=3.705 $Y2=1.465
r496 242 243 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=3.255 $Y=1.465
+ $X2=3.52 $Y2=1.465
r497 241 242 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=1.465
+ $X2=3.255 $Y2=1.465
r498 239 241 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=2.995 $Y=1.465
+ $X2=3.09 $Y2=1.465
r499 239 240 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.995
+ $Y=1.465 $X2=2.995 $Y2=1.465
r500 237 239 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=2.805 $Y=1.465
+ $X2=2.995 $Y2=1.465
r501 236 237 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=2.66 $Y=1.465
+ $X2=2.805 $Y2=1.465
r502 235 236 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=2.355 $Y=1.465
+ $X2=2.66 $Y2=1.465
r503 234 235 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=2.23 $Y=1.465
+ $X2=2.355 $Y2=1.465
r504 232 234 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=2.035 $Y=1.465
+ $X2=2.23 $Y2=1.465
r505 232 233 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.035
+ $Y=1.465 $X2=2.035 $Y2=1.465
r506 230 232 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.855 $Y=1.465
+ $X2=2.035 $Y2=1.465
r507 229 230 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=1.8 $Y=1.465
+ $X2=1.855 $Y2=1.465
r508 228 229 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=1.405 $Y=1.465
+ $X2=1.8 $Y2=1.465
r509 227 228 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=1.37 $Y=1.465
+ $X2=1.405 $Y2=1.465
r510 225 227 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=1.15 $Y=1.465
+ $X2=1.37 $Y2=1.465
r511 225 226 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.465 $X2=1.15 $Y2=1.465
r512 223 225 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.955 $Y=1.465
+ $X2=1.15 $Y2=1.465
r513 222 223 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.94 $Y=1.465
+ $X2=0.955 $Y2=1.465
r514 221 222 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.51 $Y=1.465
+ $X2=0.94 $Y2=1.465
r515 219 221 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=0.505 $Y=1.465
+ $X2=0.51 $Y2=1.465
r516 216 217 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.505 $Y=1.665
+ $X2=7.505 $Y2=1.665
r517 214 268 7.43512 $w=3.08e-07 $l=2e-07 $layer=LI1_cond $X=6.655 $Y=1.665
+ $X2=6.655 $Y2=1.465
r518 213 216 0.548572 $w=2.3e-07 $l=8.55e-07 $layer=MET1_cond $X=6.65 $Y=1.665
+ $X2=7.505 $Y2=1.665
r519 213 214 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.65 $Y=1.665
+ $X2=6.65 $Y2=1.665
r520 211 261 7.43512 $w=3.08e-07 $l=2e-07 $layer=LI1_cond $X=5.735 $Y=1.665
+ $X2=5.735 $Y2=1.465
r521 210 213 0.587068 $w=2.3e-07 $l=9.15e-07 $layer=MET1_cond $X=5.735 $Y=1.665
+ $X2=6.65 $Y2=1.665
r522 210 211 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.735 $Y=1.665
+ $X2=5.735 $Y2=1.665
r523 208 254 8.21549 $w=2.97e-07 $l=2e-07 $layer=LI1_cond $X=4.71 $Y=1.665
+ $X2=4.71 $Y2=1.465
r524 207 210 0.622356 $w=2.3e-07 $l=9.7e-07 $layer=MET1_cond $X=4.765 $Y=1.665
+ $X2=5.735 $Y2=1.665
r525 207 208 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.765 $Y=1.665
+ $X2=4.765 $Y2=1.665
r526 205 247 6.61247 $w=3.69e-07 $l=2e-07 $layer=LI1_cond $X=3.85 $Y=1.665
+ $X2=3.85 $Y2=1.465
r527 204 207 0.564612 $w=2.3e-07 $l=8.8e-07 $layer=MET1_cond $X=3.885 $Y=1.665
+ $X2=4.765 $Y2=1.665
r528 204 205 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.885 $Y=1.665
+ $X2=3.885 $Y2=1.665
r529 202 240 7.81317 $w=2.93e-07 $l=2e-07 $layer=LI1_cond $X=2.992 $Y=1.665
+ $X2=2.992 $Y2=1.465
r530 201 204 0.571028 $w=2.3e-07 $l=8.9e-07 $layer=MET1_cond $X=2.995 $Y=1.665
+ $X2=3.885 $Y2=1.665
r531 201 202 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.995 $Y=1.665
+ $X2=2.995 $Y2=1.665
r532 199 233 8.08732 $w=2.83e-07 $l=2e-07 $layer=LI1_cond $X=2.032 $Y=1.665
+ $X2=2.032 $Y2=1.465
r533 198 201 0.61594 $w=2.3e-07 $l=9.6e-07 $layer=MET1_cond $X=2.035 $Y=1.665
+ $X2=2.995 $Y2=1.665
r534 198 199 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.035 $Y=1.665
+ $X2=2.035 $Y2=1.665
r535 195 226 7.43512 $w=3.08e-07 $l=2e-07 $layer=LI1_cond $X=1.14 $Y=1.665
+ $X2=1.14 $Y2=1.465
r536 194 198 0.574236 $w=2.3e-07 $l=8.95e-07 $layer=MET1_cond $X=1.14 $Y=1.665
+ $X2=2.035 $Y2=1.665
r537 194 195 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.14 $Y=1.665
+ $X2=1.14 $Y2=1.665
r538 184 217 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.505 $Y=1.95
+ $X2=7.505 $Y2=1.665
r539 183 217 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=7.505 $Y=1.18
+ $X2=7.505 $Y2=1.665
r540 179 181 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=9.82 $Y=1.01
+ $X2=9.82 $Y2=0.515
r541 175 192 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.83 $Y=2.12
+ $X2=9.83 $Y2=2.035
r542 175 177 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=9.83 $Y=2.12
+ $X2=9.83 $Y2=2.815
r543 174 189 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.095 $Y=2.035
+ $X2=8.93 $Y2=2.035
r544 173 192 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.665 $Y=2.035
+ $X2=9.83 $Y2=2.035
r545 173 174 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=9.665 $Y=2.035
+ $X2=9.095 $Y2=2.035
r546 172 190 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.97 $Y=1.095
+ $X2=8.885 $Y2=1.095
r547 171 179 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.695 $Y=1.095
+ $X2=9.82 $Y2=1.01
r548 171 172 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=9.695 $Y=1.095
+ $X2=8.97 $Y2=1.095
r549 167 190 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.885 $Y=1.01
+ $X2=8.885 $Y2=1.095
r550 167 169 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=8.885 $Y=1.01
+ $X2=8.885 $Y2=0.515
r551 163 189 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.93 $Y=2.12
+ $X2=8.93 $Y2=2.035
r552 163 165 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=8.93 $Y=2.12
+ $X2=8.93 $Y2=2.815
r553 162 186 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.195 $Y=2.035
+ $X2=8.03 $Y2=2.035
r554 161 189 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.765 $Y=2.035
+ $X2=8.93 $Y2=2.035
r555 161 162 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.765 $Y=2.035
+ $X2=8.195 $Y2=2.035
r556 160 187 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.11 $Y=1.095
+ $X2=8.025 $Y2=1.095
r557 159 190 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.8 $Y=1.095
+ $X2=8.885 $Y2=1.095
r558 159 160 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.8 $Y=1.095
+ $X2=8.11 $Y2=1.095
r559 155 187 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.025 $Y=1.01
+ $X2=8.025 $Y2=1.095
r560 155 157 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=8.025 $Y=1.01
+ $X2=8.025 $Y2=0.515
r561 151 186 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.03 $Y=2.12
+ $X2=8.03 $Y2=2.035
r562 151 153 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=8.03 $Y=2.12
+ $X2=8.03 $Y2=2.815
r563 150 184 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.59 $Y=2.035
+ $X2=7.505 $Y2=1.95
r564 149 186 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.865 $Y=2.035
+ $X2=8.03 $Y2=2.035
r565 149 150 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.865 $Y=2.035
+ $X2=7.59 $Y2=2.035
r566 148 183 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.59 $Y=1.095
+ $X2=7.505 $Y2=1.18
r567 147 187 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.94 $Y=1.095
+ $X2=8.025 $Y2=1.095
r568 147 148 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.94 $Y=1.095
+ $X2=7.59 $Y2=1.095
r569 143 272 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.38 $Y=1.3
+ $X2=7.38 $Y2=1.465
r570 143 145 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.38 $Y=1.3
+ $X2=7.38 $Y2=0.74
r571 139 271 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.305 $Y=1.63
+ $X2=7.305 $Y2=1.465
r572 139 141 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=7.305 $Y=1.63
+ $X2=7.305 $Y2=2.4
r573 135 270 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.95 $Y=1.3
+ $X2=6.95 $Y2=1.465
r574 135 137 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.95 $Y=1.3
+ $X2=6.95 $Y2=0.74
r575 131 269 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.855 $Y=1.63
+ $X2=6.855 $Y2=1.465
r576 131 133 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=6.855 $Y=1.63
+ $X2=6.855 $Y2=2.4
r577 127 265 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.405 $Y=1.63
+ $X2=6.405 $Y2=1.465
r578 127 129 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=6.405 $Y=1.63
+ $X2=6.405 $Y2=2.4
r579 123 264 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.38 $Y=1.3
+ $X2=6.38 $Y2=1.465
r580 123 125 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.38 $Y=1.3
+ $X2=6.38 $Y2=0.74
r581 119 262 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.95 $Y=1.3
+ $X2=5.95 $Y2=1.465
r582 119 121 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.95 $Y=1.3
+ $X2=5.95 $Y2=0.74
r583 115 263 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.955 $Y=1.63
+ $X2=5.955 $Y2=1.465
r584 115 117 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=5.955 $Y=1.63
+ $X2=5.955 $Y2=2.4
r585 111 258 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.505 $Y=1.63
+ $X2=5.505 $Y2=1.465
r586 111 113 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=5.505 $Y=1.63
+ $X2=5.505 $Y2=2.4
r587 107 257 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.38 $Y=1.3
+ $X2=5.38 $Y2=1.465
r588 107 109 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.38 $Y=1.3
+ $X2=5.38 $Y2=0.74
r589 103 256 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.055 $Y=1.63
+ $X2=5.055 $Y2=1.465
r590 103 105 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=5.055 $Y=1.63
+ $X2=5.055 $Y2=2.4
r591 99 255 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.95 $Y=1.3
+ $X2=4.95 $Y2=1.465
r592 99 101 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.95 $Y=1.3
+ $X2=4.95 $Y2=0.74
r593 95 251 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.605 $Y=1.63
+ $X2=4.605 $Y2=1.465
r594 95 97 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.605 $Y=1.63
+ $X2=4.605 $Y2=2.4
r595 91 250 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.38 $Y=1.3
+ $X2=4.38 $Y2=1.465
r596 91 93 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.38 $Y=1.3
+ $X2=4.38 $Y2=0.74
r597 87 249 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.155 $Y=1.63
+ $X2=4.155 $Y2=1.465
r598 87 89 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.155 $Y=1.63
+ $X2=4.155 $Y2=2.4
r599 83 248 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.95 $Y=1.3
+ $X2=3.95 $Y2=1.465
r600 83 85 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.95 $Y=1.3
+ $X2=3.95 $Y2=0.74
r601 79 244 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.705 $Y=1.63
+ $X2=3.705 $Y2=1.465
r602 79 81 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=3.705 $Y=1.63
+ $X2=3.705 $Y2=2.4
r603 75 243 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.52 $Y=1.3
+ $X2=3.52 $Y2=1.465
r604 75 77 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.52 $Y=1.3
+ $X2=3.52 $Y2=0.74
r605 71 242 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.255 $Y=1.63
+ $X2=3.255 $Y2=1.465
r606 71 73 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=3.255 $Y=1.63
+ $X2=3.255 $Y2=2.4
r607 67 241 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=1.3
+ $X2=3.09 $Y2=1.465
r608 67 69 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.09 $Y=1.3
+ $X2=3.09 $Y2=0.74
r609 63 237 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.805 $Y=1.63
+ $X2=2.805 $Y2=1.465
r610 63 65 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=2.805 $Y=1.63
+ $X2=2.805 $Y2=2.4
r611 59 236 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.66 $Y=1.3
+ $X2=2.66 $Y2=1.465
r612 59 61 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.66 $Y=1.3
+ $X2=2.66 $Y2=0.74
r613 55 235 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.355 $Y=1.63
+ $X2=2.355 $Y2=1.465
r614 55 57 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=2.355 $Y=1.63
+ $X2=2.355 $Y2=2.4
r615 51 234 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.3
+ $X2=2.23 $Y2=1.465
r616 51 53 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.23 $Y=1.3
+ $X2=2.23 $Y2=0.74
r617 47 230 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.63
+ $X2=1.855 $Y2=1.465
r618 47 49 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.855 $Y=1.63
+ $X2=1.855 $Y2=2.4
r619 43 229 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.8 $Y=1.3
+ $X2=1.8 $Y2=1.465
r620 43 45 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.8 $Y=1.3 $X2=1.8
+ $Y2=0.74
r621 39 228 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.63
+ $X2=1.405 $Y2=1.465
r622 39 41 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.405 $Y=1.63
+ $X2=1.405 $Y2=2.4
r623 35 227 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=1.3
+ $X2=1.37 $Y2=1.465
r624 35 37 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.37 $Y=1.3
+ $X2=1.37 $Y2=0.74
r625 31 223 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.63
+ $X2=0.955 $Y2=1.465
r626 31 33 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.955 $Y=1.63
+ $X2=0.955 $Y2=2.4
r627 27 222 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.94 $Y=1.3
+ $X2=0.94 $Y2=1.465
r628 27 29 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.94 $Y=1.3
+ $X2=0.94 $Y2=0.74
r629 23 221 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.3
+ $X2=0.51 $Y2=1.465
r630 23 25 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.51 $Y=1.3
+ $X2=0.51 $Y2=0.74
r631 19 219 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=1.465
r632 19 21 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=2.4
r633 6 192 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=9.695
+ $Y=1.84 $X2=9.83 $Y2=2.115
r634 6 177 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.695
+ $Y=1.84 $X2=9.83 $Y2=2.815
r635 5 189 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=8.795
+ $Y=1.84 $X2=8.93 $Y2=2.115
r636 5 165 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.795
+ $Y=1.84 $X2=8.93 $Y2=2.815
r637 4 186 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=7.895
+ $Y=1.84 $X2=8.03 $Y2=2.115
r638 4 153 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.895
+ $Y=1.84 $X2=8.03 $Y2=2.815
r639 3 181 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.64
+ $Y=0.37 $X2=9.78 $Y2=0.515
r640 2 169 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.745
+ $Y=0.37 $X2=8.885 $Y2=0.515
r641 1 157 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.885
+ $Y=0.37 $X2=8.025 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__BUF_16%A 3 7 11 15 19 23 27 31 35 39 43 47 49 50 51
+ 52 53 77
c123 77 0 1.32147e-19 $X=10.065 $Y=1.515
c124 3 0 1.44668e-19 $X=7.805 $Y=2.4
r125 76 77 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=10.055 $Y=1.515
+ $X2=10.065 $Y2=1.515
r126 74 76 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.98 $Y=1.515
+ $X2=10.055 $Y2=1.515
r127 74 75 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=9.98
+ $Y=1.515 $X2=9.98 $Y2=1.515
r128 72 74 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=9.605 $Y=1.515
+ $X2=9.98 $Y2=1.515
r129 71 72 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=9.565 $Y=1.515
+ $X2=9.605 $Y2=1.515
r130 70 71 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=9.155 $Y=1.515
+ $X2=9.565 $Y2=1.515
r131 69 70 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=9.1 $Y=1.515
+ $X2=9.155 $Y2=1.515
r132 68 69 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=8.705 $Y=1.515
+ $X2=9.1 $Y2=1.515
r133 67 68 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=8.67 $Y=1.515
+ $X2=8.705 $Y2=1.515
r134 66 67 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=8.255 $Y=1.515
+ $X2=8.67 $Y2=1.515
r135 65 66 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=8.24 $Y=1.515
+ $X2=8.255 $Y2=1.515
r136 63 65 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=7.94 $Y=1.515
+ $X2=8.24 $Y2=1.515
r137 63 64 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=7.94
+ $Y=1.515 $X2=7.94 $Y2=1.515
r138 61 63 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=7.81 $Y=1.515
+ $X2=7.94 $Y2=1.515
r139 59 61 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=7.805 $Y=1.515
+ $X2=7.81 $Y2=1.515
r140 53 75 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=10.32 $Y=1.565
+ $X2=9.98 $Y2=1.565
r141 52 75 3.75214 $w=4.28e-07 $l=1.4e-07 $layer=LI1_cond $X=9.84 $Y=1.565
+ $X2=9.98 $Y2=1.565
r142 51 52 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=9.36 $Y=1.565
+ $X2=9.84 $Y2=1.565
r143 50 51 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.565
+ $X2=9.36 $Y2=1.565
r144 49 50 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.4 $Y=1.565
+ $X2=8.88 $Y2=1.565
r145 49 64 12.3285 $w=4.28e-07 $l=4.6e-07 $layer=LI1_cond $X=8.4 $Y=1.565
+ $X2=7.94 $Y2=1.565
r146 45 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.065 $Y=1.35
+ $X2=10.065 $Y2=1.515
r147 45 47 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=10.065 $Y=1.35
+ $X2=10.065 $Y2=0.74
r148 41 76 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.055 $Y=1.68
+ $X2=10.055 $Y2=1.515
r149 41 43 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=10.055 $Y=1.68
+ $X2=10.055 $Y2=2.4
r150 37 72 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.605 $Y=1.68
+ $X2=9.605 $Y2=1.515
r151 37 39 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=9.605 $Y=1.68
+ $X2=9.605 $Y2=2.4
r152 33 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.565 $Y=1.35
+ $X2=9.565 $Y2=1.515
r153 33 35 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.565 $Y=1.35
+ $X2=9.565 $Y2=0.74
r154 29 70 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.155 $Y=1.68
+ $X2=9.155 $Y2=1.515
r155 29 31 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=9.155 $Y=1.68
+ $X2=9.155 $Y2=2.4
r156 25 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.1 $Y=1.35
+ $X2=9.1 $Y2=1.515
r157 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.1 $Y=1.35 $X2=9.1
+ $Y2=0.74
r158 21 68 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.705 $Y=1.68
+ $X2=8.705 $Y2=1.515
r159 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.705 $Y=1.68
+ $X2=8.705 $Y2=2.4
r160 17 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.67 $Y=1.35
+ $X2=8.67 $Y2=1.515
r161 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.67 $Y=1.35
+ $X2=8.67 $Y2=0.74
r162 13 66 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.255 $Y=1.68
+ $X2=8.255 $Y2=1.515
r163 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.255 $Y=1.68
+ $X2=8.255 $Y2=2.4
r164 9 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.24 $Y=1.35
+ $X2=8.24 $Y2=1.515
r165 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.24 $Y=1.35
+ $X2=8.24 $Y2=0.74
r166 5 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.81 $Y=1.35
+ $X2=7.81 $Y2=1.515
r167 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.81 $Y=1.35 $X2=7.81
+ $Y2=0.74
r168 1 59 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.805 $Y=1.68
+ $X2=7.805 $Y2=1.515
r169 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.805 $Y=1.68
+ $X2=7.805 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__BUF_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 37 39 45 51
+ 57 63 69 75 81 87 89 93 95 99 101 103 108 109 111 112 114 115 117 118 120 121
+ 123 124 126 127 128 129 130 157 166 169 173
c189 87 0 1.92956e-20 $X=7.53 $Y=2.455
c190 81 0 1.71822e-19 $X=6.63 $Y=2.13
c191 75 0 1.71822e-19 $X=5.73 $Y=2.13
c192 63 0 1.71822e-19 $X=3.93 $Y=2.13
c193 57 0 1.71822e-19 $X=3.03 $Y=2.13
c194 45 0 1.71822e-19 $X=1.18 $Y=2.13
r195 172 173 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r196 169 170 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r197 167 170 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r198 166 167 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r199 163 164 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r200 161 173 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r201 161 170 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r202 160 161 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r203 158 169 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.465 $Y=3.33
+ $X2=9.38 $Y2=3.33
r204 158 160 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=9.465 $Y=3.33
+ $X2=9.84 $Y2=3.33
r205 157 172 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=10.195 $Y=3.33
+ $X2=10.377 $Y2=3.33
r206 157 160 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=10.195 $Y=3.33
+ $X2=9.84 $Y2=3.33
r207 156 167 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r208 155 156 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r209 153 156 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r210 152 153 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r211 150 153 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r212 149 150 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r213 146 147 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r214 144 147 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r215 143 144 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r216 141 144 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r217 140 141 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r218 138 141 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r219 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r220 135 138 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r221 135 164 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r222 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r223 132 163 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r224 132 134 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r225 130 150 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=5.52 $Y2=3.33
r226 130 147 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=4.56 $Y2=3.33
r227 128 155 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=7.445 $Y=3.33
+ $X2=7.44 $Y2=3.33
r228 128 129 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.445 $Y=3.33
+ $X2=7.57 $Y2=3.33
r229 126 152 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.545 $Y=3.33
+ $X2=6.48 $Y2=3.33
r230 126 127 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.545 $Y=3.33
+ $X2=6.63 $Y2=3.33
r231 125 155 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=6.715 $Y=3.33
+ $X2=7.44 $Y2=3.33
r232 125 127 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.715 $Y=3.33
+ $X2=6.63 $Y2=3.33
r233 123 149 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.645 $Y=3.33
+ $X2=5.52 $Y2=3.33
r234 123 124 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.645 $Y=3.33
+ $X2=5.73 $Y2=3.33
r235 122 152 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=5.815 $Y=3.33
+ $X2=6.48 $Y2=3.33
r236 122 124 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.815 $Y=3.33
+ $X2=5.73 $Y2=3.33
r237 120 146 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.745 $Y=3.33
+ $X2=4.56 $Y2=3.33
r238 120 121 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.745 $Y=3.33
+ $X2=4.83 $Y2=3.33
r239 119 149 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.915 $Y=3.33
+ $X2=5.52 $Y2=3.33
r240 119 121 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=3.33
+ $X2=4.83 $Y2=3.33
r241 117 143 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.845 $Y=3.33
+ $X2=3.6 $Y2=3.33
r242 117 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.845 $Y=3.33
+ $X2=3.93 $Y2=3.33
r243 116 146 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=4.015 $Y=3.33
+ $X2=4.56 $Y2=3.33
r244 116 118 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.015 $Y=3.33
+ $X2=3.93 $Y2=3.33
r245 114 140 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=2.64 $Y2=3.33
r246 114 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=3.03 $Y2=3.33
r247 113 143 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.115 $Y=3.33
+ $X2=3.6 $Y2=3.33
r248 113 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=3.33
+ $X2=3.03 $Y2=3.33
r249 111 137 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.965 $Y=3.33
+ $X2=1.68 $Y2=3.33
r250 111 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.965 $Y=3.33
+ $X2=2.09 $Y2=3.33
r251 110 140 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.64 $Y2=3.33
r252 110 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.09 $Y2=3.33
r253 108 134 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.72 $Y2=3.33
r254 108 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.18 $Y2=3.33
r255 107 137 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.68 $Y2=3.33
r256 107 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.18 $Y2=3.33
r257 103 106 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=10.32 $Y=2.115
+ $X2=10.32 $Y2=2.815
r258 101 172 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.32 $Y=3.245
+ $X2=10.377 $Y2=3.33
r259 101 106 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.32 $Y=3.245
+ $X2=10.32 $Y2=2.815
r260 97 169 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.38 $Y=3.245
+ $X2=9.38 $Y2=3.33
r261 97 99 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=9.38 $Y=3.245
+ $X2=9.38 $Y2=2.455
r262 96 166 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.565 $Y=3.33
+ $X2=8.48 $Y2=3.33
r263 95 169 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.295 $Y=3.33
+ $X2=9.38 $Y2=3.33
r264 95 96 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=9.295 $Y=3.33
+ $X2=8.565 $Y2=3.33
r265 91 166 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.48 $Y=3.245
+ $X2=8.48 $Y2=3.33
r266 91 93 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=8.48 $Y=3.245
+ $X2=8.48 $Y2=2.455
r267 90 129 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.695 $Y=3.33
+ $X2=7.57 $Y2=3.33
r268 89 166 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.395 $Y=3.33
+ $X2=8.48 $Y2=3.33
r269 89 90 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=8.395 $Y=3.33
+ $X2=7.695 $Y2=3.33
r270 85 129 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.57 $Y=3.245
+ $X2=7.57 $Y2=3.33
r271 85 87 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=7.57 $Y=3.245
+ $X2=7.57 $Y2=2.455
r272 81 84 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=6.63 $Y=2.13
+ $X2=6.63 $Y2=2.815
r273 79 127 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.63 $Y=3.245
+ $X2=6.63 $Y2=3.33
r274 79 84 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=6.63 $Y=3.245
+ $X2=6.63 $Y2=2.815
r275 75 78 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.73 $Y=2.13
+ $X2=5.73 $Y2=2.81
r276 73 124 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.73 $Y=3.245
+ $X2=5.73 $Y2=3.33
r277 73 78 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=5.73 $Y=3.245
+ $X2=5.73 $Y2=2.81
r278 69 72 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=4.83 $Y=2.13
+ $X2=4.83 $Y2=2.815
r279 67 121 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.83 $Y=3.245
+ $X2=4.83 $Y2=3.33
r280 67 72 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.83 $Y=3.245
+ $X2=4.83 $Y2=2.815
r281 63 66 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.93 $Y=2.13
+ $X2=3.93 $Y2=2.81
r282 61 118 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.93 $Y=3.245
+ $X2=3.93 $Y2=3.33
r283 61 66 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.93 $Y=3.245
+ $X2=3.93 $Y2=2.81
r284 57 60 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.03 $Y=2.13
+ $X2=3.03 $Y2=2.815
r285 55 115 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=3.245
+ $X2=3.03 $Y2=3.33
r286 55 60 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.03 $Y=3.245
+ $X2=3.03 $Y2=2.815
r287 51 54 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=2.09 $Y=2.13
+ $X2=2.09 $Y2=2.81
r288 49 112 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.09 $Y=3.245
+ $X2=2.09 $Y2=3.33
r289 49 54 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=2.09 $Y=3.245
+ $X2=2.09 $Y2=2.81
r290 45 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.18 $Y=2.13
+ $X2=1.18 $Y2=2.81
r291 43 109 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r292 43 48 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.81
r293 39 42 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r294 37 163 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r295 37 42 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r296 12 106 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.145
+ $Y=1.84 $X2=10.28 $Y2=2.815
r297 12 103 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=10.145
+ $Y=1.84 $X2=10.28 $Y2=2.115
r298 11 99 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=9.245
+ $Y=1.84 $X2=9.38 $Y2=2.455
r299 10 93 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=8.345
+ $Y=1.84 $X2=8.48 $Y2=2.455
r300 9 87 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=7.395
+ $Y=1.84 $X2=7.53 $Y2=2.455
r301 8 84 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.495
+ $Y=1.84 $X2=6.63 $Y2=2.815
r302 8 81 400 $w=1.7e-07 $l=3.5107e-07 $layer=licon1_PDIFF $count=1 $X=6.495
+ $Y=1.84 $X2=6.63 $Y2=2.13
r303 7 78 400 $w=1.7e-07 $l=1.0353e-06 $layer=licon1_PDIFF $count=1 $X=5.595
+ $Y=1.84 $X2=5.73 $Y2=2.81
r304 7 75 400 $w=1.7e-07 $l=3.5107e-07 $layer=licon1_PDIFF $count=1 $X=5.595
+ $Y=1.84 $X2=5.73 $Y2=2.13
r305 6 72 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.695
+ $Y=1.84 $X2=4.83 $Y2=2.815
r306 6 69 400 $w=1.7e-07 $l=3.5107e-07 $layer=licon1_PDIFF $count=1 $X=4.695
+ $Y=1.84 $X2=4.83 $Y2=2.13
r307 5 66 400 $w=1.7e-07 $l=1.0353e-06 $layer=licon1_PDIFF $count=1 $X=3.795
+ $Y=1.84 $X2=3.93 $Y2=2.81
r308 5 63 400 $w=1.7e-07 $l=3.5107e-07 $layer=licon1_PDIFF $count=1 $X=3.795
+ $Y=1.84 $X2=3.93 $Y2=2.13
r309 4 60 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.895
+ $Y=1.84 $X2=3.03 $Y2=2.815
r310 4 57 400 $w=1.7e-07 $l=3.5107e-07 $layer=licon1_PDIFF $count=1 $X=2.895
+ $Y=1.84 $X2=3.03 $Y2=2.13
r311 3 54 400 $w=1.7e-07 $l=1.05847e-06 $layer=licon1_PDIFF $count=1 $X=1.945
+ $Y=1.84 $X2=2.13 $Y2=2.81
r312 3 51 400 $w=1.7e-07 $l=3.71147e-07 $layer=licon1_PDIFF $count=1 $X=1.945
+ $Y=1.84 $X2=2.13 $Y2=2.13
r313 2 48 400 $w=1.7e-07 $l=1.0353e-06 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.81
r314 2 45 400 $w=1.7e-07 $l=3.5107e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.13
r315 1 42 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r316 1 39 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__BUF_16%X 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 51
+ 55 61 67 71 75 77 79 83 84 85 86 87 90 92 94 97 107 117 124 131 138 145 147
+ 152 153
c259 147 0 2.08474e-19 $X=7.11 $Y=2.035
c260 145 0 1.0264e-19 $X=7.08 $Y=1.985
c261 131 0 1.02687e-19 $X=5.28 $Y=1.985
c262 117 0 1.02631e-19 $X=2.58 $Y=1.985
r263 152 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.385 $Y=2.035
+ $X2=4.385 $Y2=2.035
r264 152 153 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.38 $Y=1.985
+ $X2=4.38 $Y2=1.9
r265 145 149 36.0954 $w=2.63e-07 $l=8.3e-07 $layer=LI1_cond $X=7.112 $Y=1.985
+ $X2=7.112 $Y2=2.815
r266 145 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.11 $Y=2.035
+ $X2=7.11 $Y2=2.035
r267 140 147 0.596692 $w=2.3e-07 $l=9.3e-07 $layer=MET1_cond $X=6.18 $Y=2.035
+ $X2=7.11 $Y2=2.035
r268 138 142 35.427 $w=2.68e-07 $l=8.3e-07 $layer=LI1_cond $X=6.195 $Y=1.985
+ $X2=6.195 $Y2=2.815
r269 138 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.18 $Y=2.035
+ $X2=6.18 $Y2=2.035
r270 133 140 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=5.28 $Y=2.035
+ $X2=6.18 $Y2=2.035
r271 133 155 0.574236 $w=2.3e-07 $l=8.95e-07 $layer=MET1_cond $X=5.28 $Y=2.035
+ $X2=4.385 $Y2=2.035
r272 131 135 32.4247 $w=2.93e-07 $l=8.3e-07 $layer=LI1_cond $X=5.262 $Y=1.985
+ $X2=5.262 $Y2=2.815
r273 131 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.28 $Y=2.035
+ $X2=5.28 $Y2=2.035
r274 124 128 37.5109 $w=2.53e-07 $l=8.3e-07 $layer=LI1_cond $X=3.437 $Y=1.985
+ $X2=3.437 $Y2=2.815
r275 124 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.445 $Y=2.035
+ $X2=3.445 $Y2=2.035
r276 119 126 0.571028 $w=2.3e-07 $l=8.9e-07 $layer=MET1_cond $X=2.555 $Y=2.035
+ $X2=3.445 $Y2=2.035
r277 117 121 36.7895 $w=2.58e-07 $l=8.3e-07 $layer=LI1_cond $X=2.545 $Y=1.985
+ $X2=2.545 $Y2=2.815
r278 117 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.555 $Y=2.035
+ $X2=2.555 $Y2=2.035
r279 112 119 0.612732 $w=2.3e-07 $l=9.55e-07 $layer=MET1_cond $X=1.6 $Y=2.035
+ $X2=2.555 $Y2=2.035
r280 110 114 37.5109 $w=2.53e-07 $l=8.3e-07 $layer=LI1_cond $X=1.592 $Y=1.985
+ $X2=1.592 $Y2=2.815
r281 110 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.6 $Y=2.035
+ $X2=1.6 $Y2=2.035
r282 107 110 66.435 $w=2.53e-07 $l=1.47e-06 $layer=LI1_cond $X=1.592 $Y=0.515
+ $X2=1.592 $Y2=1.985
r283 102 112 0.564612 $w=2.3e-07 $l=8.8e-07 $layer=MET1_cond $X=0.72 $Y=2.035
+ $X2=1.6 $Y2=2.035
r284 100 104 37.5109 $w=2.53e-07 $l=8.3e-07 $layer=LI1_cond $X=0.687 $Y=1.985
+ $X2=0.687 $Y2=2.815
r285 100 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=2.035
+ $X2=0.72 $Y2=2.035
r286 97 100 66.435 $w=2.53e-07 $l=1.47e-06 $layer=LI1_cond $X=0.687 $Y=0.515
+ $X2=0.687 $Y2=1.985
r287 94 155 0.301554 $w=2.3e-07 $l=4.7e-07 $layer=MET1_cond $X=3.915 $Y=2.035
+ $X2=4.385 $Y2=2.035
r288 94 126 0.301554 $w=2.3e-07 $l=4.7e-07 $layer=MET1_cond $X=3.915 $Y=2.035
+ $X2=3.445 $Y2=2.035
r289 93 145 26.2235 $w=2.63e-07 $l=6.03e-07 $layer=LI1_cond $X=7.112 $Y=1.382
+ $X2=7.112 $Y2=1.985
r290 92 138 36.494 $w=2.68e-07 $l=8.55e-07 $layer=LI1_cond $X=6.195 $Y=1.13
+ $X2=6.195 $Y2=1.985
r291 90 131 23.8302 $w=2.93e-07 $l=6.1e-07 $layer=LI1_cond $X=5.262 $Y=1.375
+ $X2=5.262 $Y2=1.985
r292 89 90 5.22441 $w=3.73e-07 $l=1.7e-07 $layer=LI1_cond $X=5.222 $Y=1.205
+ $X2=5.222 $Y2=1.375
r293 87 153 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.3 $Y=1.13
+ $X2=4.3 $Y2=1.9
r294 85 124 1.71737 $w=2.53e-07 $l=3.8e-08 $layer=LI1_cond $X=3.437 $Y=1.947
+ $X2=3.437 $Y2=1.985
r295 85 86 7.02311 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=3.437 $Y=1.947
+ $X2=3.437 $Y2=1.82
r296 84 86 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.395 $Y=1.13
+ $X2=3.395 $Y2=1.82
r297 83 117 27.9246 $w=2.58e-07 $l=6.3e-07 $layer=LI1_cond $X=2.545 $Y=1.355
+ $X2=2.545 $Y2=1.985
r298 82 83 7.39303 $w=2.63e-07 $l=1.7e-07 $layer=LI1_cond $X=2.51 $Y=1.185
+ $X2=2.51 $Y2=1.355
r299 77 93 12.2 $w=2.57e-07 $l=2.6342e-07 $layer=LI1_cond $X=7.125 $Y=1.125
+ $X2=7.112 $Y2=1.382
r300 77 79 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=7.125 $Y=1.125
+ $X2=7.125 $Y2=0.515
r301 73 92 6.17723 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.165 $Y=0.965
+ $X2=6.165 $Y2=1.13
r302 73 75 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=6.165 $Y=0.965
+ $X2=6.165 $Y2=0.515
r303 71 89 26.9554 $w=2.93e-07 $l=6.9e-07 $layer=LI1_cond $X=5.182 $Y=0.515
+ $X2=5.182 $Y2=1.205
r304 65 152 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.38 $Y=2.065
+ $X2=4.38 $Y2=1.985
r305 65 67 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=4.38 $Y=2.065
+ $X2=4.38 $Y2=2.815
r306 59 87 9.39714 $w=3.83e-07 $l=1.92e-07 $layer=LI1_cond $X=4.192 $Y=0.938
+ $X2=4.192 $Y2=1.13
r307 59 61 12.6619 $w=3.83e-07 $l=4.23e-07 $layer=LI1_cond $X=4.192 $Y=0.938
+ $X2=4.192 $Y2=0.515
r308 53 84 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=3.35 $Y=1 $X2=3.35
+ $Y2=1.13
r309 53 55 21.4975 $w=2.58e-07 $l=4.85e-07 $layer=LI1_cond $X=3.35 $Y=1 $X2=3.35
+ $Y2=0.515
r310 51 82 29.1372 $w=2.63e-07 $l=6.7e-07 $layer=LI1_cond $X=2.477 $Y=0.515
+ $X2=2.477 $Y2=1.185
r311 16 149 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.945
+ $Y=1.84 $X2=7.08 $Y2=2.815
r312 16 145 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.945
+ $Y=1.84 $X2=7.08 $Y2=1.985
r313 15 142 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.045
+ $Y=1.84 $X2=6.18 $Y2=2.815
r314 15 138 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.045
+ $Y=1.84 $X2=6.18 $Y2=1.985
r315 14 135 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.145
+ $Y=1.84 $X2=5.28 $Y2=2.815
r316 14 131 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.145
+ $Y=1.84 $X2=5.28 $Y2=1.985
r317 13 152 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.245
+ $Y=1.84 $X2=4.38 $Y2=1.985
r318 13 67 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.245
+ $Y=1.84 $X2=4.38 $Y2=2.815
r319 12 128 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.345
+ $Y=1.84 $X2=3.48 $Y2=2.815
r320 12 124 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.345
+ $Y=1.84 $X2=3.48 $Y2=1.985
r321 11 121 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.445
+ $Y=1.84 $X2=2.58 $Y2=2.815
r322 11 117 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.445
+ $Y=1.84 $X2=2.58 $Y2=1.985
r323 10 114 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.84 $X2=1.63 $Y2=2.815
r324 10 110 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.84 $X2=1.63 $Y2=1.985
r325 9 104 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.815
r326 9 100 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=1.985
r327 8 79 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.025
+ $Y=0.37 $X2=7.165 $Y2=0.515
r328 7 75 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.025
+ $Y=0.37 $X2=6.165 $Y2=0.515
r329 6 71 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.025
+ $Y=0.37 $X2=5.165 $Y2=0.515
r330 5 61 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.025
+ $Y=0.37 $X2=4.165 $Y2=0.515
r331 4 55 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.165
+ $Y=0.37 $X2=3.305 $Y2=0.515
r332 3 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.305
+ $Y=0.37 $X2=2.445 $Y2=0.515
r333 2 107 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.445
+ $Y=0.37 $X2=1.585 $Y2=0.515
r334 1 97 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.585
+ $Y=0.37 $X2=0.725 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__BUF_16%VGND 1 2 3 4 5 6 7 8 9 10 11 12 37 39 43 47
+ 51 55 57 61 63 67 71 73 77 81 85 87 89 92 93 95 96 97 98 99 100 101 103 122
+ 127 132 141 144 147 150 153 156 160
c185 89 0 1.32147e-19 $X=10.28 $Y=0.515
r186 159 160 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r187 156 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r188 153 154 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r189 150 151 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r190 147 148 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r191 144 145 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r192 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r193 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r194 136 160 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r195 136 157 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=9.36 $Y2=0
r196 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r197 133 156 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.48 $Y=0
+ $X2=9.315 $Y2=0
r198 133 135 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=9.48 $Y=0
+ $X2=9.84 $Y2=0
r199 132 159 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=10.337 $Y2=0
r200 132 135 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=9.84 $Y2=0
r201 131 157 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r202 131 154 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=8.4 $Y2=0
r203 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r204 128 153 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.62 $Y=0
+ $X2=8.455 $Y2=0
r205 128 130 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=8.62 $Y=0
+ $X2=8.88 $Y2=0
r206 127 156 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.15 $Y=0
+ $X2=9.315 $Y2=0
r207 127 130 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.15 $Y=0 $X2=8.88
+ $Y2=0
r208 126 154 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=8.4 $Y2=0
r209 126 151 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r210 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r211 123 150 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.76 $Y=0
+ $X2=7.595 $Y2=0
r212 123 125 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.76 $Y=0
+ $X2=7.92 $Y2=0
r213 122 153 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.29 $Y=0
+ $X2=8.455 $Y2=0
r214 122 125 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=8.29 $Y=0 $X2=7.92
+ $Y2=0
r215 121 151 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=7.44 $Y2=0
r216 121 148 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=5.52 $Y2=0
r217 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r218 118 147 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.83 $Y=0
+ $X2=5.665 $Y2=0
r219 118 120 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.83 $Y=0
+ $X2=6.48 $Y2=0
r220 117 145 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0
+ $X2=4.56 $Y2=0
r221 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r222 114 117 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.6 $Y2=0
r223 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r224 111 114 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.64 $Y2=0
r225 111 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=1.2 $Y2=0
r226 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r227 108 141 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=1.285 $Y=0
+ $X2=1.137 $Y2=0
r228 108 110 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.285 $Y=0
+ $X2=1.68 $Y2=0
r229 107 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=1.2 $Y2=0
r230 107 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r231 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r232 104 138 3.99177 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.38 $Y=0 $X2=0.19
+ $Y2=0
r233 104 106 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.38 $Y=0
+ $X2=0.72 $Y2=0
r234 103 141 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.99 $Y=0
+ $X2=1.137 $Y2=0
r235 103 106 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.72
+ $Y2=0
r236 101 148 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=5.52 $Y2=0
r237 101 145 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=4.56 $Y2=0
r238 99 120 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=6.5 $Y=0 $X2=6.48
+ $Y2=0
r239 99 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.5 $Y=0 $X2=6.665
+ $Y2=0
r240 97 116 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=3.65 $Y=0 $X2=3.6
+ $Y2=0
r241 97 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.65 $Y=0 $X2=3.735
+ $Y2=0
r242 95 113 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.79 $Y=0 $X2=2.64
+ $Y2=0
r243 95 96 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.79 $Y=0 $X2=2.875
+ $Y2=0
r244 94 116 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.96 $Y=0 $X2=3.6
+ $Y2=0
r245 94 96 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.96 $Y=0 $X2=2.875
+ $Y2=0
r246 92 110 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.895 $Y=0
+ $X2=1.68 $Y2=0
r247 92 93 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=1.895 $Y=0
+ $X2=1.997 $Y2=0
r248 91 113 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.1 $Y=0 $X2=2.64
+ $Y2=0
r249 91 93 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=2.1 $Y=0 $X2=1.997
+ $Y2=0
r250 87 159 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.28 $Y=0.085
+ $X2=10.337 $Y2=0
r251 87 89 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.28 $Y=0.085
+ $X2=10.28 $Y2=0.515
r252 83 156 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.315 $Y=0.085
+ $X2=9.315 $Y2=0
r253 83 85 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=9.315 $Y=0.085
+ $X2=9.315 $Y2=0.675
r254 79 153 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.455 $Y=0.085
+ $X2=8.455 $Y2=0
r255 79 81 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=8.455 $Y=0.085
+ $X2=8.455 $Y2=0.675
r256 75 150 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.595 $Y=0.085
+ $X2=7.595 $Y2=0
r257 75 77 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=7.595 $Y=0.085
+ $X2=7.595 $Y2=0.675
r258 74 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.83 $Y=0
+ $X2=6.665 $Y2=0
r259 73 150 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.43 $Y=0
+ $X2=7.595 $Y2=0
r260 73 74 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.43 $Y=0 $X2=6.83
+ $Y2=0
r261 69 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.665 $Y=0.085
+ $X2=6.665 $Y2=0
r262 69 71 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.665 $Y=0.085
+ $X2=6.665 $Y2=0.495
r263 65 147 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.665 $Y=0.085
+ $X2=5.665 $Y2=0
r264 65 67 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=5.665 $Y=0.085
+ $X2=5.665 $Y2=0.495
r265 64 144 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=4.83 $Y=0
+ $X2=4.692 $Y2=0
r266 63 147 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.5 $Y=0 $X2=5.665
+ $Y2=0
r267 63 64 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.5 $Y=0 $X2=4.83
+ $Y2=0
r268 59 144 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=4.692 $Y=0.085
+ $X2=4.692 $Y2=0
r269 59 61 17.1819 $w=2.73e-07 $l=4.1e-07 $layer=LI1_cond $X=4.692 $Y=0.085
+ $X2=4.692 $Y2=0.495
r270 58 98 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.82 $Y=0 $X2=3.735
+ $Y2=0
r271 57 144 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=4.555 $Y=0
+ $X2=4.692 $Y2=0
r272 57 58 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=4.555 $Y=0
+ $X2=3.82 $Y2=0
r273 53 98 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.735 $Y=0.085
+ $X2=3.735 $Y2=0
r274 53 55 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.735 $Y=0.085
+ $X2=3.735 $Y2=0.495
r275 49 96 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.875 $Y=0.085
+ $X2=2.875 $Y2=0
r276 49 51 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.875 $Y=0.085
+ $X2=2.875 $Y2=0.495
r277 45 93 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.997 $Y=0.085
+ $X2=1.997 $Y2=0
r278 45 47 22.1818 $w=2.03e-07 $l=4.1e-07 $layer=LI1_cond $X=1.997 $Y=0.085
+ $X2=1.997 $Y2=0.495
r279 41 141 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.137 $Y=0.085
+ $X2=1.137 $Y2=0
r280 41 43 16.017 $w=2.93e-07 $l=4.1e-07 $layer=LI1_cond $X=1.137 $Y=0.085
+ $X2=1.137 $Y2=0.495
r281 37 138 3.1514 $w=2.5e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.19 $Y2=0
r282 37 39 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.255 $Y2=0.515
r283 12 89 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.14
+ $Y=0.37 $X2=10.28 $Y2=0.515
r284 11 85 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=9.175
+ $Y=0.37 $X2=9.315 $Y2=0.675
r285 10 81 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=8.315
+ $Y=0.37 $X2=8.455 $Y2=0.675
r286 9 77 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=7.455
+ $Y=0.37 $X2=7.595 $Y2=0.675
r287 8 71 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=6.455
+ $Y=0.37 $X2=6.665 $Y2=0.495
r288 7 67 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=5.455
+ $Y=0.37 $X2=5.665 $Y2=0.495
r289 6 61 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=4.455
+ $Y=0.37 $X2=4.665 $Y2=0.495
r290 5 55 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.595
+ $Y=0.37 $X2=3.735 $Y2=0.495
r291 4 51 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.735
+ $Y=0.37 $X2=2.875 $Y2=0.495
r292 3 47 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.875
+ $Y=0.37 $X2=2.015 $Y2=0.495
r293 2 43 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.015
+ $Y=0.37 $X2=1.155 $Y2=0.495
r294 1 39 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.37 $X2=0.295 $Y2=0.515
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_ms__dlclkp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__dlclkp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN GATE
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.470000 1.335000 1.800000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.524500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.205000 1.550000 6.605000 2.980000 ;
        RECT 6.275000 0.350000 6.605000 1.550000 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.509400 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.475000 5.155000 1.805000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 6.720000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 2.670000 1.785000 ;
        RECT -0.190000 1.785000 6.910000 3.520000 ;
        RECT  5.035000 1.660000 6.910000 1.785000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.095000  0.350000 0.445000 0.790000 ;
      RECT 0.095000  0.790000 1.215000 0.960000 ;
      RECT 0.095000  0.960000 0.445000 1.130000 ;
      RECT 0.095000  1.130000 0.265000 1.820000 ;
      RECT 0.095000  1.820000 0.445000 2.980000 ;
      RECT 0.435000  1.300000 0.785000 1.630000 ;
      RECT 0.615000  1.130000 1.555000 1.300000 ;
      RECT 0.615000  1.630000 0.785000 1.970000 ;
      RECT 0.615000  1.970000 1.555000 2.140000 ;
      RECT 0.615000  2.310000 0.945000 3.245000 ;
      RECT 0.625000  0.085000 0.875000 0.620000 ;
      RECT 1.045000  0.255000 2.955000 0.425000 ;
      RECT 1.045000  0.425000 1.215000 0.790000 ;
      RECT 1.385000  0.650000 2.260000 0.980000 ;
      RECT 1.385000  0.980000 1.555000 1.130000 ;
      RECT 1.385000  2.140000 1.555000 2.550000 ;
      RECT 1.385000  2.550000 2.285000 2.880000 ;
      RECT 1.725000  1.150000 1.995000 2.050000 ;
      RECT 1.725000  2.050000 3.200000 2.380000 ;
      RECT 2.205000  1.160000 3.775000 1.330000 ;
      RECT 2.205000  1.330000 2.535000 1.840000 ;
      RECT 2.625000  0.425000 2.955000 0.510000 ;
      RECT 2.750000  0.685000 3.295000 0.935000 ;
      RECT 2.835000  2.730000 3.165000 3.245000 ;
      RECT 3.030000  1.500000 3.435000 1.830000 ;
      RECT 3.030000  1.830000 3.200000 2.050000 ;
      RECT 3.030000  2.380000 3.200000 2.390000 ;
      RECT 3.030000  2.390000 4.260000 2.560000 ;
      RECT 3.125000  0.085000 3.295000 0.685000 ;
      RECT 3.370000  2.050000 3.775000 2.220000 ;
      RECT 3.465000  0.605000 3.775000 1.160000 ;
      RECT 3.605000  1.330000 3.775000 2.050000 ;
      RECT 3.945000  1.055000 4.205000 1.945000 ;
      RECT 3.945000  1.945000 4.260000 2.390000 ;
      RECT 3.945000  2.560000 4.260000 2.825000 ;
      RECT 4.385000  0.085000 4.715000 1.305000 ;
      RECT 4.430000  1.975000 4.760000 3.245000 ;
      RECT 4.930000  1.975000 5.535000 2.145000 ;
      RECT 4.930000  2.145000 5.260000 2.825000 ;
      RECT 5.285000  0.605000 5.615000 1.285000 ;
      RECT 5.365000  1.285000 5.615000 1.300000 ;
      RECT 5.365000  1.300000 6.035000 1.630000 ;
      RECT 5.365000  1.630000 5.535000 1.975000 ;
      RECT 5.705000  1.945000 6.035000 3.245000 ;
      RECT 5.845000  0.085000 6.095000 1.130000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_ms__dlclkp_1
END LIBRARY

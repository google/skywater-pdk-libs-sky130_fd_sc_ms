* File: sky130_fd_sc_ms__a21boi_2.spice
* Created: Fri Aug 28 16:58:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a21boi_2.pex.spice"
.subckt sky130_fd_sc_ms__a21boi_2  VNB VPB B1_N A1 A2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2	A2
* A1	A1
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_B1_N_M1003_g N_A_62_94#_M1003_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.113206 AS=0.1696 PD=1.00174 PS=1.81 NRD=11.712 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1006 N_Y_M1006_d N_A_62_94#_M1006_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.130894 PD=1.02 PS=1.15826 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1011 N_Y_M1006_d N_A_62_94#_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_436_74#_M1000_d N_A1_M1000_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1012 N_A_436_74#_M1012_d N_A1_M1012_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g N_A_436_74#_M1012_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1007_d N_A2_M1013_g N_A_436_74#_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_A_62_94#_M1010_d N_B1_N_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.18 W=1
+ AD=0.26 AS=0.26 PD=2.52 PS=2.52 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1001 N_Y_M1001_d N_A_62_94#_M1001_g N_A_241_368#_M1001_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1002 N_Y_M1001_d N_A_62_94#_M1002_g N_A_241_368#_M1002_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90002 A=0.2016 P=2.6 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g N_A_241_368#_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1005 N_VPWR_M1004_d N_A1_M1005_g N_A_241_368#_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1008 N_VPWR_M1008_d N_A2_M1008_g N_A_241_368#_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1624 AS=0.1512 PD=1.41 PS=1.39 NRD=0.8668 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1009 N_VPWR_M1008_d N_A2_M1009_g N_A_241_368#_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1624 AS=0.2912 PD=1.41 PS=2.76 NRD=0.8668 NRS=0 M=1 R=6.22222 SA=90002.4
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.742 P=13.12
c_48 VNB 0 1.97879e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__a21boi_2.pxi.spice"
*
.ends
*
*

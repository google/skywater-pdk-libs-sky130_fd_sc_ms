* File: sky130_fd_sc_ms__o211ai_1.spice
* Created: Fri Aug 28 17:53:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o211ai_1.pex.spice"
.subckt sky130_fd_sc_ms__o211ai_1  VNB VPB A1 A2 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A1_M1006_g N_A_31_74#_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1000 N_A_31_74#_M1000_d N_A2_M1000_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.11655 AS=0.1295 PD=1.055 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1001 A_311_74# N_B1_M1001_g N_A_31_74#_M1000_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.11655 PD=1.16 PS=1.055 NRD=25.128 NRS=5.664 M=1 R=4.93333
+ SA=75001.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1007 N_Y_M1007_d N_C1_M1007_g A_311_74# VNB NLOWVT L=0.15 W=0.74 AD=0.4588
+ AS=0.1554 PD=2.72 PS=1.16 NRD=0 NRS=25.128 M=1 R=4.93333 SA=75001.7 SB=75000.5
+ A=0.111 P=1.78 MULT=1
MM1004 A_119_368# N_A1_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12 AD=0.1344
+ AS=0.3136 PD=1.36 PS=2.8 NRD=11.426 NRS=0 M=1 R=6.22222 SA=90000.2 SB=90001.8
+ A=0.2016 P=2.6 MULT=1
MM1005 N_Y_M1005_d N_A2_M1005_g A_119_368# VPB PSHORT L=0.18 W=1.12 AD=0.3024
+ AS=0.1344 PD=1.66 PS=1.36 NRD=23.7385 NRS=11.426 M=1 R=6.22222 SA=90000.6
+ SB=90001.4 A=0.2016 P=2.6 MULT=1
MM1003 N_VPWR_M1003_d N_B1_M1003_g N_Y_M1005_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.3024 PD=1.44 PS=1.66 NRD=0 NRS=21.9852 M=1 R=6.22222 SA=90001.3
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1002 N_Y_M1002_d N_C1_M1002_g N_VPWR_M1003_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1792 PD=2.8 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.8
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ms__o211ai_1.pxi.spice"
*
.ends
*
*

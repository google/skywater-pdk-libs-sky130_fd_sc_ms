* File: sky130_fd_sc_ms__sdfrbp_1.pex.spice
* Created: Fri Aug 28 18:11:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SDFRBP_1%A_27_74# 1 2 7 9 12 16 19 22 23 25 27 32 34
+ 35
c79 35 0 1.29655e-19 $X=2.5 $Y=1.995
c80 25 0 2.59912e-20 $X=2.365 $Y=2.135
r81 35 43 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.5 $Y=1.995
+ $X2=2.5 $Y2=2.16
r82 34 37 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=2.53 $Y=1.995
+ $X2=2.53 $Y2=2.135
r83 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.5
+ $Y=1.995 $X2=2.5 $Y2=1.995
r84 31 32 12.4206 $w=9.23e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=2.512
+ $X2=1.055 $Y2=2.512
r85 25 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=2.135
+ $X2=2.53 $Y2=2.135
r86 25 32 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=2.365 $Y=2.135
+ $X2=1.055 $Y2=2.135
r87 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.23
+ $Y=1.145 $X2=1.23 $Y2=1.145
r88 20 27 0.221902 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=1.145
+ $X2=0.24 $Y2=1.145
r89 20 22 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=0.365 $Y=1.145
+ $X2=1.23 $Y2=1.145
r90 19 31 9.10054 $w=9.23e-07 $l=6.9e-07 $layer=LI1_cond $X=0.2 $Y=2.512
+ $X2=0.89 $Y2=2.512
r91 18 27 7.38875 $w=2.1e-07 $l=1.83916e-07 $layer=LI1_cond $X=0.2 $Y=1.31
+ $X2=0.24 $Y2=1.145
r92 18 19 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.2 $Y=1.31 $X2=0.2
+ $Y2=2.05
r93 14 27 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=0.98
+ $X2=0.24 $Y2=1.145
r94 14 16 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=0.24 $Y=0.98 $X2=0.24
+ $Y2=0.58
r95 12 43 186.581 $w=1.8e-07 $l=4.8e-07 $layer=POLY_cond $X=2.485 $Y=2.64
+ $X2=2.485 $Y2=2.16
r96 7 23 45.5222 $w=2.7e-07 $l=3.27261e-07 $layer=POLY_cond $X=1.485 $Y=0.98
+ $X2=1.23 $Y2=1.145
r97 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.485 $Y=0.98
+ $X2=1.485 $Y2=0.66
r98 2 31 150 $w=1.7e-07 $l=8.24318e-07 $layer=licon1_PDIFF $count=4 $X=0.135
+ $Y=2.32 $X2=0.89 $Y2=2.465
r99 1 16 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_1%SCE 3 7 11 17 18 19 20 21 24 25 29 30 31 36
+ 44 47 49 58 60
c87 25 0 3.50849e-19 $X=2.5 $Y=1.425
c88 20 0 1.87424e-19 $X=2.62 $Y=1.105
r89 49 58 2.36399 $w=3.88e-07 $l=8e-08 $layer=LI1_cond $X=1.6 $Y=1.685 $X2=1.68
+ $Y2=1.685
r90 42 44 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.45 $Y=1.715
+ $X2=1.615 $Y2=1.715
r91 42 43 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.45
+ $Y=1.715 $X2=1.45 $Y2=1.715
r92 40 42 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=1.115 $Y=1.715
+ $X2=1.45 $Y2=1.715
r93 36 40 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.025 $Y=1.715
+ $X2=1.115 $Y2=1.715
r94 36 38 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=1.025 $Y=1.715
+ $X2=0.77 $Y2=1.715
r95 31 60 7.07103 $w=3.88e-07 $l=1.13e-07 $layer=LI1_cond $X=1.682 $Y=1.685
+ $X2=1.795 $Y2=1.685
r96 31 58 0.0590996 $w=3.88e-07 $l=2e-09 $layer=LI1_cond $X=1.682 $Y=1.685
+ $X2=1.68 $Y2=1.685
r97 31 49 0.0886495 $w=3.88e-07 $l=3e-09 $layer=LI1_cond $X=1.597 $Y=1.685
+ $X2=1.6 $Y2=1.685
r98 31 43 4.34382 $w=3.88e-07 $l=1.47e-07 $layer=LI1_cond $X=1.597 $Y=1.685
+ $X2=1.45 $Y2=1.685
r99 30 43 7.38745 $w=3.88e-07 $l=2.5e-07 $layer=LI1_cond $X=1.2 $Y=1.685
+ $X2=1.45 $Y2=1.685
r100 29 30 14.1839 $w=3.88e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.685
+ $X2=1.2 $Y2=1.685
r101 29 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.77
+ $Y=1.715 $X2=0.77 $Y2=1.715
r102 25 47 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.5 $Y=1.425
+ $X2=2.5 $Y2=1.26
r103 24 27 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.56 $Y=1.425
+ $X2=2.56 $Y2=1.575
r104 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.5
+ $Y=1.425 $X2=2.5 $Y2=1.425
r105 21 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=1.575
+ $X2=2.56 $Y2=1.575
r106 21 60 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.395 $Y=1.575
+ $X2=1.795 $Y2=1.575
r107 20 47 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=2.59 $Y=1.105
+ $X2=2.59 $Y2=1.26
r108 19 20 39.4735 $w=2.1e-07 $l=1.25e-07 $layer=POLY_cond $X=2.62 $Y=0.98
+ $X2=2.62 $Y2=1.105
r109 18 38 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.57 $Y=1.715
+ $X2=0.77 $Y2=1.715
r110 17 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.65 $Y=0.695
+ $X2=2.65 $Y2=0.98
r111 9 44 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.615 $Y=1.88
+ $X2=1.615 $Y2=1.715
r112 9 11 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=1.615 $Y=1.88
+ $X2=1.615 $Y2=2.64
r113 5 40 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.115 $Y=1.88
+ $X2=1.115 $Y2=1.715
r114 5 7 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=1.115 $Y=1.88
+ $X2=1.115 $Y2=2.64
r115 1 18 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.495 $Y=1.55
+ $X2=0.57 $Y2=1.715
r116 1 3 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=0.495 $Y=1.55
+ $X2=0.495 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_1%D 3 6 8 11 12 13
c41 12 0 1.71349e-19 $X=1.935 $Y=1.145
r42 11 14 40.8147 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.947 $Y=1.145
+ $X2=1.947 $Y2=1.31
r43 11 13 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.947 $Y=1.145
+ $X2=1.947 $Y2=0.98
r44 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.145 $X2=1.935 $Y2=1.145
r45 8 12 6.1 $w=4.98e-07 $l=2.55e-07 $layer=LI1_cond $X=1.68 $Y=1.06 $X2=1.935
+ $Y2=1.06
r46 6 14 516.984 $w=1.8e-07 $l=1.33e-06 $layer=POLY_cond $X=2.035 $Y=2.64
+ $X2=2.035 $Y2=1.31
r47 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.99 $Y=0.66 $X2=1.99
+ $Y2=0.98
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_1%SCD 1 3 5 7 9 10 11
c43 10 0 2.86215e-19 $X=3.12 $Y=1.665
c44 5 0 7.88209e-20 $X=3.025 $Y=2.245
c45 3 0 3.39925e-20 $X=3.01 $Y=0.695
r46 10 11 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.1 $Y=1.605 $X2=3.1
+ $Y2=2.035
r47 10 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.04
+ $Y=1.605 $X2=3.04 $Y2=1.605
r48 9 15 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.04 $Y=1.945
+ $X2=3.04 $Y2=1.605
r49 5 9 50.0346 $w=2.89e-07 $l=3.07409e-07 $layer=POLY_cond $X=3.025 $Y=2.245
+ $X2=3.04 $Y2=1.945
r50 5 7 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.025 $Y=2.245
+ $X2=3.025 $Y2=2.64
r51 1 15 63.4211 $w=2.66e-07 $l=3.64692e-07 $layer=POLY_cond $X=3.01 $Y=1.255
+ $X2=3.04 $Y2=1.605
r52 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.01 $Y=1.255 $X2=3.01
+ $Y2=0.695
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_1%CLK 1 5 8 12 14 16 19 24 25
c61 24 0 3.36092e-20 $X=4.565 $Y=1.51
c62 12 0 1.67878e-19 $X=4.56 $Y=1.61
r63 24 25 35.2748 $w=3.4e-07 $l=1e-07 $layer=POLY_cond $X=4.565 $Y=1.51
+ $X2=4.565 $Y2=1.41
r64 19 22 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=3.94 $Y=1.445
+ $X2=3.94 $Y2=1.51
r65 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.94
+ $Y=1.445 $X2=3.94 $Y2=1.445
r66 16 20 3.56279 $w=4.68e-07 $l=1.4e-07 $layer=LI1_cond $X=4.08 $Y=1.415
+ $X2=3.94 $Y2=1.415
r67 14 16 8.01627 $w=4.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.395 $Y=1.415
+ $X2=4.08 $Y2=1.415
r68 13 27 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=4.565 $Y=1.61
+ $X2=4.565 $Y2=1.775
r69 13 24 16.9718 $w=3.4e-07 $l=1e-07 $layer=POLY_cond $X=4.565 $Y=1.61
+ $X2=4.565 $Y2=1.51
r70 12 14 3.87822 $w=5.93e-07 $l=1.65e-07 $layer=LI1_cond $X=4.56 $Y=1.477
+ $X2=4.395 $Y2=1.477
r71 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.56
+ $Y=1.61 $X2=4.56 $Y2=1.61
r72 8 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.645 $Y=2.495
+ $X2=4.645 $Y2=1.775
r73 5 25 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.54 $Y=0.965
+ $X2=4.54 $Y2=1.41
r74 2 22 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.105 $Y=1.51 $X2=3.94
+ $Y2=1.51
r75 1 24 15.178 $w=2e-07 $l=1.7e-07 $layer=POLY_cond $X=4.395 $Y=1.51 $X2=4.565
+ $Y2=1.51
r76 1 2 96.1574 $w=2e-07 $l=2.9e-07 $layer=POLY_cond $X=4.395 $Y=1.51 $X2=4.105
+ $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_1%A_1037_119# 1 2 9 11 15 17 19 20 21 24 29
+ 30 31 32 33 36 40 41 42 44 45 46 48 50 53 56 66 67 71 73 83
c211 67 0 1.52128e-19 $X=9.27 $Y=1.07
c212 66 0 1.89691e-19 $X=9.27 $Y=1.07
c213 31 0 1.32475e-19 $X=5.502 $Y=1.575
c214 29 0 1.7726e-19 $X=5.32 $Y=0.74
c215 15 0 1.92441e-20 $X=6.53 $Y=0.805
r216 67 79 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.27 $Y=1.07 $X2=9.27
+ $Y2=1.16
r217 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.27
+ $Y=1.07 $X2=9.27 $Y2=1.07
r218 63 66 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=8.865 $Y=0.99
+ $X2=9.27 $Y2=0.99
r219 56 58 13.1603 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=5.387 $Y=1.74
+ $X2=5.387 $Y2=2.11
r220 54 83 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=9.67 $Y=2.065
+ $X2=9.77 $Y2=2.065
r221 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.67
+ $Y=2.065 $X2=9.67 $Y2=2.065
r222 51 71 0.201461 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=9.63 $Y=1.575
+ $X2=9.63 $Y2=1.46
r223 51 53 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=9.63 $Y=1.575
+ $X2=9.63 $Y2=2.065
r224 50 71 18.0382 $w=2.28e-07 $l=3.6e-07 $layer=LI1_cond $X=9.27 $Y=1.46
+ $X2=9.63 $Y2=1.46
r225 50 66 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=9.27 $Y=1.345
+ $X2=9.27 $Y2=1.075
r226 48 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.865 $Y=0.905
+ $X2=8.865 $Y2=0.99
r227 47 48 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=8.865 $Y=0.425
+ $X2=8.865 $Y2=0.905
r228 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.78 $Y=0.34
+ $X2=8.865 $Y2=0.425
r229 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.78 $Y=0.34
+ $X2=8.11 $Y2=0.34
r230 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.025 $Y=0.425
+ $X2=8.11 $Y2=0.34
r231 43 44 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.025 $Y=0.425
+ $X2=8.025 $Y2=0.595
r232 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.94 $Y=0.68
+ $X2=8.025 $Y2=0.595
r233 41 42 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=7.94 $Y=0.68
+ $X2=7.185 $Y2=0.68
r234 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.1 $Y=0.595
+ $X2=7.185 $Y2=0.68
r235 39 40 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.1 $Y=0.425
+ $X2=7.1 $Y2=0.595
r236 37 76 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.055 $Y=1.74
+ $X2=6.055 $Y2=1.905
r237 37 73 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.055 $Y=1.74
+ $X2=6.055 $Y2=1.65
r238 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.055
+ $Y=1.74 $X2=6.055 $Y2=1.74
r239 34 56 0.950996 $w=3.3e-07 $l=2.33e-07 $layer=LI1_cond $X=5.62 $Y=1.74
+ $X2=5.387 $Y2=1.74
r240 34 36 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=5.62 $Y=1.74
+ $X2=6.055 $Y2=1.74
r241 32 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.015 $Y=0.34
+ $X2=7.1 $Y2=0.425
r242 32 33 104.059 $w=1.68e-07 $l=1.595e-06 $layer=LI1_cond $X=7.015 $Y=0.34
+ $X2=5.42 $Y2=0.34
r243 31 56 7.08745 $w=3.43e-07 $l=2.14942e-07 $layer=LI1_cond $X=5.502 $Y=1.575
+ $X2=5.387 $Y2=1.74
r244 30 31 14.712 $w=2.33e-07 $l=3e-07 $layer=LI1_cond $X=5.502 $Y=1.275
+ $X2=5.502 $Y2=1.575
r245 27 30 13.5048 $w=1.68e-07 $l=2.07e-07 $layer=LI1_cond $X=5.295 $Y=1.19
+ $X2=5.502 $Y2=1.19
r246 27 29 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=5.295 $Y=1.105
+ $X2=5.295 $Y2=0.74
r247 26 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.295 $Y=0.425
+ $X2=5.42 $Y2=0.34
r248 26 29 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=5.295 $Y=0.425
+ $X2=5.295 $Y2=0.74
r249 22 83 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.77 $Y=2.23
+ $X2=9.77 $Y2=2.065
r250 22 24 165.202 $w=1.8e-07 $l=4.25e-07 $layer=POLY_cond $X=9.77 $Y=2.23
+ $X2=9.77 $Y2=2.655
r251 20 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.105 $Y=1.16
+ $X2=9.27 $Y2=1.16
r252 20 21 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=9.105 $Y=1.16
+ $X2=8.735 $Y2=1.16
r253 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.66 $Y=1.085
+ $X2=8.735 $Y2=1.16
r254 17 19 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.66 $Y=1.085
+ $X2=8.66 $Y2=0.69
r255 13 15 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=6.53 $Y=1.575
+ $X2=6.53 $Y2=0.805
r256 12 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.22 $Y=1.65
+ $X2=6.055 $Y2=1.65
r257 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.455 $Y=1.65
+ $X2=6.53 $Y2=1.575
r258 11 12 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=6.455 $Y=1.65
+ $X2=6.22 $Y2=1.65
r259 9 76 241 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=6.115 $Y=2.525 $X2=6.115
+ $Y2=1.905
r260 2 58 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.185
+ $Y=1.935 $X2=5.32 $Y2=2.11
r261 1 29 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.185
+ $Y=0.595 $X2=5.32 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_1%A_1369_93# 1 2 9 13 17 18 20 21 24 27 28 30
+ 34
c101 34 0 1.32669e-19 $X=8.445 $Y=1.02
c102 28 0 4.00536e-20 $X=8.81 $Y=1.415
c103 24 0 1.94589e-20 $X=8.445 $Y=0.81
c104 21 0 1.11854e-19 $X=7.235 $Y=1.02
r105 39 41 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=6.92 $Y=1.615
+ $X2=6.955 $Y2=1.615
r106 30 32 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=8.81 $Y=1.88
+ $X2=8.81 $Y2=2.59
r107 28 35 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.81 $Y=1.33
+ $X2=8.525 $Y2=1.33
r108 28 30 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=8.81 $Y=1.415
+ $X2=8.81 $Y2=1.88
r109 27 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.525 $Y=1.245
+ $X2=8.525 $Y2=1.33
r110 26 34 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=8.525 $Y=1.105
+ $X2=8.445 $Y2=1.02
r111 26 27 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=8.525 $Y=1.105
+ $X2=8.525 $Y2=1.245
r112 22 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.445 $Y=0.935
+ $X2=8.445 $Y2=1.02
r113 22 24 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=8.445 $Y=0.935
+ $X2=8.445 $Y2=0.81
r114 20 34 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.28 $Y=1.02
+ $X2=8.445 $Y2=1.02
r115 20 21 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=8.28 $Y=1.02
+ $X2=7.235 $Y2=1.02
r116 18 41 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=7.125 $Y=1.615
+ $X2=6.955 $Y2=1.615
r117 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.125
+ $Y=1.615 $X2=7.125 $Y2=1.615
r118 15 21 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=7.125 $Y=1.105
+ $X2=7.235 $Y2=1.02
r119 15 17 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=7.125 $Y=1.105
+ $X2=7.125 $Y2=1.615
r120 11 41 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.955 $Y=1.78
+ $X2=6.955 $Y2=1.615
r121 11 13 289.589 $w=1.8e-07 $l=7.45e-07 $layer=POLY_cond $X=6.955 $Y=1.78
+ $X2=6.955 $Y2=2.525
r122 7 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.92 $Y=1.45
+ $X2=6.92 $Y2=1.615
r123 7 9 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=6.92 $Y=1.45
+ $X2=6.92 $Y2=0.805
r124 2 32 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.635
+ $Y=1.735 $X2=8.77 $Y2=2.59
r125 2 30 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.635
+ $Y=1.735 $X2=8.77 $Y2=1.88
r126 1 24 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=8.305
+ $Y=0.37 $X2=8.445 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_1%RESET_B 4 6 9 11 12 16 19 22 25 29 35 37 40
+ 43 46 48 49 50 51 52 53 61 64 65 68 69 72 73 74
c245 73 0 1.5378e-19 $X=10.9 $Y=1.845
c246 72 0 2.44776e-20 $X=10.9 $Y=1.845
c247 49 0 8.18368e-20 $X=10.81 $Y=2.37
c248 46 0 6.47027e-20 $X=10.81 $Y=1.335
c249 40 0 1.11854e-19 $X=7.605 $Y=1.165
c250 37 0 1.32707e-19 $X=3.415 $Y=1.82
r251 73 85 5.91795 $w=3.68e-07 $l=1.9e-07 $layer=LI1_cond $X=10.88 $Y=1.845
+ $X2=10.88 $Y2=2.035
r252 72 75 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.9 $Y=1.845
+ $X2=10.9 $Y2=2.01
r253 72 74 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.9 $Y=1.845
+ $X2=10.9 $Y2=1.68
r254 72 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.9
+ $Y=1.845 $X2=10.9 $Y2=1.845
r255 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.86
+ $Y=1.985 $X2=7.86 $Y2=1.985
r256 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.985 $X2=3.95 $Y2=1.985
r257 61 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=2.035
+ $X2=10.8 $Y2=2.035
r258 59 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r259 55 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=2.035
+ $X2=4.08 $Y2=2.035
r260 53 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.065 $Y=2.035
+ $X2=7.92 $Y2=2.035
r261 52 61 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=10.8 $Y2=2.035
r262 52 53 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=8.065 $Y2=2.035
r263 51 55 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=2.035
+ $X2=4.08 $Y2=2.035
r264 50 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r265 50 51 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=4.225 $Y2=2.035
r266 48 49 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=10.81 $Y=2.22
+ $X2=10.81 $Y2=2.37
r267 48 75 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=10.84 $Y=2.22
+ $X2=10.84 $Y2=2.01
r268 44 46 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=10.545 $Y=1.335
+ $X2=10.81 $Y2=1.335
r269 42 68 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=7.68 $Y=1.985
+ $X2=7.86 $Y2=1.985
r270 42 43 3.90195 $w=3.3e-07 $l=2.22374e-07 $layer=POLY_cond $X=7.68 $Y=1.985
+ $X2=7.465 $Y2=2
r271 38 40 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=7.31 $Y=1.165
+ $X2=7.605 $Y2=1.165
r272 36 64 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=3.685 $Y=1.985
+ $X2=3.95 $Y2=1.985
r273 36 37 3.90195 $w=3.3e-07 $l=3.4271e-07 $layer=POLY_cond $X=3.685 $Y=1.985
+ $X2=3.415 $Y2=1.82
r274 34 35 100.466 $w=1.55e-07 $l=2.1e-07 $layer=POLY_cond $X=3.487 $Y=0.935
+ $X2=3.487 $Y2=1.145
r275 30 46 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.81 $Y=1.41
+ $X2=10.81 $Y2=1.335
r276 30 74 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=10.81 $Y=1.41
+ $X2=10.81 $Y2=1.68
r277 29 49 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=10.795 $Y=2.655
+ $X2=10.795 $Y2=2.37
r278 23 44 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.545 $Y=1.26
+ $X2=10.545 $Y2=1.335
r279 23 25 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=10.545 $Y=1.26
+ $X2=10.545 $Y2=0.58
r280 22 43 34.7346 $w=1.65e-07 $l=2.4e-07 $layer=POLY_cond $X=7.605 $Y=1.82
+ $X2=7.465 $Y2=2
r281 21 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.605 $Y=1.24
+ $X2=7.605 $Y2=1.165
r282 21 22 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.605 $Y=1.24
+ $X2=7.605 $Y2=1.82
r283 17 43 34.7346 $w=1.65e-07 $l=1.89737e-07 $layer=POLY_cond $X=7.555 $Y=2.15
+ $X2=7.465 $Y2=2
r284 17 19 145.766 $w=1.8e-07 $l=3.75e-07 $layer=POLY_cond $X=7.555 $Y=2.15
+ $X2=7.555 $Y2=2.525
r285 14 38 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.31 $Y=1.09
+ $X2=7.31 $Y2=1.165
r286 14 16 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.31 $Y=1.09
+ $X2=7.31 $Y2=0.805
r287 13 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7.31 $Y=0.255
+ $X2=7.31 $Y2=0.805
r288 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.235 $Y=0.18
+ $X2=7.31 $Y2=0.255
r289 11 12 1884.41 $w=1.5e-07 $l=3.675e-06 $layer=POLY_cond $X=7.235 $Y=0.18
+ $X2=3.56 $Y2=0.18
r290 7 37 34.7346 $w=1.65e-07 $l=4.10244e-07 $layer=POLY_cond $X=3.595 $Y=2.15
+ $X2=3.415 $Y2=1.82
r291 7 9 190.468 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=3.595 $Y=2.15
+ $X2=3.595 $Y2=2.64
r292 6 37 34.7346 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=3.49 $Y=1.82
+ $X2=3.415 $Y2=1.82
r293 6 35 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=3.49 $Y=1.82
+ $X2=3.49 $Y2=1.145
r294 4 34 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.485 $Y=0.65
+ $X2=3.485 $Y2=0.935
r295 1 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.485 $Y=0.255
+ $X2=3.56 $Y2=0.18
r296 1 4 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.485 $Y=0.255
+ $X2=3.485 $Y2=0.65
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_1%A_1235_119# 1 2 3 12 16 18 22 27 28 31 32
+ 34 37 42
c111 34 0 2.05564e-20 $X=8.105 $Y=1.41
c112 22 0 1.68464e-19 $X=6.675 $Y=2.585
r113 35 42 23.6275 $w=2.55e-07 $l=1.25e-07 $layer=POLY_cond $X=8.105 $Y=1.42
+ $X2=8.23 $Y2=1.42
r114 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.105
+ $Y=1.41 $X2=8.105 $Y2=1.41
r115 32 34 22.622 $w=2.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.575 $Y=1.41
+ $X2=8.105 $Y2=1.41
r116 31 40 10.6888 $w=3.31e-07 $l=3.83445e-07 $layer=LI1_cond $X=7.49 $Y=2.32
+ $X2=7.78 $Y2=2.537
r117 30 32 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=7.49 $Y=1.545
+ $X2=7.575 $Y2=1.41
r118 30 31 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=7.49 $Y=1.545
+ $X2=7.49 $Y2=2.32
r119 29 37 3.64284 $w=2.55e-07 $l=1.69245e-07 $layer=LI1_cond $X=6.845 $Y=2.405
+ $X2=6.76 $Y2=2.537
r120 28 31 6.01027 $w=3.31e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.405 $Y=2.405
+ $X2=7.49 $Y2=2.32
r121 28 29 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.405 $Y=2.405
+ $X2=6.845 $Y2=2.405
r122 27 37 2.83584 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=6.76 $Y=2.32
+ $X2=6.76 $Y2=2.537
r123 26 27 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=6.76 $Y=0.925
+ $X2=6.76 $Y2=2.32
r124 22 37 3.64284 $w=2.55e-07 $l=1.06325e-07 $layer=LI1_cond $X=6.675 $Y=2.585
+ $X2=6.76 $Y2=2.537
r125 22 24 11.355 $w=3.38e-07 $l=3.35e-07 $layer=LI1_cond $X=6.675 $Y=2.585
+ $X2=6.34 $Y2=2.585
r126 18 26 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.675 $Y=0.76
+ $X2=6.76 $Y2=0.925
r127 18 20 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=6.675 $Y=0.76
+ $X2=6.315 $Y2=0.76
r128 14 42 59.5412 $w=2.55e-07 $l=3.92874e-07 $layer=POLY_cond $X=8.545 $Y=1.595
+ $X2=8.23 $Y2=1.42
r129 14 16 248.774 $w=1.8e-07 $l=6.4e-07 $layer=POLY_cond $X=8.545 $Y=1.595
+ $X2=8.545 $Y2=2.235
r130 10 42 15.178 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=8.23 $Y=1.245
+ $X2=8.23 $Y2=1.42
r131 10 12 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=8.23 $Y=1.245
+ $X2=8.23 $Y2=0.69
r132 3 40 600 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_PDIFF $count=1 $X=7.645
+ $Y=2.315 $X2=7.78 $Y2=2.535
r133 2 24 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=6.205
+ $Y=2.315 $X2=6.34 $Y2=2.585
r134 1 20 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=6.175
+ $Y=0.595 $X2=6.315 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_1%A_819_119# 1 2 9 12 13 16 18 19 20 21 22 23
+ 25 28 30 35 36 37 40 42 43 44 46 49 51 55 56 64 67 68 70
c190 67 0 9.8866e-20 $X=5.13 $Y=1.485
c191 51 0 1.21651e-19 $X=4.9 $Y=1.945
c192 40 0 1.87517e-19 $X=9.755 $Y=0.58
c193 37 0 6.061e-20 $X=9.085 $Y=1.585
c194 36 0 2.17443e-21 $X=9.68 $Y=1.585
c195 20 0 1.7726e-19 $X=5.68 $Y=1.165
c196 18 0 2.20311e-19 $X=5.605 $Y=3.075
c197 1 0 1.43966e-19 $X=4.095 $Y=0.595
r198 67 68 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.13 $Y=1.485
+ $X2=5.13 $Y2=1.41
r199 65 70 55.5535 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=5.13 $Y=1.61
+ $X2=5.13 $Y2=1.86
r200 65 67 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.13 $Y=1.61
+ $X2=5.13 $Y2=1.485
r201 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.13
+ $Y=1.61 $X2=5.13 $Y2=1.61
r202 61 64 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=4.9 $Y=1.61
+ $X2=5.13 $Y2=1.61
r203 56 59 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.46 $Y=2.03 $X2=4.46
+ $Y2=2.11
r204 53 55 9.12989 $w=4.13e-07 $l=1.8e-07 $layer=LI1_cond $X=4.31 $Y=0.802
+ $X2=4.49 $Y2=0.802
r205 50 61 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.9 $Y=1.775
+ $X2=4.9 $Y2=1.61
r206 50 51 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.9 $Y=1.775
+ $X2=4.9 $Y2=1.945
r207 49 61 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.9 $Y=1.445
+ $X2=4.9 $Y2=1.61
r208 48 49 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.9 $Y=1.01
+ $X2=4.9 $Y2=1.445
r209 47 56 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.585 $Y=2.03
+ $X2=4.46 $Y2=2.03
r210 46 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.815 $Y=2.03
+ $X2=4.9 $Y2=1.945
r211 46 47 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.815 $Y=2.03
+ $X2=4.585 $Y2=2.03
r212 44 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.815 $Y=0.925
+ $X2=4.9 $Y2=1.01
r213 44 55 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.815 $Y=0.925
+ $X2=4.49 $Y2=0.925
r214 38 40 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=9.755 $Y=1.51
+ $X2=9.755 $Y2=0.58
r215 36 38 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.68 $Y=1.585
+ $X2=9.755 $Y2=1.51
r216 36 37 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=9.68 $Y=1.585
+ $X2=9.085 $Y2=1.585
r217 33 35 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=8.995 $Y=3.075
+ $X2=8.995 $Y2=2.235
r218 32 37 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.995 $Y=1.66
+ $X2=9.085 $Y2=1.585
r219 32 35 223.508 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.995 $Y=1.66
+ $X2=8.995 $Y2=2.235
r220 31 43 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.655 $Y=3.15
+ $X2=6.565 $Y2=3.15
r221 30 33 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.905 $Y=3.15
+ $X2=8.995 $Y2=3.075
r222 30 31 1153.72 $w=1.5e-07 $l=2.25e-06 $layer=POLY_cond $X=8.905 $Y=3.15
+ $X2=6.655 $Y2=3.15
r223 26 43 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=6.565 $Y=3.075
+ $X2=6.565 $Y2=3.15
r224 26 28 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=6.565 $Y=3.075
+ $X2=6.565 $Y2=2.525
r225 23 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.1 $Y=1.09 $X2=6.1
+ $Y2=0.805
r226 21 43 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.475 $Y=3.15
+ $X2=6.565 $Y2=3.15
r227 21 22 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=6.475 $Y=3.15
+ $X2=5.68 $Y2=3.15
r228 19 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.025 $Y=1.165
+ $X2=6.1 $Y2=1.09
r229 19 20 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=6.025 $Y=1.165
+ $X2=5.68 $Y2=1.165
r230 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.605 $Y=3.075
+ $X2=5.68 $Y2=3.15
r231 17 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.605 $Y=1.56
+ $X2=5.605 $Y2=1.485
r232 17 18 776.84 $w=1.5e-07 $l=1.515e-06 $layer=POLY_cond $X=5.605 $Y=1.56
+ $X2=5.605 $Y2=3.075
r233 16 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.605 $Y=1.41
+ $X2=5.605 $Y2=1.485
r234 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.605 $Y=1.24
+ $X2=5.68 $Y2=1.165
r235 15 16 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=5.605 $Y=1.24
+ $X2=5.605 $Y2=1.41
r236 14 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.295 $Y=1.485
+ $X2=5.13 $Y2=1.485
r237 13 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.53 $Y=1.485
+ $X2=5.605 $Y2=1.485
r238 13 14 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=5.53 $Y=1.485
+ $X2=5.295 $Y2=1.485
r239 12 68 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.11 $Y=0.965
+ $X2=5.11 $Y2=1.41
r240 9 70 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=5.095 $Y=2.495
+ $X2=5.095 $Y2=1.86
r241 2 59 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.275
+ $Y=1.935 $X2=4.42 $Y2=2.11
r242 1 53 182 $w=1.7e-07 $l=3.40955e-07 $layer=licon1_NDIFF $count=1 $X=4.095
+ $Y=0.595 $X2=4.31 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_1%A_2008_48# 1 2 9 11 13 17 20 21 24 27 28 30
+ 31 33 34 36
c132 28 0 1.60243e-20 $X=11.675 $Y=0.665
c133 20 0 2.44776e-20 $X=10.855 $Y=2.405
c134 17 0 6.47027e-20 $X=10.36 $Y=1.815
r135 36 38 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=11.12 $Y=0.55
+ $X2=11.12 $Y2=0.665
r136 32 33 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=11.76 $Y=0.75
+ $X2=11.76 $Y2=1.63
r137 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.675 $Y=1.715
+ $X2=11.76 $Y2=1.63
r138 30 31 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=11.675 $Y=1.715
+ $X2=11.405 $Y2=1.715
r139 29 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.285 $Y=0.665
+ $X2=11.12 $Y2=0.665
r140 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.675 $Y=0.665
+ $X2=11.76 $Y2=0.75
r141 28 29 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=11.675 $Y=0.665
+ $X2=11.285 $Y2=0.665
r142 27 34 3.70735 $w=2.5e-07 $l=2.28583e-07 $layer=LI1_cond $X=11.32 $Y=2.32
+ $X2=11.13 $Y2=2.405
r143 26 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.32 $Y=1.8
+ $X2=11.405 $Y2=1.715
r144 26 27 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=11.32 $Y=1.8
+ $X2=11.32 $Y2=2.32
r145 22 34 3.70735 $w=2.5e-07 $l=1.46458e-07 $layer=LI1_cond $X=11.02 $Y=2.49
+ $X2=11.13 $Y2=2.405
r146 22 24 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=11.02 $Y=2.49
+ $X2=11.02 $Y2=2.655
r147 20 34 2.76166 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=10.855 $Y=2.405
+ $X2=11.13 $Y2=2.405
r148 20 21 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=10.855 $Y=2.405
+ $X2=10.525 $Y2=2.405
r149 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.36
+ $Y=1.815 $X2=10.36 $Y2=1.815
r150 15 21 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=10.395 $Y=2.32
+ $X2=10.525 $Y2=2.405
r151 15 17 22.384 $w=2.58e-07 $l=5.05e-07 $layer=LI1_cond $X=10.395 $Y=2.32
+ $X2=10.395 $Y2=1.815
r152 11 18 34.2225 $w=3.69e-07 $l=2.17612e-07 $layer=POLY_cond $X=10.16 $Y=1.98
+ $X2=10.282 $Y2=1.815
r153 11 13 262.379 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=10.16 $Y=1.98
+ $X2=10.16 $Y2=2.655
r154 7 18 58.6339 $w=3.69e-07 $l=3.89654e-07 $layer=POLY_cond $X=10.115 $Y=1.5
+ $X2=10.282 $Y2=1.815
r155 7 9 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=10.115 $Y=1.5
+ $X2=10.115 $Y2=0.58
r156 2 24 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=10.885
+ $Y=2.445 $X2=11.02 $Y2=2.655
r157 1 36 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=10.98
+ $Y=0.37 $X2=11.12 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_1%A_1747_74# 1 2 7 9 10 11 14 19 21 23 24 25
+ 28 32 38 39 40 43 45 49 50 54 56 57 59
c170 56 0 8.18368e-20 $X=10.01 $Y=2.425
c171 10 0 1.78926e-19 $X=11.26 $Y=1.02
c172 7 0 1.60243e-20 $X=10.905 $Y=0.87
r173 66 67 4.79602 $w=4.02e-07 $l=4e-08 $layer=POLY_cond $X=11.925 $Y=1.46
+ $X2=11.965 $Y2=1.46
r174 65 66 68.9428 $w=4.02e-07 $l=5.75e-07 $layer=POLY_cond $X=11.35 $Y=1.46
+ $X2=11.925 $Y2=1.46
r175 62 63 15.0154 $w=2.6e-07 $l=3.2e-07 $layer=LI1_cond $X=9.69 $Y=1.175
+ $X2=10.01 $Y2=1.175
r176 57 63 4.30428 $w=4.3e-07 $l=1.05119e-07 $layer=LI1_cond $X=10.095 $Y=1.22
+ $X2=10.01 $Y2=1.175
r177 57 59 31.2232 $w=4.28e-07 $l=1.165e-06 $layer=LI1_cond $X=10.095 $Y=1.22
+ $X2=11.26 $Y2=1.22
r178 55 63 3.22376 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=10.01 $Y=1.435
+ $X2=10.01 $Y2=1.175
r179 55 56 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=10.01 $Y=1.435
+ $X2=10.01 $Y2=2.425
r180 54 62 3.22376 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=9.69 $Y=1.005
+ $X2=9.69 $Y2=1.175
r181 53 54 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.69 $Y=0.735
+ $X2=9.69 $Y2=1.005
r182 50 52 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=9.325 $Y=2.59
+ $X2=9.545 $Y2=2.59
r183 49 56 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.925 $Y=2.59
+ $X2=10.01 $Y2=2.425
r184 49 52 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=9.925 $Y=2.59
+ $X2=9.545 $Y2=2.59
r185 45 53 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.605 $Y=0.57
+ $X2=9.69 $Y2=0.735
r186 45 47 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=9.605 $Y=0.57
+ $X2=9.37 $Y2=0.57
r187 41 50 7.17723 $w=3.3e-07 $l=2.13014e-07 $layer=LI1_cond $X=9.215 $Y=2.425
+ $X2=9.325 $Y2=2.59
r188 41 43 26.4538 $w=2.18e-07 $l=5.05e-07 $layer=LI1_cond $X=9.215 $Y=2.425
+ $X2=9.215 $Y2=1.92
r189 38 39 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=11.29 $Y=2.22
+ $X2=11.29 $Y2=2.37
r190 30 40 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=12.93 $Y=1.355
+ $X2=12.915 $Y2=1.52
r191 30 32 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=12.93 $Y=1.355
+ $X2=12.93 $Y2=0.645
r192 26 40 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=12.915 $Y=1.685
+ $X2=12.915 $Y2=1.52
r193 26 28 332.347 $w=1.8e-07 $l=8.55e-07 $layer=POLY_cond $X=12.915 $Y=1.685
+ $X2=12.915 $Y2=2.54
r194 25 67 10.6813 $w=4.02e-07 $l=1.00623e-07 $layer=POLY_cond $X=12.04 $Y=1.52
+ $X2=11.965 $Y2=1.46
r195 24 40 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=12.825 $Y=1.52
+ $X2=12.915 $Y2=1.52
r196 24 25 137.266 $w=3.3e-07 $l=7.85e-07 $layer=POLY_cond $X=12.825 $Y=1.52
+ $X2=12.04 $Y2=1.52
r197 21 67 25.9839 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=11.965 $Y=1.235
+ $X2=11.965 $Y2=1.46
r198 21 23 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=11.965 $Y=1.235
+ $X2=11.965 $Y2=0.74
r199 17 66 21.5811 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=11.925 $Y=1.685
+ $X2=11.925 $Y2=1.46
r200 17 19 277.927 $w=1.8e-07 $l=7.15e-07 $layer=POLY_cond $X=11.925 $Y=1.685
+ $X2=11.925 $Y2=2.4
r201 15 65 25.9839 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=11.35 $Y=1.685
+ $X2=11.35 $Y2=1.46
r202 15 38 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=11.35 $Y=1.685
+ $X2=11.35 $Y2=2.22
r203 14 39 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=11.245 $Y=2.655
+ $X2=11.245 $Y2=2.37
r204 11 65 10.791 $w=4.02e-07 $l=2.66224e-07 $layer=POLY_cond $X=11.26 $Y=1.235
+ $X2=11.35 $Y2=1.46
r205 11 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.26
+ $Y=1.27 $X2=11.26 $Y2=1.27
r206 10 34 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=11.26 $Y=0.945
+ $X2=10.905 $Y2=0.945
r207 10 11 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=11.26 $Y=1.02
+ $X2=11.26 $Y2=1.235
r208 7 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.905 $Y=0.87
+ $X2=10.905 $Y2=0.945
r209 7 9 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=10.905 $Y=0.87
+ $X2=10.905 $Y2=0.58
r210 2 52 600 $w=1.7e-07 $l=1.06034e-06 $layer=licon1_PDIFF $count=1 $X=9.085
+ $Y=1.735 $X2=9.545 $Y2=2.59
r211 2 43 300 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=2 $X=9.085
+ $Y=1.735 $X2=9.22 $Y2=1.92
r212 1 47 182 $w=1.7e-07 $l=7.28166e-07 $layer=licon1_NDIFF $count=1 $X=8.735
+ $Y=0.37 $X2=9.37 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_1%A_2513_424# 1 2 9 13 17 21 25 26 28
r50 26 31 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.38 $Y=1.465
+ $X2=13.38 $Y2=1.63
r51 26 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.38 $Y=1.465
+ $X2=13.38 $Y2=1.3
r52 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.38
+ $Y=1.465 $X2=13.38 $Y2=1.465
r53 23 28 0.820356 $w=3.3e-07 $l=1.43e-07 $layer=LI1_cond $X=12.855 $Y=1.465
+ $X2=12.712 $Y2=1.465
r54 23 25 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=12.855 $Y=1.465
+ $X2=13.38 $Y2=1.465
r55 19 28 5.82594 $w=2.85e-07 $l=1.65e-07 $layer=LI1_cond $X=12.712 $Y=1.63
+ $X2=12.712 $Y2=1.465
r56 19 21 25.6772 $w=2.83e-07 $l=6.35e-07 $layer=LI1_cond $X=12.712 $Y=1.63
+ $X2=12.712 $Y2=2.265
r57 15 28 5.82594 $w=2.85e-07 $l=1.65e-07 $layer=LI1_cond $X=12.712 $Y=1.3
+ $X2=12.712 $Y2=1.465
r58 15 17 26.486 $w=2.83e-07 $l=6.55e-07 $layer=LI1_cond $X=12.712 $Y=1.3
+ $X2=12.712 $Y2=0.645
r59 13 31 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=13.435 $Y=2.4
+ $X2=13.435 $Y2=1.63
r60 9 30 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.42 $Y=0.74
+ $X2=13.42 $Y2=1.3
r61 2 21 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=12.565
+ $Y=2.12 $X2=12.69 $Y2=2.265
r62 1 17 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=12.59
+ $Y=0.37 $X2=12.715 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_1%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 49 52
+ 55 59 64 65 67 68 70 71 73 75 84 101 105 110 115 122 123 126 129 132 135 138
c181 3 0 1.21651e-19 $X=4.735 $Y=1.935
r182 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r183 135 136 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r184 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r185 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r186 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r187 123 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=13.2 $Y2=3.33
r188 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r189 120 138 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=13.325 $Y=3.33
+ $X2=13.185 $Y2=3.33
r190 120 122 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=13.325 $Y=3.33
+ $X2=13.68 $Y2=3.33
r191 119 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r192 119 136 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=11.76 $Y2=3.33
r193 118 119 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r194 116 135 10.508 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=11.815 $Y=3.33
+ $X2=11.592 $Y2=3.33
r195 116 118 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=11.815 $Y=3.33
+ $X2=12.72 $Y2=3.33
r196 115 138 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=13.045 $Y=3.33
+ $X2=13.185 $Y2=3.33
r197 115 118 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=13.045 $Y=3.33
+ $X2=12.72 $Y2=3.33
r198 114 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r199 114 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.32 $Y2=3.33
r200 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r201 111 132 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=10.65 $Y=3.33
+ $X2=10.477 $Y2=3.33
r202 111 113 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=10.65 $Y=3.33
+ $X2=11.28 $Y2=3.33
r203 110 135 10.508 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=11.37 $Y=3.33
+ $X2=11.592 $Y2=3.33
r204 110 113 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=11.37 $Y=3.33
+ $X2=11.28 $Y2=3.33
r205 109 133 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r206 109 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r207 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r208 106 129 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.485 $Y=3.33
+ $X2=8.36 $Y2=3.33
r209 106 108 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=8.485 $Y=3.33
+ $X2=8.88 $Y2=3.33
r210 105 132 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=10.305 $Y=3.33
+ $X2=10.477 $Y2=3.33
r211 105 108 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=10.305 $Y=3.33
+ $X2=8.88 $Y2=3.33
r212 104 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r213 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r214 101 129 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.235 $Y=3.33
+ $X2=8.36 $Y2=3.33
r215 101 103 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.235 $Y=3.33
+ $X2=7.92 $Y2=3.33
r216 96 99 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r217 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r218 94 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r219 93 94 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r220 91 94 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r221 91 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r222 90 93 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r223 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r224 88 126 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.445 $Y=3.33
+ $X2=3.265 $Y2=3.33
r225 88 90 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.445 $Y=3.33
+ $X2=3.6 $Y2=3.33
r226 87 127 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r227 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r228 84 126 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.085 $Y=3.33
+ $X2=3.265 $Y2=3.33
r229 84 86 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=3.085 $Y=3.33
+ $X2=1.68 $Y2=3.33
r230 83 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r231 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r232 79 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r233 78 82 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r234 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r235 75 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r236 75 97 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=5.04 $Y2=3.33
r237 75 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r238 73 74 5.78802 $w=4.43e-07 $l=1.2e-07 $layer=LI1_cond $X=11.592 $Y=2.815
+ $X2=11.592 $Y2=2.695
r239 70 99 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=7.09 $Y=3.33
+ $X2=6.96 $Y2=3.33
r240 70 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.09 $Y=3.33
+ $X2=7.255 $Y2=3.33
r241 69 103 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=7.42 $Y=3.33
+ $X2=7.92 $Y2=3.33
r242 69 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.42 $Y=3.33
+ $X2=7.255 $Y2=3.33
r243 67 93 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.56 $Y2=3.33
r244 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.87 $Y2=3.33
r245 66 96 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=5.04 $Y2=3.33
r246 66 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=4.87 $Y2=3.33
r247 64 82 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.2 $Y2=3.33
r248 64 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.39 $Y2=3.33
r249 63 86 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.68 $Y2=3.33
r250 63 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.39 $Y2=3.33
r251 59 62 17.0809 $w=2.78e-07 $l=4.15e-07 $layer=LI1_cond $X=13.185 $Y=1.985
+ $X2=13.185 $Y2=2.4
r252 57 138 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=13.185 $Y=3.245
+ $X2=13.185 $Y2=3.33
r253 57 62 34.7791 $w=2.78e-07 $l=8.45e-07 $layer=LI1_cond $X=13.185 $Y=3.245
+ $X2=13.185 $Y2=2.4
r254 55 74 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=11.7 $Y=2.135
+ $X2=11.7 $Y2=2.695
r255 52 135 1.76584 $w=4.45e-07 $l=8.5e-08 $layer=LI1_cond $X=11.592 $Y=3.245
+ $X2=11.592 $Y2=3.33
r256 51 73 2.64155 $w=4.43e-07 $l=1.02e-07 $layer=LI1_cond $X=11.592 $Y=2.917
+ $X2=11.592 $Y2=2.815
r257 51 52 8.49441 $w=4.43e-07 $l=3.28e-07 $layer=LI1_cond $X=11.592 $Y=2.917
+ $X2=11.592 $Y2=3.245
r258 47 132 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=10.477 $Y=3.245
+ $X2=10.477 $Y2=3.33
r259 47 49 14.0297 $w=3.43e-07 $l=4.2e-07 $layer=LI1_cond $X=10.477 $Y=3.245
+ $X2=10.477 $Y2=2.825
r260 43 46 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=8.36 $Y=1.88
+ $X2=8.36 $Y2=2.59
r261 41 129 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.36 $Y=3.245
+ $X2=8.36 $Y2=3.33
r262 41 46 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=8.36 $Y=3.245
+ $X2=8.36 $Y2=2.59
r263 37 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.255 $Y=3.245
+ $X2=7.255 $Y2=3.33
r264 37 39 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=7.255 $Y=3.245
+ $X2=7.255 $Y2=2.825
r265 33 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=3.33
r266 33 35 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=2.88
r267 29 126 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.265 $Y=3.245
+ $X2=3.265 $Y2=3.33
r268 29 31 13.7653 $w=3.58e-07 $l=4.3e-07 $layer=LI1_cond $X=3.265 $Y=3.245
+ $X2=3.265 $Y2=2.815
r269 25 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.39 $Y=3.245
+ $X2=1.39 $Y2=3.33
r270 25 27 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.39 $Y=3.245
+ $X2=1.39 $Y2=2.475
r271 8 62 300 $w=1.7e-07 $l=3.54965e-07 $layer=licon1_PDIFF $count=2 $X=13.005
+ $Y=2.12 $X2=13.175 $Y2=2.4
r272 8 59 600 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_PDIFF $count=1 $X=13.005
+ $Y=2.12 $X2=13.21 $Y2=1.985
r273 7 73 600 $w=1.7e-07 $l=4.59238e-07 $layer=licon1_PDIFF $count=1 $X=11.335
+ $Y=2.445 $X2=11.535 $Y2=2.815
r274 7 55 300 $w=1.7e-07 $l=4.91121e-07 $layer=licon1_PDIFF $count=2 $X=11.335
+ $Y=2.445 $X2=11.695 $Y2=2.135
r275 6 49 600 $w=1.7e-07 $l=4.79479e-07 $layer=licon1_PDIFF $count=1 $X=10.25
+ $Y=2.445 $X2=10.475 $Y2=2.825
r276 5 46 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.185
+ $Y=1.735 $X2=8.32 $Y2=2.59
r277 5 43 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.185
+ $Y=1.735 $X2=8.32 $Y2=1.88
r278 4 39 600 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=1 $X=7.045
+ $Y=2.315 $X2=7.255 $Y2=2.825
r279 3 35 600 $w=1.7e-07 $l=1.01025e-06 $layer=licon1_PDIFF $count=1 $X=4.735
+ $Y=1.935 $X2=4.87 $Y2=2.88
r280 2 31 600 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=1 $X=3.115
+ $Y=2.32 $X2=3.265 $Y2=2.815
r281 1 27 300 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_PDIFF $count=2 $X=1.205
+ $Y=2.32 $X2=1.39 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_1%A_413_90# 1 2 3 4 5 18 20 23 26 29 32 34 35
+ 36 37 39 41 43 49
c145 49 0 7.88209e-20 $X=3.715 $Y=2.535
c146 41 0 1.29655e-19 $X=2.26 $Y=2.475
c147 39 0 5.18475e-20 $X=6.42 $Y=2.075
c148 32 0 1.92441e-20 $X=5.885 $Y=0.795
c149 26 0 2.39118e-20 $X=5.725 $Y=2.535
r150 48 49 1.45527 $w=5.03e-07 $l=6e-08 $layer=LI1_cond $X=3.715 $Y=2.475
+ $X2=3.715 $Y2=2.535
r151 43 45 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.435 $Y=0.76
+ $X2=2.435 $Y2=1.005
r152 38 39 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=6.42 $Y=1.265
+ $X2=6.42 $Y2=2.075
r153 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.335 $Y=1.18
+ $X2=6.42 $Y2=1.265
r154 36 37 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.335 $Y=1.18
+ $X2=5.98 $Y2=1.18
r155 34 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.335 $Y=2.16
+ $X2=6.42 $Y2=2.075
r156 34 35 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.335 $Y=2.16
+ $X2=5.975 $Y2=2.16
r157 30 37 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=5.89 $Y=1.095
+ $X2=5.98 $Y2=1.18
r158 30 32 18.4848 $w=1.78e-07 $l=3e-07 $layer=LI1_cond $X=5.89 $Y=1.095
+ $X2=5.89 $Y2=0.795
r159 29 51 3.38195 $w=1.85e-07 $l=1.7025e-07 $layer=LI1_cond $X=5.882 $Y=2.445
+ $X2=5.85 $Y2=2.6
r160 28 35 6.83233 $w=1.7e-07 $l=1.28662e-07 $layer=LI1_cond $X=5.882 $Y=2.245
+ $X2=5.975 $Y2=2.16
r161 28 29 11.9902 $w=1.83e-07 $l=2e-07 $layer=LI1_cond $X=5.882 $Y=2.245
+ $X2=5.882 $Y2=2.445
r162 27 49 6.83659 $w=1.8e-07 $l=2.7e-07 $layer=LI1_cond $X=3.985 $Y=2.535
+ $X2=3.715 $Y2=2.535
r163 26 51 3.43621 $w=1.8e-07 $l=1.5411e-07 $layer=LI1_cond $X=5.725 $Y=2.535
+ $X2=5.85 $Y2=2.6
r164 26 27 107.212 $w=1.78e-07 $l=1.74e-06 $layer=LI1_cond $X=5.725 $Y=2.535
+ $X2=3.985 $Y2=2.535
r165 23 48 9.48372 $w=5.03e-07 $l=2.50799e-07 $layer=LI1_cond $X=3.53 $Y=2.32
+ $X2=3.715 $Y2=2.475
r166 22 23 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=3.53 $Y=1.09
+ $X2=3.53 $Y2=2.32
r167 21 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.6 $Y=1.005
+ $X2=2.435 $Y2=1.005
r168 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.445 $Y=1.005
+ $X2=3.53 $Y2=1.09
r169 20 21 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=3.445 $Y=1.005
+ $X2=2.6 $Y2=1.005
r170 19 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.425 $Y=2.475
+ $X2=2.26 $Y2=2.475
r171 18 48 7.19425 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=3.445 $Y=2.475
+ $X2=3.715 $Y2=2.475
r172 18 19 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=3.445 $Y=2.475
+ $X2=2.425 $Y2=2.475
r173 5 51 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=5.755
+ $Y=2.315 $X2=5.89 $Y2=2.525
r174 4 48 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=3.685
+ $Y=2.32 $X2=3.82 $Y2=2.475
r175 3 41 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=2.125
+ $Y=2.32 $X2=2.26 $Y2=2.475
r176 2 32 182 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=1 $X=5.76
+ $Y=0.595 $X2=5.885 $Y2=0.795
r177 1 43 182 $w=1.7e-07 $l=5.01597e-07 $layer=licon1_NDIFF $count=1 $X=2.065
+ $Y=0.45 $X2=2.435 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_1%Q_N 1 2 7 8 9 10 11 12 13
r20 13 40 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=12.18 $Y=2.775
+ $X2=12.18 $Y2=2.815
r21 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.18 $Y=2.405
+ $X2=12.18 $Y2=2.775
r22 12 34 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=12.18 $Y=2.405
+ $X2=12.18 $Y2=2.055
r23 11 34 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=12.18 $Y=2.035
+ $X2=12.18 $Y2=2.055
r24 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.18 $Y=1.665
+ $X2=12.18 $Y2=2.035
r25 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.18 $Y=1.295
+ $X2=12.18 $Y2=1.665
r26 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.18 $Y=0.925
+ $X2=12.18 $Y2=1.295
r27 7 8 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=12.18 $Y=0.515
+ $X2=12.18 $Y2=0.925
r28 2 40 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=12.015
+ $Y=1.84 $X2=12.15 $Y2=2.815
r29 2 34 400 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=12.015
+ $Y=1.84 $X2=12.15 $Y2=2.055
r30 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.04
+ $Y=0.37 $X2=12.18 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_1%Q 1 2 9 10 11 12 13 28 32 43
r21 41 43 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=13.75 $Y=1.13
+ $X2=13.75 $Y2=1.82
r22 29 32 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=13.695 $Y=1.96
+ $X2=13.695 $Y2=1.985
r23 21 28 0.726197 $w=3.63e-07 $l=2.3e-08 $layer=LI1_cond $X=13.652 $Y=0.948
+ $X2=13.652 $Y2=0.925
r24 12 13 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=13.695 $Y=2.405
+ $X2=13.695 $Y2=2.775
r25 11 29 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=13.695 $Y=1.955
+ $X2=13.695 $Y2=1.96
r26 11 43 7.32213 $w=2.78e-07 $l=1.35e-07 $layer=LI1_cond $X=13.695 $Y=1.955
+ $X2=13.695 $Y2=1.82
r27 11 12 15.0229 $w=2.78e-07 $l=3.65e-07 $layer=LI1_cond $X=13.695 $Y=2.04
+ $X2=13.695 $Y2=2.405
r28 11 32 2.26373 $w=2.78e-07 $l=5.5e-08 $layer=LI1_cond $X=13.695 $Y=2.04
+ $X2=13.695 $Y2=1.985
r29 10 41 8.08227 $w=3.63e-07 $l=1.51e-07 $layer=LI1_cond $X=13.652 $Y=0.979
+ $X2=13.652 $Y2=1.13
r30 10 21 0.978787 $w=3.63e-07 $l=3.1e-08 $layer=LI1_cond $X=13.652 $Y=0.979
+ $X2=13.652 $Y2=0.948
r31 10 28 0.978787 $w=3.63e-07 $l=3.1e-08 $layer=LI1_cond $X=13.652 $Y=0.894
+ $X2=13.652 $Y2=0.925
r32 9 10 11.9665 $w=3.63e-07 $l=3.79e-07 $layer=LI1_cond $X=13.652 $Y=0.515
+ $X2=13.652 $Y2=0.894
r33 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=13.525
+ $Y=1.84 $X2=13.66 $Y2=2.815
r34 2 32 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=13.525
+ $Y=1.84 $X2=13.66 $Y2=1.985
r35 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.495
+ $Y=0.37 $X2=13.635 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_1%VGND 1 2 3 4 5 6 7 24 28 32 36 40 42 46 49
+ 50 51 53 58 67 71 79 86 87 90 93 96 99 103 109
c138 87 0 5.91383e-20 $X=13.68 $Y=0
r139 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r140 104 110 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=13.2 $Y2=0
r141 103 106 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=11.675 $Y=0
+ $X2=11.675 $Y2=0.325
r142 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r143 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r144 96 97 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r145 93 94 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r146 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r147 87 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r148 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r149 84 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.29 $Y=0
+ $X2=13.205 $Y2=0
r150 84 86 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=13.29 $Y=0
+ $X2=13.68 $Y2=0
r151 83 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r152 83 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.32 $Y2=0
r153 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r154 80 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.495 $Y=0
+ $X2=10.33 $Y2=0
r155 80 82 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=10.495 $Y=0
+ $X2=11.28 $Y2=0
r156 79 103 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.51 $Y=0
+ $X2=11.675 $Y2=0
r157 79 82 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=11.51 $Y=0
+ $X2=11.28 $Y2=0
r158 78 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r159 77 78 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r160 75 78 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=9.84 $Y2=0
r161 75 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r162 74 77 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=7.92 $Y=0 $X2=9.84
+ $Y2=0
r163 74 75 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r164 72 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.77 $Y=0 $X2=7.605
+ $Y2=0
r165 72 74 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=7.77 $Y=0 $X2=7.92
+ $Y2=0
r166 71 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.165 $Y=0
+ $X2=10.33 $Y2=0
r167 71 77 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=10.165 $Y=0
+ $X2=9.84 $Y2=0
r168 69 70 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r169 67 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.44 $Y=0 $X2=7.605
+ $Y2=0
r170 67 69 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=7.44 $Y=0 $X2=5.04
+ $Y2=0
r171 66 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r172 66 94 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r173 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r174 63 93 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.865 $Y=0
+ $X2=3.712 $Y2=0
r175 63 65 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.865 $Y=0
+ $X2=4.56 $Y2=0
r176 62 94 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r177 62 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r178 61 62 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r179 59 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r180 59 61 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r181 58 93 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.56 $Y=0 $X2=3.712
+ $Y2=0
r182 58 61 153.968 $w=1.68e-07 $l=2.36e-06 $layer=LI1_cond $X=3.56 $Y=0 $X2=1.2
+ $Y2=0
r183 56 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r184 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r185 53 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r186 53 55 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r187 51 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r188 51 70 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=5.04 $Y2=0
r189 49 65 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.66 $Y=0 $X2=4.56
+ $Y2=0
r190 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.66 $Y=0 $X2=4.825
+ $Y2=0
r191 48 69 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=4.99 $Y=0 $X2=5.04
+ $Y2=0
r192 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.99 $Y=0 $X2=4.825
+ $Y2=0
r193 44 109 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.205 $Y=0.085
+ $X2=13.205 $Y2=0
r194 44 46 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=13.205 $Y=0.085
+ $X2=13.205 $Y2=0.515
r195 43 103 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.84 $Y=0
+ $X2=11.675 $Y2=0
r196 42 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.12 $Y=0
+ $X2=13.205 $Y2=0
r197 42 43 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=13.12 $Y=0
+ $X2=11.84 $Y2=0
r198 38 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.33 $Y=0.085
+ $X2=10.33 $Y2=0
r199 38 40 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.33 $Y=0.085
+ $X2=10.33 $Y2=0.58
r200 34 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.605 $Y=0.085
+ $X2=7.605 $Y2=0
r201 34 36 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=7.605 $Y=0.085
+ $X2=7.605 $Y2=0.34
r202 30 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.825 $Y=0.085
+ $X2=4.825 $Y2=0
r203 30 32 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=4.825 $Y=0.085
+ $X2=4.825 $Y2=0.585
r204 26 93 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.712 $Y=0.085
+ $X2=3.712 $Y2=0
r205 26 28 18.8925 $w=3.03e-07 $l=5e-07 $layer=LI1_cond $X=3.712 $Y=0.085
+ $X2=3.712 $Y2=0.585
r206 22 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r207 22 24 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.58
r208 7 46 91 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=2 $X=13.005
+ $Y=0.37 $X2=13.205 $Y2=0.515
r209 6 106 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=11.535
+ $Y=0.18 $X2=11.675 $Y2=0.325
r210 5 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.19
+ $Y=0.37 $X2=10.33 $Y2=0.58
r211 4 36 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=7.385
+ $Y=0.595 $X2=7.605 $Y2=0.34
r212 3 32 182 $w=1.7e-07 $l=2.14942e-07 $layer=licon1_NDIFF $count=1 $X=4.615
+ $Y=0.595 $X2=4.825 $Y2=0.585
r213 2 28 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.44 $X2=3.7 $Y2=0.585
r214 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRBP_1%noxref_25 1 2 9 11 12 13
c33 11 0 1.87424e-19 $X=3.06 $Y=0.34
r34 13 16 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.225 $Y=0.34
+ $X2=3.225 $Y2=0.665
r35 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.06 $Y=0.34
+ $X2=3.225 $Y2=0.34
r36 11 12 111.235 $w=1.68e-07 $l=1.705e-06 $layer=LI1_cond $X=3.06 $Y=0.34
+ $X2=1.355 $Y2=0.34
r37 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.23 $Y=0.425
+ $X2=1.355 $Y2=0.34
r38 7 9 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=1.23 $Y=0.425
+ $X2=1.23 $Y2=0.62
r39 2 16 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.085
+ $Y=0.485 $X2=3.225 $Y2=0.665
r40 1 9 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.45 $X2=1.27 $Y2=0.62
.ends


* File: sky130_fd_sc_ms__o21ba_4.pxi.spice
* Created: Wed Sep  2 12:22:23 2020
* 
x_PM_SKY130_FD_SC_MS__O21BA_4%B1_N N_B1_N_M1010_g N_B1_N_M1020_g B1_N
+ N_B1_N_c_121_n N_B1_N_c_122_n PM_SKY130_FD_SC_MS__O21BA_4%B1_N
x_PM_SKY130_FD_SC_MS__O21BA_4%A_193_48# N_A_193_48#_M1008_d N_A_193_48#_M1017_d
+ N_A_193_48#_M1016_d N_A_193_48#_M1003_g N_A_193_48#_M1001_g
+ N_A_193_48#_M1005_g N_A_193_48#_M1002_g N_A_193_48#_M1013_g
+ N_A_193_48#_M1007_g N_A_193_48#_M1018_g N_A_193_48#_M1011_g
+ N_A_193_48#_c_160_n N_A_193_48#_c_161_n N_A_193_48#_c_162_n
+ N_A_193_48#_c_163_n N_A_193_48#_c_164_n N_A_193_48#_c_183_p
+ N_A_193_48#_c_165_n N_A_193_48#_c_172_n N_A_193_48#_c_173_n
+ N_A_193_48#_c_273_p N_A_193_48#_c_166_n N_A_193_48#_c_174_n
+ N_A_193_48#_c_167_n PM_SKY130_FD_SC_MS__O21BA_4%A_193_48#
x_PM_SKY130_FD_SC_MS__O21BA_4%A_27_368# N_A_27_368#_M1020_s N_A_27_368#_M1010_s
+ N_A_27_368#_M1017_g N_A_27_368#_M1008_g N_A_27_368#_M1019_g
+ N_A_27_368#_M1015_g N_A_27_368#_c_312_n N_A_27_368#_c_319_n
+ N_A_27_368#_c_320_n N_A_27_368#_c_330_n N_A_27_368#_c_321_n
+ N_A_27_368#_c_313_n N_A_27_368#_c_322_n N_A_27_368#_c_314_n
+ N_A_27_368#_c_324_n N_A_27_368#_c_315_n N_A_27_368#_c_316_n
+ PM_SKY130_FD_SC_MS__O21BA_4%A_27_368#
x_PM_SKY130_FD_SC_MS__O21BA_4%A2 N_A2_M1016_g N_A2_M1004_g N_A2_M1021_g
+ N_A2_M1009_g A2 A2 A2 N_A2_c_408_n PM_SKY130_FD_SC_MS__O21BA_4%A2
x_PM_SKY130_FD_SC_MS__O21BA_4%A1 N_A1_M1000_g N_A1_M1006_g N_A1_c_459_n
+ N_A1_c_460_n N_A1_c_461_n N_A1_M1014_g N_A1_M1012_g A1 N_A1_c_465_n
+ PM_SKY130_FD_SC_MS__O21BA_4%A1
x_PM_SKY130_FD_SC_MS__O21BA_4%VPWR N_VPWR_M1010_d N_VPWR_M1002_s N_VPWR_M1011_s
+ N_VPWR_M1019_s N_VPWR_M1014_d N_VPWR_c_529_n N_VPWR_c_530_n N_VPWR_c_531_n
+ N_VPWR_c_532_n N_VPWR_c_533_n VPWR N_VPWR_c_534_n N_VPWR_c_535_n
+ N_VPWR_c_536_n N_VPWR_c_537_n N_VPWR_c_538_n N_VPWR_c_539_n N_VPWR_c_540_n
+ N_VPWR_c_541_n N_VPWR_c_542_n N_VPWR_c_528_n PM_SKY130_FD_SC_MS__O21BA_4%VPWR
x_PM_SKY130_FD_SC_MS__O21BA_4%X N_X_M1003_s N_X_M1013_s N_X_M1001_d N_X_M1007_d
+ N_X_c_606_n N_X_c_612_n N_X_c_607_n N_X_c_608_n N_X_c_609_n X X N_X_c_615_n X
+ N_X_c_611_n PM_SKY130_FD_SC_MS__O21BA_4%X
x_PM_SKY130_FD_SC_MS__O21BA_4%A_895_392# N_A_895_392#_M1000_s
+ N_A_895_392#_M1021_s N_A_895_392#_c_662_n N_A_895_392#_c_658_n
+ N_A_895_392#_c_659_n N_A_895_392#_c_660_n
+ PM_SKY130_FD_SC_MS__O21BA_4%A_895_392#
x_PM_SKY130_FD_SC_MS__O21BA_4%VGND N_VGND_M1020_d N_VGND_M1005_d N_VGND_M1018_d
+ N_VGND_M1006_s N_VGND_M1009_d N_VGND_c_686_n N_VGND_c_687_n N_VGND_c_688_n
+ N_VGND_c_689_n N_VGND_c_690_n N_VGND_c_691_n N_VGND_c_692_n VGND
+ N_VGND_c_693_n N_VGND_c_694_n N_VGND_c_695_n N_VGND_c_696_n N_VGND_c_697_n
+ N_VGND_c_698_n N_VGND_c_699_n N_VGND_c_700_n N_VGND_c_701_n
+ PM_SKY130_FD_SC_MS__O21BA_4%VGND
x_PM_SKY130_FD_SC_MS__O21BA_4%A_618_94# N_A_618_94#_M1008_s N_A_618_94#_M1015_s
+ N_A_618_94#_M1004_s N_A_618_94#_M1012_d N_A_618_94#_c_786_n
+ N_A_618_94#_c_777_n N_A_618_94#_c_778_n N_A_618_94#_c_779_n
+ N_A_618_94#_c_780_n N_A_618_94#_c_781_n N_A_618_94#_c_782_n
+ N_A_618_94#_c_783_n N_A_618_94#_c_784_n N_A_618_94#_c_785_n
+ PM_SKY130_FD_SC_MS__O21BA_4%A_618_94#
cc_1 VNB N_B1_N_M1010_g 0.00699056f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB B1_N 0.00980764f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_B1_N_c_121_n 0.0368096f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_4 VNB N_B1_N_c_122_n 0.0222506f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.22
cc_5 VNB N_A_193_48#_M1003_g 0.0210367f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_6 VNB N_A_193_48#_M1001_g 0.00589833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_193_48#_M1005_g 0.0199949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_193_48#_M1002_g 0.00206447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_193_48#_M1013_g 0.020485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_193_48#_M1007_g 0.00207413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_193_48#_M1018_g 0.0235858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_193_48#_M1011_g 0.0027323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_193_48#_c_160_n 0.0209991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_193_48#_c_161_n 0.0190649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_193_48#_c_162_n 0.0166372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_193_48#_c_163_n 0.0034847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_193_48#_c_164_n 0.0206699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_193_48#_c_165_n 0.00158703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_193_48#_c_166_n 0.0112053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_193_48#_c_167_n 0.0876246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_368#_M1008_g 0.0421943f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.22
cc_22 VNB N_A_27_368#_M1015_g 0.0367602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_368#_c_312_n 0.0222049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_368#_c_313_n 0.0079873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_368#_c_314_n 0.0300772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_368#_c_315_n 5.55182e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_368#_c_316_n 0.0118623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A2_M1004_g 0.0196921f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.74
cc_29 VNB N_A2_M1009_g 0.0180242f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.365
cc_30 VNB A2 0.0144679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A2_c_408_n 0.0249586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A1_M1006_g 0.0327623f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_33 VNB N_A1_c_459_n 0.0975279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A1_c_460_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.385
cc_35 VNB N_A1_c_461_n 0.0084508f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_36 VNB N_A1_M1014_g 0.0143086f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.22
cc_37 VNB N_A1_M1012_g 0.0360452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB A1 0.00447618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A1_c_465_n 0.016405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VPWR_c_528_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_606_n 0.00202189f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.365
cc_42 VNB N_X_c_607_n 0.00629496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_X_c_608_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_X_c_609_n 0.00111459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB X 7.86953e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_X_c_611_n 0.00286244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_686_n 0.00587905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_687_n 0.00412957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_688_n 0.00722278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_689_n 0.0100107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_690_n 0.00760342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_691_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_692_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_693_n 0.0157739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_694_n 0.0469424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_695_n 0.0160823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_696_n 0.0195709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_697_n 0.350143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_698_n 0.0258092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_699_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_700_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_701_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_618_94#_c_777_n 0.00431549f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.365
cc_64 VNB N_A_618_94#_c_778_n 0.00135951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_618_94#_c_779_n 0.00127304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_618_94#_c_780_n 0.00363185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_618_94#_c_781_n 0.0020675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_618_94#_c_782_n 0.0130457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_618_94#_c_783_n 0.0231872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_618_94#_c_784_n 0.00541364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_618_94#_c_785_n 0.00177818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VPB N_B1_N_M1010_g 0.030081f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_73 VPB N_A_193_48#_M1001_g 0.0225109f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_193_48#_M1002_g 0.0215714f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_193_48#_M1007_g 0.021611f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_193_48#_M1011_g 0.0262604f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_193_48#_c_172_n 0.00952528f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_193_48#_c_173_n 0.00135978f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_193_48#_c_174_n 0.00331143f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_27_368#_M1017_g 0.0239076f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_27_368#_M1019_g 0.0215163f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.365
cc_82 VPB N_A_27_368#_c_319_n 0.0153183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_27_368#_c_320_n 0.0194384f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_27_368#_c_321_n 0.00236821f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_27_368#_c_322_n 0.0136968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_27_368#_c_314_n 0.00769959f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_27_368#_c_324_n 0.00723806f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_27_368#_c_315_n 0.00479174f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_27_368#_c_316_n 0.0443762f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A2_M1016_g 0.0217395f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_91 VPB N_A2_M1021_g 0.0217971f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.385
cc_92 VPB A2 0.0119519f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A2_c_408_n 0.013941f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A1_M1000_g 0.0241345f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_95 VPB N_A1_M1014_g 0.0356297f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.22
cc_96 VPB A1 0.00323349f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A1_c_465_n 0.0104768f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_529_n 0.00623005f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_530_n 0.00261656f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_531_n 0.00935698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_532_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_533_n 0.0515719f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_534_n 0.0189171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_535_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_536_n 0.0215473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_537_n 0.0387727f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_538_n 0.00708942f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_539_n 0.00601668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_540_n 0.017758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_541_n 0.0242507f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_542_n 0.00631788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_528_n 0.0688667f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_X_c_612_n 0.00585825f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB X 0.00146502f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_895_392#_c_658_n 0.00388794f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.385
cc_116 VPB N_A_895_392#_c_659_n 0.00196159f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.385
cc_117 VPB N_A_895_392#_c_660_n 0.00250912f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.365
cc_118 B1_N N_A_193_48#_M1003_g 0.00324428f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_119 N_B1_N_c_121_n N_A_193_48#_M1003_g 0.0212371f $X=0.59 $Y=1.385 $X2=0
+ $Y2=0
cc_120 N_B1_N_c_122_n N_A_193_48#_M1003_g 0.0168899f $X=0.585 $Y=1.22 $X2=0
+ $Y2=0
cc_121 N_B1_N_M1010_g N_A_193_48#_M1001_g 0.0434904f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_122 N_B1_N_c_122_n N_A_27_368#_c_312_n 0.00581235f $X=0.585 $Y=1.22 $X2=0
+ $Y2=0
cc_123 N_B1_N_M1010_g N_A_27_368#_c_319_n 0.00857168f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_124 N_B1_N_M1010_g N_A_27_368#_c_320_n 0.00754112f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_125 N_B1_N_M1010_g N_A_27_368#_c_330_n 0.014591f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_126 B1_N N_A_27_368#_c_313_n 0.00294872f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_127 N_B1_N_c_122_n N_A_27_368#_c_313_n 0.00232983f $X=0.585 $Y=1.22 $X2=0
+ $Y2=0
cc_128 N_B1_N_M1010_g N_A_27_368#_c_322_n 0.00497742f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_129 B1_N N_A_27_368#_c_322_n 0.00105488f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_130 B1_N N_A_27_368#_c_314_n 0.0284252f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_131 N_B1_N_c_121_n N_A_27_368#_c_314_n 0.0152991f $X=0.59 $Y=1.385 $X2=0
+ $Y2=0
cc_132 N_B1_N_c_122_n N_A_27_368#_c_314_n 0.00346495f $X=0.585 $Y=1.22 $X2=0
+ $Y2=0
cc_133 N_B1_N_M1010_g N_A_27_368#_c_324_n 4.64231e-19 $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_134 N_B1_N_M1010_g N_VPWR_c_529_n 0.00490247f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_135 N_B1_N_M1010_g N_VPWR_c_534_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_136 N_B1_N_M1010_g N_VPWR_c_528_n 0.00519477f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_137 N_B1_N_M1010_g X 0.00129836f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_138 N_B1_N_M1010_g N_X_c_615_n 0.00129375f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_139 B1_N N_X_c_611_n 0.0185939f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_140 N_B1_N_c_121_n N_X_c_611_n 2.26341e-19 $X=0.59 $Y=1.385 $X2=0 $Y2=0
cc_141 B1_N N_VGND_c_686_n 0.0160286f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_142 N_B1_N_c_121_n N_VGND_c_686_n 7.44677e-19 $X=0.59 $Y=1.385 $X2=0 $Y2=0
cc_143 N_B1_N_c_122_n N_VGND_c_686_n 0.00674192f $X=0.585 $Y=1.22 $X2=0 $Y2=0
cc_144 N_B1_N_c_122_n N_VGND_c_697_n 0.0082465f $X=0.585 $Y=1.22 $X2=0 $Y2=0
cc_145 N_B1_N_c_122_n N_VGND_c_698_n 0.00434272f $X=0.585 $Y=1.22 $X2=0 $Y2=0
cc_146 N_A_193_48#_c_174_n N_A_27_368#_M1017_g 0.00204674f $X=3.575 $Y=2.295
+ $X2=0 $Y2=0
cc_147 N_A_193_48#_c_161_n N_A_27_368#_M1008_g 0.00845542f $X=2.895 $Y=1.29
+ $X2=0 $Y2=0
cc_148 N_A_193_48#_c_162_n N_A_27_368#_M1008_g 0.00964849f $X=3.5 $Y=0.34 $X2=0
+ $Y2=0
cc_149 N_A_193_48#_c_164_n N_A_27_368#_M1008_g 0.0130363f $X=3.66 $Y=1.375 $X2=0
+ $Y2=0
cc_150 N_A_193_48#_c_183_p N_A_27_368#_M1008_g 0.00612159f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_151 N_A_193_48#_c_165_n N_A_27_368#_M1008_g 0.00364839f $X=3.745 $Y=1.95
+ $X2=0 $Y2=0
cc_152 N_A_193_48#_c_166_n N_A_27_368#_M1008_g 0.00518238f $X=2.895 $Y=1.455
+ $X2=0 $Y2=0
cc_153 N_A_193_48#_c_172_n N_A_27_368#_M1019_g 0.00994471f $X=4.975 $Y=2.125
+ $X2=0 $Y2=0
cc_154 N_A_193_48#_c_174_n N_A_27_368#_M1019_g 0.0204788f $X=3.575 $Y=2.295
+ $X2=0 $Y2=0
cc_155 N_A_193_48#_c_162_n N_A_27_368#_M1015_g 0.00312284f $X=3.5 $Y=0.34 $X2=0
+ $Y2=0
cc_156 N_A_193_48#_c_164_n N_A_27_368#_M1015_g 0.00586411f $X=3.66 $Y=1.375
+ $X2=0 $Y2=0
cc_157 N_A_193_48#_c_183_p N_A_27_368#_M1015_g 0.00621111f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_158 N_A_193_48#_c_165_n N_A_27_368#_M1015_g 0.00355214f $X=3.745 $Y=1.95
+ $X2=0 $Y2=0
cc_159 N_A_193_48#_M1001_g N_A_27_368#_c_320_n 5.75473e-19 $X=1.055 $Y=2.4 $X2=0
+ $Y2=0
cc_160 N_A_193_48#_M1001_g N_A_27_368#_c_330_n 0.0169849f $X=1.055 $Y=2.4 $X2=0
+ $Y2=0
cc_161 N_A_193_48#_M1002_g N_A_27_368#_c_330_n 0.0128378f $X=1.505 $Y=2.4 $X2=0
+ $Y2=0
cc_162 N_A_193_48#_M1007_g N_A_27_368#_c_330_n 0.0128378f $X=1.955 $Y=2.4 $X2=0
+ $Y2=0
cc_163 N_A_193_48#_M1011_g N_A_27_368#_c_330_n 0.0195354f $X=2.405 $Y=2.4 $X2=0
+ $Y2=0
cc_164 N_A_193_48#_M1011_g N_A_27_368#_c_321_n 0.0091007f $X=2.405 $Y=2.4 $X2=0
+ $Y2=0
cc_165 N_A_193_48#_c_174_n N_A_27_368#_c_321_n 0.00786728f $X=3.575 $Y=2.295
+ $X2=0 $Y2=0
cc_166 N_A_193_48#_M1001_g N_A_27_368#_c_322_n 0.00200273f $X=1.055 $Y=2.4 $X2=0
+ $Y2=0
cc_167 N_A_193_48#_M1011_g N_A_27_368#_c_315_n 0.00510089f $X=2.405 $Y=2.4 $X2=0
+ $Y2=0
cc_168 N_A_193_48#_c_164_n N_A_27_368#_c_315_n 0.025164f $X=3.66 $Y=1.375 $X2=0
+ $Y2=0
cc_169 N_A_193_48#_c_165_n N_A_27_368#_c_315_n 0.0229207f $X=3.745 $Y=1.95 $X2=0
+ $Y2=0
cc_170 N_A_193_48#_c_174_n N_A_27_368#_c_315_n 7.23724e-19 $X=3.575 $Y=2.295
+ $X2=0 $Y2=0
cc_171 N_A_193_48#_M1011_g N_A_27_368#_c_316_n 0.00412196f $X=2.405 $Y=2.4 $X2=0
+ $Y2=0
cc_172 N_A_193_48#_c_164_n N_A_27_368#_c_316_n 0.00665415f $X=3.66 $Y=1.375
+ $X2=0 $Y2=0
cc_173 N_A_193_48#_c_165_n N_A_27_368#_c_316_n 0.0148328f $X=3.745 $Y=1.95 $X2=0
+ $Y2=0
cc_174 N_A_193_48#_c_172_n N_A_27_368#_c_316_n 0.00593065f $X=4.975 $Y=2.125
+ $X2=0 $Y2=0
cc_175 N_A_193_48#_c_174_n N_A_27_368#_c_316_n 0.00334127f $X=3.575 $Y=2.295
+ $X2=0 $Y2=0
cc_176 N_A_193_48#_c_172_n N_A2_M1016_g 0.0183947f $X=4.975 $Y=2.125 $X2=0 $Y2=0
cc_177 N_A_193_48#_c_172_n A2 0.00996521f $X=4.975 $Y=2.125 $X2=0 $Y2=0
cc_178 N_A_193_48#_c_173_n A2 0.0143383f $X=5.06 $Y=2.3 $X2=0 $Y2=0
cc_179 N_A_193_48#_c_173_n N_A2_c_408_n 0.00221493f $X=5.06 $Y=2.3 $X2=0 $Y2=0
cc_180 N_A_193_48#_c_165_n N_A1_M1000_g 8.94991e-19 $X=3.745 $Y=1.95 $X2=0 $Y2=0
cc_181 N_A_193_48#_c_172_n N_A1_M1000_g 0.0254117f $X=4.975 $Y=2.125 $X2=0 $Y2=0
cc_182 N_A_193_48#_c_174_n N_A1_M1000_g 8.13122e-19 $X=3.575 $Y=2.295 $X2=0
+ $Y2=0
cc_183 N_A_193_48#_c_162_n N_A1_M1006_g 0.00179591f $X=3.5 $Y=0.34 $X2=0 $Y2=0
cc_184 N_A_193_48#_c_164_n N_A1_M1006_g 7.47639e-19 $X=3.66 $Y=1.375 $X2=0 $Y2=0
cc_185 N_A_193_48#_c_183_p N_A1_M1006_g 6.35849e-19 $X=3.665 $Y=0.615 $X2=0
+ $Y2=0
cc_186 N_A_193_48#_c_164_n A1 4.2002e-19 $X=3.66 $Y=1.375 $X2=0 $Y2=0
cc_187 N_A_193_48#_c_165_n A1 0.013357f $X=3.745 $Y=1.95 $X2=0 $Y2=0
cc_188 N_A_193_48#_c_172_n A1 0.039715f $X=4.975 $Y=2.125 $X2=0 $Y2=0
cc_189 N_A_193_48#_c_165_n N_A1_c_465_n 3.39653e-19 $X=3.745 $Y=1.95 $X2=0 $Y2=0
cc_190 N_A_193_48#_c_172_n N_A1_c_465_n 0.00342255f $X=4.975 $Y=2.125 $X2=0
+ $Y2=0
cc_191 N_A_193_48#_c_172_n N_VPWR_M1019_s 0.00400726f $X=4.975 $Y=2.125 $X2=0
+ $Y2=0
cc_192 N_A_193_48#_M1001_g N_VPWR_c_529_n 0.00957198f $X=1.055 $Y=2.4 $X2=0
+ $Y2=0
cc_193 N_A_193_48#_M1002_g N_VPWR_c_529_n 0.00105272f $X=1.505 $Y=2.4 $X2=0
+ $Y2=0
cc_194 N_A_193_48#_M1001_g N_VPWR_c_530_n 0.00105361f $X=1.055 $Y=2.4 $X2=0
+ $Y2=0
cc_195 N_A_193_48#_M1002_g N_VPWR_c_530_n 0.00937886f $X=1.505 $Y=2.4 $X2=0
+ $Y2=0
cc_196 N_A_193_48#_M1007_g N_VPWR_c_530_n 0.00935677f $X=1.955 $Y=2.4 $X2=0
+ $Y2=0
cc_197 N_A_193_48#_M1011_g N_VPWR_c_530_n 0.00105503f $X=2.405 $Y=2.4 $X2=0
+ $Y2=0
cc_198 N_A_193_48#_c_172_n N_VPWR_c_531_n 0.024886f $X=4.975 $Y=2.125 $X2=0
+ $Y2=0
cc_199 N_A_193_48#_c_174_n N_VPWR_c_531_n 0.0164809f $X=3.575 $Y=2.295 $X2=0
+ $Y2=0
cc_200 N_A_193_48#_M1001_g N_VPWR_c_535_n 0.00460063f $X=1.055 $Y=2.4 $X2=0
+ $Y2=0
cc_201 N_A_193_48#_M1002_g N_VPWR_c_535_n 0.00460063f $X=1.505 $Y=2.4 $X2=0
+ $Y2=0
cc_202 N_A_193_48#_c_174_n N_VPWR_c_536_n 0.0109793f $X=3.575 $Y=2.295 $X2=0
+ $Y2=0
cc_203 N_A_193_48#_M1007_g N_VPWR_c_540_n 0.00460063f $X=1.955 $Y=2.4 $X2=0
+ $Y2=0
cc_204 N_A_193_48#_M1011_g N_VPWR_c_540_n 0.00460063f $X=2.405 $Y=2.4 $X2=0
+ $Y2=0
cc_205 N_A_193_48#_M1007_g N_VPWR_c_541_n 0.00104752f $X=1.955 $Y=2.4 $X2=0
+ $Y2=0
cc_206 N_A_193_48#_M1011_g N_VPWR_c_541_n 0.0109968f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_207 N_A_193_48#_c_174_n N_VPWR_c_541_n 0.00114658f $X=3.575 $Y=2.295 $X2=0
+ $Y2=0
cc_208 N_A_193_48#_M1001_g N_VPWR_c_528_n 0.00443247f $X=1.055 $Y=2.4 $X2=0
+ $Y2=0
cc_209 N_A_193_48#_M1002_g N_VPWR_c_528_n 0.00443247f $X=1.505 $Y=2.4 $X2=0
+ $Y2=0
cc_210 N_A_193_48#_M1007_g N_VPWR_c_528_n 0.00443247f $X=1.955 $Y=2.4 $X2=0
+ $Y2=0
cc_211 N_A_193_48#_M1011_g N_VPWR_c_528_n 0.00441691f $X=2.405 $Y=2.4 $X2=0
+ $Y2=0
cc_212 N_A_193_48#_c_174_n N_VPWR_c_528_n 0.00901959f $X=3.575 $Y=2.295 $X2=0
+ $Y2=0
cc_213 N_A_193_48#_M1003_g N_X_c_606_n 3.77529e-19 $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A_193_48#_M1005_g N_X_c_606_n 0.00305913f $X=1.48 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A_193_48#_M1002_g N_X_c_612_n 0.0192011f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_216 N_A_193_48#_M1007_g N_X_c_612_n 0.0168661f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_217 N_A_193_48#_M1011_g N_X_c_612_n 0.0201589f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_218 N_A_193_48#_c_160_n N_X_c_612_n 0.0598377f $X=2.81 $Y=1.455 $X2=0 $Y2=0
cc_219 N_A_193_48#_c_167_n N_X_c_612_n 0.00843661f $X=2.34 $Y=1.455 $X2=0 $Y2=0
cc_220 N_A_193_48#_M1005_g N_X_c_607_n 0.0147259f $X=1.48 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A_193_48#_M1013_g N_X_c_607_n 0.0119326f $X=1.91 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A_193_48#_c_160_n N_X_c_607_n 0.0559114f $X=2.81 $Y=1.455 $X2=0 $Y2=0
cc_223 N_A_193_48#_c_167_n N_X_c_607_n 0.00496587f $X=2.34 $Y=1.455 $X2=0 $Y2=0
cc_224 N_A_193_48#_M1005_g N_X_c_608_n 6.66379e-19 $X=1.48 $Y=0.74 $X2=0 $Y2=0
cc_225 N_A_193_48#_M1013_g N_X_c_608_n 0.00849619f $X=1.91 $Y=0.74 $X2=0 $Y2=0
cc_226 N_A_193_48#_M1018_g N_X_c_608_n 3.55395e-19 $X=2.34 $Y=0.74 $X2=0 $Y2=0
cc_227 N_A_193_48#_M1003_g N_X_c_609_n 2.99553e-19 $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A_193_48#_M1001_g X 0.00793524f $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_229 N_A_193_48#_M1002_g X 0.00474284f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_230 N_A_193_48#_c_167_n X 0.00760965f $X=2.34 $Y=1.455 $X2=0 $Y2=0
cc_231 N_A_193_48#_M1001_g N_X_c_615_n 0.0102814f $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_232 N_A_193_48#_M1003_g N_X_c_611_n 0.00252852f $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A_193_48#_M1005_g N_X_c_611_n 0.0038796f $X=1.48 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A_193_48#_c_160_n N_X_c_611_n 0.0253315f $X=2.81 $Y=1.455 $X2=0 $Y2=0
cc_235 N_A_193_48#_c_167_n N_X_c_611_n 0.0134482f $X=2.34 $Y=1.455 $X2=0 $Y2=0
cc_236 N_A_193_48#_c_172_n N_A_895_392#_M1000_s 0.00169557f $X=4.975 $Y=2.125
+ $X2=-0.19 $Y2=-0.245
cc_237 N_A_193_48#_c_172_n N_A_895_392#_c_662_n 0.0177444f $X=4.975 $Y=2.125
+ $X2=0 $Y2=0
cc_238 N_A_193_48#_M1016_d N_A_895_392#_c_658_n 0.00165831f $X=4.925 $Y=1.96
+ $X2=0 $Y2=0
cc_239 N_A_193_48#_c_172_n N_A_895_392#_c_658_n 0.0037387f $X=4.975 $Y=2.125
+ $X2=0 $Y2=0
cc_240 N_A_193_48#_c_273_p N_A_895_392#_c_658_n 0.0118736f $X=5.06 $Y=2.57 $X2=0
+ $Y2=0
cc_241 N_A_193_48#_c_173_n N_A_895_392#_c_660_n 0.0119511f $X=5.06 $Y=2.3 $X2=0
+ $Y2=0
cc_242 N_A_193_48#_M1003_g N_VGND_c_686_n 0.0105578f $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_243 N_A_193_48#_M1005_g N_VGND_c_686_n 4.79292e-19 $X=1.48 $Y=0.74 $X2=0
+ $Y2=0
cc_244 N_A_193_48#_M1003_g N_VGND_c_687_n 4.62568e-19 $X=1.04 $Y=0.74 $X2=0
+ $Y2=0
cc_245 N_A_193_48#_M1005_g N_VGND_c_687_n 0.00870114f $X=1.48 $Y=0.74 $X2=0
+ $Y2=0
cc_246 N_A_193_48#_M1013_g N_VGND_c_687_n 0.00167001f $X=1.91 $Y=0.74 $X2=0
+ $Y2=0
cc_247 N_A_193_48#_M1013_g N_VGND_c_688_n 6.04497e-19 $X=1.91 $Y=0.74 $X2=0
+ $Y2=0
cc_248 N_A_193_48#_M1018_g N_VGND_c_688_n 0.014379f $X=2.34 $Y=0.74 $X2=0 $Y2=0
cc_249 N_A_193_48#_c_160_n N_VGND_c_688_n 0.0214009f $X=2.81 $Y=1.455 $X2=0
+ $Y2=0
cc_250 N_A_193_48#_c_161_n N_VGND_c_688_n 0.0528834f $X=2.895 $Y=1.29 $X2=0
+ $Y2=0
cc_251 N_A_193_48#_c_163_n N_VGND_c_688_n 0.0146661f $X=2.98 $Y=0.34 $X2=0 $Y2=0
cc_252 N_A_193_48#_c_167_n N_VGND_c_688_n 0.00217919f $X=2.34 $Y=1.455 $X2=0
+ $Y2=0
cc_253 N_A_193_48#_c_162_n N_VGND_c_689_n 0.00519468f $X=3.5 $Y=0.34 $X2=0 $Y2=0
cc_254 N_A_193_48#_c_183_p N_VGND_c_689_n 0.00482934f $X=3.665 $Y=0.615 $X2=0
+ $Y2=0
cc_255 N_A_193_48#_M1013_g N_VGND_c_691_n 0.00434272f $X=1.91 $Y=0.74 $X2=0
+ $Y2=0
cc_256 N_A_193_48#_M1018_g N_VGND_c_691_n 0.00383152f $X=2.34 $Y=0.74 $X2=0
+ $Y2=0
cc_257 N_A_193_48#_M1003_g N_VGND_c_693_n 0.00429299f $X=1.04 $Y=0.74 $X2=0
+ $Y2=0
cc_258 N_A_193_48#_M1005_g N_VGND_c_693_n 0.00383152f $X=1.48 $Y=0.74 $X2=0
+ $Y2=0
cc_259 N_A_193_48#_c_162_n N_VGND_c_694_n 0.0566428f $X=3.5 $Y=0.34 $X2=0 $Y2=0
cc_260 N_A_193_48#_c_163_n N_VGND_c_694_n 0.0121867f $X=2.98 $Y=0.34 $X2=0 $Y2=0
cc_261 N_A_193_48#_M1003_g N_VGND_c_697_n 0.00847623f $X=1.04 $Y=0.74 $X2=0
+ $Y2=0
cc_262 N_A_193_48#_M1005_g N_VGND_c_697_n 0.0075764f $X=1.48 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A_193_48#_M1013_g N_VGND_c_697_n 0.00820284f $X=1.91 $Y=0.74 $X2=0
+ $Y2=0
cc_264 N_A_193_48#_M1018_g N_VGND_c_697_n 0.0075754f $X=2.34 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A_193_48#_c_162_n N_VGND_c_697_n 0.0322874f $X=3.5 $Y=0.34 $X2=0 $Y2=0
cc_266 N_A_193_48#_c_163_n N_VGND_c_697_n 0.00660921f $X=2.98 $Y=0.34 $X2=0
+ $Y2=0
cc_267 N_A_193_48#_c_161_n N_A_618_94#_c_786_n 0.0262213f $X=2.895 $Y=1.29 $X2=0
+ $Y2=0
cc_268 N_A_193_48#_c_162_n N_A_618_94#_c_786_n 0.0127218f $X=3.5 $Y=0.34 $X2=0
+ $Y2=0
cc_269 N_A_193_48#_M1008_d N_A_618_94#_c_777_n 0.00176461f $X=3.525 $Y=0.47
+ $X2=0 $Y2=0
cc_270 N_A_193_48#_c_162_n N_A_618_94#_c_777_n 0.0042894f $X=3.5 $Y=0.34 $X2=0
+ $Y2=0
cc_271 N_A_193_48#_c_164_n N_A_618_94#_c_777_n 0.03855f $X=3.66 $Y=1.375 $X2=0
+ $Y2=0
cc_272 N_A_193_48#_c_183_p N_A_618_94#_c_777_n 0.0167224f $X=3.665 $Y=0.615
+ $X2=0 $Y2=0
cc_273 N_A_193_48#_c_161_n N_A_618_94#_c_778_n 0.0140746f $X=2.895 $Y=1.29 $X2=0
+ $Y2=0
cc_274 N_A_193_48#_c_164_n N_A_618_94#_c_778_n 0.0140592f $X=3.66 $Y=1.375 $X2=0
+ $Y2=0
cc_275 N_A_193_48#_c_172_n N_A_618_94#_c_780_n 0.00462538f $X=4.975 $Y=2.125
+ $X2=0 $Y2=0
cc_276 N_A_193_48#_c_172_n N_A_618_94#_c_784_n 0.00590868f $X=4.975 $Y=2.125
+ $X2=0 $Y2=0
cc_277 N_A_27_368#_c_316_n N_A1_M1000_g 0.0298672f $X=3.8 $Y=1.795 $X2=0 $Y2=0
cc_278 N_A_27_368#_M1015_g N_A1_M1006_g 0.0285527f $X=3.88 $Y=0.79 $X2=0 $Y2=0
cc_279 N_A_27_368#_M1015_g A1 0.00126428f $X=3.88 $Y=0.79 $X2=0 $Y2=0
cc_280 N_A_27_368#_M1015_g N_A1_c_465_n 0.0195598f $X=3.88 $Y=0.79 $X2=0 $Y2=0
cc_281 N_A_27_368#_c_330_n N_VPWR_M1010_d 0.0125285f $X=3.15 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_282 N_A_27_368#_c_330_n N_VPWR_M1002_s 0.00328796f $X=3.15 $Y=2.475 $X2=0
+ $Y2=0
cc_283 N_A_27_368#_c_330_n N_VPWR_M1011_s 0.033344f $X=3.15 $Y=2.475 $X2=0 $Y2=0
cc_284 N_A_27_368#_c_321_n N_VPWR_M1011_s 0.0047109f $X=3.235 $Y=2.39 $X2=0
+ $Y2=0
cc_285 N_A_27_368#_c_320_n N_VPWR_c_529_n 0.0103139f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_286 N_A_27_368#_c_330_n N_VPWR_c_529_n 0.022352f $X=3.15 $Y=2.475 $X2=0 $Y2=0
cc_287 N_A_27_368#_c_330_n N_VPWR_c_530_n 0.0165487f $X=3.15 $Y=2.475 $X2=0
+ $Y2=0
cc_288 N_A_27_368#_M1019_g N_VPWR_c_531_n 0.00629617f $X=3.8 $Y=2.54 $X2=0 $Y2=0
cc_289 N_A_27_368#_c_320_n N_VPWR_c_534_n 0.0158876f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_290 N_A_27_368#_M1017_g N_VPWR_c_536_n 0.00553757f $X=3.35 $Y=2.54 $X2=0
+ $Y2=0
cc_291 N_A_27_368#_M1019_g N_VPWR_c_536_n 0.005209f $X=3.8 $Y=2.54 $X2=0 $Y2=0
cc_292 N_A_27_368#_M1017_g N_VPWR_c_541_n 0.0102576f $X=3.35 $Y=2.54 $X2=0 $Y2=0
cc_293 N_A_27_368#_c_330_n N_VPWR_c_541_n 0.053712f $X=3.15 $Y=2.475 $X2=0 $Y2=0
cc_294 N_A_27_368#_M1017_g N_VPWR_c_528_n 0.0090889f $X=3.35 $Y=2.54 $X2=0 $Y2=0
cc_295 N_A_27_368#_M1019_g N_VPWR_c_528_n 0.0098363f $X=3.8 $Y=2.54 $X2=0 $Y2=0
cc_296 N_A_27_368#_c_320_n N_VPWR_c_528_n 0.0130823f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_297 N_A_27_368#_c_330_n N_VPWR_c_528_n 0.0522363f $X=3.15 $Y=2.475 $X2=0
+ $Y2=0
cc_298 N_A_27_368#_c_330_n N_X_M1001_d 0.00460584f $X=3.15 $Y=2.475 $X2=0 $Y2=0
cc_299 N_A_27_368#_c_330_n N_X_M1007_d 0.00460877f $X=3.15 $Y=2.475 $X2=0 $Y2=0
cc_300 N_A_27_368#_c_330_n N_X_c_612_n 0.0557909f $X=3.15 $Y=2.475 $X2=0 $Y2=0
cc_301 N_A_27_368#_c_330_n N_X_c_615_n 0.0137163f $X=3.15 $Y=2.475 $X2=0 $Y2=0
cc_302 N_A_27_368#_c_322_n N_X_c_615_n 0.0106105f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_303 N_A_27_368#_c_312_n N_VGND_c_686_n 0.026158f $X=0.31 $Y=0.515 $X2=0 $Y2=0
cc_304 N_A_27_368#_M1008_g N_VGND_c_694_n 7.82275e-19 $X=3.45 $Y=0.79 $X2=0
+ $Y2=0
cc_305 N_A_27_368#_M1015_g N_VGND_c_694_n 0.00435309f $X=3.88 $Y=0.79 $X2=0
+ $Y2=0
cc_306 N_A_27_368#_M1015_g N_VGND_c_697_n 0.00428698f $X=3.88 $Y=0.79 $X2=0
+ $Y2=0
cc_307 N_A_27_368#_c_312_n N_VGND_c_697_n 0.0142062f $X=0.31 $Y=0.515 $X2=0
+ $Y2=0
cc_308 N_A_27_368#_c_312_n N_VGND_c_698_n 0.0172202f $X=0.31 $Y=0.515 $X2=0
+ $Y2=0
cc_309 N_A_27_368#_M1008_g N_A_618_94#_c_777_n 0.0111584f $X=3.45 $Y=0.79 $X2=0
+ $Y2=0
cc_310 N_A_27_368#_M1015_g N_A_618_94#_c_777_n 0.0167517f $X=3.88 $Y=0.79 $X2=0
+ $Y2=0
cc_311 N_A_27_368#_c_316_n N_A_618_94#_c_777_n 2.52421e-19 $X=3.8 $Y=1.795 $X2=0
+ $Y2=0
cc_312 N_A_27_368#_M1015_g N_A_618_94#_c_784_n 0.00501111f $X=3.88 $Y=0.79 $X2=0
+ $Y2=0
cc_313 N_A2_M1016_g N_A1_M1000_g 0.0449432f $X=4.835 $Y=2.46 $X2=0 $Y2=0
cc_314 N_A2_M1004_g N_A1_M1006_g 0.0248487f $X=4.88 $Y=0.945 $X2=0 $Y2=0
cc_315 N_A2_M1004_g N_A1_c_459_n 0.00895007f $X=4.88 $Y=0.945 $X2=0 $Y2=0
cc_316 N_A2_M1009_g N_A1_c_459_n 0.00894529f $X=5.31 $Y=0.945 $X2=0 $Y2=0
cc_317 N_A2_M1009_g N_A1_c_461_n 0.00674476f $X=5.31 $Y=0.945 $X2=0 $Y2=0
cc_318 A2 N_A1_M1014_g 0.025748f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_319 N_A2_c_408_n N_A1_M1014_g 0.031121f $X=5.285 $Y=1.615 $X2=0 $Y2=0
cc_320 N_A2_M1009_g N_A1_M1012_g 0.0218553f $X=5.31 $Y=0.945 $X2=0 $Y2=0
cc_321 A2 A1 0.0285452f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_322 N_A2_c_408_n A1 0.00274698f $X=5.285 $Y=1.615 $X2=0 $Y2=0
cc_323 A2 N_A1_c_465_n 2.60921e-19 $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_324 N_A2_c_408_n N_A1_c_465_n 0.0180311f $X=5.285 $Y=1.615 $X2=0 $Y2=0
cc_325 A2 N_VPWR_c_533_n 0.0211423f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_326 N_A2_M1016_g N_VPWR_c_537_n 0.00333896f $X=4.835 $Y=2.46 $X2=0 $Y2=0
cc_327 N_A2_M1021_g N_VPWR_c_537_n 0.00333896f $X=5.285 $Y=2.46 $X2=0 $Y2=0
cc_328 N_A2_M1016_g N_VPWR_c_528_n 0.00422796f $X=4.835 $Y=2.46 $X2=0 $Y2=0
cc_329 N_A2_M1021_g N_VPWR_c_528_n 0.00422796f $X=5.285 $Y=2.46 $X2=0 $Y2=0
cc_330 N_A2_M1016_g N_A_895_392#_c_662_n 0.00763409f $X=4.835 $Y=2.46 $X2=0
+ $Y2=0
cc_331 N_A2_M1021_g N_A_895_392#_c_662_n 5.16131e-19 $X=5.285 $Y=2.46 $X2=0
+ $Y2=0
cc_332 N_A2_M1016_g N_A_895_392#_c_658_n 0.00912855f $X=4.835 $Y=2.46 $X2=0
+ $Y2=0
cc_333 N_A2_M1021_g N_A_895_392#_c_658_n 0.0135505f $X=5.285 $Y=2.46 $X2=0 $Y2=0
cc_334 N_A2_M1016_g N_A_895_392#_c_659_n 0.00255139f $X=4.835 $Y=2.46 $X2=0
+ $Y2=0
cc_335 N_A2_M1016_g N_A_895_392#_c_660_n 6.83508e-19 $X=4.835 $Y=2.46 $X2=0
+ $Y2=0
cc_336 N_A2_M1021_g N_A_895_392#_c_660_n 0.0130557f $X=5.285 $Y=2.46 $X2=0 $Y2=0
cc_337 A2 N_A_895_392#_c_660_n 0.0285144f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_338 N_A2_M1004_g N_VGND_c_689_n 0.0017139f $X=4.88 $Y=0.945 $X2=0 $Y2=0
cc_339 N_A2_M1004_g N_VGND_c_690_n 4.44858e-19 $X=4.88 $Y=0.945 $X2=0 $Y2=0
cc_340 N_A2_M1009_g N_VGND_c_690_n 0.00728275f $X=5.31 $Y=0.945 $X2=0 $Y2=0
cc_341 N_A2_M1004_g N_VGND_c_697_n 9.49986e-19 $X=4.88 $Y=0.945 $X2=0 $Y2=0
cc_342 N_A2_M1009_g N_VGND_c_697_n 7.97988e-19 $X=5.31 $Y=0.945 $X2=0 $Y2=0
cc_343 N_A2_M1004_g N_A_618_94#_c_779_n 5.46534e-19 $X=4.88 $Y=0.945 $X2=0 $Y2=0
cc_344 N_A2_M1004_g N_A_618_94#_c_780_n 0.0118831f $X=4.88 $Y=0.945 $X2=0 $Y2=0
cc_345 A2 N_A_618_94#_c_780_n 0.00603618f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_346 N_A2_c_408_n N_A_618_94#_c_780_n 0.00187709f $X=5.285 $Y=1.615 $X2=0
+ $Y2=0
cc_347 N_A2_M1004_g N_A_618_94#_c_781_n 0.00720634f $X=4.88 $Y=0.945 $X2=0 $Y2=0
cc_348 N_A2_M1009_g N_A_618_94#_c_782_n 0.0121744f $X=5.31 $Y=0.945 $X2=0 $Y2=0
cc_349 A2 N_A_618_94#_c_782_n 0.0742946f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_350 N_A2_M1009_g N_A_618_94#_c_783_n 5.70901e-19 $X=5.31 $Y=0.945 $X2=0 $Y2=0
cc_351 N_A2_M1004_g N_A_618_94#_c_785_n 9.00612e-19 $X=4.88 $Y=0.945 $X2=0 $Y2=0
cc_352 A2 N_A_618_94#_c_785_n 0.0209604f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_353 N_A2_c_408_n N_A_618_94#_c_785_n 0.00248288f $X=5.285 $Y=1.615 $X2=0
+ $Y2=0
cc_354 N_A1_M1000_g N_VPWR_c_531_n 0.00240654f $X=4.385 $Y=2.46 $X2=0 $Y2=0
cc_355 N_A1_M1014_g N_VPWR_c_533_n 0.00353586f $X=5.735 $Y=2.46 $X2=0 $Y2=0
cc_356 N_A1_M1000_g N_VPWR_c_537_n 0.00517089f $X=4.385 $Y=2.46 $X2=0 $Y2=0
cc_357 N_A1_M1014_g N_VPWR_c_537_n 0.00517089f $X=5.735 $Y=2.46 $X2=0 $Y2=0
cc_358 N_A1_M1000_g N_VPWR_c_528_n 0.00978168f $X=4.385 $Y=2.46 $X2=0 $Y2=0
cc_359 N_A1_M1014_g N_VPWR_c_528_n 0.0098133f $X=5.735 $Y=2.46 $X2=0 $Y2=0
cc_360 N_A1_M1000_g N_A_895_392#_c_662_n 0.00619441f $X=4.385 $Y=2.46 $X2=0
+ $Y2=0
cc_361 N_A1_M1014_g N_A_895_392#_c_658_n 0.00358808f $X=5.735 $Y=2.46 $X2=0
+ $Y2=0
cc_362 N_A1_M1000_g N_A_895_392#_c_659_n 0.00403165f $X=4.385 $Y=2.46 $X2=0
+ $Y2=0
cc_363 N_A1_M1014_g N_A_895_392#_c_660_n 0.01247f $X=5.735 $Y=2.46 $X2=0 $Y2=0
cc_364 N_A1_M1006_g N_VGND_c_689_n 0.0104443f $X=4.38 $Y=0.945 $X2=0 $Y2=0
cc_365 N_A1_c_459_n N_VGND_c_689_n 0.0190951f $X=5.665 $Y=0.18 $X2=0 $Y2=0
cc_366 N_A1_c_459_n N_VGND_c_690_n 0.0190272f $X=5.665 $Y=0.18 $X2=0 $Y2=0
cc_367 N_A1_M1012_g N_VGND_c_690_n 0.012705f $X=5.74 $Y=0.945 $X2=0 $Y2=0
cc_368 N_A1_c_460_n N_VGND_c_694_n 0.00730708f $X=4.455 $Y=0.18 $X2=0 $Y2=0
cc_369 N_A1_c_459_n N_VGND_c_695_n 0.0187698f $X=5.665 $Y=0.18 $X2=0 $Y2=0
cc_370 N_A1_c_459_n N_VGND_c_696_n 0.00769733f $X=5.665 $Y=0.18 $X2=0 $Y2=0
cc_371 N_A1_c_459_n N_VGND_c_697_n 0.0364405f $X=5.665 $Y=0.18 $X2=0 $Y2=0
cc_372 N_A1_c_460_n N_VGND_c_697_n 0.0106516f $X=4.455 $Y=0.18 $X2=0 $Y2=0
cc_373 N_A1_M1006_g N_A_618_94#_c_779_n 0.00490618f $X=4.38 $Y=0.945 $X2=0 $Y2=0
cc_374 N_A1_M1006_g N_A_618_94#_c_780_n 0.0120608f $X=4.38 $Y=0.945 $X2=0 $Y2=0
cc_375 A1 N_A_618_94#_c_780_n 0.0261629f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_376 N_A1_c_465_n N_A_618_94#_c_780_n 0.00119983f $X=4.34 $Y=1.615 $X2=0 $Y2=0
cc_377 N_A1_M1006_g N_A_618_94#_c_781_n 6.06182e-19 $X=4.38 $Y=0.945 $X2=0 $Y2=0
cc_378 N_A1_c_459_n N_A_618_94#_c_781_n 0.00449787f $X=5.665 $Y=0.18 $X2=0 $Y2=0
cc_379 N_A1_c_461_n N_A_618_94#_c_782_n 9.10293e-19 $X=5.735 $Y=1.43 $X2=0 $Y2=0
cc_380 N_A1_M1012_g N_A_618_94#_c_782_n 0.0121208f $X=5.74 $Y=0.945 $X2=0 $Y2=0
cc_381 N_A1_M1012_g N_A_618_94#_c_783_n 0.00753506f $X=5.74 $Y=0.945 $X2=0 $Y2=0
cc_382 N_A1_M1006_g N_A_618_94#_c_784_n 0.00691928f $X=4.38 $Y=0.945 $X2=0 $Y2=0
cc_383 A1 N_A_618_94#_c_784_n 0.0128713f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_384 N_A1_c_465_n N_A_618_94#_c_784_n 0.00306209f $X=4.34 $Y=1.615 $X2=0 $Y2=0
cc_385 N_VPWR_M1002_s N_X_c_612_n 0.00170669f $X=1.595 $Y=1.84 $X2=0 $Y2=0
cc_386 N_VPWR_c_533_n N_A_895_392#_c_658_n 0.0103534f $X=5.96 $Y=2.115 $X2=0
+ $Y2=0
cc_387 N_VPWR_c_537_n N_A_895_392#_c_658_n 0.0592384f $X=5.875 $Y=3.33 $X2=0
+ $Y2=0
cc_388 N_VPWR_c_528_n N_A_895_392#_c_658_n 0.0326137f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_389 N_VPWR_c_531_n N_A_895_392#_c_659_n 0.0119238f $X=4.11 $Y=2.635 $X2=0
+ $Y2=0
cc_390 N_VPWR_c_537_n N_A_895_392#_c_659_n 0.0232421f $X=5.875 $Y=3.33 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_528_n N_A_895_392#_c_659_n 0.0125162f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_392 N_VPWR_c_533_n N_A_895_392#_c_660_n 0.0317501f $X=5.96 $Y=2.115 $X2=0
+ $Y2=0
cc_393 N_VPWR_c_533_n N_A_618_94#_c_782_n 3.21367e-19 $X=5.96 $Y=2.115 $X2=0
+ $Y2=0
cc_394 N_X_c_607_n N_VGND_M1005_d 0.00176461f $X=1.96 $Y=1.035 $X2=0 $Y2=0
cc_395 N_X_c_606_n N_VGND_c_686_n 0.0232433f $X=1.255 $Y=0.515 $X2=0 $Y2=0
cc_396 N_X_c_606_n N_VGND_c_687_n 0.0288482f $X=1.255 $Y=0.515 $X2=0 $Y2=0
cc_397 N_X_c_607_n N_VGND_c_687_n 0.0153337f $X=1.96 $Y=1.035 $X2=0 $Y2=0
cc_398 N_X_c_608_n N_VGND_c_687_n 0.0154978f $X=2.125 $Y=0.515 $X2=0 $Y2=0
cc_399 N_X_c_607_n N_VGND_c_688_n 0.00626822f $X=1.96 $Y=1.035 $X2=0 $Y2=0
cc_400 N_X_c_608_n N_VGND_c_688_n 0.021337f $X=2.125 $Y=0.515 $X2=0 $Y2=0
cc_401 N_X_c_608_n N_VGND_c_691_n 0.0109942f $X=2.125 $Y=0.515 $X2=0 $Y2=0
cc_402 N_X_c_606_n N_VGND_c_693_n 0.00861184f $X=1.255 $Y=0.515 $X2=0 $Y2=0
cc_403 N_X_c_606_n N_VGND_c_697_n 0.00712813f $X=1.255 $Y=0.515 $X2=0 $Y2=0
cc_404 N_X_c_608_n N_VGND_c_697_n 0.00904371f $X=2.125 $Y=0.515 $X2=0 $Y2=0
cc_405 N_VGND_c_689_n N_A_618_94#_c_779_n 0.013328f $X=4.665 $Y=0.77 $X2=0 $Y2=0
cc_406 N_VGND_c_694_n N_A_618_94#_c_779_n 0.00670736f $X=4.5 $Y=0 $X2=0 $Y2=0
cc_407 N_VGND_c_697_n N_A_618_94#_c_779_n 0.0100487f $X=6 $Y=0 $X2=0 $Y2=0
cc_408 N_VGND_M1006_s N_A_618_94#_c_780_n 0.00250873f $X=4.455 $Y=0.625 $X2=0
+ $Y2=0
cc_409 N_VGND_c_689_n N_A_618_94#_c_780_n 0.0192006f $X=4.665 $Y=0.77 $X2=0
+ $Y2=0
cc_410 N_VGND_c_689_n N_A_618_94#_c_781_n 0.0122347f $X=4.665 $Y=0.77 $X2=0
+ $Y2=0
cc_411 N_VGND_c_690_n N_A_618_94#_c_781_n 0.0122347f $X=5.525 $Y=0.77 $X2=0
+ $Y2=0
cc_412 N_VGND_c_695_n N_A_618_94#_c_781_n 0.00528395f $X=5.36 $Y=0 $X2=0 $Y2=0
cc_413 N_VGND_c_697_n N_A_618_94#_c_781_n 0.00668313f $X=6 $Y=0 $X2=0 $Y2=0
cc_414 N_VGND_M1009_d N_A_618_94#_c_782_n 0.00176461f $X=5.385 $Y=0.625 $X2=0
+ $Y2=0
cc_415 N_VGND_c_690_n N_A_618_94#_c_782_n 0.0152916f $X=5.525 $Y=0.77 $X2=0
+ $Y2=0
cc_416 N_VGND_c_690_n N_A_618_94#_c_783_n 0.0127625f $X=5.525 $Y=0.77 $X2=0
+ $Y2=0
cc_417 N_VGND_c_696_n N_A_618_94#_c_783_n 0.00712528f $X=6 $Y=0 $X2=0 $Y2=0
cc_418 N_VGND_c_697_n N_A_618_94#_c_783_n 0.0102037f $X=6 $Y=0 $X2=0 $Y2=0

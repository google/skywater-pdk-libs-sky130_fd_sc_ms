* File: sky130_fd_sc_ms__dlxbn_2.pex.spice
* Created: Fri Aug 28 17:28:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLXBN_2%D 3 7 9 12
c35 12 0 1.67694e-19 $X=0.605 $Y=1.615
c36 7 0 1.17509e-19 $X=0.59 $Y=2.54
r37 12 15 40.7727 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.595 $Y=1.615
+ $X2=0.595 $Y2=1.78
r38 12 14 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.595 $Y=1.615
+ $X2=0.595 $Y2=1.45
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.605
+ $Y=1.615 $X2=0.605 $Y2=1.615
r40 9 13 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.72 $Y=1.615
+ $X2=0.605 $Y2=1.615
r41 7 15 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=0.59 $Y=2.54 $X2=0.59
+ $Y2=1.78
r42 3 14 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.495 $Y=0.955
+ $X2=0.495 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_2%GATE_N 3 7 9 12 13
c37 13 0 9.5906e-20 $X=1.15 $Y=1.795
r38 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.795
+ $X2=1.15 $Y2=1.96
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.795
+ $X2=1.15 $Y2=1.63
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.795 $X2=1.15 $Y2=1.795
r41 9 13 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.15 $Y=2.035 $X2=1.15
+ $Y2=1.795
r42 7 14 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=1.085 $Y=0.86
+ $X2=1.085 $Y2=1.63
r43 3 15 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=1.09 $Y=2.54 $X2=1.09
+ $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_2%A_232_98# 1 2 7 11 15 17 18 20 21 22 24 27
+ 29 30 33 35 38 39 42 47 55 58 60 62
c148 60 0 1.87089e-19 $X=4.19 $Y=1.585
c149 58 0 3.16539e-20 $X=4.06 $Y=1.585
c150 47 0 7.17879e-20 $X=1.72 $Y=1.425
c151 35 0 1.17509e-19 $X=1.317 $Y=2.56
c152 18 0 1.8903e-19 $X=3.16 $Y=1.11
r153 66 68 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=3.73 $Y=1.585
+ $X2=3.995 $Y2=1.585
r154 58 68 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=4.06 $Y=1.585
+ $X2=3.995 $Y2=1.585
r155 57 60 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=4.06 $Y=1.585
+ $X2=4.19 $Y2=1.585
r156 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.06
+ $Y=1.585 $X2=4.06 $Y2=1.585
r157 54 55 5.07737 $w=2.38e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=2.44
+ $X2=1.655 $Y2=2.44
r158 48 62 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.72 $Y=1.425
+ $X2=1.72 $Y2=1.335
r159 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.72
+ $Y=1.425 $X2=1.72 $Y2=1.425
r160 45 47 6.52326 $w=2.63e-07 $l=1.5e-07 $layer=LI1_cond $X=1.57 $Y=1.392
+ $X2=1.72 $Y2=1.392
r161 41 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.19 $Y=1.75
+ $X2=4.19 $Y2=1.585
r162 41 42 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=4.19 $Y=1.75
+ $X2=4.19 $Y2=2.39
r163 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.105 $Y=2.475
+ $X2=4.19 $Y2=2.39
r164 39 55 159.84 $w=1.68e-07 $l=2.45e-06 $layer=LI1_cond $X=4.105 $Y=2.475
+ $X2=1.655 $Y2=2.475
r165 38 54 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.57 $Y=2.32
+ $X2=1.57 $Y2=2.44
r166 37 45 3.33486 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=1.57 $Y=1.525
+ $X2=1.57 $Y2=1.392
r167 37 38 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=1.57 $Y=1.525
+ $X2=1.57 $Y2=2.32
r168 35 54 12.1487 $w=2.38e-07 $l=2.53e-07 $layer=LI1_cond $X=1.317 $Y=2.44
+ $X2=1.57 $Y2=2.44
r169 35 51 0.0960369 $w=2.38e-07 $l=2e-09 $layer=LI1_cond $X=1.317 $Y=2.44
+ $X2=1.315 $Y2=2.44
r170 31 45 11.7419 $w=2.63e-07 $l=2.7e-07 $layer=LI1_cond $X=1.3 $Y=1.392
+ $X2=1.57 $Y2=1.392
r171 31 33 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=1.3 $Y=1.26
+ $X2=1.3 $Y2=1.085
r172 25 68 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=1.75
+ $X2=3.995 $Y2=1.585
r173 25 27 163.258 $w=1.8e-07 $l=4.2e-07 $layer=POLY_cond $X=3.995 $Y=1.75
+ $X2=3.995 $Y2=2.17
r174 24 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=1.42
+ $X2=3.73 $Y2=1.585
r175 23 24 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=3.73 $Y=1.26
+ $X2=3.73 $Y2=1.42
r176 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.655 $Y=1.185
+ $X2=3.73 $Y2=1.26
r177 21 22 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.655 $Y=1.185
+ $X2=3.235 $Y2=1.185
r178 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.16 $Y=1.11
+ $X2=3.235 $Y2=1.185
r179 18 20 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.16 $Y=1.11
+ $X2=3.16 $Y2=0.715
r180 15 30 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.215 $Y=1.88
+ $X2=2.215 $Y2=1.79
r181 15 17 133.889 $w=1.8e-07 $l=5e-07 $layer=POLY_cond $X=2.215 $Y=1.88
+ $X2=2.215 $Y2=2.38
r182 13 29 20.4101 $w=1.5e-07 $l=8.57321e-08 $layer=POLY_cond $X=2.2 $Y=1.41
+ $X2=2.177 $Y2=1.335
r183 13 30 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.2 $Y=1.41 $X2=2.2
+ $Y2=1.79
r184 9 29 20.4101 $w=1.5e-07 $l=8.52936e-08 $layer=POLY_cond $X=2.155 $Y=1.26
+ $X2=2.177 $Y2=1.335
r185 9 11 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.155 $Y=1.26
+ $X2=2.155 $Y2=0.74
r186 8 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=1.335
+ $X2=1.72 $Y2=1.335
r187 7 29 5.30422 $w=1.5e-07 $l=9.7e-08 $layer=POLY_cond $X=2.08 $Y=1.335
+ $X2=2.177 $Y2=1.335
r188 7 8 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=2.08 $Y=1.335
+ $X2=1.885 $Y2=1.335
r189 2 51 300 $w=1.7e-07 $l=3.45977e-07 $layer=licon1_PDIFF $count=2 $X=1.18
+ $Y=2.12 $X2=1.315 $Y2=2.405
r190 1 33 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.49 $X2=1.3 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_2%A_27_136# 1 2 9 13 18 23 24 27 28 30 32 33
c79 27 0 8.07505e-20 $X=2.68 $Y=1.385
c80 23 0 1.8903e-19 $X=2.515 $Y=0.665
c81 13 0 2.97788e-19 $X=2.77 $Y=0.715
r82 32 33 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=0.272 $Y=2.265
+ $X2=0.272 $Y2=2.1
r83 30 33 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=0.185 $Y=1.25
+ $X2=0.185 $Y2=2.1
r84 28 36 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.385
+ $X2=2.68 $Y2=1.55
r85 28 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.385
+ $X2=2.68 $Y2=1.22
r86 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.385 $X2=2.68 $Y2=1.385
r87 25 27 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.68 $Y=0.75
+ $X2=2.68 $Y2=1.385
r88 23 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.515 $Y=0.665
+ $X2=2.68 $Y2=0.75
r89 23 24 135.048 $w=1.68e-07 $l=2.07e-06 $layer=LI1_cond $X=2.515 $Y=0.665
+ $X2=0.445 $Y2=0.665
r90 16 30 8.71323 $w=3.43e-07 $l=1.72e-07 $layer=LI1_cond $X=0.272 $Y=1.078
+ $X2=0.272 $Y2=1.25
r91 16 18 4.10871 $w=3.43e-07 $l=1.23e-07 $layer=LI1_cond $X=0.272 $Y=1.078
+ $X2=0.272 $Y2=0.955
r92 15 24 7.89393 $w=1.7e-07 $l=2.11268e-07 $layer=LI1_cond $X=0.272 $Y=0.75
+ $X2=0.445 $Y2=0.665
r93 15 18 6.84785 $w=3.43e-07 $l=2.05e-07 $layer=LI1_cond $X=0.272 $Y=0.75
+ $X2=0.272 $Y2=0.955
r94 13 35 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.77 $Y=0.715
+ $X2=2.77 $Y2=1.22
r95 9 36 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=2.75 $Y=2.46 $X2=2.75
+ $Y2=1.55
r96 2 32 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.265
r97 1 18 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.68 $X2=0.28 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_2%A_343_74# 1 2 9 13 15 16 22 25 26 30 32 33
+ 35 37 38 39
c110 38 0 8.07505e-20 $X=3.22 $Y=1.635
c111 32 0 6.57199e-20 $X=4.1 $Y=0.34
c112 25 0 1.29216e-19 $X=2.14 $Y=1.71
c113 16 0 1.68572e-19 $X=2.055 $Y=1.005
c114 13 0 1.87089e-19 $X=4.12 $Y=0.505
r115 38 44 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.635
+ $X2=3.22 $Y2=1.8
r116 37 40 4.98354 $w=3.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.2 $Y=1.635
+ $X2=3.2 $Y2=1.795
r117 37 39 8.53881 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.2 $Y=1.635
+ $X2=3.2 $Y2=1.47
r118 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.22
+ $Y=1.635 $X2=3.22 $Y2=1.635
r119 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.1
+ $Y=0.34 $X2=4.1 $Y2=0.34
r120 30 32 42.1794 $w=2.48e-07 $l=9.15e-07 $layer=LI1_cond $X=3.185 $Y=0.38
+ $X2=4.1 $Y2=0.38
r121 28 30 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.1 $Y=0.505
+ $X2=3.185 $Y2=0.38
r122 28 39 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=3.1 $Y=0.505
+ $X2=3.1 $Y2=1.47
r123 27 35 2.76166 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=2.225 $Y=1.795
+ $X2=2.025 $Y2=1.795
r124 26 40 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.015 $Y=1.795
+ $X2=3.2 $Y2=1.795
r125 26 27 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=3.015 $Y=1.795
+ $X2=2.225 $Y2=1.795
r126 25 35 3.70735 $w=2.5e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.14 $Y=1.71
+ $X2=2.025 $Y2=1.795
r127 24 25 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.14 $Y=1.09
+ $X2=2.14 $Y2=1.71
r128 20 35 3.70735 $w=2.5e-07 $l=1.00995e-07 $layer=LI1_cond $X=1.99 $Y=1.88
+ $X2=2.025 $Y2=1.795
r129 20 22 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.99 $Y=1.88
+ $X2=1.99 $Y2=2.12
r130 16 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.055 $Y=1.005
+ $X2=2.14 $Y2=1.09
r131 16 18 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.055 $Y=1.005
+ $X2=1.86 $Y2=1.005
r132 13 33 20.7597 $w=1.5e-07 $l=1.81659e-07 $layer=POLY_cond $X=4.12 $Y=0.505
+ $X2=4.155 $Y2=0.34
r133 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.12 $Y=0.505
+ $X2=4.12 $Y2=0.825
r134 9 44 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.17 $Y=2.46
+ $X2=3.17 $Y2=1.8
r135 2 22 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=1.845
+ $Y=1.96 $X2=1.99 $Y2=2.12
r136 1 18 182 $w=1.7e-07 $l=7.03776e-07 $layer=licon1_NDIFF $count=1 $X=1.715
+ $Y=0.37 $X2=1.86 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_2%A_887_270# 1 2 9 13 17 21 25 29 33 37 41 42
+ 44 45 49 52 55 56 60 61 65 67 68 70 80
c164 60 0 1.78677e-19 $X=6.87 $Y=1.63
c165 45 0 3.16539e-20 $X=4.775 $Y=1.805
c166 13 0 6.57199e-20 $X=4.58 $Y=0.825
r167 80 81 3.0125 $w=3.2e-07 $l=2e-08 $layer=POLY_cond $X=7.135 $Y=1.465
+ $X2=7.155 $Y2=1.465
r168 77 78 14.3094 $w=3.2e-07 $l=9.5e-08 $layer=POLY_cond $X=6.555 $Y=1.465
+ $X2=6.65 $Y2=1.465
r169 76 77 53.4719 $w=3.2e-07 $l=3.55e-07 $layer=POLY_cond $X=6.2 $Y=1.465
+ $X2=6.555 $Y2=1.465
r170 75 76 11.2969 $w=3.2e-07 $l=7.5e-08 $layer=POLY_cond $X=6.125 $Y=1.465
+ $X2=6.2 $Y2=1.465
r171 71 80 51.9656 $w=3.2e-07 $l=3.45e-07 $layer=POLY_cond $X=6.79 $Y=1.465
+ $X2=7.135 $Y2=1.465
r172 71 78 21.0875 $w=3.2e-07 $l=1.4e-07 $layer=POLY_cond $X=6.79 $Y=1.465
+ $X2=6.65 $Y2=1.465
r173 70 71 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.79
+ $Y=1.465 $X2=6.79 $Y2=1.465
r174 63 65 5.3159 $w=4.93e-07 $l=2.2e-07 $layer=LI1_cond $X=5.35 $Y=0.597
+ $X2=5.57 $Y2=0.597
r175 60 70 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.87 $Y=1.63
+ $X2=6.87 $Y2=1.465
r176 60 61 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.87 $Y=1.63
+ $X2=6.87 $Y2=2.24
r177 57 68 4.59089 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=5.655 $Y=2.325
+ $X2=5.452 $Y2=2.325
r178 56 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.785 $Y=2.325
+ $X2=6.87 $Y2=2.24
r179 56 57 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=6.785 $Y=2.325
+ $X2=5.655 $Y2=2.325
r180 55 67 3.27229 $w=2.87e-07 $l=1.54771e-07 $layer=LI1_cond $X=5.57 $Y=1.72
+ $X2=5.452 $Y2=1.805
r181 54 65 7.09362 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=5.57 $Y=0.845
+ $X2=5.57 $Y2=0.597
r182 54 55 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=5.57 $Y=0.845
+ $X2=5.57 $Y2=1.72
r183 50 68 2.39067 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.452 $Y=2.41
+ $X2=5.452 $Y2=2.325
r184 50 52 11.5244 $w=4.03e-07 $l=4.05e-07 $layer=LI1_cond $X=5.452 $Y=2.41
+ $X2=5.452 $Y2=2.815
r185 47 68 2.39067 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.452 $Y=2.24
+ $X2=5.452 $Y2=2.325
r186 47 49 7.25612 $w=4.03e-07 $l=2.55e-07 $layer=LI1_cond $X=5.452 $Y=2.24
+ $X2=5.452 $Y2=1.985
r187 46 67 3.27229 $w=2.87e-07 $l=8.5e-08 $layer=LI1_cond $X=5.452 $Y=1.89
+ $X2=5.452 $Y2=1.805
r188 46 49 2.70326 $w=4.03e-07 $l=9.5e-08 $layer=LI1_cond $X=5.452 $Y=1.89
+ $X2=5.452 $Y2=1.985
r189 44 67 3.2872 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=5.25 $Y=1.805
+ $X2=5.452 $Y2=1.805
r190 44 45 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=5.25 $Y=1.805
+ $X2=4.775 $Y2=1.805
r191 42 74 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=4.605 $Y=1.515
+ $X2=4.605 $Y2=1.68
r192 42 73 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=4.605 $Y=1.515
+ $X2=4.605 $Y2=1.35
r193 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.61
+ $Y=1.515 $X2=4.61 $Y2=1.515
r194 39 45 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.61 $Y=1.72
+ $X2=4.775 $Y2=1.805
r195 39 41 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=4.61 $Y=1.72
+ $X2=4.61 $Y2=1.515
r196 35 81 16.2157 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.155 $Y=1.63
+ $X2=7.155 $Y2=1.465
r197 35 37 322.629 $w=1.8e-07 $l=8.3e-07 $layer=POLY_cond $X=7.155 $Y=1.63
+ $X2=7.155 $Y2=2.46
r198 31 80 20.4921 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.135 $Y=1.3
+ $X2=7.135 $Y2=1.465
r199 31 33 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=7.135 $Y=1.3
+ $X2=7.135 $Y2=0.79
r200 27 78 16.2157 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.65 $Y=1.63
+ $X2=6.65 $Y2=1.465
r201 27 29 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=6.65 $Y=1.63
+ $X2=6.65 $Y2=2.4
r202 23 77 20.4921 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.555 $Y=1.3
+ $X2=6.555 $Y2=1.465
r203 23 25 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.555 $Y=1.3
+ $X2=6.555 $Y2=0.74
r204 19 76 16.2157 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.2 $Y=1.63
+ $X2=6.2 $Y2=1.465
r205 19 21 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=6.2 $Y=1.63 $X2=6.2
+ $Y2=2.4
r206 15 75 20.4921 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.125 $Y=1.3
+ $X2=6.125 $Y2=1.465
r207 15 17 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.125 $Y=1.3
+ $X2=6.125 $Y2=0.74
r208 13 73 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=4.58 $Y=0.825
+ $X2=4.58 $Y2=1.35
r209 9 74 190.468 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=4.525 $Y=2.17
+ $X2=4.525 $Y2=1.68
r210 2 52 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.28
+ $Y=1.84 $X2=5.415 $Y2=2.815
r211 2 49 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.28
+ $Y=1.84 $X2=5.415 $Y2=1.985
r212 1 63 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=5.21
+ $Y=0.37 $X2=5.35 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_2%A_647_79# 1 2 9 12 14 19 20 21 24 25 32 35
c89 25 0 1.15783e-19 $X=5.15 $Y=1.385
r90 30 32 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.64 $Y=2.135
+ $X2=3.77 $Y2=2.135
r91 27 29 7.64303 $w=4.23e-07 $l=2.65e-07 $layer=LI1_cond $X=3.64 $Y=0.955
+ $X2=3.905 $Y2=0.955
r92 25 36 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.15 $Y=1.385
+ $X2=5.15 $Y2=1.55
r93 25 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.15 $Y=1.385
+ $X2=5.15 $Y2=1.22
r94 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.15
+ $Y=1.385 $X2=5.15 $Y2=1.385
r95 22 24 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=5.15 $Y=1.185 $X2=5.15
+ $Y2=1.385
r96 21 29 9.26383 $w=4.23e-07 $l=2.26164e-07 $layer=LI1_cond $X=4.07 $Y=1.1
+ $X2=3.905 $Y2=0.955
r97 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.985 $Y=1.1
+ $X2=5.15 $Y2=1.185
r98 20 21 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=4.985 $Y=1.1
+ $X2=4.07 $Y2=1.1
r99 19 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=2.05
+ $X2=3.64 $Y2=2.135
r100 18 27 6.11956 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.64 $Y=1.185
+ $X2=3.64 $Y2=0.955
r101 18 19 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=3.64 $Y=1.185
+ $X2=3.64 $Y2=2.05
r102 14 30 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.555 $Y=2.135
+ $X2=3.64 $Y2=2.135
r103 14 16 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.555 $Y=2.135
+ $X2=3.395 $Y2=2.135
r104 12 36 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=5.19 $Y=2.4
+ $X2=5.19 $Y2=1.55
r105 9 35 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.135 $Y=0.74
+ $X2=5.135 $Y2=1.22
r106 2 32 600 $w=1.7e-07 $l=5.91058e-07 $layer=licon1_PDIFF $count=1 $X=3.26
+ $Y=1.96 $X2=3.77 $Y2=2.135
r107 2 16 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.26
+ $Y=1.96 $X2=3.395 $Y2=2.135
r108 1 29 91 $w=1.7e-07 $l=8.83487e-07 $layer=licon1_NDIFF $count=2 $X=3.235
+ $Y=0.395 $X2=3.905 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_2%A_1442_94# 1 2 9 13 15 17 21 23 30 33 36 42
+ 45 46
c65 36 0 1.28661e-19 $X=7.38 $Y=2.105
c66 23 0 1.78677e-19 $X=8.075 $Y=1.485
r67 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.99
+ $Y=1.485 $X2=7.99 $Y2=1.485
r68 40 46 1.17559 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.545 $Y=1.485
+ $X2=7.38 $Y2=1.485
r69 40 42 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=7.545 $Y=1.485
+ $X2=7.99 $Y2=1.485
r70 36 38 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=7.38 $Y=2.105
+ $X2=7.38 $Y2=2.815
r71 34 46 5.36902 $w=3.15e-07 $l=1.65e-07 $layer=LI1_cond $X=7.38 $Y=1.65
+ $X2=7.38 $Y2=1.485
r72 34 36 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=7.38 $Y=1.65
+ $X2=7.38 $Y2=2.105
r73 33 46 5.36902 $w=3.15e-07 $l=1.72337e-07 $layer=LI1_cond $X=7.365 $Y=1.32
+ $X2=7.38 $Y2=1.485
r74 33 45 7.29881 $w=2.98e-07 $l=1.9e-07 $layer=LI1_cond $X=7.365 $Y=1.32
+ $X2=7.365 $Y2=1.13
r75 28 45 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.35 $Y=0.965
+ $X2=7.35 $Y2=1.13
r76 28 30 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=7.35 $Y=0.965
+ $X2=7.35 $Y2=0.615
r77 24 25 4.44923 $w=3.25e-07 $l=3e-08 $layer=POLY_cond $X=8.165 $Y=1.485
+ $X2=8.195 $Y2=1.485
r78 23 43 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=8.075 $Y=1.485
+ $X2=7.99 $Y2=1.485
r79 23 24 13.1455 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.075 $Y=1.485
+ $X2=8.165 $Y2=1.485
r80 19 27 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.625 $Y=1.32
+ $X2=8.625 $Y2=1.485
r81 19 21 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.625 $Y=1.32
+ $X2=8.625 $Y2=0.74
r82 15 27 1.48308 $w=3.25e-07 $l=1e-08 $layer=POLY_cond $X=8.615 $Y=1.485
+ $X2=8.625 $Y2=1.485
r83 15 25 62.2892 $w=3.25e-07 $l=4.2e-07 $layer=POLY_cond $X=8.615 $Y=1.485
+ $X2=8.195 $Y2=1.485
r84 15 17 293.476 $w=1.8e-07 $l=7.55e-07 $layer=POLY_cond $X=8.615 $Y=1.645
+ $X2=8.615 $Y2=2.4
r85 11 25 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.195 $Y=1.32
+ $X2=8.195 $Y2=1.485
r86 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.195 $Y=1.32
+ $X2=8.195 $Y2=0.74
r87 7 24 16.5763 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.165 $Y=1.65
+ $X2=8.165 $Y2=1.485
r88 7 9 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=8.165 $Y=1.65
+ $X2=8.165 $Y2=2.4
r89 2 38 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.245
+ $Y=1.96 $X2=7.38 $Y2=2.815
r90 2 36 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.245
+ $Y=1.96 $X2=7.38 $Y2=2.105
r91 1 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.21
+ $Y=0.47 $X2=7.35 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_2%VPWR 1 2 3 4 5 6 7 26 30 34 40 44 48 52 54
+ 59 60 62 63 64 66 78 86 90 96 99 102 105 109
r99 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r100 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r101 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r102 99 100 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r103 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r104 94 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r105 94 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r106 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r107 91 105 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=7.9 $Y2=3.33
r108 91 93 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=8.4 $Y2=3.33
r109 90 108 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=8.755 $Y=3.33
+ $X2=8.937 $Y2=3.33
r110 90 93 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.755 $Y=3.33
+ $X2=8.4 $Y2=3.33
r111 89 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r112 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r113 86 105 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.775 $Y=3.33
+ $X2=7.9 $Y2=3.33
r114 86 88 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.775 $Y=3.33
+ $X2=7.44 $Y2=3.33
r115 85 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r116 85 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r117 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r118 82 102 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.14 $Y=3.33
+ $X2=6.015 $Y2=3.33
r119 82 84 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.14 $Y=3.33
+ $X2=6.48 $Y2=3.33
r120 81 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r121 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r122 78 102 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.89 $Y=3.33
+ $X2=6.015 $Y2=3.33
r123 78 80 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.89 $Y=3.33
+ $X2=5.52 $Y2=3.33
r124 74 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=3.33
+ $X2=2.525 $Y2=3.33
r125 74 76 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=2.69 $Y=3.33 $X2=4.56
+ $Y2=3.33
r126 73 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r127 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r128 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r129 70 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r130 69 72 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r131 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r132 67 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r133 67 69 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=1.2 $Y2=3.33
r134 66 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=3.33
+ $X2=2.525 $Y2=3.33
r135 66 72 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.36 $Y=3.33 $X2=2.16
+ $Y2=3.33
r136 64 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r137 64 100 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=2.64 $Y2=3.33
r138 64 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r139 62 84 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.71 $Y=3.33
+ $X2=6.48 $Y2=3.33
r140 62 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.71 $Y=3.33
+ $X2=6.875 $Y2=3.33
r141 61 88 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=7.04 $Y=3.33 $X2=7.44
+ $Y2=3.33
r142 61 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.04 $Y=3.33
+ $X2=6.875 $Y2=3.33
r143 59 76 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=4.67 $Y=3.33
+ $X2=4.56 $Y2=3.33
r144 59 60 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=4.67 $Y=3.33
+ $X2=4.875 $Y2=3.33
r145 58 80 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.08 $Y=3.33
+ $X2=5.52 $Y2=3.33
r146 58 60 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=5.08 $Y=3.33
+ $X2=4.875 $Y2=3.33
r147 54 57 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=8.88 $Y=1.985
+ $X2=8.88 $Y2=2.815
r148 52 108 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.88 $Y=3.245
+ $X2=8.937 $Y2=3.33
r149 52 57 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.88 $Y=3.245
+ $X2=8.88 $Y2=2.815
r150 48 51 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=7.9 $Y=1.985
+ $X2=7.9 $Y2=2.815
r151 46 105 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=3.245
+ $X2=7.9 $Y2=3.33
r152 46 51 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.9 $Y=3.245 $X2=7.9
+ $Y2=2.815
r153 42 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.875 $Y=3.245
+ $X2=6.875 $Y2=3.33
r154 42 44 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=6.875 $Y=3.245
+ $X2=6.875 $Y2=2.78
r155 38 102 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.015 $Y=3.245
+ $X2=6.015 $Y2=3.33
r156 38 40 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=6.015 $Y=3.245
+ $X2=6.015 $Y2=2.78
r157 34 37 9.55684 $w=4.08e-07 $l=3.4e-07 $layer=LI1_cond $X=4.875 $Y=2.155
+ $X2=4.875 $Y2=2.495
r158 32 60 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.875 $Y=3.245
+ $X2=4.875 $Y2=3.33
r159 32 37 21.0813 $w=4.08e-07 $l=7.5e-07 $layer=LI1_cond $X=4.875 $Y=3.245
+ $X2=4.875 $Y2=2.495
r160 28 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=3.245
+ $X2=2.525 $Y2=3.33
r161 28 30 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.525 $Y=3.245
+ $X2=2.525 $Y2=2.815
r162 24 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r163 24 26 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.405
r164 7 57 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.705
+ $Y=1.84 $X2=8.84 $Y2=2.815
r165 7 54 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.705
+ $Y=1.84 $X2=8.84 $Y2=1.985
r166 6 51 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=7.795
+ $Y=1.84 $X2=7.94 $Y2=2.815
r167 6 48 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=7.795
+ $Y=1.84 $X2=7.94 $Y2=1.985
r168 5 44 600 $w=1.7e-07 $l=1.00524e-06 $layer=licon1_PDIFF $count=1 $X=6.74
+ $Y=1.84 $X2=6.875 $Y2=2.78
r169 4 40 600 $w=1.7e-07 $l=1.0099e-06 $layer=licon1_PDIFF $count=1 $X=5.83
+ $Y=1.84 $X2=5.975 $Y2=2.78
r170 3 37 300 $w=1.7e-07 $l=6.52169e-07 $layer=licon1_PDIFF $count=2 $X=4.615
+ $Y=1.96 $X2=4.875 $Y2=2.495
r171 3 34 600 $w=1.7e-07 $l=3.43948e-07 $layer=licon1_PDIFF $count=1 $X=4.615
+ $Y=1.96 $X2=4.875 $Y2=2.155
r172 2 30 600 $w=1.7e-07 $l=9.5871e-07 $layer=licon1_PDIFF $count=1 $X=2.305
+ $Y=1.96 $X2=2.525 $Y2=2.815
r173 1 26 300 $w=1.7e-07 $l=3.45977e-07 $layer=licon1_PDIFF $count=2 $X=0.68
+ $Y=2.12 $X2=0.815 $Y2=2.405
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_2%Q 1 2 7 9 13 20 23 24
r44 23 24 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6 $Y=1.295 $X2=6
+ $Y2=1.665
r45 22 24 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=6 $Y=1.8 $X2=6
+ $Y2=1.665
r46 19 20 1.44055 $w=2.78e-07 $l=3.5e-08 $layer=LI1_cond $X=6.34 $Y=0.99
+ $X2=6.375 $Y2=0.99
r47 16 23 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6 $Y=1.13 $X2=6
+ $Y2=1.295
r48 15 19 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=6 $Y=0.99 $X2=6.34
+ $Y2=0.99
r49 15 16 1.89134 $w=2.3e-07 $l=1.4e-07 $layer=LI1_cond $X=6 $Y=0.99 $X2=6
+ $Y2=1.13
r50 11 20 1.16438 $w=2.6e-07 $l=1.4e-07 $layer=LI1_cond $X=6.375 $Y=0.85
+ $X2=6.375 $Y2=0.99
r51 11 13 14.6272 $w=2.58e-07 $l=3.3e-07 $layer=LI1_cond $X=6.375 $Y=0.85
+ $X2=6.375 $Y2=0.52
r52 7 22 6.87339 $w=2.7e-07 $l=1.83712e-07 $layer=LI1_cond $X=6.115 $Y=1.935
+ $X2=6 $Y2=1.8
r53 7 9 13.2318 $w=2.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.115 $Y=1.935
+ $X2=6.425 $Y2=1.935
r54 2 9 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.29
+ $Y=1.84 $X2=6.425 $Y2=1.985
r55 1 19 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=6.2
+ $Y=0.37 $X2=6.34 $Y2=0.95
r56 1 13 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=6.2
+ $Y=0.37 $X2=6.34 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_2%Q_N 1 2 9 13 14 15 16 24 33
r24 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.39 $Y=2.405
+ $X2=8.39 $Y2=2.775
r25 14 24 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=8.39 $Y=1.967
+ $X2=8.39 $Y2=1.985
r26 14 33 7.83357 $w=3.28e-07 $l=1.47e-07 $layer=LI1_cond $X=8.39 $Y=1.967
+ $X2=8.39 $Y2=1.82
r27 14 15 12.3276 $w=3.28e-07 $l=3.53e-07 $layer=LI1_cond $X=8.39 $Y=2.052
+ $X2=8.39 $Y2=2.405
r28 14 24 2.33981 $w=3.28e-07 $l=6.7e-08 $layer=LI1_cond $X=8.39 $Y=2.052
+ $X2=8.39 $Y2=1.985
r29 13 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.41 $Y=1.13 $X2=8.41
+ $Y2=1.82
r30 7 13 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=8.37 $Y=1.005
+ $X2=8.37 $Y2=1.13
r31 7 9 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=8.37 $Y=1.005 $X2=8.37
+ $Y2=0.515
r32 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.255
+ $Y=1.84 $X2=8.39 $Y2=2.815
r33 2 24 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.255
+ $Y=1.84 $X2=8.39 $Y2=1.985
r34 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.27
+ $Y=0.37 $X2=8.41 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_2%VGND 1 2 3 4 5 6 7 24 28 32 38 40 42 45 52
+ 53 55 56 58 59 60 62 86 90 97 103 107
c104 24 0 1.15783e-19 $X=4.82 $Y=0.76
r105 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r106 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r107 97 100 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.79 $Y=0
+ $X2=0.79 $Y2=0.325
r108 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r109 94 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r110 94 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r111 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r112 91 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.075 $Y=0
+ $X2=7.91 $Y2=0
r113 91 93 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.075 $Y=0 $X2=8.4
+ $Y2=0
r114 90 106 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=8.675 $Y=0
+ $X2=8.897 $Y2=0
r115 90 93 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.675 $Y=0 $X2=8.4
+ $Y2=0
r116 89 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r117 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r118 86 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.91 $Y2=0
r119 86 88 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.44 $Y2=0
r120 85 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r121 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r122 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r123 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r124 75 78 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r125 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r126 73 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r127 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r128 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r129 70 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r130 69 72 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r131 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r132 67 97 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r133 67 69 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r134 65 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r135 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r136 62 97 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r137 62 64 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r138 60 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r139 60 76 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=2.64 $Y2=0
r140 60 78 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r141 58 84 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.675 $Y=0
+ $X2=6.48 $Y2=0
r142 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.675 $Y=0 $X2=6.84
+ $Y2=0
r143 57 88 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.005 $Y=0
+ $X2=7.44 $Y2=0
r144 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.005 $Y=0 $X2=6.84
+ $Y2=0
r145 55 81 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.825 $Y=0
+ $X2=5.52 $Y2=0
r146 55 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.825 $Y=0 $X2=5.95
+ $Y2=0
r147 54 84 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=6.075 $Y=0
+ $X2=6.48 $Y2=0
r148 54 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.075 $Y=0 $X2=5.95
+ $Y2=0
r149 52 78 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=4.63 $Y=0 $X2=4.56
+ $Y2=0
r150 52 53 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=4.63 $Y=0 $X2=4.822
+ $Y2=0
r151 51 81 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=5.015 $Y=0
+ $X2=5.52 $Y2=0
r152 51 53 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=5.015 $Y=0
+ $X2=4.822 $Y2=0
r153 45 72 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.285 $Y=0
+ $X2=2.16 $Y2=0
r154 45 49 10.5505 $w=3.53e-07 $l=3.25e-07 $layer=LI1_cond $X=2.462 $Y=0
+ $X2=2.462 $Y2=0.325
r155 45 75 5.0588 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=2.462 $Y=0 $X2=2.64
+ $Y2=0
r156 40 106 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.84 $Y=0.085
+ $X2=8.897 $Y2=0
r157 40 42 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.84 $Y=0.085
+ $X2=8.84 $Y2=0.515
r158 36 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0
r159 36 38 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0.515
r160 32 34 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=6.84 $Y=0.515
+ $X2=6.84 $Y2=0.965
r161 30 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=0.085
+ $X2=6.84 $Y2=0
r162 30 32 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.84 $Y=0.085
+ $X2=6.84 $Y2=0.515
r163 26 56 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.95 $Y=0.085
+ $X2=5.95 $Y2=0
r164 26 28 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.95 $Y=0.085
+ $X2=5.95 $Y2=0.515
r165 22 53 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.822 $Y=0.085
+ $X2=4.822 $Y2=0
r166 22 24 20.2052 $w=3.83e-07 $l=6.75e-07 $layer=LI1_cond $X=4.822 $Y=0.085
+ $X2=4.822 $Y2=0.76
r167 7 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.7
+ $Y=0.37 $X2=8.84 $Y2=0.515
r168 6 38 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=7.765
+ $Y=0.37 $X2=7.91 $Y2=0.515
r169 5 34 182 $w=1.7e-07 $l=6.9208e-07 $layer=licon1_NDIFF $count=1 $X=6.63
+ $Y=0.37 $X2=6.84 $Y2=0.965
r170 5 32 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=6.63
+ $Y=0.37 $X2=6.84 $Y2=0.515
r171 4 28 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=5.765
+ $Y=0.37 $X2=5.91 $Y2=0.515
r172 3 24 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=4.655
+ $Y=0.615 $X2=4.82 $Y2=0.76
r173 2 49 182 $w=1.7e-07 $l=2.51496e-07 $layer=licon1_NDIFF $count=1 $X=2.23
+ $Y=0.37 $X2=2.46 $Y2=0.325
r174 1 100 182 $w=1.7e-07 $l=4.51802e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.68 $X2=0.79 $Y2=0.325
.ends


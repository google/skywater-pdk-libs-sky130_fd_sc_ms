* File: sky130_fd_sc_ms__sdfsbp_1.spice
* Created: Wed Sep  2 12:30:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdfsbp_1.pex.spice"
.subckt sky130_fd_sc_ms__sdfsbp_1  VNB VPB SCE D SCD CLK SET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1036 N_VGND_M1036_d N_SCE_M1036_g N_A_27_74#_M1036_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0882 AS=0.1197 PD=0.84 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1039 A_228_74# N_A_27_74#_M1039_g N_VGND_M1036_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0882 PD=0.66 PS=0.84 NRD=18.564 NRS=19.992 M=1 R=2.8 SA=75000.8
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1040 N_A_293_464#_M1040_d N_D_M1040_g A_228_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1015 A_392_74# N_SCE_M1015_g N_A_293_464#_M1040_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_SCD_M1016_g A_392_74# VNB NLOWVT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_CLK_M1023_g N_A_594_74#_M1023_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1019 N_A_781_74#_M1019_d N_A_594_74#_M1019_g N_VGND_M1023_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1037 N_A_995_74#_M1037_d N_A_594_74#_M1037_g N_A_293_464#_M1037_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0945 AS=0.18665 PD=0.87 PS=1.8 NRD=48.564 NRS=24.276 M=1
+ R=2.8 SA=75000.3 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1007 A_1115_74# N_A_781_74#_M1007_g N_A_995_74#_M1037_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0945 PD=0.66 PS=0.87 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_1163_48#_M1005_g A_1115_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.17255 AS=0.0504 PD=1.68 PS=0.66 NRD=25.704 NRS=18.564 M=1 R=2.8
+ SA=75001.3 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1001 A_1411_74# N_A_995_74#_M1001_g N_A_1163_48#_M1001_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.2 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_SET_B_M1014_g A_1411_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.20267 AS=0.0504 PD=1.16094 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75003.9 A=0.063 P=1.14 MULT=1
MM1024 A_1684_74# N_A_995_74#_M1024_g N_VGND_M1014_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.30883 PD=0.88 PS=1.76906 NRD=12.18 NRS=0 M=1 R=4.26667
+ SA=75001.3 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1025 N_A_1762_74#_M1025_d N_A_781_74#_M1025_g A_1684_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.144362 AS=0.0768 PD=1.28 PS=0.88 NRD=13.116 NRS=12.18 M=1
+ R=4.26667 SA=75001.7 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1003 A_1876_74# N_A_594_74#_M1003_g N_A_1762_74#_M1025_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0947377 PD=0.66 PS=0.84 NRD=18.564 NRS=20.712 M=1 R=2.8
+ SA=75002.5 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1004 A_1954_74# N_A_1924_48#_M1004_g A_1876_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0504 PD=0.81 PS=0.66 NRD=39.996 NRS=18.564 M=1 R=2.8 SA=75002.9
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_SET_B_M1012_g A_1954_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1323 AS=0.0819 PD=1.05 PS=0.81 NRD=0 NRS=39.996 M=1 R=2.8 SA=75003.5
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1006 N_A_1924_48#_M1006_d N_A_1762_74#_M1006_g N_VGND_M1012_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1197 AS=0.1323 PD=1.41 PS=1.05 NRD=0 NRS=0 M=1 R=2.8
+ SA=75004.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_Q_N_M1009_d N_A_1762_74#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.2627 PD=2.05 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1018_d N_A_1762_74#_M1018_g N_A_2556_112#_M1018_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.172973 AS=0.15675 PD=1.15543 PS=1.67 NRD=58.356 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75001 A=0.0825 P=1.4 MULT=1
MM1027 N_Q_M1027_d N_A_2556_112#_M1027_g N_VGND_M1018_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.232727 PD=2.05 PS=1.55457 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_VPWR_M1010_d N_SCE_M1010_g N_A_27_74#_M1010_s VPB PSHORT L=0.18 W=0.64
+ AD=0.0864 AS=0.1792 PD=0.91 PS=1.84 NRD=0 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90002.1 A=0.1152 P=1.64 MULT=1
MM1011 A_209_464# N_SCE_M1011_g N_VPWR_M1010_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.0864 PD=0.88 PS=0.91 NRD=19.9955 NRS=0 M=1 R=3.55556 SA=90000.6
+ SB=90001.7 A=0.1152 P=1.64 MULT=1
MM1017 N_A_293_464#_M1017_d N_D_M1017_g A_209_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.144 AS=0.0768 PD=1.09 PS=0.88 NRD=26.1616 NRS=19.9955 M=1 R=3.55556
+ SA=90001.1 SB=90001.3 A=0.1152 P=1.64 MULT=1
MM1002 A_419_464# N_A_27_74#_M1002_g N_A_293_464#_M1017_d VPB PSHORT L=0.18
+ W=0.64 AD=0.0768 AS=0.144 PD=0.88 PS=1.09 NRD=19.9955 NRS=26.1616 M=1
+ R=3.55556 SA=90001.7 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1013 N_VPWR_M1013_d N_SCD_M1013_g A_419_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.1984 AS=0.0768 PD=1.9 PS=0.88 NRD=0 NRS=19.9955 M=1 R=3.55556 SA=90002.1
+ SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1026 N_VPWR_M1026_d N_CLK_M1026_g N_A_594_74#_M1026_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.308 PD=1.39 PS=2.79 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1030 N_A_781_74#_M1030_d N_A_594_74#_M1030_g N_VPWR_M1026_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3024 AS=0.1512 PD=2.78 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1022 N_A_995_74#_M1022_d N_A_781_74#_M1022_g N_A_293_464#_M1022_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0995625 AS=0.1134 PD=0.92 PS=1.38 NRD=32.8202 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90002.6 A=0.0756 P=1.2 MULT=1
MM1020 A_1136_478# N_A_594_74#_M1020_g N_A_995_74#_M1022_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0774 AS=0.0995625 PD=0.835 PS=0.92 NRD=60.6366 NRS=35.1645 M=1
+ R=2.33333 SA=90000.7 SB=90002.1 A=0.0756 P=1.2 MULT=1
MM1021 N_VPWR_M1021_d N_A_1163_48#_M1021_g A_1136_478# VPB PSHORT L=0.18 W=0.42
+ AD=0.10605 AS=0.0774 PD=0.925 PS=0.835 NRD=0 NRS=60.6366 M=1 R=2.33333
+ SA=90001.1 SB=90002 A=0.0756 P=1.2 MULT=1
MM1038 N_A_1163_48#_M1038_d N_A_995_74#_M1038_g N_VPWR_M1021_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0861 AS=0.10605 PD=0.83 PS=0.925 NRD=0 NRS=105.533 M=1 R=2.33333
+ SA=90001.8 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1035 N_VPWR_M1035_d N_SET_B_M1035_g N_A_1163_48#_M1038_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0876085 AS=0.0861 PD=0.804507 PS=0.83 NRD=39.8531 NRS=63.3158 M=1
+ R=2.33333 SA=90002.4 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1041 N_A_1603_347#_M1041_d N_A_995_74#_M1041_g N_VPWR_M1035_d VPB PSHORT
+ L=0.18 W=1 AD=0.275 AS=0.208592 PD=2.55 PS=1.91549 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90001.3 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1033 N_A_1762_74#_M1033_d N_A_781_74#_M1033_g N_A_1712_374#_M1033_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0876085 AS=0.2463 PD=0.804507 PS=3 NRD=37.5088 NRS=249.264
+ M=1 R=2.33333 SA=90000.2 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1008 N_A_1603_347#_M1008_d N_A_594_74#_M1008_g N_A_1762_74#_M1033_d VPB PSHORT
+ L=0.18 W=1 AD=0.275 AS=0.208592 PD=2.55 PS=1.91549 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.4 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1028 N_VPWR_M1028_d N_A_1924_48#_M1028_g N_A_1712_374#_M1028_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0567 AS=0.1155 PD=0.69 PS=1.39 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1032 N_A_1762_74#_M1032_d N_SET_B_M1032_g N_VPWR_M1028_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1155 AS=0.0567 PD=1.39 PS=0.69 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1029 N_VPWR_M1029_d N_A_1762_74#_M1029_g N_A_1924_48#_M1029_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0849545 AS=0.1155 PD=0.788182 PS=1.39 NRD=0 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1000 N_Q_N_M1000_d N_A_1762_74#_M1000_g N_VPWR_M1029_d VPB PSHORT L=0.18
+ W=1.12 AD=0.308 AS=0.226545 PD=2.79 PS=2.10182 NRD=0 NRS=8.7862 M=1 R=6.22222
+ SA=90000.4 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1034 N_VPWR_M1034_d N_A_1762_74#_M1034_g N_A_2556_112#_M1034_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.147 AS=0.231 PD=1.23857 PS=2.23 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1031 N_Q_M1031_d N_A_2556_112#_M1031_g N_VPWR_M1034_d VPB PSHORT L=0.18 W=1.12
+ AD=0.308 AS=0.196 PD=2.79 PS=1.65143 NRD=0 NRS=8.7862 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX42_noxref VNB VPB NWDIODE A=27.6026 P=33.49
*
.include "sky130_fd_sc_ms__sdfsbp_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__a21bo_4.spice
* Created: Fri Aug 28 16:58:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a21bo_4.pex.spice"
.subckt sky130_fd_sc_ms__a21bo_4  VNB VPB B1_N A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_B1_N_M1009_g N_A_29_392#_M1009_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.149542 AS=0.1696 PD=1.10841 PS=1.81 NRD=15.468 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75005 A=0.096 P=1.58 MULT=1
MM1003 N_X_M1003_d N_A_184_338#_M1003_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.172908 PD=1.02 PS=1.28159 NRD=0 NRS=12.972 M=1 R=4.93333
+ SA=75000.7 SB=75004.1 A=0.111 P=1.78 MULT=1
MM1008 N_X_M1003_d N_A_184_338#_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75003.6 A=0.111 P=1.78 MULT=1
MM1011 N_X_M1011_d N_A_184_338#_M1011_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1013 N_X_M1011_d N_A_184_338#_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.132302 PD=1.02 PS=1.17435 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1013_s N_A_29_392#_M1017_g N_A_184_338#_M1017_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.114423 AS=0.0896 PD=1.01565 PS=0.92 NRD=11.244 NRS=0 M=1 R=4.26667
+ SA=75002.5 SB=75002.8 A=0.096 P=1.58 MULT=1
MM1020 N_VGND_M1020_d N_A_29_392#_M1020_g N_A_184_338#_M1017_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.2016 AS=0.0896 PD=1.27 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.9 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1012 N_VGND_M1020_d N_A2_M1012_g N_A_864_123#_M1012_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.2016 AS=0.1088 PD=1.27 PS=0.98 NRD=65.616 NRS=11.244 M=1 R=4.26667
+ SA=75003.7 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1010 N_A_864_123#_M1012_s N_A1_M1010_g N_A_184_338#_M1010_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1088 AS=0.0896 PD=0.98 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75004.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1014 N_A_864_123#_M1014_d N_A1_M1014_g N_A_184_338#_M1010_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75004.6 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1019 N_VGND_M1019_d N_A2_M1019_g N_A_864_123#_M1014_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75005.1
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1016 N_VPWR_M1016_d N_B1_N_M1016_g N_A_29_392#_M1016_s VPB PSHORT L=0.18 W=1
+ AD=0.172736 AS=0.26 PD=1.37264 PS=2.52 NRD=11.8003 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90002 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1016_d N_A_184_338#_M1001_g N_X_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.193464 AS=0.1512 PD=1.53736 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1004 N_VPWR_M1004_d N_A_184_338#_M1004_g N_X_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1006 N_VPWR_M1004_d N_A_184_338#_M1006_g N_X_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1021 N_VPWR_M1021_d N_A_184_338#_M1021_g N_X_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2912 AS=0.1512 PD=2.76 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1000 N_A_184_338#_M1000_d N_A_29_392#_M1000_g N_A_596_392#_M1000_s VPB PSHORT
+ L=0.18 W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90002.4 A=0.18 P=2.36 MULT=1
MM1002 N_A_184_338#_M1000_d N_A_29_392#_M1002_g N_A_596_392#_M1002_s VPB PSHORT
+ L=0.18 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.6 SB=90002 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_A2_M1005_g N_A_596_392#_M1002_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.1
+ SB=90001.5 A=0.18 P=2.36 MULT=1
MM1007 N_A_596_392#_M1007_d N_A1_M1007_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.5
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1015 N_A_596_392#_M1007_d N_A1_M1015_g N_VPWR_M1015_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90002
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1018 N_VPWR_M1015_s N_A2_M1018_g N_A_596_392#_M1018_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=5.55556 SA=90002.4
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX22_noxref VNB VPB NWDIODE A=12.3132 P=16.96
*
.include "sky130_fd_sc_ms__a21bo_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__sdfrtp_2.spice
* Created: Wed Sep  2 12:30:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdfrtp_2.pex.spice"
.subckt sky130_fd_sc_ms__sdfrtp_2  VNB VPB SCE D SCD CLK RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1036 N_VGND_M1036_d N_SCE_M1036_g N_A_27_74#_M1036_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1014 noxref_25 N_A_27_74#_M1014_g N_noxref_24_M1014_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1015 N_A_390_81#_M1015_d N_D_M1015_g noxref_25 VNB NLOWVT L=0.15 W=0.42
+ AD=0.13335 AS=0.0504 PD=1.055 PS=0.66 NRD=99.996 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1008 noxref_26 N_SCE_M1008_g N_A_390_81#_M1015_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.13335 PD=0.66 PS=1.055 NRD=18.564 NRS=1.428 M=1 R=2.8
+ SA=75001.4 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1035 N_noxref_24_M1035_d N_SCD_M1035_g noxref_26 VNB NLOWVT L=0.15 W=0.42
+ AD=0.06615 AS=0.0504 PD=0.735 PS=0.66 NRD=9.996 NRS=18.564 M=1 R=2.8
+ SA=75001.8 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_RESET_B_M1004_g N_noxref_24_M1035_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.1365 AS=0.06615 PD=1.49 PS=0.735 NRD=17.136 NRS=0 M=1 R=2.8
+ SA=75002.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_CLK_M1016_g N_A_837_119#_M1016_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.179025 AS=0.20225 PD=1.335 PS=2.04 NRD=12.156 NRS=2.424 M=1
+ R=4.93333 SA=75000.2 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1017 N_A_1037_119#_M1017_d N_A_837_119#_M1017_g N_VGND_M1016_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1998 AS=0.179025 PD=2.02 PS=1.335 NRD=0 NRS=12.156 M=1
+ R=4.93333 SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1031 N_A_1235_119#_M1031_d N_A_837_119#_M1031_g N_A_390_81#_M1031_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.09345 AS=0.126 PD=0.865 PS=1.44 NRD=47.136 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.3 A=0.063 P=1.14 MULT=1
MM1032 A_1354_119# N_A_1037_119#_M1032_g N_A_1235_119#_M1031_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.09345 PD=0.66 PS=0.865 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.8 SB=75003.7 A=0.063 P=1.14 MULT=1
MM1022 A_1432_119# N_A_1383_349#_M1022_g A_1354_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.2
+ SB=75003.3 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_RESET_B_M1007_g A_1432_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.266392 AS=0.0504 PD=1.33603 PS=0.66 NRD=165.504 NRS=18.564 M=1 R=2.8
+ SA=75001.6 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1040 N_A_1383_349#_M1040_d N_A_1235_119#_M1040_g N_VGND_M1007_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.13135 AS=0.469358 PD=1.095 PS=2.35397 NRD=0 NRS=93.924 M=1
+ R=4.93333 SA=75001.8 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1028 N_A_1824_74#_M1028_d N_A_1037_119#_M1028_g N_A_1383_349#_M1040_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.351117 AS=0.13135 PD=2.3731 PS=1.095 NRD=54.324
+ NRS=12.156 M=1 R=4.93333 SA=75002.3 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1009 A_2078_74# N_A_837_119#_M1009_g N_A_1824_74#_M1028_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.199283 PD=0.66 PS=1.3469 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75003.4 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_2082_446#_M1010_g A_2078_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75003.8
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1026 A_2242_74# N_RESET_B_M1026_g N_VGND_M1010_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75004.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1018 N_A_2082_446#_M1018_d N_A_1824_74#_M1018_g A_2242_74# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75004.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1029 N_A_2495_392#_M1029_d N_A_1824_74#_M1029_g N_VGND_M1029_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.1824 PD=1.85 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1003 N_Q_M1003_d N_A_2495_392#_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1030 N_Q_M1003_d N_A_2495_392#_M1030_g N_VGND_M1030_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_VPWR_M1011_d N_SCE_M1011_g N_A_27_74#_M1011_s VPB PSHORT L=0.18 W=0.64
+ AD=0.320037 AS=0.1792 PD=1.675 PS=1.84 NRD=136.994 NRS=0 M=1 R=3.55556
+ SA=90000.2 SB=90002.9 A=0.1152 P=1.64 MULT=1
MM1012 A_343_483# N_SCE_M1012_g N_VPWR_M1011_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0736 AS=0.320037 PD=0.87 PS=1.675 NRD=18.4589 NRS=136.994 M=1 R=3.55556
+ SA=90001.2 SB=90002.2 A=0.1152 P=1.64 MULT=1
MM1000 N_A_390_81#_M1000_d N_D_M1000_g A_343_483# VPB PSHORT L=0.18 W=0.64
+ AD=0.0896 AS=0.0736 PD=0.92 PS=0.87 NRD=1.5366 NRS=18.4589 M=1 R=3.55556
+ SA=90001.6 SB=90001.8 A=0.1152 P=1.64 MULT=1
MM1038 A_517_483# N_A_27_74#_M1038_g N_A_390_81#_M1000_d VPB PSHORT L=0.18
+ W=0.64 AD=0.1152 AS=0.0896 PD=1 PS=0.92 NRD=38.4741 NRS=0 M=1 R=3.55556
+ SA=90002.1 SB=90001.3 A=0.1152 P=1.64 MULT=1
MM1039 N_VPWR_M1039_d N_SCD_M1039_g A_517_483# VPB PSHORT L=0.18 W=0.64
+ AD=0.0928 AS=0.1152 PD=0.93 PS=1 NRD=0 NRS=38.4741 M=1 R=3.55556 SA=90002.6
+ SB=90000.8 A=0.1152 P=1.64 MULT=1
MM1023 N_A_390_81#_M1023_d N_RESET_B_M1023_g N_VPWR_M1039_d VPB PSHORT L=0.18
+ W=0.64 AD=0.2432 AS=0.0928 PD=2.04 PS=0.93 NRD=29.2348 NRS=4.6098 M=1
+ R=3.55556 SA=90003.1 SB=90000.3 A=0.1152 P=1.64 MULT=1
MM1027 N_VPWR_M1027_d N_CLK_M1027_g N_A_837_119#_M1027_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1034 N_A_1037_119#_M1034_d N_A_837_119#_M1034_g N_VPWR_M1027_d VPB PSHORT
+ L=0.18 W=1.12 AD=0.2912 AS=0.1512 PD=2.76 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1002 N_A_1235_119#_M1002_d N_A_1037_119#_M1002_g N_A_390_81#_M1002_s VPB
+ PSHORT L=0.18 W=0.42 AD=0.0609 AS=0.1176 PD=0.71 PS=1.4 NRD=0 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90001.7 A=0.0756 P=1.2 MULT=1
MM1025 A_1339_457# N_A_837_119#_M1025_g N_A_1235_119#_M1002_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0462 AS=0.0609 PD=0.64 PS=0.71 NRD=25.7873 NRS=7.0329 M=1
+ R=2.33333 SA=90000.7 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1033 N_VPWR_M1033_d N_A_1383_349#_M1033_g A_1339_457# VPB PSHORT L=0.18 W=0.42
+ AD=0.132537 AS=0.0462 PD=1.13 PS=0.64 NRD=122.199 NRS=25.7873 M=1 R=2.33333
+ SA=90001.1 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1013 N_A_1235_119#_M1013_d N_RESET_B_M1013_g N_VPWR_M1033_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1176 AS=0.132537 PD=1.4 PS=1.13 NRD=0 NRS=122.199 M=1 R=2.33333
+ SA=90001.7 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1006 N_A_1383_349#_M1006_d N_A_1235_119#_M1006_g N_VPWR_M1006_s VPB PSHORT
+ L=0.18 W=1 AD=0.233775 AS=0.26185 PD=1.535 PS=2.56 NRD=15.7403 NRS=0 M=1
+ R=5.55556 SA=90000.2 SB=90001.4 A=0.18 P=2.36 MULT=1
MM1020 N_A_1824_74#_M1020_d N_A_837_119#_M1020_g N_A_1383_349#_M1006_d VPB
+ PSHORT L=0.18 W=1 AD=0.299965 AS=0.233775 PD=2.53521 PS=1.535 NRD=0
+ NRS=16.0752 M=1 R=5.55556 SA=90000.7 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1021 A_2040_508# N_A_1037_119#_M1021_g N_A_1824_74#_M1020_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0441 AS=0.125985 PD=0.63 PS=1.06479 NRD=23.443 NRS=0 M=1 R=2.33333
+ SA=90001.1 SB=90002.5 A=0.0756 P=1.2 MULT=1
MM1005 N_VPWR_M1005_d N_A_2082_446#_M1005_g A_2040_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.1407 AS=0.0441 PD=1.09 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.33333 SA=90001.5
+ SB=90002.1 A=0.0756 P=1.2 MULT=1
MM1019 N_A_2082_446#_M1019_d N_RESET_B_M1019_g N_VPWR_M1005_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0567 AS=0.1407 PD=0.69 PS=1.09 NRD=0 NRS=21.0987 M=1 R=2.33333
+ SA=90002.3 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1024 N_VPWR_M1024_d N_A_1824_74#_M1024_g N_A_2082_446#_M1019_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.106923 AS=0.0567 PD=0.831127 PS=0.69 NRD=37.5088 NRS=0 M=1
+ R=2.33333 SA=90002.8 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1037 N_A_2495_392#_M1037_d N_A_1824_74#_M1037_g N_VPWR_M1024_d VPB PSHORT
+ L=0.18 W=1 AD=0.28 AS=0.254577 PD=2.56 PS=1.97887 NRD=0 NRS=8.8453 M=1
+ R=5.55556 SA=90001.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A_2495_392#_M1001_g N_Q_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1041 N_VPWR_M1041_d N_A_2495_392#_M1041_g N_Q_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3696 AS=0.1512 PD=2.9 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX42_noxref VNB VPB NWDIODE A=27.6292 P=33.52
c_290 VPB 0 1.77162e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__sdfrtp_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__sdfsbp_2.spice
* Created: Wed Sep  2 12:31:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdfsbp_2.pex.spice"
.subckt sky130_fd_sc_ms__sdfsbp_2  VNB VPB SCE D SCD CLK SET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1044 N_VGND_M1044_d N_SCE_M1044_g N_A_27_74#_M1044_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.08925 AS=0.1197 PD=0.845 PS=1.41 NRD=30 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1037 A_229_74# N_A_27_74#_M1037_g N_VGND_M1044_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.08925 PD=0.66 PS=0.845 NRD=18.564 NRS=11.424 M=1 R=2.8
+ SA=75000.8 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1038 N_A_307_74#_M1038_d N_D_M1038_g A_229_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1659 AS=0.0504 PD=1.21 PS=0.66 NRD=137.136 NRS=18.564 M=1 R=2.8
+ SA=75001.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1017 A_495_74# N_SCE_M1017_g N_A_307_74#_M1038_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1659 PD=0.66 PS=1.21 NRD=18.564 NRS=8.568 M=1 R=2.8 SA=75002.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_SCD_M1015_g A_495_74# VNB NLOWVT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1043 N_VGND_M1043_d N_CLK_M1043_g N_A_619_368#_M1043_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1035 N_A_871_74#_M1035_d N_A_619_368#_M1035_g N_VGND_M1043_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1019 N_A_1069_81#_M1019_d N_A_619_368#_M1019_g N_A_307_74#_M1019_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.18375 AS=0.1197 PD=1.295 PS=1.41 NRD=142.848 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1026 A_1274_81# N_A_871_74#_M1026_g N_A_1069_81#_M1019_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.18375 PD=0.66 PS=1.295 NRD=18.564 NRS=27.132 M=1 R=2.8
+ SA=75001.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_A_1252_376#_M1024_g A_1274_81# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1554 AS=0.0504 PD=1.58 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.6
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1013 A_1567_74# N_A_1069_81#_M1013_g N_A_1252_376#_M1013_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_SET_B_M1014_g A_1567_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.189 AS=0.0504 PD=1.74 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.4 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_1069_81#_M1005_g N_A_1794_74#_M1005_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.096 AS=0.2144 PD=0.94 PS=1.95 NRD=3.744 NRS=9.372 M=1
+ R=4.26667 SA=75000.3 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1011 N_VGND_M1005_d N_A_1069_81#_M1011_g N_A_1794_74#_M1011_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.096 AS=0.0896 PD=0.94 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1032 N_A_1794_74#_M1011_s N_A_871_74#_M1032_g N_A_2067_74#_M1032_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=13.116 M=1
+ R=4.26667 SA=75001.1 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1039 N_A_1794_74#_M1039_d N_A_871_74#_M1039_g N_A_2067_74#_M1032_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.2272 AS=0.112 PD=1.99 PS=0.99 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75001.6 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1008 A_2501_74# N_A_619_368#_M1008_g N_A_2067_74#_M1008_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.3759 PD=0.66 PS=2.63 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.8 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1020 A_2579_74# N_A_2513_258#_M1020_g A_2501_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_SET_B_M1021_g A_2579_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0756 AS=0.0504 PD=0.78 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.6
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1040 N_A_2513_258#_M1040_d N_A_2067_74#_M1040_g N_VGND_M1021_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1197 AS=0.0756 PD=1.41 PS=0.78 NRD=0 NRS=22.848 M=1 R=2.8
+ SA=75002.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 N_Q_N_M1023_d N_A_2067_74#_M1023_g N_VGND_M1023_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.111 AS=0.2479 PD=1.04 PS=2.15 NRD=3.24 NRS=8.1 M=1 R=4.93333
+ SA=75000.3 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1025 N_Q_N_M1023_d N_A_2067_74#_M1025_g N_VGND_M1025_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.111 AS=0.2442 PD=1.04 PS=2.14 NRD=0 NRS=7.296 M=1 R=4.93333
+ SA=75000.7 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_A_2067_74#_M1012_g N_A_3177_368#_M1012_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.136394 AS=0.1824 PD=1.0713 PS=1.85 NRD=25.776 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1012_d N_A_3177_368#_M1001_g N_Q_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.157706 AS=0.1036 PD=1.2387 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1022_d N_A_3177_368#_M1022_g N_Q_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_VPWR_M1009_d N_SCE_M1009_g N_A_27_74#_M1009_s VPB PSHORT L=0.18 W=0.64
+ AD=0.1024 AS=0.1792 PD=0.96 PS=1.84 NRD=13.8491 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90002.1 A=0.1152 P=1.64 MULT=1
MM1007 A_223_464# N_SCE_M1007_g N_VPWR_M1009_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.1024 PD=0.88 PS=0.96 NRD=19.9955 NRS=0 M=1 R=3.55556 SA=90000.7
+ SB=90001.6 A=0.1152 P=1.64 MULT=1
MM1033 N_A_307_74#_M1033_d N_D_M1033_g A_223_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.1248 AS=0.0768 PD=1.03 PS=0.88 NRD=16.9223 NRS=19.9955 M=1 R=3.55556
+ SA=90001.1 SB=90001.2 A=0.1152 P=1.64 MULT=1
MM1027 A_421_464# N_A_27_74#_M1027_g N_A_307_74#_M1033_d VPB PSHORT L=0.18
+ W=0.64 AD=0.0768 AS=0.1248 PD=0.88 PS=1.03 NRD=19.9955 NRS=16.9223 M=1
+ R=3.55556 SA=90001.7 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1041 N_VPWR_M1041_d N_SCD_M1041_g A_421_464# VPB PSHORT L=0.18 W=0.64 AD=0.192
+ AS=0.0768 PD=1.88 PS=0.88 NRD=1.5366 NRS=19.9955 M=1 R=3.55556 SA=90002.1
+ SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1036 N_VPWR_M1036_d N_CLK_M1036_g N_A_619_368#_M1036_s VPB PSHORT L=0.18
+ W=1.12 AD=0.364 AS=0.3136 PD=1.77 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1046 N_A_871_74#_M1046_d N_A_619_368#_M1046_g N_VPWR_M1036_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3528 AS=0.364 PD=2.87 PS=1.77 NRD=5.2599 NRS=1.7533 M=1 R=6.22222
+ SA=90001 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1006 N_A_1069_81#_M1006_d N_A_871_74#_M1006_g N_A_307_74#_M1006_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0672 AS=0.1176 PD=0.74 PS=1.4 NRD=21.0987 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90003 A=0.0756 P=1.2 MULT=1
MM1002 A_1204_463# N_A_619_368#_M1002_g N_A_1069_81#_M1006_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0672 PD=0.66 PS=0.74 NRD=30.4759 NRS=0 M=1 R=2.33333
+ SA=90000.7 SB=90002.5 A=0.0756 P=1.2 MULT=1
MM1030 N_VPWR_M1030_d N_A_1252_376#_M1030_g A_1204_463# VPB PSHORT L=0.18 W=0.42
+ AD=0.19005 AS=0.0504 PD=1.325 PS=0.66 NRD=53.9386 NRS=30.4759 M=1 R=2.33333
+ SA=90001.1 SB=90002.1 A=0.0756 P=1.2 MULT=1
MM1042 N_A_1252_376#_M1042_d N_A_1069_81#_M1042_g N_VPWR_M1030_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.0777 AS=0.19005 PD=0.79 PS=1.325 NRD=0 NRS=239.197 M=1
+ R=2.33333 SA=90002.2 SB=90001 A=0.0756 P=1.2 MULT=1
MM1034 N_VPWR_M1034_d N_SET_B_M1034_g N_A_1252_376#_M1042_d VPB PSHORT L=0.18
+ W=0.42 AD=0.2394 AS=0.0777 PD=1.98 PS=0.79 NRD=133.665 NRS=44.5417 M=1
+ R=2.33333 SA=90002.7 SB=90000.5 A=0.0756 P=1.2 MULT=1
MM1003 N_A_1789_424#_M1003_d N_A_1069_81#_M1003_g N_VPWR_M1003_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.2772 AS=0.1134 PD=2.34 PS=1.11 NRD=10.5395 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90001.5 A=0.1512 P=2.04 MULT=1
MM1048 N_A_1789_424#_M1048_d N_A_1069_81#_M1048_g N_VPWR_M1003_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1134 AS=0.1134 PD=1.11 PS=1.11 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90000.7 SB=90001.1 A=0.1512 P=2.04 MULT=1
MM1028 N_A_2067_74#_M1028_d N_A_619_368#_M1028_g N_A_1789_424#_M1048_d VPB
+ PSHORT L=0.18 W=0.84 AD=0.1134 AS=0.1134 PD=1.11 PS=1.11 NRD=0 NRS=0 M=1
+ R=4.66667 SA=90001.1 SB=90000.6 A=0.1512 P=2.04 MULT=1
MM1031 N_A_2067_74#_M1028_d N_A_619_368#_M1031_g N_A_1789_424#_M1031_s VPB
+ PSHORT L=0.18 W=0.84 AD=0.1134 AS=0.2352 PD=1.11 PS=2.24 NRD=0 NRS=0 M=1
+ R=4.66667 SA=90001.6 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1010 N_A_2067_74#_M1010_d N_A_871_74#_M1010_g N_A_2277_455#_M1010_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.1176 AS=0.1197 PD=1.4 PS=1.41 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1016 N_VPWR_M1016_d N_A_2513_258#_M1016_g N_A_2277_455#_M1016_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0567 AS=0.1176 PD=0.69 PS=1.4 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1018 N_A_2067_74#_M1018_d N_SET_B_M1018_g N_VPWR_M1016_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1176 AS=0.0567 PD=1.4 PS=0.69 NRD=0 NRS=0 M=1 R=2.33333 SA=90000.6
+ SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1045 N_VPWR_M1045_d N_A_2067_74#_M1045_g N_A_2513_258#_M1045_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0941182 AS=0.1176 PD=0.804545 PS=1.4 NRD=105.533 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1004 N_Q_N_M1004_d N_A_2067_74#_M1004_g N_VPWR_M1045_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.250982 PD=1.39 PS=2.14545 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.4 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1029 N_Q_N_M1004_d N_A_2067_74#_M1029_g N_VPWR_M1029_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.8
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_2067_74#_M1000_g N_A_3177_368#_M1000_s VPB PSHORT
+ L=0.18 W=1 AD=0.190377 AS=0.28 PD=1.40566 PS=2.56 NRD=19.0302 NRS=0 M=1
+ R=5.55556 SA=90000.2 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1047 N_Q_M1047_d N_A_3177_368#_M1047_g N_VPWR_M1000_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.213223 PD=1.39 PS=1.57434 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.7
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1049 N_Q_M1047_d N_A_3177_368#_M1049_g N_VPWR_M1049_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX50_noxref VNB VPB NWDIODE A=33.7404 P=40
c_356 VPB 0 1.49424e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__sdfsbp_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__a221o_4.spice
* Created: Fri Aug 28 17:00:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a221o_4.pex.spice"
.subckt sky130_fd_sc_ms__a221o_4  VNB VPB A1 A2 C1 B2 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* B2	B2
* C1	C1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1009 N_A_154_135#_M1009_d N_A1_M1009_g N_A_71_135#_M1009_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1011 N_A_154_135#_M1009_d N_A1_M1011_g N_A_71_135#_M1011_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1022 N_A_71_135#_M1022_d N_A2_M1022_g N_VGND_M1022_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75004.7 A=0.096 P=1.58 MULT=1
MM1027 N_A_71_135#_M1022_d N_A2_M1027_g N_VGND_M1027_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.114423 PD=0.92 PS=1.01565 NRD=0 NRS=12.18 M=1 R=4.26667
+ SA=75000.6 SB=75004.3 A=0.096 P=1.58 MULT=1
MM1005 N_X_M1005_d N_A_154_135#_M1005_g N_VGND_M1027_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.132302 PD=1.02 PS=1.17435 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1015 N_X_M1005_d N_A_154_135#_M1015_g N_VGND_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.4
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1021 N_X_M1021_d N_A_154_135#_M1021_g N_VGND_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.8
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1023 N_X_M1021_d N_A_154_135#_M1023_g N_VGND_M1023_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.26817 PD=1.02 PS=1.58725 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1024 N_A_154_135#_M1024_d N_C1_M1024_g N_VGND_M1023_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.23193 PD=0.92 PS=1.37275 NRD=0 NRS=0 M=1 R=4.26667 SA=75003.3
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1025 N_A_154_135#_M1024_d N_C1_M1025_g N_VGND_M1025_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1648 PD=0.92 PS=1.17 NRD=0 NRS=30.468 M=1 R=4.26667 SA=75003.7
+ SB=75001.3 A=0.096 P=1.58 MULT=1
MM1017 N_A_1346_123#_M1017_d N_B2_M1017_g N_VGND_M1025_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1648 PD=0.92 PS=1.17 NRD=0 NRS=13.584 M=1 R=4.26667
+ SA=75004.3 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1019 N_A_1346_123#_M1017_d N_B2_M1019_g N_VGND_M1019_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75004.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1012 N_A_154_135#_M1012_d N_B1_M1012_g N_A_1346_123#_M1012_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1020 N_A_154_135#_M1012_d N_B1_M1020_g N_A_1346_123#_M1020_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.2144 PD=0.92 PS=1.95 NRD=0 NRS=4.68 M=1 R=4.26667
+ SA=75000.6 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1016 N_VPWR_M1016_d N_A1_M1016_g N_A_160_376#_M1016_s VPB PSHORT L=0.18 W=1
+ AD=0.26 AS=0.195 PD=2.52 PS=1.39 NRD=0 NRS=22.6353 M=1 R=5.55556 SA=90000.2
+ SB=90004 A=0.18 P=2.36 MULT=1
MM1018 N_VPWR_M1018_d N_A1_M1018_g N_A_160_376#_M1016_s VPB PSHORT L=0.18 W=1
+ AD=0.3575 AS=0.195 PD=1.715 PS=1.39 NRD=9.8303 NRS=0 M=1 R=5.55556 SA=90000.7
+ SB=90003.5 A=0.18 P=2.36 MULT=1
MM1001 N_A_160_376#_M1001_d N_A2_M1001_g N_VPWR_M1018_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.3575 PD=1.27 PS=1.715 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90001.6
+ SB=90002.6 A=0.18 P=2.36 MULT=1
MM1003 N_A_160_376#_M1001_d N_A2_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.217547 PD=1.27 PS=1.46226 NRD=0 NRS=31.52 M=1 R=5.55556
+ SA=90002.1 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1006 N_X_M1006_d N_A_154_135#_M1006_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.243653 PD=1.39 PS=1.63774 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.4
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1008 N_X_M1006_d N_A_154_135#_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.9
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1010 N_X_M1010_d N_A_154_135#_M1010_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.3
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1013 N_X_M1010_d N_A_154_135#_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.8
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1000 N_A_1102_392#_M1000_d N_C1_M1000_g N_A_154_135#_M1000_s VPB PSHORT L=0.18
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90002.7 A=0.18 P=2.36 MULT=1
MM1026 N_A_1102_392#_M1026_d N_C1_M1026_g N_A_154_135#_M1000_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.6
+ SB=90002.3 A=0.18 P=2.36 MULT=1
MM1002 N_A_160_376#_M1002_d N_B2_M1002_g N_A_1102_392#_M1026_d VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.1
+ SB=90001.8 A=0.18 P=2.36 MULT=1
MM1004 N_A_160_376#_M1002_d N_B2_M1004_g N_A_1102_392#_M1004_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.28 PD=1.27 PS=1.56 NRD=0 NRS=29.55 M=1 R=5.55556 SA=90001.5
+ SB=90001.4 A=0.18 P=2.36 MULT=1
MM1007 N_A_160_376#_M1007_d N_B1_M1007_g N_A_1102_392#_M1004_s VPB PSHORT L=0.18
+ W=1 AD=0.155 AS=0.28 PD=1.31 PS=1.56 NRD=2.9353 NRS=25.5903 M=1 R=5.55556
+ SA=90002.3 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1014 N_A_160_376#_M1007_d N_B1_M1014_g N_A_1102_392#_M1014_s VPB PSHORT L=0.18
+ W=1 AD=0.155 AS=0.26 PD=1.31 PS=2.52 NRD=2.9353 NRS=0 M=1 R=5.55556 SA=90002.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX28_noxref VNB VPB NWDIODE A=18.5628 P=23.68
c_155 VPB 0 2.11319e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__a221o_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__maj3_2.pxi.spice
* Created: Wed Sep  2 12:11:25 2020
* 
x_PM_SKY130_FD_SC_MS__MAJ3_2%A_87_264# N_A_87_264#_M1009_d N_A_87_264#_M1013_d
+ N_A_87_264#_M1007_d N_A_87_264#_M1015_d N_A_87_264#_M1004_g
+ N_A_87_264#_M1011_g N_A_87_264#_M1014_g N_A_87_264#_M1005_g N_A_87_264#_c_91_n
+ N_A_87_264#_c_83_n N_A_87_264#_c_84_n N_A_87_264#_c_102_p N_A_87_264#_c_85_n
+ N_A_87_264#_c_93_n N_A_87_264#_c_94_n N_A_87_264#_c_86_n N_A_87_264#_c_87_n
+ N_A_87_264#_c_88_n N_A_87_264#_c_96_n PM_SKY130_FD_SC_MS__MAJ3_2%A_87_264#
x_PM_SKY130_FD_SC_MS__MAJ3_2%B N_B_M1009_g N_B_M1007_g N_B_M1002_g N_B_M1010_g B
+ N_B_c_215_n N_B_c_216_n PM_SKY130_FD_SC_MS__MAJ3_2%B
x_PM_SKY130_FD_SC_MS__MAJ3_2%C N_C_M1003_g N_C_M1001_g N_C_M1013_g N_C_M1015_g
+ N_C_c_261_n N_C_c_262_n C N_C_c_263_n N_C_c_264_n PM_SKY130_FD_SC_MS__MAJ3_2%C
x_PM_SKY130_FD_SC_MS__MAJ3_2%A N_A_M1000_g N_A_c_321_n N_A_M1008_g N_A_c_328_n
+ N_A_c_329_n N_A_c_322_n N_A_M1006_g N_A_M1012_g N_A_c_324_n N_A_c_325_n A
+ PM_SKY130_FD_SC_MS__MAJ3_2%A
x_PM_SKY130_FD_SC_MS__MAJ3_2%VPWR N_VPWR_M1004_d N_VPWR_M1005_d N_VPWR_M1001_d
+ N_VPWR_c_391_n N_VPWR_c_392_n N_VPWR_c_393_n N_VPWR_c_394_n VPWR
+ N_VPWR_c_395_n N_VPWR_c_396_n N_VPWR_c_397_n N_VPWR_c_390_n N_VPWR_c_399_n
+ N_VPWR_c_400_n PM_SKY130_FD_SC_MS__MAJ3_2%VPWR
x_PM_SKY130_FD_SC_MS__MAJ3_2%X N_X_M1011_s N_X_M1004_s N_X_c_438_n N_X_c_439_n X
+ X X X N_X_c_440_n PM_SKY130_FD_SC_MS__MAJ3_2%X
x_PM_SKY130_FD_SC_MS__MAJ3_2%VGND N_VGND_M1011_d N_VGND_M1014_d N_VGND_M1003_d
+ N_VGND_c_473_n N_VGND_c_474_n N_VGND_c_475_n N_VGND_c_476_n VGND
+ N_VGND_c_477_n N_VGND_c_478_n N_VGND_c_479_n N_VGND_c_480_n N_VGND_c_481_n
+ N_VGND_c_482_n PM_SKY130_FD_SC_MS__MAJ3_2%VGND
cc_1 VNB N_A_87_264#_M1004_g 7.19436e-19 $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.4
cc_2 VNB N_A_87_264#_M1011_g 0.0275446f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_3 VNB N_A_87_264#_M1014_g 0.0258102f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=0.74
cc_4 VNB N_A_87_264#_M1005_g 5.17345e-19 $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.4
cc_5 VNB N_A_87_264#_c_83_n 0.00315813f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=1.78
cc_6 VNB N_A_87_264#_c_84_n 0.0153736f $X=-0.19 $Y=-0.245 $X2=4.33 $Y2=0.99
cc_7 VNB N_A_87_264#_c_85_n 0.0237216f $X=-0.19 $Y=-0.245 $X2=4.495 $Y2=0.515
cc_8 VNB N_A_87_264#_c_86_n 0.00814668f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.485
cc_9 VNB N_A_87_264#_c_87_n 0.0662865f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.485
cc_10 VNB N_A_87_264#_c_88_n 0.00446828f $X=-0.19 $Y=-0.245 $X2=2.76 $Y2=0.712
cc_11 VNB N_B_M1009_g 0.0182529f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=1.735
cc_12 VNB N_B_M1002_g 0.0193109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B_c_215_n 0.00176754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B_c_216_n 0.0387324f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.65
cc_15 VNB N_C_M1003_g 0.020459f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=1.735
cc_16 VNB N_C_M1013_g 0.0299104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_C_M1015_g 0.00245727f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.4
cc_18 VNB N_C_c_261_n 0.0202004f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_19 VNB N_C_c_262_n 0.0328125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_C_c_263_n 0.0255377f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.65
cc_21 VNB N_C_c_264_n 0.00433354f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.4
cc_22 VNB N_A_M1000_g 0.00402508f $X=-0.19 $Y=-0.245 $X2=4.385 $Y2=1.84
cc_23 VNB N_A_c_321_n 0.0193072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_c_322_n 0.00137966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_M1012_g 0.0343707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_c_324_n 0.0375928f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_27 VNB N_A_c_325_n 0.021884f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_28 VNB A 0.0072112f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.32
cc_29 VNB N_VPWR_c_390_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_X_c_438_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_439_n 0.00429968f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.65
cc_32 VNB N_X_c_440_n 0.00139976f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=1.78
cc_33 VNB N_VGND_c_473_n 0.011316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_474_n 0.0505285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_475_n 0.0141402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_476_n 0.00492322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_477_n 0.0192531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_478_n 0.042745f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=1.865
cc_39 VNB N_VGND_c_479_n 0.0299721f $X=-0.19 $Y=-0.245 $X2=4.495 $Y2=0.515
cc_40 VNB N_VGND_c_480_n 0.29124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_481_n 0.013849f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.485
cc_42 VNB N_VGND_c_482_n 0.00923827f $X=-0.19 $Y=-0.245 $X2=2.595 $Y2=0.712
cc_43 VPB N_A_87_264#_M1004_g 0.0274013f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.4
cc_44 VPB N_A_87_264#_M1005_g 0.0238269f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=2.4
cc_45 VPB N_A_87_264#_c_91_n 0.0100301f $X=-0.19 $Y=1.66 $X2=1.965 $Y2=1.865
cc_46 VPB N_A_87_264#_c_83_n 0.00108141f $X=-0.19 $Y=1.66 $X2=2.05 $Y2=1.78
cc_47 VPB N_A_87_264#_c_93_n 0.0191391f $X=-0.19 $Y=1.66 $X2=4.52 $Y2=2.12
cc_48 VPB N_A_87_264#_c_94_n 0.0312613f $X=-0.19 $Y=1.66 $X2=4.52 $Y2=2.695
cc_49 VPB N_A_87_264#_c_86_n 0.00311091f $X=-0.19 $Y=1.66 $X2=1.06 $Y2=1.485
cc_50 VPB N_A_87_264#_c_96_n 0.00280657f $X=-0.19 $Y=1.66 $X2=2.375 $Y2=2.035
cc_51 VPB N_B_M1007_g 0.0185435f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_B_M1010_g 0.0173313f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.4
cc_53 VPB N_B_c_215_n 0.00113295f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_B_c_216_n 0.00590114f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.65
cc_55 VPB N_C_M1001_g 0.019787f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_C_M1015_g 0.0304773f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.4
cc_57 VPB N_C_c_261_n 9.84389e-19 $X=-0.19 $Y=1.66 $X2=0.515 $Y2=0.74
cc_58 VPB N_C_c_263_n 0.00560401f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.65
cc_59 VPB N_C_c_264_n 0.00235698f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=2.4
cc_60 VPB N_A_M1000_g 0.0341458f $X=-0.19 $Y=1.66 $X2=4.385 $Y2=1.84
cc_61 VPB N_A_c_328_n 0.146924f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_c_329_n 0.0139998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_c_322_n 0.00465897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_M1006_g 0.0261431f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.65
cc_65 VPB N_A_M1012_g 0.00103027f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_391_n 0.0112901f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_392_n 0.0644823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_393_n 0.0168953f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=0.74
cc_69 VPB N_VPWR_c_394_n 0.00880679f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_395_n 0.0194151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_396_n 0.049034f $X=-0.19 $Y=1.66 $X2=4.33 $Y2=0.99
cc_72 VPB N_VPWR_c_397_n 0.0304171f $X=-0.19 $Y=1.66 $X2=4.52 $Y2=2.695
cc_73 VPB N_VPWR_c_390_n 0.0675307f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_399_n 0.0133423f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_400_n 0.00435574f $X=-0.19 $Y=1.66 $X2=2.76 $Y2=0.712
cc_76 VPB X 0.00446143f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.4
cc_77 VPB X 0.00231613f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=0.74
cc_78 VPB N_X_c_440_n 8.5093e-19 $X=-0.19 $Y=1.66 $X2=2.05 $Y2=1.78
cc_79 N_A_87_264#_c_83_n N_B_M1009_g 0.00680221f $X=2.05 $Y=1.78 $X2=0 $Y2=0
cc_80 N_A_87_264#_c_88_n N_B_M1009_g 0.0214115f $X=2.76 $Y=0.712 $X2=0 $Y2=0
cc_81 N_A_87_264#_c_96_n N_B_M1007_g 0.0351229f $X=2.375 $Y=2.035 $X2=0 $Y2=0
cc_82 N_A_87_264#_c_84_n N_B_M1002_g 0.0112064f $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_83 N_A_87_264#_c_88_n N_B_M1002_g 0.0119906f $X=2.76 $Y=0.712 $X2=0 $Y2=0
cc_84 N_A_87_264#_c_102_p N_B_M1010_g 0.0129464f $X=4.355 $Y=2.035 $X2=0 $Y2=0
cc_85 N_A_87_264#_c_96_n N_B_M1010_g 0.0156821f $X=2.375 $Y=2.035 $X2=0 $Y2=0
cc_86 N_A_87_264#_M1007_d N_B_c_215_n 0.00171375f $X=2.485 $Y=1.735 $X2=0 $Y2=0
cc_87 N_A_87_264#_c_83_n N_B_c_215_n 0.0423661f $X=2.05 $Y=1.78 $X2=0 $Y2=0
cc_88 N_A_87_264#_c_102_p N_B_c_215_n 0.0111658f $X=4.355 $Y=2.035 $X2=0 $Y2=0
cc_89 N_A_87_264#_c_88_n N_B_c_215_n 0.0472156f $X=2.76 $Y=0.712 $X2=0 $Y2=0
cc_90 N_A_87_264#_c_96_n N_B_c_215_n 0.0311098f $X=2.375 $Y=2.035 $X2=0 $Y2=0
cc_91 N_A_87_264#_c_84_n N_B_c_216_n 4.98325e-19 $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_92 N_A_87_264#_c_88_n N_B_c_216_n 7.88032e-19 $X=2.76 $Y=0.712 $X2=0 $Y2=0
cc_93 N_A_87_264#_c_96_n N_B_c_216_n 4.43633e-19 $X=2.375 $Y=2.035 $X2=0 $Y2=0
cc_94 N_A_87_264#_c_84_n N_C_M1003_g 0.0151982f $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_95 N_A_87_264#_c_88_n N_C_M1003_g 0.0020622f $X=2.76 $Y=0.712 $X2=0 $Y2=0
cc_96 N_A_87_264#_c_102_p N_C_M1001_g 0.0177071f $X=4.355 $Y=2.035 $X2=0 $Y2=0
cc_97 N_A_87_264#_c_96_n N_C_M1001_g 0.00298595f $X=2.375 $Y=2.035 $X2=0 $Y2=0
cc_98 N_A_87_264#_c_84_n N_C_M1013_g 0.0130655f $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_99 N_A_87_264#_c_85_n N_C_M1013_g 0.0112749f $X=4.495 $Y=0.515 $X2=0 $Y2=0
cc_100 N_A_87_264#_c_102_p N_C_M1015_g 0.0135388f $X=4.355 $Y=2.035 $X2=0 $Y2=0
cc_101 N_A_87_264#_c_93_n N_C_M1015_g 0.00374487f $X=4.52 $Y=2.12 $X2=0 $Y2=0
cc_102 N_A_87_264#_c_94_n N_C_M1015_g 0.0144609f $X=4.52 $Y=2.695 $X2=0 $Y2=0
cc_103 N_A_87_264#_c_84_n N_C_c_261_n 0.0494717f $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_104 N_A_87_264#_c_102_p N_C_c_261_n 0.0256836f $X=4.355 $Y=2.035 $X2=0 $Y2=0
cc_105 N_A_87_264#_c_93_n N_C_c_261_n 0.0138249f $X=4.52 $Y=2.12 $X2=0 $Y2=0
cc_106 N_A_87_264#_c_84_n N_C_c_262_n 0.00431154f $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_107 N_A_87_264#_c_93_n N_C_c_262_n 0.00345942f $X=4.52 $Y=2.12 $X2=0 $Y2=0
cc_108 N_A_87_264#_c_84_n N_C_c_263_n 0.00114171f $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_109 N_A_87_264#_c_102_p N_C_c_263_n 5.69919e-19 $X=4.355 $Y=2.035 $X2=0 $Y2=0
cc_110 N_A_87_264#_c_84_n N_C_c_264_n 0.0366919f $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_111 N_A_87_264#_c_102_p N_C_c_264_n 0.0343866f $X=4.355 $Y=2.035 $X2=0 $Y2=0
cc_112 N_A_87_264#_c_91_n N_A_M1000_g 0.0208764f $X=1.965 $Y=1.865 $X2=0 $Y2=0
cc_113 N_A_87_264#_c_83_n N_A_M1000_g 0.0110075f $X=2.05 $Y=1.78 $X2=0 $Y2=0
cc_114 N_A_87_264#_c_86_n N_A_M1000_g 0.00480836f $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_115 N_A_87_264#_c_87_n N_A_M1000_g 0.00154813f $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_116 N_A_87_264#_c_96_n N_A_M1000_g 0.0276851f $X=2.375 $Y=2.035 $X2=0 $Y2=0
cc_117 N_A_87_264#_c_83_n N_A_c_321_n 0.00640847f $X=2.05 $Y=1.78 $X2=0 $Y2=0
cc_118 N_A_87_264#_c_88_n N_A_c_321_n 0.0224413f $X=2.76 $Y=0.712 $X2=0 $Y2=0
cc_119 N_A_87_264#_c_96_n N_A_c_328_n 0.0108552f $X=2.375 $Y=2.035 $X2=0 $Y2=0
cc_120 N_A_87_264#_c_102_p N_A_M1006_g 0.0176459f $X=4.355 $Y=2.035 $X2=0 $Y2=0
cc_121 N_A_87_264#_c_93_n N_A_M1006_g 6.25758e-19 $X=4.52 $Y=2.12 $X2=0 $Y2=0
cc_122 N_A_87_264#_c_94_n N_A_M1006_g 0.00243009f $X=4.52 $Y=2.695 $X2=0 $Y2=0
cc_123 N_A_87_264#_c_84_n N_A_M1012_g 0.0152913f $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_124 N_A_87_264#_c_85_n N_A_M1012_g 0.00204644f $X=4.495 $Y=0.515 $X2=0 $Y2=0
cc_125 N_A_87_264#_M1014_g N_A_c_324_n 0.00312895f $X=0.945 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A_87_264#_c_91_n N_A_c_324_n 0.00236155f $X=1.965 $Y=1.865 $X2=0 $Y2=0
cc_127 N_A_87_264#_c_86_n N_A_c_324_n 0.00152219f $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_128 N_A_87_264#_c_87_n N_A_c_324_n 0.0128112f $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_129 N_A_87_264#_c_83_n N_A_c_325_n 0.0111192f $X=2.05 $Y=1.78 $X2=0 $Y2=0
cc_130 N_A_87_264#_M1014_g A 0.00166385f $X=0.945 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A_87_264#_c_91_n A 0.0199019f $X=1.965 $Y=1.865 $X2=0 $Y2=0
cc_132 N_A_87_264#_c_83_n A 0.0265523f $X=2.05 $Y=1.78 $X2=0 $Y2=0
cc_133 N_A_87_264#_c_86_n A 0.0157135f $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_134 N_A_87_264#_c_87_n A 2.7436e-19 $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_135 N_A_87_264#_c_91_n N_VPWR_M1005_d 0.00737298f $X=1.965 $Y=1.865 $X2=0
+ $Y2=0
cc_136 N_A_87_264#_c_86_n N_VPWR_M1005_d 0.00227816f $X=1.06 $Y=1.485 $X2=0
+ $Y2=0
cc_137 N_A_87_264#_c_102_p N_VPWR_M1001_d 0.00693378f $X=4.355 $Y=2.035 $X2=0
+ $Y2=0
cc_138 N_A_87_264#_M1004_g N_VPWR_c_392_n 0.00647357f $X=0.525 $Y=2.4 $X2=0
+ $Y2=0
cc_139 N_A_87_264#_M1005_g N_VPWR_c_393_n 0.00863415f $X=0.975 $Y=2.4 $X2=0
+ $Y2=0
cc_140 N_A_87_264#_c_91_n N_VPWR_c_393_n 0.0396665f $X=1.965 $Y=1.865 $X2=0
+ $Y2=0
cc_141 N_A_87_264#_c_86_n N_VPWR_c_393_n 0.011924f $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_142 N_A_87_264#_c_87_n N_VPWR_c_393_n 5.13368e-19 $X=1.06 $Y=1.485 $X2=0
+ $Y2=0
cc_143 N_A_87_264#_c_102_p N_VPWR_c_394_n 0.0218557f $X=4.355 $Y=2.035 $X2=0
+ $Y2=0
cc_144 N_A_87_264#_c_94_n N_VPWR_c_394_n 0.0165748f $X=4.52 $Y=2.695 $X2=0 $Y2=0
cc_145 N_A_87_264#_M1004_g N_VPWR_c_395_n 0.0048691f $X=0.525 $Y=2.4 $X2=0 $Y2=0
cc_146 N_A_87_264#_M1005_g N_VPWR_c_395_n 0.005209f $X=0.975 $Y=2.4 $X2=0 $Y2=0
cc_147 N_A_87_264#_c_96_n N_VPWR_c_396_n 0.0174863f $X=2.375 $Y=2.035 $X2=0
+ $Y2=0
cc_148 N_A_87_264#_c_94_n N_VPWR_c_397_n 0.00975961f $X=4.52 $Y=2.695 $X2=0
+ $Y2=0
cc_149 N_A_87_264#_M1004_g N_VPWR_c_390_n 0.00876015f $X=0.525 $Y=2.4 $X2=0
+ $Y2=0
cc_150 N_A_87_264#_M1005_g N_VPWR_c_390_n 0.00986727f $X=0.975 $Y=2.4 $X2=0
+ $Y2=0
cc_151 N_A_87_264#_c_94_n N_VPWR_c_390_n 0.0111753f $X=4.52 $Y=2.695 $X2=0 $Y2=0
cc_152 N_A_87_264#_c_96_n N_VPWR_c_390_n 0.0224582f $X=2.375 $Y=2.035 $X2=0
+ $Y2=0
cc_153 N_A_87_264#_M1011_g N_X_c_438_n 0.0081896f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A_87_264#_M1014_g N_X_c_438_n 0.00783249f $X=0.945 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A_87_264#_M1011_g N_X_c_439_n 0.00215589f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A_87_264#_M1014_g N_X_c_439_n 0.00723846f $X=0.945 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A_87_264#_c_87_n N_X_c_439_n 0.00239209f $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_158 N_A_87_264#_M1004_g X 0.00270934f $X=0.525 $Y=2.4 $X2=0 $Y2=0
cc_159 N_A_87_264#_M1005_g X 0.00476645f $X=0.975 $Y=2.4 $X2=0 $Y2=0
cc_160 N_A_87_264#_c_86_n X 0.00737712f $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_161 N_A_87_264#_c_87_n X 0.00317005f $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_162 N_A_87_264#_M1004_g X 0.0149161f $X=0.525 $Y=2.4 $X2=0 $Y2=0
cc_163 N_A_87_264#_M1005_g X 0.0164918f $X=0.975 $Y=2.4 $X2=0 $Y2=0
cc_164 N_A_87_264#_M1004_g N_X_c_440_n 0.00894847f $X=0.525 $Y=2.4 $X2=0 $Y2=0
cc_165 N_A_87_264#_M1011_g N_X_c_440_n 0.00963174f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A_87_264#_M1014_g N_X_c_440_n 0.00298176f $X=0.945 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A_87_264#_M1005_g N_X_c_440_n 9.33303e-19 $X=0.975 $Y=2.4 $X2=0 $Y2=0
cc_168 N_A_87_264#_c_86_n N_X_c_440_n 0.0292291f $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_169 N_A_87_264#_c_87_n N_X_c_440_n 0.0238411f $X=1.06 $Y=1.485 $X2=0 $Y2=0
cc_170 N_A_87_264#_c_83_n A_396_368# 3.68242e-19 $X=2.05 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_171 N_A_87_264#_c_96_n A_396_368# 0.0100999f $X=2.375 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_172 N_A_87_264#_c_102_p A_587_347# 0.0126676f $X=4.355 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_173 N_A_87_264#_c_102_p A_793_368# 0.00660859f $X=4.355 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_174 N_A_87_264#_c_84_n N_VGND_M1003_d 0.00817304f $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_175 N_A_87_264#_M1011_g N_VGND_c_474_n 0.00646793f $X=0.515 $Y=0.74 $X2=0
+ $Y2=0
cc_176 N_A_87_264#_M1014_g N_VGND_c_475_n 0.00552888f $X=0.945 $Y=0.74 $X2=0
+ $Y2=0
cc_177 N_A_87_264#_c_86_n N_VGND_c_475_n 0.00986737f $X=1.06 $Y=1.485 $X2=0
+ $Y2=0
cc_178 N_A_87_264#_c_87_n N_VGND_c_475_n 0.00109081f $X=1.06 $Y=1.485 $X2=0
+ $Y2=0
cc_179 N_A_87_264#_c_88_n N_VGND_c_475_n 0.0576083f $X=2.76 $Y=0.712 $X2=0 $Y2=0
cc_180 N_A_87_264#_c_84_n N_VGND_c_476_n 0.0251177f $X=4.33 $Y=0.99 $X2=0 $Y2=0
cc_181 N_A_87_264#_c_85_n N_VGND_c_476_n 0.0107976f $X=4.495 $Y=0.515 $X2=0
+ $Y2=0
cc_182 N_A_87_264#_c_88_n N_VGND_c_476_n 0.00980679f $X=2.76 $Y=0.712 $X2=0
+ $Y2=0
cc_183 N_A_87_264#_M1011_g N_VGND_c_477_n 0.00422942f $X=0.515 $Y=0.74 $X2=0
+ $Y2=0
cc_184 N_A_87_264#_M1014_g N_VGND_c_477_n 0.00434272f $X=0.945 $Y=0.74 $X2=0
+ $Y2=0
cc_185 N_A_87_264#_c_88_n N_VGND_c_478_n 0.0345112f $X=2.76 $Y=0.712 $X2=0 $Y2=0
cc_186 N_A_87_264#_c_85_n N_VGND_c_479_n 0.0145639f $X=4.495 $Y=0.515 $X2=0
+ $Y2=0
cc_187 N_A_87_264#_M1011_g N_VGND_c_480_n 0.00787322f $X=0.515 $Y=0.74 $X2=0
+ $Y2=0
cc_188 N_A_87_264#_M1014_g N_VGND_c_480_n 0.00825283f $X=0.945 $Y=0.74 $X2=0
+ $Y2=0
cc_189 N_A_87_264#_c_85_n N_VGND_c_480_n 0.0119984f $X=4.495 $Y=0.515 $X2=0
+ $Y2=0
cc_190 N_A_87_264#_c_88_n N_VGND_c_480_n 0.0280173f $X=2.76 $Y=0.712 $X2=0 $Y2=0
cc_191 N_A_87_264#_c_83_n A_413_74# 4.41425e-19 $X=2.05 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_192 N_A_87_264#_c_88_n A_413_74# 0.00517808f $X=2.76 $Y=0.712 $X2=-0.19
+ $Y2=-0.245
cc_193 N_A_87_264#_c_84_n A_577_74# 0.0155294f $X=4.33 $Y=0.99 $X2=-0.19
+ $Y2=-0.245
cc_194 N_A_87_264#_c_84_n A_793_74# 0.00632546f $X=4.33 $Y=0.99 $X2=-0.19
+ $Y2=-0.245
cc_195 N_B_M1002_g N_C_M1003_g 0.0375136f $X=2.81 $Y=0.74 $X2=0 $Y2=0
cc_196 N_B_M1010_g N_C_M1001_g 0.058442f $X=2.845 $Y=2.235 $X2=0 $Y2=0
cc_197 N_B_c_215_n N_C_M1001_g 0.00119256f $X=2.81 $Y=1.41 $X2=0 $Y2=0
cc_198 N_B_c_215_n N_C_c_263_n 0.00121114f $X=2.81 $Y=1.41 $X2=0 $Y2=0
cc_199 N_B_c_216_n N_C_c_263_n 0.0180484f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_200 N_B_M1010_g N_C_c_264_n 2.46331e-19 $X=2.845 $Y=2.235 $X2=0 $Y2=0
cc_201 N_B_c_215_n N_C_c_264_n 0.0324723f $X=2.81 $Y=1.41 $X2=0 $Y2=0
cc_202 N_B_c_216_n N_C_c_264_n 0.00138848f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_203 N_B_c_215_n N_A_M1000_g 2.30641e-19 $X=2.81 $Y=1.41 $X2=0 $Y2=0
cc_204 N_B_c_216_n N_A_M1000_g 0.0478998f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_205 N_B_M1009_g N_A_c_321_n 0.0355006f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_206 N_B_M1007_g N_A_c_328_n 0.0116292f $X=2.395 $Y=2.235 $X2=0 $Y2=0
cc_207 N_B_M1010_g N_A_c_328_n 0.0123546f $X=2.845 $Y=2.235 $X2=0 $Y2=0
cc_208 N_B_c_215_n N_A_c_325_n 3.322e-19 $X=2.81 $Y=1.41 $X2=0 $Y2=0
cc_209 N_B_c_216_n N_A_c_325_n 0.0355006f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_210 N_B_M1007_g N_VPWR_c_390_n 0.00112709f $X=2.395 $Y=2.235 $X2=0 $Y2=0
cc_211 N_B_M1010_g N_VPWR_c_390_n 0.00112709f $X=2.845 $Y=2.235 $X2=0 $Y2=0
cc_212 N_B_M1002_g N_VGND_c_476_n 0.00153831f $X=2.81 $Y=0.74 $X2=0 $Y2=0
cc_213 N_B_M1009_g N_VGND_c_478_n 0.00291649f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_214 N_B_M1002_g N_VGND_c_478_n 0.00433162f $X=2.81 $Y=0.74 $X2=0 $Y2=0
cc_215 N_B_M1009_g N_VGND_c_480_n 0.00358831f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_216 N_B_M1002_g N_VGND_c_480_n 0.00818163f $X=2.81 $Y=0.74 $X2=0 $Y2=0
cc_217 N_C_M1001_g N_A_c_328_n 0.0124996f $X=3.305 $Y=2.235 $X2=0 $Y2=0
cc_218 N_C_M1001_g N_A_c_322_n 0.0268814f $X=3.305 $Y=2.235 $X2=0 $Y2=0
cc_219 N_C_c_261_n N_A_c_322_n 0.00467468f $X=4.37 $Y=1.465 $X2=0 $Y2=0
cc_220 N_C_c_262_n N_A_c_322_n 0.0484282f $X=4.37 $Y=1.465 $X2=0 $Y2=0
cc_221 N_C_c_264_n N_A_c_322_n 0.00462228f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_222 N_C_M1015_g N_A_M1006_g 0.0484282f $X=4.295 $Y=2.34 $X2=0 $Y2=0
cc_223 N_C_M1003_g N_A_M1012_g 0.027073f $X=3.29 $Y=0.74 $X2=0 $Y2=0
cc_224 N_C_M1001_g N_A_M1012_g 0.00100202f $X=3.305 $Y=2.235 $X2=0 $Y2=0
cc_225 N_C_M1013_g N_A_M1012_g 0.0484282f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_226 N_C_c_261_n N_A_M1012_g 0.0120146f $X=4.37 $Y=1.465 $X2=0 $Y2=0
cc_227 N_C_c_263_n N_A_M1012_g 0.0153368f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_228 N_C_c_264_n N_A_M1012_g 0.00200531f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_229 N_C_c_264_n N_VPWR_M1001_d 0.00216694f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_230 N_C_M1001_g N_VPWR_c_394_n 0.0157974f $X=3.305 $Y=2.235 $X2=0 $Y2=0
cc_231 N_C_M1015_g N_VPWR_c_394_n 0.00214461f $X=4.295 $Y=2.34 $X2=0 $Y2=0
cc_232 N_C_M1015_g N_VPWR_c_397_n 0.00567889f $X=4.295 $Y=2.34 $X2=0 $Y2=0
cc_233 N_C_M1001_g N_VPWR_c_390_n 0.00112709f $X=3.305 $Y=2.235 $X2=0 $Y2=0
cc_234 N_C_M1015_g N_VPWR_c_390_n 0.00610055f $X=4.295 $Y=2.34 $X2=0 $Y2=0
cc_235 N_C_M1003_g N_VGND_c_476_n 0.0164979f $X=3.29 $Y=0.74 $X2=0 $Y2=0
cc_236 N_C_M1013_g N_VGND_c_476_n 0.00149046f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_237 N_C_M1003_g N_VGND_c_478_n 0.00383152f $X=3.29 $Y=0.74 $X2=0 $Y2=0
cc_238 N_C_M1013_g N_VGND_c_479_n 0.00434272f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_239 N_C_M1003_g N_VGND_c_480_n 0.00758084f $X=3.29 $Y=0.74 $X2=0 $Y2=0
cc_240 N_C_M1013_g N_VGND_c_480_n 0.0082472f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_241 N_A_M1000_g N_VPWR_c_393_n 0.0187961f $X=1.89 $Y=2.34 $X2=0 $Y2=0
cc_242 N_A_c_328_n N_VPWR_c_394_n 0.0226039f $X=3.785 $Y=3.15 $X2=0 $Y2=0
cc_243 N_A_M1006_g N_VPWR_c_394_n 0.0221327f $X=3.875 $Y=2.34 $X2=0 $Y2=0
cc_244 N_A_c_329_n N_VPWR_c_396_n 0.0511764f $X=1.98 $Y=3.15 $X2=0 $Y2=0
cc_245 N_A_c_328_n N_VPWR_c_397_n 0.00583607f $X=3.785 $Y=3.15 $X2=0 $Y2=0
cc_246 N_A_c_328_n N_VPWR_c_390_n 0.0631216f $X=3.785 $Y=3.15 $X2=0 $Y2=0
cc_247 N_A_c_329_n N_VPWR_c_390_n 0.0127316f $X=1.98 $Y=3.15 $X2=0 $Y2=0
cc_248 N_A_c_321_n N_VGND_c_475_n 0.0187277f $X=1.99 $Y=1.22 $X2=0 $Y2=0
cc_249 N_A_c_324_n N_VGND_c_475_n 0.00232901f $X=1.8 $Y=1.385 $X2=0 $Y2=0
cc_250 A N_VGND_c_475_n 0.0288088f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_251 N_A_M1012_g N_VGND_c_476_n 0.0157197f $X=3.89 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A_c_321_n N_VGND_c_478_n 0.00348254f $X=1.99 $Y=1.22 $X2=0 $Y2=0
cc_253 N_A_M1012_g N_VGND_c_479_n 0.00383152f $X=3.89 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A_c_321_n N_VGND_c_480_n 0.00547229f $X=1.99 $Y=1.22 $X2=0 $Y2=0
cc_255 N_A_M1012_g N_VGND_c_480_n 0.0075725f $X=3.89 $Y=0.74 $X2=0 $Y2=0
cc_256 N_VPWR_c_392_n X 0.0455874f $X=0.3 $Y=1.985 $X2=0 $Y2=0
cc_257 N_VPWR_c_393_n X 0.0335865f $X=1.205 $Y=2.285 $X2=0 $Y2=0
cc_258 N_VPWR_c_395_n X 0.0157112f $X=1.085 $Y=3.33 $X2=0 $Y2=0
cc_259 N_VPWR_c_390_n X 0.0127977f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_260 N_X_c_438_n N_VGND_c_474_n 0.0308798f $X=0.73 $Y=0.515 $X2=0 $Y2=0
cc_261 N_X_c_438_n N_VGND_c_475_n 0.0245818f $X=0.73 $Y=0.515 $X2=0 $Y2=0
cc_262 N_X_c_438_n N_VGND_c_477_n 0.0149085f $X=0.73 $Y=0.515 $X2=0 $Y2=0
cc_263 N_X_c_438_n N_VGND_c_480_n 0.0122037f $X=0.73 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__dfxtp_4.spice
* Created: Wed Sep  2 12:04:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dfxtp_4.pex.spice"
.subckt sky130_fd_sc_ms__dfxtp_4  VNB VPB CLK D VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1028 N_VGND_M1028_d N_CLK_M1028_g N_A_27_74#_M1028_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.17575 AS=0.2109 PD=1.215 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1025 N_A_209_368#_M1025_d N_A_27_74#_M1025_g N_VGND_M1028_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2516 AS=0.17575 PD=2.16 PS=1.215 NRD=8.916 NRS=31.62 M=1 R=4.93333
+ SA=75000.8 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1022 N_A_440_503#_M1022_d N_D_M1022_g N_VGND_M1022_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.355025 PD=0.7 PS=2.6 NRD=0 NRS=225.792 M=1 R=2.8 SA=75000.5
+ SB=75003.1 A=0.063 P=1.14 MULT=1
MM1023 N_A_547_485#_M1023_d N_A_27_74#_M1023_g N_A_440_503#_M1022_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0756875 AS=0.0588 PD=0.83 PS=0.7 NRD=4.284 NRS=0 M=1 R=2.8
+ SA=75001 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1021 A_735_102# N_A_209_368#_M1021_g N_A_547_485#_M1023_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0756875 PD=0.63 PS=0.83 NRD=14.28 NRS=8.568 M=1 R=2.8
+ SA=75001.2 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_696_458#_M1016_g A_735_102# VNB NLOWVT L=0.15 W=0.42
+ AD=0.170728 AS=0.0441 PD=1.18206 PS=0.63 NRD=100.416 NRS=14.28 M=1 R=2.8
+ SA=75001.5 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1011 N_A_696_458#_M1011_d N_A_547_485#_M1011_g N_VGND_M1016_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.099 AS=0.223572 PD=0.985 PS=1.54794 NRD=0 NRS=76.68 M=1
+ R=3.66667 SA=75001.9 SB=75001.2 A=0.0825 P=1.4 MULT=1
MM1024 N_A_1037_424#_M1024_d N_A_209_368#_M1024_g N_A_696_458#_M1011_d VNB
+ NLOWVT L=0.15 W=0.55 AD=0.122021 AS=0.099 PD=1.11701 PS=0.985 NRD=24 NRS=0 M=1
+ R=3.66667 SA=75002.2 SB=75001 A=0.0825 P=1.4 MULT=1
MM1030 A_1178_124# N_A_27_74#_M1030_g N_A_1037_424#_M1024_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.06615 AS=0.0931794 PD=0.735 PS=0.85299 NRD=29.28 NRS=12.852 M=1
+ R=2.8 SA=75002.9 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_1226_296#_M1020_g A_1178_124# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.06615 PD=1.41 PS=0.735 NRD=0 NRS=29.28 M=1 R=2.8 SA=75003.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_A_1037_424#_M1026_g N_A_1226_296#_M1026_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1147 AS=0.2109 PD=1.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1026_d N_A_1226_296#_M1002_g N_Q_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1147 AS=0.1184 PD=1.05 PS=1.06 NRD=4.86 NRS=6.48 M=1 R=4.93333 SA=75000.7
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A_1226_296#_M1003_g N_Q_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.111 AS=0.1184 PD=1.04 PS=1.06 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1003_d N_A_1226_296#_M1008_g N_Q_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.111 AS=0.1036 PD=1.04 PS=1.02 NRD=3.24 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_A_1226_296#_M1017_g N_Q_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1012 N_VPWR_M1012_d N_CLK_M1012_g N_A_27_74#_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1013 N_A_209_368#_M1013_d N_A_27_74#_M1013_g N_VPWR_M1012_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1009 N_A_440_503#_M1009_d N_D_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=0.42
+ AD=0.082425 AS=0.2481 PD=0.865 PS=2.17 NRD=39.8531 NRS=251.274 M=1 R=2.33333
+ SA=90000.3 SB=90005.4 A=0.0756 P=1.2 MULT=1
MM1014 N_A_547_485#_M1014_d N_A_209_368#_M1014_g N_A_440_503#_M1009_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.082425 AS=0.082425 PD=0.865 PS=0.865 NRD=0 NRS=0 M=1
+ R=2.33333 SA=90000.7 SB=90005 A=0.0756 P=1.2 MULT=1
MM1005 A_654_503# N_A_27_74#_M1005_g N_A_547_485#_M1014_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0441 AS=0.082425 PD=0.63 PS=0.865 NRD=23.443 NRS=37.5088 M=1
+ R=2.33333 SA=90001.1 SB=90005.9 A=0.0756 P=1.2 MULT=1
MM1027 N_VPWR_M1027_d N_A_696_458#_M1027_g A_654_503# VPB PSHORT L=0.18 W=0.42
+ AD=0.1536 AS=0.0441 PD=1.13667 PS=0.63 NRD=145.721 NRS=23.443 M=1 R=2.33333
+ SA=90001.5 SB=90005.5 A=0.0756 P=1.2 MULT=1
MM1029 N_A_696_458#_M1029_d N_A_547_485#_M1029_g N_VPWR_M1027_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.21 AS=0.3072 PD=1.34 PS=2.27333 NRD=0 NRS=72.8506 M=1
+ R=4.66667 SA=90001.3 SB=90002.9 A=0.1512 P=2.04 MULT=1
MM1018 N_A_1037_424#_M1018_d N_A_27_74#_M1018_g N_A_696_458#_M1029_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.1778 AS=0.21 PD=1.59333 PS=1.34 NRD=0 NRS=52.7566 M=1
+ R=4.66667 SA=90002 SB=90002.2 A=0.1512 P=2.04 MULT=1
MM1006 A_1144_508# N_A_209_368#_M1006_g N_A_1037_424#_M1018_d VPB PSHORT L=0.18
+ W=0.42 AD=0.09345 AS=0.0889 PD=0.865 PS=0.796667 NRD=78.5636 NRS=73.481 M=1
+ R=2.33333 SA=90003.5 SB=90003.7 A=0.0756 P=1.2 MULT=1
MM1000 N_VPWR_M1000_d N_A_1226_296#_M1000_g A_1144_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.0805 AS=0.09345 PD=0.776667 PS=0.865 NRD=0 NRS=78.5636 M=1 R=2.33333
+ SA=90004.1 SB=90003 A=0.0756 P=1.2 MULT=1
MM1015 N_A_1226_296#_M1015_d N_A_1037_424#_M1015_g N_VPWR_M1000_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.1134 AS=0.161 PD=1.11 PS=1.55333 NRD=0 NRS=10.5395 M=1
+ R=4.66667 SA=90002.4 SB=90002.5 A=0.1512 P=2.04 MULT=1
MM1019 N_A_1226_296#_M1015_d N_A_1037_424#_M1019_g N_VPWR_M1019_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1134 AS=0.1614 PD=1.11 PS=1.26429 NRD=0 NRS=18.7544 M=1
+ R=4.66667 SA=90002.8 SB=90002.1 A=0.1512 P=2.04 MULT=1
MM1001 N_Q_M1001_d N_A_1226_296#_M1001_g N_VPWR_M1019_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2152 PD=1.39 PS=1.68571 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.6
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1004 N_Q_M1001_d N_A_1226_296#_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1007 N_Q_M1007_d N_A_1226_296#_M1007_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.5
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1010 N_Q_M1007_d N_A_1226_296#_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.9
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX31_noxref VNB VPB NWDIODE A=18.5628 P=23.68
c_217 VPB 0 1.17955e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__dfxtp_4.pxi.spice"
*
.ends
*
*

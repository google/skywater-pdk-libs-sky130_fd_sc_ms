* NGSPICE file created from sky130_fd_sc_ms__nand3_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__nand3_2 A B C VGND VNB VPB VPWR Y
M1000 a_27_74# C VGND VNB nlowvt w=740000u l=150000u
+  ad=6.068e+11p pd=6.08e+06u as=2.072e+11p ps=2.04e+06u
M1001 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=1.3384e+12p pd=1.135e+07u as=9.128e+11p ps=8.35e+06u
M1002 a_283_74# A Y VNB nlowvt w=740000u l=150000u
+  ad=7.123e+11p pd=5.5e+06u as=2.072e+11p ps=2.04e+06u
M1003 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y C VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR C Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_283_74# B a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_74# B a_283_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND C a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A a_283_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


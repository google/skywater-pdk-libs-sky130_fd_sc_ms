* NGSPICE file created from sky130_fd_sc_ms__edfxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__edfxbp_1 CLK D DE VGND VNB VPB VPWR Q Q_N
M1000 a_1198_97# a_1008_74# a_27_74# VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=4.349e+11p ps=4.69e+06u
M1001 a_527_74# a_161_446# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.908e+12p ps=1.641e+07u
M1002 a_27_74# a_575_48# a_527_74# VNB nlowvt w=420000u l=150000u
+  ad=4.158e+11p pd=4.5e+06u as=0p ps=0u
M1003 a_2209_443# a_1008_74# a_1879_74# VPB pshort w=420000u l=180000u
+  ad=1.26e+11p pd=1.44e+06u as=3.262e+11p ps=2.78e+06u
M1004 a_1807_74# a_1419_71# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.554e+11p pd=1.9e+06u as=0p ps=0u
M1005 a_1419_71# a_1198_97# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=2.42065e+12p ps=2.12e+07u
M1006 a_1879_74# a_1008_74# a_1807_74# VNB nlowvt w=740000u l=150000u
+  ad=7.478e+11p pd=4.66e+06u as=0p ps=0u
M1007 a_1426_508# a_818_74# a_1198_97# VPB pshort w=420000u l=180000u
+  ad=1.386e+11p pd=1.5e+06u as=0p ps=0u
M1008 VPWR DE a_161_446# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1009 a_559_504# DE VPWR VPB pshort w=420000u l=180000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1010 VGND a_575_48# a_2227_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1011 VPWR a_161_446# a_119_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1012 a_2011_392# a_1419_71# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1013 a_575_48# a_1879_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1014 a_1334_97# a_1008_74# a_1198_97# VNB nlowvt w=420000u l=150000u
+  ad=1.785e+11p pd=1.69e+06u as=2.226e+11p ps=1.9e+06u
M1015 a_1419_71# a_1198_97# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1016 a_575_48# a_1879_74# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1017 VGND a_1879_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1018 VGND DE a_145_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1019 VGND a_1419_71# a_1334_97# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Q_N a_575_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1021 a_2227_118# a_818_74# a_1879_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_575_48# a_2209_443# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR a_1419_71# a_1426_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND DE a_161_446# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.281e+11p ps=1.45e+06u
M1025 a_818_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1026 VPWR a_1879_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1027 a_119_508# D a_27_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1008_74# a_818_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1029 a_1008_74# a_818_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1030 Q_N a_575_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1031 a_818_74# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1032 a_145_74# D a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_27_74# a_575_48# a_559_504# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1198_97# a_818_74# a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1879_74# a_818_74# a_2011_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__o32a_2.pxi.spice
* Created: Wed Sep  2 12:26:16 2020
* 
x_PM_SKY130_FD_SC_MS__O32A_2%A_83_264# N_A_83_264#_M1001_d N_A_83_264#_M1006_d
+ N_A_83_264#_M1004_g N_A_83_264#_M1010_g N_A_83_264#_M1005_g
+ N_A_83_264#_M1013_g N_A_83_264#_c_87_n N_A_83_264#_c_102_p N_A_83_264#_c_146_p
+ N_A_83_264#_c_94_n N_A_83_264#_c_95_n N_A_83_264#_c_139_p N_A_83_264#_c_88_n
+ N_A_83_264#_c_89_n N_A_83_264#_c_90_n N_A_83_264#_c_118_p N_A_83_264#_c_122_p
+ PM_SKY130_FD_SC_MS__O32A_2%A_83_264#
x_PM_SKY130_FD_SC_MS__O32A_2%A1 N_A1_M1012_g N_A1_M1007_g A1 N_A1_c_197_n
+ N_A1_c_198_n N_A1_c_201_n PM_SKY130_FD_SC_MS__O32A_2%A1
x_PM_SKY130_FD_SC_MS__O32A_2%A2 N_A2_M1000_g N_A2_M1011_g A2 N_A2_c_236_n
+ N_A2_c_237_n PM_SKY130_FD_SC_MS__O32A_2%A2
x_PM_SKY130_FD_SC_MS__O32A_2%A3 N_A3_M1006_g N_A3_M1002_g A3 N_A3_c_273_n
+ N_A3_c_274_n PM_SKY130_FD_SC_MS__O32A_2%A3
x_PM_SKY130_FD_SC_MS__O32A_2%B2 N_B2_M1001_g N_B2_M1003_g B2 N_B2_c_311_n
+ PM_SKY130_FD_SC_MS__O32A_2%B2
x_PM_SKY130_FD_SC_MS__O32A_2%B1 N_B1_M1008_g N_B1_c_346_n N_B1_c_347_n
+ N_B1_c_348_n N_B1_M1009_g N_B1_c_349_n B1 B1 B1 B1 B1 N_B1_c_351_n
+ PM_SKY130_FD_SC_MS__O32A_2%B1
x_PM_SKY130_FD_SC_MS__O32A_2%VPWR N_VPWR_M1004_s N_VPWR_M1005_s N_VPWR_M1008_d
+ N_VPWR_c_382_n N_VPWR_c_383_n N_VPWR_c_384_n N_VPWR_c_385_n N_VPWR_c_386_n
+ N_VPWR_c_387_n VPWR N_VPWR_c_388_n N_VPWR_c_389_n N_VPWR_c_381_n
+ N_VPWR_c_391_n PM_SKY130_FD_SC_MS__O32A_2%VPWR
x_PM_SKY130_FD_SC_MS__O32A_2%X N_X_M1010_d N_X_M1004_d N_X_c_431_n N_X_c_432_n X
+ X X X N_X_c_433_n PM_SKY130_FD_SC_MS__O32A_2%X
x_PM_SKY130_FD_SC_MS__O32A_2%VGND N_VGND_M1010_s N_VGND_M1013_s N_VGND_M1011_d
+ N_VGND_c_473_n N_VGND_c_474_n N_VGND_c_475_n N_VGND_c_476_n N_VGND_c_477_n
+ N_VGND_c_478_n N_VGND_c_479_n N_VGND_c_480_n N_VGND_c_481_n N_VGND_c_482_n
+ VGND N_VGND_c_483_n N_VGND_c_484_n PM_SKY130_FD_SC_MS__O32A_2%VGND
x_PM_SKY130_FD_SC_MS__O32A_2%A_349_74# N_A_349_74#_M1007_d N_A_349_74#_M1002_d
+ N_A_349_74#_M1009_d N_A_349_74#_c_533_n N_A_349_74#_c_534_n
+ N_A_349_74#_c_535_n N_A_349_74#_c_536_n N_A_349_74#_c_553_n
+ N_A_349_74#_c_537_n N_A_349_74#_c_538_n PM_SKY130_FD_SC_MS__O32A_2%A_349_74#
cc_1 VNB N_A_83_264#_M1004_g 0.0150953f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A_83_264#_M1010_g 0.0249445f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.74
cc_3 VNB N_A_83_264#_M1005_g 5.20588e-19 $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_4 VNB N_A_83_264#_M1013_g 0.0241735f $X=-0.19 $Y=-0.245 $X2=1.1 $Y2=0.74
cc_5 VNB N_A_83_264#_c_87_n 2.18704e-19 $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.95
cc_6 VNB N_A_83_264#_c_88_n 0.0105334f $X=-0.19 $Y=-0.245 $X2=4.1 $Y2=1.95
cc_7 VNB N_A_83_264#_c_89_n 0.0516301f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.485
cc_8 VNB N_A_83_264#_c_90_n 0.00302828f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.485
cc_9 VNB N_A1_M1007_g 0.0261215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A1_c_197_n 0.0247502f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.32
cc_11 VNB N_A1_c_198_n 0.00555649f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.74
cc_12 VNB N_A2_M1011_g 0.0257807f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.47
cc_13 VNB N_A2_c_236_n 0.0266114f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.74
cc_14 VNB N_A2_c_237_n 0.00165774f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.74
cc_15 VNB N_A3_M1002_g 0.0267316f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.47
cc_16 VNB N_A3_c_273_n 0.0266032f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.74
cc_17 VNB N_A3_c_274_n 0.00165645f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.74
cc_18 VNB N_B2_M1001_g 0.0357125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB B2 0.00601402f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_20 VNB N_B2_c_311_n 0.0236905f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.74
cc_21 VNB N_B1_M1008_g 0.00582472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B1_c_346_n 0.0218972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B1_c_347_n 0.00989991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B1_c_348_n 0.0274572f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.47
cc_25 VNB N_B1_c_349_n 0.0180432f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.32
cc_26 VNB B1 0.0118942f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.74
cc_27 VNB N_B1_c_351_n 0.0543697f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.65
cc_28 VNB N_VPWR_c_381_n 0.203486f $X=-0.19 $Y=-0.245 $X2=2.892 $Y2=2.035
cc_29 VNB N_X_c_431_n 0.00500933f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_30 VNB N_X_c_432_n 0.00239713f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.32
cc_31 VNB N_X_c_433_n 0.00759022f $X=-0.19 $Y=-0.245 $X2=4.1 $Y2=1.045
cc_32 VNB N_VGND_c_473_n 0.0140441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_474_n 0.0226334f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.74
cc_34 VNB N_VGND_c_475_n 0.0175838f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_35 VNB N_VGND_c_476_n 0.0178579f $X=-0.19 $Y=-0.245 $X2=1.1 $Y2=0.74
cc_36 VNB N_VGND_c_477_n 0.00899389f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.95
cc_37 VNB N_VGND_c_478_n 0.00829839f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=2.035
cc_38 VNB N_VGND_c_479_n 0.019013f $X=-0.19 $Y=-0.245 $X2=2.892 $Y2=2.715
cc_39 VNB N_VGND_c_480_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.9 $Y2=2.715
cc_40 VNB N_VGND_c_481_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=4.015 $Y2=2.035
cc_41 VNB N_VGND_c_482_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=3.11 $Y2=2.035
cc_42 VNB N_VGND_c_483_n 0.0589592f $X=-0.19 $Y=-0.245 $X2=4.02 $Y2=0.88
cc_43 VNB N_VGND_c_484_n 0.27806f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.47
cc_44 VNB N_A_349_74#_c_533_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.74
cc_45 VNB N_A_349_74#_c_534_n 0.0183106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_349_74#_c_535_n 0.00851793f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.65
cc_47 VNB N_A_349_74#_c_536_n 0.00261637f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_48 VNB N_A_349_74#_c_537_n 0.00879016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_349_74#_c_538_n 0.00311899f $X=-0.19 $Y=-0.245 $X2=2.675 $Y2=2.035
cc_50 VPB N_A_83_264#_M1004_g 0.0274013f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_51 VPB N_A_83_264#_M1005_g 0.0243899f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_52 VPB N_A_83_264#_c_87_n 0.00278836f $X=-0.19 $Y=1.66 $X2=1.15 $Y2=1.95
cc_53 VPB N_A_83_264#_c_94_n 0.00399457f $X=-0.19 $Y=1.66 $X2=2.9 $Y2=2.715
cc_54 VPB N_A_83_264#_c_95_n 0.00378081f $X=-0.19 $Y=1.66 $X2=4.015 $Y2=2.035
cc_55 VPB N_A_83_264#_c_88_n 0.00500212f $X=-0.19 $Y=1.66 $X2=4.1 $Y2=1.95
cc_56 VPB N_A1_c_197_n 0.00874992f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.32
cc_57 VPB N_A1_c_198_n 0.00298783f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=0.74
cc_58 VPB N_A1_c_201_n 0.0190646f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A2_M1000_g 0.0214855f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A2_c_236_n 0.00564792f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=0.74
cc_61 VPB N_A2_c_237_n 0.00205011f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=0.74
cc_62 VPB N_A3_M1006_g 0.0227919f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A3_c_273_n 0.00564713f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=0.74
cc_64 VPB N_A3_c_274_n 0.00208094f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=0.74
cc_65 VPB N_B2_M1003_g 0.0225579f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.47
cc_66 VPB B2 0.00454059f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_67 VPB N_B2_c_311_n 0.00545272f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=0.74
cc_68 VPB N_B1_M1008_g 0.0251101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB B1 0.0735816f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=0.74
cc_70 VPB N_VPWR_c_382_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_383_n 0.0587144f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=0.74
cc_72 VPB N_VPWR_c_384_n 0.0142926f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_385_n 0.0247234f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_386_n 0.0676428f $X=-0.19 $Y=1.66 $X2=2.675 $Y2=2.035
cc_75 VPB N_VPWR_c_387_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.235 $Y2=2.035
cc_76 VPB N_VPWR_c_388_n 0.0194151f $X=-0.19 $Y=1.66 $X2=2.9 $Y2=2.715
cc_77 VPB N_VPWR_c_389_n 0.0208395f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_381_n 0.120852f $X=-0.19 $Y=1.66 $X2=2.892 $Y2=2.035
cc_79 VPB N_VPWR_c_391_n 0.0102647f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.47
cc_80 VPB X 0.00459114f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_81 VPB X 0.00231613f $X=-0.19 $Y=1.66 $X2=1.235 $Y2=2.035
cc_82 VPB N_X_c_433_n 0.00123129f $X=-0.19 $Y=1.66 $X2=4.1 $Y2=1.045
cc_83 N_A_83_264#_M1013_g N_A1_M1007_g 0.0233513f $X=1.1 $Y=0.74 $X2=0 $Y2=0
cc_84 N_A_83_264#_c_89_n N_A1_M1007_g 8.1421e-19 $X=1.04 $Y=1.485 $X2=0 $Y2=0
cc_85 N_A_83_264#_c_90_n N_A1_M1007_g 5.77738e-19 $X=1.15 $Y=1.485 $X2=0 $Y2=0
cc_86 N_A_83_264#_M1005_g N_A1_c_197_n 0.00189768f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_87 N_A_83_264#_c_87_n N_A1_c_197_n 5.4577e-19 $X=1.15 $Y=1.95 $X2=0 $Y2=0
cc_88 N_A_83_264#_c_102_p N_A1_c_197_n 7.901e-19 $X=2.675 $Y=2.035 $X2=0 $Y2=0
cc_89 N_A_83_264#_c_89_n N_A1_c_197_n 0.0188248f $X=1.04 $Y=1.485 $X2=0 $Y2=0
cc_90 N_A_83_264#_c_90_n N_A1_c_197_n 0.00170854f $X=1.15 $Y=1.485 $X2=0 $Y2=0
cc_91 N_A_83_264#_c_87_n N_A1_c_198_n 0.00969328f $X=1.15 $Y=1.95 $X2=0 $Y2=0
cc_92 N_A_83_264#_c_102_p N_A1_c_198_n 0.0251787f $X=2.675 $Y=2.035 $X2=0 $Y2=0
cc_93 N_A_83_264#_c_89_n N_A1_c_198_n 3.50433e-19 $X=1.04 $Y=1.485 $X2=0 $Y2=0
cc_94 N_A_83_264#_c_90_n N_A1_c_198_n 0.0231673f $X=1.15 $Y=1.485 $X2=0 $Y2=0
cc_95 N_A_83_264#_M1005_g N_A1_c_201_n 0.0148269f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_96 N_A_83_264#_c_87_n N_A1_c_201_n 0.0033687f $X=1.15 $Y=1.95 $X2=0 $Y2=0
cc_97 N_A_83_264#_c_102_p N_A1_c_201_n 0.0168407f $X=2.675 $Y=2.035 $X2=0 $Y2=0
cc_98 N_A_83_264#_c_102_p N_A2_M1000_g 0.0173173f $X=2.675 $Y=2.035 $X2=0 $Y2=0
cc_99 N_A_83_264#_c_94_n N_A2_M1000_g 0.00348338f $X=2.9 $Y=2.715 $X2=0 $Y2=0
cc_100 N_A_83_264#_c_102_p N_A2_c_236_n 7.07929e-19 $X=2.675 $Y=2.035 $X2=0
+ $Y2=0
cc_101 N_A_83_264#_c_102_p N_A2_c_237_n 0.0229716f $X=2.675 $Y=2.035 $X2=0 $Y2=0
cc_102 N_A_83_264#_c_102_p N_A3_M1006_g 0.0133177f $X=2.675 $Y=2.035 $X2=0 $Y2=0
cc_103 N_A_83_264#_c_94_n N_A3_M1006_g 0.0168861f $X=2.9 $Y=2.715 $X2=0 $Y2=0
cc_104 N_A_83_264#_c_118_p N_A3_M1006_g 8.8334e-19 $X=2.9 $Y=2.035 $X2=0 $Y2=0
cc_105 N_A_83_264#_c_118_p N_A3_c_273_n 7.71396e-19 $X=2.9 $Y=2.035 $X2=0 $Y2=0
cc_106 N_A_83_264#_c_102_p N_A3_c_274_n 0.0108932f $X=2.675 $Y=2.035 $X2=0 $Y2=0
cc_107 N_A_83_264#_c_118_p N_A3_c_274_n 0.0130747f $X=2.9 $Y=2.035 $X2=0 $Y2=0
cc_108 N_A_83_264#_c_122_p N_B2_M1001_g 0.00419034f $X=4.02 $Y=0.88 $X2=0 $Y2=0
cc_109 N_A_83_264#_c_94_n N_B2_M1003_g 0.0162401f $X=2.9 $Y=2.715 $X2=0 $Y2=0
cc_110 N_A_83_264#_c_95_n N_B2_M1003_g 0.0146269f $X=4.015 $Y=2.035 $X2=0 $Y2=0
cc_111 N_A_83_264#_c_118_p N_B2_M1003_g 4.27055e-19 $X=2.9 $Y=2.035 $X2=0 $Y2=0
cc_112 N_A_83_264#_c_95_n B2 0.042577f $X=4.015 $Y=2.035 $X2=0 $Y2=0
cc_113 N_A_83_264#_c_88_n B2 0.0217679f $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_114 N_A_83_264#_c_118_p B2 0.00117862f $X=2.9 $Y=2.035 $X2=0 $Y2=0
cc_115 N_A_83_264#_c_122_p B2 0.0247412f $X=4.02 $Y=0.88 $X2=0 $Y2=0
cc_116 N_A_83_264#_c_95_n N_B2_c_311_n 7.14995e-19 $X=4.015 $Y=2.035 $X2=0 $Y2=0
cc_117 N_A_83_264#_c_88_n N_B2_c_311_n 2.63846e-19 $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_118 N_A_83_264#_c_122_p N_B2_c_311_n 0.00366748f $X=4.02 $Y=0.88 $X2=0 $Y2=0
cc_119 N_A_83_264#_c_94_n N_B1_M1008_g 0.00335433f $X=2.9 $Y=2.715 $X2=0 $Y2=0
cc_120 N_A_83_264#_c_95_n N_B1_M1008_g 0.0220977f $X=4.015 $Y=2.035 $X2=0 $Y2=0
cc_121 N_A_83_264#_c_88_n N_B1_M1008_g 0.010813f $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_122 N_A_83_264#_c_95_n N_B1_c_346_n 0.00376079f $X=4.015 $Y=2.035 $X2=0 $Y2=0
cc_123 N_A_83_264#_c_88_n N_B1_c_346_n 0.0113712f $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_124 N_A_83_264#_c_122_p N_B1_c_347_n 0.0101883f $X=4.02 $Y=0.88 $X2=0 $Y2=0
cc_125 N_A_83_264#_c_139_p N_B1_c_348_n 0.00517368f $X=4.1 $Y=1.045 $X2=0 $Y2=0
cc_126 N_A_83_264#_c_88_n N_B1_c_348_n 0.00830667f $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_127 N_A_83_264#_c_88_n N_B1_c_349_n 0.00891863f $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_128 N_A_83_264#_c_95_n B1 0.0150384f $X=4.015 $Y=2.035 $X2=0 $Y2=0
cc_129 N_A_83_264#_c_88_n B1 0.0582284f $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_130 N_A_83_264#_c_87_n N_VPWR_M1005_s 0.00223621f $X=1.15 $Y=1.95 $X2=0 $Y2=0
cc_131 N_A_83_264#_c_102_p N_VPWR_M1005_s 0.0119287f $X=2.675 $Y=2.035 $X2=0
+ $Y2=0
cc_132 N_A_83_264#_c_146_p N_VPWR_M1005_s 0.00269585f $X=1.235 $Y=2.035 $X2=0
+ $Y2=0
cc_133 N_A_83_264#_c_95_n N_VPWR_M1008_d 0.00491466f $X=4.015 $Y=2.035 $X2=0
+ $Y2=0
cc_134 N_A_83_264#_c_88_n N_VPWR_M1008_d 0.00186754f $X=4.1 $Y=1.95 $X2=0 $Y2=0
cc_135 N_A_83_264#_M1004_g N_VPWR_c_383_n 0.00647357f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_136 N_A_83_264#_M1005_g N_VPWR_c_384_n 0.00773607f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_137 N_A_83_264#_c_102_p N_VPWR_c_384_n 0.0247222f $X=2.675 $Y=2.035 $X2=0
+ $Y2=0
cc_138 N_A_83_264#_c_146_p N_VPWR_c_384_n 0.0116292f $X=1.235 $Y=2.035 $X2=0
+ $Y2=0
cc_139 N_A_83_264#_c_89_n N_VPWR_c_384_n 3.82399e-19 $X=1.04 $Y=1.485 $X2=0
+ $Y2=0
cc_140 N_A_83_264#_c_95_n N_VPWR_c_385_n 0.022977f $X=4.015 $Y=2.035 $X2=0 $Y2=0
cc_141 N_A_83_264#_c_94_n N_VPWR_c_386_n 0.0136324f $X=2.9 $Y=2.715 $X2=0 $Y2=0
cc_142 N_A_83_264#_M1004_g N_VPWR_c_388_n 0.0048691f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_143 N_A_83_264#_M1005_g N_VPWR_c_388_n 0.005209f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A_83_264#_M1004_g N_VPWR_c_381_n 0.00875947f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_145 N_A_83_264#_M1005_g N_VPWR_c_381_n 0.00986727f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_146 N_A_83_264#_c_94_n N_VPWR_c_381_n 0.0149529f $X=2.9 $Y=2.715 $X2=0 $Y2=0
cc_147 N_A_83_264#_M1010_g N_X_c_431_n 0.0127873f $X=0.67 $Y=0.74 $X2=0 $Y2=0
cc_148 N_A_83_264#_M1013_g N_X_c_431_n 0.002387f $X=1.1 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A_83_264#_c_89_n N_X_c_431_n 0.00344849f $X=1.04 $Y=1.485 $X2=0 $Y2=0
cc_150 N_A_83_264#_c_90_n N_X_c_431_n 0.0120032f $X=1.15 $Y=1.485 $X2=0 $Y2=0
cc_151 N_A_83_264#_M1010_g N_X_c_432_n 0.00875007f $X=0.67 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A_83_264#_M1013_g N_X_c_432_n 0.00755147f $X=1.1 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A_83_264#_M1004_g X 0.00270934f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_154 N_A_83_264#_M1005_g X 0.00304813f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_155 N_A_83_264#_c_87_n X 0.00565814f $X=1.15 $Y=1.95 $X2=0 $Y2=0
cc_156 N_A_83_264#_c_89_n X 0.00279675f $X=1.04 $Y=1.485 $X2=0 $Y2=0
cc_157 N_A_83_264#_c_90_n X 0.00151667f $X=1.15 $Y=1.485 $X2=0 $Y2=0
cc_158 N_A_83_264#_M1004_g X 0.0149161f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_159 N_A_83_264#_M1005_g X 0.0143207f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_160 N_A_83_264#_M1004_g N_X_c_433_n 0.0172943f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_161 N_A_83_264#_M1010_g N_X_c_433_n 0.00770058f $X=0.67 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A_83_264#_M1013_g N_X_c_433_n 0.00109865f $X=1.1 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A_83_264#_c_87_n N_X_c_433_n 0.00756879f $X=1.15 $Y=1.95 $X2=0 $Y2=0
cc_164 N_A_83_264#_c_89_n N_X_c_433_n 0.0141153f $X=1.04 $Y=1.485 $X2=0 $Y2=0
cc_165 N_A_83_264#_c_90_n N_X_c_433_n 0.0243803f $X=1.15 $Y=1.485 $X2=0 $Y2=0
cc_166 N_A_83_264#_c_102_p A_349_368# 0.0096152f $X=2.675 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_167 N_A_83_264#_c_102_p A_433_368# 0.01606f $X=2.675 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_168 N_A_83_264#_c_95_n A_655_368# 0.0135682f $X=4.015 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_169 N_A_83_264#_M1010_g N_VGND_c_474_n 0.00671933f $X=0.67 $Y=0.74 $X2=0
+ $Y2=0
cc_170 N_A_83_264#_M1010_g N_VGND_c_475_n 0.00453882f $X=0.67 $Y=0.74 $X2=0
+ $Y2=0
cc_171 N_A_83_264#_M1013_g N_VGND_c_476_n 0.00806966f $X=1.1 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A_83_264#_c_90_n N_VGND_c_476_n 0.00114473f $X=1.15 $Y=1.485 $X2=0
+ $Y2=0
cc_173 N_A_83_264#_c_89_n N_VGND_c_478_n 0.00401809f $X=1.04 $Y=1.485 $X2=0
+ $Y2=0
cc_174 N_A_83_264#_M1010_g N_VGND_c_479_n 0.00434272f $X=0.67 $Y=0.74 $X2=0
+ $Y2=0
cc_175 N_A_83_264#_M1013_g N_VGND_c_479_n 0.00434272f $X=1.1 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A_83_264#_M1010_g N_VGND_c_484_n 0.00824408f $X=0.67 $Y=0.74 $X2=0
+ $Y2=0
cc_177 N_A_83_264#_M1013_g N_VGND_c_484_n 0.00821312f $X=1.1 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A_83_264#_M1013_g N_A_349_74#_c_535_n 2.49809e-19 $X=1.1 $Y=0.74 $X2=0
+ $Y2=0
cc_179 N_A_83_264#_M1001_d N_A_349_74#_c_537_n 0.0136122f $X=3.245 $Y=0.37 $X2=0
+ $Y2=0
cc_180 N_A_83_264#_c_139_p N_A_349_74#_c_537_n 0.0076481f $X=4.1 $Y=1.045 $X2=0
+ $Y2=0
cc_181 N_A_83_264#_c_122_p N_A_349_74#_c_537_n 0.0478533f $X=4.02 $Y=0.88 $X2=0
+ $Y2=0
cc_182 N_A1_c_201_n N_A2_M1000_g 0.0448317f $X=1.58 $Y=1.725 $X2=0 $Y2=0
cc_183 N_A1_M1007_g N_A2_M1011_g 0.019972f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_184 N_A1_c_197_n N_A2_c_236_n 0.0448317f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_185 N_A1_c_198_n N_A2_c_236_n 0.00260109f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_186 N_A1_c_197_n N_A2_c_237_n 4.97174e-19 $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_187 N_A1_c_198_n N_A2_c_237_n 0.0316293f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_188 N_A1_c_201_n N_VPWR_c_384_n 0.0215558f $X=1.58 $Y=1.725 $X2=0 $Y2=0
cc_189 N_A1_c_201_n N_VPWR_c_386_n 0.00476448f $X=1.58 $Y=1.725 $X2=0 $Y2=0
cc_190 N_A1_c_201_n N_VPWR_c_381_n 0.00494823f $X=1.58 $Y=1.725 $X2=0 $Y2=0
cc_191 N_A1_c_201_n X 7.38946e-19 $X=1.58 $Y=1.725 $X2=0 $Y2=0
cc_192 N_A1_M1007_g N_VGND_c_476_n 0.00666787f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_193 N_A1_c_197_n N_VGND_c_476_n 0.00101787f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_194 N_A1_c_198_n N_VGND_c_476_n 0.00945165f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_195 N_A1_M1007_g N_VGND_c_481_n 0.00434272f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A1_M1007_g N_VGND_c_484_n 0.0082141f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A1_M1007_g N_A_349_74#_c_533_n 0.00795429f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_198 N_A1_M1007_g N_A_349_74#_c_535_n 0.00350994f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A1_c_198_n N_A_349_74#_c_535_n 0.00648331f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_200 N_A2_M1000_g N_A3_M1006_g 0.0469345f $X=2.075 $Y=2.34 $X2=0 $Y2=0
cc_201 N_A2_c_237_n N_A3_M1006_g 6.85212e-19 $X=2.15 $Y=1.515 $X2=0 $Y2=0
cc_202 N_A2_M1011_g N_A3_M1002_g 0.0260254f $X=2.1 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A2_c_236_n N_A3_c_273_n 0.0201104f $X=2.15 $Y=1.515 $X2=0 $Y2=0
cc_204 N_A2_c_237_n N_A3_c_273_n 0.00114936f $X=2.15 $Y=1.515 $X2=0 $Y2=0
cc_205 N_A2_c_236_n N_A3_c_274_n 0.00114936f $X=2.15 $Y=1.515 $X2=0 $Y2=0
cc_206 N_A2_c_237_n N_A3_c_274_n 0.0276388f $X=2.15 $Y=1.515 $X2=0 $Y2=0
cc_207 N_A2_M1000_g N_VPWR_c_384_n 0.0032754f $X=2.075 $Y=2.34 $X2=0 $Y2=0
cc_208 N_A2_M1000_g N_VPWR_c_386_n 0.0059286f $X=2.075 $Y=2.34 $X2=0 $Y2=0
cc_209 N_A2_M1000_g N_VPWR_c_381_n 0.00610055f $X=2.075 $Y=2.34 $X2=0 $Y2=0
cc_210 N_A2_M1011_g N_VGND_c_477_n 0.00484409f $X=2.1 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A2_M1011_g N_VGND_c_481_n 0.00434272f $X=2.1 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A2_M1011_g N_VGND_c_484_n 0.0082141f $X=2.1 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A2_M1011_g N_A_349_74#_c_533_n 0.00966073f $X=2.1 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A2_M1011_g N_A_349_74#_c_534_n 0.0117933f $X=2.1 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A2_c_236_n N_A_349_74#_c_534_n 9.79877e-19 $X=2.15 $Y=1.515 $X2=0 $Y2=0
cc_216 N_A2_c_237_n N_A_349_74#_c_534_n 0.019847f $X=2.15 $Y=1.515 $X2=0 $Y2=0
cc_217 N_A2_M1011_g N_A_349_74#_c_535_n 0.0015571f $X=2.1 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A2_c_236_n N_A_349_74#_c_535_n 3.0499e-19 $X=2.15 $Y=1.515 $X2=0 $Y2=0
cc_219 N_A2_c_237_n N_A_349_74#_c_535_n 0.00541082f $X=2.15 $Y=1.515 $X2=0 $Y2=0
cc_220 N_A2_M1011_g N_A_349_74#_c_553_n 5.94859e-19 $X=2.1 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A3_M1002_g N_B2_M1001_g 0.0247403f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A3_M1006_g N_B2_M1003_g 0.00980851f $X=2.615 $Y=2.34 $X2=0 $Y2=0
cc_223 N_A3_c_274_n N_B2_M1003_g 3.99374e-19 $X=2.69 $Y=1.515 $X2=0 $Y2=0
cc_224 N_A3_c_273_n B2 0.00120971f $X=2.69 $Y=1.515 $X2=0 $Y2=0
cc_225 N_A3_c_274_n B2 0.0260963f $X=2.69 $Y=1.515 $X2=0 $Y2=0
cc_226 N_A3_c_273_n N_B2_c_311_n 0.017626f $X=2.69 $Y=1.515 $X2=0 $Y2=0
cc_227 N_A3_c_274_n N_B2_c_311_n 4.20763e-19 $X=2.69 $Y=1.515 $X2=0 $Y2=0
cc_228 N_A3_M1006_g N_VPWR_c_386_n 0.0056753f $X=2.615 $Y=2.34 $X2=0 $Y2=0
cc_229 N_A3_M1006_g N_VPWR_c_381_n 0.00610055f $X=2.615 $Y=2.34 $X2=0 $Y2=0
cc_230 N_A3_M1002_g N_VGND_c_477_n 0.00622568f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A3_M1002_g N_VGND_c_483_n 0.00433139f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A3_M1002_g N_VGND_c_484_n 0.00818355f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A3_M1002_g N_A_349_74#_c_533_n 6.28869e-19 $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A3_M1002_g N_A_349_74#_c_534_n 0.0133747f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A3_c_273_n N_A_349_74#_c_534_n 0.00134262f $X=2.69 $Y=1.515 $X2=0 $Y2=0
cc_236 N_A3_c_274_n N_A_349_74#_c_534_n 0.0259036f $X=2.69 $Y=1.515 $X2=0 $Y2=0
cc_237 N_A3_M1002_g N_A_349_74#_c_536_n 0.00227367f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A3_M1002_g N_A_349_74#_c_553_n 0.00745726f $X=2.67 $Y=0.74 $X2=0 $Y2=0
cc_239 N_B2_M1003_g N_B1_M1008_g 0.0399904f $X=3.185 $Y=2.34 $X2=0 $Y2=0
cc_240 B2 N_B1_M1008_g 0.0073182f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_241 B2 N_B1_c_347_n 0.00597337f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_242 N_B2_c_311_n N_B1_c_347_n 0.0153847f $X=3.26 $Y=1.515 $X2=0 $Y2=0
cc_243 B2 N_B1_c_349_n 2.68126e-19 $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_244 N_B2_M1003_g N_VPWR_c_385_n 0.00308866f $X=3.185 $Y=2.34 $X2=0 $Y2=0
cc_245 N_B2_M1003_g N_VPWR_c_386_n 0.00580632f $X=3.185 $Y=2.34 $X2=0 $Y2=0
cc_246 N_B2_M1003_g N_VPWR_c_381_n 0.00610055f $X=3.185 $Y=2.34 $X2=0 $Y2=0
cc_247 N_B2_M1001_g N_VGND_c_483_n 0.00291649f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_248 N_B2_M1001_g N_VGND_c_484_n 0.00364831f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_249 N_B2_M1001_g N_A_349_74#_c_534_n 0.0028014f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_250 N_B2_M1001_g N_A_349_74#_c_537_n 0.0161408f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_251 N_B1_M1008_g N_VPWR_c_385_n 0.0178572f $X=3.755 $Y=2.34 $X2=0 $Y2=0
cc_252 B1 N_VPWR_c_385_n 0.0430854f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_253 N_B1_M1008_g N_VPWR_c_386_n 0.00492916f $X=3.755 $Y=2.34 $X2=0 $Y2=0
cc_254 B1 N_VPWR_c_389_n 0.0107254f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_255 N_B1_M1008_g N_VPWR_c_381_n 0.00511769f $X=3.755 $Y=2.34 $X2=0 $Y2=0
cc_256 B1 N_VPWR_c_381_n 0.0114362f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_257 N_B1_c_348_n N_VGND_c_483_n 0.00291649f $X=4.235 $Y=1.22 $X2=0 $Y2=0
cc_258 N_B1_c_348_n N_VGND_c_484_n 0.00367994f $X=4.235 $Y=1.22 $X2=0 $Y2=0
cc_259 N_B1_c_348_n N_A_349_74#_c_537_n 0.0141061f $X=4.235 $Y=1.22 $X2=0 $Y2=0
cc_260 B1 N_A_349_74#_c_538_n 0.0231725f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_261 N_B1_c_351_n N_A_349_74#_c_538_n 0.00178757f $X=4.52 $Y=1.385 $X2=0 $Y2=0
cc_262 N_VPWR_c_383_n X 0.0455874f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_263 N_VPWR_c_384_n X 0.0270879f $X=1.425 $Y=2.385 $X2=0 $Y2=0
cc_264 N_VPWR_c_388_n X 0.0157112f $X=1.065 $Y=3.33 $X2=0 $Y2=0
cc_265 N_VPWR_c_381_n X 0.0127977f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_266 N_VPWR_c_383_n N_VGND_c_475_n 0.00876255f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_267 N_X_c_431_n N_VGND_M1010_s 0.00163897f $X=0.885 $Y=0.96 $X2=-0.19
+ $Y2=-0.245
cc_268 N_X_c_432_n N_VGND_c_474_n 0.016559f $X=0.885 $Y=0.515 $X2=0 $Y2=0
cc_269 N_X_c_431_n N_VGND_c_475_n 0.013787f $X=0.885 $Y=0.96 $X2=0 $Y2=0
cc_270 N_X_c_432_n N_VGND_c_475_n 0.0073154f $X=0.885 $Y=0.515 $X2=0 $Y2=0
cc_271 N_X_c_433_n N_VGND_c_475_n 7.75603e-19 $X=0.715 $Y=1.82 $X2=0 $Y2=0
cc_272 N_X_c_431_n N_VGND_c_476_n 0.00753583f $X=0.885 $Y=0.96 $X2=0 $Y2=0
cc_273 N_X_c_432_n N_VGND_c_476_n 0.0236791f $X=0.885 $Y=0.515 $X2=0 $Y2=0
cc_274 N_X_c_432_n N_VGND_c_479_n 0.014379f $X=0.885 $Y=0.515 $X2=0 $Y2=0
cc_275 N_X_c_432_n N_VGND_c_484_n 0.0118382f $X=0.885 $Y=0.515 $X2=0 $Y2=0
cc_276 N_VGND_c_476_n N_A_349_74#_c_533_n 0.0255177f $X=1.385 $Y=0.515 $X2=0
+ $Y2=0
cc_277 N_VGND_c_477_n N_A_349_74#_c_533_n 0.0191765f $X=2.385 $Y=0.675 $X2=0
+ $Y2=0
cc_278 N_VGND_c_481_n N_A_349_74#_c_533_n 0.0144922f $X=2.22 $Y=0 $X2=0 $Y2=0
cc_279 N_VGND_c_484_n N_A_349_74#_c_533_n 0.0118826f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_280 N_VGND_M1011_d N_A_349_74#_c_534_n 0.00358162f $X=2.175 $Y=0.37 $X2=0
+ $Y2=0
cc_281 N_VGND_c_477_n N_A_349_74#_c_534_n 0.0248957f $X=2.385 $Y=0.675 $X2=0
+ $Y2=0
cc_282 N_VGND_c_476_n N_A_349_74#_c_535_n 0.00584871f $X=1.385 $Y=0.515 $X2=0
+ $Y2=0
cc_283 N_VGND_c_477_n N_A_349_74#_c_536_n 0.00795492f $X=2.385 $Y=0.675 $X2=0
+ $Y2=0
cc_284 N_VGND_c_483_n N_A_349_74#_c_536_n 0.0146502f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_285 N_VGND_c_484_n N_A_349_74#_c_536_n 0.0120674f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_286 N_VGND_c_483_n N_A_349_74#_c_537_n 0.0518789f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_287 N_VGND_c_484_n N_A_349_74#_c_537_n 0.0447063f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_288 N_VGND_c_483_n N_A_349_74#_c_538_n 0.0115764f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_289 N_VGND_c_484_n N_A_349_74#_c_538_n 0.00959296f $X=4.56 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__dlxbn_2.spice
* Created: Fri Aug 28 17:28:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dlxbn_2.pex.spice"
.subckt sky130_fd_sc_ms__dlxbn_2  VNB VPB D GATE_N VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1018 N_VGND_M1018_d N_D_M1018_g N_A_27_136#_M1018_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.171076 AS=0.15675 PD=1.27054 PS=1.67 NRD=55.86 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1001 N_A_232_98#_M1001_d N_GATE_N_M1001_g N_VGND_M1018_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.230174 PD=2.05 PS=1.70946 NRD=0 NRS=41.52 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A_232_98#_M1004_g N_A_343_74#_M1004_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.206959 AS=0.2817 PD=1.49609 PS=2.29 NRD=36.432 NRS=2.016 M=1
+ R=4.93333 SA=75000.3 SB=75002.2 A=0.111 P=1.78 MULT=1
MM1012 A_569_79# N_A_27_136#_M1012_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.178991 PD=0.88 PS=1.29391 NRD=12.18 NRS=18.744 M=1 R=4.26667
+ SA=75000.9 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1013 N_A_647_79#_M1013_d N_A_232_98#_M1013_g A_569_79# VNB NLOWVT L=0.15
+ W=0.64 AD=0.238611 AS=0.0768 PD=1.75094 PS=0.88 NRD=27.18 NRS=12.18 M=1
+ R=4.26667 SA=75001.3 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1025 A_839_123# N_A_343_74#_M1025_g N_A_647_79#_M1013_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0651 AS=0.156589 PD=0.73 PS=1.14906 NRD=28.56 NRS=0 M=1 R=2.8
+ SA=75002.3 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_A_887_270#_M1022_g A_839_123# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0905534 AS=0.0651 PD=0.829138 PS=0.73 NRD=7.14 NRS=28.56 M=1 R=2.8
+ SA=75002.7 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1015 N_A_887_270#_M1015_d N_A_647_79#_M1015_g N_VGND_M1022_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.159547 PD=2.05 PS=1.46086 NRD=0 NRS=16.212 M=1 R=4.93333
+ SA=75001.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_Q_M1002_d N_A_887_270#_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1008 N_Q_M1002_d N_A_887_270#_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.166607 PD=1.02 PS=1.25478 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.6 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1016 N_A_1442_94#_M1016_d N_A_887_270#_M1016_g N_VGND_M1008_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.144093 PD=1.85 PS=1.08522 NRD=0 NRS=15.468 M=1
+ R=4.26667 SA=75001.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_Q_N_M1007_d N_A_1442_94#_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.3 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1014 N_Q_N_M1007_d N_A_1442_94#_M1014_g N_VGND_M1014_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1020 N_VPWR_M1020_d N_D_M1020_g N_A_27_136#_M1020_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1344 AS=0.3066 PD=1.16 PS=2.41 NRD=0 NRS=18.7544 M=1 R=4.66667 SA=90000.3
+ SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1019 N_A_232_98#_M1019_d N_GATE_N_M1019_g N_VPWR_M1020_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.1344 PD=2.24 PS=1.16 NRD=0 NRS=10.5395 M=1 R=4.66667
+ SA=90000.8 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1023 N_VPWR_M1023_d N_A_232_98#_M1023_g N_A_343_74#_M1023_s VPB PSHORT L=0.18
+ W=0.84 AD=0.156587 AS=0.2352 PD=1.23717 PS=2.24 NRD=19.9167 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90002.1 A=0.1512 P=2.04 MULT=1
MM1011 A_568_392# N_A_27_136#_M1011_g N_VPWR_M1023_d VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.186413 PD=1.24 PS=1.47283 NRD=12.7853 NRS=0 M=1 R=5.55556
+ SA=90000.6 SB=90001.4 A=0.18 P=2.36 MULT=1
MM1017 N_A_647_79#_M1017_d N_A_343_74#_M1017_g A_568_392# VPB PSHORT L=0.18 W=1
+ AD=0.292887 AS=0.12 PD=2.3169 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556
+ SA=90001.1 SB=90001 A=0.18 P=2.36 MULT=1
MM1006 A_817_392# N_A_232_98#_M1006_g N_A_647_79#_M1017_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0735 AS=0.123013 PD=0.77 PS=0.973099 NRD=56.2829 NRS=0 M=1
+ R=2.33333 SA=90002 SB=90001.4 A=0.0756 P=1.2 MULT=1
MM1021 N_VPWR_M1021_d N_A_887_270#_M1021_g A_817_392# VPB PSHORT L=0.18 W=0.42
+ AD=0.128591 AS=0.0735 PD=0.875455 PS=0.77 NRD=56.2829 NRS=56.2829 M=1
+ R=2.33333 SA=90002.5 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1009 N_A_887_270#_M1009_d N_A_647_79#_M1009_g N_VPWR_M1021_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.342909 PD=2.8 PS=2.33455 NRD=0 NRS=14.9326 M=1 R=6.22222
+ SA=90001.4 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_887_270#_M1000_g N_Q_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1024 N_VPWR_M1024_d N_A_887_270#_M1024_g N_Q_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.187547 AS=0.1512 PD=1.52679 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1010 N_A_1442_94#_M1010_d N_A_887_270#_M1010_g N_VPWR_M1024_d VPB PSHORT
+ L=0.18 W=1 AD=0.28 AS=0.167453 PD=2.56 PS=1.36321 NRD=0 NRS=9.8303 M=1
+ R=5.55556 SA=90001.1 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1003 N_Q_N_M1003_d N_A_1442_94#_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1005 N_Q_N_M1003_d N_A_1442_94#_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX26_noxref VNB VPB NWDIODE A=17.67 P=22.72
c_94 VNB 0 1.28661e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__dlxbn_2.pxi.spice"
*
.ends
*
*

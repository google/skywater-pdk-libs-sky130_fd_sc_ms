* File: sky130_fd_sc_ms__o21ba_1.pex.spice
* Created: Wed Sep  2 12:22:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O21BA_1%A1 2 3 5 8 9 10 14 16
r29 14 16 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.395 $Y=1.295
+ $X2=0.395 $Y2=1.13
r30 9 10 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.665
r31 9 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.295 $X2=0.385 $Y2=1.295
r32 8 16 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=0.495 $Y=0.69
+ $X2=0.495 $Y2=1.13
r33 3 5 152.633 $w=1.8e-07 $l=5.7e-07 $layer=POLY_cond $X=0.505 $Y=1.89
+ $X2=0.505 $Y2=2.46
r34 2 3 43.7431 $w=2.92e-07 $l=3.15238e-07 $layer=POLY_cond $X=0.395 $Y=1.625
+ $X2=0.505 $Y2=1.89
r35 1 14 1.64869 $w=3.5e-07 $l=1e-08 $layer=POLY_cond $X=0.395 $Y=1.305
+ $X2=0.395 $Y2=1.295
r36 1 2 52.7581 $w=3.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.395 $Y=1.305
+ $X2=0.395 $Y2=1.625
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_1%A2 3 7 9 10 11 12 13 17
r39 12 13 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.075 $Y=1.295
+ $X2=1.075 $Y2=1.665
r40 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1 $Y=1.295
+ $X2=1 $Y2=1.295
r41 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1 $Y=1.635 $X2=1
+ $Y2=1.295
r42 10 11 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.635 $X2=1
+ $Y2=1.8
r43 9 17 42.4377 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.13 $X2=1
+ $Y2=1.295
r44 7 9 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.065 $Y=0.69
+ $X2=1.065 $Y2=1.13
r45 3 11 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=0.925 $Y=2.46
+ $X2=0.925 $Y2=1.8
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_1%A_281_244# 1 2 9 13 17 19 21 22 25 27 29 33
+ 36
c58 9 0 1.91607e-19 $X=1.495 $Y=2.46
r59 30 33 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.22 $Y=0.845
+ $X2=2.555 $Y2=0.845
r60 25 27 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.305 $Y=1.985
+ $X2=2.52 $Y2=1.985
r61 23 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=1.01
+ $X2=2.22 $Y2=0.845
r62 23 29 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.22 $Y=1.01
+ $X2=2.22 $Y2=1.22
r63 22 36 29.847 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.14 $Y=1.385
+ $X2=1.975 $Y2=1.385
r64 21 29 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.14 $Y=1.385
+ $X2=2.14 $Y2=1.22
r65 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.385 $X2=2.14 $Y2=1.385
r66 19 25 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=2.14 $Y=1.82
+ $X2=2.305 $Y2=1.985
r67 19 21 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=2.14 $Y=1.82
+ $X2=2.14 $Y2=1.385
r68 16 17 2.30962 $w=2.9e-07 $l=9e-08 $layer=POLY_cond $X=1.585 $Y=1.365
+ $X2=1.495 $Y2=1.365
r69 16 36 80.672 $w=2.9e-07 $l=3.9e-07 $layer=POLY_cond $X=1.585 $Y=1.365
+ $X2=1.975 $Y2=1.365
r70 11 17 31.696 $w=1.65e-07 $l=1.52315e-07 $layer=POLY_cond $X=1.51 $Y=1.22
+ $X2=1.495 $Y2=1.365
r71 11 13 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.51 $Y=1.22
+ $X2=1.51 $Y2=0.69
r72 7 17 31.696 $w=1.65e-07 $l=1.45e-07 $layer=POLY_cond $X=1.495 $Y=1.51
+ $X2=1.495 $Y2=1.365
r73 7 9 369.274 $w=1.8e-07 $l=9.5e-07 $layer=POLY_cond $X=1.495 $Y=1.51
+ $X2=1.495 $Y2=2.46
r74 2 27 600 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=1 $X=2.305
+ $Y=1.84 $X2=2.52 $Y2=1.985
r75 1 33 182 $w=1.7e-07 $l=4.81871e-07 $layer=licon1_NDIFF $count=1 $X=2.195
+ $Y=0.56 $X2=2.555 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_1%B1_N 3 7 8 11 13
c36 3 0 9.93607e-20 $X=2.75 $Y=2.26
r37 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.385
+ $X2=2.68 $Y2=1.55
r38 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.385
+ $X2=2.68 $Y2=1.22
r39 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.385 $X2=2.68 $Y2=1.385
r40 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.68 $Y=1.295 $X2=2.68
+ $Y2=1.385
r41 7 13 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=2.77 $Y=0.835
+ $X2=2.77 $Y2=1.22
r42 3 14 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=2.75 $Y=2.26 $X2=2.75
+ $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_1%A_203_392# 1 2 9 13 19 22 23 26 28 32 33 37
+ 38
c82 28 0 1.91607e-19 $X=1.22 $Y=2.135
r83 38 42 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=3.255 $Y=1.485
+ $X2=3.255 $Y2=1.65
r84 38 41 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=3.255 $Y=1.485
+ $X2=3.255 $Y2=1.32
r85 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.25
+ $Y=1.485 $X2=3.25 $Y2=1.485
r86 34 37 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.14 $Y=1.485
+ $X2=3.25 $Y2=1.485
r87 31 32 7.80118 $w=5.18e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=2.23
+ $X2=1.785 $Y2=2.23
r88 28 31 11.0407 $w=5.18e-07 $l=4.8e-07 $layer=LI1_cond $X=1.22 $Y=2.23 $X2=1.7
+ $Y2=2.23
r89 25 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=1.65
+ $X2=3.14 $Y2=1.485
r90 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.14 $Y=1.65
+ $X2=3.14 $Y2=2.32
r91 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.055 $Y=2.405
+ $X2=3.14 $Y2=2.32
r92 23 32 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=3.055 $Y=2.405
+ $X2=1.785 $Y2=2.405
r93 22 31 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=1.7 $Y=1.97 $X2=1.7
+ $Y2=2.23
r94 22 33 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.7 $Y=1.97 $X2=1.7
+ $Y2=1.03
r95 17 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.78 $Y=0.865
+ $X2=1.78 $Y2=1.03
r96 17 19 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=1.78 $Y=0.865
+ $X2=1.78 $Y2=0.515
r97 13 41 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.34 $Y=0.74
+ $X2=3.34 $Y2=1.32
r98 9 42 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=3.335 $Y=2.4
+ $X2=3.335 $Y2=1.65
r99 2 28 300 $w=1.7e-07 $l=6.08933e-07 $layer=licon1_PDIFF $count=2 $X=1.015
+ $Y=1.96 $X2=1.22 $Y2=2.475
r100 2 28 600 $w=1.7e-07 $l=2.79106e-07 $layer=licon1_PDIFF $count=1 $X=1.015
+ $Y=1.96 $X2=1.22 $Y2=2.135
r101 1 19 91 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=2 $X=1.585
+ $Y=0.37 $X2=1.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_1%VPWR 1 2 3 10 12 18 22 24 26 31 38 39 45 48
r45 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 39 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r50 36 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.225 $Y=3.33
+ $X2=3.06 $Y2=3.33
r51 36 38 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.225 $Y=3.33
+ $X2=3.6 $Y2=3.33
r52 35 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r53 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.885 $Y=3.33
+ $X2=1.72 $Y2=3.33
r55 32 34 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.885 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 31 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=3.06 $Y2=3.33
r57 31 34 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=2.64 $Y2=3.33
r58 30 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r59 30 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r60 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r61 27 42 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r62 27 29 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=1.2 $Y2=3.33
r63 26 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.72 $Y2=3.33
r64 26 29 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.2 $Y2=3.33
r65 24 35 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r66 24 46 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r67 20 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.06 $Y=3.245
+ $X2=3.06 $Y2=3.33
r68 20 22 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.06 $Y=3.245
+ $X2=3.06 $Y2=2.78
r69 16 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=3.245
+ $X2=1.72 $Y2=3.33
r70 16 18 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.72 $Y=3.245
+ $X2=1.72 $Y2=2.78
r71 12 15 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.28 $Y=2.135
+ $X2=0.28 $Y2=2.815
r72 10 42 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r73 10 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r74 3 22 600 $w=1.7e-07 $l=1.04422e-06 $layer=licon1_PDIFF $count=1 $X=2.84
+ $Y=1.84 $X2=3.06 $Y2=2.78
r75 2 18 600 $w=1.7e-07 $l=8.84929e-07 $layer=licon1_PDIFF $count=1 $X=1.585
+ $Y=1.96 $X2=1.72 $Y2=2.78
r76 1 15 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r77 1 12 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_1%X 1 2 9 13 14 15 16 23 32
c26 14 0 9.93607e-20 $X=3.515 $Y=1.95
r27 21 23 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=3.575 $Y=2 $X2=3.575
+ $Y2=2.035
r28 15 16 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.575 $Y=2.405
+ $X2=3.575 $Y2=2.775
r29 14 21 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=3.575 $Y=1.975
+ $X2=3.575 $Y2=2
r30 14 32 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=3.575 $Y=1.975
+ $X2=3.575 $Y2=1.82
r31 14 15 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=3.575 $Y=2.06
+ $X2=3.575 $Y2=2.405
r32 14 23 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=3.575 $Y=2.06
+ $X2=3.575 $Y2=2.035
r33 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.67 $Y=1.13 $X2=3.67
+ $Y2=1.82
r34 7 13 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=3.572 $Y=0.948
+ $X2=3.572 $Y2=1.13
r35 7 9 13.6714 $w=3.63e-07 $l=4.33e-07 $layer=LI1_cond $X=3.572 $Y=0.948
+ $X2=3.572 $Y2=0.515
r36 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=1.84 $X2=3.56 $Y2=1.985
r37 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=1.84 $X2=3.56 $Y2=2.815
r38 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.415
+ $Y=0.37 $X2=3.555 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_1%A_27_74# 1 2 9 11 12 15
r27 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.28 $Y=0.79
+ $X2=1.28 $Y2=0.515
r28 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.115 $Y=0.875
+ $X2=1.28 $Y2=0.79
r29 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=0.875
+ $X2=0.445 $Y2=0.875
r30 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.79
+ $X2=0.445 $Y2=0.875
r31 7 9 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.28 $Y=0.79 $X2=0.28
+ $Y2=0.515
r32 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.14
+ $Y=0.37 $X2=1.28 $Y2=0.515
r33 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O21BA_1%VGND 1 2 9 13 15 17 22 32 33 36 39
r40 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r41 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r42 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r43 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r44 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.22 $Y=0 $X2=3.055
+ $Y2=0
r45 30 32 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.22 $Y=0 $X2=3.6
+ $Y2=0
r46 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r47 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r48 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r49 25 28 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r50 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r51 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r52 23 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r53 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=3.055
+ $Y2=0
r54 22 28 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=2.64
+ $Y2=0
r55 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r56 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r57 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r58 17 19 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r59 15 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r60 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r61 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.055 $Y=0.085
+ $X2=3.055 $Y2=0
r62 11 13 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.055 $Y=0.085
+ $X2=3.055 $Y2=0.495
r63 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0
r64 7 9 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0.525
r65 2 13 91 $w=1.7e-07 $l=3.10805e-07 $layer=licon1_NDIFF $count=2 $X=2.845
+ $Y=0.56 $X2=3.125 $Y2=0.495
r66 1 9 182 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.525
.ends


* File: sky130_fd_sc_ms__nand3b_4.spice
* Created: Wed Sep  2 12:14:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nand3b_4.pex.spice"
.subckt sky130_fd_sc_ms__nand3b_4  VNB VPB A_N C B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* C	C
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_N_M1000_g N_A_89_172#_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.203425 AS=0.19515 PD=1.425 PS=2.05 NRD=35.652 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1006 N_A_297_82#_M1006_d N_C_M1006_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.203425 PD=1.02 PS=1.425 NRD=0 NRS=35.652 M=1 R=4.93333
+ SA=75000.8 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1010 N_A_297_82#_M1006_d N_C_M1010_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2715 PD=1.02 PS=1.56 NRD=0 NRS=50.568 M=1 R=4.93333 SA=75001.2
+ SB=75001.4 A=0.111 P=1.78 MULT=1
MM1011 N_A_297_82#_M1011_d N_C_M1011_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2715 PD=1.09 PS=1.56 NRD=0 NRS=50.568 M=1 R=4.93333 SA=75002
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1012 N_A_297_82#_M1011_d N_C_M1012_g N_VGND_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.19935 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_A_744_74#_M1005_d N_A_89_172#_M1005_g N_Y_M1005_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1962 AS=0.11285 PD=2.05 PS=1.045 NRD=0 NRS=1.62 M=1 R=4.93333
+ SA=75000.2 SB=75003.3 A=0.111 P=1.78 MULT=1
MM1013 N_A_744_74#_M1013_d N_A_89_172#_M1013_g N_Y_M1005_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.11285 PD=1.02 PS=1.045 NRD=0 NRS=2.424 M=1 R=4.93333
+ SA=75000.6 SB=75002.8 A=0.111 P=1.78 MULT=1
MM1014 N_A_744_74#_M1013_d N_A_89_172#_M1014_g N_Y_M1014_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75002.4 A=0.111 P=1.78 MULT=1
MM1019 N_A_744_74#_M1019_d N_A_89_172#_M1019_g N_Y_M1014_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75002 A=0.111 P=1.78 MULT=1
MM1003 N_A_744_74#_M1019_d N_B_M1003_g N_A_297_82#_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1007 N_A_744_74#_M1007_d N_B_M1007_g N_A_297_82#_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1015 N_A_744_74#_M1007_d N_B_M1015_g N_A_297_82#_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.9 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1016 N_A_744_74#_M1016_d N_B_M1016_g N_A_297_82#_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1976 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1017 N_A_89_172#_M1017_d N_A_N_M1017_g N_VPWR_M1017_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.5628 PD=1.11 PS=3.02 NRD=0 NRS=90.2851 M=1 R=4.66667 SA=90000.6
+ SB=90006.5 A=0.1512 P=2.04 MULT=1
MM1020 N_A_89_172#_M1017_d N_A_N_M1020_g N_VPWR_M1020_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.519 PD=1.11 PS=1.90286 NRD=0 NRS=131.99 M=1 R=4.66667 SA=90001
+ SB=90006 A=0.1512 P=2.04 MULT=1
MM1001 N_VPWR_M1020_s N_C_M1001_g N_Y_M1001_s VPB PSHORT L=0.18 W=1.12 AD=0.692
+ AS=0.1512 PD=2.53714 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002 SB=90004.7
+ A=0.2016 P=2.6 MULT=1
MM1018 N_VPWR_M1018_d N_C_M1018_g N_Y_M1001_s VPB PSHORT L=0.18 W=1.12 AD=0.2436
+ AS=0.1512 PD=1.555 PS=1.39 NRD=13.1793 NRS=0 M=1 R=6.22222 SA=90002.4
+ SB=90004.3 A=0.2016 P=2.6 MULT=1
MM1008 N_VPWR_M1018_d N_A_89_172#_M1008_g N_Y_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2436 AS=0.364 PD=1.555 PS=1.77 NRD=14.0658 NRS=0 M=1 R=6.22222 SA=90003
+ SB=90003.7 A=0.2016 P=2.6 MULT=1
MM1009 N_VPWR_M1009_d N_A_89_172#_M1009_g N_Y_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.4256 AS=0.364 PD=1.88 PS=1.77 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.9
+ SB=90002.8 A=0.2016 P=2.6 MULT=1
MM1002 N_Y_M1002_d N_B_M1002_g N_VPWR_M1009_d VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.4256 PD=1.39 PS=1.88 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.8 SB=90001.9
+ A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1002_d N_B_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=1.7304 PD=1.39 PS=5.33 NRD=0 NRS=36.051 M=1 R=6.22222 SA=90005.3 SB=90001.5
+ A=0.2016 P=2.6 MULT=1
DX21_noxref VNB VPB NWDIODE A=14.9916 P=19.84
c_99 VPB 0 1.70138e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__nand3b_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__xnor2_4.pxi.spice
* Created: Fri Aug 28 18:17:51 2020
* 
x_PM_SKY130_FD_SC_MS__XNOR2_4%A N_A_M1012_g N_A_M1019_g N_A_M1013_g N_A_M1028_g
+ N_A_M1002_g N_A_M1000_g N_A_M1009_g N_A_M1004_g N_A_M1021_g N_A_c_163_n
+ N_A_M1006_g N_A_c_151_n N_A_M1023_g N_A_c_165_n N_A_M1007_g A N_A_c_153_n
+ N_A_c_167_n N_A_c_154_n N_A_c_155_n N_A_c_156_n N_A_c_157_n N_A_c_158_n
+ PM_SKY130_FD_SC_MS__XNOR2_4%A
x_PM_SKY130_FD_SC_MS__XNOR2_4%B N_B_M1018_g N_B_M1022_g N_B_M1020_g N_B_M1026_g
+ N_B_c_335_n N_B_M1001_g N_B_M1003_g N_B_M1015_g N_B_M1005_g N_B_M1016_g
+ N_B_M1008_g N_B_c_338_n N_B_c_339_n N_B_M1011_g N_B_M1024_g N_B_c_342_n
+ N_B_c_343_n N_B_c_354_n N_B_c_355_n N_B_c_432_p N_B_c_344_n N_B_c_357_n
+ N_B_c_390_n N_B_c_345_n B B B B N_B_c_346_n PM_SKY130_FD_SC_MS__XNOR2_4%B
x_PM_SKY130_FD_SC_MS__XNOR2_4%A_119_368# N_A_119_368#_M1022_s
+ N_A_119_368#_M1012_d N_A_119_368#_M1018_d N_A_119_368#_M1025_g
+ N_A_119_368#_M1010_g N_A_119_368#_M1027_g N_A_119_368#_M1014_g
+ N_A_119_368#_M1017_g N_A_119_368#_c_549_n N_A_119_368#_c_538_n
+ N_A_119_368#_M1029_g N_A_119_368#_c_540_n N_A_119_368#_c_541_n
+ N_A_119_368#_c_552_n N_A_119_368#_c_553_n N_A_119_368#_c_573_n
+ N_A_119_368#_c_578_n N_A_119_368#_c_579_n N_A_119_368#_c_554_n
+ N_A_119_368#_c_542_n N_A_119_368#_c_543_n N_A_119_368#_c_544_n
+ N_A_119_368#_c_555_n N_A_119_368#_c_556_n N_A_119_368#_c_557_n
+ N_A_119_368#_c_558_n N_A_119_368#_c_545_n N_A_119_368#_c_559_n
+ N_A_119_368#_c_546_n PM_SKY130_FD_SC_MS__XNOR2_4%A_119_368#
x_PM_SKY130_FD_SC_MS__XNOR2_4%VPWR N_VPWR_M1012_s N_VPWR_M1013_s N_VPWR_M1020_s
+ N_VPWR_M1027_s N_VPWR_M1000_s N_VPWR_M1006_s N_VPWR_c_708_n N_VPWR_c_709_n
+ N_VPWR_c_710_n N_VPWR_c_711_n N_VPWR_c_712_n N_VPWR_c_713_n N_VPWR_c_714_n
+ N_VPWR_c_715_n VPWR N_VPWR_c_716_n N_VPWR_c_717_n N_VPWR_c_718_n
+ N_VPWR_c_707_n N_VPWR_c_720_n N_VPWR_c_721_n N_VPWR_c_722_n
+ PM_SKY130_FD_SC_MS__XNOR2_4%VPWR
x_PM_SKY130_FD_SC_MS__XNOR2_4%Y N_Y_M1010_s N_Y_M1017_s N_Y_M1025_d N_Y_M1003_d
+ N_Y_M1008_d N_Y_c_823_n N_Y_c_884_n N_Y_c_818_n N_Y_c_819_n N_Y_c_832_n
+ N_Y_c_820_n N_Y_c_857_n N_Y_c_821_n N_Y_c_822_n N_Y_c_867_n Y N_Y_c_843_n
+ PM_SKY130_FD_SC_MS__XNOR2_4%Y
x_PM_SKY130_FD_SC_MS__XNOR2_4%A_950_368# N_A_950_368#_M1000_d
+ N_A_950_368#_M1004_d N_A_950_368#_M1007_d N_A_950_368#_M1005_s
+ N_A_950_368#_M1011_s N_A_950_368#_c_952_n N_A_950_368#_c_945_n
+ N_A_950_368#_c_1005_n N_A_950_368#_c_946_n N_A_950_368#_c_947_n
+ N_A_950_368#_c_948_n N_A_950_368#_c_956_n N_A_950_368#_c_949_n
+ N_A_950_368#_c_950_n N_A_950_368#_c_951_n
+ PM_SKY130_FD_SC_MS__XNOR2_4%A_950_368#
x_PM_SKY130_FD_SC_MS__XNOR2_4%A_27_74# N_A_27_74#_M1019_d N_A_27_74#_M1028_d
+ N_A_27_74#_M1026_d N_A_27_74#_c_1011_n N_A_27_74#_c_1012_n N_A_27_74#_c_1013_n
+ N_A_27_74#_c_1014_n N_A_27_74#_c_1024_n N_A_27_74#_c_1015_n
+ PM_SKY130_FD_SC_MS__XNOR2_4%A_27_74#
x_PM_SKY130_FD_SC_MS__XNOR2_4%VGND N_VGND_M1019_s N_VGND_M1002_s N_VGND_M1021_s
+ N_VGND_M1001_d N_VGND_M1016_d N_VGND_c_1051_n N_VGND_c_1052_n N_VGND_c_1053_n
+ N_VGND_c_1054_n N_VGND_c_1055_n N_VGND_c_1056_n N_VGND_c_1057_n
+ N_VGND_c_1058_n N_VGND_c_1059_n N_VGND_c_1060_n N_VGND_c_1061_n VGND
+ N_VGND_c_1062_n N_VGND_c_1063_n N_VGND_c_1064_n N_VGND_c_1065_n
+ N_VGND_c_1066_n N_VGND_c_1067_n PM_SKY130_FD_SC_MS__XNOR2_4%VGND
x_PM_SKY130_FD_SC_MS__XNOR2_4%A_511_74# N_A_511_74#_M1010_d N_A_511_74#_M1014_d
+ N_A_511_74#_M1029_d N_A_511_74#_M1009_d N_A_511_74#_M1023_d
+ N_A_511_74#_M1015_s N_A_511_74#_M1024_s N_A_511_74#_c_1168_n
+ N_A_511_74#_c_1169_n N_A_511_74#_c_1170_n N_A_511_74#_c_1217_n
+ N_A_511_74#_c_1171_n N_A_511_74#_c_1178_n N_A_511_74#_c_1180_n
+ N_A_511_74#_c_1182_n N_A_511_74#_c_1183_n N_A_511_74#_c_1193_n
+ N_A_511_74#_c_1195_n N_A_511_74#_c_1172_n N_A_511_74#_c_1173_n
+ N_A_511_74#_c_1174_n N_A_511_74#_c_1175_n N_A_511_74#_c_1176_n
+ PM_SKY130_FD_SC_MS__XNOR2_4%A_511_74#
cc_1 VNB N_A_M1012_g 7.56802e-19 $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_2 VNB N_A_M1019_g 0.0371038f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_3 VNB N_A_M1013_g 4.9236e-19 $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.26
cc_4 VNB N_A_M1028_g 0.0276926f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.69
cc_5 VNB N_A_M1002_g 0.0260416f $X=-0.19 $Y=-0.245 $X2=4.94 $Y2=0.74
cc_6 VNB N_A_M1009_g 0.0251608f $X=-0.19 $Y=-0.245 $X2=5.53 $Y2=0.74
cc_7 VNB N_A_M1021_g 0.0251608f $X=-0.19 $Y=-0.245 $X2=5.96 $Y2=0.74
cc_8 VNB N_A_c_151_n 0.0977967f $X=-0.19 $Y=-0.245 $X2=6.55 $Y2=1.425
cc_9 VNB N_A_M1023_g 0.0298944f $X=-0.19 $Y=-0.245 $X2=6.55 $Y2=0.74
cc_10 VNB N_A_c_153_n 0.00561281f $X=-0.19 $Y=-0.245 $X2=4.415 $Y2=1.665
cc_11 VNB N_A_c_154_n 0.00326505f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.665
cc_12 VNB N_A_c_155_n 6.78237e-19 $X=-0.19 $Y=-0.245 $X2=4.56 $Y2=1.665
cc_13 VNB N_A_c_156_n 0.051872f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.485
cc_14 VNB N_A_c_157_n 0.00506297f $X=-0.19 $Y=-0.245 $X2=5.67 $Y2=1.515
cc_15 VNB N_A_c_158_n 4.06206e-19 $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.55
cc_16 VNB N_B_M1022_g 0.0297891f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_17 VNB N_B_M1026_g 0.0343393f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.69
cc_18 VNB N_B_c_335_n 0.0161782f $X=-0.19 $Y=-0.245 $X2=4.94 $Y2=1.35
cc_19 VNB N_B_M1015_g 0.0240473f $X=-0.19 $Y=-0.245 $X2=5.53 $Y2=0.74
cc_20 VNB N_B_M1016_g 0.0250428f $X=-0.19 $Y=-0.245 $X2=5.96 $Y2=0.74
cc_21 VNB N_B_c_338_n 0.012483f $X=-0.19 $Y=-0.245 $X2=6.55 $Y2=1.425
cc_22 VNB N_B_c_339_n 0.0784379f $X=-0.19 $Y=-0.245 $X2=6.55 $Y2=0.74
cc_23 VNB N_B_M1011_g 0.0133284f $X=-0.19 $Y=-0.245 $X2=6.815 $Y2=1.725
cc_24 VNB N_B_M1024_g 0.0358145f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.485
cc_25 VNB N_B_c_342_n 0.0112911f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.485
cc_26 VNB N_B_c_343_n 0.00348803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B_c_344_n 0.00178818f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.665
cc_28 VNB N_B_c_345_n 0.0447275f $X=-0.19 $Y=-0.245 $X2=4.56 $Y2=1.665
cc_29 VNB N_B_c_346_n 0.0042237f $X=-0.19 $Y=-0.245 $X2=5.67 $Y2=1.562
cc_30 VNB N_A_119_368#_M1010_g 0.0274838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_119_368#_M1014_g 0.0253545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_119_368#_M1017_g 0.0243566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_119_368#_c_538_n 0.0241313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_119_368#_M1029_g 0.0234833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_119_368#_c_540_n 0.0209789f $X=-0.19 $Y=-0.245 $X2=6.195 $Y2=2.4
cc_36 VNB N_A_119_368#_c_541_n 0.00693272f $X=-0.19 $Y=-0.245 $X2=6.195 $Y2=2.4
cc_37 VNB N_A_119_368#_c_542_n 0.0201514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_119_368#_c_543_n 0.00574833f $X=-0.19 $Y=-0.245 $X2=4.415
+ $Y2=1.665
cc_39 VNB N_A_119_368#_c_544_n 4.66653e-19 $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.665
cc_40 VNB N_A_119_368#_c_545_n 0.00385626f $X=-0.19 $Y=-0.245 $X2=4.99 $Y2=1.537
cc_41 VNB N_A_119_368#_c_546_n 0.0575257f $X=-0.19 $Y=-0.245 $X2=4.56 $Y2=1.562
cc_42 VNB N_VPWR_c_707_n 0.382608f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.485
cc_43 VNB N_Y_c_818_n 0.00312983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_Y_c_819_n 0.00294709f $X=-0.19 $Y=-0.245 $X2=5.53 $Y2=1.35
cc_45 VNB N_Y_c_820_n 0.0279518f $X=-0.19 $Y=-0.245 $X2=5.745 $Y2=2.4
cc_46 VNB N_Y_c_821_n 0.00558427f $X=-0.19 $Y=-0.245 $X2=6.195 $Y2=1.725
cc_47 VNB N_Y_c_822_n 0.0034915f $X=-0.19 $Y=-0.245 $X2=6.195 $Y2=2.4
cc_48 VNB N_A_27_74#_c_1011_n 0.0255089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_27_74#_c_1012_n 0.00664623f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.69
cc_50 VNB N_A_27_74#_c_1013_n 0.0118921f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.69
cc_51 VNB N_A_27_74#_c_1014_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_27_74#_c_1015_n 0.00808886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_1051_n 0.00640788f $X=-0.19 $Y=-0.245 $X2=4.94 $Y2=0.74
cc_54 VNB N_VGND_c_1052_n 0.00752608f $X=-0.19 $Y=-0.245 $X2=5.12 $Y2=2.4
cc_55 VNB N_VGND_c_1053_n 0.00790334f $X=-0.19 $Y=-0.245 $X2=5.53 $Y2=0.74
cc_56 VNB N_VGND_c_1054_n 0.00806735f $X=-0.19 $Y=-0.245 $X2=5.745 $Y2=2.4
cc_57 VNB N_VGND_c_1055_n 0.00790334f $X=-0.19 $Y=-0.245 $X2=5.96 $Y2=0.74
cc_58 VNB N_VGND_c_1056_n 0.100013f $X=-0.19 $Y=-0.245 $X2=6.195 $Y2=1.725
cc_59 VNB N_VGND_c_1057_n 0.00631651f $X=-0.19 $Y=-0.245 $X2=6.195 $Y2=2.4
cc_60 VNB N_VGND_c_1058_n 0.0178221f $X=-0.19 $Y=-0.245 $X2=6.55 $Y2=1.425
cc_61 VNB N_VGND_c_1059_n 0.00631651f $X=-0.19 $Y=-0.245 $X2=6.55 $Y2=0.74
cc_62 VNB N_VGND_c_1060_n 0.0178221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1061_n 0.00698918f $X=-0.19 $Y=-0.245 $X2=6.815 $Y2=1.725
cc_64 VNB N_VGND_c_1062_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.485
cc_65 VNB N_VGND_c_1063_n 0.0178221f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.485
cc_66 VNB N_VGND_c_1064_n 0.0187151f $X=-0.19 $Y=-0.245 $X2=4.99 $Y2=1.515
cc_67 VNB N_VGND_c_1065_n 0.477298f $X=-0.19 $Y=-0.245 $X2=4.99 $Y2=1.515
cc_68 VNB N_VGND_c_1066_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=5.67 $Y2=1.537
cc_69 VNB N_VGND_c_1067_n 0.00631651f $X=-0.19 $Y=-0.245 $X2=5.745 $Y2=1.537
cc_70 VNB N_A_511_74#_c_1168_n 0.00516301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_511_74#_c_1169_n 0.00280532f $X=-0.19 $Y=-0.245 $X2=5.53 $Y2=0.74
cc_72 VNB N_A_511_74#_c_1170_n 0.00489319f $X=-0.19 $Y=-0.245 $X2=5.53 $Y2=0.74
cc_73 VNB N_A_511_74#_c_1171_n 0.00501279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_511_74#_c_1172_n 0.00274314f $X=-0.19 $Y=-0.245 $X2=6.815 $Y2=2.4
cc_75 VNB N_A_511_74#_c_1173_n 0.00238751f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.485
cc_76 VNB N_A_511_74#_c_1174_n 0.00238751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_511_74#_c_1175_n 0.00238751f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.665
cc_78 VNB N_A_511_74#_c_1176_n 0.0446173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VPB N_A_M1012_g 0.0275985f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_80 VPB N_A_M1013_g 0.022431f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.26
cc_81 VPB N_A_M1000_g 0.0293978f $X=-0.19 $Y=1.66 $X2=5.12 $Y2=2.4
cc_82 VPB N_A_M1004_g 0.0222675f $X=-0.19 $Y=1.66 $X2=5.745 $Y2=2.4
cc_83 VPB N_A_c_163_n 0.0202756f $X=-0.19 $Y=1.66 $X2=6.195 $Y2=1.725
cc_84 VPB N_A_c_151_n 0.0312124f $X=-0.19 $Y=1.66 $X2=6.55 $Y2=1.425
cc_85 VPB N_A_c_165_n 0.0197759f $X=-0.19 $Y=1.66 $X2=6.815 $Y2=1.725
cc_86 VPB N_A_c_153_n 0.0163331f $X=-0.19 $Y=1.66 $X2=4.415 $Y2=1.665
cc_87 VPB N_A_c_167_n 0.00371688f $X=-0.19 $Y=1.66 $X2=1.345 $Y2=1.665
cc_88 VPB N_A_c_154_n 0.00264396f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.665
cc_89 VPB N_A_c_155_n 0.00286931f $X=-0.19 $Y=1.66 $X2=4.56 $Y2=1.665
cc_90 VPB N_A_c_157_n 0.0112353f $X=-0.19 $Y=1.66 $X2=5.67 $Y2=1.515
cc_91 VPB N_B_M1018_g 0.0202511f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_92 VPB N_B_M1020_g 0.0215392f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.26
cc_93 VPB N_B_M1003_g 0.019868f $X=-0.19 $Y=1.66 $X2=5.12 $Y2=2.4
cc_94 VPB N_B_M1005_g 0.0197619f $X=-0.19 $Y=1.66 $X2=5.745 $Y2=2.4
cc_95 VPB N_B_M1008_g 0.0200662f $X=-0.19 $Y=1.66 $X2=6.195 $Y2=2.4
cc_96 VPB N_B_c_339_n 0.00892093f $X=-0.19 $Y=1.66 $X2=6.55 $Y2=0.74
cc_97 VPB N_B_M1011_g 0.0293141f $X=-0.19 $Y=1.66 $X2=6.815 $Y2=1.725
cc_98 VPB N_B_c_354_n 0.00321634f $X=-0.19 $Y=1.66 $X2=4.415 $Y2=1.665
cc_99 VPB N_B_c_355_n 0.021855f $X=-0.19 $Y=1.66 $X2=1.345 $Y2=1.665
cc_100 VPB N_B_c_344_n 3.59843e-19 $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.665
cc_101 VPB N_B_c_357_n 0.00139419f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.665
cc_102 VPB N_B_c_345_n 0.011487f $X=-0.19 $Y=1.66 $X2=4.56 $Y2=1.665
cc_103 VPB N_B_c_346_n 0.01195f $X=-0.19 $Y=1.66 $X2=5.67 $Y2=1.562
cc_104 VPB N_A_119_368#_M1025_g 0.0229774f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_119_368#_M1027_g 0.0262012f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_119_368#_c_549_n 0.0772741f $X=-0.19 $Y=1.66 $X2=5.745 $Y2=2.4
cc_107 VPB N_A_119_368#_c_540_n 0.0129525f $X=-0.19 $Y=1.66 $X2=6.195 $Y2=2.4
cc_108 VPB N_A_119_368#_c_541_n 8.60627e-19 $X=-0.19 $Y=1.66 $X2=6.195 $Y2=2.4
cc_109 VPB N_A_119_368#_c_552_n 0.0372463f $X=-0.19 $Y=1.66 $X2=6.55 $Y2=0.74
cc_110 VPB N_A_119_368#_c_553_n 0.00950794f $X=-0.19 $Y=1.66 $X2=6.55 $Y2=0.74
cc_111 VPB N_A_119_368#_c_554_n 0.00311731f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.485
cc_112 VPB N_A_119_368#_c_555_n 0.0025368f $X=-0.19 $Y=1.66 $X2=4.56 $Y2=1.665
cc_113 VPB N_A_119_368#_c_556_n 0.00253374f $X=-0.19 $Y=1.66 $X2=4.56 $Y2=1.665
cc_114 VPB N_A_119_368#_c_557_n 0.0491514f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_119_368#_c_558_n 0.00579457f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.485
cc_116 VPB N_A_119_368#_c_559_n 0.00461368f $X=-0.19 $Y=1.66 $X2=6.195 $Y2=1.537
cc_117 VPB N_A_119_368#_c_546_n 0.0183485f $X=-0.19 $Y=1.66 $X2=4.56 $Y2=1.562
cc_118 VPB N_VPWR_c_708_n 0.0106521f $X=-0.19 $Y=1.66 $X2=4.94 $Y2=0.74
cc_119 VPB N_VPWR_c_709_n 0.0710817f $X=-0.19 $Y=1.66 $X2=5.12 $Y2=1.68
cc_120 VPB N_VPWR_c_710_n 0.0284114f $X=-0.19 $Y=1.66 $X2=5.53 $Y2=1.35
cc_121 VPB N_VPWR_c_711_n 0.0195396f $X=-0.19 $Y=1.66 $X2=5.53 $Y2=0.74
cc_122 VPB N_VPWR_c_712_n 0.0216916f $X=-0.19 $Y=1.66 $X2=5.745 $Y2=2.4
cc_123 VPB N_VPWR_c_713_n 0.00324402f $X=-0.19 $Y=1.66 $X2=5.745 $Y2=2.4
cc_124 VPB N_VPWR_c_714_n 0.0140797f $X=-0.19 $Y=1.66 $X2=5.96 $Y2=1.35
cc_125 VPB N_VPWR_c_715_n 0.0475504f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_716_n 0.0204556f $X=-0.19 $Y=1.66 $X2=6.815 $Y2=2.4
cc_127 VPB N_VPWR_c_717_n 0.0187544f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.665
cc_128 VPB N_VPWR_c_718_n 0.0583481f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.485
cc_129 VPB N_VPWR_c_707_n 0.108109f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.485
cc_130 VPB N_VPWR_c_720_n 0.0175982f $X=-0.19 $Y=1.66 $X2=4.99 $Y2=1.515
cc_131 VPB N_VPWR_c_721_n 0.0173161f $X=-0.19 $Y=1.66 $X2=5.96 $Y2=1.537
cc_132 VPB N_VPWR_c_722_n 0.0136173f $X=-0.19 $Y=1.66 $X2=4.99 $Y2=1.562
cc_133 VPB N_Y_c_823_n 0.0271881f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_Y_c_821_n 0.00335454f $X=-0.19 $Y=1.66 $X2=6.195 $Y2=1.725
cc_135 VPB N_A_950_368#_c_945_n 0.00284344f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_950_368#_c_946_n 0.0119149f $X=-0.19 $Y=1.66 $X2=5.53 $Y2=0.74
cc_137 VPB N_A_950_368#_c_947_n 0.0363596f $X=-0.19 $Y=1.66 $X2=5.745 $Y2=2.4
cc_138 VPB N_A_950_368#_c_948_n 0.00260564f $X=-0.19 $Y=1.66 $X2=5.96 $Y2=0.74
cc_139 VPB N_A_950_368#_c_949_n 0.0022923f $X=-0.19 $Y=1.66 $X2=6.55 $Y2=0.74
cc_140 VPB N_A_950_368#_c_950_n 0.0017942f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_950_368#_c_951_n 0.00123754f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=1.485
cc_142 N_A_M1013_g N_B_M1018_g 0.0217143f $X=0.955 $Y=2.26 $X2=0 $Y2=0
cc_143 N_A_c_153_n N_B_M1018_g 0.00171963f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_144 N_A_c_167_n N_B_M1018_g 0.00107433f $X=1.345 $Y=1.665 $X2=0 $Y2=0
cc_145 N_A_M1028_g N_B_M1022_g 0.0219955f $X=0.995 $Y=0.69 $X2=0 $Y2=0
cc_146 N_A_c_154_n N_B_M1022_g 9.36198e-19 $X=1.2 $Y=1.665 $X2=0 $Y2=0
cc_147 N_A_c_153_n N_B_M1020_g 0.00726585f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_148 N_A_c_167_n N_B_M1020_g 2.02663e-19 $X=1.345 $Y=1.665 $X2=0 $Y2=0
cc_149 N_A_c_154_n N_B_M1020_g 3.47757e-19 $X=1.2 $Y=1.665 $X2=0 $Y2=0
cc_150 N_A_M1023_g N_B_c_335_n 0.0338967f $X=6.55 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A_c_151_n N_B_M1003_g 0.0507496f $X=6.55 $Y=1.425 $X2=0 $Y2=0
cc_152 N_A_c_151_n N_B_c_339_n 0.00582193f $X=6.55 $Y=1.425 $X2=0 $Y2=0
cc_153 N_A_M1023_g N_B_c_339_n 0.00452214f $X=6.55 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A_c_153_n N_B_c_343_n 0.00530645f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_155 N_A_c_153_n N_B_c_354_n 0.0122757f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_156 N_A_c_154_n N_B_c_354_n 0.00142845f $X=1.2 $Y=1.665 $X2=0 $Y2=0
cc_157 N_A_M1000_g N_B_c_355_n 0.0146568f $X=5.12 $Y=2.4 $X2=0 $Y2=0
cc_158 N_A_M1004_g N_B_c_355_n 0.0125087f $X=5.745 $Y=2.4 $X2=0 $Y2=0
cc_159 N_A_c_163_n N_B_c_355_n 0.0169867f $X=6.195 $Y=1.725 $X2=0 $Y2=0
cc_160 N_A_c_151_n N_B_c_355_n 0.00548353f $X=6.55 $Y=1.425 $X2=0 $Y2=0
cc_161 N_A_c_165_n N_B_c_355_n 0.00487002f $X=6.815 $Y=1.725 $X2=0 $Y2=0
cc_162 N_A_c_153_n N_B_c_355_n 0.065691f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_163 N_A_c_155_n N_B_c_355_n 0.00862409f $X=4.56 $Y=1.665 $X2=0 $Y2=0
cc_164 N_A_c_157_n N_B_c_355_n 0.0987207f $X=5.67 $Y=1.515 $X2=0 $Y2=0
cc_165 N_A_c_163_n N_B_c_344_n 6.31572e-19 $X=6.195 $Y=1.725 $X2=0 $Y2=0
cc_166 N_A_c_151_n N_B_c_344_n 0.0163714f $X=6.55 $Y=1.425 $X2=0 $Y2=0
cc_167 N_A_M1023_g N_B_c_344_n 0.00198641f $X=6.55 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A_c_157_n N_B_c_344_n 0.0142188f $X=5.67 $Y=1.515 $X2=0 $Y2=0
cc_169 N_A_c_163_n N_B_c_357_n 0.00441147f $X=6.195 $Y=1.725 $X2=0 $Y2=0
cc_170 N_A_c_165_n N_B_c_357_n 0.00391365f $X=6.815 $Y=1.725 $X2=0 $Y2=0
cc_171 N_A_c_157_n N_B_c_357_n 2.84442e-19 $X=5.67 $Y=1.515 $X2=0 $Y2=0
cc_172 N_A_c_153_n N_B_c_390_n 0.0195253f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_173 N_A_c_167_n N_B_c_390_n 0.00117519f $X=1.345 $Y=1.665 $X2=0 $Y2=0
cc_174 N_A_c_154_n N_B_c_390_n 0.0254288f $X=1.2 $Y=1.665 $X2=0 $Y2=0
cc_175 N_A_c_156_n N_B_c_390_n 2.33407e-19 $X=0.955 $Y=1.485 $X2=0 $Y2=0
cc_176 N_A_c_153_n N_B_c_345_n 0.00646557f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_177 N_A_c_167_n N_B_c_345_n 7.41198e-19 $X=1.345 $Y=1.665 $X2=0 $Y2=0
cc_178 N_A_c_154_n N_B_c_345_n 0.00477684f $X=1.2 $Y=1.665 $X2=0 $Y2=0
cc_179 N_A_c_156_n N_B_c_345_n 0.0281974f $X=0.955 $Y=1.485 $X2=0 $Y2=0
cc_180 N_A_c_151_n N_B_c_346_n 0.0175838f $X=6.55 $Y=1.425 $X2=0 $Y2=0
cc_181 N_A_M1023_g N_B_c_346_n 0.00317485f $X=6.55 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A_c_165_n N_B_c_346_n 0.00636874f $X=6.815 $Y=1.725 $X2=0 $Y2=0
cc_183 N_A_c_153_n N_A_119_368#_M1025_g 0.00249111f $X=4.415 $Y=1.665 $X2=0
+ $Y2=0
cc_184 N_A_c_153_n N_A_119_368#_M1027_g 0.00287541f $X=4.415 $Y=1.665 $X2=0
+ $Y2=0
cc_185 N_A_c_153_n N_A_119_368#_c_549_n 0.00218275f $X=4.415 $Y=1.665 $X2=0
+ $Y2=0
cc_186 N_A_c_155_n N_A_119_368#_c_549_n 0.0011884f $X=4.56 $Y=1.665 $X2=0 $Y2=0
cc_187 N_A_c_151_n N_A_119_368#_c_538_n 0.00603888f $X=6.55 $Y=1.425 $X2=0 $Y2=0
cc_188 N_A_c_153_n N_A_119_368#_c_538_n 0.00886514f $X=4.415 $Y=1.665 $X2=0
+ $Y2=0
cc_189 N_A_c_155_n N_A_119_368#_c_538_n 9.53184e-19 $X=4.56 $Y=1.665 $X2=0 $Y2=0
cc_190 N_A_c_157_n N_A_119_368#_c_538_n 0.00855692f $X=5.67 $Y=1.515 $X2=0 $Y2=0
cc_191 N_A_M1002_g N_A_119_368#_M1029_g 0.030803f $X=4.94 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A_c_153_n N_A_119_368#_c_540_n 0.00314716f $X=4.415 $Y=1.665 $X2=0
+ $Y2=0
cc_193 N_A_c_153_n N_A_119_368#_c_541_n 0.00121497f $X=4.415 $Y=1.665 $X2=0
+ $Y2=0
cc_194 N_A_c_157_n N_A_119_368#_c_541_n 0.00299094f $X=5.67 $Y=1.515 $X2=0 $Y2=0
cc_195 N_A_M1013_g N_A_119_368#_c_573_n 0.0136267f $X=0.955 $Y=2.26 $X2=0 $Y2=0
cc_196 N_A_c_153_n N_A_119_368#_c_573_n 0.00429022f $X=4.415 $Y=1.665 $X2=0
+ $Y2=0
cc_197 N_A_c_167_n N_A_119_368#_c_573_n 0.00840921f $X=1.345 $Y=1.665 $X2=0
+ $Y2=0
cc_198 N_A_c_154_n N_A_119_368#_c_573_n 0.0129635f $X=1.2 $Y=1.665 $X2=0 $Y2=0
cc_199 N_A_c_158_n N_A_119_368#_c_573_n 0.00765793f $X=1.085 $Y=1.55 $X2=0 $Y2=0
cc_200 N_A_c_153_n N_A_119_368#_c_578_n 0.00893565f $X=4.415 $Y=1.665 $X2=0
+ $Y2=0
cc_201 N_A_M1013_g N_A_119_368#_c_579_n 6.01608e-19 $X=0.955 $Y=2.26 $X2=0 $Y2=0
cc_202 N_A_c_153_n N_A_119_368#_c_542_n 0.00978895f $X=4.415 $Y=1.665 $X2=0
+ $Y2=0
cc_203 N_A_c_153_n N_A_119_368#_c_543_n 0.012739f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_204 N_A_c_153_n N_A_119_368#_c_544_n 0.0622782f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_205 N_A_c_155_n N_A_119_368#_c_544_n 0.001203f $X=4.56 $Y=1.665 $X2=0 $Y2=0
cc_206 N_A_c_157_n N_A_119_368#_c_544_n 0.0134513f $X=5.67 $Y=1.515 $X2=0 $Y2=0
cc_207 N_A_M1012_g N_A_119_368#_c_558_n 0.0142427f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_208 N_A_M1013_g N_A_119_368#_c_558_n 0.0142844f $X=0.955 $Y=2.26 $X2=0 $Y2=0
cc_209 N_A_c_156_n N_A_119_368#_c_558_n 0.00209661f $X=0.955 $Y=1.485 $X2=0
+ $Y2=0
cc_210 N_A_c_158_n N_A_119_368#_c_558_n 0.0275631f $X=1.085 $Y=1.55 $X2=0 $Y2=0
cc_211 N_A_c_153_n N_A_119_368#_c_545_n 0.00158684f $X=4.415 $Y=1.665 $X2=0
+ $Y2=0
cc_212 N_A_c_153_n N_A_119_368#_c_546_n 0.0046128f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_213 N_A_M1012_g N_VPWR_c_709_n 0.00873548f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_214 N_A_M1013_g N_VPWR_c_710_n 0.00283706f $X=0.955 $Y=2.26 $X2=0 $Y2=0
cc_215 N_A_M1012_g N_VPWR_c_712_n 0.00465228f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_216 N_A_M1013_g N_VPWR_c_712_n 0.00465228f $X=0.955 $Y=2.26 $X2=0 $Y2=0
cc_217 N_A_M1000_g N_VPWR_c_714_n 0.00336946f $X=5.12 $Y=2.4 $X2=0 $Y2=0
cc_218 N_A_M1004_g N_VPWR_c_714_n 0.00338835f $X=5.745 $Y=2.4 $X2=0 $Y2=0
cc_219 N_A_M1000_g N_VPWR_c_715_n 0.00374396f $X=5.12 $Y=2.4 $X2=0 $Y2=0
cc_220 N_A_M1004_g N_VPWR_c_717_n 0.0037329f $X=5.745 $Y=2.4 $X2=0 $Y2=0
cc_221 N_A_c_163_n N_VPWR_c_717_n 0.0037329f $X=6.195 $Y=1.725 $X2=0 $Y2=0
cc_222 N_A_c_165_n N_VPWR_c_718_n 0.00371808f $X=6.815 $Y=1.725 $X2=0 $Y2=0
cc_223 N_A_M1012_g N_VPWR_c_707_n 0.00555093f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_224 N_A_M1013_g N_VPWR_c_707_n 0.00555093f $X=0.955 $Y=2.26 $X2=0 $Y2=0
cc_225 N_A_M1000_g N_VPWR_c_707_n 0.00465707f $X=5.12 $Y=2.4 $X2=0 $Y2=0
cc_226 N_A_M1004_g N_VPWR_c_707_n 0.00461542f $X=5.745 $Y=2.4 $X2=0 $Y2=0
cc_227 N_A_c_163_n N_VPWR_c_707_n 0.00461505f $X=6.195 $Y=1.725 $X2=0 $Y2=0
cc_228 N_A_c_165_n N_VPWR_c_707_n 0.00459566f $X=6.815 $Y=1.725 $X2=0 $Y2=0
cc_229 N_A_c_163_n N_VPWR_c_722_n 0.00337218f $X=6.195 $Y=1.725 $X2=0 $Y2=0
cc_230 N_A_c_165_n N_VPWR_c_722_n 0.00154259f $X=6.815 $Y=1.725 $X2=0 $Y2=0
cc_231 N_A_M1000_g N_Y_c_823_n 0.0146556f $X=5.12 $Y=2.4 $X2=0 $Y2=0
cc_232 N_A_M1004_g N_Y_c_823_n 0.0125474f $X=5.745 $Y=2.4 $X2=0 $Y2=0
cc_233 N_A_c_163_n N_Y_c_823_n 0.0125275f $X=6.195 $Y=1.725 $X2=0 $Y2=0
cc_234 N_A_c_151_n N_Y_c_823_n 0.00100839f $X=6.55 $Y=1.425 $X2=0 $Y2=0
cc_235 N_A_c_165_n N_Y_c_823_n 0.0153314f $X=6.815 $Y=1.725 $X2=0 $Y2=0
cc_236 N_A_c_153_n N_Y_c_818_n 0.00304231f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_237 N_A_c_153_n N_Y_c_819_n 0.00164873f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_238 N_A_M1002_g N_Y_c_832_n 8.81742e-19 $X=4.94 $Y=0.74 $X2=0 $Y2=0
cc_239 N_A_M1002_g N_Y_c_820_n 0.0116256f $X=4.94 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A_M1009_g N_Y_c_820_n 0.0112794f $X=5.53 $Y=0.74 $X2=0 $Y2=0
cc_241 N_A_M1021_g N_Y_c_820_n 0.0155633f $X=5.96 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A_c_151_n N_Y_c_820_n 0.0205991f $X=6.55 $Y=1.425 $X2=0 $Y2=0
cc_243 N_A_M1023_g N_Y_c_820_n 0.0112304f $X=6.55 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A_c_153_n N_Y_c_820_n 7.74234e-19 $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_245 N_A_c_155_n N_Y_c_820_n 0.00229058f $X=4.56 $Y=1.665 $X2=0 $Y2=0
cc_246 N_A_c_157_n N_Y_c_820_n 0.105415f $X=5.67 $Y=1.515 $X2=0 $Y2=0
cc_247 N_A_c_153_n N_Y_c_822_n 0.0124755f $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_248 N_A_c_165_n Y 8.51526e-19 $X=6.815 $Y=1.725 $X2=0 $Y2=0
cc_249 N_A_c_165_n N_Y_c_843_n 8.01936e-19 $X=6.815 $Y=1.725 $X2=0 $Y2=0
cc_250 N_A_c_163_n N_A_950_368#_c_952_n 0.00987883f $X=6.195 $Y=1.725 $X2=0
+ $Y2=0
cc_251 N_A_c_165_n N_A_950_368#_c_952_n 0.0104237f $X=6.815 $Y=1.725 $X2=0 $Y2=0
cc_252 N_A_M1000_g N_A_950_368#_c_948_n 0.00579977f $X=5.12 $Y=2.4 $X2=0 $Y2=0
cc_253 N_A_M1004_g N_A_950_368#_c_948_n 8.35113e-19 $X=5.745 $Y=2.4 $X2=0 $Y2=0
cc_254 N_A_M1000_g N_A_950_368#_c_956_n 0.0104582f $X=5.12 $Y=2.4 $X2=0 $Y2=0
cc_255 N_A_M1004_g N_A_950_368#_c_956_n 0.00989875f $X=5.745 $Y=2.4 $X2=0 $Y2=0
cc_256 N_A_M1000_g N_A_950_368#_c_949_n 7.56466e-19 $X=5.12 $Y=2.4 $X2=0 $Y2=0
cc_257 N_A_M1004_g N_A_950_368#_c_949_n 0.00521412f $X=5.745 $Y=2.4 $X2=0 $Y2=0
cc_258 N_A_c_163_n N_A_950_368#_c_949_n 0.00520106f $X=6.195 $Y=1.725 $X2=0
+ $Y2=0
cc_259 N_A_c_165_n N_A_950_368#_c_949_n 7.58362e-19 $X=6.815 $Y=1.725 $X2=0
+ $Y2=0
cc_260 N_A_c_163_n N_A_950_368#_c_950_n 8.57558e-19 $X=6.195 $Y=1.725 $X2=0
+ $Y2=0
cc_261 N_A_c_165_n N_A_950_368#_c_950_n 0.00745278f $X=6.815 $Y=1.725 $X2=0
+ $Y2=0
cc_262 N_A_M1019_g N_A_27_74#_c_1011_n 4.43891e-19 $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_263 N_A_M1019_g N_A_27_74#_c_1012_n 0.0192715f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_264 N_A_M1028_g N_A_27_74#_c_1012_n 0.0139223f $X=0.995 $Y=0.69 $X2=0 $Y2=0
cc_265 N_A_c_153_n N_A_27_74#_c_1012_n 9.94348e-19 $X=4.415 $Y=1.665 $X2=0 $Y2=0
cc_266 N_A_c_167_n N_A_27_74#_c_1012_n 0.00253611f $X=1.345 $Y=1.665 $X2=0 $Y2=0
cc_267 N_A_c_156_n N_A_27_74#_c_1012_n 0.00433422f $X=0.955 $Y=1.485 $X2=0 $Y2=0
cc_268 N_A_c_158_n N_A_27_74#_c_1012_n 0.0599098f $X=1.085 $Y=1.55 $X2=0 $Y2=0
cc_269 N_A_M1028_g N_A_27_74#_c_1014_n 0.00303571f $X=0.995 $Y=0.69 $X2=0 $Y2=0
cc_270 N_A_M1019_g N_A_27_74#_c_1024_n 8.66511e-19 $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_271 N_A_M1028_g N_A_27_74#_c_1024_n 0.00539747f $X=0.995 $Y=0.69 $X2=0 $Y2=0
cc_272 N_A_M1019_g N_VGND_c_1051_n 0.0126947f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_273 N_A_M1028_g N_VGND_c_1051_n 0.00555362f $X=0.995 $Y=0.69 $X2=0 $Y2=0
cc_274 N_A_M1002_g N_VGND_c_1052_n 0.00231005f $X=4.94 $Y=0.74 $X2=0 $Y2=0
cc_275 N_A_M1009_g N_VGND_c_1052_n 0.00416335f $X=5.53 $Y=0.74 $X2=0 $Y2=0
cc_276 N_A_M1021_g N_VGND_c_1053_n 0.00416335f $X=5.96 $Y=0.74 $X2=0 $Y2=0
cc_277 N_A_M1023_g N_VGND_c_1053_n 0.00416335f $X=6.55 $Y=0.74 $X2=0 $Y2=0
cc_278 N_A_M1028_g N_VGND_c_1056_n 0.00433139f $X=0.995 $Y=0.69 $X2=0 $Y2=0
cc_279 N_A_M1002_g N_VGND_c_1056_n 0.00321293f $X=4.94 $Y=0.74 $X2=0 $Y2=0
cc_280 N_A_M1009_g N_VGND_c_1058_n 0.00324657f $X=5.53 $Y=0.74 $X2=0 $Y2=0
cc_281 N_A_M1021_g N_VGND_c_1058_n 0.00324657f $X=5.96 $Y=0.74 $X2=0 $Y2=0
cc_282 N_A_M1023_g N_VGND_c_1060_n 0.00324657f $X=6.55 $Y=0.74 $X2=0 $Y2=0
cc_283 N_A_M1019_g N_VGND_c_1062_n 0.00383152f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_284 N_A_M1019_g N_VGND_c_1065_n 0.00761198f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_285 N_A_M1028_g N_VGND_c_1065_n 0.00817147f $X=0.995 $Y=0.69 $X2=0 $Y2=0
cc_286 N_A_M1002_g N_VGND_c_1065_n 0.00411864f $X=4.94 $Y=0.74 $X2=0 $Y2=0
cc_287 N_A_M1009_g N_VGND_c_1065_n 0.0041114f $X=5.53 $Y=0.74 $X2=0 $Y2=0
cc_288 N_A_M1021_g N_VGND_c_1065_n 0.0041114f $X=5.96 $Y=0.74 $X2=0 $Y2=0
cc_289 N_A_M1023_g N_VGND_c_1065_n 0.00411237f $X=6.55 $Y=0.74 $X2=0 $Y2=0
cc_290 N_A_M1002_g N_A_511_74#_c_1171_n 0.00396171f $X=4.94 $Y=0.74 $X2=0 $Y2=0
cc_291 N_A_M1002_g N_A_511_74#_c_1178_n 0.0042743f $X=4.94 $Y=0.74 $X2=0 $Y2=0
cc_292 N_A_M1009_g N_A_511_74#_c_1178_n 7.80342e-19 $X=5.53 $Y=0.74 $X2=0 $Y2=0
cc_293 N_A_M1002_g N_A_511_74#_c_1180_n 0.00927675f $X=4.94 $Y=0.74 $X2=0 $Y2=0
cc_294 N_A_M1009_g N_A_511_74#_c_1180_n 0.00982687f $X=5.53 $Y=0.74 $X2=0 $Y2=0
cc_295 N_A_M1002_g N_A_511_74#_c_1182_n 0.00134994f $X=4.94 $Y=0.74 $X2=0 $Y2=0
cc_296 N_A_M1021_g N_A_511_74#_c_1183_n 0.00982687f $X=5.96 $Y=0.74 $X2=0 $Y2=0
cc_297 N_A_M1023_g N_A_511_74#_c_1183_n 0.00982687f $X=6.55 $Y=0.74 $X2=0 $Y2=0
cc_298 N_A_M1002_g N_A_511_74#_c_1173_n 8.79578e-19 $X=4.94 $Y=0.74 $X2=0 $Y2=0
cc_299 N_A_M1009_g N_A_511_74#_c_1173_n 0.00777472f $X=5.53 $Y=0.74 $X2=0 $Y2=0
cc_300 N_A_M1021_g N_A_511_74#_c_1173_n 0.00777472f $X=5.96 $Y=0.74 $X2=0 $Y2=0
cc_301 N_A_M1023_g N_A_511_74#_c_1173_n 8.79578e-19 $X=6.55 $Y=0.74 $X2=0 $Y2=0
cc_302 N_A_M1021_g N_A_511_74#_c_1174_n 8.79578e-19 $X=5.96 $Y=0.74 $X2=0 $Y2=0
cc_303 N_A_M1023_g N_A_511_74#_c_1174_n 0.00774728f $X=6.55 $Y=0.74 $X2=0 $Y2=0
cc_304 N_B_M1020_g N_A_119_368#_M1025_g 0.0272618f $X=1.855 $Y=2.26 $X2=0 $Y2=0
cc_305 N_B_c_354_n N_A_119_368#_M1025_g 0.00516554f $X=2.07 $Y=1.945 $X2=0 $Y2=0
cc_306 N_B_c_355_n N_A_119_368#_M1025_g 0.0144424f $X=6.365 $Y=2.03 $X2=0 $Y2=0
cc_307 N_B_c_355_n N_A_119_368#_M1027_g 0.0143082f $X=6.365 $Y=2.03 $X2=0 $Y2=0
cc_308 N_B_c_355_n N_A_119_368#_c_549_n 0.0150083f $X=6.365 $Y=2.03 $X2=0 $Y2=0
cc_309 N_B_c_355_n N_A_119_368#_c_538_n 0.0108663f $X=6.365 $Y=2.03 $X2=0 $Y2=0
cc_310 N_B_M1018_g N_A_119_368#_c_573_n 0.0132431f $X=1.405 $Y=2.26 $X2=0 $Y2=0
cc_311 N_B_M1018_g N_A_119_368#_c_578_n 0.00100736f $X=1.405 $Y=2.26 $X2=0 $Y2=0
cc_312 N_B_M1020_g N_A_119_368#_c_578_n 0.0025966f $X=1.855 $Y=2.26 $X2=0 $Y2=0
cc_313 N_B_c_390_n N_A_119_368#_c_578_n 0.0101037f $X=1.99 $Y=1.515 $X2=0 $Y2=0
cc_314 N_B_c_345_n N_A_119_368#_c_578_n 0.00147245f $X=1.99 $Y=1.515 $X2=0 $Y2=0
cc_315 N_B_M1018_g N_A_119_368#_c_579_n 0.00755332f $X=1.405 $Y=2.26 $X2=0 $Y2=0
cc_316 N_B_M1020_g N_A_119_368#_c_579_n 0.0113195f $X=1.855 $Y=2.26 $X2=0 $Y2=0
cc_317 N_B_M1018_g N_A_119_368#_c_554_n 0.00370781f $X=1.405 $Y=2.26 $X2=0 $Y2=0
cc_318 N_B_M1020_g N_A_119_368#_c_554_n 0.00214545f $X=1.855 $Y=2.26 $X2=0 $Y2=0
cc_319 N_B_M1026_g N_A_119_368#_c_542_n 0.0109028f $X=1.925 $Y=0.69 $X2=0 $Y2=0
cc_320 N_B_c_343_n N_A_119_368#_c_542_n 0.0129304f $X=2.07 $Y=1.68 $X2=0 $Y2=0
cc_321 N_B_c_390_n N_A_119_368#_c_542_n 0.00746228f $X=1.99 $Y=1.515 $X2=0 $Y2=0
cc_322 N_B_c_345_n N_A_119_368#_c_542_n 0.00109267f $X=1.99 $Y=1.515 $X2=0 $Y2=0
cc_323 N_B_M1026_g N_A_119_368#_c_543_n 0.00454544f $X=1.925 $Y=0.69 $X2=0 $Y2=0
cc_324 N_B_c_343_n N_A_119_368#_c_543_n 0.0195139f $X=2.07 $Y=1.68 $X2=0 $Y2=0
cc_325 N_B_c_355_n N_A_119_368#_c_543_n 0.00614033f $X=6.365 $Y=2.03 $X2=0 $Y2=0
cc_326 N_B_c_345_n N_A_119_368#_c_543_n 4.8736e-19 $X=1.99 $Y=1.515 $X2=0 $Y2=0
cc_327 N_B_c_355_n N_A_119_368#_c_544_n 0.0538853f $X=6.365 $Y=2.03 $X2=0 $Y2=0
cc_328 N_B_M1018_g N_A_119_368#_c_558_n 0.00124553f $X=1.405 $Y=2.26 $X2=0 $Y2=0
cc_329 N_B_M1022_g N_A_119_368#_c_545_n 0.00328898f $X=1.425 $Y=0.69 $X2=0 $Y2=0
cc_330 N_B_M1026_g N_A_119_368#_c_545_n 0.0125638f $X=1.925 $Y=0.69 $X2=0 $Y2=0
cc_331 N_B_c_390_n N_A_119_368#_c_545_n 0.0251134f $X=1.99 $Y=1.515 $X2=0 $Y2=0
cc_332 N_B_c_345_n N_A_119_368#_c_545_n 0.00423307f $X=1.99 $Y=1.515 $X2=0 $Y2=0
cc_333 N_B_M1020_g N_A_119_368#_c_559_n 0.0134811f $X=1.855 $Y=2.26 $X2=0 $Y2=0
cc_334 N_B_c_355_n N_A_119_368#_c_559_n 0.0100177f $X=6.365 $Y=2.03 $X2=0 $Y2=0
cc_335 N_B_c_432_p N_A_119_368#_c_559_n 0.00547814f $X=2.155 $Y=2.03 $X2=0 $Y2=0
cc_336 N_B_c_343_n N_A_119_368#_c_546_n 4.86818e-19 $X=2.07 $Y=1.68 $X2=0 $Y2=0
cc_337 N_B_c_355_n N_A_119_368#_c_546_n 0.0129307f $X=6.365 $Y=2.03 $X2=0 $Y2=0
cc_338 N_B_c_345_n N_A_119_368#_c_546_n 0.0182975f $X=1.99 $Y=1.515 $X2=0 $Y2=0
cc_339 N_B_c_354_n N_VPWR_M1020_s 0.00197747f $X=2.07 $Y=1.945 $X2=0 $Y2=0
cc_340 N_B_c_355_n N_VPWR_M1020_s 0.00632717f $X=6.365 $Y=2.03 $X2=0 $Y2=0
cc_341 N_B_c_432_p N_VPWR_M1020_s 0.0043466f $X=2.155 $Y=2.03 $X2=0 $Y2=0
cc_342 N_B_c_355_n N_VPWR_M1027_s 0.00796575f $X=6.365 $Y=2.03 $X2=0 $Y2=0
cc_343 N_B_c_355_n N_VPWR_M1000_s 0.00731925f $X=6.365 $Y=2.03 $X2=0 $Y2=0
cc_344 N_B_c_355_n N_VPWR_M1006_s 0.00595801f $X=6.365 $Y=2.03 $X2=0 $Y2=0
cc_345 N_B_c_357_n N_VPWR_M1006_s 0.00252309f $X=6.45 $Y=1.945 $X2=0 $Y2=0
cc_346 N_B_M1018_g N_VPWR_c_710_n 0.00126695f $X=1.405 $Y=2.26 $X2=0 $Y2=0
cc_347 N_B_M1018_g N_VPWR_c_716_n 0.00463504f $X=1.405 $Y=2.26 $X2=0 $Y2=0
cc_348 N_B_M1020_g N_VPWR_c_716_n 0.00366756f $X=1.855 $Y=2.26 $X2=0 $Y2=0
cc_349 N_B_M1003_g N_VPWR_c_718_n 0.00333926f $X=7.265 $Y=2.4 $X2=0 $Y2=0
cc_350 N_B_M1005_g N_VPWR_c_718_n 0.00333926f $X=7.715 $Y=2.4 $X2=0 $Y2=0
cc_351 N_B_M1008_g N_VPWR_c_718_n 0.00333926f $X=8.165 $Y=2.4 $X2=0 $Y2=0
cc_352 N_B_M1011_g N_VPWR_c_718_n 0.00333926f $X=8.615 $Y=2.4 $X2=0 $Y2=0
cc_353 N_B_M1018_g N_VPWR_c_707_n 0.00555093f $X=1.405 $Y=2.26 $X2=0 $Y2=0
cc_354 N_B_M1020_g N_VPWR_c_707_n 0.00555093f $X=1.855 $Y=2.26 $X2=0 $Y2=0
cc_355 N_B_M1003_g N_VPWR_c_707_n 0.00422798f $X=7.265 $Y=2.4 $X2=0 $Y2=0
cc_356 N_B_M1005_g N_VPWR_c_707_n 0.00422687f $X=7.715 $Y=2.4 $X2=0 $Y2=0
cc_357 N_B_M1008_g N_VPWR_c_707_n 0.00422687f $X=8.165 $Y=2.4 $X2=0 $Y2=0
cc_358 N_B_M1011_g N_VPWR_c_707_n 0.00426429f $X=8.615 $Y=2.4 $X2=0 $Y2=0
cc_359 N_B_c_355_n N_Y_M1025_d 0.00328051f $X=6.365 $Y=2.03 $X2=0 $Y2=0
cc_360 N_B_M1020_g N_Y_c_823_n 7.36526e-19 $X=1.855 $Y=2.26 $X2=0 $Y2=0
cc_361 N_B_M1003_g N_Y_c_823_n 0.0178867f $X=7.265 $Y=2.4 $X2=0 $Y2=0
cc_362 N_B_M1005_g N_Y_c_823_n 0.0067118f $X=7.715 $Y=2.4 $X2=0 $Y2=0
cc_363 N_B_c_355_n N_Y_c_823_n 0.248288f $X=6.365 $Y=2.03 $X2=0 $Y2=0
cc_364 N_B_c_346_n N_Y_c_823_n 0.0233129f $X=7.99 $Y=1.515 $X2=0 $Y2=0
cc_365 N_B_c_335_n N_Y_c_820_n 0.0106974f $X=6.98 $Y=1.185 $X2=0 $Y2=0
cc_366 N_B_M1015_g N_Y_c_820_n 0.0114133f $X=7.605 $Y=0.74 $X2=0 $Y2=0
cc_367 N_B_M1016_g N_Y_c_820_n 0.010959f $X=8.035 $Y=0.74 $X2=0 $Y2=0
cc_368 N_B_c_339_n N_Y_c_820_n 0.0204787f $X=8.255 $Y=1.425 $X2=0 $Y2=0
cc_369 N_B_M1024_g N_Y_c_820_n 0.00250202f $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_370 N_B_c_344_n N_Y_c_820_n 0.013861f $X=6.45 $Y=1.765 $X2=0 $Y2=0
cc_371 N_B_c_346_n N_Y_c_820_n 0.124065f $X=7.99 $Y=1.515 $X2=0 $Y2=0
cc_372 N_B_M1005_g N_Y_c_857_n 0.012931f $X=7.715 $Y=2.4 $X2=0 $Y2=0
cc_373 N_B_M1008_g N_Y_c_857_n 0.0149936f $X=8.165 $Y=2.4 $X2=0 $Y2=0
cc_374 N_B_c_339_n N_Y_c_857_n 5.01604e-19 $X=8.255 $Y=1.425 $X2=0 $Y2=0
cc_375 N_B_c_346_n N_Y_c_857_n 0.0340021f $X=7.99 $Y=1.515 $X2=0 $Y2=0
cc_376 N_B_M1016_g N_Y_c_821_n 0.0035594f $X=8.035 $Y=0.74 $X2=0 $Y2=0
cc_377 N_B_c_338_n N_Y_c_821_n 0.0152156f $X=8.525 $Y=1.425 $X2=0 $Y2=0
cc_378 N_B_c_339_n N_Y_c_821_n 0.0059337f $X=8.255 $Y=1.425 $X2=0 $Y2=0
cc_379 N_B_M1011_g N_Y_c_821_n 0.00865837f $X=8.615 $Y=2.4 $X2=0 $Y2=0
cc_380 N_B_M1024_g N_Y_c_821_n 0.00436712f $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_381 N_B_c_346_n N_Y_c_821_n 0.0324034f $X=7.99 $Y=1.515 $X2=0 $Y2=0
cc_382 N_B_M1005_g N_Y_c_867_n 5.7779e-19 $X=7.715 $Y=2.4 $X2=0 $Y2=0
cc_383 N_B_M1008_g N_Y_c_867_n 0.0119305f $X=8.165 $Y=2.4 $X2=0 $Y2=0
cc_384 N_B_M1011_g N_Y_c_867_n 0.0128516f $X=8.615 $Y=2.4 $X2=0 $Y2=0
cc_385 N_B_M1003_g Y 0.00339706f $X=7.265 $Y=2.4 $X2=0 $Y2=0
cc_386 N_B_M1005_g Y 0.00334408f $X=7.715 $Y=2.4 $X2=0 $Y2=0
cc_387 N_B_M1008_g Y 4.35184e-19 $X=8.165 $Y=2.4 $X2=0 $Y2=0
cc_388 N_B_M1003_g N_Y_c_843_n 0.00392468f $X=7.265 $Y=2.4 $X2=0 $Y2=0
cc_389 N_B_M1005_g N_Y_c_843_n 8.84614e-19 $X=7.715 $Y=2.4 $X2=0 $Y2=0
cc_390 N_B_c_339_n N_Y_c_843_n 5.73741e-19 $X=8.255 $Y=1.425 $X2=0 $Y2=0
cc_391 N_B_c_346_n N_Y_c_843_n 0.0234738f $X=7.99 $Y=1.515 $X2=0 $Y2=0
cc_392 N_B_c_355_n N_A_950_368#_M1000_d 0.00538903f $X=6.365 $Y=2.03 $X2=-0.19
+ $Y2=-0.245
cc_393 N_B_c_355_n N_A_950_368#_M1004_d 0.0054135f $X=6.365 $Y=2.03 $X2=0 $Y2=0
cc_394 N_B_M1003_g N_A_950_368#_c_945_n 0.0100488f $X=7.265 $Y=2.4 $X2=0 $Y2=0
cc_395 N_B_M1005_g N_A_950_368#_c_945_n 0.0139528f $X=7.715 $Y=2.4 $X2=0 $Y2=0
cc_396 N_B_M1008_g N_A_950_368#_c_946_n 0.0140221f $X=8.165 $Y=2.4 $X2=0 $Y2=0
cc_397 N_B_M1011_g N_A_950_368#_c_946_n 0.0149887f $X=8.615 $Y=2.4 $X2=0 $Y2=0
cc_398 N_B_M1003_g N_A_950_368#_c_950_n 2.29065e-19 $X=7.265 $Y=2.4 $X2=0 $Y2=0
cc_399 N_B_M1022_g N_A_27_74#_c_1012_n 0.00399373f $X=1.425 $Y=0.69 $X2=0 $Y2=0
cc_400 N_B_c_345_n N_A_27_74#_c_1012_n 0.0016396f $X=1.99 $Y=1.515 $X2=0 $Y2=0
cc_401 N_B_M1022_g N_A_27_74#_c_1014_n 0.00103489f $X=1.425 $Y=0.69 $X2=0 $Y2=0
cc_402 N_B_M1022_g N_A_27_74#_c_1024_n 0.00539747f $X=1.425 $Y=0.69 $X2=0 $Y2=0
cc_403 N_B_M1026_g N_A_27_74#_c_1024_n 5.54947e-19 $X=1.925 $Y=0.69 $X2=0 $Y2=0
cc_404 N_B_M1022_g N_A_27_74#_c_1015_n 0.0134011f $X=1.425 $Y=0.69 $X2=0 $Y2=0
cc_405 N_B_M1026_g N_A_27_74#_c_1015_n 0.0120063f $X=1.925 $Y=0.69 $X2=0 $Y2=0
cc_406 N_B_c_335_n N_VGND_c_1054_n 0.00432496f $X=6.98 $Y=1.185 $X2=0 $Y2=0
cc_407 N_B_M1015_g N_VGND_c_1054_n 0.00432496f $X=7.605 $Y=0.74 $X2=0 $Y2=0
cc_408 N_B_M1016_g N_VGND_c_1055_n 0.00416335f $X=8.035 $Y=0.74 $X2=0 $Y2=0
cc_409 N_B_M1024_g N_VGND_c_1055_n 0.00416335f $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_410 N_B_M1022_g N_VGND_c_1056_n 0.00291626f $X=1.425 $Y=0.69 $X2=0 $Y2=0
cc_411 N_B_M1026_g N_VGND_c_1056_n 0.00291649f $X=1.925 $Y=0.69 $X2=0 $Y2=0
cc_412 N_B_c_335_n N_VGND_c_1060_n 0.00324657f $X=6.98 $Y=1.185 $X2=0 $Y2=0
cc_413 N_B_M1015_g N_VGND_c_1063_n 0.00324657f $X=7.605 $Y=0.74 $X2=0 $Y2=0
cc_414 N_B_M1016_g N_VGND_c_1063_n 0.00324657f $X=8.035 $Y=0.74 $X2=0 $Y2=0
cc_415 N_B_M1024_g N_VGND_c_1064_n 0.00324657f $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_416 N_B_M1022_g N_VGND_c_1065_n 0.00359859f $X=1.425 $Y=0.69 $X2=0 $Y2=0
cc_417 N_B_M1026_g N_VGND_c_1065_n 0.00364778f $X=1.925 $Y=0.69 $X2=0 $Y2=0
cc_418 N_B_c_335_n N_VGND_c_1065_n 0.00411487f $X=6.98 $Y=1.185 $X2=0 $Y2=0
cc_419 N_B_M1015_g N_VGND_c_1065_n 0.0041139f $X=7.605 $Y=0.74 $X2=0 $Y2=0
cc_420 N_B_M1016_g N_VGND_c_1065_n 0.0041114f $X=8.035 $Y=0.74 $X2=0 $Y2=0
cc_421 N_B_M1024_g N_VGND_c_1065_n 0.00414797f $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_422 N_B_M1026_g N_A_511_74#_c_1168_n 0.00416658f $X=1.925 $Y=0.69 $X2=0 $Y2=0
cc_423 N_B_M1026_g N_A_511_74#_c_1170_n 0.00288917f $X=1.925 $Y=0.69 $X2=0 $Y2=0
cc_424 N_B_c_335_n N_A_511_74#_c_1193_n 0.00996083f $X=6.98 $Y=1.185 $X2=0 $Y2=0
cc_425 N_B_M1015_g N_A_511_74#_c_1193_n 0.00996083f $X=7.605 $Y=0.74 $X2=0 $Y2=0
cc_426 N_B_M1016_g N_A_511_74#_c_1195_n 0.00982687f $X=8.035 $Y=0.74 $X2=0 $Y2=0
cc_427 N_B_c_338_n N_A_511_74#_c_1195_n 6.23126e-19 $X=8.525 $Y=1.425 $X2=0
+ $Y2=0
cc_428 N_B_M1024_g N_A_511_74#_c_1195_n 0.0136762f $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_429 N_B_c_335_n N_A_511_74#_c_1174_n 0.00784562f $X=6.98 $Y=1.185 $X2=0 $Y2=0
cc_430 N_B_M1015_g N_A_511_74#_c_1174_n 8.61714e-19 $X=7.605 $Y=0.74 $X2=0 $Y2=0
cc_431 N_B_c_335_n N_A_511_74#_c_1175_n 8.61714e-19 $X=6.98 $Y=1.185 $X2=0 $Y2=0
cc_432 N_B_M1015_g N_A_511_74#_c_1175_n 0.00787306f $X=7.605 $Y=0.74 $X2=0 $Y2=0
cc_433 N_B_M1016_g N_A_511_74#_c_1175_n 0.00777472f $X=8.035 $Y=0.74 $X2=0 $Y2=0
cc_434 N_B_M1024_g N_A_511_74#_c_1175_n 8.79578e-19 $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_435 N_B_M1016_g N_A_511_74#_c_1176_n 0.00173277f $X=8.035 $Y=0.74 $X2=0 $Y2=0
cc_436 N_B_M1024_g N_A_511_74#_c_1176_n 0.0142624f $X=8.625 $Y=0.74 $X2=0 $Y2=0
cc_437 N_B_c_342_n N_A_511_74#_c_1176_n 2.29254e-19 $X=8.615 $Y=1.425 $X2=0
+ $Y2=0
cc_438 N_A_119_368#_c_573_n N_VPWR_M1013_s 0.00316737f $X=1.465 $Y=2.035 $X2=0
+ $Y2=0
cc_439 N_A_119_368#_c_559_n N_VPWR_M1020_s 0.0101251f $X=3.58 $Y=2.79 $X2=0
+ $Y2=0
cc_440 N_A_119_368#_c_559_n N_VPWR_M1027_s 0.00807841f $X=3.58 $Y=2.79 $X2=0
+ $Y2=0
cc_441 N_A_119_368#_c_558_n N_VPWR_c_709_n 0.0310168f $X=0.73 $Y=1.985 $X2=0
+ $Y2=0
cc_442 N_A_119_368#_c_573_n N_VPWR_c_710_n 0.0122197f $X=1.465 $Y=2.035 $X2=0
+ $Y2=0
cc_443 N_A_119_368#_c_554_n N_VPWR_c_710_n 0.0101219f $X=1.795 $Y=2.71 $X2=0
+ $Y2=0
cc_444 N_A_119_368#_c_558_n N_VPWR_c_710_n 0.0141452f $X=0.73 $Y=1.985 $X2=0
+ $Y2=0
cc_445 N_A_119_368#_M1025_g N_VPWR_c_711_n 0.00377953f $X=2.485 $Y=2.4 $X2=0
+ $Y2=0
cc_446 N_A_119_368#_M1027_g N_VPWR_c_711_n 0.00377953f $X=2.935 $Y=2.4 $X2=0
+ $Y2=0
cc_447 N_A_119_368#_c_559_n N_VPWR_c_711_n 0.0138438f $X=3.58 $Y=2.79 $X2=0
+ $Y2=0
cc_448 N_A_119_368#_c_558_n N_VPWR_c_712_n 0.00657675f $X=0.73 $Y=1.985 $X2=0
+ $Y2=0
cc_449 N_A_119_368#_c_552_n N_VPWR_c_715_n 0.0205254f $X=3.935 $Y=2.79 $X2=0
+ $Y2=0
cc_450 N_A_119_368#_c_555_n N_VPWR_c_715_n 0.0360898f $X=3.91 $Y=2.79 $X2=0
+ $Y2=0
cc_451 N_A_119_368#_c_559_n N_VPWR_c_715_n 0.00388367f $X=3.58 $Y=2.79 $X2=0
+ $Y2=0
cc_452 N_A_119_368#_c_554_n N_VPWR_c_716_n 0.00821095f $X=1.795 $Y=2.71 $X2=0
+ $Y2=0
cc_453 N_A_119_368#_c_559_n N_VPWR_c_716_n 0.00438681f $X=3.58 $Y=2.79 $X2=0
+ $Y2=0
cc_454 N_A_119_368#_M1025_g N_VPWR_c_707_n 0.0047145f $X=2.485 $Y=2.4 $X2=0
+ $Y2=0
cc_455 N_A_119_368#_M1027_g N_VPWR_c_707_n 0.0047145f $X=2.935 $Y=2.4 $X2=0
+ $Y2=0
cc_456 N_A_119_368#_c_552_n N_VPWR_c_707_n 0.0306241f $X=3.935 $Y=2.79 $X2=0
+ $Y2=0
cc_457 N_A_119_368#_c_554_n N_VPWR_c_707_n 0.0107033f $X=1.795 $Y=2.71 $X2=0
+ $Y2=0
cc_458 N_A_119_368#_c_555_n N_VPWR_c_707_n 0.0349577f $X=3.91 $Y=2.79 $X2=0
+ $Y2=0
cc_459 N_A_119_368#_c_558_n N_VPWR_c_707_n 0.00992028f $X=0.73 $Y=1.985 $X2=0
+ $Y2=0
cc_460 N_A_119_368#_c_559_n N_VPWR_c_707_n 0.0362835f $X=3.58 $Y=2.79 $X2=0
+ $Y2=0
cc_461 N_A_119_368#_M1025_g N_VPWR_c_720_n 0.00533815f $X=2.485 $Y=2.4 $X2=0
+ $Y2=0
cc_462 N_A_119_368#_c_559_n N_VPWR_c_720_n 0.024929f $X=3.58 $Y=2.79 $X2=0 $Y2=0
cc_463 N_A_119_368#_M1027_g N_VPWR_c_721_n 0.00531893f $X=2.935 $Y=2.4 $X2=0
+ $Y2=0
cc_464 N_A_119_368#_c_559_n N_VPWR_c_721_n 0.024193f $X=3.58 $Y=2.79 $X2=0 $Y2=0
cc_465 N_A_119_368#_c_559_n N_Y_M1025_d 0.00405446f $X=3.58 $Y=2.79 $X2=0 $Y2=0
cc_466 N_A_119_368#_M1025_g N_Y_c_823_n 0.00475326f $X=2.485 $Y=2.4 $X2=0 $Y2=0
cc_467 N_A_119_368#_M1027_g N_Y_c_823_n 0.0117897f $X=2.935 $Y=2.4 $X2=0 $Y2=0
cc_468 N_A_119_368#_c_549_n N_Y_c_823_n 0.0145656f $X=4.01 $Y=2.625 $X2=0 $Y2=0
cc_469 N_A_119_368#_c_552_n N_Y_c_823_n 0.00793907f $X=3.935 $Y=2.79 $X2=0 $Y2=0
cc_470 N_A_119_368#_c_557_n N_Y_c_823_n 0.0113022f $X=4.425 $Y=2.79 $X2=0 $Y2=0
cc_471 N_A_119_368#_c_559_n N_Y_c_823_n 0.137372f $X=3.58 $Y=2.79 $X2=0 $Y2=0
cc_472 N_A_119_368#_M1014_g N_Y_c_884_n 0.0072257f $X=3.415 $Y=0.74 $X2=0 $Y2=0
cc_473 N_A_119_368#_M1017_g N_Y_c_884_n 8.09439e-19 $X=4.01 $Y=0.74 $X2=0 $Y2=0
cc_474 N_A_119_368#_M1014_g N_Y_c_818_n 0.00980971f $X=3.415 $Y=0.74 $X2=0 $Y2=0
cc_475 N_A_119_368#_M1017_g N_Y_c_818_n 0.00980971f $X=4.01 $Y=0.74 $X2=0 $Y2=0
cc_476 N_A_119_368#_c_540_n N_Y_c_818_n 0.00594145f $X=3.935 $Y=1.515 $X2=0
+ $Y2=0
cc_477 N_A_119_368#_c_544_n N_Y_c_818_n 0.0487586f $X=3.92 $Y=1.515 $X2=0 $Y2=0
cc_478 N_A_119_368#_M1010_g N_Y_c_819_n 0.00154617f $X=2.915 $Y=0.74 $X2=0 $Y2=0
cc_479 N_A_119_368#_M1014_g N_Y_c_819_n 0.00224059f $X=3.415 $Y=0.74 $X2=0 $Y2=0
cc_480 N_A_119_368#_c_542_n N_Y_c_819_n 0.00530643f $X=2.395 $Y=1.095 $X2=0
+ $Y2=0
cc_481 N_A_119_368#_c_544_n N_Y_c_819_n 0.0259696f $X=3.92 $Y=1.515 $X2=0 $Y2=0
cc_482 N_A_119_368#_c_546_n N_Y_c_819_n 0.00407434f $X=3.49 $Y=1.515 $X2=0 $Y2=0
cc_483 N_A_119_368#_M1014_g N_Y_c_832_n 8.15756e-19 $X=3.415 $Y=0.74 $X2=0 $Y2=0
cc_484 N_A_119_368#_M1017_g N_Y_c_832_n 0.00736932f $X=4.01 $Y=0.74 $X2=0 $Y2=0
cc_485 N_A_119_368#_M1029_g N_Y_c_832_n 0.0069444f $X=4.44 $Y=0.74 $X2=0 $Y2=0
cc_486 N_A_119_368#_M1029_g N_Y_c_820_n 0.00955794f $X=4.44 $Y=0.74 $X2=0 $Y2=0
cc_487 N_A_119_368#_M1017_g N_Y_c_822_n 0.00223114f $X=4.01 $Y=0.74 $X2=0 $Y2=0
cc_488 N_A_119_368#_c_538_n N_Y_c_822_n 0.00399889f $X=4.365 $Y=1.425 $X2=0
+ $Y2=0
cc_489 N_A_119_368#_M1029_g N_Y_c_822_n 0.00239941f $X=4.44 $Y=0.74 $X2=0 $Y2=0
cc_490 N_A_119_368#_c_544_n N_Y_c_822_n 0.00187548f $X=3.92 $Y=1.515 $X2=0 $Y2=0
cc_491 N_A_119_368#_c_556_n N_A_950_368#_c_948_n 0.0216952f $X=4.425 $Y=2.79
+ $X2=0 $Y2=0
cc_492 N_A_119_368#_c_557_n N_A_950_368#_c_948_n 0.00127602f $X=4.425 $Y=2.79
+ $X2=0 $Y2=0
cc_493 N_A_119_368#_c_545_n N_A_27_74#_c_1012_n 0.0129684f $X=1.71 $Y=0.86 $X2=0
+ $Y2=0
cc_494 N_A_119_368#_M1022_s N_A_27_74#_c_1015_n 0.00253871f $X=1.5 $Y=0.37 $X2=0
+ $Y2=0
cc_495 N_A_119_368#_M1010_g N_A_27_74#_c_1015_n 6.20634e-19 $X=2.915 $Y=0.74
+ $X2=0 $Y2=0
cc_496 N_A_119_368#_c_542_n N_A_27_74#_c_1015_n 0.0155485f $X=2.395 $Y=1.095
+ $X2=0 $Y2=0
cc_497 N_A_119_368#_c_545_n N_A_27_74#_c_1015_n 0.0200266f $X=1.71 $Y=0.86 $X2=0
+ $Y2=0
cc_498 N_A_119_368#_M1010_g N_VGND_c_1056_n 0.00278247f $X=2.915 $Y=0.74 $X2=0
+ $Y2=0
cc_499 N_A_119_368#_M1014_g N_VGND_c_1056_n 0.00278271f $X=3.415 $Y=0.74 $X2=0
+ $Y2=0
cc_500 N_A_119_368#_M1017_g N_VGND_c_1056_n 0.00278271f $X=4.01 $Y=0.74 $X2=0
+ $Y2=0
cc_501 N_A_119_368#_M1029_g N_VGND_c_1056_n 0.00278271f $X=4.44 $Y=0.74 $X2=0
+ $Y2=0
cc_502 N_A_119_368#_M1010_g N_VGND_c_1065_n 0.00359084f $X=2.915 $Y=0.74 $X2=0
+ $Y2=0
cc_503 N_A_119_368#_M1014_g N_VGND_c_1065_n 0.00355508f $X=3.415 $Y=0.74 $X2=0
+ $Y2=0
cc_504 N_A_119_368#_M1017_g N_VGND_c_1065_n 0.00354849f $X=4.01 $Y=0.74 $X2=0
+ $Y2=0
cc_505 N_A_119_368#_M1029_g N_VGND_c_1065_n 0.0035414f $X=4.44 $Y=0.74 $X2=0
+ $Y2=0
cc_506 N_A_119_368#_c_542_n N_A_511_74#_M1010_d 0.00155395f $X=2.395 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_507 N_A_119_368#_M1010_g N_A_511_74#_c_1168_n 0.00752841f $X=2.915 $Y=0.74
+ $X2=0 $Y2=0
cc_508 N_A_119_368#_M1014_g N_A_511_74#_c_1168_n 6.23275e-19 $X=3.415 $Y=0.74
+ $X2=0 $Y2=0
cc_509 N_A_119_368#_c_542_n N_A_511_74#_c_1168_n 0.00264903f $X=2.395 $Y=1.095
+ $X2=0 $Y2=0
cc_510 N_A_119_368#_c_544_n N_A_511_74#_c_1168_n 0.00919438f $X=3.92 $Y=1.515
+ $X2=0 $Y2=0
cc_511 N_A_119_368#_c_545_n N_A_511_74#_c_1168_n 0.00197495f $X=1.71 $Y=0.86
+ $X2=0 $Y2=0
cc_512 N_A_119_368#_c_546_n N_A_511_74#_c_1168_n 0.00543335f $X=3.49 $Y=1.515
+ $X2=0 $Y2=0
cc_513 N_A_119_368#_M1010_g N_A_511_74#_c_1169_n 0.0104643f $X=2.915 $Y=0.74
+ $X2=0 $Y2=0
cc_514 N_A_119_368#_M1014_g N_A_511_74#_c_1169_n 0.0120431f $X=3.415 $Y=0.74
+ $X2=0 $Y2=0
cc_515 N_A_119_368#_M1010_g N_A_511_74#_c_1170_n 0.00344571f $X=2.915 $Y=0.74
+ $X2=0 $Y2=0
cc_516 N_A_119_368#_M1017_g N_A_511_74#_c_1217_n 0.00719113f $X=4.01 $Y=0.74
+ $X2=0 $Y2=0
cc_517 N_A_119_368#_M1017_g N_A_511_74#_c_1171_n 0.0116499f $X=4.01 $Y=0.74
+ $X2=0 $Y2=0
cc_518 N_A_119_368#_M1029_g N_A_511_74#_c_1171_n 0.011161f $X=4.44 $Y=0.74 $X2=0
+ $Y2=0
cc_519 N_VPWR_M1027_s N_Y_c_823_n 0.00798432f $X=3.025 $Y=1.84 $X2=0 $Y2=0
cc_520 N_VPWR_M1000_s N_Y_c_823_n 0.00760622f $X=5.21 $Y=1.84 $X2=0 $Y2=0
cc_521 N_VPWR_M1006_s N_Y_c_823_n 0.00828316f $X=6.285 $Y=1.84 $X2=0 $Y2=0
cc_522 N_VPWR_M1006_s N_A_950_368#_c_952_n 0.0074523f $X=6.285 $Y=1.84 $X2=0
+ $Y2=0
cc_523 N_VPWR_c_717_n N_A_950_368#_c_952_n 0.00383176f $X=6.34 $Y=3.33 $X2=0
+ $Y2=0
cc_524 N_VPWR_c_718_n N_A_950_368#_c_952_n 0.00383985f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_525 N_VPWR_c_707_n N_A_950_368#_c_952_n 0.01304f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_526 N_VPWR_c_722_n N_A_950_368#_c_952_n 0.0241399f $X=6.505 $Y=3.05 $X2=0
+ $Y2=0
cc_527 N_VPWR_c_718_n N_A_950_368#_c_945_n 0.0459483f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_528 N_VPWR_c_707_n N_A_950_368#_c_945_n 0.0258042f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_529 N_VPWR_c_718_n N_A_950_368#_c_946_n 0.0638408f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_530 N_VPWR_c_707_n N_A_950_368#_c_946_n 0.0355196f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_531 N_VPWR_c_714_n N_A_950_368#_c_948_n 0.00101269f $X=5.43 $Y=3.05 $X2=0
+ $Y2=0
cc_532 N_VPWR_c_715_n N_A_950_368#_c_948_n 0.0104857f $X=5.265 $Y=3.33 $X2=0
+ $Y2=0
cc_533 N_VPWR_c_707_n N_A_950_368#_c_948_n 0.00882882f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_534 N_VPWR_M1000_s N_A_950_368#_c_956_n 0.00762332f $X=5.21 $Y=1.84 $X2=0
+ $Y2=0
cc_535 N_VPWR_c_714_n N_A_950_368#_c_956_n 0.0245079f $X=5.43 $Y=3.05 $X2=0
+ $Y2=0
cc_536 N_VPWR_c_715_n N_A_950_368#_c_956_n 0.00383985f $X=5.265 $Y=3.33 $X2=0
+ $Y2=0
cc_537 N_VPWR_c_717_n N_A_950_368#_c_956_n 0.00383176f $X=6.34 $Y=3.33 $X2=0
+ $Y2=0
cc_538 N_VPWR_c_707_n N_A_950_368#_c_956_n 0.0130673f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_539 N_VPWR_c_714_n N_A_950_368#_c_949_n 9.67958e-19 $X=5.43 $Y=3.05 $X2=0
+ $Y2=0
cc_540 N_VPWR_c_717_n N_A_950_368#_c_949_n 0.0138332f $X=6.34 $Y=3.33 $X2=0
+ $Y2=0
cc_541 N_VPWR_c_707_n N_A_950_368#_c_949_n 0.0116354f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_542 N_VPWR_c_722_n N_A_950_368#_c_949_n 9.66792e-19 $X=6.505 $Y=3.05 $X2=0
+ $Y2=0
cc_543 N_VPWR_c_718_n N_A_950_368#_c_950_n 0.0171415f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_544 N_VPWR_c_707_n N_A_950_368#_c_950_n 0.00940804f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_545 N_VPWR_c_722_n N_A_950_368#_c_950_n 0.00741728f $X=6.505 $Y=3.05 $X2=0
+ $Y2=0
cc_546 N_VPWR_c_718_n N_A_950_368#_c_951_n 0.0121867f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_547 N_VPWR_c_707_n N_A_950_368#_c_951_n 0.00660921f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_548 N_VPWR_c_709_n N_A_27_74#_c_1013_n 0.00886035f $X=0.28 $Y=1.985 $X2=0
+ $Y2=0
cc_549 N_Y_c_823_n N_A_950_368#_M1000_d 0.0072137f $X=7.325 $Y=2.37 $X2=-0.19
+ $Y2=-0.245
cc_550 N_Y_c_823_n N_A_950_368#_M1004_d 0.00332471f $X=7.325 $Y=2.37 $X2=0 $Y2=0
cc_551 N_Y_c_823_n N_A_950_368#_M1007_d 0.0045357f $X=7.325 $Y=2.37 $X2=0 $Y2=0
cc_552 N_Y_c_857_n N_A_950_368#_M1005_s 0.00313909f $X=8.225 $Y=2.02 $X2=0 $Y2=0
cc_553 N_Y_M1003_d N_A_950_368#_c_945_n 0.00165831f $X=7.355 $Y=1.84 $X2=0 $Y2=0
cc_554 N_Y_c_823_n N_A_950_368#_c_945_n 0.0206639f $X=7.325 $Y=2.37 $X2=0 $Y2=0
cc_555 N_Y_c_857_n N_A_950_368#_c_1005_n 0.0126919f $X=8.225 $Y=2.02 $X2=0 $Y2=0
cc_556 N_Y_M1008_d N_A_950_368#_c_946_n 0.00165831f $X=8.255 $Y=1.84 $X2=0 $Y2=0
cc_557 N_Y_c_867_n N_A_950_368#_c_946_n 0.0159318f $X=8.39 $Y=2.1 $X2=0 $Y2=0
cc_558 N_Y_c_823_n N_A_950_368#_c_948_n 0.0145678f $X=7.325 $Y=2.37 $X2=0 $Y2=0
cc_559 N_Y_c_823_n N_A_950_368#_c_956_n 0.104545f $X=7.325 $Y=2.37 $X2=0 $Y2=0
cc_560 N_Y_c_823_n N_A_950_368#_c_950_n 0.0143712f $X=7.325 $Y=2.37 $X2=0 $Y2=0
cc_561 N_Y_c_820_n N_VGND_M1002_s 0.00391227f $X=8.325 $Y=1.095 $X2=0 $Y2=0
cc_562 N_Y_c_820_n N_VGND_M1021_s 0.00391227f $X=8.325 $Y=1.095 $X2=0 $Y2=0
cc_563 N_Y_c_820_n N_VGND_M1001_d 0.00447702f $X=8.325 $Y=1.095 $X2=0 $Y2=0
cc_564 N_Y_c_820_n N_VGND_M1016_d 0.00459163f $X=8.325 $Y=1.095 $X2=0 $Y2=0
cc_565 N_Y_c_818_n N_A_511_74#_M1014_d 0.00409088f $X=4.06 $Y=1.095 $X2=0 $Y2=0
cc_566 N_Y_c_820_n N_A_511_74#_M1029_d 0.00250873f $X=8.325 $Y=1.095 $X2=0 $Y2=0
cc_567 N_Y_c_820_n N_A_511_74#_M1009_d 0.00176461f $X=8.325 $Y=1.095 $X2=0 $Y2=0
cc_568 N_Y_c_820_n N_A_511_74#_M1023_d 0.00176461f $X=8.325 $Y=1.095 $X2=0 $Y2=0
cc_569 N_Y_c_820_n N_A_511_74#_M1015_s 0.00176461f $X=8.325 $Y=1.095 $X2=0 $Y2=0
cc_570 N_Y_M1010_s N_A_511_74#_c_1169_n 0.00250873f $X=2.99 $Y=0.37 $X2=0 $Y2=0
cc_571 N_Y_c_884_n N_A_511_74#_c_1169_n 0.019446f $X=3.2 $Y=0.86 $X2=0 $Y2=0
cc_572 N_Y_c_818_n N_A_511_74#_c_1169_n 0.00304353f $X=4.06 $Y=1.095 $X2=0 $Y2=0
cc_573 N_Y_c_818_n N_A_511_74#_c_1217_n 0.0254766f $X=4.06 $Y=1.095 $X2=0 $Y2=0
cc_574 N_Y_c_832_n N_A_511_74#_c_1217_n 0.0171106f $X=4.225 $Y=0.86 $X2=0 $Y2=0
cc_575 N_Y_M1017_s N_A_511_74#_c_1171_n 0.00176461f $X=4.085 $Y=0.37 $X2=0 $Y2=0
cc_576 N_Y_c_818_n N_A_511_74#_c_1171_n 0.0034045f $X=4.06 $Y=1.095 $X2=0 $Y2=0
cc_577 N_Y_c_832_n N_A_511_74#_c_1171_n 0.0158692f $X=4.225 $Y=0.86 $X2=0 $Y2=0
cc_578 N_Y_c_820_n N_A_511_74#_c_1171_n 0.00304353f $X=8.325 $Y=1.095 $X2=0
+ $Y2=0
cc_579 N_Y_c_820_n N_A_511_74#_c_1180_n 0.0405897f $X=8.325 $Y=1.095 $X2=0 $Y2=0
cc_580 N_Y_c_820_n N_A_511_74#_c_1182_n 0.0208474f $X=8.325 $Y=1.095 $X2=0 $Y2=0
cc_581 N_Y_c_820_n N_A_511_74#_c_1183_n 0.0406235f $X=8.325 $Y=1.095 $X2=0 $Y2=0
cc_582 N_Y_c_820_n N_A_511_74#_c_1193_n 0.0431657f $X=8.325 $Y=1.095 $X2=0 $Y2=0
cc_583 N_Y_c_820_n N_A_511_74#_c_1195_n 0.0335805f $X=8.325 $Y=1.095 $X2=0 $Y2=0
cc_584 N_Y_c_820_n N_A_511_74#_c_1173_n 0.0167101f $X=8.325 $Y=1.095 $X2=0 $Y2=0
cc_585 N_Y_c_820_n N_A_511_74#_c_1174_n 0.0167101f $X=8.325 $Y=1.095 $X2=0 $Y2=0
cc_586 N_Y_c_820_n N_A_511_74#_c_1175_n 0.0167101f $X=8.325 $Y=1.095 $X2=0 $Y2=0
cc_587 N_Y_c_820_n N_A_511_74#_c_1176_n 0.00517071f $X=8.325 $Y=1.095 $X2=0
+ $Y2=0
cc_588 N_A_27_74#_c_1012_n N_VGND_M1019_s 0.00250873f $X=1.045 $Y=1.065
+ $X2=-0.19 $Y2=-0.245
cc_589 N_A_27_74#_c_1011_n N_VGND_c_1051_n 0.017215f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_590 N_A_27_74#_c_1012_n N_VGND_c_1051_n 0.0210288f $X=1.045 $Y=1.065 $X2=0
+ $Y2=0
cc_591 N_A_27_74#_c_1014_n N_VGND_c_1051_n 0.0113248f $X=1.21 $Y=0.6 $X2=0 $Y2=0
cc_592 N_A_27_74#_c_1014_n N_VGND_c_1056_n 0.0145754f $X=1.21 $Y=0.6 $X2=0 $Y2=0
cc_593 N_A_27_74#_c_1015_n N_VGND_c_1056_n 0.0377744f $X=2.14 $Y=0.515 $X2=0
+ $Y2=0
cc_594 N_A_27_74#_c_1011_n N_VGND_c_1062_n 0.011066f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_595 N_A_27_74#_c_1011_n N_VGND_c_1065_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_596 N_A_27_74#_c_1014_n N_VGND_c_1065_n 0.0119468f $X=1.21 $Y=0.6 $X2=0 $Y2=0
cc_597 N_A_27_74#_c_1015_n N_VGND_c_1065_n 0.031928f $X=2.14 $Y=0.515 $X2=0
+ $Y2=0
cc_598 N_A_27_74#_c_1015_n N_A_511_74#_c_1168_n 0.012414f $X=2.14 $Y=0.515 $X2=0
+ $Y2=0
cc_599 N_A_27_74#_c_1015_n N_A_511_74#_c_1170_n 0.00560069f $X=2.14 $Y=0.515
+ $X2=0 $Y2=0
cc_600 N_VGND_c_1056_n N_A_511_74#_c_1169_n 0.0423044f $X=5.07 $Y=0 $X2=0 $Y2=0
cc_601 N_VGND_c_1065_n N_A_511_74#_c_1169_n 0.0239316f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_602 N_VGND_c_1056_n N_A_511_74#_c_1170_n 0.0233048f $X=5.07 $Y=0 $X2=0 $Y2=0
cc_603 N_VGND_c_1065_n N_A_511_74#_c_1170_n 0.0126653f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_604 N_VGND_c_1052_n N_A_511_74#_c_1171_n 0.0114117f $X=5.235 $Y=0.335 $X2=0
+ $Y2=0
cc_605 N_VGND_c_1056_n N_A_511_74#_c_1171_n 0.0671424f $X=5.07 $Y=0 $X2=0 $Y2=0
cc_606 N_VGND_c_1065_n N_A_511_74#_c_1171_n 0.0374222f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_607 N_VGND_M1002_s N_A_511_74#_c_1180_n 0.00726893f $X=5.015 $Y=0.37 $X2=0
+ $Y2=0
cc_608 N_VGND_c_1052_n N_A_511_74#_c_1180_n 0.0251188f $X=5.235 $Y=0.335 $X2=0
+ $Y2=0
cc_609 N_VGND_c_1056_n N_A_511_74#_c_1180_n 0.00236055f $X=5.07 $Y=0 $X2=0 $Y2=0
cc_610 N_VGND_c_1058_n N_A_511_74#_c_1180_n 0.0023667f $X=6.09 $Y=0 $X2=0 $Y2=0
cc_611 N_VGND_c_1065_n N_A_511_74#_c_1180_n 0.0102151f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_612 N_VGND_M1021_s N_A_511_74#_c_1183_n 0.00732248f $X=6.035 $Y=0.37 $X2=0
+ $Y2=0
cc_613 N_VGND_c_1053_n N_A_511_74#_c_1183_n 0.0251188f $X=6.255 $Y=0.335 $X2=0
+ $Y2=0
cc_614 N_VGND_c_1058_n N_A_511_74#_c_1183_n 0.0023667f $X=6.09 $Y=0 $X2=0 $Y2=0
cc_615 N_VGND_c_1060_n N_A_511_74#_c_1183_n 0.0023667f $X=7.11 $Y=0 $X2=0 $Y2=0
cc_616 N_VGND_c_1065_n N_A_511_74#_c_1183_n 0.0102196f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_617 N_VGND_M1001_d N_A_511_74#_c_1193_n 0.00811089f $X=7.055 $Y=0.37 $X2=0
+ $Y2=0
cc_618 N_VGND_c_1054_n N_A_511_74#_c_1193_n 0.0278156f $X=7.29 $Y=0.335 $X2=0
+ $Y2=0
cc_619 N_VGND_c_1060_n N_A_511_74#_c_1193_n 0.0023667f $X=7.11 $Y=0 $X2=0 $Y2=0
cc_620 N_VGND_c_1063_n N_A_511_74#_c_1193_n 0.0023667f $X=8.165 $Y=0 $X2=0 $Y2=0
cc_621 N_VGND_c_1065_n N_A_511_74#_c_1193_n 0.0103668f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_622 N_VGND_M1016_d N_A_511_74#_c_1195_n 0.00725567f $X=8.11 $Y=0.37 $X2=0
+ $Y2=0
cc_623 N_VGND_c_1055_n N_A_511_74#_c_1195_n 0.0251188f $X=8.33 $Y=0.335 $X2=0
+ $Y2=0
cc_624 N_VGND_c_1063_n N_A_511_74#_c_1195_n 0.0023667f $X=8.165 $Y=0 $X2=0 $Y2=0
cc_625 N_VGND_c_1064_n N_A_511_74#_c_1195_n 0.0023667f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_626 N_VGND_c_1065_n N_A_511_74#_c_1195_n 0.0102196f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_627 N_VGND_c_1056_n N_A_511_74#_c_1172_n 0.023391f $X=5.07 $Y=0 $X2=0 $Y2=0
cc_628 N_VGND_c_1065_n N_A_511_74#_c_1172_n 0.0127797f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_629 N_VGND_c_1052_n N_A_511_74#_c_1173_n 0.00613542f $X=5.235 $Y=0.335 $X2=0
+ $Y2=0
cc_630 N_VGND_c_1053_n N_A_511_74#_c_1173_n 0.00613542f $X=6.255 $Y=0.335 $X2=0
+ $Y2=0
cc_631 N_VGND_c_1058_n N_A_511_74#_c_1173_n 0.0141563f $X=6.09 $Y=0 $X2=0 $Y2=0
cc_632 N_VGND_c_1065_n N_A_511_74#_c_1173_n 0.0117515f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_633 N_VGND_c_1053_n N_A_511_74#_c_1174_n 0.00613542f $X=6.255 $Y=0.335 $X2=0
+ $Y2=0
cc_634 N_VGND_c_1054_n N_A_511_74#_c_1174_n 0.00614709f $X=7.29 $Y=0.335 $X2=0
+ $Y2=0
cc_635 N_VGND_c_1060_n N_A_511_74#_c_1174_n 0.0141563f $X=7.11 $Y=0 $X2=0 $Y2=0
cc_636 N_VGND_c_1065_n N_A_511_74#_c_1174_n 0.0117515f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_637 N_VGND_c_1054_n N_A_511_74#_c_1175_n 0.00614709f $X=7.29 $Y=0.335 $X2=0
+ $Y2=0
cc_638 N_VGND_c_1055_n N_A_511_74#_c_1175_n 0.00613542f $X=8.33 $Y=0.335 $X2=0
+ $Y2=0
cc_639 N_VGND_c_1063_n N_A_511_74#_c_1175_n 0.0141563f $X=8.165 $Y=0 $X2=0 $Y2=0
cc_640 N_VGND_c_1065_n N_A_511_74#_c_1175_n 0.0117515f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_641 N_VGND_c_1055_n N_A_511_74#_c_1176_n 0.00613542f $X=8.33 $Y=0.335 $X2=0
+ $Y2=0
cc_642 N_VGND_c_1064_n N_A_511_74#_c_1176_n 0.0145639f $X=8.88 $Y=0 $X2=0 $Y2=0
cc_643 N_VGND_c_1065_n N_A_511_74#_c_1176_n 0.0119984f $X=8.88 $Y=0 $X2=0 $Y2=0

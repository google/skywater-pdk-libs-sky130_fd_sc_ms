* File: sky130_fd_sc_ms__dlxtp_1.pex.spice
* Created: Fri Aug 28 17:30:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLXTP_1%D 3 7 11 12 13 14 18
r30 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.43
+ $Y=1.345 $X2=0.43 $Y2=1.345
r31 14 19 8.14351 $w=4.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.36 $Y=1.665
+ $X2=0.36 $Y2=1.345
r32 13 19 1.27242 $w=4.68e-07 $l=5e-08 $layer=LI1_cond $X=0.36 $Y=1.295 $X2=0.36
+ $Y2=1.345
r33 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.43 $Y=1.685
+ $X2=0.43 $Y2=1.345
r34 11 12 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.43 $Y=1.685
+ $X2=0.43 $Y2=1.85
r35 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.43 $Y=1.18
+ $X2=0.43 $Y2=1.345
r36 7 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.52 $Y=0.715
+ $X2=0.52 $Y2=1.18
r37 3 12 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=0.505 $Y=2.54
+ $X2=0.505 $Y2=1.85
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTP_1%A_119_88# 1 2 9 13 15 17 18 21 23 25 27 28
+ 33 34 35
r69 34 35 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.86 $Y=2.1 $X2=0.86
+ $Y2=1.77
r70 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1 $Y=1.265
+ $X2=1 $Y2=1.265
r71 28 35 9.49412 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=0.97 $Y=1.575
+ $X2=0.97 $Y2=1.77
r72 27 32 1.32389 $w=3.9e-07 $l=9.38083e-08 $layer=LI1_cond $X=0.97 $Y=1.295
+ $X2=0.89 $Y2=1.265
r73 27 28 8.27395 $w=3.88e-07 $l=2.8e-07 $layer=LI1_cond $X=0.97 $Y=1.295
+ $X2=0.97 $Y2=1.575
r74 23 34 7.90841 $w=2.98e-07 $l=1.5e-07 $layer=LI1_cond $X=0.795 $Y=2.25
+ $X2=0.795 $Y2=2.1
r75 23 25 0.576222 $w=2.98e-07 $l=1.5e-08 $layer=LI1_cond $X=0.795 $Y=2.25
+ $X2=0.795 $Y2=2.265
r76 19 32 15.5273 $w=3.3e-07 $l=4.71805e-07 $layer=LI1_cond $X=0.78 $Y=0.845
+ $X2=0.89 $Y2=1.265
r77 19 21 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.78 $Y=0.845
+ $X2=0.78 $Y2=0.715
r78 15 18 18.8402 $w=1.65e-07 $l=9.68246e-08 $layer=POLY_cond $X=1.6 $Y=1.24
+ $X2=1.55 $Y2=1.315
r79 15 17 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.6 $Y=1.24 $X2=1.6
+ $Y2=0.795
r80 11 18 18.8402 $w=1.65e-07 $l=9.08295e-08 $layer=POLY_cond $X=1.515 $Y=1.39
+ $X2=1.55 $Y2=1.315
r81 11 13 415.919 $w=1.8e-07 $l=1.07e-06 $layer=POLY_cond $X=1.515 $Y=1.39
+ $X2=1.515 $Y2=2.46
r82 10 33 19.8992 $w=1.5e-07 $l=1.96914e-07 $layer=POLY_cond $X=1.165 $Y=1.315
+ $X2=1 $Y2=1.245
r83 9 18 6.66866 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=1.425 $Y=1.315
+ $X2=1.55 $Y2=1.315
r84 9 10 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.425 $Y=1.315
+ $X2=1.165 $Y2=1.315
r85 2 25 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=2.12 $X2=0.73 $Y2=2.265
r86 1 21 182 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.44 $X2=0.78 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTP_1%A_386_326# 1 2 9 11 12 16 19 23 25 30 32 33
+ 36 37 46 48 52 53 57
c142 46 0 2.34272e-19 $X=4.69 $Y=1.83
c143 25 0 1.23079e-19 $X=4.565 $Y=0.34
r144 53 61 40.6969 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=7.092 $Y=1.485
+ $X2=7.092 $Y2=1.65
r145 53 60 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=7.092 $Y=1.485
+ $X2=7.092 $Y2=1.32
r146 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.09
+ $Y=1.485 $X2=7.09 $Y2=1.485
r147 49 52 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=6.98 $Y=1.485
+ $X2=7.09 $Y2=1.485
r148 44 46 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=4.45 $Y=1.83
+ $X2=4.69 $Y2=1.83
r149 41 57 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=2.34 $Y=0.42
+ $X2=2.495 $Y2=0.42
r150 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.34
+ $Y=0.42 $X2=2.34 $Y2=0.42
r151 37 40 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.34 $Y=0.34 $X2=2.34
+ $Y2=0.42
r152 36 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.98 $Y=1.32
+ $X2=6.98 $Y2=1.485
r153 35 36 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=6.98 $Y=0.75
+ $X2=6.98 $Y2=1.32
r154 34 48 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.815 $Y=0.665
+ $X2=4.69 $Y2=0.665
r155 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.895 $Y=0.665
+ $X2=6.98 $Y2=0.75
r156 33 34 135.701 $w=1.68e-07 $l=2.08e-06 $layer=LI1_cond $X=6.895 $Y=0.665
+ $X2=4.815 $Y2=0.665
r157 32 46 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=4.69 $Y=1.665
+ $X2=4.69 $Y2=1.83
r158 31 48 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.69 $Y=0.75
+ $X2=4.69 $Y2=0.665
r159 31 32 42.1794 $w=2.48e-07 $l=9.15e-07 $layer=LI1_cond $X=4.69 $Y=0.75
+ $X2=4.69 $Y2=1.665
r160 28 48 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.69 $Y=0.58
+ $X2=4.69 $Y2=0.665
r161 28 30 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=4.69 $Y=0.58
+ $X2=4.69 $Y2=0.555
r162 27 30 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=4.69 $Y=0.425
+ $X2=4.69 $Y2=0.555
r163 26 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=0.34
+ $X2=2.34 $Y2=0.34
r164 25 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.565 $Y=0.34
+ $X2=4.69 $Y2=0.425
r165 25 26 134.396 $w=1.68e-07 $l=2.06e-06 $layer=LI1_cond $X=4.565 $Y=0.34
+ $X2=2.505 $Y2=0.34
r166 23 60 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=7.185 $Y=0.78
+ $X2=7.185 $Y2=1.32
r167 19 61 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=7.17 $Y=2.4
+ $X2=7.17 $Y2=1.65
r168 14 16 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.495 $Y=1.63
+ $X2=2.495 $Y2=0.955
r169 13 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.495 $Y=0.585
+ $X2=2.495 $Y2=0.42
r170 13 16 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.495 $Y=0.585
+ $X2=2.495 $Y2=0.955
r171 11 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.42 $Y=1.705
+ $X2=2.495 $Y2=1.63
r172 11 12 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=2.42 $Y=1.705
+ $X2=2.11 $Y2=1.705
r173 7 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.02 $Y=1.78
+ $X2=2.11 $Y2=1.705
r174 7 9 151.597 $w=1.8e-07 $l=3.9e-07 $layer=POLY_cond $X=2.02 $Y=1.78 $X2=2.02
+ $Y2=2.17
r175 2 44 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=4.29
+ $Y=1.685 $X2=4.45 $Y2=1.83
r176 1 30 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.505
+ $Y=0.41 $X2=4.65 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTP_1%A_562_123# 1 2 9 13 17 21 23 24 28 29 31 32
+ 33 35 37 43 44 47 51 56
c134 43 0 1.01851e-19 $X=3.02 $Y=1.6
c135 21 0 9.26936e-20 $X=5.455 $Y=0.78
c136 17 0 7.64129e-20 $X=5.315 $Y=2.105
c137 9 0 1.72744e-19 $X=2.885 $Y=0.955
r138 48 51 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=6.09 $Y=1.045
+ $X2=6.235 $Y2=1.045
r139 44 46 8.32359 $w=5.13e-07 $l=3.5e-07 $layer=LI1_cond $X=6.01 $Y=2.325
+ $X2=6.36 $Y2=2.325
r140 43 55 39.5669 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=2.997 $Y=1.6
+ $X2=2.997 $Y2=1.765
r141 43 54 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=2.997 $Y=1.6
+ $X2=2.997 $Y2=1.435
r142 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.02
+ $Y=1.6 $X2=3.02 $Y2=1.6
r143 39 48 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.09 $Y=1.17
+ $X2=6.09 $Y2=1.045
r144 39 47 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.09 $Y=1.17
+ $X2=6.09 $Y2=1.35
r145 38 56 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.01 $Y=1.515
+ $X2=6.01 $Y2=1.425
r146 37 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.01 $Y=1.515
+ $X2=6.01 $Y2=1.35
r147 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.01
+ $Y=1.515 $X2=6.01 $Y2=1.515
r148 35 44 3.31882 $w=3.3e-07 $l=3.75e-07 $layer=LI1_cond $X=6.01 $Y=1.95
+ $X2=6.01 $Y2=2.325
r149 35 37 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=6.01 $Y=1.95
+ $X2=6.01 $Y2=1.515
r150 32 44 21.7992 $w=5.13e-07 $l=7.91486e-07 $layer=LI1_cond $X=5.34 $Y=2.59
+ $X2=6.01 $Y2=2.325
r151 32 33 103.08 $w=1.68e-07 $l=1.58e-06 $layer=LI1_cond $X=5.34 $Y=2.59
+ $X2=3.76 $Y2=2.59
r152 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.675 $Y=2.505
+ $X2=3.76 $Y2=2.59
r153 30 31 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.675 $Y=1.885
+ $X2=3.675 $Y2=2.505
r154 29 42 14.6448 $w=3.7e-07 $l=3.98905e-07 $layer=LI1_cond $X=3.355 $Y=1.8
+ $X2=3.02 $Y2=1.66
r155 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.59 $Y=1.8
+ $X2=3.675 $Y2=1.885
r156 28 29 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.59 $Y=1.8
+ $X2=3.355 $Y2=1.8
r157 24 27 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.53 $Y=1.425
+ $X2=5.455 $Y2=1.425
r158 23 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.845 $Y=1.425
+ $X2=6.01 $Y2=1.425
r159 23 24 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=5.845 $Y=1.425
+ $X2=5.53 $Y2=1.425
r160 19 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.455 $Y=1.35
+ $X2=5.455 $Y2=1.425
r161 19 21 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=5.455 $Y=1.35
+ $X2=5.455 $Y2=0.78
r162 15 27 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=5.315 $Y=1.425
+ $X2=5.455 $Y2=1.425
r163 15 17 235.169 $w=1.8e-07 $l=6.05e-07 $layer=POLY_cond $X=5.315 $Y=1.5
+ $X2=5.315 $Y2=2.105
r164 13 55 270.153 $w=1.8e-07 $l=6.95e-07 $layer=POLY_cond $X=3.03 $Y=2.46
+ $X2=3.03 $Y2=1.765
r165 9 54 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.885 $Y=0.955
+ $X2=2.885 $Y2=1.435
r166 2 46 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=6.215
+ $Y=1.84 $X2=6.36 $Y2=2.115
r167 1 51 182 $w=1.7e-07 $l=6.65789e-07 $layer=licon1_NDIFF $count=1 $X=6.085
+ $Y=0.41 $X2=6.235 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTP_1%A_685_59# 1 2 9 12 15 16 19 20 23 26 27 28
+ 32 36
c87 32 0 9.36104e-20 $X=5.54 $Y=1.83
c88 20 0 1.01851e-19 $X=3.93 $Y=1.41
c89 19 0 8.54063e-20 $X=3.665 $Y=1.78
c90 12 0 1.15446e-19 $X=3.565 $Y=2.75
r91 33 36 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=5.5 $Y=1.045
+ $X2=5.67 $Y2=1.045
r92 30 32 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.5 $Y=2.165
+ $X2=5.5 $Y2=1.83
r93 29 33 0.716491 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=5.5 $Y=1.17 $X2=5.5
+ $Y2=1.045
r94 29 32 30.4245 $w=2.48e-07 $l=6.6e-07 $layer=LI1_cond $X=5.5 $Y=1.17 $X2=5.5
+ $Y2=1.83
r95 27 30 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.375 $Y=2.25
+ $X2=5.5 $Y2=2.165
r96 27 28 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=5.375 $Y=2.25
+ $X2=4.1 $Y2=2.25
r97 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.015 $Y=2.165
+ $X2=4.1 $Y2=2.25
r98 25 26 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.015 $Y=1.545
+ $X2=4.015 $Y2=2.165
r99 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.69
+ $Y=1.44 $X2=3.69 $Y2=1.44
r100 20 25 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=3.93 $Y=1.41
+ $X2=4.015 $Y2=1.545
r101 20 22 10.2439 $w=2.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.93 $Y=1.41
+ $X2=3.69 $Y2=1.41
r102 18 23 31.3252 $w=3.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.68 $Y=1.63
+ $X2=3.68 $Y2=1.44
r103 18 19 38.2996 $w=3.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.665 $Y=1.63
+ $X2=3.665 $Y2=1.78
r104 16 23 8.24346 $w=3.5e-07 $l=5e-08 $layer=POLY_cond $X=3.68 $Y=1.39 $X2=3.68
+ $Y2=1.44
r105 15 16 43.9584 $w=3.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.64 $Y=1.24
+ $X2=3.64 $Y2=1.39
r106 12 19 377.048 $w=1.8e-07 $l=9.7e-07 $layer=POLY_cond $X=3.565 $Y=2.75
+ $X2=3.565 $Y2=1.78
r107 9 15 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.5 $Y=0.795
+ $X2=3.5 $Y2=1.24
r108 2 32 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=5.405
+ $Y=1.685 $X2=5.54 $Y2=1.83
r109 1 36 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=5.53
+ $Y=0.41 $X2=5.67 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTP_1%A_592_149# 1 2 7 8 11 13 15 18 21 23 24 26
+ 28 33 34 36 37
c103 28 0 8.54063e-20 $X=4.065 $Y=1.02
c104 24 0 3.11805e-20 $X=3.015 $Y=2.14
c105 23 0 3.03849e-20 $X=2.685 $Y=1.18
c106 18 0 1.92762e-19 $X=4.865 $Y=1.3
c107 7 0 1.3512e-19 $X=4.605 $Y=1.3
r108 36 39 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.23 $Y=0.94 $X2=4.23
+ $Y2=1.02
r109 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.23
+ $Y=0.94 $X2=4.23 $Y2=0.94
r110 32 34 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.185 $Y=1.1
+ $X2=3.355 $Y2=1.1
r111 32 33 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.185 $Y=1.1
+ $X2=3.015 $Y2=1.1
r112 28 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.065 $Y=1.02
+ $X2=4.23 $Y2=1.02
r113 28 34 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.065 $Y=1.02
+ $X2=3.355 $Y2=1.02
r114 24 30 24.5879 $w=2.1e-07 $l=4.43988e-07 $layer=LI1_cond $X=3.015 $Y=2.14
+ $X2=2.6 $Y2=2.08
r115 24 26 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.015 $Y=2.14
+ $X2=3.255 $Y2=2.14
r116 23 33 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.685 $Y=1.18
+ $X2=3.015 $Y2=1.18
r117 21 30 1.9771 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.6 $Y=1.935 $X2=2.6
+ $Y2=2.08
r118 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.6 $Y=1.265
+ $X2=2.685 $Y2=1.18
r119 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.6 $Y=1.265
+ $X2=2.6 $Y2=1.935
r120 16 37 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=4.23 $Y=1.225
+ $X2=4.23 $Y2=0.94
r121 13 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.865 $Y=1.225
+ $X2=4.865 $Y2=1.3
r122 13 15 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.865 $Y=1.225
+ $X2=4.865 $Y2=0.78
r123 9 18 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.695 $Y=1.3
+ $X2=4.865 $Y2=1.3
r124 9 11 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=4.695 $Y=1.375
+ $X2=4.695 $Y2=2.245
r125 8 16 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.395 $Y=1.3
+ $X2=4.23 $Y2=1.225
r126 7 9 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.605 $Y=1.3 $X2=4.695
+ $Y2=1.3
r127 7 8 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.605 $Y=1.3
+ $X2=4.395 $Y2=1.3
r128 2 26 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=3.12
+ $Y=1.96 $X2=3.255 $Y2=2.14
r129 1 32 182 $w=1.7e-07 $l=3.7081e-07 $layer=licon1_NDIFF $count=1 $X=2.96
+ $Y=0.745 $X2=3.185 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTP_1%GATE 3 7 9 12 13
r38 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.55 $Y=1.515
+ $X2=6.55 $Y2=1.68
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.55 $Y=1.515
+ $X2=6.55 $Y2=1.35
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.55
+ $Y=1.515 $X2=6.55 $Y2=1.515
r41 9 13 4.93904 $w=3.48e-07 $l=1.5e-07 $layer=LI1_cond $X=6.54 $Y=1.665
+ $X2=6.54 $Y2=1.515
r42 7 15 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=6.585 $Y=2.26
+ $X2=6.585 $Y2=1.68
r43 3 14 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=6.46 $Y=0.78 $X2=6.46
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTP_1%VPWR 1 2 3 4 13 15 19 23 25 27 32 40 50 51
+ 57 64 67
r68 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r69 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r70 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r71 51 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r72 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r73 48 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.06 $Y=3.33
+ $X2=6.895 $Y2=3.33
r74 48 50 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=7.06 $Y=3.33
+ $X2=7.44 $Y2=3.33
r75 47 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r76 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r77 44 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r78 44 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r79 43 46 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.52 $Y=3.33 $X2=6.48
+ $Y2=3.33
r80 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r81 41 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.17 $Y=3.33
+ $X2=5.005 $Y2=3.33
r82 41 43 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5.17 $Y=3.33
+ $X2=5.52 $Y2=3.33
r83 40 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.73 $Y=3.33
+ $X2=6.895 $Y2=3.33
r84 40 46 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.73 $Y=3.33
+ $X2=6.48 $Y2=3.33
r85 39 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r86 38 39 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r87 36 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r88 35 38 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=4.56 $Y2=3.33
r89 35 36 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r90 33 35 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=2.16 $Y2=3.33
r91 32 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.84 $Y=3.33
+ $X2=5.005 $Y2=3.33
r92 32 38 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.84 $Y=3.33
+ $X2=4.56 $Y2=3.33
r93 31 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r94 31 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r95 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r96 28 54 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r97 28 30 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r98 27 33 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=1.827 $Y=3.33
+ $X2=1.995 $Y2=3.33
r99 27 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r100 27 57 9.97637 $w=3.33e-07 $l=2.9e-07 $layer=LI1_cond $X=1.827 $Y=3.33
+ $X2=1.827 $Y2=3.04
r101 27 30 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.66 $Y=3.33
+ $X2=0.72 $Y2=3.33
r102 25 39 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.56 $Y2=3.33
r103 25 36 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=2.16 $Y2=3.33
r104 21 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.895 $Y=3.245
+ $X2=6.895 $Y2=3.33
r105 21 23 39.4624 $w=3.28e-07 $l=1.13e-06 $layer=LI1_cond $X=6.895 $Y=3.245
+ $X2=6.895 $Y2=2.115
r106 17 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=3.245
+ $X2=5.005 $Y2=3.33
r107 17 19 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=5.005 $Y=3.245
+ $X2=5.005 $Y2=3.01
r108 13 54 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r109 13 15 34.2241 $w=3.28e-07 $l=9.8e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.265
r110 4 23 300 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_PDIFF $count=2 $X=6.675
+ $Y=1.84 $X2=6.895 $Y2=2.115
r111 3 19 600 $w=1.7e-07 $l=1.43078e-06 $layer=licon1_PDIFF $count=1 $X=4.785
+ $Y=1.685 $X2=5.005 $Y2=3.01
r112 2 57 600 $w=1.7e-07 $l=1.18491e-06 $layer=licon1_PDIFF $count=1 $X=1.605
+ $Y=1.96 $X2=1.825 $Y2=3.04
r113 1 15 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.265
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTP_1%A_229_392# 1 2 9 15 17 21 22
c41 15 0 1.46626e-19 $X=2.805 $Y=2.82
r42 21 22 9.02376 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=2.165 $Y=2.8
+ $X2=2.335 $Y2=2.8
r43 17 19 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.29 $Y=2.7
+ $X2=1.29 $Y2=2.815
r44 15 22 21.6659 $w=2.48e-07 $l=4.7e-07 $layer=LI1_cond $X=2.805 $Y=2.86
+ $X2=2.335 $Y2=2.86
r45 12 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=2.7
+ $X2=1.29 $Y2=2.7
r46 12 21 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.455 $Y=2.7
+ $X2=2.165 $Y2=2.7
r47 7 17 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.29 $Y=2.615
+ $X2=1.29 $Y2=2.7
r48 7 9 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=1.29 $Y=2.615 $X2=1.29
+ $Y2=2.105
r49 2 15 600 $w=1.7e-07 $l=9.29677e-07 $layer=licon1_PDIFF $count=1 $X=2.66
+ $Y=1.96 $X2=2.805 $Y2=2.82
r50 1 19 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.96 $X2=1.29 $Y2=2.815
r51 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.96 $X2=1.29 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTP_1%A_422_392# 1 2 9 11 12 13 16 17 19 21
r54 21 23 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.59 $Y=2.36
+ $X2=2.59 $Y2=2.48
r55 17 19 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.31 $Y=2.93
+ $X2=3.875 $Y2=2.93
r56 16 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.225 $Y=2.845
+ $X2=3.31 $Y2=2.93
r57 15 16 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.225 $Y=2.565
+ $X2=3.225 $Y2=2.845
r58 14 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.675 $Y=2.48
+ $X2=2.59 $Y2=2.48
r59 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.14 $Y=2.48
+ $X2=3.225 $Y2=2.565
r60 13 14 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.14 $Y=2.48
+ $X2=2.675 $Y2=2.48
r61 11 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=2.36
+ $X2=2.59 $Y2=2.36
r62 11 12 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.505 $Y=2.36
+ $X2=2.33 $Y2=2.36
r63 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.205 $Y=2.275
+ $X2=2.33 $Y2=2.36
r64 7 9 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=2.205 $Y=2.275
+ $X2=2.205 $Y2=2.17
r65 2 19 600 $w=1.7e-07 $l=4.8775e-07 $layer=licon1_PDIFF $count=1 $X=3.655
+ $Y=2.54 $X2=3.875 $Y2=2.93
r66 1 9 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=2.11
+ $Y=1.96 $X2=2.245 $Y2=2.17
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTP_1%Q 1 2 9 13 14 15 16 23 32
r22 21 23 1.04193 $w=3.63e-07 $l=3.3e-08 $layer=LI1_cond $X=7.412 $Y=2.002
+ $X2=7.412 $Y2=2.035
r23 15 16 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=7.412 $Y=2.405
+ $X2=7.412 $Y2=2.775
r24 14 21 0.820918 $w=3.63e-07 $l=2.6e-08 $layer=LI1_cond $X=7.412 $Y=1.976
+ $X2=7.412 $Y2=2.002
r25 14 32 8.24014 $w=3.63e-07 $l=1.56e-07 $layer=LI1_cond $X=7.412 $Y=1.976
+ $X2=7.412 $Y2=1.82
r26 14 15 10.8614 $w=3.63e-07 $l=3.44e-07 $layer=LI1_cond $X=7.412 $Y=2.061
+ $X2=7.412 $Y2=2.405
r27 14 23 0.820918 $w=3.63e-07 $l=2.6e-08 $layer=LI1_cond $X=7.412 $Y=2.061
+ $X2=7.412 $Y2=2.035
r28 13 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.51 $Y=1.15
+ $X2=7.51 $Y2=1.82
r29 7 13 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=7.415 $Y=0.97
+ $X2=7.415 $Y2=1.15
r30 7 9 13.2851 $w=3.58e-07 $l=4.15e-07 $layer=LI1_cond $X=7.415 $Y=0.97
+ $X2=7.415 $Y2=0.555
r31 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.26
+ $Y=1.84 $X2=7.395 $Y2=1.985
r32 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.26
+ $Y=1.84 $X2=7.395 $Y2=2.815
r33 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.26
+ $Y=0.41 $X2=7.4 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTP_1%VGND 1 2 3 4 13 15 19 21 23 28 33 43 44 50
+ 54
c66 28 0 2.76589e-20 $X=4.995 $Y=0
r67 54 57 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=5.16 $Y=0 $X2=5.16
+ $Y2=0.325
r68 54 55 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r69 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r70 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r71 44 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r72 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r73 41 43 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=7.055 $Y=0 $X2=7.44
+ $Y2=0
r74 40 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r75 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r76 37 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r77 37 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r78 36 39 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r79 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r80 34 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.325 $Y=0 $X2=5.16
+ $Y2=0
r81 34 36 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.325 $Y=0 $X2=5.52
+ $Y2=0
r82 33 64 8.35969 $w=4.63e-07 $l=3.25e-07 $layer=LI1_cond $X=6.822 $Y=0
+ $X2=6.822 $Y2=0.325
r83 33 41 6.7035 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=6.822 $Y=0 $X2=7.055
+ $Y2=0
r84 33 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r85 33 39 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.59 $Y=0 $X2=6.48
+ $Y2=0
r86 32 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r87 31 32 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r88 29 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=1.84
+ $Y2=0
r89 29 31 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=2.16
+ $Y2=0
r90 28 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.995 $Y=0 $X2=5.16
+ $Y2=0
r91 28 31 184.957 $w=1.68e-07 $l=2.835e-06 $layer=LI1_cond $X=4.995 $Y=0
+ $X2=2.16 $Y2=0
r92 27 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r93 27 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r94 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r95 24 47 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r96 24 26 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r97 23 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.675 $Y=0 $X2=1.84
+ $Y2=0
r98 23 26 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.675 $Y=0 $X2=0.72
+ $Y2=0
r99 21 55 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.84 $Y=0 $X2=5.04
+ $Y2=0
r100 21 32 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=2.16 $Y2=0
r101 17 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.84 $Y=0.085
+ $X2=1.84 $Y2=0
r102 17 19 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=1.84 $Y=0.085
+ $X2=1.84 $Y2=0.955
r103 13 47 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r104 13 15 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.715
r105 4 64 182 $w=1.7e-07 $l=3.24731e-07 $layer=licon1_NDIFF $count=1 $X=6.535
+ $Y=0.41 $X2=6.82 $Y2=0.325
r106 3 57 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=4.94
+ $Y=0.41 $X2=5.16 $Y2=0.325
r107 2 19 182 $w=1.7e-07 $l=6.06918e-07 $layer=licon1_NDIFF $count=1 $X=1.675
+ $Y=0.425 $X2=1.84 $Y2=0.955
r108 1 15 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.44 $X2=0.28 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_MS__DLXTP_1%A_239_85# 1 2 9 12 13 14 16 17 18 21 23 24
c71 18 0 1.51199e-20 $X=2.345 $Y=0.84
c72 17 0 1.85283e-19 $X=2.675 $Y=0.84
r73 24 26 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.76 $Y=0.68
+ $X2=2.76 $Y2=0.84
r74 19 24 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.845 $Y=0.68
+ $X2=2.76 $Y2=0.68
r75 19 21 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=2.845 $Y=0.68
+ $X2=3.72 $Y2=0.68
r76 17 26 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.675 $Y=0.84
+ $X2=2.76 $Y2=0.84
r77 17 18 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.675 $Y=0.84
+ $X2=2.345 $Y2=0.84
r78 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.26 $Y=0.925
+ $X2=2.345 $Y2=0.84
r79 15 16 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.26 $Y=0.925
+ $X2=2.26 $Y2=1.355
r80 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.175 $Y=1.44
+ $X2=2.26 $Y2=1.355
r81 13 14 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.175 $Y=1.44
+ $X2=1.505 $Y2=1.44
r82 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.42 $Y=1.355
+ $X2=1.505 $Y2=1.44
r83 12 23 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.42 $Y=1.355
+ $X2=1.42 $Y2=0.93
r84 7 23 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.34 $Y=0.765
+ $X2=1.34 $Y2=0.93
r85 7 9 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.34 $Y=0.765 $X2=1.34
+ $Y2=0.665
r86 2 21 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=3.575
+ $Y=0.425 $X2=3.72 $Y2=0.68
r87 1 9 182 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_NDIFF $count=1 $X=1.195
+ $Y=0.425 $X2=1.34 $Y2=0.665
.ends


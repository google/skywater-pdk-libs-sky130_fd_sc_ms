* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or2b_2 A B_N VGND VNB VPB VPWR X
X0 VGND A a_187_48# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X1 a_473_368# a_27_368# a_187_48# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X2 VPWR a_187_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 X a_187_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X4 VPWR A a_473_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X5 VGND a_187_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 X a_187_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_27_368# B_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X8 a_27_368# B_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X9 a_187_48# a_27_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends

* File: sky130_fd_sc_ms__sdfstp_4.spice
* Created: Fri Aug 28 18:13:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdfstp_4.pex.spice"
.subckt sky130_fd_sc_ms__sdfstp_4  VNB VPB SCE D SCD CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1045 N_VGND_M1045_d N_SCE_M1045_g N_A_27_74#_M1045_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0819 AS=0.1197 PD=0.81 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1040 A_222_74# N_A_27_74#_M1040_g N_VGND_M1045_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0819 PD=0.66 PS=0.81 NRD=18.564 NRS=11.424 M=1 R=2.8 SA=75000.7
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1041 N_A_291_464#_M1041_d N_D_M1041_g A_222_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.09135 AS=0.0504 PD=0.855 PS=0.66 NRD=21.42 NRS=18.564 M=1 R=2.8
+ SA=75001.1 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1016 A_417_74# N_SCE_M1016_g N_A_291_464#_M1041_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.09135 PD=0.66 PS=0.855 NRD=18.564 NRS=22.848 M=1 R=2.8
+ SA=75001.7 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_SCD_M1017_g A_417_74# VNB NLOWVT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_CLK_M1025_g N_A_616_74#_M1025_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1020 N_A_803_74#_M1020_d N_A_616_74#_M1020_g N_VGND_M1025_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_A_1017_81#_M1002_d N_A_616_74#_M1002_g N_A_291_464#_M1002_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1765 PD=0.95 PS=1.73 NRD=71.424 NRS=24.276 M=1
+ R=2.8 SA=75000.3 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1019 A_1153_81# N_A_803_74#_M1019_g N_A_1017_81#_M1002_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.1113 PD=0.66 PS=0.95 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_A_1201_55#_M1018_g A_1153_81# VNB NLOWVT L=0.15 W=0.42
+ AD=0.2084 AS=0.0504 PD=1.95 PS=0.66 NRD=24.276 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1022 A_1445_74# N_A_1017_81#_M1022_g N_A_1201_55#_M1022_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_SET_B_M1003_g A_1445_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.136302 AS=0.0504 PD=0.998491 PS=0.66 NRD=98.568 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1003_d N_A_1017_81#_M1012_g N_A_1677_74#_M1012_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.207698 AS=0.0896 PD=1.52151 PS=0.92 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75001 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1049 N_VGND_M1049_d N_A_1017_81#_M1049_g N_A_1677_74#_M1012_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1006 N_A_1823_524#_M1006_d N_A_803_74#_M1006_g N_A_1677_74#_M1006_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002 A=0.096 P=1.58 MULT=1
MM1036 N_A_1823_524#_M1036_d N_A_803_74#_M1036_g N_A_1677_74#_M1006_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.129147 AS=0.0896 PD=1.20755 PS=0.92 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.6 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1026 A_2149_74# N_A_616_74#_M1026_g N_A_1823_524#_M1036_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0847528 PD=0.66 PS=0.792453 NRD=18.564 NRS=23.568 M=1
+ R=2.8 SA=75001.1 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1004 A_2227_74# N_A_2191_180#_M1004_g A_2149_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0504 PD=0.81 PS=0.66 NRD=39.996 NRS=18.564 M=1 R=2.8 SA=75001.5
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1038 N_VGND_M1038_d N_SET_B_M1038_g A_2227_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1092 AS=0.0819 PD=0.94 PS=0.81 NRD=24.276 NRS=39.996 M=1 R=2.8 SA=75002.1
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1039 N_A_2191_180#_M1039_d N_A_1823_524#_M1039_g N_VGND_M1038_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1197 AS=0.1092 PD=1.41 PS=0.94 NRD=0 NRS=44.28 M=1 R=2.8
+ SA=75002.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_1823_524#_M1005_g N_A_2580_74#_M1005_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1
+ R=4.93333 SA=75000.2 SB=75002.3 A=0.111 P=1.78 MULT=1
MM1001 N_Q_M1001_d N_A_2580_74#_M1001_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.16095 AS=0.1295 PD=1.175 PS=1.09 NRD=13.776 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1015 N_Q_M1001_d N_A_2580_74#_M1015_g N_VGND_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.16095 AS=0.1295 PD=1.175 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.3
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1021 N_Q_M1021_d N_A_2580_74#_M1021_g N_VGND_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.8
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1031 N_Q_M1021_d N_A_2580_74#_M1031_g N_VGND_M1031_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.25955 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.2
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1033 N_VPWR_M1033_d N_SCE_M1033_g N_A_27_74#_M1033_s VPB PSHORT L=0.18 W=0.64
+ AD=0.0864 AS=0.1728 PD=0.91 PS=1.82 NRD=0 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90002.2 A=0.1152 P=1.64 MULT=1
MM1034 A_207_464# N_SCE_M1034_g N_VPWR_M1033_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.0864 PD=0.88 PS=0.91 NRD=19.9955 NRS=0 M=1 R=3.55556 SA=90000.6
+ SB=90001.7 A=0.1152 P=1.64 MULT=1
MM1044 N_A_291_464#_M1044_d N_D_M1044_g A_207_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.144 AS=0.0768 PD=1.09 PS=0.88 NRD=26.1616 NRS=19.9955 M=1 R=3.55556
+ SA=90001 SB=90001.3 A=0.1152 P=1.64 MULT=1
MM1027 A_417_464# N_A_27_74#_M1027_g N_A_291_464#_M1044_d VPB PSHORT L=0.18
+ W=0.64 AD=0.0768 AS=0.144 PD=0.88 PS=1.09 NRD=19.9955 NRS=26.1616 M=1
+ R=3.55556 SA=90001.7 SB=90000.7 A=0.1152 P=1.64 MULT=1
MM1035 N_VPWR_M1035_d N_SCD_M1035_g A_417_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.2858 AS=0.0768 PD=2.37 PS=0.88 NRD=26.1616 NRS=19.9955 M=1 R=3.55556
+ SA=90002.1 SB=90000.3 A=0.1152 P=1.64 MULT=1
MM1042 N_VPWR_M1042_d N_CLK_M1042_g N_A_616_74#_M1042_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1048 N_A_803_74#_M1048_d N_A_616_74#_M1048_g N_VPWR_M1042_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3088 AS=0.1512 PD=2.9 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1008 N_A_1017_81#_M1008_d N_A_803_74#_M1008_g N_A_291_464#_M1008_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.091175 AS=0.1176 PD=0.965 PS=1.4 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90002 A=0.0756 P=1.2 MULT=1
MM1013 A_1143_495# N_A_616_74#_M1013_g N_A_1017_81#_M1008_d VPB PSHORT L=0.18
+ W=0.42 AD=0.084875 AS=0.091175 PD=0.935 PS=0.965 NRD=68.9697 NRS=39.8531 M=1
+ R=2.33333 SA=90000.5 SB=90001.7 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1010_d N_A_1201_55#_M1010_g A_1143_495# VPB PSHORT L=0.18 W=0.42
+ AD=0.150625 AS=0.084875 PD=1.21 PS=0.935 NRD=142.411 NRS=68.9697 M=1 R=2.33333
+ SA=90000.7 SB=90002.5 A=0.0756 P=1.2 MULT=1
MM1028 N_A_1201_55#_M1028_d N_A_1017_81#_M1028_g N_VPWR_M1010_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.063 AS=0.150625 PD=0.72 PS=1.21 NRD=11.7215 NRS=142.411 M=1
+ R=2.33333 SA=90001.5 SB=90001.8 A=0.0756 P=1.2 MULT=1
MM1023 N_VPWR_M1023_d N_SET_B_M1023_g N_A_1201_55#_M1028_d VPB PSHORT L=0.18
+ W=0.42 AD=0.105 AS=0.063 PD=0.893333 PS=0.72 NRD=105.533 NRS=0 M=1 R=2.33333
+ SA=90002 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1024 N_A_1623_373#_M1024_d N_A_1017_81#_M1024_g N_VPWR_M1023_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.1134 AS=0.21 PD=1.11 PS=1.78667 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90001.4 SB=90000.6 A=0.1512 P=2.04 MULT=1
MM1029 N_A_1623_373#_M1024_d N_A_1017_81#_M1029_g N_VPWR_M1029_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1134 AS=0.21915 PD=1.11 PS=2.24 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90001.9 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1043 N_A_1623_373#_M1043_d N_A_616_74#_M1043_g N_A_1823_524#_M1043_s VPB
+ PSHORT L=0.18 W=0.84 AD=0.1134 AS=0.2202 PD=1.11 PS=2.24 NRD=0 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90001.4 A=0.1512 P=2.04 MULT=1
MM1047 N_A_1623_373#_M1043_d N_A_616_74#_M1047_g N_A_1823_524#_M1047_s VPB
+ PSHORT L=0.18 W=0.84 AD=0.1134 AS=0.161 PD=1.11 PS=1.55333 NRD=0 NRS=10.5395
+ M=1 R=4.66667 SA=90000.6 SB=90001 A=0.1512 P=2.04 MULT=1
MM1032 A_2106_508# N_A_803_74#_M1032_g N_A_1823_524#_M1047_s VPB PSHORT L=0.18
+ W=0.42 AD=0.09345 AS=0.0805 PD=0.865 PS=0.776667 NRD=37.5088 NRS=0 M=1
+ R=2.33333 SA=90001.1 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1007 N_VPWR_M1007_d N_A_2191_180#_M1007_g A_2106_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.0567 AS=0.09345 PD=0.69 PS=0.865 NRD=0 NRS=39.8531 M=1 R=2.33333
+ SA=90001.8 SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1011 N_A_1823_524#_M1011_d N_SET_B_M1011_g N_VPWR_M1007_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1176 AS=0.0567 PD=1.4 PS=0.69 NRD=0 NRS=0 M=1 R=2.33333 SA=90002.2
+ SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1037 N_VPWR_M1037_d N_A_1823_524#_M1037_g N_A_2191_180#_M1037_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0805 AS=0.1176 PD=0.776667 PS=1.4 NRD=23.443 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90003 A=0.0756 P=1.2 MULT=1
MM1009 N_A_2580_74#_M1009_d N_A_1823_524#_M1009_g N_VPWR_M1037_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.1134 AS=0.161 PD=1.11 PS=1.55333 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90000.4 SB=90002.5 A=0.1512 P=2.04 MULT=1
MM1014 N_A_2580_74#_M1009_d N_A_1823_524#_M1014_g N_VPWR_M1014_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1134 AS=0.147 PD=1.11 PS=1.23857 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90000.9 SB=90002 A=0.1512 P=2.04 MULT=1
MM1000 N_Q_M1000_d N_A_2580_74#_M1000_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.196 PD=1.39 PS=1.65143 NRD=0 NRS=8.7862 M=1 R=6.22222
+ SA=90001.1 SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1030 N_Q_M1000_d N_A_2580_74#_M1030_g N_VPWR_M1030_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1046 N_Q_M1046_d N_A_2580_74#_M1046_g N_VPWR_M1030_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1050 N_Q_M1046_d N_A_2580_74#_M1050_g N_VPWR_M1050_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.4
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX51_noxref VNB VPB NWDIODE A=30.1692 P=36.16
c_169 VNB 0 7.95967e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__sdfstp_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__o22ai_1.spice
* Created: Wed Sep  2 12:23:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o22ai_1.pex.spice"
.subckt sky130_fd_sc_ms__o22ai_1  VNB VPB B1 B2 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1006 N_Y_M1006_d N_B1_M1006_g N_A_27_74#_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.21275 AS=0.2109 PD=1.315 PS=2.05 NRD=23.508 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002 A=0.111 P=1.78 MULT=1
MM1003 N_A_27_74#_M1003_d N_B2_M1003_g N_Y_M1006_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.21275 PD=1.09 PS=1.315 NRD=11.34 NRS=24.324 M=1 R=4.93333
+ SA=75000.9 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_A2_M1002_g N_A_27_74#_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1295 PD=1.16 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.4
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1004 N_A_27_74#_M1004_d N_A1_M1004_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 A_145_368# N_B1_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12 AD=0.1344
+ AS=0.448 PD=1.36 PS=3.04 NRD=11.426 NRS=20.2122 M=1 R=6.22222 SA=90000.3
+ SB=90001.8 A=0.2016 P=2.6 MULT=1
MM1000 N_Y_M1000_d N_B2_M1000_g A_145_368# VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.1344 PD=1.51 PS=1.36 NRD=8.7862 NRS=11.426 M=1 R=6.22222 SA=90000.7
+ SB=90001.3 A=0.2016 P=2.6 MULT=1
MM1007 A_343_368# N_A2_M1007_g N_Y_M1000_d VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.2184 PD=1.51 PS=1.51 NRD=24.6053 NRS=10.5395 M=1 R=6.22222 SA=90001.3
+ SB=90000.8 A=0.2016 P=2.6 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g A_343_368# VPB PSHORT L=0.18 W=1.12 AD=0.3136
+ AS=0.2184 PD=2.8 PS=1.51 NRD=0 NRS=24.6053 M=1 R=6.22222 SA=90001.9 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ms__o22ai_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__a2111o_4.spice
* Created: Fri Aug 28 16:55:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a2111o_4.pex.spice"
.subckt sky130_fd_sc_ms__a2111o_4  VNB VPB D1 C1 B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_137_260#_M1003_g N_X_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.8 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A_137_260#_M1010_g N_X_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75003.3 A=0.111 P=1.78 MULT=1
MM1020 N_VGND_M1010_d N_A_137_260#_M1020_g N_X_M1020_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1024 N_VGND_M1024_d N_A_137_260#_M1024_g N_X_M1020_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.124942 AS=0.1036 PD=1.14217 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1011 N_A_137_260#_M1011_d N_D1_M1011_g N_VGND_M1024_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.108058 PD=0.92 PS=0.987826 NRD=0 NRS=8.436 M=1 R=4.26667
+ SA=75002 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1021 N_A_137_260#_M1011_d N_D1_M1021_g N_VGND_M1021_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0928 PD=0.92 PS=0.93 NRD=0 NRS=0.936 M=1 R=4.26667 SA=75002.4
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1004 N_VGND_M1021_s N_C1_M1004_g N_A_137_260#_M1004_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0928 AS=0.0896 PD=0.93 PS=0.92 NRD=0.936 NRS=0 M=1 R=4.26667 SA=75002.8
+ SB=75001.5 A=0.096 P=1.58 MULT=1
MM1022 N_VGND_M1022_d N_C1_M1022_g N_A_137_260#_M1004_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0928 AS=0.0896 PD=0.93 PS=0.92 NRD=0.936 NRS=0 M=1 R=4.26667 SA=75003.3
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1009 N_VGND_M1022_d N_B1_M1009_g N_A_137_260#_M1009_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0928 AS=0.0896 PD=0.93 PS=0.92 NRD=0.936 NRS=0 M=1 R=4.26667 SA=75003.7
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1026 N_VGND_M1026_d N_B1_M1026_g N_A_137_260#_M1009_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75004.1
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_A_137_260#_M1001_d N_A1_M1001_g N_A_1210_74#_M1001_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1012 N_A_137_260#_M1001_d N_A1_M1012_g N_A_1210_74#_M1012_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1007 N_A_1210_74#_M1012_s N_A2_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1027 N_A_1210_74#_M1027_d N_A2_M1027_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1014 N_X_M1014_d N_A_137_260#_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1016 N_X_M1014_d N_A_137_260#_M1016_g N_VPWR_M1016_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1018 N_X_M1018_d N_A_137_260#_M1018_g N_VPWR_M1016_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1023 N_X_M1018_d N_A_137_260#_M1023_g N_VPWR_M1023_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1002 N_A_137_260#_M1002_d N_D1_M1002_g N_A_549_392#_M1002_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.5 A=0.18 P=2.36 MULT=1
MM1005 N_A_137_260#_M1002_d N_D1_M1005_g N_A_549_392#_M1005_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.6
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1006 N_A_817_392#_M1006_d N_C1_M1006_g N_A_549_392#_M1005_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.1
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1008 N_A_817_392#_M1006_d N_C1_M1008_g N_A_549_392#_M1008_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.5
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1013 N_A_817_392#_M1013_d N_B1_M1013_g N_A_1013_392#_M1013_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90002.4 A=0.18 P=2.36 MULT=1
MM1015 N_A_817_392#_M1013_d N_B1_M1015_g N_A_1013_392#_M1015_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.6
+ SB=90002 A=0.18 P=2.36 MULT=1
MM1017 N_VPWR_M1017_d N_A1_M1017_g N_A_1013_392#_M1015_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.1
+ SB=90001.5 A=0.18 P=2.36 MULT=1
MM1019 N_VPWR_M1017_d N_A1_M1019_g N_A_1013_392#_M1019_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.5
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1000 N_A_1013_392#_M1019_s N_A2_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90002
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1025 N_A_1013_392#_M1025_d N_A2_M1025_g N_VPWR_M1000_s VPB PSHORT L=0.18 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90002.4
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.8844 P=20.8
c_88 VNB 0 1.80394e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__a2111o_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__einvp_8.pex.spice
* Created: Wed Sep  2 12:08:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__EINVP_8%A 3 5 7 8 10 13 17 19 21 24 26 28 31 33 35
+ 38 40 42 45 47 49 52 54 56 57 58 59 60 61 97 99
c162 99 0 5.65346e-20 $X=3.65 $Y=1.385
c163 54 0 1.9142e-19 $X=3.925 $Y=1.22
c164 52 0 1.88192e-19 $X=3.65 $Y=2.4
c165 47 0 8.60601e-20 $X=3.425 $Y=1.22
c166 33 0 8.60601e-20 $X=2.425 $Y=1.22
c167 19 0 8.60869e-20 $X=1.425 $Y=1.22
r168 98 99 34.3196 $w=3.16e-07 $l=2.25e-07 $layer=POLY_cond $X=3.425 $Y=1.385
+ $X2=3.65 $Y2=1.385
r169 96 98 19.8291 $w=3.16e-07 $l=1.3e-07 $layer=POLY_cond $X=3.295 $Y=1.385
+ $X2=3.425 $Y2=1.385
r170 96 97 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.295
+ $Y=1.385 $X2=3.295 $Y2=1.385
r171 94 96 14.4905 $w=3.16e-07 $l=9.5e-08 $layer=POLY_cond $X=3.2 $Y=1.385
+ $X2=3.295 $Y2=1.385
r172 93 94 41.9462 $w=3.16e-07 $l=2.75e-07 $layer=POLY_cond $X=2.925 $Y=1.385
+ $X2=3.2 $Y2=1.385
r173 92 93 26.693 $w=3.16e-07 $l=1.75e-07 $layer=POLY_cond $X=2.75 $Y=1.385
+ $X2=2.925 $Y2=1.385
r174 90 92 20.5918 $w=3.16e-07 $l=1.35e-07 $layer=POLY_cond $X=2.615 $Y=1.385
+ $X2=2.75 $Y2=1.385
r175 90 91 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.615
+ $Y=1.385 $X2=2.615 $Y2=1.385
r176 88 90 28.981 $w=3.16e-07 $l=1.9e-07 $layer=POLY_cond $X=2.425 $Y=1.385
+ $X2=2.615 $Y2=1.385
r177 87 88 19.0665 $w=3.16e-07 $l=1.25e-07 $layer=POLY_cond $X=2.3 $Y=1.385
+ $X2=2.425 $Y2=1.385
r178 86 91 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.275 $Y=1.365
+ $X2=2.615 $Y2=1.365
r179 85 87 3.81329 $w=3.16e-07 $l=2.5e-08 $layer=POLY_cond $X=2.275 $Y=1.385
+ $X2=2.3 $Y2=1.385
r180 85 86 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.275
+ $Y=1.385 $X2=2.275 $Y2=1.385
r181 83 85 53.3861 $w=3.16e-07 $l=3.5e-07 $layer=POLY_cond $X=1.925 $Y=1.385
+ $X2=2.275 $Y2=1.385
r182 82 83 11.4399 $w=3.16e-07 $l=7.5e-08 $layer=POLY_cond $X=1.85 $Y=1.385
+ $X2=1.925 $Y2=1.385
r183 80 82 38.8956 $w=3.16e-07 $l=2.55e-07 $layer=POLY_cond $X=1.595 $Y=1.385
+ $X2=1.85 $Y2=1.385
r184 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.595
+ $Y=1.385 $X2=1.595 $Y2=1.385
r185 78 80 25.9304 $w=3.16e-07 $l=1.7e-07 $layer=POLY_cond $X=1.425 $Y=1.385
+ $X2=1.595 $Y2=1.385
r186 77 78 3.81329 $w=3.16e-07 $l=2.5e-08 $layer=POLY_cond $X=1.4 $Y=1.385
+ $X2=1.425 $Y2=1.385
r187 76 81 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.255 $Y=1.365
+ $X2=1.595 $Y2=1.365
r188 75 77 22.1171 $w=3.16e-07 $l=1.45e-07 $layer=POLY_cond $X=1.255 $Y=1.385
+ $X2=1.4 $Y2=1.385
r189 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.255
+ $Y=1.385 $X2=1.255 $Y2=1.385
r190 73 75 46.5222 $w=3.16e-07 $l=3.05e-07 $layer=POLY_cond $X=0.95 $Y=1.385
+ $X2=1.255 $Y2=1.385
r191 72 73 3.81329 $w=3.16e-07 $l=2.5e-08 $layer=POLY_cond $X=0.925 $Y=1.385
+ $X2=0.95 $Y2=1.385
r192 70 72 1.52532 $w=3.16e-07 $l=1e-08 $layer=POLY_cond $X=0.915 $Y=1.385
+ $X2=0.925 $Y2=1.385
r193 70 71 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.915
+ $Y=1.385 $X2=0.915 $Y2=1.385
r194 68 70 63.3006 $w=3.16e-07 $l=4.15e-07 $layer=POLY_cond $X=0.5 $Y=1.385
+ $X2=0.915 $Y2=1.385
r195 67 68 0.762658 $w=3.16e-07 $l=5e-09 $layer=POLY_cond $X=0.495 $Y=1.385
+ $X2=0.5 $Y2=1.385
r196 61 97 5.45074 $w=3.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.12 $Y=1.365
+ $X2=3.295 $Y2=1.365
r197 60 61 14.9506 $w=3.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.365
+ $X2=3.12 $Y2=1.365
r198 60 91 0.778678 $w=3.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.64 $Y=1.365
+ $X2=2.615 $Y2=1.365
r199 59 86 3.58192 $w=3.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.16 $Y=1.365
+ $X2=2.275 $Y2=1.365
r200 58 59 14.9506 $w=3.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=2.16 $Y2=1.365
r201 58 81 2.6475 $w=3.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=1.595 $Y2=1.365
r202 57 76 1.71309 $w=3.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.2 $Y=1.365
+ $X2=1.255 $Y2=1.365
r203 57 71 8.87693 $w=3.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.2 $Y=1.365
+ $X2=0.915 $Y2=1.365
r204 54 99 41.9462 $w=3.16e-07 $l=3.47851e-07 $layer=POLY_cond $X=3.925 $Y=1.22
+ $X2=3.65 $Y2=1.385
r205 54 56 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.925 $Y=1.22
+ $X2=3.925 $Y2=0.74
r206 50 99 15.9236 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.65 $Y=1.55
+ $X2=3.65 $Y2=1.385
r207 50 52 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.65 $Y=1.55
+ $X2=3.65 $Y2=2.4
r208 47 98 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.425 $Y=1.22
+ $X2=3.425 $Y2=1.385
r209 47 49 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.425 $Y=1.22
+ $X2=3.425 $Y2=0.74
r210 43 94 15.9236 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.2 $Y=1.55
+ $X2=3.2 $Y2=1.385
r211 43 45 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.2 $Y=1.55 $X2=3.2
+ $Y2=2.4
r212 40 93 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.925 $Y=1.22
+ $X2=2.925 $Y2=1.385
r213 40 42 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.925 $Y=1.22
+ $X2=2.925 $Y2=0.74
r214 36 92 15.9236 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.75 $Y=1.55
+ $X2=2.75 $Y2=1.385
r215 36 38 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.75 $Y=1.55
+ $X2=2.75 $Y2=2.4
r216 33 88 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.425 $Y=1.22
+ $X2=2.425 $Y2=1.385
r217 33 35 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.425 $Y=1.22
+ $X2=2.425 $Y2=0.74
r218 29 87 15.9236 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.3 $Y=1.55
+ $X2=2.3 $Y2=1.385
r219 29 31 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.3 $Y=1.55 $X2=2.3
+ $Y2=2.4
r220 26 83 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.22
+ $X2=1.925 $Y2=1.385
r221 26 28 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.925 $Y=1.22
+ $X2=1.925 $Y2=0.74
r222 22 82 15.9236 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.85 $Y=1.55
+ $X2=1.85 $Y2=1.385
r223 22 24 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.85 $Y=1.55
+ $X2=1.85 $Y2=2.4
r224 19 78 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.22
+ $X2=1.425 $Y2=1.385
r225 19 21 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.425 $Y=1.22
+ $X2=1.425 $Y2=0.74
r226 15 77 15.9236 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.4 $Y=1.55
+ $X2=1.4 $Y2=1.385
r227 15 17 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.4 $Y=1.55 $X2=1.4
+ $Y2=2.4
r228 11 73 15.9236 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=1.55
+ $X2=0.95 $Y2=1.385
r229 11 13 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.95 $Y=1.55
+ $X2=0.95 $Y2=2.4
r230 8 72 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.22
+ $X2=0.925 $Y2=1.385
r231 8 10 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.925 $Y=1.22
+ $X2=0.925 $Y2=0.74
r232 5 67 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.495 $Y2=1.385
r233 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.495 $Y2=0.74
r234 1 68 15.9236 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.55 $X2=0.5
+ $Y2=1.385
r235 1 3 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.5 $Y=1.55 $X2=0.5
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__EINVP_8%A_802_323# 1 2 7 9 10 11 12 14 15 17 19 20
+ 22 24 25 27 29 30 32 34 35 37 39 40 42 44 45 47 48 49 50 51 52 53 56 59 63 68
c179 56 0 3.05834e-20 $X=8.14 $Y=1.615
r180 68 70 17.9954 $w=4.48e-07 $l=4.95e-07 $layer=LI1_cond $X=8.28 $Y=0.515
+ $X2=8.28 $Y2=1.01
r181 63 66 0.249659 $w=7.33e-07 $l=1.5e-08 $layer=LI1_cond $X=8.17 $Y=2.8
+ $X2=8.17 $Y2=2.815
r182 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.94
+ $Y=2.8 $X2=7.94 $Y2=2.8
r183 61 63 13.5648 $w=7.33e-07 $l=8.15e-07 $layer=LI1_cond $X=8.17 $Y=1.985
+ $X2=8.17 $Y2=2.8
r184 59 64 178.359 $w=3.3e-07 $l=1.02e-06 $layer=POLY_cond $X=7.94 $Y=1.78
+ $X2=7.94 $Y2=2.8
r185 58 61 3.41201 $w=7.33e-07 $l=2.05e-07 $layer=LI1_cond $X=8.17 $Y=1.78
+ $X2=8.17 $Y2=1.985
r186 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.94
+ $Y=1.78 $X2=7.94 $Y2=1.78
r187 56 58 11.2359 $w=7.33e-07 $l=1.79374e-07 $layer=LI1_cond $X=8.14 $Y=1.615
+ $X2=8.17 $Y2=1.78
r188 56 70 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=8.14 $Y=1.615
+ $X2=8.14 $Y2=1.01
r189 54 59 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.94 $Y=1.765
+ $X2=7.94 $Y2=1.78
r190 46 53 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.34 $Y=1.69 $X2=7.25
+ $Y2=1.69
r191 45 54 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=7.775 $Y=1.69
+ $X2=7.94 $Y2=1.765
r192 45 46 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.775 $Y=1.69
+ $X2=7.34 $Y2=1.69
r193 42 53 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=7.25 $Y=1.765
+ $X2=7.25 $Y2=1.69
r194 42 44 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=7.25 $Y=1.765
+ $X2=7.25 $Y2=2.4
r195 41 52 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.89 $Y=1.69 $X2=6.8
+ $Y2=1.69
r196 40 53 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.16 $Y=1.69 $X2=7.25
+ $Y2=1.69
r197 40 41 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=7.16 $Y=1.69
+ $X2=6.89 $Y2=1.69
r198 37 52 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=6.8 $Y=1.765 $X2=6.8
+ $Y2=1.69
r199 37 39 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=6.8 $Y=1.765
+ $X2=6.8 $Y2=2.4
r200 36 51 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.44 $Y=1.69 $X2=6.35
+ $Y2=1.69
r201 35 52 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.71 $Y=1.69 $X2=6.8
+ $Y2=1.69
r202 35 36 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=6.71 $Y=1.69
+ $X2=6.44 $Y2=1.69
r203 32 51 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=6.35 $Y=1.765
+ $X2=6.35 $Y2=1.69
r204 32 34 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=6.35 $Y=1.765
+ $X2=6.35 $Y2=2.4
r205 31 50 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.99 $Y=1.69 $X2=5.9
+ $Y2=1.69
r206 30 51 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.26 $Y=1.69 $X2=6.35
+ $Y2=1.69
r207 30 31 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=6.26 $Y=1.69
+ $X2=5.99 $Y2=1.69
r208 27 50 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=5.9 $Y=1.765 $X2=5.9
+ $Y2=1.69
r209 27 29 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=5.9 $Y=1.765
+ $X2=5.9 $Y2=2.4
r210 26 49 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.54 $Y=1.69 $X2=5.45
+ $Y2=1.69
r211 25 50 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.81 $Y=1.69 $X2=5.9
+ $Y2=1.69
r212 25 26 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.81 $Y=1.69
+ $X2=5.54 $Y2=1.69
r213 22 49 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=5.45 $Y=1.765
+ $X2=5.45 $Y2=1.69
r214 22 24 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=5.45 $Y=1.765
+ $X2=5.45 $Y2=2.4
r215 21 48 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.09 $Y=1.69 $X2=5
+ $Y2=1.69
r216 20 49 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.36 $Y=1.69 $X2=5.45
+ $Y2=1.69
r217 20 21 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.36 $Y=1.69
+ $X2=5.09 $Y2=1.69
r218 17 48 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=5 $Y=1.765 $X2=5
+ $Y2=1.69
r219 17 19 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=5 $Y=1.765 $X2=5
+ $Y2=2.4
r220 16 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.64 $Y=1.69 $X2=4.55
+ $Y2=1.69
r221 15 48 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.91 $Y=1.69 $X2=5
+ $Y2=1.69
r222 15 16 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.91 $Y=1.69
+ $X2=4.64 $Y2=1.69
r223 12 47 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.55 $Y=1.765
+ $X2=4.55 $Y2=1.69
r224 12 14 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=4.55 $Y=1.765
+ $X2=4.55 $Y2=2.4
r225 10 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.46 $Y=1.69 $X2=4.55
+ $Y2=1.69
r226 10 11 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.46 $Y=1.69
+ $X2=4.19 $Y2=1.69
r227 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.1 $Y=1.765
+ $X2=4.19 $Y2=1.69
r228 7 9 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=4.1 $Y=1.765 $X2=4.1
+ $Y2=2.4
r229 2 66 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.265
+ $Y=1.84 $X2=8.4 $Y2=2.815
r230 2 61 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.265
+ $Y=1.84 $X2=8.4 $Y2=1.985
r231 1 68 91 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=2 $X=8.19
+ $Y=0.37 $X2=8.34 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__EINVP_8%TE 1 3 4 5 6 8 9 11 13 14 16 18 19 21 23 24
+ 26 28 29 31 33 34 36 38 39 43 46 48 49 50 51 52 53 54 55 57 58
c152 36 0 3.05834e-20 $X=7.505 $Y=1.22
c153 31 0 1.07496e-19 $X=7.005 $Y=1.22
c154 6 0 1.07496e-19 $X=4.855 $Y=1.22
c155 1 0 3.03515e-19 $X=4.355 $Y=1.22
r156 60 62 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.6 $Y=1.385
+ $X2=8.6 $Y2=1.55
r157 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.6
+ $Y=1.385 $X2=8.6 $Y2=1.385
r158 57 60 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.6 $Y=1.295 $X2=8.6
+ $Y2=1.385
r159 57 58 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.6 $Y=1.295 $X2=8.6
+ $Y2=1.22
r160 55 61 10.9487 $w=3.12e-07 $l=2.8e-07 $layer=LI1_cond $X=8.88 $Y=1.365
+ $X2=8.6 $Y2=1.365
r161 46 62 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=8.625 $Y=2.4
+ $X2=8.625 $Y2=1.55
r162 43 58 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.555 $Y=0.74
+ $X2=8.555 $Y2=1.22
r163 40 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.58 $Y=1.295
+ $X2=7.505 $Y2=1.295
r164 39 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.435 $Y=1.295
+ $X2=8.6 $Y2=1.295
r165 39 40 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=8.435 $Y=1.295
+ $X2=7.58 $Y2=1.295
r166 36 54 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.505 $Y=1.22
+ $X2=7.505 $Y2=1.295
r167 36 38 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.505 $Y=1.22
+ $X2=7.505 $Y2=0.74
r168 35 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.08 $Y=1.295
+ $X2=7.005 $Y2=1.295
r169 34 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.43 $Y=1.295
+ $X2=7.505 $Y2=1.295
r170 34 35 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=7.43 $Y=1.295
+ $X2=7.08 $Y2=1.295
r171 31 53 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.005 $Y=1.22
+ $X2=7.005 $Y2=1.295
r172 31 33 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.005 $Y=1.22
+ $X2=7.005 $Y2=0.74
r173 30 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.65 $Y=1.295
+ $X2=6.575 $Y2=1.295
r174 29 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.93 $Y=1.295
+ $X2=7.005 $Y2=1.295
r175 29 30 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.93 $Y=1.295
+ $X2=6.65 $Y2=1.295
r176 26 52 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.575 $Y=1.22
+ $X2=6.575 $Y2=1.295
r177 26 28 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.575 $Y=1.22
+ $X2=6.575 $Y2=0.74
r178 25 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.22 $Y=1.295
+ $X2=6.145 $Y2=1.295
r179 24 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.5 $Y=1.295
+ $X2=6.575 $Y2=1.295
r180 24 25 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.5 $Y=1.295
+ $X2=6.22 $Y2=1.295
r181 21 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.145 $Y=1.22
+ $X2=6.145 $Y2=1.295
r182 21 23 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.145 $Y=1.22
+ $X2=6.145 $Y2=0.74
r183 20 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.79 $Y=1.295
+ $X2=5.715 $Y2=1.295
r184 19 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.07 $Y=1.295
+ $X2=6.145 $Y2=1.295
r185 19 20 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.07 $Y=1.295
+ $X2=5.79 $Y2=1.295
r186 16 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.715 $Y=1.22
+ $X2=5.715 $Y2=1.295
r187 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.715 $Y=1.22
+ $X2=5.715 $Y2=0.74
r188 15 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.36 $Y=1.295
+ $X2=5.285 $Y2=1.295
r189 14 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.64 $Y=1.295
+ $X2=5.715 $Y2=1.295
r190 14 15 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.64 $Y=1.295
+ $X2=5.36 $Y2=1.295
r191 11 49 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.285 $Y=1.22
+ $X2=5.285 $Y2=1.295
r192 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.285 $Y=1.22
+ $X2=5.285 $Y2=0.74
r193 10 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.93 $Y=1.295
+ $X2=4.855 $Y2=1.295
r194 9 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.21 $Y=1.295
+ $X2=5.285 $Y2=1.295
r195 9 10 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.21 $Y=1.295
+ $X2=4.93 $Y2=1.295
r196 6 48 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.855 $Y=1.22
+ $X2=4.855 $Y2=1.295
r197 6 8 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.855 $Y=1.22
+ $X2=4.855 $Y2=0.74
r198 4 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.78 $Y=1.295
+ $X2=4.855 $Y2=1.295
r199 4 5 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.78 $Y=1.295
+ $X2=4.43 $Y2=1.295
r200 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.355 $Y=1.22
+ $X2=4.43 $Y2=1.295
r201 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.355 $Y=1.22
+ $X2=4.355 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__EINVP_8%A_27_368# 1 2 3 4 5 6 7 8 9 30 34 35 38 40
+ 44 46 50 52 54 56 61 64 66 67 70 74 78 82 86 90 91 92 95 96 97
r156 86 88 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=7.435 $Y=1.985
+ $X2=7.435 $Y2=2.815
r157 84 86 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=7.435 $Y=1.72
+ $X2=7.435 $Y2=1.985
r158 83 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.66 $Y=1.635
+ $X2=6.535 $Y2=1.635
r159 82 84 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.31 $Y=1.635
+ $X2=7.435 $Y2=1.72
r160 82 83 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=7.31 $Y=1.635
+ $X2=6.66 $Y2=1.635
r161 78 80 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=6.535 $Y=1.985
+ $X2=6.535 $Y2=2.815
r162 76 97 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.535 $Y=1.72
+ $X2=6.535 $Y2=1.635
r163 76 78 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=6.535 $Y=1.72
+ $X2=6.535 $Y2=1.985
r164 75 96 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.76 $Y=1.635
+ $X2=5.635 $Y2=1.635
r165 74 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.41 $Y=1.635
+ $X2=6.535 $Y2=1.635
r166 74 75 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.41 $Y=1.635
+ $X2=5.76 $Y2=1.635
r167 70 72 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=5.635 $Y=1.985
+ $X2=5.635 $Y2=2.815
r168 68 96 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.635 $Y=1.72
+ $X2=5.635 $Y2=1.635
r169 68 70 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=5.635 $Y=1.72
+ $X2=5.635 $Y2=1.985
r170 66 96 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.51 $Y=1.635
+ $X2=5.635 $Y2=1.635
r171 66 67 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.51 $Y=1.635
+ $X2=4.94 $Y2=1.635
r172 62 95 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.815 $Y=2.23
+ $X2=4.815 $Y2=2.145
r173 62 64 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=4.815 $Y=2.23
+ $X2=4.815 $Y2=2.4
r174 59 95 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.815 $Y=2.06
+ $X2=4.815 $Y2=2.145
r175 59 61 3.45733 $w=2.48e-07 $l=7.5e-08 $layer=LI1_cond $X=4.815 $Y=2.06
+ $X2=4.815 $Y2=1.985
r176 58 67 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.815 $Y=1.72
+ $X2=4.94 $Y2=1.635
r177 58 61 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=4.815 $Y=1.72
+ $X2=4.815 $Y2=1.985
r178 57 94 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.96 $Y=2.145
+ $X2=3.875 $Y2=2.145
r179 56 95 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.69 $Y=2.145
+ $X2=4.815 $Y2=2.145
r180 56 57 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.69 $Y=2.145
+ $X2=3.96 $Y2=2.145
r181 54 94 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.875 $Y=2.23
+ $X2=3.875 $Y2=2.145
r182 54 55 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=3.875 $Y=2.23
+ $X2=3.875 $Y2=2.905
r183 53 92 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.075 $Y=2.99
+ $X2=2.975 $Y2=2.99
r184 52 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.79 $Y=2.99
+ $X2=3.875 $Y2=2.905
r185 52 53 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=3.79 $Y=2.99
+ $X2=3.075 $Y2=2.99
r186 48 92 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=2.905
+ $X2=2.975 $Y2=2.99
r187 48 50 37.7091 $w=1.98e-07 $l=6.8e-07 $layer=LI1_cond $X=2.975 $Y=2.905
+ $X2=2.975 $Y2=2.225
r188 47 91 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.19 $Y=2.99
+ $X2=2.08 $Y2=2.99
r189 46 92 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.875 $Y=2.99
+ $X2=2.975 $Y2=2.99
r190 46 47 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=2.875 $Y=2.99
+ $X2=2.19 $Y2=2.99
r191 42 91 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=2.905
+ $X2=2.08 $Y2=2.99
r192 42 44 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=2.08 $Y=2.905
+ $X2=2.08 $Y2=2.225
r193 41 90 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=1.275 $Y=2.99
+ $X2=1.172 $Y2=2.99
r194 40 91 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.97 $Y=2.99
+ $X2=2.08 $Y2=2.99
r195 40 41 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.97 $Y=2.99
+ $X2=1.275 $Y2=2.99
r196 36 90 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.172 $Y=2.905
+ $X2=1.172 $Y2=2.99
r197 36 38 36.7894 $w=2.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.172 $Y=2.905
+ $X2=1.172 $Y2=2.225
r198 34 90 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=1.07 $Y=2.99
+ $X2=1.172 $Y2=2.99
r199 34 35 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.07 $Y=2.99
+ $X2=0.375 $Y2=2.99
r200 30 33 36.0954 $w=2.63e-07 $l=8.3e-07 $layer=LI1_cond $X=0.242 $Y=1.985
+ $X2=0.242 $Y2=2.815
r201 28 35 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=0.242 $Y=2.905
+ $X2=0.375 $Y2=2.99
r202 28 33 3.91396 $w=2.63e-07 $l=9e-08 $layer=LI1_cond $X=0.242 $Y=2.905
+ $X2=0.242 $Y2=2.815
r203 9 88 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.34
+ $Y=1.84 $X2=7.475 $Y2=2.815
r204 9 86 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.34
+ $Y=1.84 $X2=7.475 $Y2=1.985
r205 8 80 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.44
+ $Y=1.84 $X2=6.575 $Y2=2.815
r206 8 78 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.44
+ $Y=1.84 $X2=6.575 $Y2=1.985
r207 7 72 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.54
+ $Y=1.84 $X2=5.675 $Y2=2.815
r208 7 70 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.54
+ $Y=1.84 $X2=5.675 $Y2=1.985
r209 6 64 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=4.64
+ $Y=1.84 $X2=4.775 $Y2=2.4
r210 6 61 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.64
+ $Y=1.84 $X2=4.775 $Y2=1.985
r211 5 94 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=3.74
+ $Y=1.84 $X2=3.875 $Y2=2.225
r212 4 50 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=2.84
+ $Y=1.84 $X2=2.975 $Y2=2.225
r213 3 44 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=1.94
+ $Y=1.84 $X2=2.075 $Y2=2.225
r214 2 38 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=1.04
+ $Y=1.84 $X2=1.175 $Y2=2.225
r215 1 33 400 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.275 $Y2=2.815
r216 1 30 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.275 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__EINVP_8%Z 1 2 3 4 5 6 7 8 27 33 34 37 41 47 51 53 57
+ 62 64 68 71 72 73 76 77 79 83
c128 79 0 1.86694e-19 $X=3.71 $Y=0.76
c129 62 0 1.16821e-19 $X=3.79 $Y=1.55
r130 83 86 13.6602 $w=2.59e-07 $l=2.9e-07 $layer=LI1_cond $X=4.08 $Y=1.72
+ $X2=3.79 $Y2=1.72
r131 81 82 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.71 $Y=0.925
+ $X2=3.71 $Y2=1.01
r132 79 81 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.71 $Y=0.76
+ $X2=3.71 $Y2=0.925
r133 75 77 8.6272 $w=3.93e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=0.812
+ $X2=2.875 $Y2=0.812
r134 75 76 8.6272 $w=3.93e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=0.812
+ $X2=2.545 $Y2=0.812
r135 72 76 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.875 $Y=0.925
+ $X2=2.545 $Y2=0.925
r136 70 72 8.6272 $w=3.93e-07 $l=1.65e-07 $layer=LI1_cond $X=1.71 $Y=0.812
+ $X2=1.875 $Y2=0.812
r137 70 71 8.6272 $w=3.93e-07 $l=1.65e-07 $layer=LI1_cond $X=1.71 $Y=0.812
+ $X2=1.545 $Y2=0.812
r138 64 66 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=0.75 $Y=0.78
+ $X2=0.75 $Y2=0.925
r139 62 86 3.20129 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.79 $Y=1.55
+ $X2=3.79 $Y2=1.72
r140 62 82 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.79 $Y=1.55
+ $X2=3.79 $Y2=1.01
r141 57 59 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.425 $Y=1.97
+ $X2=3.425 $Y2=2.65
r142 55 86 17.1931 $w=2.59e-07 $l=3.65e-07 $layer=LI1_cond $X=3.425 $Y=1.72
+ $X2=3.79 $Y2=1.72
r143 55 57 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.425 $Y=1.89
+ $X2=3.425 $Y2=1.97
r144 53 81 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.545 $Y=0.925
+ $X2=3.71 $Y2=0.925
r145 53 77 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.545 $Y=0.925
+ $X2=2.875 $Y2=0.925
r146 52 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=1.805
+ $X2=2.525 $Y2=1.805
r147 51 55 9.21269 $w=2.59e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.26 $Y=1.805
+ $X2=3.425 $Y2=1.72
r148 51 52 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.26 $Y=1.805
+ $X2=2.69 $Y2=1.805
r149 47 49 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.525 $Y=1.97
+ $X2=2.525 $Y2=2.65
r150 45 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=1.89
+ $X2=2.525 $Y2=1.805
r151 45 47 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.525 $Y=1.89
+ $X2=2.525 $Y2=1.97
r152 42 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.79 $Y=1.805
+ $X2=1.625 $Y2=1.805
r153 41 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=1.805
+ $X2=2.525 $Y2=1.805
r154 41 42 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.36 $Y=1.805
+ $X2=1.79 $Y2=1.805
r155 37 39 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.625 $Y=1.97
+ $X2=1.625 $Y2=2.65
r156 35 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=1.89
+ $X2=1.625 $Y2=1.805
r157 35 37 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.625 $Y=1.89
+ $X2=1.625 $Y2=1.97
r158 33 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.46 $Y=1.805
+ $X2=1.625 $Y2=1.805
r159 33 34 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.46 $Y=1.805
+ $X2=0.89 $Y2=1.805
r160 32 66 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=0.925
+ $X2=0.75 $Y2=0.925
r161 32 71 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.875 $Y=0.925
+ $X2=1.545 $Y2=0.925
r162 27 29 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.725 $Y=1.97
+ $X2=0.725 $Y2=2.65
r163 25 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.725 $Y=1.89
+ $X2=0.89 $Y2=1.805
r164 25 27 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=0.725 $Y=1.89
+ $X2=0.725 $Y2=1.97
r165 8 59 400 $w=1.7e-07 $l=8.749e-07 $layer=licon1_PDIFF $count=1 $X=3.29
+ $Y=1.84 $X2=3.425 $Y2=2.65
r166 8 57 400 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_PDIFF $count=1 $X=3.29
+ $Y=1.84 $X2=3.425 $Y2=1.97
r167 7 49 400 $w=1.7e-07 $l=8.749e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=1.84 $X2=2.525 $Y2=2.65
r168 7 47 400 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=1.84 $X2=2.525 $Y2=1.97
r169 6 39 400 $w=1.7e-07 $l=8.749e-07 $layer=licon1_PDIFF $count=1 $X=1.49
+ $Y=1.84 $X2=1.625 $Y2=2.65
r170 6 37 400 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_PDIFF $count=1 $X=1.49
+ $Y=1.84 $X2=1.625 $Y2=1.97
r171 5 29 400 $w=1.7e-07 $l=8.749e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.84 $X2=0.725 $Y2=2.65
r172 5 27 400 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.84 $X2=0.725 $Y2=1.97
r173 4 79 182 $w=1.7e-07 $l=4.83735e-07 $layer=licon1_NDIFF $count=1 $X=3.5
+ $Y=0.37 $X2=3.71 $Y2=0.76
r174 3 75 182 $w=1.7e-07 $l=5.04182e-07 $layer=licon1_NDIFF $count=1 $X=2.5
+ $Y=0.37 $X2=2.71 $Y2=0.78
r175 2 70 182 $w=1.7e-07 $l=5.04182e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.71 $Y2=0.78
r176 1 64 182 $w=1.7e-07 $l=4.74868e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_MS__EINVP_8%VPWR 1 2 3 4 5 18 22 26 30 36 40 42 47 48 49
+ 50 51 63 68 77 80 84
c108 18 0 1.88192e-19 $X=4.325 $Y=2.485
r109 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r110 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r111 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r112 75 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r113 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r114 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r115 72 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r116 71 74 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=7.44 $Y=3.33 $X2=8.4
+ $Y2=3.33
r117 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r118 69 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.11 $Y=3.33
+ $X2=6.985 $Y2=3.33
r119 69 71 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.11 $Y=3.33
+ $X2=7.44 $Y2=3.33
r120 68 83 4.02656 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=8.765 $Y=3.33
+ $X2=8.942 $Y2=3.33
r121 68 74 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.765 $Y=3.33
+ $X2=8.4 $Y2=3.33
r122 67 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r123 67 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r124 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r125 64 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.21 $Y=3.33
+ $X2=6.085 $Y2=3.33
r126 64 66 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.21 $Y=3.33
+ $X2=6.48 $Y2=3.33
r127 63 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.86 $Y=3.33
+ $X2=6.985 $Y2=3.33
r128 63 66 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.86 $Y=3.33
+ $X2=6.48 $Y2=3.33
r129 62 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r130 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r131 58 59 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r132 55 59 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=4.08 $Y2=3.33
r133 54 58 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=4.08 $Y2=3.33
r134 54 55 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r135 51 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r136 51 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r137 49 61 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=5.14 $Y=3.33 $X2=5.04
+ $Y2=3.33
r138 49 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.14 $Y=3.33
+ $X2=5.225 $Y2=3.33
r139 47 58 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=4.16 $Y=3.33 $X2=4.08
+ $Y2=3.33
r140 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.16 $Y=3.33
+ $X2=4.325 $Y2=3.33
r141 46 61 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=4.49 $Y=3.33
+ $X2=5.04 $Y2=3.33
r142 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.49 $Y=3.33
+ $X2=4.325 $Y2=3.33
r143 42 45 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=8.89 $Y=1.985
+ $X2=8.89 $Y2=2.815
r144 40 83 3.1166 $w=2.5e-07 $l=1.07912e-07 $layer=LI1_cond $X=8.89 $Y=3.245
+ $X2=8.942 $Y2=3.33
r145 40 45 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.89 $Y=3.245
+ $X2=8.89 $Y2=2.815
r146 36 39 35.0343 $w=2.48e-07 $l=7.6e-07 $layer=LI1_cond $X=6.985 $Y=2.055
+ $X2=6.985 $Y2=2.815
r147 34 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.985 $Y=3.245
+ $X2=6.985 $Y2=3.33
r148 34 39 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6.985 $Y=3.245
+ $X2=6.985 $Y2=2.815
r149 30 33 35.0343 $w=2.48e-07 $l=7.6e-07 $layer=LI1_cond $X=6.085 $Y=2.055
+ $X2=6.085 $Y2=2.815
r150 28 77 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.085 $Y=3.245
+ $X2=6.085 $Y2=3.33
r151 28 33 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6.085 $Y=3.245
+ $X2=6.085 $Y2=2.815
r152 27 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.31 $Y=3.33
+ $X2=5.225 $Y2=3.33
r153 26 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.96 $Y=3.33
+ $X2=6.085 $Y2=3.33
r154 26 27 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.96 $Y=3.33
+ $X2=5.31 $Y2=3.33
r155 22 25 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=5.225 $Y=2.055
+ $X2=5.225 $Y2=2.815
r156 20 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=3.245
+ $X2=5.225 $Y2=3.33
r157 20 25 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=5.225 $Y=3.245
+ $X2=5.225 $Y2=2.815
r158 16 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.325 $Y=3.245
+ $X2=4.325 $Y2=3.33
r159 16 18 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=4.325 $Y=3.245
+ $X2=4.325 $Y2=2.485
r160 5 45 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.715
+ $Y=1.84 $X2=8.85 $Y2=2.815
r161 5 42 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.715
+ $Y=1.84 $X2=8.85 $Y2=1.985
r162 4 39 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.89
+ $Y=1.84 $X2=7.025 $Y2=2.815
r163 4 36 400 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=6.89
+ $Y=1.84 $X2=7.025 $Y2=2.055
r164 3 33 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.99
+ $Y=1.84 $X2=6.125 $Y2=2.815
r165 3 30 400 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=5.99
+ $Y=1.84 $X2=6.125 $Y2=2.055
r166 2 25 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.09
+ $Y=1.84 $X2=5.225 $Y2=2.815
r167 2 22 400 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=5.09
+ $Y=1.84 $X2=5.225 $Y2=2.055
r168 1 18 300 $w=1.7e-07 $l=7.09295e-07 $layer=licon1_PDIFF $count=2 $X=4.19
+ $Y=1.84 $X2=4.325 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_MS__EINVP_8%A_27_74# 1 2 3 4 5 6 7 8 9 30 32 33 34 36 38
+ 43 44 45 48 50 54 56 60 62 66 68 73 78 83 84 85
c172 85 0 1.07496e-19 $X=6.83 $Y=1.295
c173 83 0 1.07496e-19 $X=5.03 $Y=1.295
c174 45 0 5.65346e-20 $X=4.225 $Y=1.295
c175 36 0 8.60601e-20 $X=3.045 $Y=0.34
c176 34 0 8.60601e-20 $X=2.045 $Y=0.34
c177 32 0 8.60869e-20 $X=1.045 $Y=0.34
r178 78 81 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=3.21 $Y=0.34
+ $X2=3.21 $Y2=0.55
r179 73 76 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.21 $Y=0.34
+ $X2=2.21 $Y2=0.55
r180 68 71 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.21 $Y=0.34
+ $X2=1.21 $Y2=0.55
r181 64 66 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=7.76 $Y=1.21
+ $X2=7.76 $Y2=0.515
r182 63 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.955 $Y=1.295
+ $X2=6.83 $Y2=1.295
r183 62 64 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.635 $Y=1.295
+ $X2=7.76 $Y2=1.21
r184 62 63 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.635 $Y=1.295
+ $X2=6.955 $Y2=1.295
r185 58 85 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.83 $Y=1.21
+ $X2=6.83 $Y2=1.295
r186 58 60 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=6.83 $Y=1.21
+ $X2=6.83 $Y2=0.515
r187 57 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.015 $Y=1.295
+ $X2=5.93 $Y2=1.295
r188 56 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.705 $Y=1.295
+ $X2=6.83 $Y2=1.295
r189 56 57 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.705 $Y=1.295
+ $X2=6.015 $Y2=1.295
r190 52 84 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.93 $Y=1.21
+ $X2=5.93 $Y2=1.295
r191 52 54 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=5.93 $Y=1.21
+ $X2=5.93 $Y2=0.515
r192 51 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.155 $Y=1.295
+ $X2=5.03 $Y2=1.295
r193 50 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.845 $Y=1.295
+ $X2=5.93 $Y2=1.295
r194 50 51 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.845 $Y=1.295
+ $X2=5.155 $Y2=1.295
r195 46 83 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=1.21
+ $X2=5.03 $Y2=1.295
r196 46 48 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=5.03 $Y=1.21
+ $X2=5.03 $Y2=0.515
r197 44 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.905 $Y=1.295
+ $X2=5.03 $Y2=1.295
r198 44 45 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.905 $Y=1.295
+ $X2=4.225 $Y2=1.295
r199 41 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.14 $Y=1.21
+ $X2=4.225 $Y2=1.295
r200 41 43 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.14 $Y=1.21
+ $X2=4.14 $Y2=0.515
r201 40 43 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.14 $Y=0.425
+ $X2=4.14 $Y2=0.515
r202 39 78 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=0.34
+ $X2=3.21 $Y2=0.34
r203 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.055 $Y=0.34
+ $X2=4.14 $Y2=0.425
r204 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.055 $Y=0.34
+ $X2=3.375 $Y2=0.34
r205 37 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=0.34
+ $X2=2.21 $Y2=0.34
r206 36 78 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.045 $Y=0.34
+ $X2=3.21 $Y2=0.34
r207 36 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.045 $Y=0.34
+ $X2=2.375 $Y2=0.34
r208 35 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.34
+ $X2=1.21 $Y2=0.34
r209 34 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.045 $Y=0.34
+ $X2=2.21 $Y2=0.34
r210 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.045 $Y=0.34
+ $X2=1.375 $Y2=0.34
r211 32 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=1.21 $Y2=0.34
r212 32 33 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=0.445 $Y2=0.34
r213 28 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.425
+ $X2=0.445 $Y2=0.34
r214 28 30 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=0.28 $Y=0.425
+ $X2=0.28 $Y2=0.55
r215 9 66 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.58
+ $Y=0.37 $X2=7.72 $Y2=0.515
r216 8 60 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.65
+ $Y=0.37 $X2=6.79 $Y2=0.515
r217 7 54 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.79
+ $Y=0.37 $X2=5.93 $Y2=0.515
r218 6 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.93
+ $Y=0.37 $X2=5.07 $Y2=0.515
r219 5 43 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4 $Y=0.37
+ $X2=4.14 $Y2=0.515
r220 4 81 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=3
+ $Y=0.37 $X2=3.21 $Y2=0.55
r221 3 76 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=2
+ $Y=0.37 $X2=2.21 $Y2=0.55
r222 2 71 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.37 $X2=1.21 $Y2=0.55
r223 1 30 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_MS__EINVP_8%VGND 1 2 3 4 5 18 22 26 30 32 34 37 38 39 41
+ 49 58 62 68 71 74 78
c111 18 0 1.9142e-19 $X=4.57 $Y=0.515
r112 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r113 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r114 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r115 66 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r116 66 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.44
+ $Y2=0
r117 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r118 63 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.455 $Y=0 $X2=7.29
+ $Y2=0
r119 63 65 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=7.455 $Y=0 $X2=8.4
+ $Y2=0
r120 62 77 4.01281 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=8.675 $Y=0
+ $X2=8.897 $Y2=0
r121 62 65 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.675 $Y=0 $X2=8.4
+ $Y2=0
r122 61 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r123 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r124 58 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.125 $Y=0 $X2=7.29
+ $Y2=0
r125 58 60 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.125 $Y=0
+ $X2=6.96 $Y2=0
r126 57 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r127 57 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r128 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r129 54 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.665 $Y=0 $X2=5.5
+ $Y2=0
r130 54 56 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.665 $Y=0 $X2=6
+ $Y2=0
r131 53 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r132 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r133 50 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.735 $Y=0 $X2=4.57
+ $Y2=0
r134 50 52 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.735 $Y=0
+ $X2=5.04 $Y2=0
r135 49 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=0 $X2=5.5
+ $Y2=0
r136 49 52 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.335 $Y=0 $X2=5.04
+ $Y2=0
r137 47 48 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r138 44 48 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=4.08
+ $Y2=0
r139 43 47 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=4.08
+ $Y2=0
r140 43 44 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r141 41 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.405 $Y=0 $X2=4.57
+ $Y2=0
r142 41 47 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.405 $Y=0
+ $X2=4.08 $Y2=0
r143 39 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r144 39 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r145 39 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r146 37 56 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.195 $Y=0 $X2=6
+ $Y2=0
r147 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.195 $Y=0 $X2=6.36
+ $Y2=0
r148 36 60 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=6.525 $Y=0
+ $X2=6.96 $Y2=0
r149 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.525 $Y=0 $X2=6.36
+ $Y2=0
r150 32 77 3.19941 $w=2.6e-07 $l=1.27609e-07 $layer=LI1_cond $X=8.805 $Y=0.085
+ $X2=8.897 $Y2=0
r151 32 34 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=8.805 $Y=0.085
+ $X2=8.805 $Y2=0.505
r152 28 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.29 $Y=0.085
+ $X2=7.29 $Y2=0
r153 28 30 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.29 $Y=0.085
+ $X2=7.29 $Y2=0.515
r154 24 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.36 $Y=0.085
+ $X2=6.36 $Y2=0
r155 24 26 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.36 $Y=0.085
+ $X2=6.36 $Y2=0.515
r156 20 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.5 $Y=0.085 $X2=5.5
+ $Y2=0
r157 20 22 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.5 $Y=0.085
+ $X2=5.5 $Y2=0.515
r158 16 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.57 $Y=0.085
+ $X2=4.57 $Y2=0
r159 16 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.57 $Y=0.085
+ $X2=4.57 $Y2=0.515
r160 5 34 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=8.63
+ $Y=0.37 $X2=8.77 $Y2=0.505
r161 4 30 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=7.08
+ $Y=0.37 $X2=7.29 $Y2=0.515
r162 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.22
+ $Y=0.37 $X2=6.36 $Y2=0.515
r163 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.36
+ $Y=0.37 $X2=5.5 $Y2=0.515
r164 1 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.43
+ $Y=0.37 $X2=4.57 $Y2=0.515
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfrtn_1 CLK_N D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 VPWR a_859_347# a_1069_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X1 a_2492_424# a_1827_144# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X2 a_1273_131# a_859_347# a_1409_131# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 a_287_464# a_859_347# a_1273_131# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X4 a_2045_508# a_2087_410# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X5 a_324_81# D a_287_464# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X6 a_287_464# SCE a_538_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X7 VGND a_1273_131# a_1417_294# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_209_464# D a_287_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X9 a_474_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X10 a_859_347# CLK_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 VGND a_859_347# a_1069_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VPWR a_1273_131# a_1417_294# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X13 a_287_464# a_1069_74# a_1273_131# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X14 a_1827_144# a_1069_74# a_2073_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X15 VPWR RESET_B a_2087_410# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X16 a_27_88# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X17 a_859_347# CLK_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X18 a_1273_131# a_1069_74# a_1381_457# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X19 a_2492_424# a_1827_144# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X20 VPWR RESET_B a_1273_131# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X21 a_2265_74# a_1827_144# a_2087_410# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X22 VGND a_2492_424# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 a_1381_457# a_1417_294# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X24 VGND RESET_B a_2265_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X25 a_1409_131# a_1417_294# a_1483_131# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X26 a_1483_131# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X27 VPWR RESET_B a_287_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X28 a_1417_294# a_1069_74# a_1827_144# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X29 a_1417_294# a_859_347# a_1827_144# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X30 a_1827_144# a_859_347# a_2045_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X31 a_239_81# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X32 a_2087_410# a_1827_144# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X33 a_239_81# a_27_88# a_324_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X34 a_538_81# SCD a_239_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X35 a_27_88# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X36 VPWR a_2492_424# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X37 a_2073_74# a_2087_410# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X38 VPWR SCE a_209_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X39 a_287_464# a_27_88# a_474_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
.ends

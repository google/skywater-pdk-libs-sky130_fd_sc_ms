# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__dlxbn_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__dlxbn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.233700 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.440000 1.450000 0.815000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 0.850000 6.505000 1.130000 ;
        RECT 5.885000 1.130000 6.115000 1.800000 ;
        RECT 5.885000 1.800000 6.590000 2.070000 ;
        RECT 6.245000 0.355000 6.505000 0.850000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.225000 1.820000 8.555000 2.980000 ;
        RECT 8.245000 0.350000 8.495000 1.130000 ;
        RECT 8.325000 1.130000 8.495000 1.820000 ;
    END
  END Q_N
  PIN GATE_N
    ANTENNAGATEAREA  0.262200 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.695000 1.315000 2.150000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.100000  0.580000 2.845000 0.750000 ;
      RECT 0.100000  0.750000 0.445000 1.250000 ;
      RECT 0.100000  1.250000 0.270000 2.100000 ;
      RECT 0.100000  2.100000 0.445000 2.980000 ;
      RECT 0.625000  0.085000 0.955000 0.410000 ;
      RECT 0.650000  2.320000 0.980000 3.245000 ;
      RECT 1.135000  0.920000 1.465000 1.260000 ;
      RECT 1.135000  1.260000 1.885000 1.525000 ;
      RECT 1.150000  2.320000 1.655000 2.390000 ;
      RECT 1.150000  2.390000 4.275000 2.560000 ;
      RECT 1.150000  2.560000 1.485000 2.980000 ;
      RECT 1.485000  1.525000 1.655000 2.320000 ;
      RECT 1.695000  0.920000 2.225000 1.090000 ;
      RECT 1.825000  1.710000 3.385000 1.880000 ;
      RECT 1.825000  1.880000 2.155000 2.220000 ;
      RECT 2.055000  1.090000 2.225000 1.710000 ;
      RECT 2.285000  0.085000 2.640000 0.410000 ;
      RECT 2.360000  2.730000 2.690000 3.245000 ;
      RECT 2.515000  0.750000 2.845000 1.540000 ;
      RECT 3.015000  0.255000 4.265000 0.505000 ;
      RECT 3.015000  0.505000 3.185000 1.470000 ;
      RECT 3.015000  1.470000 3.385000 1.710000 ;
      RECT 3.230000  2.050000 3.935000 2.220000 ;
      RECT 3.355000  0.725000 4.070000 1.015000 ;
      RECT 3.355000  1.015000 5.315000 1.055000 ;
      RECT 3.555000  1.055000 5.315000 1.185000 ;
      RECT 3.555000  1.185000 3.725000 2.050000 ;
      RECT 3.895000  1.420000 4.275000 1.750000 ;
      RECT 4.105000  1.750000 4.275000 2.390000 ;
      RECT 4.445000  1.355000 4.775000 1.720000 ;
      RECT 4.445000  1.720000 5.655000 1.890000 ;
      RECT 4.630000  0.085000 5.015000 0.845000 ;
      RECT 4.670000  2.070000 5.080000 3.245000 ;
      RECT 4.985000  1.185000 5.315000 1.550000 ;
      RECT 5.185000  0.350000 5.655000 0.845000 ;
      RECT 5.250000  1.890000 5.655000 2.240000 ;
      RECT 5.250000  2.240000 6.955000 2.410000 ;
      RECT 5.250000  2.410000 5.655000 2.980000 ;
      RECT 5.485000  0.845000 5.655000 1.720000 ;
      RECT 5.825000  0.085000 6.075000 0.680000 ;
      RECT 5.890000  2.580000 6.140000 3.245000 ;
      RECT 6.285000  1.300000 6.955000 1.630000 ;
      RECT 6.675000  0.085000 7.005000 1.130000 ;
      RECT 6.710000  2.580000 7.040000 3.245000 ;
      RECT 6.785000  1.630000 6.955000 2.240000 ;
      RECT 7.185000  0.450000 7.515000 1.130000 ;
      RECT 7.215000  1.130000 7.515000 1.320000 ;
      RECT 7.215000  1.320000 8.155000 1.650000 ;
      RECT 7.215000  1.650000 7.545000 2.980000 ;
      RECT 7.745000  0.085000 8.075000 1.130000 ;
      RECT 7.775000  1.820000 8.025000 3.245000 ;
      RECT 8.675000  0.085000 9.005000 1.130000 ;
      RECT 8.755000  1.820000 9.005000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_ms__dlxbn_2
END LIBRARY

* File: sky130_fd_sc_ms__dlrtp_4.spice
* Created: Wed Sep  2 12:05:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dlrtp_4.pex.spice"
.subckt sky130_fd_sc_ms__dlrtp_4  VNB VPB D GATE RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_D_M1017_g N_A_27_126#_M1017_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.165874 AS=0.15675 PD=1.09574 PS=1.67 NRD=29.448 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.9 A=0.0825 P=1.4 MULT=1
MM1005 N_A_243_394#_M1005_d N_GATE_M1005_g N_VGND_M1017_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.223176 PD=2.05 PS=1.47426 NRD=0 NRS=21.072 M=1 R=4.93333
+ SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1021_d N_A_243_394#_M1021_g N_A_364_120#_M1021_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.160253 AS=0.2294 PD=1.43174 PS=2.1 NRD=26.196 NRS=2.424 M=1
+ R=4.93333 SA=75000.2 SB=75001 A=0.111 P=1.78 MULT=1
MM1002 A_559_74# N_A_27_126#_M1002_g N_VGND_M1021_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0816 AS=0.138597 PD=0.895 PS=1.23826 NRD=13.584 NRS=0.936 M=1 R=4.26667
+ SA=75000.6 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1026 N_A_640_74#_M1026_d N_A_364_120#_M1026_g A_559_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.154264 AS=0.0816 PD=1.28604 PS=0.895 NRD=5.616 NRS=13.584 M=1
+ R=4.26667 SA=75001 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1003 A_755_74# N_A_243_394#_M1003_g N_A_640_74#_M1026_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.101236 PD=0.63 PS=0.843962 NRD=14.28 NRS=34.284 M=1
+ R=2.8 SA=75001.4 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_A_797_48#_M1023_g A_755_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_A_938_74#_M1001_d N_A_640_74#_M1001_g N_A_797_48#_M1001_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.0912 PD=1.85 PS=0.925 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1007 N_A_938_74#_M1007_d N_A_640_74#_M1007_g N_A_797_48#_M1001_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0912 PD=0.92 PS=0.925 NRD=0 NRS=0.936 M=1
+ R=4.26667 SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1018 N_VGND_M1018_d N_RESET_B_M1018_g N_A_938_74#_M1007_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1028 N_VGND_M1018_d N_RESET_B_M1028_g N_A_938_74#_M1028_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1009 N_Q_M1009_d N_A_797_48#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1010 N_Q_M1009_d N_A_797_48#_M1010_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1020 N_Q_M1020_d N_A_797_48#_M1020_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1029 N_Q_M1020_d N_A_797_48#_M1029_g N_VGND_M1029_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_D_M1000_g N_A_27_126#_M1000_s VPB PSHORT L=0.18 W=0.84
+ AD=0.21525 AS=0.2352 PD=1.49 PS=2.24 NRD=47.1815 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90000.9 A=0.1512 P=2.04 MULT=1
MM1016 N_A_243_394#_M1016_d N_GATE_M1016_g N_VPWR_M1000_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2814 AS=0.21525 PD=2.35 PS=1.49 NRD=0 NRS=47.1815 M=1 R=4.66667
+ SA=90000.8 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1006 N_VPWR_M1006_d N_A_243_394#_M1006_g N_A_364_120#_M1006_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.161152 AS=0.2352 PD=1.2463 PS=2.24 NRD=19.9167 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90002.2 A=0.1512 P=2.04 MULT=1
MM1027 A_565_392# N_A_27_126#_M1027_g N_VPWR_M1006_d VPB PSHORT L=0.18 W=1
+ AD=0.105 AS=0.191848 PD=1.21 PS=1.4837 NRD=9.8303 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1015 N_A_640_74#_M1015_d N_A_243_394#_M1015_g A_565_392# VPB PSHORT L=0.18 W=1
+ AD=0.219366 AS=0.105 PD=1.90845 PS=1.21 NRD=0 NRS=9.8303 M=1 R=5.55556
+ SA=90001 SB=90001.3 A=0.18 P=2.36 MULT=1
MM1025 A_750_508# N_A_364_120#_M1025_g N_A_640_74#_M1015_d VPB PSHORT L=0.18
+ W=0.42 AD=0.09345 AS=0.0921338 PD=0.865 PS=0.801549 NRD=78.5636 NRS=39.8531
+ M=1 R=2.33333 SA=90001.5 SB=90002.4 A=0.0756 P=1.2 MULT=1
MM1014 N_VPWR_M1014_d N_A_797_48#_M1014_g A_750_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.133233 AS=0.09345 PD=1.13667 PS=0.865 NRD=51.5943 NRS=78.5636 M=1
+ R=2.33333 SA=90002.1 SB=90001.8 A=0.0756 P=1.2 MULT=1
MM1008 N_A_797_48#_M1008_d N_A_640_74#_M1008_g N_VPWR_M1014_d VPB PSHORT L=0.18
+ W=0.84 AD=0.1134 AS=0.266467 PD=1.11 PS=2.27333 NRD=0 NRS=61.4837 M=1
+ R=4.66667 SA=90000.6 SB=90003.7 A=0.1512 P=2.04 MULT=1
MM1012 N_A_797_48#_M1008_d N_A_640_74#_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1134 AS=0.1344 PD=1.11 PS=1.16 NRD=0 NRS=10.5395 M=1 R=4.66667
+ SA=90001.1 SB=90003.2 A=0.1512 P=2.04 MULT=1
MM1011 N_VPWR_M1012_s N_RESET_B_M1011_g N_A_797_48#_M1011_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1344 AS=0.1344 PD=1.16 PS=1.16 NRD=0 NRS=10.5395 M=1 R=4.66667
+ SA=90001.6 SB=90002.7 A=0.1512 P=2.04 MULT=1
MM1013 N_VPWR_M1013_d N_RESET_B_M1013_g N_A_797_48#_M1011_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1614 AS=0.1344 PD=1.26429 PS=1.16 NRD=18.7544 NRS=0 M=1 R=4.66667
+ SA=90002.1 SB=90002.2 A=0.1512 P=2.04 MULT=1
MM1004 N_VPWR_M1013_d N_A_797_48#_M1004_g N_Q_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2152 AS=0.1512 PD=1.68571 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1019 N_VPWR_M1019_d N_A_797_48#_M1019_g N_Q_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90002.5
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1022 N_VPWR_M1019_d N_A_797_48#_M1022_g N_Q_M1022_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1904 PD=1.44 PS=1.46 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1024 N_VPWR_M1024_d N_A_797_48#_M1024_g N_Q_M1022_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3472 AS=0.1904 PD=2.86 PS=1.46 NRD=4.3931 NRS=2.6201 M=1 R=6.22222
+ SA=90003.5 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX30_noxref VNB VPB NWDIODE A=17.5032 P=22.96
c_1074 A_565_392# 0 1.67587e-19 $X=2.825 $Y=1.96
c_1277 A_559_74# 0 5.47968e-20 $X=2.795 $Y=0.37
*
.include "sky130_fd_sc_ms__dlrtp_4.pxi.spice"
*
.ends
*
*

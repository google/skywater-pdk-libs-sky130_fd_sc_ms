* File: sky130_fd_sc_ms__o311a_4.pex.spice
* Created: Wed Sep  2 12:25:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O311A_4%A_83_244# 1 2 3 4 15 17 19 22 24 26 29 31 33
+ 36 38 40 41 46 47 48 49 52 54 58 60 62 65 69 75 77 81 94
c187 94 0 1.56333e-19 $X=2.19 $Y=1.385
c188 58 0 1.72297e-19 $X=4.255 $Y=2.815
c189 54 0 9.87938e-21 $X=4.09 $Y=2.035
c190 24 0 4.74979e-20 $X=0.995 $Y=1.22
c191 22 0 5.8386e-20 $X=0.955 $Y=2.4
c192 15 0 7.10079e-20 $X=0.505 $Y=2.4
r193 91 92 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=1.69 $Y=1.385
+ $X2=2.09 $Y2=1.385
r194 90 91 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=1.455 $Y=1.385
+ $X2=1.69 $Y2=1.385
r195 87 88 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=0.955 $Y=1.385
+ $X2=0.995 $Y2=1.385
r196 86 87 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=0.565 $Y=1.385
+ $X2=0.955 $Y2=1.385
r197 84 86 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=0.505 $Y=1.385
+ $X2=0.565 $Y2=1.385
r198 81 83 16.7345 $w=2.26e-07 $l=3.1e-07 $layer=LI1_cond $X=5.615 $Y=2.075
+ $X2=5.925 $Y2=2.075
r199 77 79 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=4.46 $Y=1.1
+ $X2=4.46 $Y2=1.215
r200 71 73 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=2.82 $Y=2.035
+ $X2=2.82 $Y2=2.105
r201 69 71 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.82 $Y=1.805
+ $X2=2.82 $Y2=2.035
r202 68 94 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.1 $Y=1.385 $X2=2.19
+ $Y2=1.385
r203 68 92 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=2.1 $Y=1.385 $X2=2.09
+ $Y2=1.385
r204 67 68 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.1
+ $Y=1.385 $X2=2.1 $Y2=1.385
r205 65 81 2.4068 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.615 $Y=1.95
+ $X2=5.615 $Y2=2.075
r206 64 65 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.615 $Y=1.3
+ $X2=5.615 $Y2=1.95
r207 63 79 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.585 $Y=1.215
+ $X2=4.46 $Y2=1.215
r208 62 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.53 $Y=1.215
+ $X2=5.615 $Y2=1.3
r209 62 63 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=5.53 $Y=1.215
+ $X2=4.585 $Y2=1.215
r210 61 75 8.61065 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=4.42 $Y=2.055
+ $X2=4.255 $Y2=2.04
r211 60 81 5.36542 $w=2.26e-07 $l=9.44722e-08 $layer=LI1_cond $X=5.53 $Y=2.055
+ $X2=5.615 $Y2=2.075
r212 60 61 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=5.53 $Y=2.055
+ $X2=4.42 $Y2=2.055
r213 56 75 0.89609 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=4.255 $Y=2.14
+ $X2=4.255 $Y2=2.04
r214 56 58 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.255 $Y=2.14
+ $X2=4.255 $Y2=2.815
r215 55 71 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.985 $Y=2.035
+ $X2=2.82 $Y2=2.035
r216 54 75 8.61065 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=4.09 $Y=2.035
+ $X2=4.255 $Y2=2.04
r217 54 55 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=4.09 $Y=2.035
+ $X2=2.985 $Y2=2.035
r218 50 73 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.82 $Y=2.12
+ $X2=2.82 $Y2=2.105
r219 50 52 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.82 $Y=2.12
+ $X2=2.82 $Y2=2.815
r220 48 69 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=1.805
+ $X2=2.82 $Y2=1.805
r221 48 49 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.655 $Y=1.805
+ $X2=2.265 $Y2=1.805
r222 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.18 $Y=1.72
+ $X2=2.265 $Y2=1.805
r223 46 67 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.18 $Y=1.55
+ $X2=2.18 $Y2=1.385
r224 46 47 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.18 $Y=1.55
+ $X2=2.18 $Y2=1.72
r225 44 90 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=1.42 $Y=1.385
+ $X2=1.455 $Y2=1.385
r226 44 88 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=1.42 $Y=1.385
+ $X2=0.995 $Y2=1.385
r227 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.42
+ $Y=1.385 $X2=1.42 $Y2=1.385
r228 41 67 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.095 $Y=1.385
+ $X2=2.18 $Y2=1.385
r229 41 43 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.095 $Y=1.385
+ $X2=1.42 $Y2=1.385
r230 38 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.19 $Y=1.22
+ $X2=2.19 $Y2=1.385
r231 38 40 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.19 $Y=1.22
+ $X2=2.19 $Y2=0.74
r232 34 92 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.09 $Y=1.55
+ $X2=2.09 $Y2=1.385
r233 34 36 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.09 $Y=1.55
+ $X2=2.09 $Y2=2.4
r234 31 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.22
+ $X2=1.69 $Y2=1.385
r235 31 33 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.69 $Y=1.22
+ $X2=1.69 $Y2=0.74
r236 27 90 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.455 $Y=1.55
+ $X2=1.455 $Y2=1.385
r237 27 29 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.455 $Y=1.55
+ $X2=1.455 $Y2=2.4
r238 24 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.22
+ $X2=0.995 $Y2=1.385
r239 24 26 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.995 $Y=1.22
+ $X2=0.995 $Y2=0.74
r240 20 87 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.55
+ $X2=0.955 $Y2=1.385
r241 20 22 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.955 $Y=1.55
+ $X2=0.955 $Y2=2.4
r242 17 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=1.22
+ $X2=0.565 $Y2=1.385
r243 17 19 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.565 $Y=1.22
+ $X2=0.565 $Y2=0.74
r244 13 84 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.55
+ $X2=0.505 $Y2=1.385
r245 13 15 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.505 $Y=1.55
+ $X2=0.505 $Y2=2.4
r246 4 83 600 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=5.78
+ $Y=1.96 $X2=5.925 $Y2=2.115
r247 3 75 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.12
+ $Y=1.96 $X2=4.255 $Y2=2.105
r248 3 58 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.12
+ $Y=1.96 $X2=4.255 $Y2=2.815
r249 2 73 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.685
+ $Y=1.96 $X2=2.82 $Y2=2.105
r250 2 52 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.685
+ $Y=1.96 $X2=2.82 $Y2=2.815
r251 1 77 182 $w=1.7e-07 $l=8.12588e-07 $layer=licon1_NDIFF $count=1 $X=4.2
+ $Y=0.39 $X2=4.42 $Y2=1.1
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_4%B1 3 5 9 11 13 14 15 18 20 21 23 25 30 32 37
+ 38 43
c103 23 0 1.03664e-19 $X=4.08 $Y=1.47
c104 11 0 1.72297e-19 $X=4.53 $Y=1.86
c105 3 0 9.87938e-21 $X=2.595 $Y=2.46
r106 37 40 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=5.195 $Y=1.635
+ $X2=5.195 $Y2=1.785
r107 37 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.195 $Y=1.635
+ $X2=5.195 $Y2=1.47
r108 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.195
+ $Y=1.635 $X2=5.195 $Y2=1.635
r109 30 38 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=5.04 $Y=1.635
+ $X2=5.195 $Y2=1.635
r110 30 43 6.71605 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=5.04 $Y=1.635
+ $X2=4.925 $Y2=1.635
r111 29 35 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.385
+ $X2=2.67 $Y2=1.55
r112 29 32 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.67 $Y=1.385
+ $X2=2.67 $Y2=1.295
r113 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.385 $X2=2.67 $Y2=1.385
r114 25 43 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=4.165 $Y=1.555
+ $X2=4.925 $Y2=1.555
r115 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.08 $Y=1.47
+ $X2=4.165 $Y2=1.555
r116 22 23 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.08 $Y=1.265
+ $X2=4.08 $Y2=1.47
r117 21 28 7.35588 $w=3.4e-07 $l=2.89206e-07 $layer=LI1_cond $X=2.91 $Y=1.18
+ $X2=2.707 $Y2=1.385
r118 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.995 $Y=1.18
+ $X2=4.08 $Y2=1.265
r119 20 21 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=3.995 $Y=1.18
+ $X2=2.91 $Y2=1.18
r120 18 39 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=5.145 $Y=0.71
+ $X2=5.145 $Y2=1.47
r121 14 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.03 $Y=1.785
+ $X2=5.195 $Y2=1.785
r122 14 15 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=5.03 $Y=1.785
+ $X2=4.62 $Y2=1.785
r123 11 15 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.53 $Y=1.86
+ $X2=4.62 $Y2=1.785
r124 11 13 160.667 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=4.53 $Y=1.86 $X2=4.53
+ $Y2=2.46
r125 7 9 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=3.18 $Y=1.22 $X2=3.18
+ $Y2=0.71
r126 6 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=1.295
+ $X2=2.67 $Y2=1.295
r127 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.105 $Y=1.295
+ $X2=3.18 $Y2=1.22
r128 5 6 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.105 $Y=1.295
+ $X2=2.835 $Y2=1.295
r129 3 35 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=2.595 $Y=2.46
+ $X2=2.595 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_4%C1 3 6 9 13 15 19 21 26 29
c71 19 0 1.03664e-19 $X=4.715 $Y=0.71
r72 24 27 46.242 $w=4.45e-07 $l=3.7e-07 $layer=POLY_cond $X=3.66 $Y=1.542
+ $X2=4.03 $Y2=1.542
r73 24 26 46.8028 $w=4.45e-07 $l=1.65e-07 $layer=POLY_cond $X=3.66 $Y=1.542
+ $X2=3.495 $Y2=1.542
r74 21 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.66
+ $Y=1.6 $X2=3.66 $Y2=1.6
r75 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.715 $Y=1.32
+ $X2=4.715 $Y2=0.71
r76 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.64 $Y=1.395
+ $X2=4.715 $Y2=1.32
r77 15 29 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=4.64 $Y=1.395
+ $X2=4.2 $Y2=1.395
r78 11 29 35.5547 $w=4.45e-07 $l=7.5e-08 $layer=POLY_cond $X=4.125 $Y=1.542
+ $X2=4.2 $Y2=1.542
r79 11 27 11.8729 $w=4.45e-07 $l=9.5e-08 $layer=POLY_cond $X=4.125 $Y=1.542
+ $X2=4.03 $Y2=1.542
r80 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.125 $Y=1.32
+ $X2=4.125 $Y2=0.71
r81 7 27 24.0211 $w=1.8e-07 $l=2.23e-07 $layer=POLY_cond $X=4.03 $Y=1.765
+ $X2=4.03 $Y2=1.542
r82 7 9 270.153 $w=1.8e-07 $l=6.95e-07 $layer=POLY_cond $X=4.03 $Y=1.765
+ $X2=4.03 $Y2=2.46
r83 6 26 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.255 $Y=1.69
+ $X2=3.495 $Y2=1.69
r84 1 6 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.165 $Y=1.765
+ $X2=3.255 $Y2=1.69
r85 1 3 270.153 $w=1.8e-07 $l=6.95e-07 $layer=POLY_cond $X=3.165 $Y=1.765
+ $X2=3.165 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_4%A3 3 7 11 15 17 24
c58 17 0 1.46209e-19 $X=6 $Y=1.665
r59 24 25 7.53125 $w=3.2e-07 $l=5e-08 $layer=POLY_cond $X=6.16 $Y=1.585 $X2=6.21
+ $Y2=1.585
r60 22 24 18.8281 $w=3.2e-07 $l=1.25e-07 $layer=POLY_cond $X=6.035 $Y=1.585
+ $X2=6.16 $Y2=1.585
r61 20 22 51.9656 $w=3.2e-07 $l=3.45e-07 $layer=POLY_cond $X=5.69 $Y=1.585
+ $X2=6.035 $Y2=1.585
r62 19 20 2.25938 $w=3.2e-07 $l=1.5e-08 $layer=POLY_cond $X=5.675 $Y=1.585
+ $X2=5.69 $Y2=1.585
r63 17 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.035
+ $Y=1.585 $X2=6.035 $Y2=1.585
r64 13 25 20.4921 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.21 $Y=1.42
+ $X2=6.21 $Y2=1.585
r65 13 15 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.21 $Y=1.42
+ $X2=6.21 $Y2=0.71
r66 9 24 16.2157 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.16 $Y=1.75
+ $X2=6.16 $Y2=1.585
r67 9 11 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=6.16 $Y=1.75 $X2=6.16
+ $Y2=2.46
r68 5 20 16.2157 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.69 $Y=1.75
+ $X2=5.69 $Y2=1.585
r69 5 7 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=5.69 $Y=1.75 $X2=5.69
+ $Y2=2.46
r70 1 19 20.4921 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.675 $Y=1.42
+ $X2=5.675 $Y2=1.585
r71 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.675 $Y=1.42
+ $X2=5.675 $Y2=0.71
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_4%A2 3 7 11 13 15 16 17 21 22 23 31 35
c75 21 0 2.29863e-19 $X=6.69 $Y=1.385
c76 11 0 1.43398e-19 $X=8.105 $Y=2.46
r77 31 33 31.7105 $w=3.42e-07 $l=2.25e-07 $layer=POLY_cond $X=8.145 $Y=1.35
+ $X2=8.37 $Y2=1.35
r78 30 31 5.63743 $w=3.42e-07 $l=4e-08 $layer=POLY_cond $X=8.105 $Y=1.35
+ $X2=8.145 $Y2=1.35
r79 22 35 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.37 $Y=1.215 $X2=8.37
+ $Y2=1.3
r80 22 23 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=8.37 $Y=1.305
+ $X2=8.37 $Y2=1.665
r81 22 35 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=8.37 $Y=1.305
+ $X2=8.37 $Y2=1.3
r82 22 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.37
+ $Y=1.305 $X2=8.37 $Y2=1.305
r83 21 29 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.69 $Y=1.385
+ $X2=6.69 $Y2=1.55
r84 21 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.69 $Y=1.385
+ $X2=6.69 $Y2=1.22
r85 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.69
+ $Y=1.385 $X2=6.69 $Y2=1.385
r86 17 20 5.7933 $w=3.58e-07 $l=2.77263e-07 $layer=LI1_cond $X=6.935 $Y=1.215
+ $X2=6.73 $Y2=1.385
r87 16 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.205 $Y=1.215
+ $X2=8.37 $Y2=1.215
r88 16 17 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=8.205 $Y=1.215
+ $X2=6.935 $Y2=1.215
r89 13 31 22.0749 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=8.145 $Y=1.14
+ $X2=8.145 $Y2=1.35
r90 13 15 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.145 $Y=1.14
+ $X2=8.145 $Y2=0.71
r91 9 30 17.7656 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=8.105 $Y=1.56
+ $X2=8.105 $Y2=1.35
r92 9 11 349.839 $w=1.8e-07 $l=9e-07 $layer=POLY_cond $X=8.105 $Y=1.56 $X2=8.105
+ $Y2=2.46
r93 7 28 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=6.645 $Y=0.71
+ $X2=6.645 $Y2=1.22
r94 3 29 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=6.615 $Y=2.46
+ $X2=6.615 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_4%A1 3 7 11 15 17 18 28
c54 18 0 8.3654e-20 $X=7.92 $Y=1.665
r55 27 28 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=7.635 $Y=1.635
+ $X2=7.7 $Y2=1.635
r56 25 27 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=7.61 $Y=1.635
+ $X2=7.635 $Y2=1.635
r57 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.61
+ $Y=1.635 $X2=7.61 $Y2=1.635
r58 23 25 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=7.185 $Y=1.635
+ $X2=7.61 $Y2=1.635
r59 21 23 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.17 $Y=1.635
+ $X2=7.185 $Y2=1.635
r60 18 26 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=7.92 $Y=1.635
+ $X2=7.61 $Y2=1.635
r61 17 26 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.44 $Y=1.635
+ $X2=7.61 $Y2=1.635
r62 13 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.7 $Y=1.47 $X2=7.7
+ $Y2=1.635
r63 13 15 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=7.7 $Y=1.47 $X2=7.7
+ $Y2=0.71
r64 9 27 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.635 $Y=1.8
+ $X2=7.635 $Y2=1.635
r65 9 11 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=7.635 $Y=1.8
+ $X2=7.635 $Y2=2.46
r66 5 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.185 $Y=1.8
+ $X2=7.185 $Y2=1.635
r67 5 7 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=7.185 $Y=1.8 $X2=7.185
+ $Y2=2.46
r68 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.17 $Y=1.47
+ $X2=7.17 $Y2=1.635
r69 1 3 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=7.17 $Y=1.47 $X2=7.17
+ $Y2=0.71
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_4%VPWR 1 2 3 4 5 6 19 21 27 31 35 41 43 44 49
+ 54 55 56 57 58 60 65 78 79 85 88 91
c126 49 0 1.43398e-19 $X=7.41 $Y=2.18
r127 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r128 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r129 86 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r130 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r131 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r132 78 79 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r133 76 79 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=8.4 $Y2=3.33
r134 75 78 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=8.4 $Y2=3.33
r135 75 76 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r136 73 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r137 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r138 70 91 13.6095 $w=1.7e-07 $l=3.48e-07 $layer=LI1_cond $X=3.92 $Y=3.33
+ $X2=3.572 $Y2=3.33
r139 70 72 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.92 $Y=3.33
+ $X2=4.56 $Y2=3.33
r140 69 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r141 69 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r142 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r143 66 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.48 $Y=3.33
+ $X2=2.315 $Y2=3.33
r144 66 68 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.48 $Y=3.33
+ $X2=3.12 $Y2=3.33
r145 65 91 13.6095 $w=1.7e-07 $l=3.47e-07 $layer=LI1_cond $X=3.225 $Y=3.33
+ $X2=3.572 $Y2=3.33
r146 65 68 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.225 $Y=3.33
+ $X2=3.12 $Y2=3.33
r147 64 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r148 64 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r149 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r150 61 82 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r151 61 63 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r152 60 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.23 $Y2=3.33
r153 60 63 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.72 $Y2=3.33
r154 58 73 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r155 58 92 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=3.6 $Y2=3.33
r156 56 57 8.89604 $w=4.23e-07 $l=1.7e-07 $layer=LI1_cond $X=6.38 $Y=2.255
+ $X2=6.55 $Y2=2.255
r157 54 72 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=4.59 $Y=3.33 $X2=4.56
+ $Y2=3.33
r158 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.59 $Y=3.33
+ $X2=4.755 $Y2=3.33
r159 53 75 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.92 $Y=3.33
+ $X2=5.04 $Y2=3.33
r160 53 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.92 $Y=3.33
+ $X2=4.755 $Y2=3.33
r161 49 57 23.32 $w=4.23e-07 $l=8.6e-07 $layer=LI1_cond $X=7.41 $Y=2.182
+ $X2=6.55 $Y2=2.182
r162 46 52 4.88517 $w=1.7e-07 $l=1.79374e-07 $layer=LI1_cond $X=4.92 $Y=2.455
+ $X2=4.755 $Y2=2.425
r163 46 56 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=4.92 $Y=2.455
+ $X2=6.38 $Y2=2.455
r164 44 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.755 $Y=3.245
+ $X2=4.755 $Y2=3.33
r165 43 52 2.881 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=4.755 $Y=2.54
+ $X2=4.755 $Y2=2.425
r166 43 44 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=4.755 $Y=2.54
+ $X2=4.755 $Y2=3.245
r167 39 91 2.84707 $w=6.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.572 $Y=3.245
+ $X2=3.572 $Y2=3.33
r168 39 41 13.5957 $w=6.93e-07 $l=7.9e-07 $layer=LI1_cond $X=3.572 $Y=3.245
+ $X2=3.572 $Y2=2.455
r169 35 38 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.315 $Y=2.145
+ $X2=2.315 $Y2=2.825
r170 33 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.315 $Y=3.245
+ $X2=2.315 $Y2=3.33
r171 33 38 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=2.315 $Y=3.245
+ $X2=2.315 $Y2=2.825
r172 32 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.23 $Y2=3.33
r173 31 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.15 $Y=3.33
+ $X2=2.315 $Y2=3.33
r174 31 32 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.15 $Y=3.33
+ $X2=1.395 $Y2=3.33
r175 27 30 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.23 $Y=2.145
+ $X2=1.23 $Y2=2.825
r176 25 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=3.33
r177 25 30 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=2.825
r178 21 24 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r179 19 82 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r180 19 24 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r181 6 49 600 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_PDIFF $count=1 $X=7.275
+ $Y=1.96 $X2=7.41 $Y2=2.18
r182 5 52 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.62
+ $Y=1.96 $X2=4.755 $Y2=2.475
r183 4 41 150 $w=1.7e-07 $l=7.58123e-07 $layer=licon1_PDIFF $count=4 $X=3.255
+ $Y=1.96 $X2=3.805 $Y2=2.455
r184 3 38 400 $w=1.7e-07 $l=1.05033e-06 $layer=licon1_PDIFF $count=1 $X=2.18
+ $Y=1.84 $X2=2.315 $Y2=2.825
r185 3 35 400 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_PDIFF $count=1 $X=2.18
+ $Y=1.84 $X2=2.315 $Y2=2.145
r186 2 30 400 $w=1.7e-07 $l=1.07352e-06 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.23 $Y2=2.825
r187 2 27 400 $w=1.7e-07 $l=3.86588e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.23 $Y2=2.145
r188 1 24 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r189 1 21 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_4%X 1 2 3 4 13 15 16 19 25 27 29 33 39 42 45
+ 48 51
c70 27 0 7.10079e-20 $X=1.565 $Y=1.805
c71 15 0 5.8386e-20 $X=0.565 $Y=1.565
c72 13 0 4.74979e-20 $X=0.615 $Y=1.225
r73 48 51 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=1.225 $X2=0.24
+ $Y2=1.31
r74 48 51 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.24 $Y=1.345
+ $X2=0.24 $Y2=1.31
r75 45 46 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=0.78 $Y=0.965
+ $X2=0.78 $Y2=1.225
r76 42 44 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.73 $Y=1.565
+ $X2=0.73 $Y2=1.805
r77 41 48 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.24 $Y=1.48
+ $X2=0.24 $Y2=1.345
r78 37 39 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.905 $Y=0.88
+ $X2=1.905 $Y2=0.515
r79 33 35 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.73 $Y=1.985
+ $X2=1.73 $Y2=2.815
r80 31 33 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.73 $Y=1.89
+ $X2=1.73 $Y2=1.985
r81 30 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0.965
+ $X2=0.78 $Y2=0.965
r82 29 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.74 $Y=0.965
+ $X2=1.905 $Y2=0.88
r83 29 30 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=1.74 $Y=0.965
+ $X2=0.945 $Y2=0.965
r84 28 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=1.805
+ $X2=0.73 $Y2=1.805
r85 27 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.565 $Y=1.805
+ $X2=1.73 $Y2=1.89
r86 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.565 $Y=1.805
+ $X2=0.895 $Y2=1.805
r87 23 45 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.88
+ $X2=0.78 $Y2=0.965
r88 23 25 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.78 $Y=0.88
+ $X2=0.78 $Y2=0.515
r89 19 21 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.73 $Y=1.985
+ $X2=0.73 $Y2=2.815
r90 17 44 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.89
+ $X2=0.73 $Y2=1.805
r91 17 19 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.73 $Y=1.89
+ $X2=0.73 $Y2=1.985
r92 16 41 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.565
+ $X2=0.24 $Y2=1.48
r93 15 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=1.565
+ $X2=0.73 $Y2=1.565
r94 15 16 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.565 $Y=1.565
+ $X2=0.355 $Y2=1.565
r95 14 48 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.355 $Y=1.225
+ $X2=0.24 $Y2=1.225
r96 13 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=1.225
+ $X2=0.78 $Y2=1.225
r97 13 14 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.615 $Y=1.225
+ $X2=0.355 $Y2=1.225
r98 4 35 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.84 $X2=1.73 $Y2=2.815
r99 4 33 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.84 $X2=1.73 $Y2=1.985
r100 3 21 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.815
r101 3 19 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=1.985
r102 2 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.765
+ $Y=0.37 $X2=1.905 $Y2=0.515
r103 1 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.64
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_4%A_1034_392# 1 2 3 14 18 24 25
r38 23 25 8.52431 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=6.385 $Y=2.892
+ $X2=6.55 $Y2=2.892
r39 23 24 6.36223 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=6.385 $Y=2.892
+ $X2=6.22 $Y2=2.892
r40 18 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=8.36 $Y=2.135
+ $X2=8.36 $Y2=2.815
r41 16 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=8.36 $Y=2.905 $X2=8.36
+ $Y2=2.815
r42 14 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.195 $Y=2.99
+ $X2=8.36 $Y2=2.905
r43 14 25 107.321 $w=1.68e-07 $l=1.645e-06 $layer=LI1_cond $X=8.195 $Y=2.99
+ $X2=6.55 $Y2=2.99
r44 12 24 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=5.39 $Y=2.835
+ $X2=6.22 $Y2=2.835
r45 3 21 400 $w=1.7e-07 $l=9.33863e-07 $layer=licon1_PDIFF $count=1 $X=8.195
+ $Y=1.96 $X2=8.36 $Y2=2.815
r46 3 18 400 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_PDIFF $count=1 $X=8.195
+ $Y=1.96 $X2=8.36 $Y2=2.135
r47 2 23 600 $w=1.7e-07 $l=9.1e-07 $layer=licon1_PDIFF $count=1 $X=6.25 $Y=1.96
+ $X2=6.385 $Y2=2.805
r48 1 12 600 $w=1.7e-07 $l=9.38576e-07 $layer=licon1_PDIFF $count=1 $X=5.17
+ $Y=1.96 $X2=5.39 $Y2=2.795
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_4%A_1341_392# 1 2 7 13
r13 11 13 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.9 $Y=2.565 $X2=7.9
+ $Y2=2.135
r14 7 11 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.775 $Y=2.65
+ $X2=7.9 $Y2=2.565
r15 7 9 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=7.775 $Y=2.65
+ $X2=6.92 $Y2=2.65
r16 2 13 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=7.725
+ $Y=1.96 $X2=7.86 $Y2=2.135
r17 1 9 600 $w=1.7e-07 $l=7.90221e-07 $layer=licon1_PDIFF $count=1 $X=6.705
+ $Y=1.96 $X2=6.92 $Y2=2.65
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_4%VGND 1 2 3 4 5 6 19 21 25 29 33 37 41 44 45
+ 46 48 57 64 69 76 77 83 86 89 92
c99 21 0 1.56333e-19 $X=0.35 $Y=0.515
r100 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r101 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r102 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r103 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r104 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r105 77 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r106 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r107 74 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.095 $Y=0 $X2=7.93
+ $Y2=0
r108 74 76 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.095 $Y=0 $X2=8.4
+ $Y2=0
r109 73 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r110 73 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r111 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r112 70 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.095 $Y=0 $X2=6.93
+ $Y2=0
r113 70 72 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.095 $Y=0 $X2=7.44
+ $Y2=0
r114 69 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.765 $Y=0 $X2=7.93
+ $Y2=0
r115 69 72 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.765 $Y=0
+ $X2=7.44 $Y2=0
r116 68 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r117 68 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r118 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r119 65 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.095 $Y=0 $X2=5.93
+ $Y2=0
r120 65 67 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.095 $Y=0
+ $X2=6.48 $Y2=0
r121 64 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.765 $Y=0 $X2=6.93
+ $Y2=0
r122 64 67 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.765 $Y=0
+ $X2=6.48 $Y2=0
r123 63 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r124 62 63 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r125 59 62 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=5.52
+ $Y2=0
r126 59 60 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r127 57 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.765 $Y=0 $X2=5.93
+ $Y2=0
r128 57 62 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.765 $Y=0 $X2=5.52
+ $Y2=0
r129 56 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r130 56 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r131 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r132 53 83 10.6558 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=1.57 $Y=0 $X2=1.342
+ $Y2=0
r133 53 55 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.57 $Y=0 $X2=2.16
+ $Y2=0
r134 52 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r135 52 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r136 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r137 49 80 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r138 49 51 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r139 48 83 10.6558 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=1.115 $Y=0
+ $X2=1.342 $Y2=0
r140 48 51 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=0
+ $X2=0.72 $Y2=0
r141 46 63 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.32 $Y=0 $X2=5.52
+ $Y2=0
r142 46 60 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=2.64 $Y2=0
r143 44 55 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.24 $Y=0 $X2=2.16
+ $Y2=0
r144 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=0 $X2=2.405
+ $Y2=0
r145 43 59 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.57 $Y=0 $X2=2.64
+ $Y2=0
r146 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.57 $Y=0 $X2=2.405
+ $Y2=0
r147 39 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.93 $Y=0.085
+ $X2=7.93 $Y2=0
r148 39 41 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=7.93 $Y=0.085
+ $X2=7.93 $Y2=0.535
r149 35 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.93 $Y=0.085
+ $X2=6.93 $Y2=0
r150 35 37 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=6.93 $Y=0.085
+ $X2=6.93 $Y2=0.535
r151 31 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.93 $Y=0.085
+ $X2=5.93 $Y2=0
r152 31 33 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=5.93 $Y=0.085
+ $X2=5.93 $Y2=0.535
r153 27 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.405 $Y=0.085
+ $X2=2.405 $Y2=0
r154 27 29 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.405 $Y=0.085
+ $X2=2.405 $Y2=0.515
r155 23 83 1.82608 $w=4.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.342 $Y=0.085
+ $X2=1.342 $Y2=0
r156 23 25 11.3036 $w=4.53e-07 $l=4.3e-07 $layer=LI1_cond $X=1.342 $Y=0.085
+ $X2=1.342 $Y2=0.515
r157 19 80 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r158 19 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.515
r159 6 41 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=7.775
+ $Y=0.39 $X2=7.93 $Y2=0.535
r160 5 37 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=6.72
+ $Y=0.39 $X2=6.93 $Y2=0.535
r161 4 33 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=5.75
+ $Y=0.39 $X2=5.93 $Y2=0.535
r162 3 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.265
+ $Y=0.37 $X2=2.405 $Y2=0.515
r163 2 25 182 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.34 $Y2=0.515
r164 1 21 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.35 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_4%A_564_78# 1 2 3 4 5 18 20 21 23 26 30 32 36
+ 38 40 42 46 48
r83 40 50 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.4 $Y=0.79 $X2=8.4
+ $Y2=0.875
r84 40 42 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=8.4 $Y=0.79 $X2=8.4
+ $Y2=0.515
r85 39 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.595 $Y=0.875
+ $X2=7.43 $Y2=0.875
r86 38 50 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.275 $Y=0.875
+ $X2=8.4 $Y2=0.875
r87 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.275 $Y=0.875
+ $X2=7.595 $Y2=0.875
r88 34 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.43 $Y=0.79 $X2=7.43
+ $Y2=0.875
r89 34 36 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=7.43 $Y=0.79
+ $X2=7.43 $Y2=0.515
r90 33 46 8.61065 $w=1.7e-07 $l=1.86145e-07 $layer=LI1_cond $X=6.595 $Y=0.875
+ $X2=6.43 $Y2=0.92
r91 32 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.265 $Y=0.875
+ $X2=7.43 $Y2=0.875
r92 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.265 $Y=0.875
+ $X2=6.595 $Y2=0.875
r93 28 46 0.89609 $w=3.3e-07 $l=1.3e-07 $layer=LI1_cond $X=6.43 $Y=0.79 $X2=6.43
+ $Y2=0.92
r94 28 30 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=6.43 $Y=0.79
+ $X2=6.43 $Y2=0.535
r95 27 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.595 $Y=0.875
+ $X2=5.43 $Y2=0.875
r96 26 46 8.61065 $w=1.7e-07 $l=1.86145e-07 $layer=LI1_cond $X=6.265 $Y=0.875
+ $X2=6.43 $Y2=0.92
r97 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.265 $Y=0.875
+ $X2=5.595 $Y2=0.875
r98 23 45 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.43 $Y=0.79 $X2=5.43
+ $Y2=0.875
r99 23 25 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.43 $Y=0.79
+ $X2=5.43 $Y2=0.535
r100 22 25 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=5.43 $Y=0.425
+ $X2=5.43 $Y2=0.535
r101 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.265 $Y=0.34
+ $X2=5.43 $Y2=0.425
r102 20 21 139.289 $w=1.68e-07 $l=2.135e-06 $layer=LI1_cond $X=5.265 $Y=0.34
+ $X2=3.13 $Y2=0.34
r103 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.965 $Y=0.425
+ $X2=3.13 $Y2=0.34
r104 16 18 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.965 $Y=0.425
+ $X2=2.965 $Y2=0.67
r105 5 50 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=8.22
+ $Y=0.39 $X2=8.36 $Y2=0.875
r106 5 42 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=8.22
+ $Y=0.39 $X2=8.36 $Y2=0.515
r107 4 48 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=7.245
+ $Y=0.39 $X2=7.43 $Y2=0.875
r108 4 36 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=7.245
+ $Y=0.39 $X2=7.43 $Y2=0.515
r109 3 30 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=6.285
+ $Y=0.39 $X2=6.43 $Y2=0.535
r110 2 45 182 $w=1.7e-07 $l=5.80582e-07 $layer=licon1_NDIFF $count=1 $X=5.22
+ $Y=0.39 $X2=5.43 $Y2=0.875
r111 2 25 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.22
+ $Y=0.39 $X2=5.43 $Y2=0.535
r112 1 18 182 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_NDIFF $count=1 $X=2.82
+ $Y=0.39 $X2=2.965 $Y2=0.67
.ends

.subckt PM_SKY130_FD_SC_MS__O311A_4%A_651_78# 1 2 9 12 13 14
r20 14 17 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=4.93 $Y=0.68
+ $X2=4.93 $Y2=0.775
r21 12 13 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.91 $Y=0.76
+ $X2=4.075 $Y2=0.76
r22 9 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.765 $Y=0.68
+ $X2=4.93 $Y2=0.68
r23 9 13 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.765 $Y=0.68
+ $X2=4.075 $Y2=0.68
r24 2 17 182 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_NDIFF $count=1 $X=4.79
+ $Y=0.39 $X2=4.93 $Y2=0.775
r25 1 12 91 $w=1.7e-07 $l=8.19375e-07 $layer=licon1_NDIFF $count=2 $X=3.255
+ $Y=0.39 $X2=3.91 $Y2=0.76
.ends


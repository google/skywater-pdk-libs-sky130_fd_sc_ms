* File: sky130_fd_sc_ms__a2111oi_2.pxi.spice
* Created: Fri Aug 28 16:55:58 2020
* 
x_PM_SKY130_FD_SC_MS__A2111OI_2%D1 N_D1_M1003_g N_D1_M1007_g N_D1_M1004_g D1 D1
+ N_D1_c_92_n PM_SKY130_FD_SC_MS__A2111OI_2%D1
x_PM_SKY130_FD_SC_MS__A2111OI_2%C1 N_C1_M1000_g N_C1_c_132_n N_C1_M1006_g
+ N_C1_c_133_n N_C1_M1008_g C1 C1 C1 N_C1_c_131_n
+ PM_SKY130_FD_SC_MS__A2111OI_2%C1
x_PM_SKY130_FD_SC_MS__A2111OI_2%B1 N_B1_c_171_n N_B1_M1009_g N_B1_c_172_n
+ N_B1_M1010_g N_B1_M1011_g B1 B1 N_B1_c_176_n N_B1_c_177_n
+ PM_SKY130_FD_SC_MS__A2111OI_2%B1
x_PM_SKY130_FD_SC_MS__A2111OI_2%A1 N_A1_M1012_g N_A1_M1001_g N_A1_M1015_g
+ N_A1_M1014_g A1 A1 N_A1_c_223_n PM_SKY130_FD_SC_MS__A2111OI_2%A1
x_PM_SKY130_FD_SC_MS__A2111OI_2%A2 N_A2_M1002_g N_A2_M1005_g N_A2_M1013_g
+ N_A2_M1016_g A2 N_A2_c_277_n N_A2_c_278_n PM_SKY130_FD_SC_MS__A2111OI_2%A2
x_PM_SKY130_FD_SC_MS__A2111OI_2%A_69_368# N_A_69_368#_M1003_s
+ N_A_69_368#_M1004_s N_A_69_368#_M1008_s N_A_69_368#_c_313_n
+ N_A_69_368#_c_314_n N_A_69_368#_c_315_n N_A_69_368#_c_321_n
+ N_A_69_368#_c_316_n N_A_69_368#_c_317_n N_A_69_368#_c_318_n
+ PM_SKY130_FD_SC_MS__A2111OI_2%A_69_368#
x_PM_SKY130_FD_SC_MS__A2111OI_2%Y N_Y_M1007_d N_Y_M1009_d N_Y_M1001_s
+ N_Y_M1003_d N_Y_c_345_n N_Y_c_346_n N_Y_c_360_n N_Y_c_355_n N_Y_c_347_n
+ N_Y_c_348_n N_Y_c_349_n N_Y_c_350_n N_Y_c_363_n N_Y_c_351_n N_Y_c_352_n
+ N_Y_c_353_n Y Y PM_SKY130_FD_SC_MS__A2111OI_2%Y
x_PM_SKY130_FD_SC_MS__A2111OI_2%A_337_368# N_A_337_368#_M1006_d
+ N_A_337_368#_M1010_d N_A_337_368#_c_416_n N_A_337_368#_c_420_n
+ N_A_337_368#_c_417_n PM_SKY130_FD_SC_MS__A2111OI_2%A_337_368#
x_PM_SKY130_FD_SC_MS__A2111OI_2%A_533_368# N_A_533_368#_M1010_s
+ N_A_533_368#_M1011_s N_A_533_368#_M1015_s N_A_533_368#_M1016_d
+ N_A_533_368#_c_439_n N_A_533_368#_c_440_n N_A_533_368#_c_441_n
+ N_A_533_368#_c_448_n N_A_533_368#_c_450_n N_A_533_368#_c_456_n
+ N_A_533_368#_c_442_n N_A_533_368#_c_465_n N_A_533_368#_c_443_n
+ N_A_533_368#_c_444_n N_A_533_368#_c_462_n
+ PM_SKY130_FD_SC_MS__A2111OI_2%A_533_368#
x_PM_SKY130_FD_SC_MS__A2111OI_2%VPWR N_VPWR_M1012_d N_VPWR_M1002_s
+ N_VPWR_c_495_n N_VPWR_c_496_n VPWR N_VPWR_c_497_n N_VPWR_c_498_n
+ N_VPWR_c_499_n N_VPWR_c_494_n N_VPWR_c_501_n N_VPWR_c_502_n
+ PM_SKY130_FD_SC_MS__A2111OI_2%VPWR
x_PM_SKY130_FD_SC_MS__A2111OI_2%VGND N_VGND_M1007_s N_VGND_M1000_d
+ N_VGND_M1005_s N_VGND_c_552_n N_VGND_c_553_n N_VGND_c_554_n N_VGND_c_555_n
+ VGND N_VGND_c_556_n N_VGND_c_557_n N_VGND_c_558_n N_VGND_c_559_n
+ N_VGND_c_560_n N_VGND_c_561_n PM_SKY130_FD_SC_MS__A2111OI_2%VGND
x_PM_SKY130_FD_SC_MS__A2111OI_2%A_722_74# N_A_722_74#_M1001_d
+ N_A_722_74#_M1014_d N_A_722_74#_M1013_d N_A_722_74#_c_605_n
+ N_A_722_74#_c_606_n N_A_722_74#_c_607_n N_A_722_74#_c_608_n
+ N_A_722_74#_c_609_n PM_SKY130_FD_SC_MS__A2111OI_2%A_722_74#
cc_1 VNB N_D1_M1007_g 0.0296222f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.74
cc_2 VNB D1 0.00551793f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_3 VNB N_D1_c_92_n 0.0484877f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.515
cc_4 VNB N_C1_M1000_g 0.0273389f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.4
cc_5 VNB C1 0.0165977f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_6 VNB N_C1_c_131_n 0.0371835f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.515
cc_7 VNB N_B1_c_171_n 0.0201467f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.68
cc_8 VNB N_B1_c_172_n 0.00913645f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.35
cc_9 VNB N_B1_M1010_g 0.0064155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B1_M1011_g 0.00598961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB B1 0.0124371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B1_c_176_n 0.0446588f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.515
cc_13 VNB N_B1_c_177_n 0.0556069f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.515
cc_14 VNB N_A1_M1001_g 0.0295402f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.74
cc_15 VNB N_A1_M1014_g 0.024081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB A1 0.00589944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_c_223_n 0.0347619f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.565
cc_18 VNB N_A2_M1005_g 0.023157f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.74
cc_19 VNB N_A2_M1013_g 0.0320221f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=2.4
cc_20 VNB N_A2_c_277_n 0.00102489f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.515
cc_21 VNB N_A2_c_278_n 0.0473252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_345_n 0.0238079f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_23 VNB N_Y_c_346_n 0.0177372f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_24 VNB N_Y_c_347_n 0.00327056f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.515
cc_25 VNB N_Y_c_348_n 0.00305444f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.515
cc_26 VNB N_Y_c_349_n 0.0188906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_350_n 0.0355113f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_28 VNB N_Y_c_351_n 0.00821167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_352_n 0.0108587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_353_n 0.00250929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB Y 0.025793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_494_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_552_n 0.0274256f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_34 VNB N_VGND_c_553_n 0.0184856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_554_n 0.00917051f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.515
cc_36 VNB N_VGND_c_555_n 0.00396562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_556_n 0.0795701f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.565
cc_38 VNB N_VGND_c_557_n 0.0178682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_558_n 0.348653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_559_n 0.0293037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_560_n 0.00653982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_561_n 0.00622543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_722_74#_c_605_n 0.016287f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=2.4
cc_44 VNB N_A_722_74#_c_606_n 0.0016059f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_45 VNB N_A_722_74#_c_607_n 0.0172894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_722_74#_c_608_n 0.00250711f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.515
cc_47 VNB N_A_722_74#_c_609_n 0.0270834f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.515
cc_48 VPB N_D1_M1003_g 0.0238279f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=2.4
cc_49 VPB N_D1_M1004_g 0.0197881f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=2.4
cc_50 VPB D1 0.00679131f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_51 VPB N_D1_c_92_n 0.00652678f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=1.515
cc_52 VPB N_C1_c_132_n 0.0177675f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.35
cc_53 VPB N_C1_c_133_n 0.0225686f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB C1 0.0123734f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_55 VPB N_C1_c_131_n 0.00955879f $X=-0.19 $Y=1.66 $X2=1.13 $Y2=1.515
cc_56 VPB N_B1_M1010_g 0.0262613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_B1_M1011_g 0.0219145f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A1_M1012_g 0.0208333f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=2.4
cc_59 VPB N_A1_M1015_g 0.0208092f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=2.4
cc_60 VPB A1 0.00542803f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A1_c_223_n 0.00455847f $X=-0.19 $Y=1.66 $X2=1.13 $Y2=1.565
cc_62 VPB N_A2_M1002_g 0.0207899f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=2.4
cc_63 VPB N_A2_M1016_g 0.028131f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A2_c_277_n 0.00251564f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=1.515
cc_65 VPB N_A2_c_278_n 0.00538531f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_69_368#_c_313_n 0.0233684f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_69_368#_c_314_n 0.0026202f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_68 VPB N_A_69_368#_c_315_n 0.00933537f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_69_368#_c_316_n 0.00629773f $X=-0.19 $Y=1.66 $X2=1.13 $Y2=1.515
cc_70 VPB N_A_69_368#_c_317_n 0.0058157f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_69_368#_c_318_n 0.00123754f $X=-0.19 $Y=1.66 $X2=1.13 $Y2=1.565
cc_72 VPB N_Y_c_355_n 0.0160034f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB Y 0.0141982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_337_368#_c_416_n 0.0110263f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=1.68
cc_75 VPB N_A_337_368#_c_417_n 0.0023439f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_533_368#_c_439_n 0.00582476f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_533_368#_c_440_n 0.00402322f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.515
cc_78 VPB N_A_533_368#_c_441_n 0.00389592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_533_368#_c_442_n 0.00202354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_533_368#_c_443_n 0.0171219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_533_368#_c_444_n 0.0345796f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_495_n 0.0070415f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=1.68
cc_83 VPB N_VPWR_c_496_n 0.00339119f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_84 VPB N_VPWR_c_497_n 0.0986435f $X=-0.19 $Y=1.66 $X2=0.695 $Y2=1.515
cc_85 VPB N_VPWR_c_498_n 0.0185125f $X=-0.19 $Y=1.66 $X2=1.13 $Y2=1.515
cc_86 VPB N_VPWR_c_499_n 0.0177091f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_87 VPB N_VPWR_c_494_n 0.0892464f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_501_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_502_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 N_D1_M1007_g N_C1_M1000_g 0.0207626f $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_91 D1 C1 0.0351515f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_92 N_D1_c_92_n C1 3.90301e-19 $X=1.145 $Y=1.515 $X2=0 $Y2=0
cc_93 N_D1_M1004_g N_C1_c_131_n 0.0184903f $X=1.145 $Y=2.4 $X2=0 $Y2=0
cc_94 D1 N_C1_c_131_n 0.00168672f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_95 N_D1_c_92_n N_C1_c_131_n 0.0215303f $X=1.145 $Y=1.515 $X2=0 $Y2=0
cc_96 N_D1_M1003_g N_A_69_368#_c_314_n 0.0149887f $X=0.695 $Y=2.4 $X2=0 $Y2=0
cc_97 N_D1_M1004_g N_A_69_368#_c_314_n 0.0139961f $X=1.145 $Y=2.4 $X2=0 $Y2=0
cc_98 D1 N_A_69_368#_c_321_n 0.00229424f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_99 N_D1_M1007_g N_Y_c_345_n 0.0169004f $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_100 D1 N_Y_c_345_n 0.0419733f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_101 N_D1_c_92_n N_Y_c_345_n 0.0103192f $X=1.145 $Y=1.515 $X2=0 $Y2=0
cc_102 N_D1_M1003_g N_Y_c_360_n 0.0147399f $X=0.695 $Y=2.4 $X2=0 $Y2=0
cc_103 D1 N_Y_c_360_n 0.0109106f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_104 N_D1_M1007_g N_Y_c_347_n 0.00383226f $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_105 N_D1_M1003_g N_Y_c_363_n 0.0150733f $X=0.695 $Y=2.4 $X2=0 $Y2=0
cc_106 N_D1_M1004_g N_Y_c_363_n 0.010896f $X=1.145 $Y=2.4 $X2=0 $Y2=0
cc_107 D1 N_Y_c_363_n 0.0235495f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_108 N_D1_c_92_n N_Y_c_363_n 5.54777e-19 $X=1.145 $Y=1.515 $X2=0 $Y2=0
cc_109 D1 N_Y_c_351_n 0.0133987f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_110 N_D1_c_92_n N_Y_c_351_n 0.00344073f $X=1.145 $Y=1.515 $X2=0 $Y2=0
cc_111 N_D1_M1003_g Y 0.0056647f $X=0.695 $Y=2.4 $X2=0 $Y2=0
cc_112 N_D1_M1007_g Y 0.00380025f $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_113 D1 Y 0.0262077f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_114 N_D1_c_92_n Y 0.00284307f $X=1.145 $Y=1.515 $X2=0 $Y2=0
cc_115 N_D1_M1003_g N_VPWR_c_497_n 0.00333926f $X=0.695 $Y=2.4 $X2=0 $Y2=0
cc_116 N_D1_M1004_g N_VPWR_c_497_n 0.00333926f $X=1.145 $Y=2.4 $X2=0 $Y2=0
cc_117 N_D1_M1003_g N_VPWR_c_494_n 0.00426932f $X=0.695 $Y=2.4 $X2=0 $Y2=0
cc_118 N_D1_M1004_g N_VPWR_c_494_n 0.00422798f $X=1.145 $Y=2.4 $X2=0 $Y2=0
cc_119 N_D1_M1007_g N_VGND_c_552_n 0.0129243f $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_120 N_D1_M1007_g N_VGND_c_553_n 0.00383152f $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_121 N_D1_M1007_g N_VGND_c_558_n 0.00758569f $X=1.04 $Y=0.74 $X2=0 $Y2=0
cc_122 N_C1_M1000_g N_B1_c_171_n 0.0247539f $X=1.58 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_123 C1 N_B1_c_172_n 0.0170771f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_124 N_C1_c_131_n N_B1_c_172_n 0.00496204f $X=1.67 $Y=1.515 $X2=0 $Y2=0
cc_125 C1 B1 0.0132423f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_126 C1 N_B1_c_177_n 0.0151105f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_127 N_C1_c_132_n N_A_69_368#_c_316_n 0.0139518f $X=1.595 $Y=1.725 $X2=0 $Y2=0
cc_128 N_C1_c_133_n N_A_69_368#_c_316_n 0.0149887f $X=2.045 $Y=1.725 $X2=0 $Y2=0
cc_129 N_C1_M1000_g N_Y_c_347_n 5.52855e-19 $X=1.58 $Y=0.74 $X2=0 $Y2=0
cc_130 N_C1_M1000_g N_Y_c_348_n 0.0145564f $X=1.58 $Y=0.74 $X2=0 $Y2=0
cc_131 C1 N_Y_c_348_n 0.0514073f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_132 N_C1_c_131_n N_Y_c_348_n 0.00548075f $X=1.67 $Y=1.515 $X2=0 $Y2=0
cc_133 N_C1_M1000_g N_Y_c_349_n 8.24518e-19 $X=1.58 $Y=0.74 $X2=0 $Y2=0
cc_134 C1 N_Y_c_350_n 0.0120661f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_135 C1 N_Y_c_352_n 0.0294457f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_136 N_C1_c_133_n N_A_337_368#_c_416_n 0.0150161f $X=2.045 $Y=1.725 $X2=0
+ $Y2=0
cc_137 C1 N_A_337_368#_c_416_n 0.0585844f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_138 N_C1_c_132_n N_A_337_368#_c_420_n 0.010896f $X=1.595 $Y=1.725 $X2=0 $Y2=0
cc_139 N_C1_c_133_n N_A_337_368#_c_420_n 0.0150733f $X=2.045 $Y=1.725 $X2=0
+ $Y2=0
cc_140 C1 N_A_337_368#_c_420_n 0.0235494f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_141 N_C1_c_131_n N_A_337_368#_c_420_n 6.18429e-19 $X=1.67 $Y=1.515 $X2=0
+ $Y2=0
cc_142 N_C1_c_133_n N_A_533_368#_c_441_n 5.81668e-19 $X=2.045 $Y=1.725 $X2=0
+ $Y2=0
cc_143 N_C1_c_132_n N_VPWR_c_497_n 0.00333926f $X=1.595 $Y=1.725 $X2=0 $Y2=0
cc_144 N_C1_c_133_n N_VPWR_c_497_n 0.00333926f $X=2.045 $Y=1.725 $X2=0 $Y2=0
cc_145 N_C1_c_132_n N_VPWR_c_494_n 0.00422798f $X=1.595 $Y=1.725 $X2=0 $Y2=0
cc_146 N_C1_c_133_n N_VPWR_c_494_n 0.0042782f $X=2.045 $Y=1.725 $X2=0 $Y2=0
cc_147 N_C1_M1000_g N_VGND_c_552_n 4.50149e-19 $X=1.58 $Y=0.74 $X2=0 $Y2=0
cc_148 N_C1_M1000_g N_VGND_c_553_n 0.00461464f $X=1.58 $Y=0.74 $X2=0 $Y2=0
cc_149 N_C1_M1000_g N_VGND_c_554_n 0.00279591f $X=1.58 $Y=0.74 $X2=0 $Y2=0
cc_150 N_C1_M1000_g N_VGND_c_558_n 0.0090927f $X=1.58 $Y=0.74 $X2=0 $Y2=0
cc_151 N_B1_M1011_g N_A1_M1012_g 0.0158122f $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_152 B1 N_A1_M1001_g 0.00481817f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_153 N_B1_c_177_n N_A1_M1001_g 0.00561135f $X=3.465 $Y=1.367 $X2=0 $Y2=0
cc_154 B1 A1 0.0132858f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_155 N_B1_c_177_n A1 0.00126148f $X=3.465 $Y=1.367 $X2=0 $Y2=0
cc_156 B1 N_A1_c_223_n 0.00199478f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_157 N_B1_c_177_n N_A1_c_223_n 0.0158122f $X=3.465 $Y=1.367 $X2=0 $Y2=0
cc_158 N_B1_M1010_g N_A_69_368#_c_316_n 5.81668e-19 $X=3.015 $Y=2.4 $X2=0 $Y2=0
cc_159 N_B1_c_171_n N_Y_c_348_n 0.0116603f $X=2.12 $Y=1.185 $X2=0 $Y2=0
cc_160 N_B1_c_171_n N_Y_c_349_n 0.00612384f $X=2.12 $Y=1.185 $X2=0 $Y2=0
cc_161 B1 N_Y_c_350_n 0.0503328f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_162 N_B1_c_176_n N_Y_c_350_n 0.0141472f $X=2.925 $Y=1.367 $X2=0 $Y2=0
cc_163 N_B1_c_177_n N_Y_c_350_n 0.00370226f $X=3.465 $Y=1.367 $X2=0 $Y2=0
cc_164 N_B1_c_171_n N_Y_c_352_n 0.00662344f $X=2.12 $Y=1.185 $X2=0 $Y2=0
cc_165 N_B1_c_176_n N_Y_c_352_n 0.00744713f $X=2.925 $Y=1.367 $X2=0 $Y2=0
cc_166 N_B1_M1010_g N_A_337_368#_c_416_n 0.0180631f $X=3.015 $Y=2.4 $X2=0 $Y2=0
cc_167 B1 N_A_337_368#_c_416_n 0.00251507f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_168 N_B1_c_176_n N_A_337_368#_c_416_n 0.00358973f $X=2.925 $Y=1.367 $X2=0
+ $Y2=0
cc_169 N_B1_M1010_g N_A_337_368#_c_417_n 0.0213497f $X=3.015 $Y=2.4 $X2=0 $Y2=0
cc_170 N_B1_M1011_g N_A_337_368#_c_417_n 4.97677e-19 $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_171 B1 N_A_337_368#_c_417_n 0.0149146f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_172 N_B1_c_177_n N_A_337_368#_c_417_n 0.00202078f $X=3.465 $Y=1.367 $X2=0
+ $Y2=0
cc_173 N_B1_M1010_g N_A_533_368#_c_440_n 0.0149887f $X=3.015 $Y=2.4 $X2=0 $Y2=0
cc_174 N_B1_M1011_g N_A_533_368#_c_440_n 0.0135505f $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_175 N_B1_M1011_g N_A_533_368#_c_448_n 0.00269738f $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_176 B1 N_A_533_368#_c_448_n 0.00740358f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_177 N_B1_M1010_g N_A_533_368#_c_450_n 7.18074e-19 $X=3.015 $Y=2.4 $X2=0 $Y2=0
cc_178 N_B1_M1011_g N_A_533_368#_c_450_n 0.0108836f $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_179 N_B1_M1010_g N_VPWR_c_497_n 0.00333926f $X=3.015 $Y=2.4 $X2=0 $Y2=0
cc_180 N_B1_M1011_g N_VPWR_c_497_n 0.00333896f $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_181 N_B1_M1010_g N_VPWR_c_494_n 0.0042782f $X=3.015 $Y=2.4 $X2=0 $Y2=0
cc_182 N_B1_M1011_g N_VPWR_c_494_n 0.00422796f $X=3.465 $Y=2.4 $X2=0 $Y2=0
cc_183 N_B1_c_171_n N_VGND_c_554_n 0.00602646f $X=2.12 $Y=1.185 $X2=0 $Y2=0
cc_184 N_B1_c_171_n N_VGND_c_556_n 0.00434272f $X=2.12 $Y=1.185 $X2=0 $Y2=0
cc_185 N_B1_c_171_n N_VGND_c_558_n 0.00826088f $X=2.12 $Y=1.185 $X2=0 $Y2=0
cc_186 N_A1_M1015_g N_A2_M1002_g 0.0147666f $X=4.365 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A1_M1014_g N_A2_M1005_g 0.019323f $X=4.38 $Y=0.74 $X2=0 $Y2=0
cc_188 A1 N_A2_c_277_n 0.0353991f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_189 N_A1_c_223_n N_A2_c_277_n 3.141e-19 $X=4.38 $Y=1.515 $X2=0 $Y2=0
cc_190 A1 N_A2_c_278_n 0.00400504f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_191 N_A1_c_223_n N_A2_c_278_n 0.0147666f $X=4.38 $Y=1.515 $X2=0 $Y2=0
cc_192 N_A1_M1001_g N_Y_c_350_n 0.0149884f $X=3.95 $Y=0.74 $X2=0 $Y2=0
cc_193 A1 N_Y_c_350_n 0.00137046f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_194 N_A1_M1001_g N_Y_c_353_n 0.00878264f $X=3.95 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A1_M1014_g N_Y_c_353_n 0.00464929f $X=4.38 $Y=0.74 $X2=0 $Y2=0
cc_196 A1 N_Y_c_353_n 0.0218587f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_197 N_A1_c_223_n N_Y_c_353_n 0.00233006f $X=4.38 $Y=1.515 $X2=0 $Y2=0
cc_198 N_A1_M1012_g N_A_533_368#_c_440_n 0.00347836f $X=3.915 $Y=2.4 $X2=0 $Y2=0
cc_199 N_A1_M1012_g N_A_533_368#_c_448_n 0.00190089f $X=3.915 $Y=2.4 $X2=0 $Y2=0
cc_200 N_A1_M1012_g N_A_533_368#_c_450_n 0.0107569f $X=3.915 $Y=2.4 $X2=0 $Y2=0
cc_201 N_A1_M1015_g N_A_533_368#_c_450_n 6.26485e-19 $X=4.365 $Y=2.4 $X2=0 $Y2=0
cc_202 N_A1_M1012_g N_A_533_368#_c_456_n 0.0162265f $X=3.915 $Y=2.4 $X2=0 $Y2=0
cc_203 N_A1_M1015_g N_A_533_368#_c_456_n 0.012931f $X=4.365 $Y=2.4 $X2=0 $Y2=0
cc_204 A1 N_A_533_368#_c_456_n 0.0311948f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_205 N_A1_c_223_n N_A_533_368#_c_456_n 4.89356e-19 $X=4.38 $Y=1.515 $X2=0
+ $Y2=0
cc_206 N_A1_M1012_g N_A_533_368#_c_442_n 6.52999e-19 $X=3.915 $Y=2.4 $X2=0 $Y2=0
cc_207 N_A1_M1015_g N_A_533_368#_c_442_n 0.0120602f $X=4.365 $Y=2.4 $X2=0 $Y2=0
cc_208 N_A1_M1015_g N_A_533_368#_c_462_n 8.84614e-19 $X=4.365 $Y=2.4 $X2=0 $Y2=0
cc_209 A1 N_A_533_368#_c_462_n 0.0189744f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_210 N_A1_M1012_g N_VPWR_c_495_n 0.00120619f $X=3.915 $Y=2.4 $X2=0 $Y2=0
cc_211 N_A1_M1015_g N_VPWR_c_495_n 0.00156821f $X=4.365 $Y=2.4 $X2=0 $Y2=0
cc_212 N_A1_M1015_g N_VPWR_c_496_n 5.60169e-19 $X=4.365 $Y=2.4 $X2=0 $Y2=0
cc_213 N_A1_M1012_g N_VPWR_c_497_n 0.00517089f $X=3.915 $Y=2.4 $X2=0 $Y2=0
cc_214 N_A1_M1015_g N_VPWR_c_498_n 0.005209f $X=4.365 $Y=2.4 $X2=0 $Y2=0
cc_215 N_A1_M1012_g N_VPWR_c_494_n 0.00977588f $X=3.915 $Y=2.4 $X2=0 $Y2=0
cc_216 N_A1_M1015_g N_VPWR_c_494_n 0.00982376f $X=4.365 $Y=2.4 $X2=0 $Y2=0
cc_217 N_A1_M1014_g N_VGND_c_555_n 6.35092e-19 $X=4.38 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A1_M1001_g N_VGND_c_556_n 0.00291649f $X=3.95 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A1_M1014_g N_VGND_c_556_n 0.00291649f $X=4.38 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A1_M1001_g N_VGND_c_558_n 0.00363173f $X=3.95 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A1_M1014_g N_VGND_c_558_n 0.00359219f $X=4.38 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A1_M1001_g N_A_722_74#_c_605_n 0.010283f $X=3.95 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A1_M1014_g N_A_722_74#_c_605_n 0.0142063f $X=4.38 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A1_M1014_g N_A_722_74#_c_608_n 0.00174382f $X=4.38 $Y=0.74 $X2=0 $Y2=0
cc_225 A1 N_A_722_74#_c_608_n 0.0148778f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_226 N_A2_M1002_g N_A_533_368#_c_442_n 2.39324e-19 $X=4.815 $Y=2.4 $X2=0 $Y2=0
cc_227 N_A2_M1002_g N_A_533_368#_c_465_n 0.0180558f $X=4.815 $Y=2.4 $X2=0 $Y2=0
cc_228 N_A2_M1016_g N_A_533_368#_c_465_n 0.0194091f $X=5.265 $Y=2.4 $X2=0 $Y2=0
cc_229 N_A2_c_277_n N_A_533_368#_c_465_n 0.0217013f $X=5.015 $Y=1.515 $X2=0
+ $Y2=0
cc_230 N_A2_c_278_n N_A_533_368#_c_465_n 4.89879e-19 $X=5.25 $Y=1.515 $X2=0
+ $Y2=0
cc_231 N_A2_M1016_g N_A_533_368#_c_443_n 8.13654e-19 $X=5.265 $Y=2.4 $X2=0 $Y2=0
cc_232 N_A2_M1016_g N_A_533_368#_c_444_n 0.00147311f $X=5.265 $Y=2.4 $X2=0 $Y2=0
cc_233 N_A2_M1002_g N_VPWR_c_496_n 0.0131455f $X=4.815 $Y=2.4 $X2=0 $Y2=0
cc_234 N_A2_M1016_g N_VPWR_c_496_n 0.0160814f $X=5.265 $Y=2.4 $X2=0 $Y2=0
cc_235 N_A2_M1002_g N_VPWR_c_498_n 0.00460063f $X=4.815 $Y=2.4 $X2=0 $Y2=0
cc_236 N_A2_M1016_g N_VPWR_c_499_n 0.00460063f $X=5.265 $Y=2.4 $X2=0 $Y2=0
cc_237 N_A2_M1002_g N_VPWR_c_494_n 0.00908665f $X=4.815 $Y=2.4 $X2=0 $Y2=0
cc_238 N_A2_M1016_g N_VPWR_c_494_n 0.00912261f $X=5.265 $Y=2.4 $X2=0 $Y2=0
cc_239 N_A2_M1005_g N_VGND_c_555_n 0.0108748f $X=4.81 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A2_M1013_g N_VGND_c_555_n 0.0137776f $X=5.25 $Y=0.74 $X2=0 $Y2=0
cc_241 N_A2_M1005_g N_VGND_c_556_n 0.00383152f $X=4.81 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A2_M1013_g N_VGND_c_557_n 0.00383152f $X=5.25 $Y=0.74 $X2=0 $Y2=0
cc_243 N_A2_M1005_g N_VGND_c_558_n 0.00757637f $X=4.81 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A2_M1013_g N_VGND_c_558_n 0.00761248f $X=5.25 $Y=0.74 $X2=0 $Y2=0
cc_245 N_A2_M1005_g N_A_722_74#_c_607_n 0.0164989f $X=4.81 $Y=0.74 $X2=0 $Y2=0
cc_246 N_A2_M1013_g N_A_722_74#_c_607_n 0.0180697f $X=5.25 $Y=0.74 $X2=0 $Y2=0
cc_247 N_A2_c_277_n N_A_722_74#_c_607_n 0.0251424f $X=5.015 $Y=1.515 $X2=0 $Y2=0
cc_248 N_A2_c_278_n N_A_722_74#_c_607_n 0.00224972f $X=5.25 $Y=1.515 $X2=0 $Y2=0
cc_249 N_A2_M1013_g N_A_722_74#_c_609_n 0.00159319f $X=5.25 $Y=0.74 $X2=0 $Y2=0
cc_250 N_A_69_368#_c_314_n N_Y_M1003_d 0.00165831f $X=1.285 $Y=2.99 $X2=0 $Y2=0
cc_251 N_A_69_368#_M1003_s N_Y_c_360_n 0.0100085f $X=0.345 $Y=1.84 $X2=0 $Y2=0
cc_252 N_A_69_368#_c_313_n N_Y_c_360_n 0.0156657f $X=0.47 $Y=2.455 $X2=0 $Y2=0
cc_253 N_A_69_368#_c_313_n N_Y_c_355_n 0.00451074f $X=0.47 $Y=2.455 $X2=0 $Y2=0
cc_254 N_A_69_368#_c_314_n N_Y_c_363_n 0.0159318f $X=1.285 $Y=2.99 $X2=0 $Y2=0
cc_255 N_A_69_368#_M1003_s Y 0.00144714f $X=0.345 $Y=1.84 $X2=0 $Y2=0
cc_256 N_A_69_368#_c_316_n N_A_337_368#_M1006_d 0.00165831f $X=2.185 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_257 N_A_69_368#_M1008_s N_A_337_368#_c_416_n 0.00488721f $X=2.135 $Y=1.84
+ $X2=0 $Y2=0
cc_258 N_A_69_368#_c_317_n N_A_337_368#_c_416_n 0.0198097f $X=2.27 $Y=2.455
+ $X2=0 $Y2=0
cc_259 N_A_69_368#_c_316_n N_A_337_368#_c_420_n 0.0159318f $X=2.185 $Y=2.99
+ $X2=0 $Y2=0
cc_260 N_A_69_368#_c_317_n N_A_533_368#_c_439_n 0.0457256f $X=2.27 $Y=2.455
+ $X2=0 $Y2=0
cc_261 N_A_69_368#_c_316_n N_A_533_368#_c_441_n 0.0147157f $X=2.185 $Y=2.99
+ $X2=0 $Y2=0
cc_262 N_A_69_368#_c_314_n N_VPWR_c_497_n 0.0459191f $X=1.285 $Y=2.99 $X2=0
+ $Y2=0
cc_263 N_A_69_368#_c_315_n N_VPWR_c_497_n 0.0179217f $X=0.555 $Y=2.99 $X2=0
+ $Y2=0
cc_264 N_A_69_368#_c_316_n N_VPWR_c_497_n 0.0638408f $X=2.185 $Y=2.99 $X2=0
+ $Y2=0
cc_265 N_A_69_368#_c_318_n N_VPWR_c_497_n 0.0121867f $X=1.37 $Y=2.99 $X2=0 $Y2=0
cc_266 N_A_69_368#_c_314_n N_VPWR_c_494_n 0.0258001f $X=1.285 $Y=2.99 $X2=0
+ $Y2=0
cc_267 N_A_69_368#_c_315_n N_VPWR_c_494_n 0.00971942f $X=0.555 $Y=2.99 $X2=0
+ $Y2=0
cc_268 N_A_69_368#_c_316_n N_VPWR_c_494_n 0.0355196f $X=2.185 $Y=2.99 $X2=0
+ $Y2=0
cc_269 N_A_69_368#_c_318_n N_VPWR_c_494_n 0.00660921f $X=1.37 $Y=2.99 $X2=0
+ $Y2=0
cc_270 N_Y_c_345_n N_VGND_M1007_s 0.00299905f $X=1.16 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_271 N_Y_c_348_n N_VGND_M1000_d 0.00309832f $X=2.17 $Y=1.095 $X2=0 $Y2=0
cc_272 N_Y_c_345_n N_VGND_c_552_n 0.0219406f $X=1.16 $Y=1.095 $X2=0 $Y2=0
cc_273 N_Y_c_347_n N_VGND_c_552_n 0.0191765f $X=1.325 $Y=0.515 $X2=0 $Y2=0
cc_274 N_Y_c_347_n N_VGND_c_553_n 0.0146357f $X=1.325 $Y=0.515 $X2=0 $Y2=0
cc_275 N_Y_c_347_n N_VGND_c_554_n 0.00158453f $X=1.325 $Y=0.515 $X2=0 $Y2=0
cc_276 N_Y_c_348_n N_VGND_c_554_n 0.022455f $X=2.17 $Y=1.095 $X2=0 $Y2=0
cc_277 N_Y_c_349_n N_VGND_c_554_n 0.0191425f $X=2.335 $Y=0.515 $X2=0 $Y2=0
cc_278 N_Y_c_349_n N_VGND_c_556_n 0.0145639f $X=2.335 $Y=0.515 $X2=0 $Y2=0
cc_279 N_Y_c_347_n N_VGND_c_558_n 0.0121141f $X=1.325 $Y=0.515 $X2=0 $Y2=0
cc_280 N_Y_c_349_n N_VGND_c_558_n 0.0119984f $X=2.335 $Y=0.515 $X2=0 $Y2=0
cc_281 N_Y_c_350_n N_VGND_c_558_n 0.0406621f $X=4 $Y=0.872 $X2=0 $Y2=0
cc_282 N_Y_c_350_n N_A_722_74#_M1001_d 0.00838011f $X=4 $Y=0.872 $X2=-0.19
+ $Y2=-0.245
cc_283 N_Y_M1001_s N_A_722_74#_c_605_n 0.00178571f $X=4.025 $Y=0.37 $X2=0 $Y2=0
cc_284 N_Y_c_350_n N_A_722_74#_c_605_n 0.0268535f $X=4 $Y=0.872 $X2=0 $Y2=0
cc_285 N_Y_c_353_n N_A_722_74#_c_605_n 0.0161432f $X=4.165 $Y=0.872 $X2=0 $Y2=0
cc_286 N_Y_c_353_n N_A_722_74#_c_608_n 0.00517071f $X=4.165 $Y=0.872 $X2=0 $Y2=0
cc_287 N_A_337_368#_c_416_n N_A_533_368#_M1010_s 0.00569965f $X=3.075 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_288 N_A_337_368#_c_416_n N_A_533_368#_c_439_n 0.0198097f $X=3.075 $Y=2.035
+ $X2=0 $Y2=0
cc_289 N_A_337_368#_M1010_d N_A_533_368#_c_440_n 0.00165831f $X=3.105 $Y=1.84
+ $X2=0 $Y2=0
cc_290 N_A_337_368#_c_417_n N_A_533_368#_c_440_n 0.0139027f $X=3.24 $Y=1.985
+ $X2=0 $Y2=0
cc_291 N_A_533_368#_c_456_n N_VPWR_M1012_d 0.00314376f $X=4.425 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_292 N_A_533_368#_c_465_n N_VPWR_M1002_s 0.00314031f $X=5.405 $Y=2.035 $X2=0
+ $Y2=0
cc_293 N_A_533_368#_c_440_n N_VPWR_c_495_n 0.0101219f $X=3.525 $Y=2.99 $X2=0
+ $Y2=0
cc_294 N_A_533_368#_c_456_n N_VPWR_c_495_n 0.0126919f $X=4.425 $Y=2.035 $X2=0
+ $Y2=0
cc_295 N_A_533_368#_c_442_n N_VPWR_c_495_n 0.022423f $X=4.59 $Y=2.445 $X2=0
+ $Y2=0
cc_296 N_A_533_368#_c_442_n N_VPWR_c_496_n 0.0234083f $X=4.59 $Y=2.445 $X2=0
+ $Y2=0
cc_297 N_A_533_368#_c_465_n N_VPWR_c_496_n 0.0170259f $X=5.405 $Y=2.035 $X2=0
+ $Y2=0
cc_298 N_A_533_368#_c_444_n N_VPWR_c_496_n 0.0234083f $X=5.49 $Y=2.4 $X2=0 $Y2=0
cc_299 N_A_533_368#_c_440_n N_VPWR_c_497_n 0.0623691f $X=3.525 $Y=2.99 $X2=0
+ $Y2=0
cc_300 N_A_533_368#_c_441_n N_VPWR_c_497_n 0.0200723f $X=2.905 $Y=2.99 $X2=0
+ $Y2=0
cc_301 N_A_533_368#_c_442_n N_VPWR_c_498_n 0.0109793f $X=4.59 $Y=2.445 $X2=0
+ $Y2=0
cc_302 N_A_533_368#_c_444_n N_VPWR_c_499_n 0.011066f $X=5.49 $Y=2.4 $X2=0 $Y2=0
cc_303 N_A_533_368#_c_440_n N_VPWR_c_494_n 0.0343566f $X=3.525 $Y=2.99 $X2=0
+ $Y2=0
cc_304 N_A_533_368#_c_441_n N_VPWR_c_494_n 0.0108858f $X=2.905 $Y=2.99 $X2=0
+ $Y2=0
cc_305 N_A_533_368#_c_442_n N_VPWR_c_494_n 0.00901959f $X=4.59 $Y=2.445 $X2=0
+ $Y2=0
cc_306 N_A_533_368#_c_444_n N_VPWR_c_494_n 0.00915947f $X=5.49 $Y=2.4 $X2=0
+ $Y2=0
cc_307 N_A_533_368#_c_443_n N_A_722_74#_c_607_n 0.00831718f $X=5.53 $Y=2.12
+ $X2=0 $Y2=0
cc_308 N_VGND_c_556_n N_A_722_74#_c_605_n 0.038121f $X=4.86 $Y=0 $X2=0 $Y2=0
cc_309 N_VGND_c_558_n N_A_722_74#_c_605_n 0.0321651f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_310 N_VGND_c_555_n N_A_722_74#_c_606_n 0.00989215f $X=5.03 $Y=0.675 $X2=0
+ $Y2=0
cc_311 N_VGND_c_556_n N_A_722_74#_c_606_n 0.00758556f $X=4.86 $Y=0 $X2=0 $Y2=0
cc_312 N_VGND_c_558_n N_A_722_74#_c_606_n 0.00627867f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_313 N_VGND_M1005_s N_A_722_74#_c_607_n 0.00187091f $X=4.885 $Y=0.37 $X2=0
+ $Y2=0
cc_314 N_VGND_c_555_n N_A_722_74#_c_607_n 0.0178913f $X=5.03 $Y=0.675 $X2=0
+ $Y2=0
cc_315 N_VGND_c_555_n N_A_722_74#_c_609_n 0.0183707f $X=5.03 $Y=0.675 $X2=0
+ $Y2=0
cc_316 N_VGND_c_557_n N_A_722_74#_c_609_n 0.011066f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_317 N_VGND_c_558_n N_A_722_74#_c_609_n 0.00915947f $X=5.52 $Y=0 $X2=0 $Y2=0

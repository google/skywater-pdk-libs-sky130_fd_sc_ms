* NGSPICE file created from sky130_fd_sc_ms__a221o_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 VPWR a_148_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=6.262e+11p pd=5.43e+06u as=2.912e+11p ps=2.76e+06u
M1001 a_313_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=0p ps=0u
M1002 VPWR A1 a_313_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_148_260# C1 VGND VNB nlowvt w=640000u l=150000u
+  ad=4.192e+11p pd=3.87e+06u as=8.64875e+11p ps=5.71e+06u
M1004 a_417_79# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1005 a_148_260# A1 a_417_79# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_148_260# C1 a_509_392# VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=5.6e+11p ps=5.12e+06u
M1007 VGND a_148_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.961e+11p ps=2.01e+06u
M1008 a_597_79# B1 a_148_260# VNB nlowvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1009 VGND B2 a_597_79# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_313_392# B1 a_509_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_509_392# B2 a_313_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__o2bb2a_4.pxi.spice
* Created: Fri Aug 28 17:59:47 2020
* 
x_PM_SKY130_FD_SC_MS__O2BB2A_4%B1 N_B1_M1022_g N_B1_M1000_g N_B1_M1001_g
+ N_B1_M1023_g B1 B1 N_B1_c_131_n N_B1_c_132_n PM_SKY130_FD_SC_MS__O2BB2A_4%B1
x_PM_SKY130_FD_SC_MS__O2BB2A_4%B2 N_B2_M1006_g N_B2_M1014_g N_B2_M1009_g
+ N_B2_M1016_g B2 B2 N_B2_c_186_n PM_SKY130_FD_SC_MS__O2BB2A_4%B2
x_PM_SKY130_FD_SC_MS__O2BB2A_4%A_476_48# N_A_476_48#_M1020_s N_A_476_48#_M1002_d
+ N_A_476_48#_M1005_g N_A_476_48#_M1019_g N_A_476_48#_M1010_g
+ N_A_476_48#_c_249_n N_A_476_48#_M1021_g N_A_476_48#_c_242_n
+ N_A_476_48#_c_243_n N_A_476_48#_c_244_n N_A_476_48#_c_245_n
+ N_A_476_48#_c_251_n N_A_476_48#_c_285_p N_A_476_48#_c_261_p
+ N_A_476_48#_c_246_n N_A_476_48#_c_247_n PM_SKY130_FD_SC_MS__O2BB2A_4%A_476_48#
x_PM_SKY130_FD_SC_MS__O2BB2A_4%A2_N N_A2_N_M1002_g N_A2_N_M1020_g A2_N
+ N_A2_N_c_325_n N_A2_N_c_326_n PM_SKY130_FD_SC_MS__O2BB2A_4%A2_N
x_PM_SKY130_FD_SC_MS__O2BB2A_4%A1_N N_A1_N_M1017_g N_A1_N_M1007_g A1_N
+ N_A1_N_c_365_n N_A1_N_c_366_n PM_SKY130_FD_SC_MS__O2BB2A_4%A1_N
x_PM_SKY130_FD_SC_MS__O2BB2A_4%A_313_392# N_A_313_392#_M1005_s
+ N_A_313_392#_M1006_d N_A_313_392#_M1010_s N_A_313_392#_c_403_n
+ N_A_313_392#_M1004_g N_A_313_392#_M1003_g N_A_313_392#_c_405_n
+ N_A_313_392#_M1011_g N_A_313_392#_c_407_n N_A_313_392#_M1008_g
+ N_A_313_392#_M1013_g N_A_313_392#_c_409_n N_A_313_392#_M1012_g
+ N_A_313_392#_c_410_n N_A_313_392#_c_411_n N_A_313_392#_M1018_g
+ N_A_313_392#_M1015_g N_A_313_392#_c_413_n N_A_313_392#_c_414_n
+ N_A_313_392#_c_440_n N_A_313_392#_c_441_n N_A_313_392#_c_445_n
+ N_A_313_392#_c_415_n N_A_313_392#_c_416_n N_A_313_392#_c_417_n
+ N_A_313_392#_c_418_n N_A_313_392#_c_419_n N_A_313_392#_c_512_p
+ N_A_313_392#_c_428_n N_A_313_392#_c_420_n N_A_313_392#_c_429_n
+ N_A_313_392#_c_430_n N_A_313_392#_c_421_n N_A_313_392#_c_422_n
+ PM_SKY130_FD_SC_MS__O2BB2A_4%A_313_392#
x_PM_SKY130_FD_SC_MS__O2BB2A_4%A_41_392# N_A_41_392#_M1000_s N_A_41_392#_M1001_s
+ N_A_41_392#_M1009_s N_A_41_392#_c_580_n N_A_41_392#_c_581_n
+ N_A_41_392#_c_582_n N_A_41_392#_c_583_n N_A_41_392#_c_599_n
+ N_A_41_392#_c_584_n N_A_41_392#_c_585_n N_A_41_392#_c_586_n
+ PM_SKY130_FD_SC_MS__O2BB2A_4%A_41_392#
x_PM_SKY130_FD_SC_MS__O2BB2A_4%VPWR N_VPWR_M1000_d N_VPWR_M1010_d N_VPWR_M1021_d
+ N_VPWR_M1007_d N_VPWR_M1011_d N_VPWR_M1015_d N_VPWR_c_629_n N_VPWR_c_630_n
+ N_VPWR_c_631_n N_VPWR_c_632_n N_VPWR_c_633_n N_VPWR_c_634_n N_VPWR_c_635_n
+ N_VPWR_c_636_n N_VPWR_c_637_n N_VPWR_c_638_n VPWR N_VPWR_c_639_n
+ N_VPWR_c_640_n N_VPWR_c_641_n N_VPWR_c_642_n N_VPWR_c_643_n N_VPWR_c_644_n
+ N_VPWR_c_645_n N_VPWR_c_628_n PM_SKY130_FD_SC_MS__O2BB2A_4%VPWR
x_PM_SKY130_FD_SC_MS__O2BB2A_4%X N_X_M1004_d N_X_M1012_d N_X_M1003_s N_X_M1013_s
+ N_X_c_731_n N_X_c_725_n N_X_c_727_n N_X_c_728_n N_X_c_729_n N_X_c_726_n
+ N_X_c_748_n N_X_c_730_n N_X_c_761_n N_X_c_765_n N_X_c_767_n X X
+ PM_SKY130_FD_SC_MS__O2BB2A_4%X
x_PM_SKY130_FD_SC_MS__O2BB2A_4%A_27_74# N_A_27_74#_M1022_s N_A_27_74#_M1023_s
+ N_A_27_74#_M1016_d N_A_27_74#_M1019_d N_A_27_74#_c_792_n N_A_27_74#_c_793_n
+ N_A_27_74#_c_794_n N_A_27_74#_c_795_n N_A_27_74#_c_796_n N_A_27_74#_c_797_n
+ N_A_27_74#_c_798_n PM_SKY130_FD_SC_MS__O2BB2A_4%A_27_74#
x_PM_SKY130_FD_SC_MS__O2BB2A_4%VGND N_VGND_M1022_d N_VGND_M1014_s N_VGND_M1017_d
+ N_VGND_M1008_s N_VGND_M1018_s N_VGND_c_845_n N_VGND_c_846_n N_VGND_c_847_n
+ N_VGND_c_848_n N_VGND_c_849_n N_VGND_c_850_n N_VGND_c_851_n VGND
+ N_VGND_c_852_n N_VGND_c_853_n N_VGND_c_854_n N_VGND_c_855_n N_VGND_c_856_n
+ N_VGND_c_857_n N_VGND_c_858_n N_VGND_c_859_n N_VGND_c_860_n
+ PM_SKY130_FD_SC_MS__O2BB2A_4%VGND
cc_1 VNB N_B1_M1022_g 0.0351242f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_2 VNB N_B1_M1000_g 0.00418093f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.46
cc_3 VNB N_B1_M1001_g 0.00309826f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=2.46
cc_4 VNB N_B1_M1023_g 0.0258723f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.69
cc_5 VNB N_B1_c_131_n 0.0184978f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.425
cc_6 VNB N_B1_c_132_n 0.0787933f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.425
cc_7 VNB N_B2_M1014_g 0.0354936f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.46
cc_8 VNB N_B2_M1016_g 0.0355932f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.69
cc_9 VNB B2 0.00338057f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_10 VNB N_B2_c_186_n 0.0323306f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.425
cc_11 VNB N_A_476_48#_M1005_g 0.0267856f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.59
cc_12 VNB N_A_476_48#_M1019_g 0.030921f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.26
cc_13 VNB N_A_476_48#_M1010_g 0.00203907f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_14 VNB N_A_476_48#_c_242_n 0.0463001f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.425
cc_15 VNB N_A_476_48#_c_243_n 0.00129542f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.425
cc_16 VNB N_A_476_48#_c_244_n 0.0182277f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.515
cc_17 VNB N_A_476_48#_c_245_n 0.00405041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_476_48#_c_246_n 0.00238033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_476_48#_c_247_n 0.0442713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A2_N_M1020_g 0.026815f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.46
cc_21 VNB N_A2_N_c_325_n 0.0260861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A2_N_c_326_n 0.00465481f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.26
cc_23 VNB N_A1_N_M1017_g 0.0250549f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_24 VNB N_A1_N_c_365_n 0.0278334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A1_N_c_366_n 0.00186123f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.26
cc_26 VNB N_A_313_392#_c_403_n 0.0197713f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=2.46
cc_27 VNB N_A_313_392#_M1003_g 0.00595357f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.69
cc_28 VNB N_A_313_392#_c_405_n 0.0235051f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_29 VNB N_A_313_392#_M1011_g 0.00643297f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.425
cc_30 VNB N_A_313_392#_c_407_n 0.0184166f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.425
cc_31 VNB N_A_313_392#_M1013_g 0.0055873f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.425
cc_32 VNB N_A_313_392#_c_409_n 0.0172383f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.425
cc_33 VNB N_A_313_392#_c_410_n 0.00993014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_313_392#_c_411_n 0.0199243f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.515
cc_35 VNB N_A_313_392#_M1015_g 0.0231638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_313_392#_c_413_n 0.0128144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_313_392#_c_414_n 0.028216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_313_392#_c_415_n 6.46475e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_313_392#_c_416_n 0.00866423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_313_392#_c_417_n 0.00697079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_313_392#_c_418_n 6.54855e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_313_392#_c_419_n 0.0117907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_313_392#_c_420_n 0.00239894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_313_392#_c_421_n 0.00379973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_313_392#_c_422_n 0.033721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VPWR_c_628_n 0.302998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_X_c_725_n 0.00327262f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.69
cc_48 VNB N_X_c_726_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.425
cc_49 VNB N_A_27_74#_c_792_n 0.0242911f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=0.69
cc_50 VNB N_A_27_74#_c_793_n 0.00325303f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_51 VNB N_A_27_74#_c_794_n 0.00919114f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_52 VNB N_A_27_74#_c_795_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.425
cc_53 VNB N_A_27_74#_c_796_n 0.0129155f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.425
cc_54 VNB N_A_27_74#_c_797_n 0.0104454f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.425
cc_55 VNB N_A_27_74#_c_798_n 0.00829653f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.425
cc_56 VNB N_VGND_c_845_n 0.00900728f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_57 VNB N_VGND_c_846_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_847_n 0.00571618f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.425
cc_59 VNB N_VGND_c_848_n 0.00682834f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.425
cc_60 VNB N_VGND_c_849_n 0.00517079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_850_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.515
cc_62 VNB N_VGND_c_851_n 0.0551317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_852_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_853_n 0.0645768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_854_n 0.0185379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_855_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_856_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_857_n 0.00613276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_858_n 0.0101972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_859_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_860_n 0.388386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VPB N_B1_M1000_g 0.0387008f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=2.46
cc_73 VPB N_B1_M1001_g 0.0277206f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=2.46
cc_74 VPB N_B1_c_131_n 0.0138762f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.425
cc_75 VPB N_B2_M1006_g 0.0217971f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.69
cc_76 VPB N_B2_M1009_g 0.0288064f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=2.46
cc_77 VPB B2 0.00317786f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_78 VPB N_B2_c_186_n 0.0201019f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.425
cc_79 VPB N_A_476_48#_M1010_g 0.0278439f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_80 VPB N_A_476_48#_c_249_n 0.0207897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_476_48#_c_242_n 0.00336932f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.425
cc_82 VPB N_A_476_48#_c_251_n 0.00141245f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.515
cc_83 VPB N_A2_N_M1002_g 0.0226102f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.69
cc_84 VPB N_A2_N_c_325_n 0.00559309f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A2_N_c_326_n 0.00303521f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=1.26
cc_86 VPB N_A1_N_M1007_g 0.0226023f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=2.46
cc_87 VPB N_A1_N_c_365_n 0.0056959f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A1_N_c_366_n 0.00373149f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=1.26
cc_89 VPB N_A_313_392#_M1003_g 0.0245816f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.69
cc_90 VPB N_A_313_392#_M1011_g 0.0225739f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.425
cc_91 VPB N_A_313_392#_M1013_g 0.0217989f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.425
cc_92 VPB N_A_313_392#_M1015_g 0.0274594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_313_392#_c_418_n 0.00140298f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_313_392#_c_428_n 0.00135969f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_313_392#_c_429_n 0.018068f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_313_392#_c_430_n 0.00265213f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_41_392#_c_580_n 0.00953141f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=2.46
cc_98 VPB N_A_41_392#_c_581_n 0.0352562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_41_392#_c_582_n 0.00229495f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=0.69
cc_100 VPB N_A_41_392#_c_583_n 0.0103719f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_41_392#_c_584_n 0.00643964f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_41_392#_c_585_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.425
cc_103 VPB N_A_41_392#_c_586_n 0.00599433f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.425
cc_104 VPB N_VPWR_c_629_n 0.00768638f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.425
cc_105 VPB N_VPWR_c_630_n 0.0254753f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.425
cc_106 VPB N_VPWR_c_631_n 0.0213455f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=1.425
cc_107 VPB N_VPWR_c_632_n 0.0275115f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_633_n 0.0179357f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.515
cc_109 VPB N_VPWR_c_634_n 0.00565985f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_635_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_636_n 0.0695549f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_637_n 0.020661f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_638_n 0.00631873f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_639_n 0.0407783f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_640_n 0.0209196f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_641_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_642_n 0.0255777f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_643_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_644_n 0.00631873f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_645_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_628_n 0.101746f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_X_c_727_n 0.00328511f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_X_c_728_n 0.00290991f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.425
cc_124 VPB N_X_c_729_n 0.00384241f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.425
cc_125 VPB N_X_c_730_n 0.00235902f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 N_B1_M1001_g N_B2_M1006_g 0.016003f $X=1.025 $Y=2.46 $X2=0 $Y2=0
cc_127 N_B1_M1023_g N_B2_M1014_g 0.0254685f $X=1.065 $Y=0.69 $X2=0 $Y2=0
cc_128 N_B1_c_131_n N_B2_M1014_g 0.00111826f $X=0.95 $Y=1.425 $X2=0 $Y2=0
cc_129 N_B1_c_132_n N_B2_M1014_g 0.00148703f $X=1.025 $Y=1.425 $X2=0 $Y2=0
cc_130 N_B1_c_131_n B2 0.0148123f $X=0.95 $Y=1.425 $X2=0 $Y2=0
cc_131 N_B1_c_132_n B2 3.55107e-19 $X=1.025 $Y=1.425 $X2=0 $Y2=0
cc_132 N_B1_c_131_n N_B2_c_186_n 0.00147947f $X=0.95 $Y=1.425 $X2=0 $Y2=0
cc_133 N_B1_c_132_n N_B2_c_186_n 0.016003f $X=1.025 $Y=1.425 $X2=0 $Y2=0
cc_134 N_B1_M1000_g N_A_41_392#_c_580_n 0.0014751f $X=0.575 $Y=2.46 $X2=0 $Y2=0
cc_135 N_B1_c_131_n N_A_41_392#_c_580_n 0.0298625f $X=0.95 $Y=1.425 $X2=0 $Y2=0
cc_136 N_B1_c_132_n N_A_41_392#_c_580_n 0.00155726f $X=1.025 $Y=1.425 $X2=0
+ $Y2=0
cc_137 N_B1_M1000_g N_A_41_392#_c_581_n 0.0121004f $X=0.575 $Y=2.46 $X2=0 $Y2=0
cc_138 N_B1_M1001_g N_A_41_392#_c_581_n 6.50516e-19 $X=1.025 $Y=2.46 $X2=0 $Y2=0
cc_139 N_B1_M1000_g N_A_41_392#_c_582_n 0.0129919f $X=0.575 $Y=2.46 $X2=0 $Y2=0
cc_140 N_B1_M1001_g N_A_41_392#_c_582_n 0.0129919f $X=1.025 $Y=2.46 $X2=0 $Y2=0
cc_141 N_B1_c_131_n N_A_41_392#_c_582_n 0.042435f $X=0.95 $Y=1.425 $X2=0 $Y2=0
cc_142 N_B1_c_132_n N_A_41_392#_c_582_n 4.12623e-19 $X=1.025 $Y=1.425 $X2=0
+ $Y2=0
cc_143 N_B1_M1001_g N_A_41_392#_c_583_n 0.00101522f $X=1.025 $Y=2.46 $X2=0 $Y2=0
cc_144 N_B1_c_131_n N_A_41_392#_c_583_n 0.00236117f $X=0.95 $Y=1.425 $X2=0 $Y2=0
cc_145 N_B1_c_132_n N_A_41_392#_c_583_n 8.21866e-19 $X=1.025 $Y=1.425 $X2=0
+ $Y2=0
cc_146 N_B1_M1000_g N_A_41_392#_c_599_n 6.26485e-19 $X=0.575 $Y=2.46 $X2=0 $Y2=0
cc_147 N_B1_M1001_g N_A_41_392#_c_599_n 0.0105282f $X=1.025 $Y=2.46 $X2=0 $Y2=0
cc_148 N_B1_M1001_g N_A_41_392#_c_585_n 0.00347836f $X=1.025 $Y=2.46 $X2=0 $Y2=0
cc_149 N_B1_M1000_g N_VPWR_c_629_n 0.0027763f $X=0.575 $Y=2.46 $X2=0 $Y2=0
cc_150 N_B1_M1001_g N_VPWR_c_629_n 0.00120619f $X=1.025 $Y=2.46 $X2=0 $Y2=0
cc_151 N_B1_M1001_g N_VPWR_c_639_n 0.00517089f $X=1.025 $Y=2.46 $X2=0 $Y2=0
cc_152 N_B1_M1000_g N_VPWR_c_642_n 0.005209f $X=0.575 $Y=2.46 $X2=0 $Y2=0
cc_153 N_B1_M1000_g N_VPWR_c_628_n 0.00986227f $X=0.575 $Y=2.46 $X2=0 $Y2=0
cc_154 N_B1_M1001_g N_VPWR_c_628_n 0.00977588f $X=1.025 $Y=2.46 $X2=0 $Y2=0
cc_155 N_B1_M1022_g N_A_27_74#_c_792_n 0.00818668f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_156 N_B1_M1023_g N_A_27_74#_c_792_n 6.10854e-19 $X=1.065 $Y=0.69 $X2=0 $Y2=0
cc_157 N_B1_M1022_g N_A_27_74#_c_793_n 0.0118691f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_158 N_B1_M1023_g N_A_27_74#_c_793_n 0.0118691f $X=1.065 $Y=0.69 $X2=0 $Y2=0
cc_159 N_B1_c_131_n N_A_27_74#_c_793_n 0.0510846f $X=0.95 $Y=1.425 $X2=0 $Y2=0
cc_160 N_B1_c_132_n N_A_27_74#_c_793_n 0.00597192f $X=1.025 $Y=1.425 $X2=0 $Y2=0
cc_161 N_B1_M1022_g N_A_27_74#_c_794_n 0.00235019f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_162 N_B1_c_131_n N_A_27_74#_c_794_n 0.0285737f $X=0.95 $Y=1.425 $X2=0 $Y2=0
cc_163 N_B1_c_132_n N_A_27_74#_c_794_n 0.00710517f $X=1.025 $Y=1.425 $X2=0 $Y2=0
cc_164 N_B1_M1023_g N_A_27_74#_c_795_n 0.00517605f $X=1.065 $Y=0.69 $X2=0 $Y2=0
cc_165 N_B1_M1022_g N_A_27_74#_c_797_n 4.37003e-19 $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_166 N_B1_M1023_g N_A_27_74#_c_797_n 0.00535077f $X=1.065 $Y=0.69 $X2=0 $Y2=0
cc_167 N_B1_M1022_g N_VGND_c_845_n 0.00567941f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_168 N_B1_M1023_g N_VGND_c_845_n 0.00429749f $X=1.065 $Y=0.69 $X2=0 $Y2=0
cc_169 N_B1_M1023_g N_VGND_c_846_n 0.00434272f $X=1.065 $Y=0.69 $X2=0 $Y2=0
cc_170 N_B1_M1022_g N_VGND_c_852_n 0.00434272f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_171 N_B1_M1022_g N_VGND_c_860_n 0.00824951f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_172 N_B1_M1023_g N_VGND_c_860_n 0.00821391f $X=1.065 $Y=0.69 $X2=0 $Y2=0
cc_173 N_B2_M1016_g N_A_476_48#_M1005_g 0.0360783f $X=1.995 $Y=0.69 $X2=0 $Y2=0
cc_174 B2 N_A_476_48#_M1010_g 0.00294262f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_175 N_B2_c_186_n N_A_476_48#_M1010_g 0.00161561f $X=1.995 $Y=1.615 $X2=0
+ $Y2=0
cc_176 N_B2_M1016_g N_A_476_48#_c_243_n 7.28417e-19 $X=1.995 $Y=0.69 $X2=0 $Y2=0
cc_177 B2 N_A_476_48#_c_243_n 0.0132888f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_178 B2 N_A_476_48#_c_247_n 7.85605e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_179 N_B2_c_186_n N_A_476_48#_c_247_n 0.00615356f $X=1.995 $Y=1.615 $X2=0
+ $Y2=0
cc_180 B2 N_A_313_392#_c_428_n 0.0143383f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_181 N_B2_c_186_n N_A_313_392#_c_428_n 0.00211633f $X=1.995 $Y=1.615 $X2=0
+ $Y2=0
cc_182 N_B2_M1016_g N_A_313_392#_c_420_n 0.00106797f $X=1.995 $Y=0.69 $X2=0
+ $Y2=0
cc_183 N_B2_M1009_g N_A_313_392#_c_429_n 0.0164637f $X=1.925 $Y=2.46 $X2=0 $Y2=0
cc_184 B2 N_A_313_392#_c_429_n 0.0366734f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_185 N_B2_c_186_n N_A_313_392#_c_429_n 0.00301926f $X=1.995 $Y=1.615 $X2=0
+ $Y2=0
cc_186 N_B2_M1006_g N_A_41_392#_c_583_n 0.00357165f $X=1.475 $Y=2.46 $X2=0 $Y2=0
cc_187 N_B2_M1006_g N_A_41_392#_c_599_n 0.0105282f $X=1.475 $Y=2.46 $X2=0 $Y2=0
cc_188 N_B2_M1009_g N_A_41_392#_c_599_n 6.26485e-19 $X=1.925 $Y=2.46 $X2=0 $Y2=0
cc_189 N_B2_M1006_g N_A_41_392#_c_584_n 0.0116345f $X=1.475 $Y=2.46 $X2=0 $Y2=0
cc_190 N_B2_M1009_g N_A_41_392#_c_584_n 0.014552f $X=1.925 $Y=2.46 $X2=0 $Y2=0
cc_191 N_B2_M1006_g N_A_41_392#_c_585_n 0.001916f $X=1.475 $Y=2.46 $X2=0 $Y2=0
cc_192 N_B2_M1006_g N_A_41_392#_c_586_n 5.73047e-19 $X=1.475 $Y=2.46 $X2=0 $Y2=0
cc_193 N_B2_M1009_g N_A_41_392#_c_586_n 0.00892729f $X=1.925 $Y=2.46 $X2=0 $Y2=0
cc_194 N_B2_M1009_g N_VPWR_c_630_n 0.00190837f $X=1.925 $Y=2.46 $X2=0 $Y2=0
cc_195 N_B2_M1006_g N_VPWR_c_639_n 0.00333896f $X=1.475 $Y=2.46 $X2=0 $Y2=0
cc_196 N_B2_M1009_g N_VPWR_c_639_n 0.00333896f $X=1.925 $Y=2.46 $X2=0 $Y2=0
cc_197 N_B2_M1006_g N_VPWR_c_628_n 0.00422796f $X=1.475 $Y=2.46 $X2=0 $Y2=0
cc_198 N_B2_M1009_g N_VPWR_c_628_n 0.00427818f $X=1.925 $Y=2.46 $X2=0 $Y2=0
cc_199 N_B2_M1014_g N_A_27_74#_c_795_n 0.00637865f $X=1.495 $Y=0.69 $X2=0 $Y2=0
cc_200 N_B2_M1016_g N_A_27_74#_c_795_n 6.25537e-19 $X=1.995 $Y=0.69 $X2=0 $Y2=0
cc_201 N_B2_M1014_g N_A_27_74#_c_796_n 0.0141322f $X=1.495 $Y=0.69 $X2=0 $Y2=0
cc_202 N_B2_M1016_g N_A_27_74#_c_796_n 0.0161338f $X=1.995 $Y=0.69 $X2=0 $Y2=0
cc_203 B2 N_A_27_74#_c_796_n 0.0358207f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_204 N_B2_c_186_n N_A_27_74#_c_796_n 0.00507416f $X=1.995 $Y=1.615 $X2=0 $Y2=0
cc_205 N_B2_M1014_g N_A_27_74#_c_797_n 0.00292768f $X=1.495 $Y=0.69 $X2=0 $Y2=0
cc_206 N_B2_c_186_n N_A_27_74#_c_797_n 0.00138383f $X=1.995 $Y=1.615 $X2=0 $Y2=0
cc_207 N_B2_M1014_g N_VGND_c_846_n 0.00434272f $X=1.495 $Y=0.69 $X2=0 $Y2=0
cc_208 N_B2_M1014_g N_VGND_c_847_n 0.00312943f $X=1.495 $Y=0.69 $X2=0 $Y2=0
cc_209 N_B2_M1016_g N_VGND_c_847_n 0.00910301f $X=1.995 $Y=0.69 $X2=0 $Y2=0
cc_210 N_B2_M1016_g N_VGND_c_853_n 0.00383152f $X=1.995 $Y=0.69 $X2=0 $Y2=0
cc_211 N_B2_M1014_g N_VGND_c_860_n 0.00433099f $X=1.495 $Y=0.69 $X2=0 $Y2=0
cc_212 N_B2_M1016_g N_VGND_c_860_n 0.00371743f $X=1.995 $Y=0.69 $X2=0 $Y2=0
cc_213 N_A_476_48#_c_242_n N_A2_N_M1002_g 0.0294959f $X=3.365 $Y=1.465 $X2=0
+ $Y2=0
cc_214 N_A_476_48#_c_251_n N_A2_N_M1002_g 0.00345537f $X=3.59 $Y=1.95 $X2=0
+ $Y2=0
cc_215 N_A_476_48#_c_261_p N_A2_N_M1002_g 0.0159042f $X=4.3 $Y=2.115 $X2=0 $Y2=0
cc_216 N_A_476_48#_c_242_n N_A2_N_M1020_g 8.73622e-19 $X=3.365 $Y=1.465 $X2=0
+ $Y2=0
cc_217 N_A_476_48#_c_244_n N_A2_N_M1020_g 0.0075272f $X=3.59 $Y=1.13 $X2=0 $Y2=0
cc_218 N_A_476_48#_c_245_n N_A2_N_M1020_g 0.0047775f $X=3.59 $Y=1.3 $X2=0 $Y2=0
cc_219 N_A_476_48#_c_246_n N_A2_N_M1020_g 0.00119678f $X=3.59 $Y=1.465 $X2=0
+ $Y2=0
cc_220 N_A_476_48#_c_242_n N_A2_N_c_325_n 0.0116234f $X=3.365 $Y=1.465 $X2=0
+ $Y2=0
cc_221 N_A_476_48#_c_244_n N_A2_N_c_325_n 0.0013179f $X=3.59 $Y=1.13 $X2=0 $Y2=0
cc_222 N_A_476_48#_c_251_n N_A2_N_c_325_n 3.20056e-19 $X=3.59 $Y=1.95 $X2=0
+ $Y2=0
cc_223 N_A_476_48#_c_261_p N_A2_N_c_325_n 6.7849e-19 $X=4.3 $Y=2.115 $X2=0 $Y2=0
cc_224 N_A_476_48#_c_246_n N_A2_N_c_325_n 0.00215032f $X=3.59 $Y=1.465 $X2=0
+ $Y2=0
cc_225 N_A_476_48#_c_242_n N_A2_N_c_326_n 6.17993e-19 $X=3.365 $Y=1.465 $X2=0
+ $Y2=0
cc_226 N_A_476_48#_c_244_n N_A2_N_c_326_n 0.012719f $X=3.59 $Y=1.13 $X2=0 $Y2=0
cc_227 N_A_476_48#_c_251_n N_A2_N_c_326_n 0.0117018f $X=3.59 $Y=1.95 $X2=0 $Y2=0
cc_228 N_A_476_48#_c_261_p N_A2_N_c_326_n 0.0244388f $X=4.3 $Y=2.115 $X2=0 $Y2=0
cc_229 N_A_476_48#_c_246_n N_A2_N_c_326_n 0.0237088f $X=3.59 $Y=1.465 $X2=0
+ $Y2=0
cc_230 N_A_476_48#_c_244_n N_A1_N_M1017_g 2.65127e-19 $X=3.59 $Y=1.13 $X2=0
+ $Y2=0
cc_231 N_A_476_48#_c_261_p N_A1_N_M1007_g 0.00665754f $X=4.3 $Y=2.115 $X2=0
+ $Y2=0
cc_232 N_A_476_48#_c_261_p N_A1_N_c_366_n 0.00309929f $X=4.3 $Y=2.115 $X2=0
+ $Y2=0
cc_233 N_A_476_48#_c_261_p N_A_313_392#_M1003_g 2.82705e-19 $X=4.3 $Y=2.115
+ $X2=0 $Y2=0
cc_234 N_A_476_48#_M1019_g N_A_313_392#_c_414_n 0.0106608f $X=2.92 $Y=0.69 $X2=0
+ $Y2=0
cc_235 N_A_476_48#_c_244_n N_A_313_392#_c_414_n 0.0264525f $X=3.59 $Y=1.13 $X2=0
+ $Y2=0
cc_236 N_A_476_48#_M1010_g N_A_313_392#_c_440_n 0.00471494f $X=2.935 $Y=2.26
+ $X2=0 $Y2=0
cc_237 N_A_476_48#_M1002_d N_A_313_392#_c_441_n 0.00460881f $X=4.165 $Y=1.84
+ $X2=0 $Y2=0
cc_238 N_A_476_48#_c_249_n N_A_313_392#_c_441_n 0.0175651f $X=3.455 $Y=1.72
+ $X2=0 $Y2=0
cc_239 N_A_476_48#_c_285_p N_A_313_392#_c_441_n 0.00889918f $X=3.675 $Y=2.115
+ $X2=0 $Y2=0
cc_240 N_A_476_48#_c_261_p N_A_313_392#_c_441_n 0.046138f $X=4.3 $Y=2.115 $X2=0
+ $Y2=0
cc_241 N_A_476_48#_M1010_g N_A_313_392#_c_445_n 0.00163952f $X=2.935 $Y=2.26
+ $X2=0 $Y2=0
cc_242 N_A_476_48#_c_244_n N_A_313_392#_c_417_n 0.00731399f $X=3.59 $Y=1.13
+ $X2=0 $Y2=0
cc_243 N_A_476_48#_c_261_p N_A_313_392#_c_418_n 0.0120728f $X=4.3 $Y=2.115 $X2=0
+ $Y2=0
cc_244 N_A_476_48#_M1005_g N_A_313_392#_c_420_n 0.00814829f $X=2.455 $Y=0.69
+ $X2=0 $Y2=0
cc_245 N_A_476_48#_M1019_g N_A_313_392#_c_420_n 5.51117e-19 $X=2.92 $Y=0.69
+ $X2=0 $Y2=0
cc_246 N_A_476_48#_M1010_g N_A_313_392#_c_429_n 0.0150392f $X=2.935 $Y=2.26
+ $X2=0 $Y2=0
cc_247 N_A_476_48#_c_243_n N_A_313_392#_c_429_n 0.0213716f $X=3.505 $Y=1.465
+ $X2=0 $Y2=0
cc_248 N_A_476_48#_c_247_n N_A_313_392#_c_429_n 0.0109604f $X=3.025 $Y=1.465
+ $X2=0 $Y2=0
cc_249 N_A_476_48#_M1010_g N_A_313_392#_c_430_n 0.00947676f $X=2.935 $Y=2.26
+ $X2=0 $Y2=0
cc_250 N_A_476_48#_c_249_n N_A_313_392#_c_430_n 0.00185905f $X=3.455 $Y=1.72
+ $X2=0 $Y2=0
cc_251 N_A_476_48#_c_242_n N_A_313_392#_c_430_n 0.0036026f $X=3.365 $Y=1.465
+ $X2=0 $Y2=0
cc_252 N_A_476_48#_c_243_n N_A_313_392#_c_430_n 0.024598f $X=3.505 $Y=1.465
+ $X2=0 $Y2=0
cc_253 N_A_476_48#_c_251_n N_A_313_392#_c_430_n 0.00511463f $X=3.59 $Y=1.95
+ $X2=0 $Y2=0
cc_254 N_A_476_48#_M1010_g N_A_41_392#_c_586_n 0.00186151f $X=2.935 $Y=2.26
+ $X2=0 $Y2=0
cc_255 N_A_476_48#_c_251_n N_VPWR_M1021_d 0.00141422f $X=3.59 $Y=1.95 $X2=0
+ $Y2=0
cc_256 N_A_476_48#_c_285_p N_VPWR_M1021_d 7.9873e-19 $X=3.675 $Y=2.115 $X2=0
+ $Y2=0
cc_257 N_A_476_48#_c_261_p N_VPWR_M1021_d 0.0119464f $X=4.3 $Y=2.115 $X2=0 $Y2=0
cc_258 N_A_476_48#_M1010_g N_VPWR_c_630_n 0.01175f $X=2.935 $Y=2.26 $X2=0 $Y2=0
cc_259 N_A_476_48#_c_249_n N_VPWR_c_630_n 0.00107061f $X=3.455 $Y=1.72 $X2=0
+ $Y2=0
cc_260 N_A_476_48#_M1010_g N_VPWR_c_631_n 0.00401533f $X=2.935 $Y=2.26 $X2=0
+ $Y2=0
cc_261 N_A_476_48#_c_249_n N_VPWR_c_631_n 0.00378791f $X=3.455 $Y=1.72 $X2=0
+ $Y2=0
cc_262 N_A_476_48#_c_249_n N_VPWR_c_632_n 5.86893e-19 $X=3.455 $Y=1.72 $X2=0
+ $Y2=0
cc_263 N_A_476_48#_M1010_g N_VPWR_c_628_n 0.00465661f $X=2.935 $Y=2.26 $X2=0
+ $Y2=0
cc_264 N_A_476_48#_c_249_n N_VPWR_c_628_n 0.00555093f $X=3.455 $Y=1.72 $X2=0
+ $Y2=0
cc_265 N_A_476_48#_M1005_g N_A_27_74#_c_796_n 0.0179232f $X=2.455 $Y=0.69 $X2=0
+ $Y2=0
cc_266 N_A_476_48#_M1019_g N_A_27_74#_c_796_n 0.015014f $X=2.92 $Y=0.69 $X2=0
+ $Y2=0
cc_267 N_A_476_48#_c_243_n N_A_27_74#_c_796_n 0.0338384f $X=3.505 $Y=1.465 $X2=0
+ $Y2=0
cc_268 N_A_476_48#_c_247_n N_A_27_74#_c_796_n 0.00325692f $X=3.025 $Y=1.465
+ $X2=0 $Y2=0
cc_269 N_A_476_48#_M1019_g N_A_27_74#_c_798_n 0.00159024f $X=2.92 $Y=0.69 $X2=0
+ $Y2=0
cc_270 N_A_476_48#_c_243_n N_A_27_74#_c_798_n 0.0229645f $X=3.505 $Y=1.465 $X2=0
+ $Y2=0
cc_271 N_A_476_48#_c_244_n N_A_27_74#_c_798_n 0.0272649f $X=3.59 $Y=1.13 $X2=0
+ $Y2=0
cc_272 N_A_476_48#_c_247_n N_A_27_74#_c_798_n 0.00800385f $X=3.025 $Y=1.465
+ $X2=0 $Y2=0
cc_273 N_A_476_48#_M1005_g N_VGND_c_847_n 0.00115316f $X=2.455 $Y=0.69 $X2=0
+ $Y2=0
cc_274 N_A_476_48#_M1005_g N_VGND_c_853_n 0.0043213f $X=2.455 $Y=0.69 $X2=0
+ $Y2=0
cc_275 N_A_476_48#_M1019_g N_VGND_c_853_n 0.00278271f $X=2.92 $Y=0.69 $X2=0
+ $Y2=0
cc_276 N_A_476_48#_M1005_g N_VGND_c_860_n 0.00434917f $X=2.455 $Y=0.69 $X2=0
+ $Y2=0
cc_277 N_A_476_48#_M1019_g N_VGND_c_860_n 0.00358767f $X=2.92 $Y=0.69 $X2=0
+ $Y2=0
cc_278 N_A2_N_M1020_g N_A1_N_M1017_g 0.0330395f $X=4.1 $Y=0.79 $X2=0 $Y2=0
cc_279 N_A2_N_M1002_g N_A1_N_M1007_g 0.0379102f $X=4.075 $Y=2.26 $X2=0 $Y2=0
cc_280 N_A2_N_c_326_n N_A1_N_M1007_g 3.57706e-19 $X=4.01 $Y=1.515 $X2=0 $Y2=0
cc_281 N_A2_N_c_325_n N_A1_N_c_365_n 0.0330395f $X=4.01 $Y=1.515 $X2=0 $Y2=0
cc_282 N_A2_N_c_326_n N_A1_N_c_365_n 0.00202352f $X=4.01 $Y=1.515 $X2=0 $Y2=0
cc_283 N_A2_N_M1002_g N_A1_N_c_366_n 3.46097e-19 $X=4.075 $Y=2.26 $X2=0 $Y2=0
cc_284 N_A2_N_c_325_n N_A1_N_c_366_n 4.06701e-19 $X=4.01 $Y=1.515 $X2=0 $Y2=0
cc_285 N_A2_N_c_326_n N_A1_N_c_366_n 0.0286239f $X=4.01 $Y=1.515 $X2=0 $Y2=0
cc_286 N_A2_N_M1020_g N_A_313_392#_c_414_n 0.0127071f $X=4.1 $Y=0.79 $X2=0 $Y2=0
cc_287 N_A2_N_M1002_g N_A_313_392#_c_441_n 0.0135494f $X=4.075 $Y=2.26 $X2=0
+ $Y2=0
cc_288 N_A2_N_M1020_g N_A_313_392#_c_415_n 0.00292575f $X=4.1 $Y=0.79 $X2=0
+ $Y2=0
cc_289 N_A2_N_M1020_g N_A_313_392#_c_417_n 7.02683e-19 $X=4.1 $Y=0.79 $X2=0
+ $Y2=0
cc_290 N_A2_N_M1002_g N_VPWR_c_632_n 5.86893e-19 $X=4.075 $Y=2.26 $X2=0 $Y2=0
cc_291 N_A2_N_M1002_g N_VPWR_c_637_n 0.00378791f $X=4.075 $Y=2.26 $X2=0 $Y2=0
cc_292 N_A2_N_M1002_g N_VPWR_c_628_n 0.00555093f $X=4.075 $Y=2.26 $X2=0 $Y2=0
cc_293 N_A2_N_M1020_g N_A_27_74#_c_798_n 0.0015342f $X=4.1 $Y=0.79 $X2=0 $Y2=0
cc_294 N_A2_N_M1020_g N_VGND_c_853_n 7.64118e-19 $X=4.1 $Y=0.79 $X2=0 $Y2=0
cc_295 N_A1_N_M1017_g N_A_313_392#_c_403_n 0.020147f $X=4.49 $Y=0.79 $X2=0 $Y2=0
cc_296 N_A1_N_M1007_g N_A_313_392#_M1003_g 0.0267922f $X=4.525 $Y=2.26 $X2=0
+ $Y2=0
cc_297 N_A1_N_c_366_n N_A_313_392#_M1003_g 2.83492e-19 $X=4.58 $Y=1.515 $X2=0
+ $Y2=0
cc_298 N_A1_N_M1017_g N_A_313_392#_c_414_n 6.54318e-19 $X=4.49 $Y=0.79 $X2=0
+ $Y2=0
cc_299 N_A1_N_M1007_g N_A_313_392#_c_441_n 0.0158247f $X=4.525 $Y=2.26 $X2=0
+ $Y2=0
cc_300 N_A1_N_c_366_n N_A_313_392#_c_441_n 0.00656442f $X=4.58 $Y=1.515 $X2=0
+ $Y2=0
cc_301 N_A1_N_M1017_g N_A_313_392#_c_415_n 0.00208925f $X=4.49 $Y=0.79 $X2=0
+ $Y2=0
cc_302 N_A1_N_M1017_g N_A_313_392#_c_416_n 0.0143138f $X=4.49 $Y=0.79 $X2=0
+ $Y2=0
cc_303 N_A1_N_c_365_n N_A_313_392#_c_416_n 0.00117988f $X=4.58 $Y=1.515 $X2=0
+ $Y2=0
cc_304 N_A1_N_c_366_n N_A_313_392#_c_416_n 0.0195571f $X=4.58 $Y=1.515 $X2=0
+ $Y2=0
cc_305 N_A1_N_M1007_g N_A_313_392#_c_418_n 0.00945892f $X=4.525 $Y=2.26 $X2=0
+ $Y2=0
cc_306 N_A1_N_c_365_n N_A_313_392#_c_419_n 0.0123767f $X=4.58 $Y=1.515 $X2=0
+ $Y2=0
cc_307 N_A1_N_c_366_n N_A_313_392#_c_419_n 3.32121e-19 $X=4.58 $Y=1.515 $X2=0
+ $Y2=0
cc_308 N_A1_N_M1017_g N_A_313_392#_c_421_n 0.00435133f $X=4.49 $Y=0.79 $X2=0
+ $Y2=0
cc_309 N_A1_N_c_365_n N_A_313_392#_c_421_n 0.00216596f $X=4.58 $Y=1.515 $X2=0
+ $Y2=0
cc_310 N_A1_N_c_366_n N_A_313_392#_c_421_n 0.0326915f $X=4.58 $Y=1.515 $X2=0
+ $Y2=0
cc_311 N_A1_N_M1007_g N_VPWR_c_633_n 5.86893e-19 $X=4.525 $Y=2.26 $X2=0 $Y2=0
cc_312 N_A1_N_M1007_g N_VPWR_c_637_n 0.00378791f $X=4.525 $Y=2.26 $X2=0 $Y2=0
cc_313 N_A1_N_M1007_g N_VPWR_c_628_n 0.00555093f $X=4.525 $Y=2.26 $X2=0 $Y2=0
cc_314 N_A1_N_M1017_g N_VGND_c_848_n 0.0129587f $X=4.49 $Y=0.79 $X2=0 $Y2=0
cc_315 N_A1_N_M1017_g N_VGND_c_853_n 0.00421418f $X=4.49 $Y=0.79 $X2=0 $Y2=0
cc_316 N_A1_N_M1017_g N_VGND_c_860_n 0.00432128f $X=4.49 $Y=0.79 $X2=0 $Y2=0
cc_317 N_A_313_392#_c_429_n N_A_41_392#_M1009_s 0.0032506f $X=2.995 $Y=1.985
+ $X2=0 $Y2=0
cc_318 N_A_313_392#_c_428_n N_A_41_392#_c_583_n 0.00668359f $X=1.7 $Y=2.115
+ $X2=0 $Y2=0
cc_319 N_A_313_392#_M1006_d N_A_41_392#_c_584_n 0.00165831f $X=1.565 $Y=1.96
+ $X2=0 $Y2=0
cc_320 N_A_313_392#_c_428_n N_A_41_392#_c_584_n 0.0118736f $X=1.7 $Y=2.115 $X2=0
+ $Y2=0
cc_321 N_A_313_392#_c_429_n N_A_41_392#_c_586_n 0.0219147f $X=2.995 $Y=1.985
+ $X2=0 $Y2=0
cc_322 N_A_313_392#_c_429_n N_VPWR_M1010_d 0.00604501f $X=2.995 $Y=1.985 $X2=0
+ $Y2=0
cc_323 N_A_313_392#_c_441_n N_VPWR_M1021_d 0.00757752f $X=4.915 $Y=2.535 $X2=0
+ $Y2=0
cc_324 N_A_313_392#_c_441_n N_VPWR_M1007_d 0.012135f $X=4.915 $Y=2.535 $X2=0
+ $Y2=0
cc_325 N_A_313_392#_c_418_n N_VPWR_M1007_d 0.00797294f $X=5 $Y=2.45 $X2=0 $Y2=0
cc_326 N_A_313_392#_c_440_n N_VPWR_c_630_n 0.00634453f $X=3.25 $Y=2.45 $X2=0
+ $Y2=0
cc_327 N_A_313_392#_c_445_n N_VPWR_c_630_n 0.0093134f $X=3.335 $Y=2.535 $X2=0
+ $Y2=0
cc_328 N_A_313_392#_c_429_n N_VPWR_c_630_n 0.0194052f $X=2.995 $Y=1.985 $X2=0
+ $Y2=0
cc_329 N_A_313_392#_c_441_n N_VPWR_c_631_n 0.00316105f $X=4.915 $Y=2.535 $X2=0
+ $Y2=0
cc_330 N_A_313_392#_c_445_n N_VPWR_c_631_n 0.00251418f $X=3.335 $Y=2.535 $X2=0
+ $Y2=0
cc_331 N_A_313_392#_c_441_n N_VPWR_c_632_n 0.0255558f $X=4.915 $Y=2.535 $X2=0
+ $Y2=0
cc_332 N_A_313_392#_M1003_g N_VPWR_c_633_n 0.00828811f $X=5.145 $Y=2.4 $X2=0
+ $Y2=0
cc_333 N_A_313_392#_c_441_n N_VPWR_c_633_n 0.0260806f $X=4.915 $Y=2.535 $X2=0
+ $Y2=0
cc_334 N_A_313_392#_M1003_g N_VPWR_c_634_n 7.08086e-19 $X=5.145 $Y=2.4 $X2=0
+ $Y2=0
cc_335 N_A_313_392#_M1011_g N_VPWR_c_634_n 0.0151804f $X=5.695 $Y=2.4 $X2=0
+ $Y2=0
cc_336 N_A_313_392#_M1013_g N_VPWR_c_634_n 0.00194999f $X=6.195 $Y=2.4 $X2=0
+ $Y2=0
cc_337 N_A_313_392#_M1015_g N_VPWR_c_636_n 0.00550375f $X=6.65 $Y=2.4 $X2=0
+ $Y2=0
cc_338 N_A_313_392#_c_441_n N_VPWR_c_637_n 0.0090807f $X=4.915 $Y=2.535 $X2=0
+ $Y2=0
cc_339 N_A_313_392#_M1003_g N_VPWR_c_640_n 0.00528256f $X=5.145 $Y=2.4 $X2=0
+ $Y2=0
cc_340 N_A_313_392#_M1011_g N_VPWR_c_640_n 0.00460063f $X=5.695 $Y=2.4 $X2=0
+ $Y2=0
cc_341 N_A_313_392#_c_441_n N_VPWR_c_640_n 8.84959e-19 $X=4.915 $Y=2.535 $X2=0
+ $Y2=0
cc_342 N_A_313_392#_M1013_g N_VPWR_c_641_n 0.005209f $X=6.195 $Y=2.4 $X2=0 $Y2=0
cc_343 N_A_313_392#_M1015_g N_VPWR_c_641_n 0.00526565f $X=6.65 $Y=2.4 $X2=0
+ $Y2=0
cc_344 N_A_313_392#_M1003_g N_VPWR_c_628_n 0.00999343f $X=5.145 $Y=2.4 $X2=0
+ $Y2=0
cc_345 N_A_313_392#_M1011_g N_VPWR_c_628_n 0.00909486f $X=5.695 $Y=2.4 $X2=0
+ $Y2=0
cc_346 N_A_313_392#_M1013_g N_VPWR_c_628_n 0.00982133f $X=6.195 $Y=2.4 $X2=0
+ $Y2=0
cc_347 N_A_313_392#_M1015_g N_VPWR_c_628_n 0.0100376f $X=6.65 $Y=2.4 $X2=0 $Y2=0
cc_348 N_A_313_392#_c_441_n N_VPWR_c_628_n 0.0315436f $X=4.915 $Y=2.535 $X2=0
+ $Y2=0
cc_349 N_A_313_392#_c_445_n N_VPWR_c_628_n 0.00479577f $X=3.335 $Y=2.535 $X2=0
+ $Y2=0
cc_350 N_A_313_392#_c_405_n N_X_c_731_n 0.00591958f $X=5.605 $Y=1.385 $X2=0
+ $Y2=0
cc_351 N_A_313_392#_c_512_p N_X_c_731_n 0.0264591f $X=5.9 $Y=1.385 $X2=0 $Y2=0
cc_352 N_A_313_392#_c_403_n N_X_c_725_n 0.00285666f $X=5.13 $Y=1.22 $X2=0 $Y2=0
cc_353 N_A_313_392#_c_407_n N_X_c_725_n 0.00288393f $X=5.705 $Y=1.22 $X2=0 $Y2=0
cc_354 N_A_313_392#_M1003_g N_X_c_727_n 5.15122e-19 $X=5.145 $Y=2.4 $X2=0 $Y2=0
cc_355 N_A_313_392#_M1011_g N_X_c_727_n 4.86047e-19 $X=5.695 $Y=2.4 $X2=0 $Y2=0
cc_356 N_A_313_392#_M1011_g N_X_c_728_n 0.0161211f $X=5.695 $Y=2.4 $X2=0 $Y2=0
cc_357 N_A_313_392#_M1013_g N_X_c_728_n 0.0154236f $X=6.195 $Y=2.4 $X2=0 $Y2=0
cc_358 N_A_313_392#_c_512_p N_X_c_728_n 0.0353287f $X=5.9 $Y=1.385 $X2=0 $Y2=0
cc_359 N_A_313_392#_c_422_n N_X_c_728_n 0.00313888f $X=6.285 $Y=1.385 $X2=0
+ $Y2=0
cc_360 N_A_313_392#_M1003_g N_X_c_729_n 0.00121619f $X=5.145 $Y=2.4 $X2=0 $Y2=0
cc_361 N_A_313_392#_c_405_n N_X_c_729_n 0.00442617f $X=5.605 $Y=1.385 $X2=0
+ $Y2=0
cc_362 N_A_313_392#_c_418_n N_X_c_729_n 0.0113363f $X=5 $Y=2.45 $X2=0 $Y2=0
cc_363 N_A_313_392#_c_512_p N_X_c_729_n 0.0278328f $X=5.9 $Y=1.385 $X2=0 $Y2=0
cc_364 N_A_313_392#_c_407_n N_X_c_726_n 3.99786e-19 $X=5.705 $Y=1.22 $X2=0 $Y2=0
cc_365 N_A_313_392#_c_409_n N_X_c_726_n 0.00752662f $X=6.205 $Y=1.22 $X2=0 $Y2=0
cc_366 N_A_313_392#_c_411_n N_X_c_726_n 0.00607717f $X=6.635 $Y=1.22 $X2=0 $Y2=0
cc_367 N_A_313_392#_M1011_g N_X_c_748_n 7.87895e-19 $X=5.695 $Y=2.4 $X2=0 $Y2=0
cc_368 N_A_313_392#_c_407_n N_X_c_748_n 7.96256e-19 $X=5.705 $Y=1.22 $X2=0 $Y2=0
cc_369 N_A_313_392#_M1013_g N_X_c_748_n 0.00532275f $X=6.195 $Y=2.4 $X2=0 $Y2=0
cc_370 N_A_313_392#_c_409_n N_X_c_748_n 0.00454277f $X=6.205 $Y=1.22 $X2=0 $Y2=0
cc_371 N_A_313_392#_c_410_n N_X_c_748_n 0.00855884f $X=6.56 $Y=1.295 $X2=0 $Y2=0
cc_372 N_A_313_392#_c_411_n N_X_c_748_n 0.00599906f $X=6.635 $Y=1.22 $X2=0 $Y2=0
cc_373 N_A_313_392#_M1015_g N_X_c_748_n 0.0193406f $X=6.65 $Y=2.4 $X2=0 $Y2=0
cc_374 N_A_313_392#_c_413_n N_X_c_748_n 0.00657255f $X=6.65 $Y=1.295 $X2=0 $Y2=0
cc_375 N_A_313_392#_c_512_p N_X_c_748_n 0.0239381f $X=5.9 $Y=1.385 $X2=0 $Y2=0
cc_376 N_A_313_392#_c_422_n N_X_c_748_n 0.00790034f $X=6.285 $Y=1.385 $X2=0
+ $Y2=0
cc_377 N_A_313_392#_M1011_g N_X_c_730_n 5.00939e-19 $X=5.695 $Y=2.4 $X2=0 $Y2=0
cc_378 N_A_313_392#_M1013_g N_X_c_730_n 0.015006f $X=6.195 $Y=2.4 $X2=0 $Y2=0
cc_379 N_A_313_392#_M1015_g N_X_c_730_n 0.01346f $X=6.65 $Y=2.4 $X2=0 $Y2=0
cc_380 N_A_313_392#_c_407_n N_X_c_761_n 0.0155444f $X=5.705 $Y=1.22 $X2=0 $Y2=0
cc_381 N_A_313_392#_c_409_n N_X_c_761_n 0.0125913f $X=6.205 $Y=1.22 $X2=0 $Y2=0
cc_382 N_A_313_392#_c_512_p N_X_c_761_n 0.0320524f $X=5.9 $Y=1.385 $X2=0 $Y2=0
cc_383 N_A_313_392#_c_422_n N_X_c_761_n 0.00396053f $X=6.285 $Y=1.385 $X2=0
+ $Y2=0
cc_384 N_A_313_392#_c_409_n N_X_c_765_n 5.42387e-19 $X=6.205 $Y=1.22 $X2=0 $Y2=0
cc_385 N_A_313_392#_c_411_n N_X_c_765_n 0.00256692f $X=6.635 $Y=1.22 $X2=0 $Y2=0
cc_386 N_A_313_392#_M1013_g N_X_c_767_n 0.0018749f $X=6.195 $Y=2.4 $X2=0 $Y2=0
cc_387 N_A_313_392#_M1015_g N_X_c_767_n 0.00695925f $X=6.65 $Y=2.4 $X2=0 $Y2=0
cc_388 N_A_313_392#_c_414_n N_A_27_74#_M1019_d 0.00321419f $X=4.2 $Y=0.34 $X2=0
+ $Y2=0
cc_389 N_A_313_392#_M1005_s N_A_27_74#_c_796_n 0.00213583f $X=2.53 $Y=0.37 $X2=0
+ $Y2=0
cc_390 N_A_313_392#_c_414_n N_A_27_74#_c_796_n 0.00505884f $X=4.2 $Y=0.34 $X2=0
+ $Y2=0
cc_391 N_A_313_392#_c_420_n N_A_27_74#_c_796_n 0.0174411f $X=2.67 $Y=0.34 $X2=0
+ $Y2=0
cc_392 N_A_313_392#_c_414_n N_A_27_74#_c_798_n 0.0210028f $X=4.2 $Y=0.34 $X2=0
+ $Y2=0
cc_393 N_A_313_392#_c_416_n N_VGND_M1017_d 0.00463969f $X=4.915 $Y=1.035 $X2=0
+ $Y2=0
cc_394 N_A_313_392#_c_421_n N_VGND_M1017_d 0.00131647f $X=5 $Y=1.035 $X2=0 $Y2=0
cc_395 N_A_313_392#_c_420_n N_VGND_c_847_n 0.00999258f $X=2.67 $Y=0.34 $X2=0
+ $Y2=0
cc_396 N_A_313_392#_c_403_n N_VGND_c_848_n 0.017509f $X=5.13 $Y=1.22 $X2=0 $Y2=0
cc_397 N_A_313_392#_c_407_n N_VGND_c_848_n 4.29376e-19 $X=5.705 $Y=1.22 $X2=0
+ $Y2=0
cc_398 N_A_313_392#_c_414_n N_VGND_c_848_n 0.0152116f $X=4.2 $Y=0.34 $X2=0 $Y2=0
cc_399 N_A_313_392#_c_415_n N_VGND_c_848_n 0.01598f $X=4.285 $Y=0.95 $X2=0 $Y2=0
cc_400 N_A_313_392#_c_416_n N_VGND_c_848_n 0.0256663f $X=4.915 $Y=1.035 $X2=0
+ $Y2=0
cc_401 N_A_313_392#_c_421_n N_VGND_c_848_n 0.00942489f $X=5 $Y=1.035 $X2=0 $Y2=0
cc_402 N_A_313_392#_c_403_n N_VGND_c_849_n 4.011e-19 $X=5.13 $Y=1.22 $X2=0 $Y2=0
cc_403 N_A_313_392#_c_407_n N_VGND_c_849_n 0.00760292f $X=5.705 $Y=1.22 $X2=0
+ $Y2=0
cc_404 N_A_313_392#_c_409_n N_VGND_c_849_n 0.00328582f $X=6.205 $Y=1.22 $X2=0
+ $Y2=0
cc_405 N_A_313_392#_c_411_n N_VGND_c_851_n 0.0184907f $X=6.635 $Y=1.22 $X2=0
+ $Y2=0
cc_406 N_A_313_392#_c_414_n N_VGND_c_853_n 0.0996519f $X=4.2 $Y=0.34 $X2=0 $Y2=0
cc_407 N_A_313_392#_c_420_n N_VGND_c_853_n 0.0223303f $X=2.67 $Y=0.34 $X2=0
+ $Y2=0
cc_408 N_A_313_392#_c_403_n N_VGND_c_854_n 0.00383152f $X=5.13 $Y=1.22 $X2=0
+ $Y2=0
cc_409 N_A_313_392#_c_407_n N_VGND_c_854_n 0.00383152f $X=5.705 $Y=1.22 $X2=0
+ $Y2=0
cc_410 N_A_313_392#_c_409_n N_VGND_c_855_n 0.00434272f $X=6.205 $Y=1.22 $X2=0
+ $Y2=0
cc_411 N_A_313_392#_c_411_n N_VGND_c_855_n 0.00434272f $X=6.635 $Y=1.22 $X2=0
+ $Y2=0
cc_412 N_A_313_392#_c_403_n N_VGND_c_860_n 0.00758812f $X=5.13 $Y=1.22 $X2=0
+ $Y2=0
cc_413 N_A_313_392#_c_407_n N_VGND_c_860_n 0.0037895f $X=5.705 $Y=1.22 $X2=0
+ $Y2=0
cc_414 N_A_313_392#_c_409_n N_VGND_c_860_n 0.00439256f $X=6.205 $Y=1.22 $X2=0
+ $Y2=0
cc_415 N_A_313_392#_c_411_n N_VGND_c_860_n 0.00823934f $X=6.635 $Y=1.22 $X2=0
+ $Y2=0
cc_416 N_A_313_392#_c_414_n N_VGND_c_860_n 0.0572436f $X=4.2 $Y=0.34 $X2=0 $Y2=0
cc_417 N_A_313_392#_c_420_n N_VGND_c_860_n 0.0124365f $X=2.67 $Y=0.34 $X2=0
+ $Y2=0
cc_418 N_A_313_392#_c_415_n A_835_94# 0.00121649f $X=4.285 $Y=0.95 $X2=-0.19
+ $Y2=-0.245
cc_419 N_A_41_392#_c_582_n N_VPWR_M1000_d 0.00165831f $X=1.085 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_420 N_A_41_392#_c_581_n N_VPWR_c_629_n 0.0233699f $X=0.35 $Y=2.815 $X2=0
+ $Y2=0
cc_421 N_A_41_392#_c_582_n N_VPWR_c_629_n 0.0126919f $X=1.085 $Y=2.035 $X2=0
+ $Y2=0
cc_422 N_A_41_392#_c_585_n N_VPWR_c_629_n 0.0101219f $X=1.415 $Y=2.99 $X2=0
+ $Y2=0
cc_423 N_A_41_392#_c_584_n N_VPWR_c_630_n 0.0121618f $X=1.985 $Y=2.99 $X2=0
+ $Y2=0
cc_424 N_A_41_392#_c_586_n N_VPWR_c_630_n 0.0394061f $X=2.15 $Y=2.455 $X2=0
+ $Y2=0
cc_425 N_A_41_392#_c_584_n N_VPWR_c_639_n 0.0593439f $X=1.985 $Y=2.99 $X2=0
+ $Y2=0
cc_426 N_A_41_392#_c_585_n N_VPWR_c_639_n 0.0234458f $X=1.415 $Y=2.99 $X2=0
+ $Y2=0
cc_427 N_A_41_392#_c_581_n N_VPWR_c_642_n 0.014549f $X=0.35 $Y=2.815 $X2=0 $Y2=0
cc_428 N_A_41_392#_c_581_n N_VPWR_c_628_n 0.0119743f $X=0.35 $Y=2.815 $X2=0
+ $Y2=0
cc_429 N_A_41_392#_c_584_n N_VPWR_c_628_n 0.032751f $X=1.985 $Y=2.99 $X2=0 $Y2=0
cc_430 N_A_41_392#_c_585_n N_VPWR_c_628_n 0.0125551f $X=1.415 $Y=2.99 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_633_n N_X_c_727_n 0.00119078f $X=4.835 $Y=2.955 $X2=0 $Y2=0
cc_432 N_VPWR_c_634_n N_X_c_727_n 0.0353111f $X=5.92 $Y=2.145 $X2=0 $Y2=0
cc_433 N_VPWR_c_640_n N_X_c_727_n 0.0146357f $X=5.755 $Y=3.33 $X2=0 $Y2=0
cc_434 N_VPWR_c_628_n N_X_c_727_n 0.0121141f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_435 N_VPWR_M1011_d N_X_c_728_n 0.00218982f $X=5.785 $Y=1.84 $X2=0 $Y2=0
cc_436 N_VPWR_c_634_n N_X_c_728_n 0.0189268f $X=5.92 $Y=2.145 $X2=0 $Y2=0
cc_437 N_VPWR_c_634_n N_X_c_730_n 0.0353111f $X=5.92 $Y=2.145 $X2=0 $Y2=0
cc_438 N_VPWR_c_636_n N_X_c_730_n 0.0416523f $X=6.92 $Y=1.985 $X2=0 $Y2=0
cc_439 N_VPWR_c_641_n N_X_c_730_n 0.0144772f $X=6.755 $Y=3.33 $X2=0 $Y2=0
cc_440 N_VPWR_c_628_n N_X_c_730_n 0.0118585f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_441 N_VPWR_c_636_n N_X_c_767_n 0.00374248f $X=6.92 $Y=1.985 $X2=0 $Y2=0
cc_442 N_X_c_761_n N_VGND_M1008_s 0.00471803f $X=6.255 $Y=0.93 $X2=0 $Y2=0
cc_443 N_X_c_725_n N_VGND_c_848_n 0.017771f $X=5.42 $Y=0.515 $X2=0 $Y2=0
cc_444 N_X_c_725_n N_VGND_c_849_n 0.011672f $X=5.42 $Y=0.515 $X2=0 $Y2=0
cc_445 N_X_c_726_n N_VGND_c_849_n 0.011672f $X=6.42 $Y=0.515 $X2=0 $Y2=0
cc_446 N_X_c_761_n N_VGND_c_849_n 0.020944f $X=6.255 $Y=0.93 $X2=0 $Y2=0
cc_447 N_X_c_726_n N_VGND_c_851_n 0.0180133f $X=6.42 $Y=0.515 $X2=0 $Y2=0
cc_448 N_X_c_748_n N_VGND_c_851_n 0.00375477f $X=6.42 $Y=1.72 $X2=0 $Y2=0
cc_449 N_X_c_725_n N_VGND_c_854_n 0.0146668f $X=5.42 $Y=0.515 $X2=0 $Y2=0
cc_450 N_X_c_726_n N_VGND_c_855_n 0.0144922f $X=6.42 $Y=0.515 $X2=0 $Y2=0
cc_451 N_X_c_725_n N_VGND_c_860_n 0.0121262f $X=5.42 $Y=0.515 $X2=0 $Y2=0
cc_452 N_X_c_726_n N_VGND_c_860_n 0.0118826f $X=6.42 $Y=0.515 $X2=0 $Y2=0
cc_453 N_X_c_761_n N_VGND_c_860_n 0.0117654f $X=6.255 $Y=0.93 $X2=0 $Y2=0
cc_454 N_A_27_74#_c_793_n N_VGND_M1022_d 0.00354841f $X=1.115 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_455 N_A_27_74#_c_796_n N_VGND_M1014_s 0.00250774f $X=3.005 $Y=0.935 $X2=0
+ $Y2=0
cc_456 N_A_27_74#_c_792_n N_VGND_c_845_n 0.0157994f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_457 N_A_27_74#_c_793_n N_VGND_c_845_n 0.0248957f $X=1.115 $Y=1.005 $X2=0
+ $Y2=0
cc_458 N_A_27_74#_c_795_n N_VGND_c_845_n 0.0157994f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_459 N_A_27_74#_c_795_n N_VGND_c_846_n 0.0144922f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_460 N_A_27_74#_c_795_n N_VGND_c_847_n 0.0105463f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_461 N_A_27_74#_c_796_n N_VGND_c_847_n 0.021281f $X=3.005 $Y=0.935 $X2=0 $Y2=0
cc_462 N_A_27_74#_c_792_n N_VGND_c_852_n 0.0145639f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_463 N_A_27_74#_c_792_n N_VGND_c_860_n 0.0119984f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_464 N_A_27_74#_c_795_n N_VGND_c_860_n 0.0118826f $X=1.28 $Y=0.515 $X2=0 $Y2=0
cc_465 N_A_27_74#_c_796_n N_VGND_c_860_n 0.0275803f $X=3.005 $Y=0.935 $X2=0
+ $Y2=0

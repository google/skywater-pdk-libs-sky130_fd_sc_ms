* File: sky130_fd_sc_ms__or4b_2.pex.spice
* Created: Fri Aug 28 18:09:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__OR4B_2%D_N 1 3 6 8 12
c27 6 0 2.4196e-19 $X=0.51 $Y=0.835
c28 1 0 1.43922e-19 $X=0.505 $Y=1.77
r29 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.515 $X2=0.385 $Y2=1.515
r30 8 12 4.06745 $w=4.23e-07 $l=1.5e-07 $layer=LI1_cond $X=0.337 $Y=1.665
+ $X2=0.337 $Y2=1.515
r31 4 11 38.571 $w=3.25e-07 $l=2.10286e-07 $layer=POLY_cond $X=0.51 $Y=1.35
+ $X2=0.407 $Y2=1.515
r32 4 6 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=0.51 $Y=1.35 $X2=0.51
+ $Y2=0.835
r33 1 11 47.3393 $w=3.25e-07 $l=3.00025e-07 $layer=POLY_cond $X=0.505 $Y=1.77
+ $X2=0.407 $Y2=1.515
r34 1 3 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=0.505 $Y=1.77
+ $X2=0.505 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_2%A_190_48# 1 2 3 12 16 18 22 26 28 30 31 32 35
+ 41 43 47 55 57 59 60 62 63 64
c127 57 0 1.3676e-19 $X=2.34 $Y=1.045
c128 41 0 1.69342e-19 $X=3.54 $Y=0.615
c129 32 0 1.7764e-19 $X=1.745 $Y=1.045
r130 64 65 31.5932 $w=3.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.555 $Y=1.375
+ $X2=1.555 $Y2=1.3
r131 62 63 8.53881 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.05 $Y=2.105
+ $X2=4.05 $Y2=1.94
r132 58 60 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=3.54 $Y=1.115
+ $X2=3.705 $Y2=1.115
r133 58 59 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=3.54 $Y=1.115
+ $X2=3.375 $Y2=1.115
r134 53 67 40.7727 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.555 $Y=1.465
+ $X2=1.555 $Y2=1.63
r135 53 64 14.8382 $w=3.5e-07 $l=9e-08 $layer=POLY_cond $X=1.555 $Y=1.465
+ $X2=1.555 $Y2=1.375
r136 52 55 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.565 $Y=1.465
+ $X2=1.66 $Y2=1.465
r137 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.565
+ $Y=1.465 $X2=1.565 $Y2=1.465
r138 49 63 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.15 $Y=1.27
+ $X2=4.15 $Y2=1.94
r139 45 62 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=4.05 $Y=2.125
+ $X2=4.05 $Y2=2.105
r140 45 47 21.4915 $w=3.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.05 $Y=2.125
+ $X2=4.05 $Y2=2.815
r141 43 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.065 $Y=1.185
+ $X2=4.15 $Y2=1.27
r142 43 60 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.065 $Y=1.185
+ $X2=3.705 $Y2=1.185
r143 39 58 0.331605 $w=3.3e-07 $l=1.55e-07 $layer=LI1_cond $X=3.54 $Y=0.96
+ $X2=3.54 $Y2=1.115
r144 39 41 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.54 $Y=0.96
+ $X2=3.54 $Y2=0.615
r145 38 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=1.045
+ $X2=2.34 $Y2=1.045
r146 38 59 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=2.505 $Y=1.045
+ $X2=3.375 $Y2=1.045
r147 33 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=0.96
+ $X2=2.34 $Y2=1.045
r148 33 35 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.34 $Y=0.96
+ $X2=2.34 $Y2=0.615
r149 31 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.175 $Y=1.045
+ $X2=2.34 $Y2=1.045
r150 31 32 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.175 $Y=1.045
+ $X2=1.745 $Y2=1.045
r151 30 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.66 $Y=1.3
+ $X2=1.66 $Y2=1.465
r152 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.66 $Y=1.13
+ $X2=1.745 $Y2=1.045
r153 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.66 $Y=1.13
+ $X2=1.66 $Y2=1.3
r154 26 67 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.49 $Y=2.4
+ $X2=1.49 $Y2=1.63
r155 22 65 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.455 $Y=0.74
+ $X2=1.455 $Y2=1.3
r156 19 28 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.13 $Y=1.375
+ $X2=1.04 $Y2=1.375
r157 18 64 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.38 $Y=1.375
+ $X2=1.555 $Y2=1.375
r158 18 19 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.38 $Y=1.375
+ $X2=1.13 $Y2=1.375
r159 14 28 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=1.04 $Y=1.45
+ $X2=1.04 $Y2=1.375
r160 14 16 369.274 $w=1.8e-07 $l=9.5e-07 $layer=POLY_cond $X=1.04 $Y=1.45
+ $X2=1.04 $Y2=2.4
r161 10 28 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=1.025 $Y=1.3
+ $X2=1.04 $Y2=1.375
r162 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.025 $Y=1.3
+ $X2=1.025 $Y2=0.74
r163 3 62 400 $w=1.7e-07 $l=3.50071e-07 $layer=licon1_PDIFF $count=1 $X=3.745
+ $Y=1.96 $X2=4.03 $Y2=2.105
r164 3 47 400 $w=1.7e-07 $l=9.87269e-07 $layer=licon1_PDIFF $count=1 $X=3.745
+ $Y=1.96 $X2=4.03 $Y2=2.815
r165 2 41 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=3.355
+ $Y=0.47 $X2=3.54 $Y2=0.615
r166 1 35 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=2.12
+ $Y=0.47 $X2=2.34 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_2%A 3 7 9 10 14 15
c47 3 0 1.08939e-19 $X=2.045 $Y=0.79
r48 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.11 $Y=1.515
+ $X2=2.11 $Y2=1.68
r49 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.11 $Y=1.515
+ $X2=2.11 $Y2=1.35
r50 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.11
+ $Y=1.515 $X2=2.11 $Y2=1.515
r51 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.11 $Y=1.665
+ $X2=2.11 $Y2=2.035
r52 9 15 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.11 $Y=1.665
+ $X2=2.11 $Y2=1.515
r53 7 17 303.194 $w=1.8e-07 $l=7.8e-07 $layer=POLY_cond $X=2.185 $Y=2.46
+ $X2=2.185 $Y2=1.68
r54 3 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.045 $Y=0.79
+ $X2=2.045 $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_2%B 3 7 9 10 14
c39 14 0 1.3676e-19 $X=2.65 $Y=1.635
r40 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.65 $Y=1.635
+ $X2=2.65 $Y2=1.8
r41 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.65 $Y=1.635
+ $X2=2.65 $Y2=1.47
r42 9 10 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=2.65 $Y=1.635 $X2=2.65
+ $Y2=2.035
r43 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.65
+ $Y=1.635 $X2=2.65 $Y2=1.635
r44 7 16 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.635 $Y=0.79
+ $X2=2.635 $Y2=1.47
r45 3 17 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.605 $Y=2.46
+ $X2=2.605 $Y2=1.8
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_2%C 3 7 9 10 11 16
c36 16 0 1.58197e-19 $X=3.19 $Y=1.635
c37 7 0 1.69342e-19 $X=3.28 $Y=0.79
r38 16 19 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.19 $Y=1.635
+ $X2=3.19 $Y2=1.8
r39 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.19 $Y=1.635
+ $X2=3.19 $Y2=1.47
r40 10 11 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.18 $Y=2.035
+ $X2=3.18 $Y2=2.405
r41 9 10 13.1708 $w=3.48e-07 $l=4e-07 $layer=LI1_cond $X=3.18 $Y=1.635 $X2=3.18
+ $Y2=2.035
r42 9 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.19
+ $Y=1.635 $X2=3.19 $Y2=1.635
r43 7 18 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.28 $Y=0.79 $X2=3.28
+ $Y2=1.47
r44 3 19 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.115 $Y=2.46
+ $X2=3.115 $Y2=1.8
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_2%A_27_368# 1 2 9 13 17 19 20 22 23 24 27 28 30
+ 37 38
c98 30 0 1.58197e-19 $X=3.61 $Y=2.69
r99 38 42 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=1.605
+ $X2=3.73 $Y2=1.77
r100 38 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=1.605
+ $X2=3.73 $Y2=1.44
r101 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.73
+ $Y=1.605 $X2=3.73 $Y2=1.605
r102 34 37 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=3.61 $Y=1.605
+ $X2=3.73 $Y2=1.605
r103 32 33 10.1828 $w=6.29e-07 $l=5.25e-07 $layer=LI1_cond $X=0.28 $Y=2.325
+ $X2=0.805 $Y2=2.325
r104 29 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.61 $Y=1.77
+ $X2=3.61 $Y2=1.605
r105 29 30 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.61 $Y=1.77
+ $X2=3.61 $Y2=2.69
r106 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.525 $Y=2.775
+ $X2=3.61 $Y2=2.69
r107 27 28 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=3.525 $Y=2.775
+ $X2=2.465 $Y2=2.775
r108 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.38 $Y=2.69
+ $X2=2.465 $Y2=2.775
r109 25 26 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.38 $Y=2.49 $X2=2.38
+ $Y2=2.69
r110 24 33 9.00042 $w=6.29e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.89 $Y=2.405
+ $X2=0.805 $Y2=2.325
r111 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.295 $Y=2.405
+ $X2=2.38 $Y2=2.49
r112 23 24 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=2.295 $Y=2.405
+ $X2=0.89 $Y2=2.405
r113 22 33 8.62214 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=0.805 $Y=1.95
+ $X2=0.805 $Y2=2.325
r114 21 22 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.805 $Y=1.18
+ $X2=0.805 $Y2=1.95
r115 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.72 $Y=1.095
+ $X2=0.805 $Y2=1.18
r116 19 20 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.72 $Y=1.095
+ $X2=0.46 $Y2=1.095
r117 15 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.295 $Y=1.01
+ $X2=0.46 $Y2=1.095
r118 15 17 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=0.295 $Y=1.01
+ $X2=0.295 $Y2=0.835
r119 13 41 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=3.755 $Y=0.79
+ $X2=3.755 $Y2=1.44
r120 9 42 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=3.655 $Y=2.46
+ $X2=3.655 $Y2=1.77
r121 2 32 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r122 1 17 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.56 $X2=0.295 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_2%VPWR 1 2 11 13 15 25 26 29 32
r44 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r46 22 25 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r47 20 22 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.125 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 19 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r49 19 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 16 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r52 16 18 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33 $X2=1.2
+ $Y2=3.33
r53 15 20 8.04321 $w=1.7e-07 $l=2.88e-07 $layer=LI1_cond $X=1.837 $Y=3.33
+ $X2=2.125 $Y2=3.33
r54 15 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 15 32 10.7127 $w=5.73e-07 $l=5.15e-07 $layer=LI1_cond $X=1.837 $Y=3.33
+ $X2=1.837 $Y2=2.815
r56 15 18 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.55 $Y=3.33 $X2=1.2
+ $Y2=3.33
r57 13 26 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r58 13 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r59 13 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r60 9 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r61 9 11 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.78
r62 2 32 600 $w=1.7e-07 $l=1.0951e-06 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.84 $X2=1.835 $Y2=2.815
r63 1 11 600 $w=1.7e-07 $l=1.04422e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.815 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_2%X 1 2 9 13 14 18
c39 18 0 1.22068e-19 $X=1.245 $Y=1.82
c40 14 0 1.43922e-19 $X=1.2 $Y=2.035
c41 13 0 2.2883e-19 $X=1.232 $Y=1.13
r42 14 18 8.53881 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.245 $Y=1.985
+ $X2=1.245 $Y2=1.82
r43 13 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.145 $Y=1.13
+ $X2=1.145 $Y2=1.82
r44 7 13 8.71323 $w=3.43e-07 $l=1.72e-07 $layer=LI1_cond $X=1.232 $Y=0.958
+ $X2=1.232 $Y2=1.13
r45 7 9 14.798 $w=3.43e-07 $l=4.43e-07 $layer=LI1_cond $X=1.232 $Y=0.958
+ $X2=1.232 $Y2=0.515
r46 2 14 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=1.84 $X2=1.265 $Y2=1.985
r47 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.1 $Y=0.37
+ $X2=1.24 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_2%VGND 1 2 3 4 17 21 25 27 29 31 33 38 43 49 52
+ 55 59
r61 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r62 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r63 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r64 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r65 47 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r66 47 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r67 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r68 44 55 11.5608 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=3.205 $Y=0 $X2=2.945
+ $Y2=0
r69 44 46 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.205 $Y=0 $X2=3.6
+ $Y2=0
r70 43 58 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=3.875 $Y=0 $X2=4.097
+ $Y2=0
r71 43 46 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.875 $Y=0 $X2=3.6
+ $Y2=0
r72 42 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r73 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r74 39 52 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=1.995 $Y=0 $X2=1.785
+ $Y2=0
r75 39 41 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.995 $Y=0 $X2=2.64
+ $Y2=0
r76 38 55 11.5608 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=2.685 $Y=0 $X2=2.945
+ $Y2=0
r77 38 41 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.685 $Y=0 $X2=2.64
+ $Y2=0
r78 37 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r79 37 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r80 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r81 34 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.89 $Y=0 $X2=0.765
+ $Y2=0
r82 34 36 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.89 $Y=0 $X2=1.2
+ $Y2=0
r83 33 52 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=1.575 $Y=0 $X2=1.785
+ $Y2=0
r84 33 36 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.575 $Y=0 $X2=1.2
+ $Y2=0
r85 31 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r86 31 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r87 27 58 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.097 $Y2=0
r88 27 29 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0.69
r89 23 55 2.17428 $w=5.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=0.085
+ $X2=2.945 $Y2=0
r90 23 25 12.1908 $w=5.18e-07 $l=5.3e-07 $layer=LI1_cond $X=2.945 $Y=0.085
+ $X2=2.945 $Y2=0.615
r91 19 52 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=0.085
+ $X2=1.785 $Y2=0
r92 19 21 14.5427 $w=4.18e-07 $l=5.3e-07 $layer=LI1_cond $X=1.785 $Y=0.085
+ $X2=1.785 $Y2=0.615
r93 15 49 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0.085
+ $X2=0.765 $Y2=0
r94 15 17 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=0.765 $Y=0.085
+ $X2=0.765 $Y2=0.595
r95 4 29 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=3.83
+ $Y=0.47 $X2=4.04 $Y2=0.69
r96 3 25 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=2.71
+ $Y=0.47 $X2=2.945 $Y2=0.615
r97 2 21 182 $w=1.7e-07 $l=3.57071e-07 $layer=licon1_NDIFF $count=1 $X=1.53
+ $Y=0.37 $X2=1.785 $Y2=0.615
r98 1 17 182 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_NDIFF $count=1 $X=0.585
+ $Y=0.56 $X2=0.805 $Y2=0.595
.ends


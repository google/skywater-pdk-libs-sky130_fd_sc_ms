* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or4b_1 A B C D_N VGND VNB VPB VPWR X
X0 VPWR a_228_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 a_27_74# D_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X2 VGND B a_228_74# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X3 a_228_74# a_27_74# a_359_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X4 a_527_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X5 VGND a_27_74# a_228_74# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X6 a_359_368# C a_443_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X7 a_228_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X8 VGND a_228_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_443_368# B a_527_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X10 a_228_74# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X11 a_27_74# D_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
.ends

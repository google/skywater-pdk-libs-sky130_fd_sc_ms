* NGSPICE file created from sky130_fd_sc_ms__einvn_4.ext - technology: sky130A

.subckt sky130_fd_sc_ms__einvn_4 A TE_B VGND VNB VPB VPWR Z
M1000 VPWR TE_B a_241_368# VPB pshort w=1.12e+06u l=180000u
+  ad=9.744e+11p pd=8.46e+06u as=1.5344e+12p ps=1.394e+07u
M1001 a_281_74# A Z VNB nlowvt w=740000u l=150000u
+  ad=1.0508e+12p pd=1.024e+07u as=4.144e+11p ps=4.08e+06u
M1002 a_241_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_281_74# a_114_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=6.253e+11p ps=6.13e+06u
M1004 VPWR TE_B a_241_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_241_368# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_114_74# a_281_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_281_74# A Z VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Z A a_241_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1009 a_241_368# A Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Z A a_241_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_241_368# A Z VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Z A a_281_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_281_74# a_114_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_114_74# TE_B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1015 a_114_74# TE_B VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1016 Z A a_281_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_114_74# a_281_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__sdfxtp_1.pex.spice
* Created: Wed Sep  2 12:31:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SDFXTP_1%A_35_74# 1 2 9 13 16 18 21 23 27 28 33 40
+ 41
c95 41 0 1.8681e-19 $X=0.825 $Y=1.825
c96 40 0 1.63729e-19 $X=0.66 $Y=1.69
r97 39 41 10.1561 $w=5.98e-07 $l=1.65e-07 $layer=LI1_cond $X=0.66 $Y=1.825
+ $X2=0.825 $Y2=1.825
r98 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.66
+ $Y=1.69 $X2=0.66 $Y2=1.69
r99 37 39 6.77778 $w=5.98e-07 $l=3.4e-07 $layer=LI1_cond $X=0.32 $Y=1.825
+ $X2=0.66 $Y2=1.825
r100 35 37 2.9902 $w=5.98e-07 $l=1.5e-07 $layer=LI1_cond $X=0.17 $Y=1.825
+ $X2=0.32 $Y2=1.825
r101 30 33 3.97394 $w=4.33e-07 $l=1.5e-07 $layer=LI1_cond $X=0.17 $Y=0.567
+ $X2=0.32 $Y2=0.567
r102 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.03
+ $Y=1.635 $X2=2.03 $Y2=1.635
r103 25 27 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=2.03 $Y=1.955
+ $X2=2.03 $Y2=1.635
r104 23 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.865 $Y=2.04
+ $X2=2.03 $Y2=1.955
r105 23 41 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=1.865 $Y=2.04
+ $X2=0.825 $Y2=2.04
r106 19 37 2.16985 $w=4.7e-07 $l=3e-07 $layer=LI1_cond $X=0.32 $Y=2.125 $X2=0.32
+ $Y2=1.825
r107 19 21 8.65248 $w=4.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.32 $Y=2.125
+ $X2=0.32 $Y2=2.465
r108 18 35 8.31678 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=0.17 $Y=1.525 $X2=0.17
+ $Y2=1.825
r109 17 30 6.29128 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.17 $Y=0.785
+ $X2=0.17 $Y2=0.567
r110 17 18 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.17 $Y=0.785
+ $X2=0.17 $Y2=1.525
r111 15 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.03 $Y=1.975
+ $X2=2.03 $Y2=1.635
r112 15 16 37.308 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.03 $Y=1.975
+ $X2=2.03 $Y2=2.14
r113 13 16 194.355 $w=1.8e-07 $l=5e-07 $layer=POLY_cond $X=1.985 $Y=2.64
+ $X2=1.985 $Y2=2.14
r114 7 40 74.7592 $w=2.45e-07 $l=4.55082e-07 $layer=POLY_cond $X=1.04 $Y=1.525
+ $X2=0.66 $Y2=1.69
r115 7 9 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=1.04 $Y=1.525
+ $X2=1.04 $Y2=0.58
r116 2 21 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.245
+ $Y=2.32 $X2=0.39 $Y2=2.465
r117 1 33 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.37 $X2=0.32 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_1%SCE 2 3 4 5 6 9 11 13 14 16 18 21 22 26 30
+ 31 33 40 43 45
r87 33 45 3.36024 $w=4.73e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.047
+ $X2=1.315 $Y2=1.047
r88 33 43 4.02225 $w=4.73e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.047
+ $X2=1.085 $Y2=1.047
r89 31 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.085 $Y=1.065
+ $X2=2.085 $Y2=0.9
r90 30 45 23.0489 $w=3.83e-07 $l=7.7e-07 $layer=LI1_cond $X=2.085 $Y=1.092
+ $X2=1.315 $Y2=1.092
r91 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.085
+ $Y=1.065 $X2=2.085 $Y2=1.065
r92 26 37 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.59 $Y=1.12 $X2=0.59
+ $Y2=1.21
r93 26 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.12
+ $X2=0.59 $Y2=0.955
r94 25 43 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.59 $Y=1.12
+ $X2=1.085 $Y2=1.12
r95 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.12 $X2=0.59 $Y2=1.12
r96 21 40 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.175 $Y=0.58
+ $X2=2.175 $Y2=0.9
r97 16 18 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.115 $Y=2.245
+ $X2=1.115 $Y2=2.64
r98 15 22 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.705 $Y=2.17
+ $X2=0.615 $Y2=2.17
r99 14 16 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.025 $Y=2.17
+ $X2=1.115 $Y2=2.245
r100 14 15 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.025 $Y=2.17
+ $X2=0.705 $Y2=2.17
r101 11 22 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=0.615 $Y=2.245
+ $X2=0.615 $Y2=2.17
r102 11 13 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.615 $Y=2.245
+ $X2=0.615 $Y2=2.64
r103 9 36 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=0.535 $Y=0.58
+ $X2=0.535 $Y2=0.955
r104 5 22 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.525 $Y=2.17
+ $X2=0.615 $Y2=2.17
r105 5 6 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.525 $Y=2.17
+ $X2=0.255 $Y2=2.17
r106 3 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.425 $Y=1.21
+ $X2=0.59 $Y2=1.21
r107 3 4 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.425 $Y=1.21
+ $X2=0.255 $Y2=1.21
r108 2 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.18 $Y=2.095
+ $X2=0.255 $Y2=2.17
r109 1 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.18 $Y=1.285
+ $X2=0.255 $Y2=1.21
r110 1 2 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.18 $Y=1.285 $X2=0.18
+ $Y2=2.095
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_1%D 3 7 9 12 13
c39 12 0 1.8681e-19 $X=1.49 $Y=1.62
r40 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.49 $Y=1.62
+ $X2=1.49 $Y2=1.785
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.49 $Y=1.62
+ $X2=1.49 $Y2=1.455
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.49
+ $Y=1.62 $X2=1.49 $Y2=1.62
r43 9 13 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.2 $Y=1.62 $X2=1.49
+ $Y2=1.62
r44 7 15 332.347 $w=1.8e-07 $l=8.55e-07 $layer=POLY_cond $X=1.535 $Y=2.64
+ $X2=1.535 $Y2=1.785
r45 3 14 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=1.43 $Y=0.58 $X2=1.43
+ $Y2=1.455
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_1%SCD 3 7 11 12 13 16
c46 7 0 7.17504e-20 $X=2.565 $Y=0.58
r47 13 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.57
+ $Y=1.635 $X2=2.57 $Y2=1.635
r48 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.57 $Y=1.975
+ $X2=2.57 $Y2=1.635
r49 11 12 37.308 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.975
+ $X2=2.57 $Y2=2.14
r50 10 16 37.7798 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.47
+ $X2=2.57 $Y2=1.635
r51 7 10 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=2.565 $Y=0.58
+ $X2=2.565 $Y2=1.47
r52 3 12 194.355 $w=1.8e-07 $l=5e-07 $layer=POLY_cond $X=2.525 $Y=2.64 $X2=2.525
+ $Y2=2.14
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_1%CLK 1 3 6 8 11
c43 8 0 7.17504e-20 $X=3.6 $Y=1.295
r44 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.415
+ $Y=1.385 $X2=3.415 $Y2=1.385
r45 11 13 30.4421 $w=2.85e-07 $l=1.8e-07 $layer=POLY_cond $X=3.235 $Y=1.385
+ $X2=3.415 $Y2=1.385
r46 8 14 5.76222 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.6 $Y=1.365
+ $X2=3.415 $Y2=1.365
r47 4 11 13.5351 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.235 $Y=1.55
+ $X2=3.235 $Y2=1.385
r48 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.235 $Y=1.55
+ $X2=3.235 $Y2=2.4
r49 1 11 27.0596 $w=2.85e-07 $l=2.31571e-07 $layer=POLY_cond $X=3.075 $Y=1.22
+ $X2=3.235 $Y2=1.385
r50 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.075 $Y=1.22 $X2=3.075
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_1%A_828_74# 1 2 9 11 13 16 19 21 24 26 27 29
+ 30 33 36 37 39 42 43 44 47 51 52 57 58 60 61 63 64 65 78
c197 64 0 7.65965e-20 $X=7.57 $Y=1.195
c198 58 0 7.022e-20 $X=5.12 $Y=2.215
c199 57 0 4.72498e-21 $X=5.12 $Y=2.215
c200 47 0 7.308e-20 $X=8.07 $Y=1.275
c201 33 0 1.68607e-19 $X=5.82 $Y=0.69
c202 19 0 1.46857e-19 $X=8.365 $Y=2.75
r203 64 78 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.57 $Y=1.195
+ $X2=7.57 $Y2=1.03
r204 63 66 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.65 $Y=1.195 $X2=7.65
+ $Y2=1.275
r205 63 65 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.65 $Y=1.195
+ $X2=7.65 $Y2=1.03
r206 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.57
+ $Y=1.195 $X2=7.57 $Y2=1.195
r207 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.12
+ $Y=2.215 $X2=5.12 $Y2=2.215
r208 55 57 17.8075 $w=3.22e-07 $l=4.7e-07 $layer=LI1_cond $X=4.65 $Y=2.1
+ $X2=5.12 $Y2=2.1
r209 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.47
+ $Y=1.57 $X2=8.47 $Y2=1.57
r210 49 51 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=8.43 $Y=1.49 $X2=8.43
+ $Y2=1.57
r211 48 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.815 $Y=1.275
+ $X2=7.65 $Y2=1.275
r212 47 49 20.9966 $w=2.15e-07 $l=3.91152e-07 $layer=LI1_cond $X=8.07 $Y=1.275
+ $X2=8.43 $Y2=1.34
r213 47 48 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.07 $Y=1.275
+ $X2=7.815 $Y2=1.275
r214 45 65 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=7.73 $Y=0.425
+ $X2=7.73 $Y2=1.03
r215 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.645 $Y=0.34
+ $X2=7.73 $Y2=0.425
r216 43 44 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.645 $Y=0.34
+ $X2=6.975 $Y2=0.34
r217 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.89 $Y=0.425
+ $X2=6.975 $Y2=0.34
r218 41 42 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.89 $Y=0.425
+ $X2=6.89 $Y2=0.69
r219 40 61 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.985 $Y=0.775
+ $X2=5.86 $Y2=0.775
r220 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.805 $Y=0.775
+ $X2=6.89 $Y2=0.69
r221 39 40 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=6.805 $Y=0.775
+ $X2=5.985 $Y2=0.775
r222 37 73 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.82 $Y=1.195
+ $X2=5.695 $Y2=1.195
r223 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.82
+ $Y=1.195 $X2=5.82 $Y2=1.195
r224 34 61 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.86 $Y=0.86 $X2=5.86
+ $Y2=0.775
r225 34 36 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.86 $Y=0.86
+ $X2=5.86 $Y2=1.195
r226 33 61 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=5.82 $Y=0.69
+ $X2=5.86 $Y2=0.775
r227 32 33 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.82 $Y=0.425
+ $X2=5.82 $Y2=0.69
r228 31 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.225 $Y=0.34
+ $X2=5.14 $Y2=0.34
r229 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.735 $Y=0.34
+ $X2=5.82 $Y2=0.425
r230 30 31 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.735 $Y=0.34
+ $X2=5.225 $Y2=0.34
r231 29 57 0.757764 $w=3.22e-07 $l=2e-08 $layer=LI1_cond $X=5.14 $Y=2.1 $X2=5.12
+ $Y2=2.1
r232 28 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.14 $Y=0.425
+ $X2=5.14 $Y2=0.34
r233 28 29 106.016 $w=1.68e-07 $l=1.625e-06 $layer=LI1_cond $X=5.14 $Y=0.425
+ $X2=5.14 $Y2=2.05
r234 26 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.055 $Y=0.34
+ $X2=5.14 $Y2=0.34
r235 26 27 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.055 $Y=0.34
+ $X2=4.445 $Y2=0.34
r236 22 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.32 $Y=0.425
+ $X2=4.445 $Y2=0.34
r237 22 24 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.32 $Y=0.425
+ $X2=4.32 $Y2=0.515
r238 21 52 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.47 $Y=1.91
+ $X2=8.47 $Y2=1.57
r239 17 21 44.3718 $w=2.77e-07 $l=3.02985e-07 $layer=POLY_cond $X=8.365 $Y=2.165
+ $X2=8.47 $Y2=1.91
r240 17 19 227.395 $w=1.8e-07 $l=5.85e-07 $layer=POLY_cond $X=8.365 $Y=2.165
+ $X2=8.365 $Y2=2.75
r241 16 78 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=7.525 $Y=0.645
+ $X2=7.525 $Y2=1.03
r242 11 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.695 $Y=1.03
+ $X2=5.695 $Y2=1.195
r243 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.695 $Y=1.03
+ $X2=5.695 $Y2=0.71
r244 7 58 59.7756 $w=2.54e-07 $l=3.88844e-07 $layer=POLY_cond $X=5.435 $Y=2.38
+ $X2=5.12 $Y2=2.215
r245 7 9 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=5.435 $Y=2.38
+ $X2=5.435 $Y2=2.75
r246 2 55 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=4.515
+ $Y=1.84 $X2=4.65 $Y2=2.02
r247 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.14
+ $Y=0.37 $X2=4.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_1%A_630_74# 1 2 9 11 15 17 21 23 29 33 36 37
+ 38 39 41 42 43 48 50 54 55 58 61 62 64 65 66 68 69 72 74 79 80 87
c212 68 0 1.8193e-19 $X=7.63 $Y=2.52
c213 66 0 1.11961e-19 $X=6.215 $Y=2.605
c214 43 0 1.89404e-19 $X=5.015 $Y=1.555
c215 37 0 1.41929e-19 $X=8.29 $Y=1.09
c216 29 0 8.19904e-20 $X=5.935 $Y=2.75
c217 21 0 1.68607e-19 $X=5.015 $Y=0.71
r218 80 88 13.7452 $w=2.63e-07 $l=7.5e-08 $layer=POLY_cond $X=7.735 $Y=1.765
+ $X2=7.66 $Y2=1.765
r219 79 80 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.735
+ $Y=1.765 $X2=7.735 $Y2=1.765
r220 76 79 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=7.63 $Y=1.765
+ $X2=7.735 $Y2=1.765
r221 72 87 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.9 $Y=2.035
+ $X2=5.9 $Y2=2.2
r222 71 74 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=5.9 $Y=2.035
+ $X2=6.13 $Y2=2.035
r223 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.9
+ $Y=2.035 $X2=5.9 $Y2=2.035
r224 67 76 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.63 $Y=1.93
+ $X2=7.63 $Y2=1.765
r225 67 68 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.63 $Y=1.93
+ $X2=7.63 $Y2=2.52
r226 65 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.545 $Y=2.605
+ $X2=7.63 $Y2=2.52
r227 65 66 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=7.545 $Y=2.605
+ $X2=6.215 $Y2=2.605
r228 64 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.13 $Y=2.52
+ $X2=6.215 $Y2=2.605
r229 63 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.13 $Y=2.2
+ $X2=6.13 $Y2=2.035
r230 63 64 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.13 $Y=2.2 $X2=6.13
+ $Y2=2.52
r231 62 84 14.8382 $w=3.5e-07 $l=9e-08 $layer=POLY_cond $X=3.965 $Y=1.465
+ $X2=3.965 $Y2=1.555
r232 62 83 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.965 $Y=1.465
+ $X2=3.965 $Y2=1.3
r233 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.955
+ $Y=1.465 $X2=3.955 $Y2=1.465
r234 59 61 19.6864 $w=1.98e-07 $l=3.55e-07 $layer=LI1_cond $X=3.955 $Y=1.82
+ $X2=3.955 $Y2=1.465
r235 58 69 5.8268 $w=1.98e-07 $l=1e-07 $layer=LI1_cond $X=3.955 $Y=1.4 $X2=3.955
+ $Y2=1.3
r236 58 61 3.60455 $w=1.98e-07 $l=6.5e-08 $layer=LI1_cond $X=3.955 $Y=1.4
+ $X2=3.955 $Y2=1.465
r237 56 69 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.94 $Y=0.96
+ $X2=3.94 $Y2=1.3
r238 54 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.855 $Y=0.875
+ $X2=3.94 $Y2=0.96
r239 54 55 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.855 $Y=0.875
+ $X2=3.455 $Y2=0.875
r240 50 59 7.29955 $w=3.2e-07 $l=2.03961e-07 $layer=LI1_cond $X=3.855 $Y=1.98
+ $X2=3.955 $Y2=1.82
r241 50 52 14.2255 $w=3.18e-07 $l=3.95e-07 $layer=LI1_cond $X=3.855 $Y=1.98
+ $X2=3.46 $Y2=1.98
r242 46 55 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.29 $Y=0.79
+ $X2=3.455 $Y2=0.875
r243 46 48 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.29 $Y=0.79
+ $X2=3.29 $Y2=0.515
r244 43 44 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.015 $Y=1.555
+ $X2=5.015 $Y2=1.765
r245 39 41 98.0067 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=8.365 $Y=1.015
+ $X2=8.365 $Y2=0.71
r246 37 39 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.29 $Y=1.09
+ $X2=8.365 $Y2=1.015
r247 37 38 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=8.29 $Y=1.09
+ $X2=8.095 $Y2=1.09
r248 36 80 52.2319 $w=2.63e-07 $l=3.5812e-07 $layer=POLY_cond $X=8.02 $Y=1.6
+ $X2=7.735 $Y2=1.765
r249 35 38 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.02 $Y=1.165
+ $X2=8.095 $Y2=1.09
r250 35 36 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.02 $Y=1.165
+ $X2=8.02 $Y2=1.6
r251 31 88 11.6845 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.66 $Y=1.93
+ $X2=7.66 $Y2=1.765
r252 31 33 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=7.66 $Y=1.93
+ $X2=7.66 $Y2=2.54
r253 29 87 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=5.935 $Y=2.75
+ $X2=5.935 $Y2=2.2
r254 25 72 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=5.9 $Y=1.84
+ $X2=5.9 $Y2=2.035
r255 24 44 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.09 $Y=1.765
+ $X2=5.015 $Y2=1.765
r256 23 25 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.735 $Y=1.765
+ $X2=5.9 $Y2=1.84
r257 23 24 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=5.735 $Y=1.765
+ $X2=5.09 $Y2=1.765
r258 19 43 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.015 $Y=1.48
+ $X2=5.015 $Y2=1.555
r259 19 21 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=5.015 $Y=1.48
+ $X2=5.015 $Y2=0.71
r260 18 42 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.515 $Y=1.555
+ $X2=4.425 $Y2=1.555
r261 17 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.94 $Y=1.555
+ $X2=5.015 $Y2=1.555
r262 17 18 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=4.94 $Y=1.555
+ $X2=4.515 $Y2=1.555
r263 13 42 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.425 $Y=1.63
+ $X2=4.425 $Y2=1.555
r264 13 15 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.425 $Y=1.63
+ $X2=4.425 $Y2=2.4
r265 12 84 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.14 $Y=1.555
+ $X2=3.965 $Y2=1.555
r266 11 42 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.335 $Y=1.555
+ $X2=4.425 $Y2=1.555
r267 11 12 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=4.335 $Y=1.555
+ $X2=4.14 $Y2=1.555
r268 9 83 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.065 $Y=0.74
+ $X2=4.065 $Y2=1.3
r269 2 52 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=3.325
+ $Y=1.84 $X2=3.46 $Y2=2.02
r270 1 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.15
+ $Y=0.37 $X2=3.29 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_1%A_1239_74# 1 2 9 10 12 16 17 20 23 27 28 31
+ 34 36
c77 12 0 1.67177e-19 $X=6.335 $Y=2.75
r78 31 33 8.8114 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=7.31 $Y=0.685
+ $X2=7.31 $Y2=0.86
r79 27 28 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=7.195 $Y=2.265
+ $X2=7.195 $Y2=2.1
r80 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.23 $Y=1.36
+ $X2=7.23 $Y2=1.195
r81 24 28 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=7.23 $Y=1.36
+ $X2=7.23 $Y2=2.1
r82 23 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.23 $Y=1.03
+ $X2=7.23 $Y2=1.195
r83 23 33 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.23 $Y=1.03
+ $X2=7.23 $Y2=0.86
r84 20 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.36 $Y=1.195
+ $X2=6.36 $Y2=1.36
r85 20 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.36 $Y=1.195
+ $X2=6.36 $Y2=1.03
r86 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.36
+ $Y=1.195 $X2=6.36 $Y2=1.195
r87 17 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.145 $Y=1.195
+ $X2=7.23 $Y2=1.195
r88 17 19 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=7.145 $Y=1.195
+ $X2=6.36 $Y2=1.195
r89 16 37 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=6.35 $Y=2.315
+ $X2=6.35 $Y2=1.36
r90 10 16 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.335 $Y=2.405
+ $X2=6.335 $Y2=2.315
r91 10 12 134.105 $w=1.8e-07 $l=3.45e-07 $layer=POLY_cond $X=6.335 $Y=2.405
+ $X2=6.335 $Y2=2.75
r92 9 36 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.27 $Y=0.71 $X2=6.27
+ $Y2=1.03
r93 2 27 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=7.045
+ $Y=2.12 $X2=7.195 $Y2=2.265
r94 1 31 182 $w=1.7e-07 $l=3.80657e-07 $layer=licon1_NDIFF $count=1 $X=7.165
+ $Y=0.37 $X2=7.31 $Y2=0.685
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_1%A_1018_100# 1 2 9 13 17 23 25 27 28 29 30
+ 39
c90 29 0 1.67177e-19 $X=5.635 $Y=2.54
c91 27 0 1.97671e-19 $X=5.48 $Y=1.615
c92 9 0 3.50729e-20 $X=6.955 $Y=2.54
r93 38 39 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6.955 $Y=1.765
+ $X2=7.09 $Y2=1.765
r94 34 38 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=6.81 $Y=1.765
+ $X2=6.955 $Y2=1.765
r95 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.81
+ $Y=1.765 $X2=6.81 $Y2=1.765
r96 30 33 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=6.81 $Y=1.615
+ $X2=6.81 $Y2=1.765
r97 28 29 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.635 $Y=2.37
+ $X2=5.635 $Y2=2.54
r98 26 27 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=1.615
+ $X2=5.48 $Y2=1.615
r99 25 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.645 $Y=1.615
+ $X2=6.81 $Y2=1.615
r100 25 26 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=6.645 $Y=1.615
+ $X2=5.565 $Y2=1.615
r101 23 29 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=5.71 $Y=2.75
+ $X2=5.71 $Y2=2.54
r102 19 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=1.7 $X2=5.48
+ $Y2=1.615
r103 19 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.48 $Y=1.7
+ $X2=5.48 $Y2=2.37
r104 15 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=1.53
+ $X2=5.48 $Y2=1.615
r105 15 17 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=5.48 $Y=1.53
+ $X2=5.48 $Y2=0.765
r106 11 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.09 $Y=1.6
+ $X2=7.09 $Y2=1.765
r107 11 13 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=7.09 $Y=1.6
+ $X2=7.09 $Y2=0.645
r108 7 38 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.955 $Y=1.93
+ $X2=6.955 $Y2=1.765
r109 7 9 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=6.955 $Y=1.93
+ $X2=6.955 $Y2=2.54
r110 2 23 600 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_PDIFF $count=1 $X=5.525
+ $Y=2.54 $X2=5.71 $Y2=2.75
r111 1 17 182 $w=1.7e-07 $l=5.05421e-07 $layer=licon1_NDIFF $count=1 $X=5.09
+ $Y=0.5 $X2=5.48 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_1%A_1736_74# 1 2 7 9 10 12 14 17 21 25 27 28
+ 29 38 40 43 44 52
c86 44 0 1.61732e-19 $X=9.762 $Y=2.1
c87 29 0 4.59464e-20 $X=9.65 $Y=1.195
c88 27 0 4.09155e-20 $X=10.45 $Y=1.485
c89 14 0 7.308e-20 $X=8.95 $Y=2.315
r90 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.08
+ $Y=1.485 $X2=10.08 $Y2=1.485
r91 45 47 8.48441 $w=4.17e-07 $l=2.9e-07 $layer=LI1_cond $X=9.947 $Y=1.195
+ $X2=9.947 $Y2=1.485
r92 43 44 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=9.762 $Y=2.265
+ $X2=9.762 $Y2=2.1
r93 40 47 9.23389 $w=4.17e-07 $l=2.07918e-07 $layer=LI1_cond $X=9.85 $Y=1.65
+ $X2=9.947 $Y2=1.485
r94 40 44 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=9.85 $Y=1.65
+ $X2=9.85 $Y2=2.1
r95 36 45 5.39268 $w=4.17e-07 $l=2.21371e-07 $layer=LI1_cond $X=9.815 $Y=1.03
+ $X2=9.947 $Y2=1.195
r96 36 38 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=9.815 $Y=1.03
+ $X2=9.815 $Y2=0.645
r97 32 52 33.8246 $w=2.85e-07 $l=2e-07 $layer=POLY_cond $X=9.15 $Y=1.187
+ $X2=8.95 $Y2=1.187
r98 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.15
+ $Y=1.195 $X2=9.15 $Y2=1.195
r99 29 45 2.11011 $w=3.3e-07 $l=2.97e-07 $layer=LI1_cond $X=9.65 $Y=1.195
+ $X2=9.947 $Y2=1.195
r100 29 31 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=9.65 $Y=1.195
+ $X2=9.15 $Y2=1.195
r101 27 48 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=10.45 $Y=1.485
+ $X2=10.08 $Y2=1.485
r102 27 28 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=10.45 $Y=1.485
+ $X2=10.54 $Y2=1.485
r103 19 28 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=10.555 $Y=1.32
+ $X2=10.54 $Y2=1.485
r104 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=10.555 $Y=1.32
+ $X2=10.555 $Y2=0.76
r105 15 28 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=10.54 $Y=1.65
+ $X2=10.54 $Y2=1.485
r106 15 17 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=10.54 $Y=1.65
+ $X2=10.54 $Y2=2.4
r107 14 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.95 $Y=2.315
+ $X2=8.95 $Y2=2.39
r108 13 52 17.7656 $w=1.5e-07 $l=1.73e-07 $layer=POLY_cond $X=8.95 $Y=1.36
+ $X2=8.95 $Y2=1.187
r109 13 14 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=8.95 $Y=1.36
+ $X2=8.95 $Y2=2.315
r110 10 25 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.785 $Y=2.39
+ $X2=8.95 $Y2=2.39
r111 10 12 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=8.785 $Y=2.465
+ $X2=8.785 $Y2=2.75
r112 7 52 32.9789 $w=2.85e-07 $l=2.67516e-07 $layer=POLY_cond $X=8.755 $Y=1.015
+ $X2=8.95 $Y2=1.187
r113 7 9 98.0067 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=8.755 $Y=1.015
+ $X2=8.755 $Y2=0.71
r114 2 43 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=9.62
+ $Y=2.12 $X2=9.755 $Y2=2.265
r115 1 38 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=9.675
+ $Y=0.37 $X2=9.815 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_1%A_1520_74# 1 2 9 13 15 17 19 22 24 27 28 33
+ 35
c89 33 0 7.65965e-20 $X=8.15 $Y=0.71
c90 27 0 4.09155e-20 $X=9.43 $Y=1.765
c91 22 0 9.5983e-20 $X=8.81 $Y=1.6
r92 28 38 40.172 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=9.47 $Y=1.765
+ $X2=9.47 $Y2=1.93
r93 28 37 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=9.47 $Y=1.765
+ $X2=9.47 $Y2=1.6
r94 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.43
+ $Y=1.765 $X2=9.43 $Y2=1.765
r95 25 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.895 $Y=1.765
+ $X2=8.81 $Y2=1.765
r96 25 27 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=8.895 $Y=1.765
+ $X2=9.43 $Y2=1.765
r97 23 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.81 $Y=1.93
+ $X2=8.81 $Y2=1.765
r98 23 24 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.81 $Y=1.93
+ $X2=8.81 $Y2=2.245
r99 22 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.81 $Y=1.6 $X2=8.81
+ $Y2=1.765
r100 21 33 25.6433 $w=3.14e-07 $l=8.1037e-07 $layer=LI1_cond $X=8.81 $Y=1.15
+ $X2=8.15 $Y2=0.815
r101 21 22 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=8.81 $Y=1.15
+ $X2=8.81 $Y2=1.6
r102 20 31 3.97288 $w=1.7e-07 $l=1.57321e-07 $layer=LI1_cond $X=8.135 $Y=2.33
+ $X2=8.01 $Y2=2.257
r103 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.725 $Y=2.33
+ $X2=8.81 $Y2=2.245
r104 19 20 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.725 $Y=2.33
+ $X2=8.135 $Y2=2.33
r105 15 31 3.17028 $w=2.5e-07 $l=1.58e-07 $layer=LI1_cond $X=8.01 $Y=2.415
+ $X2=8.01 $Y2=2.257
r106 15 17 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=8.01 $Y=2.415
+ $X2=8.01 $Y2=2.815
r107 13 37 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=9.6 $Y=0.645
+ $X2=9.6 $Y2=1.6
r108 9 38 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=9.53 $Y=2.54
+ $X2=9.53 $Y2=1.93
r109 2 31 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=7.75
+ $Y=2.12 $X2=7.97 $Y2=2.265
r110 2 17 600 $w=1.7e-07 $l=7.97449e-07 $layer=licon1_PDIFF $count=1 $X=7.75
+ $Y=2.12 $X2=7.97 $Y2=2.815
r111 1 33 182 $w=1.7e-07 $l=6.99643e-07 $layer=licon1_NDIFF $count=1 $X=7.6
+ $Y=0.37 $X2=8.15 $Y2=0.71
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_1%VPWR 1 2 3 4 5 6 21 25 29 33 37 41 46 47 49
+ 50 52 53 54 66 70 75 85 86 89 92 95
c120 21 0 1.63729e-19 $X=0.89 $Y=2.465
r121 95 96 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r122 92 93 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r123 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r124 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r125 83 86 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.8 $Y2=3.33
r126 83 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=8.88 $Y2=3.33
r127 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r128 80 95 12.2593 $w=1.7e-07 $l=2.88e-07 $layer=LI1_cond $X=9.42 $Y=3.33
+ $X2=9.132 $Y2=3.33
r129 80 82 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=9.42 $Y=3.33
+ $X2=9.84 $Y2=3.33
r130 79 96 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.88 $Y2=3.33
r131 79 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r132 78 79 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r133 76 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.81 $Y=3.33
+ $X2=6.645 $Y2=3.33
r134 76 78 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=6.81 $Y=3.33
+ $X2=6.96 $Y2=3.33
r135 75 95 12.2593 $w=1.7e-07 $l=2.87e-07 $layer=LI1_cond $X=8.845 $Y=3.33
+ $X2=9.132 $Y2=3.33
r136 75 78 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=8.845 $Y=3.33
+ $X2=6.96 $Y2=3.33
r137 74 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r138 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r139 71 89 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=4.365 $Y=3.33
+ $X2=4.11 $Y2=3.33
r140 71 73 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=4.365 $Y=3.33
+ $X2=4.56 $Y2=3.33
r141 70 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=6.645 $Y2=3.33
r142 70 73 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=4.56 $Y2=3.33
r143 69 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r144 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r145 66 89 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=4.11 $Y2=3.33
r146 66 68 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=3.6 $Y2=3.33
r147 65 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r148 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r149 62 65 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r150 61 64 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r151 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r152 58 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r153 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r154 54 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r155 54 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r156 52 82 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.15 $Y=3.33
+ $X2=9.84 $Y2=3.33
r157 52 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.15 $Y=3.33
+ $X2=10.275 $Y2=3.33
r158 51 85 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=10.4 $Y=3.33 $X2=10.8
+ $Y2=3.33
r159 51 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.4 $Y=3.33
+ $X2=10.275 $Y2=3.33
r160 49 64 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.67 $Y=3.33 $X2=2.64
+ $Y2=3.33
r161 49 50 11.3601 $w=1.7e-07 $l=2.52e-07 $layer=LI1_cond $X=2.67 $Y=3.33
+ $X2=2.922 $Y2=3.33
r162 48 68 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.175 $Y=3.33
+ $X2=3.6 $Y2=3.33
r163 48 50 11.3601 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=3.175 $Y=3.33
+ $X2=2.922 $Y2=3.33
r164 46 57 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.72 $Y2=3.33
r165 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.89 $Y2=3.33
r166 45 61 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.2 $Y2=3.33
r167 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.89 $Y2=3.33
r168 41 44 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=10.275 $Y=1.985
+ $X2=10.275 $Y2=2.815
r169 39 53 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.275 $Y=3.245
+ $X2=10.275 $Y2=3.33
r170 39 44 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.275 $Y=3.245
+ $X2=10.275 $Y2=2.815
r171 35 95 2.42056 $w=5.75e-07 $l=8.5e-08 $layer=LI1_cond $X=9.132 $Y=3.245
+ $X2=9.132 $Y2=3.33
r172 35 37 8.94459 $w=5.73e-07 $l=4.3e-07 $layer=LI1_cond $X=9.132 $Y=3.245
+ $X2=9.132 $Y2=2.815
r173 31 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.645 $Y=3.245
+ $X2=6.645 $Y2=3.33
r174 31 33 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=6.645 $Y=3.245
+ $X2=6.645 $Y2=3.025
r175 27 89 2.12513 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=3.245
+ $X2=4.11 $Y2=3.33
r176 27 29 10.0846 $w=5.08e-07 $l=4.3e-07 $layer=LI1_cond $X=4.11 $Y=3.245
+ $X2=4.11 $Y2=2.815
r177 23 50 2.09999 $w=5.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.922 $Y=3.245
+ $X2=2.922 $Y2=3.33
r178 23 25 10.1844 $w=5.03e-07 $l=4.3e-07 $layer=LI1_cond $X=2.922 $Y=3.245
+ $X2=2.922 $Y2=2.815
r179 19 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=3.245
+ $X2=0.89 $Y2=3.33
r180 19 21 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=0.89 $Y=3.245
+ $X2=0.89 $Y2=2.465
r181 6 44 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=10.17
+ $Y=1.84 $X2=10.315 $Y2=2.815
r182 6 41 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.17
+ $Y=1.84 $X2=10.315 $Y2=1.985
r183 5 37 600 $w=1.7e-07 $l=3.81772e-07 $layer=licon1_PDIFF $count=1 $X=8.875
+ $Y=2.54 $X2=9.13 $Y2=2.815
r184 4 33 600 $w=1.7e-07 $l=5.84744e-07 $layer=licon1_PDIFF $count=1 $X=6.425
+ $Y=2.54 $X2=6.645 $Y2=3.025
r185 3 29 600 $w=1.7e-07 $l=1.08616e-06 $layer=licon1_PDIFF $count=1 $X=3.875
+ $Y=1.84 $X2=4.11 $Y2=2.815
r186 2 25 600 $w=1.7e-07 $l=6.29285e-07 $layer=licon1_PDIFF $count=1 $X=2.615
+ $Y=2.32 $X2=2.92 $Y2=2.815
r187 1 21 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=0.705
+ $Y=2.32 $X2=0.89 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_1%A_301_74# 1 2 3 4 13 19 22 23 24 26 27 30
+ 31 32 34 36 37 39 42 43 44 49
c134 44 0 7.022e-20 $X=4.31 $Y=2.435
c135 39 0 7.72654e-20 $X=5.21 $Y=2.805
c136 31 0 1.89404e-19 $X=4.615 $Y=1.565
c137 30 0 8.2679e-20 $X=4.31 $Y=2.31
r138 46 49 3.34041 $w=3.43e-07 $l=1e-07 $layer=LI1_cond $X=4.7 $Y=0.767 $X2=4.8
+ $Y2=0.767
r139 44 45 16.3723 $w=2.31e-07 $l=3.1e-07 $layer=LI1_cond $X=4.31 $Y=2.435
+ $X2=4.62 $Y2=2.435
r140 37 39 21.555 $w=2.68e-07 $l=5.05e-07 $layer=LI1_cond $X=4.705 $Y=2.845
+ $X2=5.21 $Y2=2.845
r141 35 46 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=4.7 $Y=0.94 $X2=4.7
+ $Y2=0.767
r142 35 36 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=4.7 $Y=0.94 $X2=4.7
+ $Y2=1.48
r143 34 37 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=4.62 $Y=2.71
+ $X2=4.705 $Y2=2.845
r144 33 45 2.5345 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.62 $Y=2.56
+ $X2=4.62 $Y2=2.435
r145 33 34 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=4.62 $Y=2.56
+ $X2=4.62 $Y2=2.71
r146 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.615 $Y=1.565
+ $X2=4.7 $Y2=1.48
r147 31 32 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.615 $Y=1.565
+ $X2=4.395 $Y2=1.565
r148 30 44 2.5345 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.31 $Y=2.31
+ $X2=4.31 $Y2=2.435
r149 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.31 $Y=1.65
+ $X2=4.395 $Y2=1.565
r150 29 30 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=4.31 $Y=1.65
+ $X2=4.31 $Y2=2.31
r151 28 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.395
+ $X2=2.995 $Y2=2.395
r152 27 44 51.8401 $w=2.31e-07 $l=9.84797e-07 $layer=LI1_cond $X=3.345 $Y=2.395
+ $X2=4.31 $Y2=2.435
r153 27 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.345 $Y=2.395
+ $X2=3.08 $Y2=2.395
r154 26 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=2.31
+ $X2=2.995 $Y2=2.395
r155 25 26 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=2.995 $Y=1.3
+ $X2=2.995 $Y2=2.31
r156 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.91 $Y=1.215
+ $X2=2.995 $Y2=1.3
r157 23 24 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.91 $Y=1.215
+ $X2=2.59 $Y2=1.215
r158 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.505 $Y=1.13
+ $X2=2.59 $Y2=1.215
r159 21 22 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.505 $Y=0.73
+ $X2=2.505 $Y2=1.13
r160 20 42 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.925 $Y=2.395
+ $X2=1.76 $Y2=2.395
r161 19 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.91 $Y=2.395
+ $X2=2.995 $Y2=2.395
r162 19 20 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=2.91 $Y=2.395
+ $X2=1.925 $Y2=2.395
r163 13 21 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.42 $Y=0.565
+ $X2=2.505 $Y2=0.73
r164 13 15 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=2.42 $Y=0.565
+ $X2=1.815 $Y2=0.565
r165 4 39 600 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_PDIFF $count=1 $X=5.065
+ $Y=2.54 $X2=5.21 $Y2=2.805
r166 3 42 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=1.625
+ $Y=2.32 $X2=1.76 $Y2=2.475
r167 2 49 182 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=1 $X=4.675
+ $Y=0.5 $X2=4.8 $Y2=0.765
r168 1 15 182 $w=1.7e-07 $l=3.95664e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.37 $X2=1.815 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_1%Q 1 2 7 8 9 10 11 12 13
r13 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=10.767 $Y=2.405
+ $X2=10.767 $Y2=2.775
r14 11 12 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=10.767 $Y=1.985
+ $X2=10.767 $Y2=2.405
r15 10 11 11.0084 $w=3.33e-07 $l=3.2e-07 $layer=LI1_cond $X=10.767 $Y=1.665
+ $X2=10.767 $Y2=1.985
r16 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=10.767 $Y=1.295
+ $X2=10.767 $Y2=1.665
r17 8 9 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=10.767 $Y=0.925
+ $X2=10.767 $Y2=1.295
r18 7 8 13.4165 $w=3.33e-07 $l=3.9e-07 $layer=LI1_cond $X=10.767 $Y=0.535
+ $X2=10.767 $Y2=0.925
r19 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.63
+ $Y=1.84 $X2=10.765 $Y2=2.815
r20 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.63
+ $Y=1.84 $X2=10.765 $Y2=1.985
r21 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.63
+ $Y=0.39 $X2=10.77 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_1%VGND 1 2 3 4 5 6 21 25 29 33 37 41 44 45 47
+ 48 49 51 66 73 78 85 86 89 92 95 100
r124 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r125 96 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=8.88
+ $Y2=0
r126 95 98 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r127 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r128 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r129 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r130 86 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r131 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r132 83 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.425 $Y=0
+ $X2=10.3 $Y2=0
r133 83 85 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=10.425 $Y=0
+ $X2=10.8 $Y2=0
r134 82 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r135 82 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r136 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r137 79 95 13.399 $w=1.7e-07 $l=3.38e-07 $layer=LI1_cond $X=9.48 $Y=0 $X2=9.142
+ $Y2=0
r138 79 81 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=9.48 $Y=0 $X2=9.84
+ $Y2=0
r139 78 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.175 $Y=0
+ $X2=10.3 $Y2=0
r140 78 81 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=10.175 $Y=0
+ $X2=9.84 $Y2=0
r141 77 98 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=8.88 $Y2=0
r142 77 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r143 76 77 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r144 74 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.635 $Y=0 $X2=6.51
+ $Y2=0
r145 74 76 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.635 $Y=0
+ $X2=6.96 $Y2=0
r146 73 95 13.399 $w=1.7e-07 $l=3.37e-07 $layer=LI1_cond $X=8.805 $Y=0 $X2=9.142
+ $Y2=0
r147 73 76 120.369 $w=1.68e-07 $l=1.845e-06 $layer=LI1_cond $X=8.805 $Y=0
+ $X2=6.96 $Y2=0
r148 72 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r149 71 72 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r150 68 71 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r151 68 69 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r152 66 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.385 $Y=0 $X2=6.51
+ $Y2=0
r153 66 71 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.385 $Y=0 $X2=6
+ $Y2=0
r154 65 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r155 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r156 62 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r157 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r158 59 62 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r159 59 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r160 58 61 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r161 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r162 56 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.75
+ $Y2=0
r163 56 58 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.2
+ $Y2=0
r164 54 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r165 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r166 51 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.75
+ $Y2=0
r167 51 53 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r168 49 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r169 49 69 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=4.08 $Y2=0
r170 47 64 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.6
+ $Y2=0
r171 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.85
+ $Y2=0
r172 46 68 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.015 $Y=0 $X2=4.08
+ $Y2=0
r173 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.015 $Y=0 $X2=3.85
+ $Y2=0
r174 44 61 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.775 $Y=0
+ $X2=2.64 $Y2=0
r175 44 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.86
+ $Y2=0
r176 43 64 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.945 $Y=0 $X2=3.6
+ $Y2=0
r177 43 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=0 $X2=2.86
+ $Y2=0
r178 39 100 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.3 $Y=0.085
+ $X2=10.3 $Y2=0
r179 39 41 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=10.3 $Y=0.085
+ $X2=10.3 $Y2=0.535
r180 35 95 2.78459 $w=6.75e-07 $l=8.5e-08 $layer=LI1_cond $X=9.142 $Y=0.085
+ $X2=9.142 $Y2=0
r181 35 37 9.92302 $w=6.73e-07 $l=5.6e-07 $layer=LI1_cond $X=9.142 $Y=0.085
+ $X2=9.142 $Y2=0.645
r182 31 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.51 $Y=0.085
+ $X2=6.51 $Y2=0
r183 31 33 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=6.51 $Y=0.085
+ $X2=6.51 $Y2=0.355
r184 27 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=0.085
+ $X2=3.85 $Y2=0
r185 27 29 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.85 $Y=0.085
+ $X2=3.85 $Y2=0.525
r186 23 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=0.085
+ $X2=2.86 $Y2=0
r187 23 25 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.86 $Y=0.085
+ $X2=2.86 $Y2=0.625
r188 19 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r189 19 21 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.565
r190 6 41 91 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_NDIFF $count=2 $X=10.21
+ $Y=0.39 $X2=10.34 $Y2=0.535
r191 5 37 91 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_NDIFF $count=2 $X=8.83
+ $Y=0.5 $X2=9.315 $Y2=0.645
r192 4 33 182 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=1 $X=6.345
+ $Y=0.5 $X2=6.55 $Y2=0.355
r193 3 29 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=3.705
+ $Y=0.37 $X2=3.85 $Y2=0.525
r194 2 25 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=2.64
+ $Y=0.37 $X2=2.86 $Y2=0.625
r195 1 21 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.61
+ $Y=0.37 $X2=0.75 $Y2=0.565
.ends


* File: sky130_fd_sc_ms__o311a_1.spice
* Created: Wed Sep  2 12:24:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o311a_1.pex.spice"
.subckt sky130_fd_sc_ms__o311a_1  VNB VPB C1 B1 A2 A3 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A3	A3
* A2	A2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1004 A_131_74# N_C1_M1004_g N_A_31_387#_M1004_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1824 PD=0.88 PS=1.85 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75003.4 A=0.096 P=1.58 MULT=1
MM1002 N_A_209_74#_M1002_d N_B1_M1002_g A_131_74# VNB NLOWVT L=0.15 W=0.64
+ AD=0.1248 AS=0.0768 PD=1.03 PS=0.88 NRD=7.488 NRS=12.18 M=1 R=4.26667
+ SA=75000.6 SB=75003.1 A=0.096 P=1.58 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g N_A_209_74#_M1002_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.1248 PD=1.21 PS=1.03 NRD=27.18 NRS=13.116 M=1 R=4.26667
+ SA=75001.1 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1005 N_A_209_74#_M1005_d N_A3_M1005_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.2976 AS=0.1824 PD=1.57 PS=1.21 NRD=0 NRS=27.18 M=1 R=4.26667 SA=75001.9
+ SB=75001.8 A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1000_d N_A1_M1000_g N_A_209_74#_M1005_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.118446 AS=0.2976 PD=1.02029 PS=1.57 NRD=0 NRS=14.988 M=1 R=4.26667
+ SA=75002.9 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1006 N_X_M1006_d N_A_31_387#_M1006_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.136954 PD=2.05 PS=1.17971 NRD=0 NRS=12.972 M=1 R=4.93333
+ SA=75003 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_VPWR_M1010_d N_C1_M1010_g N_A_31_387#_M1010_s VPB PSHORT L=0.18 W=1
+ AD=0.185 AS=0.28 PD=1.37 PS=2.56 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90003.5 A=0.18 P=2.36 MULT=1
MM1008 N_A_31_387#_M1008_d N_B1_M1008_g N_VPWR_M1010_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.185 PD=1.27 PS=1.37 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90000.7
+ SB=90002.9 A=0.18 P=2.36 MULT=1
MM1009 A_323_387# N_A3_M1009_g N_A_31_387#_M1008_d VPB PSHORT L=0.18 W=1 AD=0.45
+ AS=0.135 PD=1.9 PS=1.27 NRD=77.7953 NRS=0 M=1 R=5.55556 SA=90001.2 SB=90002.5
+ A=0.18 P=2.36 MULT=1
MM1003 A_539_387# N_A2_M1003_g A_323_387# VPB PSHORT L=0.18 W=1 AD=0.195 AS=0.45
+ PD=1.39 PS=1.9 NRD=27.5603 NRS=77.7953 M=1 R=5.55556 SA=90002.3 SB=90001.4
+ A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g A_539_387# VPB PSHORT L=0.18 W=1 AD=0.222642
+ AS=0.195 PD=1.4717 PS=1.39 NRD=22.6353 NRS=27.5603 M=1 R=5.55556 SA=90002.8
+ SB=90000.8 A=0.18 P=2.36 MULT=1
MM1011 N_X_M1011_d N_A_31_387#_M1011_g N_VPWR_M1001_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.249358 PD=2.8 PS=1.6483 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90003.1 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__o311a_1.pxi.spice"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nand3b_4 A_N B C VGND VNB VPB VPWR Y
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 Y a_89_172# a_744_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 a_297_82# B a_744_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VGND C a_297_82# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_297_82# B a_744_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_744_74# a_89_172# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_297_82# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_89_172# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_744_74# a_89_172# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_89_172# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X10 a_297_82# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 VPWR B Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X12 Y a_89_172# a_744_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 VPWR C Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X14 Y C VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 VPWR a_89_172# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X16 VGND C a_297_82# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 Y a_89_172# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X18 a_744_74# B a_297_82# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 VPWR A_N a_89_172# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X20 a_744_74# B a_297_82# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__sedfxtp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__sedfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.36000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.110000 0.805000 1.780000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.515000 1.320000 1.845000 1.780000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.502100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.475000 0.350000 14.815000 2.980000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.180000 5.280000 1.745000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.400000 1.180000 4.730000 1.510000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 6.330000 1.180000 6.660000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 15.360000 0.085000 ;
        RECT  1.080000  0.085000  1.410000 0.810000 ;
        RECT  2.070000  0.085000  2.400000 0.995000 ;
        RECT  4.755000  0.085000  5.005000 1.010000 ;
        RECT  6.020000  0.085000  6.280000 0.905000 ;
        RECT  7.005000  0.085000  7.335000 0.670000 ;
        RECT  9.750000  0.085000 10.000000 0.680000 ;
        RECT 11.190000  0.085000 11.440000 0.685000 ;
        RECT 12.800000  0.085000 13.755000 0.600000 ;
        RECT 14.995000  0.085000 15.245000 1.130000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
        RECT 15.035000 -0.085000 15.205000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 15.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 15.360000 3.415000 ;
        RECT  0.945000 2.630000  1.195000 3.245000 ;
        RECT  2.385000 2.630000  2.635000 3.245000 ;
        RECT  4.880000 2.595000  5.130000 3.245000 ;
        RECT  6.160000 2.670000  6.490000 3.245000 ;
        RECT  7.510000 2.670000  7.840000 3.245000 ;
        RECT  9.865000 2.730000 10.195000 3.245000 ;
        RECT 10.905000 2.730000 11.235000 3.245000 ;
        RECT 13.330000 2.650000 13.785000 3.245000 ;
        RECT 15.005000 1.820000 15.255000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
        RECT 14.555000 3.245000 14.725000 3.415000 ;
        RECT 15.035000 3.245000 15.205000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 15.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.085000 0.480000  0.590000 0.810000 ;
      RECT  0.085000 0.810000  0.255000 2.290000 ;
      RECT  0.085000 2.290000  1.535000 2.460000 ;
      RECT  0.085000 2.460000  0.435000 2.980000 ;
      RECT  0.975000 0.980000  1.890000 0.995000 ;
      RECT  0.975000 0.995000  1.810000 1.150000 ;
      RECT  0.975000 1.150000  1.305000 1.950000 ;
      RECT  0.975000 1.950000  2.385000 2.120000 ;
      RECT  1.365000 2.460000  1.535000 2.905000 ;
      RECT  1.365000 2.905000  2.215000 3.075000 ;
      RECT  1.640000 0.535000  1.890000 0.980000 ;
      RECT  1.705000 2.120000  1.875000 2.735000 ;
      RECT  2.045000 2.290000  3.395000 2.460000 ;
      RECT  2.045000 2.460000  2.215000 2.905000 ;
      RECT  2.055000 1.520000  2.385000 1.950000 ;
      RECT  2.555000 1.505000  3.055000 1.835000 ;
      RECT  2.890000 0.535000  3.220000 1.165000 ;
      RECT  2.890000 1.165000  3.395000 1.335000 ;
      RECT  3.145000 2.460000  3.395000 2.975000 ;
      RECT  3.225000 1.335000  3.395000 2.290000 ;
      RECT  3.390000 0.535000  3.735000 0.995000 ;
      RECT  3.565000 0.995000  3.735000 2.295000 ;
      RECT  3.565000 2.295000  3.845000 2.905000 ;
      RECT  3.565000 2.905000  4.710000 3.075000 ;
      RECT  3.905000 0.255000  4.185000 0.605000 ;
      RECT  3.905000 0.605000  4.575000 1.010000 ;
      RECT  3.905000 1.010000  4.185000 1.915000 ;
      RECT  3.905000 1.915000  5.820000 2.085000 ;
      RECT  4.015000 2.085000  4.185000 2.255000 ;
      RECT  4.015000 2.255000  4.370000 2.735000 ;
      RECT  4.540000 2.255000  6.160000 2.330000 ;
      RECT  4.540000 2.330000  8.180000 2.425000 ;
      RECT  4.540000 2.425000  4.710000 2.905000 ;
      RECT  5.465000 0.605000  5.795000 1.075000 ;
      RECT  5.465000 1.075000  6.160000 1.245000 ;
      RECT  5.490000 1.415000  5.820000 1.915000 ;
      RECT  5.640000 2.425000  8.180000 2.500000 ;
      RECT  5.640000 2.500000  5.990000 2.935000 ;
      RECT  5.990000 1.245000  6.160000 2.255000 ;
      RECT  6.450000 0.350000  6.780000 0.840000 ;
      RECT  6.450000 0.840000  7.000000 1.010000 ;
      RECT  6.610000 1.760000  7.000000 1.830000 ;
      RECT  6.610000 1.830000  7.390000 2.160000 ;
      RECT  6.830000 1.010000  7.000000 1.760000 ;
      RECT  7.515000 0.255000  9.255000 0.425000 ;
      RECT  7.515000 0.425000  7.765000 1.130000 ;
      RECT  7.620000 1.480000  8.235000 1.650000 ;
      RECT  7.620000 1.650000  7.790000 2.330000 ;
      RECT  7.960000 1.820000  8.575000 1.990000 ;
      RECT  7.960000 1.990000  8.665000 2.160000 ;
      RECT  7.985000 0.595000  8.235000 1.480000 ;
      RECT  8.010000 2.500000  8.180000 2.730000 ;
      RECT  8.010000 2.730000  8.815000 2.980000 ;
      RECT  8.405000 0.425000  8.575000 1.820000 ;
      RECT  8.405000 2.160000  8.665000 2.335000 ;
      RECT  8.745000 0.595000  8.915000 1.620000 ;
      RECT  8.745000 1.620000 10.465000 1.790000 ;
      RECT  8.835000 1.790000  9.005000 2.390000 ;
      RECT  8.835000 2.390000  9.315000 2.560000 ;
      RECT  8.985000 2.560000  9.315000 2.980000 ;
      RECT  9.085000 0.425000  9.255000 0.850000 ;
      RECT  9.085000 0.850000 10.340000 1.020000 ;
      RECT  9.085000 1.020000  9.340000 1.345000 ;
      RECT  9.175000 1.960000  9.655000 2.220000 ;
      RECT  9.485000 2.220000  9.655000 2.390000 ;
      RECT  9.485000 2.390000 12.200000 2.560000 ;
      RECT  9.565000 1.190000  9.895000 1.195000 ;
      RECT  9.565000 1.195000 11.385000 1.365000 ;
      RECT  9.565000 1.365000  9.895000 1.450000 ;
      RECT 10.135000 1.535000 10.465000 1.620000 ;
      RECT 10.135000 1.790000 10.465000 1.795000 ;
      RECT 10.170000 0.255000 11.020000 0.425000 ;
      RECT 10.170000 0.425000 10.340000 0.850000 ;
      RECT 10.385000 1.970000 10.805000 2.220000 ;
      RECT 10.510000 0.595000 10.680000 1.195000 ;
      RECT 10.635000 1.365000 11.385000 1.525000 ;
      RECT 10.635000 1.525000 10.805000 1.970000 ;
      RECT 10.850000 0.425000 11.020000 0.855000 ;
      RECT 10.850000 0.855000 11.730000 1.025000 ;
      RECT 11.560000 1.025000 11.730000 1.110000 ;
      RECT 11.560000 1.110000 13.005000 1.280000 ;
      RECT 11.560000 1.280000 11.860000 1.800000 ;
      RECT 11.900000 0.350000 12.230000 0.770000 ;
      RECT 11.900000 0.770000 13.345000 0.940000 ;
      RECT 12.030000 1.450000 12.465000 1.735000 ;
      RECT 12.030000 1.735000 12.200000 2.390000 ;
      RECT 12.370000 1.940000 12.805000 2.980000 ;
      RECT 12.635000 1.735000 13.785000 1.905000 ;
      RECT 12.635000 1.905000 12.805000 1.940000 ;
      RECT 12.675000 1.280000 13.005000 1.555000 ;
      RECT 13.065000 2.075000 14.285000 2.380000 ;
      RECT 13.175000 0.940000 13.345000 1.735000 ;
      RECT 13.615000 1.050000 13.945000 1.380000 ;
      RECT 13.615000 1.380000 13.785000 1.735000 ;
      RECT 13.925000 0.350000 14.285000 0.810000 ;
      RECT 13.955000 2.380000 14.285000 2.980000 ;
      RECT 14.045000 1.550000 14.285000 2.075000 ;
      RECT 14.115000 0.810000 14.285000 1.550000 ;
    LAYER mcon ;
      RECT  2.555000 1.580000  2.725000 1.750000 ;
      RECT 14.075000 1.580000 14.245000 1.750000 ;
    LAYER met1 ;
      RECT  2.495000 1.550000  2.785000 1.595000 ;
      RECT  2.495000 1.595000 14.305000 1.735000 ;
      RECT  2.495000 1.735000  2.785000 1.780000 ;
      RECT 14.015000 1.550000 14.305000 1.595000 ;
      RECT 14.015000 1.735000 14.305000 1.780000 ;
  END
END sky130_fd_sc_ms__sedfxtp_1

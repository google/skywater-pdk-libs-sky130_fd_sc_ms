* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__xnor2_2 A B VGND VNB VPB VPWR Y
M1000 Y B a_641_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=8.894e+11p ps=6.2e+06u
M1001 a_340_107# B VGND VNB nlowvt w=740000u l=150000u
+  ad=8.30525e+11p pd=8.22e+06u as=1.024e+12p ps=7.92e+06u
M1002 VPWR A a_641_368# VPB pshort w=1.12e+06u l=180000u
+  ad=2.16185e+12p pd=1.301e+07u as=0p ps=0u
M1003 a_641_368# B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y a_136_368# a_340_107# VNB nlowvt w=740000u l=150000u
+  ad=4.008e+11p pd=2.67e+06u as=0p ps=0u
M1005 VGND B a_340_107# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A a_340_107# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_340_107# A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_641_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_136_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_136_368# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_136_368# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=3.15e+11p pd=2.63e+06u as=0p ps=0u
M1012 VPWR B a_136_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_136_368# B a_151_74# VNB nlowvt w=740000u l=150000u
+  ad=2.06875e+11p pd=2.05e+06u as=1.776e+11p ps=1.96e+06u
M1014 a_151_74# A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_340_107# a_136_368# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

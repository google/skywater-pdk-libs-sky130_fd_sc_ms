* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfstp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
X0 VPWR a_599_74# a_800_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 a_998_81# a_599_74# a_1131_457# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X2 VPWR a_998_81# a_1613_341# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X3 VPWR SCE a_208_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X4 a_2395_112# a_1764_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X5 a_599_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VGND a_2395_112# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_292_464# a_27_464# a_418_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X8 VPWR SET_B a_1764_74# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X9 a_1686_74# a_800_74# a_1764_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X10 a_208_464# D a_292_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X11 a_238_74# D a_292_464# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X12 a_1198_55# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X13 a_1721_374# a_800_74# a_1764_74# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X14 a_292_464# a_800_74# a_998_81# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X15 a_998_81# a_800_74# a_1150_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X16 VGND a_998_81# a_1686_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X17 VPWR a_2395_112# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X18 a_418_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X19 VPWR a_998_81# a_1198_55# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X20 a_1910_74# a_1958_48# a_1988_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X21 a_1426_118# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X22 a_1988_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X23 a_402_74# SCD VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X24 a_1958_48# a_1764_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X25 a_27_464# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X26 a_292_464# SCE a_402_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X27 a_599_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X28 a_292_464# a_599_74# a_998_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X29 VGND a_27_464# a_238_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X30 a_1150_81# a_1198_55# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X31 a_1721_374# a_1958_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X32 VGND a_1764_74# a_1958_48# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X33 a_1131_457# a_1198_55# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X34 a_1764_74# a_599_74# a_1910_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X35 a_1764_74# a_599_74# a_1613_341# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X36 a_1198_55# a_998_81# a_1426_118# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X37 VGND a_599_74# a_800_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X38 a_2395_112# a_1764_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X39 a_27_464# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
.ends

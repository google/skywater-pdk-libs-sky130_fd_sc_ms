* NGSPICE file created from sky130_fd_sc_ms__a21boi_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 a_436_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=5.994e+11p pd=6.06e+06u as=4.144e+11p ps=4.08e+06u
M1001 Y a_62_94# a_241_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.1872e+12p ps=1.108e+07u
M1002 a_241_368# a_62_94# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND B1_N a_62_94# VNB nlowvt w=640000u l=150000u
+  ad=6.474e+11p pd=6.21e+06u as=1.696e+11p ps=1.81e+06u
M1004 VPWR A1 a_241_368# VPB pshort w=1.12e+06u l=180000u
+  ad=8.872e+11p pd=8.12e+06u as=0p ps=0u
M1005 a_241_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y a_62_94# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_436_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A2 a_241_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_241_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_62_94# B1_N VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1011 VGND a_62_94# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A1 a_436_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_436_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__nand2b_1.pxi.spice
* Created: Wed Sep  2 12:13:09 2020
* 
x_PM_SKY130_FD_SC_MS__NAND2B_1%A_N N_A_N_M1002_g N_A_N_M1003_g A_N A_N
+ N_A_N_c_47_n PM_SKY130_FD_SC_MS__NAND2B_1%A_N
x_PM_SKY130_FD_SC_MS__NAND2B_1%B N_B_M1004_g N_B_M1001_g B N_B_c_80_n N_B_c_81_n
+ PM_SKY130_FD_SC_MS__NAND2B_1%B
x_PM_SKY130_FD_SC_MS__NAND2B_1%A_27_112# N_A_27_112#_M1003_s N_A_27_112#_M1002_s
+ N_A_27_112#_M1000_g N_A_27_112#_M1005_g N_A_27_112#_c_123_n
+ N_A_27_112#_c_124_n N_A_27_112#_c_125_n N_A_27_112#_c_138_n
+ N_A_27_112#_c_130_n N_A_27_112#_c_131_n N_A_27_112#_c_126_n
+ N_A_27_112#_c_127_n N_A_27_112#_c_128_n PM_SKY130_FD_SC_MS__NAND2B_1%A_27_112#
x_PM_SKY130_FD_SC_MS__NAND2B_1%VPWR N_VPWR_M1002_d N_VPWR_M1005_d N_VPWR_c_196_n
+ N_VPWR_c_197_n N_VPWR_c_198_n N_VPWR_c_199_n VPWR N_VPWR_c_200_n
+ N_VPWR_c_195_n N_VPWR_c_202_n PM_SKY130_FD_SC_MS__NAND2B_1%VPWR
x_PM_SKY130_FD_SC_MS__NAND2B_1%Y N_Y_M1000_d N_Y_M1004_d N_Y_c_228_n N_Y_c_225_n
+ N_Y_c_226_n N_Y_c_227_n Y Y N_Y_c_232_n PM_SKY130_FD_SC_MS__NAND2B_1%Y
x_PM_SKY130_FD_SC_MS__NAND2B_1%VGND N_VGND_M1003_d N_VGND_c_261_n VGND
+ N_VGND_c_262_n N_VGND_c_263_n N_VGND_c_264_n N_VGND_c_265_n
+ PM_SKY130_FD_SC_MS__NAND2B_1%VGND
cc_1 VNB N_A_N_M1002_g 0.00191101f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_2 VNB N_A_N_M1003_g 0.031967f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_3 VNB A_N 0.0177819f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_A_N_c_47_n 0.0638847f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.465
cc_5 VNB N_B_M1001_g 0.0274125f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_6 VNB N_B_c_80_n 0.0271913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_B_c_81_n 0.00182951f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_8 VNB N_A_27_112#_M1000_g 0.0248499f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_9 VNB N_A_27_112#_M1005_g 0.001621f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_10 VNB N_A_27_112#_c_123_n 0.0188303f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.465
cc_11 VNB N_A_27_112#_c_124_n 0.0153597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_112#_c_125_n 0.00869634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_112#_c_126_n 0.00981133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_112#_c_127_n 0.0327357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_112#_c_128_n 0.00161243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_195_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_225_n 0.027835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_226_n 0.0250664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_227_n 0.0158601f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_20 VNB N_VGND_c_261_n 0.0155608f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_21 VNB N_VGND_c_262_n 0.0182319f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_22 VNB N_VGND_c_263_n 0.0364261f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.465
cc_23 VNB N_VGND_c_264_n 0.175015f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.465
cc_24 VNB N_VGND_c_265_n 0.0126977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VPB N_A_N_M1002_g 0.0309988f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_26 VPB A_N 0.0110509f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_27 VPB N_B_M1004_g 0.0233901f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_28 VPB N_B_c_80_n 0.00576405f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_29 VPB N_B_c_81_n 0.00270771f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.465
cc_30 VPB N_A_27_112#_M1005_g 0.0253282f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.465
cc_31 VPB N_A_27_112#_c_130_n 0.00135795f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB N_A_27_112#_c_131_n 0.0331749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_196_n 0.0193212f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_197_n 0.021977f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.465
cc_35 VPB N_VPWR_c_198_n 0.0221255f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.54
cc_36 VPB N_VPWR_c_199_n 0.00622357f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_200_n 0.0126445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_195_n 0.0726209f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_202_n 0.0264241f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_Y_c_228_n 0.0169104f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.835
cc_41 VPB N_Y_c_226_n 0.0313588f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB Y 0.00275815f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.465
cc_43 N_A_N_M1002_g N_B_M1004_g 0.0237085f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_44 A_N N_B_M1004_g 3.87236e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_45 N_A_N_M1003_g N_B_M1001_g 0.00900688f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_46 A_N N_B_M1001_g 0.00113012f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_47 N_A_N_c_47_n N_B_M1001_g 0.00121331f $X=0.61 $Y=1.465 $X2=0 $Y2=0
cc_48 N_A_N_M1002_g N_B_c_80_n 0.00119089f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_49 A_N N_B_c_80_n 0.00227619f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_50 N_A_N_c_47_n N_B_c_80_n 0.014832f $X=0.61 $Y=1.465 $X2=0 $Y2=0
cc_51 N_A_N_M1002_g N_B_c_81_n 2.81447e-19 $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_52 A_N N_B_c_81_n 0.0350659f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_53 N_A_N_c_47_n N_B_c_81_n 3.13222e-19 $X=0.61 $Y=1.465 $X2=0 $Y2=0
cc_54 N_A_N_M1003_g N_A_27_112#_c_123_n 0.0020078f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_55 N_A_N_M1003_g N_A_27_112#_c_124_n 0.015445f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_56 A_N N_A_27_112#_c_124_n 0.0348645f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_57 N_A_N_c_47_n N_A_27_112#_c_124_n 0.00560904f $X=0.61 $Y=1.465 $X2=0 $Y2=0
cc_58 A_N N_A_27_112#_c_125_n 0.0226786f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_59 N_A_N_c_47_n N_A_27_112#_c_125_n 0.00613776f $X=0.61 $Y=1.465 $X2=0 $Y2=0
cc_60 N_A_N_M1002_g N_A_27_112#_c_138_n 0.0139134f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_61 A_N N_A_27_112#_c_138_n 0.0282304f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_62 N_A_N_c_47_n N_A_27_112#_c_138_n 7.85743e-19 $X=0.61 $Y=1.465 $X2=0 $Y2=0
cc_63 N_A_N_M1002_g N_A_27_112#_c_131_n 0.0111437f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_64 A_N N_A_27_112#_c_131_n 0.0266342f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_65 N_A_N_c_47_n N_A_27_112#_c_131_n 0.00152954f $X=0.61 $Y=1.465 $X2=0 $Y2=0
cc_66 N_A_N_M1002_g N_VPWR_c_196_n 0.00612139f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_67 N_A_N_M1002_g N_VPWR_c_195_n 0.00555093f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_68 N_A_N_M1002_g N_VPWR_c_202_n 0.00465228f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_69 N_A_N_M1003_g N_VGND_c_261_n 0.010935f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_70 N_A_N_M1003_g N_VGND_c_262_n 0.003901f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_71 N_A_N_M1003_g N_VGND_c_264_n 0.00425985f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_72 N_B_M1001_g N_A_27_112#_M1000_g 0.0373316f $X=1.27 $Y=0.74 $X2=0 $Y2=0
cc_73 N_B_M1004_g N_A_27_112#_M1005_g 0.027494f $X=1.175 $Y=2.4 $X2=0 $Y2=0
cc_74 N_B_c_81_n N_A_27_112#_M1005_g 3.06787e-19 $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_75 N_B_M1001_g N_A_27_112#_c_124_n 0.0156214f $X=1.27 $Y=0.74 $X2=0 $Y2=0
cc_76 N_B_c_80_n N_A_27_112#_c_124_n 0.00118587f $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_77 N_B_c_81_n N_A_27_112#_c_124_n 0.0202397f $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_78 N_B_M1004_g N_A_27_112#_c_138_n 0.0128784f $X=1.175 $Y=2.4 $X2=0 $Y2=0
cc_79 N_B_c_80_n N_A_27_112#_c_138_n 5.95231e-19 $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_80 N_B_c_81_n N_A_27_112#_c_138_n 0.0208858f $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_81 N_B_M1004_g N_A_27_112#_c_130_n 0.00352936f $X=1.175 $Y=2.4 $X2=0 $Y2=0
cc_82 N_B_M1004_g N_A_27_112#_c_131_n 7.33428e-19 $X=1.175 $Y=2.4 $X2=0 $Y2=0
cc_83 N_B_c_80_n N_A_27_112#_c_126_n 0.00330428f $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_84 N_B_c_81_n N_A_27_112#_c_126_n 0.0341497f $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_85 N_B_c_80_n N_A_27_112#_c_127_n 0.0373316f $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_86 N_B_c_81_n N_A_27_112#_c_127_n 3.65128e-19 $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_87 N_B_M1001_g N_A_27_112#_c_128_n 0.00330428f $X=1.27 $Y=0.74 $X2=0 $Y2=0
cc_88 N_B_M1004_g N_VPWR_c_196_n 0.0109164f $X=1.175 $Y=2.4 $X2=0 $Y2=0
cc_89 N_B_M1004_g N_VPWR_c_197_n 6.13365e-19 $X=1.175 $Y=2.4 $X2=0 $Y2=0
cc_90 N_B_M1004_g N_VPWR_c_198_n 0.00350949f $X=1.175 $Y=2.4 $X2=0 $Y2=0
cc_91 N_B_M1004_g N_VPWR_c_195_n 0.00434146f $X=1.175 $Y=2.4 $X2=0 $Y2=0
cc_92 N_B_M1004_g Y 0.0130729f $X=1.175 $Y=2.4 $X2=0 $Y2=0
cc_93 N_B_M1004_g N_Y_c_232_n 0.00544733f $X=1.175 $Y=2.4 $X2=0 $Y2=0
cc_94 N_B_M1001_g N_VGND_c_261_n 0.0172792f $X=1.27 $Y=0.74 $X2=0 $Y2=0
cc_95 N_B_M1001_g N_VGND_c_263_n 0.00383152f $X=1.27 $Y=0.74 $X2=0 $Y2=0
cc_96 N_B_M1001_g N_VGND_c_264_n 0.0075725f $X=1.27 $Y=0.74 $X2=0 $Y2=0
cc_97 N_A_27_112#_c_138_n N_VPWR_M1002_d 0.0170839f $X=1.515 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_98 N_A_27_112#_c_138_n N_VPWR_c_196_n 0.0213159f $X=1.515 $Y=2.035 $X2=0
+ $Y2=0
cc_99 N_A_27_112#_c_131_n N_VPWR_c_196_n 0.0139143f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_100 N_A_27_112#_M1005_g N_VPWR_c_197_n 0.00955692f $X=1.675 $Y=2.4 $X2=0
+ $Y2=0
cc_101 N_A_27_112#_M1005_g N_VPWR_c_198_n 0.00460063f $X=1.675 $Y=2.4 $X2=0
+ $Y2=0
cc_102 N_A_27_112#_M1005_g N_VPWR_c_195_n 0.00909121f $X=1.675 $Y=2.4 $X2=0
+ $Y2=0
cc_103 N_A_27_112#_c_131_n N_VPWR_c_195_n 0.00995531f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_104 N_A_27_112#_c_131_n N_VPWR_c_202_n 0.0066444f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_105 N_A_27_112#_c_138_n N_Y_M1004_d 0.008851f $X=1.515 $Y=2.035 $X2=0 $Y2=0
cc_106 N_A_27_112#_c_130_n N_Y_M1004_d 0.00134282f $X=1.6 $Y=1.95 $X2=0 $Y2=0
cc_107 N_A_27_112#_M1005_g N_Y_c_228_n 0.0170459f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_108 N_A_27_112#_c_138_n N_Y_c_228_n 0.00754135f $X=1.515 $Y=2.035 $X2=0 $Y2=0
cc_109 N_A_27_112#_c_126_n N_Y_c_228_n 0.00485682f $X=1.75 $Y=1.465 $X2=0 $Y2=0
cc_110 N_A_27_112#_c_127_n N_Y_c_228_n 5.46639e-19 $X=1.75 $Y=1.465 $X2=0 $Y2=0
cc_111 N_A_27_112#_M1000_g N_Y_c_225_n 0.0221957f $X=1.66 $Y=0.74 $X2=0 $Y2=0
cc_112 N_A_27_112#_M1000_g N_Y_c_226_n 0.00292854f $X=1.66 $Y=0.74 $X2=0 $Y2=0
cc_113 N_A_27_112#_M1005_g N_Y_c_226_n 0.0141327f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_114 N_A_27_112#_c_138_n N_Y_c_226_n 0.00712876f $X=1.515 $Y=2.035 $X2=0 $Y2=0
cc_115 N_A_27_112#_c_130_n N_Y_c_226_n 0.0120688f $X=1.6 $Y=1.95 $X2=0 $Y2=0
cc_116 N_A_27_112#_c_126_n N_Y_c_226_n 0.0251716f $X=1.75 $Y=1.465 $X2=0 $Y2=0
cc_117 N_A_27_112#_c_127_n N_Y_c_226_n 0.00739878f $X=1.75 $Y=1.465 $X2=0 $Y2=0
cc_118 N_A_27_112#_c_128_n N_Y_c_226_n 0.00637596f $X=1.715 $Y=1.3 $X2=0 $Y2=0
cc_119 N_A_27_112#_c_124_n N_Y_c_227_n 0.0142393f $X=1.515 $Y=1.045 $X2=0 $Y2=0
cc_120 N_A_27_112#_c_126_n N_Y_c_227_n 0.0049152f $X=1.75 $Y=1.465 $X2=0 $Y2=0
cc_121 N_A_27_112#_c_127_n N_Y_c_227_n 4.59055e-19 $X=1.75 $Y=1.465 $X2=0 $Y2=0
cc_122 N_A_27_112#_c_138_n N_Y_c_232_n 0.0304989f $X=1.515 $Y=2.035 $X2=0 $Y2=0
cc_123 N_A_27_112#_c_124_n N_VGND_M1003_d 0.00761754f $X=1.515 $Y=1.045
+ $X2=-0.19 $Y2=-0.245
cc_124 N_A_27_112#_M1000_g N_VGND_c_261_n 0.00188096f $X=1.66 $Y=0.74 $X2=0
+ $Y2=0
cc_125 N_A_27_112#_c_123_n N_VGND_c_261_n 0.0112176f $X=0.28 $Y=0.835 $X2=0
+ $Y2=0
cc_126 N_A_27_112#_c_124_n N_VGND_c_261_n 0.0447655f $X=1.515 $Y=1.045 $X2=0
+ $Y2=0
cc_127 N_A_27_112#_c_123_n N_VGND_c_262_n 0.00651231f $X=0.28 $Y=0.835 $X2=0
+ $Y2=0
cc_128 N_A_27_112#_M1000_g N_VGND_c_263_n 0.00461464f $X=1.66 $Y=0.74 $X2=0
+ $Y2=0
cc_129 N_A_27_112#_M1000_g N_VGND_c_264_n 0.00913279f $X=1.66 $Y=0.74 $X2=0
+ $Y2=0
cc_130 N_A_27_112#_c_123_n N_VGND_c_264_n 0.00849993f $X=0.28 $Y=0.835 $X2=0
+ $Y2=0
cc_131 N_A_27_112#_c_124_n A_269_74# 0.00485986f $X=1.515 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_132 N_VPWR_M1005_d N_Y_c_228_n 0.0103861f $X=1.765 $Y=1.84 $X2=0 $Y2=0
cc_133 N_VPWR_c_197_n N_Y_c_228_n 0.0205361f $X=1.9 $Y=2.815 $X2=0 $Y2=0
cc_134 N_VPWR_c_196_n Y 0.0408335f $X=0.82 $Y=2.455 $X2=0 $Y2=0
cc_135 N_VPWR_c_197_n Y 0.0132475f $X=1.9 $Y=2.815 $X2=0 $Y2=0
cc_136 N_VPWR_c_198_n Y 0.0208154f $X=1.735 $Y=3.33 $X2=0 $Y2=0
cc_137 N_VPWR_c_195_n Y 0.0167995f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_138 N_VPWR_c_196_n N_Y_c_232_n 0.0137881f $X=0.82 $Y=2.455 $X2=0 $Y2=0
cc_139 N_Y_c_225_n N_VGND_c_261_n 0.0128668f $X=1.94 $Y=0.515 $X2=0 $Y2=0
cc_140 N_Y_c_225_n N_VGND_c_263_n 0.0177591f $X=1.94 $Y=0.515 $X2=0 $Y2=0
cc_141 N_Y_c_225_n N_VGND_c_264_n 0.0146995f $X=1.94 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__o2111a_2.pxi.spice
* Created: Fri Aug 28 17:51:37 2020
* 
x_PM_SKY130_FD_SC_MS__O2111A_2%A1 N_A1_M1006_g N_A1_c_78_n N_A1_M1007_g A1 A1
+ N_A1_c_80_n PM_SKY130_FD_SC_MS__O2111A_2%A1
x_PM_SKY130_FD_SC_MS__O2111A_2%A2 N_A2_M1011_g N_A2_M1003_g A2 N_A2_c_103_n
+ N_A2_c_104_n PM_SKY130_FD_SC_MS__O2111A_2%A2
x_PM_SKY130_FD_SC_MS__O2111A_2%B1 N_B1_M1010_g N_B1_M1013_g B1 N_B1_c_134_n
+ N_B1_c_135_n PM_SKY130_FD_SC_MS__O2111A_2%B1
x_PM_SKY130_FD_SC_MS__O2111A_2%C1 N_C1_M1005_g N_C1_M1002_g C1 N_C1_c_171_n
+ PM_SKY130_FD_SC_MS__O2111A_2%C1
x_PM_SKY130_FD_SC_MS__O2111A_2%D1 N_D1_M1008_g N_D1_M1000_g D1 N_D1_c_212_n
+ N_D1_c_213_n PM_SKY130_FD_SC_MS__O2111A_2%D1
x_PM_SKY130_FD_SC_MS__O2111A_2%A_239_368# N_A_239_368#_M1008_d
+ N_A_239_368#_M1011_d N_A_239_368#_M1002_d N_A_239_368#_M1001_g
+ N_A_239_368#_M1004_g N_A_239_368#_M1012_g N_A_239_368#_M1009_g
+ N_A_239_368#_c_262_n N_A_239_368#_c_263_n N_A_239_368#_c_273_n
+ N_A_239_368#_c_264_n N_A_239_368#_c_283_n N_A_239_368#_c_254_n
+ N_A_239_368#_c_255_n N_A_239_368#_c_256_n N_A_239_368#_c_257_n
+ N_A_239_368#_c_258_n N_A_239_368#_c_286_n N_A_239_368#_c_259_n
+ PM_SKY130_FD_SC_MS__O2111A_2%A_239_368#
x_PM_SKY130_FD_SC_MS__O2111A_2%VPWR N_VPWR_M1006_s N_VPWR_M1010_d N_VPWR_M1000_d
+ N_VPWR_M1012_d N_VPWR_c_364_n N_VPWR_c_365_n N_VPWR_c_366_n N_VPWR_c_367_n
+ N_VPWR_c_368_n N_VPWR_c_369_n N_VPWR_c_370_n N_VPWR_c_371_n N_VPWR_c_372_n
+ VPWR N_VPWR_c_373_n N_VPWR_c_374_n N_VPWR_c_375_n N_VPWR_c_363_n
+ PM_SKY130_FD_SC_MS__O2111A_2%VPWR
x_PM_SKY130_FD_SC_MS__O2111A_2%X N_X_M1004_s N_X_M1001_s N_X_c_424_n N_X_c_425_n
+ N_X_c_421_n X X X PM_SKY130_FD_SC_MS__O2111A_2%X
x_PM_SKY130_FD_SC_MS__O2111A_2%A_54_74# N_A_54_74#_M1007_s N_A_54_74#_M1003_d
+ N_A_54_74#_c_453_n N_A_54_74#_c_454_n N_A_54_74#_c_459_n N_A_54_74#_c_465_n
+ N_A_54_74#_c_455_n PM_SKY130_FD_SC_MS__O2111A_2%A_54_74#
x_PM_SKY130_FD_SC_MS__O2111A_2%VGND N_VGND_M1007_d N_VGND_M1004_d N_VGND_M1009_d
+ N_VGND_c_480_n N_VGND_c_481_n N_VGND_c_482_n N_VGND_c_483_n VGND
+ N_VGND_c_484_n N_VGND_c_485_n N_VGND_c_486_n N_VGND_c_487_n N_VGND_c_488_n
+ N_VGND_c_489_n PM_SKY130_FD_SC_MS__O2111A_2%VGND
cc_1 VNB N_A1_M1006_g 0.00923934f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=2.34
cc_2 VNB N_A1_c_78_n 0.023452f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.22
cc_3 VNB A1 0.0291142f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_A1_c_80_n 0.0688992f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_5 VNB N_A2_M1011_g 0.00654075f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.55
cc_6 VNB A2 0.00596829f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.74
cc_7 VNB N_A2_c_103_n 0.0326603f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_8 VNB N_A2_c_104_n 0.0186009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B1_M1010_g 0.00712091f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.55
cc_10 VNB B1 0.00892781f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.74
cc_11 VNB N_B1_c_134_n 0.0306617f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_12 VNB N_B1_c_135_n 0.0183068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_C1_M1005_g 0.026905f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.55
cc_14 VNB C1 0.0121385f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.74
cc_15 VNB N_C1_c_171_n 0.0282571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_D1_M1008_g 0.030729f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.55
cc_17 VNB N_D1_c_212_n 0.0377416f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_18 VNB N_D1_c_213_n 0.00305137f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_19 VNB N_A_239_368#_M1001_g 0.00174353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_239_368#_M1004_g 0.0223898f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_21 VNB N_A_239_368#_M1012_g 0.00231818f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.365
cc_22 VNB N_A_239_368#_M1009_g 0.0266858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_239_368#_c_254_n 0.00994708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_239_368#_c_255_n 0.0187701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_239_368#_c_256_n 0.00248805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_239_368#_c_257_n 0.0094184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_239_368#_c_258_n 4.18697e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_239_368#_c_259_n 0.0719033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_363_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_X_c_421_n 0.00270411f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_31 VNB X 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_32 VNB X 0.00448002f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_33 VNB N_A_54_74#_c_453_n 0.00716827f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.22
cc_34 VNB N_A_54_74#_c_454_n 0.0217137f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.74
cc_35 VNB N_A_54_74#_c_455_n 0.00280313f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_36 VNB N_VGND_c_480_n 0.00460613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_481_n 0.0145024f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_38 VNB N_VGND_c_482_n 0.0109665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_483_n 0.0516149f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.365
cc_40 VNB N_VGND_c_484_n 0.0232895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_485_n 0.0643439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_486_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_487_n 0.00866122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_488_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_489_n 0.308027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VPB N_A1_M1006_g 0.0283462f $X=-0.19 $Y=1.66 $X2=0.685 $Y2=2.34
cc_47 VPB N_A2_M1011_g 0.0236104f $X=-0.19 $Y=1.66 $X2=0.685 $Y2=1.55
cc_48 VPB N_B1_M1010_g 0.0255736f $X=-0.19 $Y=1.66 $X2=0.685 $Y2=1.55
cc_49 VPB N_C1_M1002_g 0.0223716f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.22
cc_50 VPB C1 0.0052439f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=0.74
cc_51 VPB N_C1_c_171_n 0.00556231f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_D1_M1000_g 0.0236449f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.22
cc_53 VPB N_D1_c_212_n 0.0117843f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_54 VPB N_D1_c_213_n 0.00444735f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_55 VPB N_A_239_368#_M1001_g 0.0238771f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_239_368#_M1012_g 0.0273944f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.365
cc_57 VPB N_A_239_368#_c_262_n 0.00998062f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_239_368#_c_263_n 0.00340823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_239_368#_c_264_n 0.00341904f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_239_368#_c_258_n 0.00339199f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_364_n 0.0610756f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_62 VPB N_VPWR_c_365_n 0.0198717f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.365
cc_63 VPB N_VPWR_c_366_n 0.017832f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_367_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_368_n 0.0693112f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_369_n 0.0115308f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_370_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_371_n 0.0348258f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_372_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_373_n 0.0220157f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_374_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_375_n 0.0155543f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_363_n 0.0958345f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_X_c_424_n 0.00412671f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=0.74
cc_75 VPB N_X_c_425_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_76 VPB N_X_c_421_n 8.13921e-19 $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_77 N_A1_M1006_g N_A2_M1011_g 0.0466303f $X=0.685 $Y=2.34 $X2=0 $Y2=0
cc_78 A1 A2 0.029889f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_79 N_A1_c_80_n A2 3.68035e-19 $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_80 A1 N_A2_c_103_n 0.00216087f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_81 N_A1_c_80_n N_A2_c_103_n 0.0466303f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_82 N_A1_c_78_n N_A2_c_104_n 0.0268292f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_83 N_A1_M1006_g N_VPWR_c_364_n 0.0272975f $X=0.685 $Y=2.34 $X2=0 $Y2=0
cc_84 A1 N_VPWR_c_364_n 0.0195859f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_85 N_A1_c_80_n N_VPWR_c_364_n 0.00656875f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_86 N_A1_M1006_g N_VPWR_c_371_n 0.00492916f $X=0.685 $Y=2.34 $X2=0 $Y2=0
cc_87 N_A1_M1006_g N_VPWR_c_363_n 0.00511769f $X=0.685 $Y=2.34 $X2=0 $Y2=0
cc_88 A1 N_A_54_74#_c_453_n 0.0282818f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_89 N_A1_c_80_n N_A_54_74#_c_453_n 0.00229697f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_90 N_A1_c_78_n N_A_54_74#_c_454_n 8.37507e-19 $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_91 N_A1_c_78_n N_A_54_74#_c_459_n 0.0102656f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_92 A1 N_A_54_74#_c_459_n 0.0153343f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_93 N_A1_c_78_n N_VGND_c_480_n 0.0159254f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_94 N_A1_c_78_n N_VGND_c_484_n 0.00383152f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_95 N_A1_c_78_n N_VGND_c_489_n 0.00388149f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_96 N_A2_M1011_g N_B1_M1010_g 0.0262179f $X=1.105 $Y=2.34 $X2=0 $Y2=0
cc_97 A2 B1 0.0242365f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_98 N_A2_c_104_n B1 0.00228667f $X=1.18 $Y=1.22 $X2=0 $Y2=0
cc_99 A2 N_B1_c_134_n 4.06701e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_100 N_A2_c_103_n N_B1_c_134_n 0.0175474f $X=1.18 $Y=1.385 $X2=0 $Y2=0
cc_101 N_A2_c_104_n N_B1_c_135_n 0.0198524f $X=1.18 $Y=1.22 $X2=0 $Y2=0
cc_102 N_A2_M1011_g N_A_239_368#_c_262_n 0.0048092f $X=1.105 $Y=2.34 $X2=0 $Y2=0
cc_103 A2 N_A_239_368#_c_262_n 0.00356336f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_104 N_A2_c_103_n N_A_239_368#_c_262_n 4.37254e-19 $X=1.18 $Y=1.385 $X2=0
+ $Y2=0
cc_105 N_A2_M1011_g N_A_239_368#_c_263_n 0.0110517f $X=1.105 $Y=2.34 $X2=0 $Y2=0
cc_106 N_A2_M1011_g N_VPWR_c_364_n 0.00362989f $X=1.105 $Y=2.34 $X2=0 $Y2=0
cc_107 N_A2_M1011_g N_VPWR_c_371_n 0.0059286f $X=1.105 $Y=2.34 $X2=0 $Y2=0
cc_108 N_A2_M1011_g N_VPWR_c_363_n 0.00610055f $X=1.105 $Y=2.34 $X2=0 $Y2=0
cc_109 A2 N_A_54_74#_c_459_n 0.0228656f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_110 N_A2_c_103_n N_A_54_74#_c_459_n 9.98643e-19 $X=1.18 $Y=1.385 $X2=0 $Y2=0
cc_111 N_A2_c_104_n N_A_54_74#_c_459_n 0.0126376f $X=1.18 $Y=1.22 $X2=0 $Y2=0
cc_112 N_A2_c_104_n N_A_54_74#_c_455_n 0.0026172f $X=1.18 $Y=1.22 $X2=0 $Y2=0
cc_113 N_A2_c_104_n N_VGND_c_480_n 0.0131556f $X=1.18 $Y=1.22 $X2=0 $Y2=0
cc_114 N_A2_c_104_n N_VGND_c_485_n 0.00383152f $X=1.18 $Y=1.22 $X2=0 $Y2=0
cc_115 N_A2_c_104_n N_VGND_c_489_n 0.00384679f $X=1.18 $Y=1.22 $X2=0 $Y2=0
cc_116 B1 N_C1_M1005_g 0.00173356f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_117 N_B1_c_134_n N_C1_M1005_g 0.0179214f $X=1.75 $Y=1.385 $X2=0 $Y2=0
cc_118 N_B1_c_135_n N_C1_M1005_g 0.0415061f $X=1.75 $Y=1.22 $X2=0 $Y2=0
cc_119 N_B1_M1010_g N_C1_M1002_g 0.0205753f $X=1.675 $Y=2.34 $X2=0 $Y2=0
cc_120 N_B1_M1010_g C1 0.00293713f $X=1.675 $Y=2.34 $X2=0 $Y2=0
cc_121 B1 C1 0.0119739f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_122 N_B1_c_134_n C1 7.31814e-19 $X=1.75 $Y=1.385 $X2=0 $Y2=0
cc_123 N_B1_M1010_g N_C1_c_171_n 0.00356318f $X=1.675 $Y=2.34 $X2=0 $Y2=0
cc_124 B1 N_C1_c_171_n 2.54315e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_125 N_B1_M1010_g N_A_239_368#_c_262_n 0.00413137f $X=1.675 $Y=2.34 $X2=0
+ $Y2=0
cc_126 B1 N_A_239_368#_c_262_n 0.00290148f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_127 N_B1_M1010_g N_A_239_368#_c_263_n 0.0108548f $X=1.675 $Y=2.34 $X2=0 $Y2=0
cc_128 N_B1_M1010_g N_A_239_368#_c_273_n 0.0150233f $X=1.675 $Y=2.34 $X2=0 $Y2=0
cc_129 B1 N_A_239_368#_c_273_n 0.0100691f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_130 N_B1_c_134_n N_A_239_368#_c_273_n 6.88201e-19 $X=1.75 $Y=1.385 $X2=0
+ $Y2=0
cc_131 N_B1_M1010_g N_A_239_368#_c_264_n 6.20636e-19 $X=1.675 $Y=2.34 $X2=0
+ $Y2=0
cc_132 N_B1_M1010_g N_VPWR_c_365_n 0.00361649f $X=1.675 $Y=2.34 $X2=0 $Y2=0
cc_133 N_B1_M1010_g N_VPWR_c_371_n 0.00567889f $X=1.675 $Y=2.34 $X2=0 $Y2=0
cc_134 N_B1_M1010_g N_VPWR_c_363_n 0.00610055f $X=1.675 $Y=2.34 $X2=0 $Y2=0
cc_135 B1 N_A_54_74#_c_465_n 0.0107224f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_136 N_B1_c_134_n N_A_54_74#_c_465_n 6.09387e-19 $X=1.75 $Y=1.385 $X2=0 $Y2=0
cc_137 N_B1_c_135_n N_A_54_74#_c_465_n 0.00377406f $X=1.75 $Y=1.22 $X2=0 $Y2=0
cc_138 N_B1_c_135_n N_A_54_74#_c_455_n 0.00985605f $X=1.75 $Y=1.22 $X2=0 $Y2=0
cc_139 N_B1_c_135_n N_VGND_c_480_n 6.14068e-19 $X=1.75 $Y=1.22 $X2=0 $Y2=0
cc_140 N_B1_c_135_n N_VGND_c_485_n 0.00434272f $X=1.75 $Y=1.22 $X2=0 $Y2=0
cc_141 N_B1_c_135_n N_VGND_c_489_n 0.00822352f $X=1.75 $Y=1.22 $X2=0 $Y2=0
cc_142 N_C1_M1005_g N_D1_M1008_g 0.034788f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_143 N_C1_M1002_g N_D1_M1000_g 0.0112311f $X=2.315 $Y=2.34 $X2=0 $Y2=0
cc_144 C1 N_D1_M1000_g 0.00287029f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_145 C1 N_D1_c_212_n 0.0105656f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_146 N_C1_c_171_n N_D1_c_212_n 0.0182087f $X=2.32 $Y=1.515 $X2=0 $Y2=0
cc_147 C1 N_D1_c_213_n 0.0341872f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_148 N_C1_c_171_n N_D1_c_213_n 2.00281e-19 $X=2.32 $Y=1.515 $X2=0 $Y2=0
cc_149 N_C1_M1002_g N_A_239_368#_c_262_n 5.719e-19 $X=2.315 $Y=2.34 $X2=0 $Y2=0
cc_150 N_C1_M1002_g N_A_239_368#_c_263_n 8.42462e-19 $X=2.315 $Y=2.34 $X2=0
+ $Y2=0
cc_151 N_C1_M1002_g N_A_239_368#_c_273_n 0.0138062f $X=2.315 $Y=2.34 $X2=0 $Y2=0
cc_152 C1 N_A_239_368#_c_273_n 0.0144161f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_153 N_C1_c_171_n N_A_239_368#_c_273_n 2.7382e-19 $X=2.32 $Y=1.515 $X2=0 $Y2=0
cc_154 N_C1_M1002_g N_A_239_368#_c_264_n 0.0125423f $X=2.315 $Y=2.34 $X2=0 $Y2=0
cc_155 C1 N_A_239_368#_c_283_n 0.0030217f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_156 N_C1_M1005_g N_A_239_368#_c_254_n 0.00300965f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_157 N_C1_M1005_g N_A_239_368#_c_256_n 7.70038e-19 $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_158 N_C1_M1002_g N_A_239_368#_c_286_n 8.84614e-19 $X=2.315 $Y=2.34 $X2=0
+ $Y2=0
cc_159 C1 N_A_239_368#_c_286_n 0.0246997f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_160 N_C1_c_171_n N_A_239_368#_c_286_n 3.50164e-19 $X=2.32 $Y=1.515 $X2=0
+ $Y2=0
cc_161 N_C1_M1002_g N_VPWR_c_365_n 0.00852005f $X=2.315 $Y=2.34 $X2=0 $Y2=0
cc_162 N_C1_M1002_g N_VPWR_c_366_n 5.72044e-19 $X=2.315 $Y=2.34 $X2=0 $Y2=0
cc_163 N_C1_M1002_g N_VPWR_c_373_n 0.0056753f $X=2.315 $Y=2.34 $X2=0 $Y2=0
cc_164 N_C1_M1002_g N_VPWR_c_363_n 0.00610055f $X=2.315 $Y=2.34 $X2=0 $Y2=0
cc_165 N_C1_M1005_g N_A_54_74#_c_465_n 8.11227e-19 $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_166 N_C1_M1005_g N_A_54_74#_c_455_n 0.00235594f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_167 N_C1_M1005_g N_VGND_c_485_n 0.00461464f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_168 N_C1_M1005_g N_VGND_c_489_n 0.00910941f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_169 N_D1_c_212_n N_A_239_368#_M1001_g 9.94734e-19 $X=3.09 $Y=1.515 $X2=0
+ $Y2=0
cc_170 N_D1_M1000_g N_A_239_368#_c_264_n 3.48084e-19 $X=2.815 $Y=2.34 $X2=0
+ $Y2=0
cc_171 N_D1_M1000_g N_A_239_368#_c_283_n 0.0209075f $X=2.815 $Y=2.34 $X2=0 $Y2=0
cc_172 N_D1_c_212_n N_A_239_368#_c_283_n 0.00172067f $X=3.09 $Y=1.515 $X2=0
+ $Y2=0
cc_173 N_D1_c_213_n N_A_239_368#_c_283_n 0.0249341f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_174 N_D1_M1008_g N_A_239_368#_c_254_n 0.015254f $X=2.8 $Y=0.74 $X2=0 $Y2=0
cc_175 N_D1_c_212_n N_A_239_368#_c_255_n 5.19479e-19 $X=3.09 $Y=1.515 $X2=0
+ $Y2=0
cc_176 N_D1_c_213_n N_A_239_368#_c_255_n 0.00566599f $X=3.09 $Y=1.515 $X2=0
+ $Y2=0
cc_177 N_D1_M1008_g N_A_239_368#_c_256_n 0.006714f $X=2.8 $Y=0.74 $X2=0 $Y2=0
cc_178 N_D1_c_212_n N_A_239_368#_c_256_n 0.00439517f $X=3.09 $Y=1.515 $X2=0
+ $Y2=0
cc_179 N_D1_c_213_n N_A_239_368#_c_256_n 0.021921f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_180 N_D1_M1008_g N_A_239_368#_c_257_n 0.00277277f $X=2.8 $Y=0.74 $X2=0 $Y2=0
cc_181 N_D1_c_212_n N_A_239_368#_c_257_n 0.00116423f $X=3.09 $Y=1.515 $X2=0
+ $Y2=0
cc_182 N_D1_c_213_n N_A_239_368#_c_257_n 0.0150172f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_183 N_D1_M1000_g N_A_239_368#_c_258_n 0.00390173f $X=2.815 $Y=2.34 $X2=0
+ $Y2=0
cc_184 N_D1_c_212_n N_A_239_368#_c_258_n 4.17225e-19 $X=3.09 $Y=1.515 $X2=0
+ $Y2=0
cc_185 N_D1_c_213_n N_A_239_368#_c_258_n 0.00860661f $X=3.09 $Y=1.515 $X2=0
+ $Y2=0
cc_186 N_D1_M1008_g N_A_239_368#_c_259_n 6.46057e-19 $X=2.8 $Y=0.74 $X2=0 $Y2=0
cc_187 N_D1_c_212_n N_A_239_368#_c_259_n 0.0140828f $X=3.09 $Y=1.515 $X2=0 $Y2=0
cc_188 N_D1_c_213_n N_A_239_368#_c_259_n 3.56038e-19 $X=3.09 $Y=1.515 $X2=0
+ $Y2=0
cc_189 N_D1_M1000_g N_VPWR_c_366_n 0.0127492f $X=2.815 $Y=2.34 $X2=0 $Y2=0
cc_190 N_D1_M1000_g N_VPWR_c_373_n 0.00492916f $X=2.815 $Y=2.34 $X2=0 $Y2=0
cc_191 N_D1_M1000_g N_VPWR_c_363_n 0.00511769f $X=2.815 $Y=2.34 $X2=0 $Y2=0
cc_192 N_D1_M1008_g N_VGND_c_481_n 0.00373386f $X=2.8 $Y=0.74 $X2=0 $Y2=0
cc_193 N_D1_M1008_g N_VGND_c_485_n 0.00434272f $X=2.8 $Y=0.74 $X2=0 $Y2=0
cc_194 N_D1_M1008_g N_VGND_c_489_n 0.00827521f $X=2.8 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A_239_368#_c_273_n N_VPWR_M1010_d 0.0166166f $X=2.375 $Y=2.035 $X2=0
+ $Y2=0
cc_196 N_A_239_368#_c_283_n N_VPWR_M1000_d 0.0250217f $X=3.515 $Y=2.035 $X2=0
+ $Y2=0
cc_197 N_A_239_368#_c_258_n N_VPWR_M1000_d 0.00263868f $X=3.6 $Y=1.95 $X2=0
+ $Y2=0
cc_198 N_A_239_368#_c_262_n N_VPWR_c_364_n 0.00823114f $X=1.45 $Y=2.12 $X2=0
+ $Y2=0
cc_199 N_A_239_368#_c_263_n N_VPWR_c_364_n 0.0195279f $X=1.45 $Y=2.695 $X2=0
+ $Y2=0
cc_200 N_A_239_368#_c_263_n N_VPWR_c_365_n 0.0221782f $X=1.45 $Y=2.695 $X2=0
+ $Y2=0
cc_201 N_A_239_368#_c_273_n N_VPWR_c_365_n 0.0237567f $X=2.375 $Y=2.035 $X2=0
+ $Y2=0
cc_202 N_A_239_368#_c_264_n N_VPWR_c_365_n 0.0331287f $X=2.54 $Y=2.375 $X2=0
+ $Y2=0
cc_203 N_A_239_368#_M1001_g N_VPWR_c_366_n 0.00523041f $X=3.795 $Y=2.4 $X2=0
+ $Y2=0
cc_204 N_A_239_368#_c_264_n N_VPWR_c_366_n 0.0263584f $X=2.54 $Y=2.375 $X2=0
+ $Y2=0
cc_205 N_A_239_368#_c_283_n N_VPWR_c_366_n 0.0590682f $X=3.515 $Y=2.035 $X2=0
+ $Y2=0
cc_206 N_A_239_368#_c_259_n N_VPWR_c_366_n 4.61822e-19 $X=4.245 $Y=1.465 $X2=0
+ $Y2=0
cc_207 N_A_239_368#_M1012_g N_VPWR_c_368_n 0.00546761f $X=4.245 $Y=2.4 $X2=0
+ $Y2=0
cc_208 N_A_239_368#_c_259_n N_VPWR_c_368_n 3.5215e-19 $X=4.245 $Y=1.465 $X2=0
+ $Y2=0
cc_209 N_A_239_368#_c_263_n N_VPWR_c_371_n 0.00975961f $X=1.45 $Y=2.695 $X2=0
+ $Y2=0
cc_210 N_A_239_368#_c_264_n N_VPWR_c_373_n 0.010336f $X=2.54 $Y=2.375 $X2=0
+ $Y2=0
cc_211 N_A_239_368#_M1001_g N_VPWR_c_374_n 0.005209f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_212 N_A_239_368#_M1012_g N_VPWR_c_374_n 0.005209f $X=4.245 $Y=2.4 $X2=0 $Y2=0
cc_213 N_A_239_368#_M1001_g N_VPWR_c_363_n 0.00986727f $X=3.795 $Y=2.4 $X2=0
+ $Y2=0
cc_214 N_A_239_368#_M1012_g N_VPWR_c_363_n 0.00985497f $X=4.245 $Y=2.4 $X2=0
+ $Y2=0
cc_215 N_A_239_368#_c_263_n N_VPWR_c_363_n 0.0111753f $X=1.45 $Y=2.695 $X2=0
+ $Y2=0
cc_216 N_A_239_368#_c_264_n N_VPWR_c_363_n 0.0113305f $X=2.54 $Y=2.375 $X2=0
+ $Y2=0
cc_217 N_A_239_368#_M1001_g N_X_c_424_n 0.003664f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_218 N_A_239_368#_M1012_g N_X_c_424_n 0.00215936f $X=4.245 $Y=2.4 $X2=0 $Y2=0
cc_219 N_A_239_368#_c_258_n N_X_c_424_n 0.00559274f $X=3.6 $Y=1.95 $X2=0 $Y2=0
cc_220 N_A_239_368#_c_259_n N_X_c_424_n 0.0018941f $X=4.245 $Y=1.465 $X2=0 $Y2=0
cc_221 N_A_239_368#_M1001_g N_X_c_425_n 0.0182659f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_222 N_A_239_368#_M1012_g N_X_c_425_n 0.0127634f $X=4.245 $Y=2.4 $X2=0 $Y2=0
cc_223 N_A_239_368#_M1001_g N_X_c_421_n 0.00111019f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_224 N_A_239_368#_M1004_g N_X_c_421_n 0.00104557f $X=3.86 $Y=0.74 $X2=0 $Y2=0
cc_225 N_A_239_368#_M1012_g N_X_c_421_n 0.00959299f $X=4.245 $Y=2.4 $X2=0 $Y2=0
cc_226 N_A_239_368#_M1009_g N_X_c_421_n 0.00455396f $X=4.29 $Y=0.74 $X2=0 $Y2=0
cc_227 N_A_239_368#_c_257_n N_X_c_421_n 0.0293979f $X=3.6 $Y=1.63 $X2=0 $Y2=0
cc_228 N_A_239_368#_c_258_n N_X_c_421_n 0.00661604f $X=3.6 $Y=1.95 $X2=0 $Y2=0
cc_229 N_A_239_368#_c_259_n N_X_c_421_n 0.0261549f $X=4.245 $Y=1.465 $X2=0 $Y2=0
cc_230 N_A_239_368#_M1004_g X 0.0122719f $X=3.86 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A_239_368#_M1009_g X 0.00788704f $X=4.29 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A_239_368#_M1004_g X 0.0048722f $X=3.86 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A_239_368#_M1009_g X 0.00327512f $X=4.29 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A_239_368#_c_257_n X 0.00802092f $X=3.6 $Y=1.63 $X2=0 $Y2=0
cc_235 N_A_239_368#_c_255_n N_VGND_M1004_d 0.00138568f $X=3.515 $Y=1.095 $X2=0
+ $Y2=0
cc_236 N_A_239_368#_c_257_n N_VGND_M1004_d 0.00384491f $X=3.6 $Y=1.63 $X2=0
+ $Y2=0
cc_237 N_A_239_368#_M1004_g N_VGND_c_481_n 0.00634966f $X=3.86 $Y=0.74 $X2=0
+ $Y2=0
cc_238 N_A_239_368#_c_254_n N_VGND_c_481_n 0.032024f $X=3.015 $Y=0.515 $X2=0
+ $Y2=0
cc_239 N_A_239_368#_c_255_n N_VGND_c_481_n 0.00796924f $X=3.515 $Y=1.095 $X2=0
+ $Y2=0
cc_240 N_A_239_368#_c_257_n N_VGND_c_481_n 0.0161682f $X=3.6 $Y=1.63 $X2=0 $Y2=0
cc_241 N_A_239_368#_c_259_n N_VGND_c_481_n 0.00103859f $X=4.245 $Y=1.465 $X2=0
+ $Y2=0
cc_242 N_A_239_368#_M1009_g N_VGND_c_483_n 0.00650681f $X=4.29 $Y=0.74 $X2=0
+ $Y2=0
cc_243 N_A_239_368#_c_254_n N_VGND_c_485_n 0.0145639f $X=3.015 $Y=0.515 $X2=0
+ $Y2=0
cc_244 N_A_239_368#_M1004_g N_VGND_c_486_n 0.00434272f $X=3.86 $Y=0.74 $X2=0
+ $Y2=0
cc_245 N_A_239_368#_M1009_g N_VGND_c_486_n 0.00434272f $X=4.29 $Y=0.74 $X2=0
+ $Y2=0
cc_246 N_A_239_368#_M1004_g N_VGND_c_489_n 0.00825059f $X=3.86 $Y=0.74 $X2=0
+ $Y2=0
cc_247 N_A_239_368#_M1009_g N_VGND_c_489_n 0.00823992f $X=4.29 $Y=0.74 $X2=0
+ $Y2=0
cc_248 N_A_239_368#_c_254_n N_VGND_c_489_n 0.0119984f $X=3.015 $Y=0.515 $X2=0
+ $Y2=0
cc_249 N_VPWR_c_368_n N_X_c_424_n 0.0450694f $X=4.52 $Y=1.985 $X2=0 $Y2=0
cc_250 N_VPWR_c_366_n N_X_c_425_n 0.0267725f $X=3.52 $Y=2.375 $X2=0 $Y2=0
cc_251 N_VPWR_c_374_n N_X_c_425_n 0.0144623f $X=4.355 $Y=3.33 $X2=0 $Y2=0
cc_252 N_VPWR_c_363_n N_X_c_425_n 0.0118344f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_253 X N_VGND_c_481_n 0.0186136f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_254 X N_VGND_c_483_n 0.0293892f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_255 X N_VGND_c_486_n 0.0144922f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_256 X N_VGND_c_489_n 0.0118826f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_257 N_A_54_74#_c_459_n N_VGND_M1007_d 0.0117062f $X=1.39 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_258 N_A_54_74#_c_454_n N_VGND_c_480_n 0.013465f $X=0.485 $Y=0.515 $X2=0 $Y2=0
cc_259 N_A_54_74#_c_459_n N_VGND_c_480_n 0.0279268f $X=1.39 $Y=0.925 $X2=0 $Y2=0
cc_260 N_A_54_74#_c_455_n N_VGND_c_480_n 0.013465f $X=1.555 $Y=0.515 $X2=0 $Y2=0
cc_261 N_A_54_74#_c_454_n N_VGND_c_484_n 0.0146038f $X=0.485 $Y=0.515 $X2=0
+ $Y2=0
cc_262 N_A_54_74#_c_455_n N_VGND_c_485_n 0.0145323f $X=1.555 $Y=0.515 $X2=0
+ $Y2=0
cc_263 N_A_54_74#_c_454_n N_VGND_c_489_n 0.0121018f $X=0.485 $Y=0.515 $X2=0
+ $Y2=0
cc_264 N_A_54_74#_c_459_n N_VGND_c_489_n 0.0114395f $X=1.39 $Y=0.925 $X2=0 $Y2=0
cc_265 N_A_54_74#_c_455_n N_VGND_c_489_n 0.0119861f $X=1.555 $Y=0.515 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__nor4b_2.spice
* Created: Wed Sep  2 12:17:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nor4b_2.pex.spice"
.subckt sky130_fd_sc_ms__nor4b_2  VNB VPB D_N C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_D_N_M1000_g N_A_27_392#_M1000_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.136255 AS=0.1824 PD=1.07594 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75004.8 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1000_d N_A_27_392#_M1006_g N_Y_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.157545 AS=0.1295 PD=1.24406 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75004.3 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_27_392#_M1009_g N_Y_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1998 AS=0.1295 PD=1.28 PS=1.09 NRD=15.396 NRS=11.34 M=1 R=4.93333
+ SA=75001.2 SB=75003.8 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1009_d N_C_M1010_g N_Y_M1010_s VNB NLOWVT L=0.15 W=0.74 AD=0.1998
+ AS=0.1036 PD=1.28 PS=1.02 NRD=26.748 NRS=0 M=1 R=4.93333 SA=75001.9 SB=75003.1
+ A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_C_M1017_g N_Y_M1010_s VNB NLOWVT L=0.15 W=0.74 AD=0.148
+ AS=0.1036 PD=1.14 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.3 SB=75002.7
+ A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_B_M1002_g N_VGND_M1017_d VNB NLOWVT L=0.15 W=0.74 AD=0.1369
+ AS=0.148 PD=1.11 PS=1.14 NRD=3.24 NRS=8.1 M=1 R=4.93333 SA=75002.9 SB=75002.1
+ A=0.111 P=1.78 MULT=1
MM1011 N_Y_M1002_d N_B_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.74 AD=0.1369
+ AS=0.26825 PD=1.11 PS=1.465 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75003.4
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1011_s N_A_M1004_g N_Y_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.26825 AS=0.12395 PD=1.465 PS=1.075 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.3
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_A_M1013_g N_Y_M1004_s VNB NLOWVT L=0.15 W=0.74 AD=0.222
+ AS=0.12395 PD=2.08 PS=1.075 NRD=2.424 NRS=8.916 M=1 R=4.93333 SA=75004.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VPWR_M1001_d N_D_N_M1001_g N_A_27_392#_M1001_s VPB PSHORT L=0.18 W=1
+ AD=0.28 AS=0.28 PD=2.56 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1012 N_Y_M1012_d N_A_27_392#_M1012_g N_A_229_368#_M1012_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1014 N_Y_M1012_d N_A_27_392#_M1014_g N_A_229_368#_M1014_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1015 N_A_501_368#_M1015_d N_C_M1015_g N_A_229_368#_M1014_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.1 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1016 N_A_501_368#_M1015_d N_C_M1016_g N_A_229_368#_M1016_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1005 N_A_501_368#_M1005_d N_B_M1005_g N_A_701_368#_M1005_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1007 N_A_501_368#_M1005_d N_B_M1007_g N_A_701_368#_M1007_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1003 N_A_701_368#_M1007_s N_A_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1568 PD=1.39 PS=1.4 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1008 N_A_701_368#_M1008_d N_A_M1008_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1568 PD=2.8 PS=1.4 NRD=0 NRS=0.8668 M=1 R=6.22222 SA=90001.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX18_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ms__nor4b_2.pxi.spice"
*
.ends
*
*

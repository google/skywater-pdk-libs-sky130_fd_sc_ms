# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__sdfrtn_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__sdfrtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.780000 1.980000 2.120000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.530100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.475000 0.350000 13.805000 2.980000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.455400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  3.405000 1.355000  3.735000 2.025000 ;
        RECT  7.655000 1.470000  8.035000 1.800000 ;
        RECT 10.995000 1.210000 11.395000 1.540000 ;
        RECT 11.195000 1.540000 11.395000 1.780000 ;
      LAYER mcon ;
        RECT  3.515000 1.580000  3.685000 1.750000 ;
        RECT  7.835000 1.580000  8.005000 1.750000 ;
        RECT 11.195000 1.580000 11.365000 1.750000 ;
      LAYER met1 ;
        RECT  3.455000 1.550000  3.745000 1.595000 ;
        RECT  3.455000 1.595000 11.425000 1.735000 ;
        RECT  3.455000 1.735000  3.745000 1.780000 ;
        RECT  7.775000 1.550000  8.065000 1.595000 ;
        RECT  7.775000 1.735000  8.065000 1.780000 ;
        RECT 11.135000 1.550000 11.425000 1.595000 ;
        RECT 11.135000 1.735000 11.425000 1.780000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.800000 1.525000 3.235000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 1.410000 2.045000 1.580000 ;
        RECT 0.535000 1.580000 0.865000 2.080000 ;
        RECT 1.875000 0.955000 2.550000 1.410000 ;
    END
  END SCE
  PIN CLK_N
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.275000 1.210000 4.675000 1.550000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 13.920000 0.085000 ;
        RECT  0.615000  0.085000  0.945000 0.880000 ;
        RECT  3.655000  0.085000  3.985000 0.780000 ;
        RECT  4.835000  0.085000  5.165000 0.640000 ;
        RECT  7.890000  0.085000  8.220000 0.620000 ;
        RECT 10.730000  0.085000 11.200000 0.680000 ;
        RECT 12.975000  0.085000 13.305000 1.130000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.920000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 13.920000 3.415000 ;
        RECT  0.565000 2.630000  0.895000 3.245000 ;
        RECT  2.815000 2.970000  3.145000 3.245000 ;
        RECT  4.840000 2.550000  5.170000 3.245000 ;
        RECT  7.295000 2.360000  7.545000 3.245000 ;
        RECT  8.295000 2.310000  8.625000 3.245000 ;
        RECT 10.605000 2.650000 11.210000 3.245000 ;
        RECT 11.880000 2.630000 12.210000 3.245000 ;
        RECT 12.975000 1.820000 13.305000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 13.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.115000 0.420000  0.445000 1.050000 ;
      RECT  0.115000 1.050000  1.620000 1.240000 ;
      RECT  0.115000 1.240000  0.365000 2.290000 ;
      RECT  0.115000 2.290000  2.545000 2.460000 ;
      RECT  0.115000 2.460000  0.365000 2.980000 ;
      RECT  1.165000 0.255000  3.390000 0.425000 ;
      RECT  1.165000 0.425000  1.495000 0.765000 ;
      RECT  1.290000 0.935000  1.620000 1.050000 ;
      RECT  1.405000 2.630000  3.680000 2.800000 ;
      RECT  1.405000 2.800000  2.220000 2.960000 ;
      RECT  1.955000 0.595000  2.890000 0.765000 ;
      RECT  2.215000 1.580000  2.545000 2.290000 ;
      RECT  2.720000 0.765000  2.890000 0.960000 ;
      RECT  2.720000 0.960000  4.075000 1.185000 ;
      RECT  3.060000 0.425000  3.390000 0.780000 ;
      RECT  3.430000 2.300000  6.235000 2.380000 ;
      RECT  3.430000 2.380000  4.515000 2.600000 ;
      RECT  3.430000 2.600000  3.680000 2.630000 ;
      RECT  3.430000 2.800000  3.680000 2.980000 ;
      RECT  3.905000 1.185000  4.075000 2.180000 ;
      RECT  3.905000 2.180000  6.235000 2.300000 ;
      RECT  4.310000 1.820000  5.190000 2.010000 ;
      RECT  4.325000 0.395000  4.660000 0.810000 ;
      RECT  4.325000 0.810000  5.270000 1.010000 ;
      RECT  4.940000 1.010000  5.270000 1.220000 ;
      RECT  4.940000 1.220000  5.300000 1.575000 ;
      RECT  4.940000 1.575000  5.190000 1.820000 ;
      RECT  5.360000 1.745000  5.735000 2.010000 ;
      RECT  5.440000 0.255000  7.260000 0.465000 ;
      RECT  5.440000 0.465000  5.735000 1.090000 ;
      RECT  5.470000 1.090000  5.735000 1.745000 ;
      RECT  5.910000 0.635000  6.160000 1.840000 ;
      RECT  5.910000 1.840000  6.235000 2.180000 ;
      RECT  5.965000 2.380000  6.235000 2.705000 ;
      RECT  6.330000 0.465000  6.500000 1.670000 ;
      RECT  6.415000 2.275000  6.850000 2.705000 ;
      RECT  6.670000 0.635000  6.920000 1.075000 ;
      RECT  6.670000 1.075000  6.850000 1.970000 ;
      RECT  6.670000 1.970000  8.490000 2.140000 ;
      RECT  6.670000 2.140000  8.125000 2.190000 ;
      RECT  6.670000 2.190000  6.850000 2.275000 ;
      RECT  7.075000 1.470000  7.415000 1.800000 ;
      RECT  7.090000 0.465000  7.260000 0.790000 ;
      RECT  7.090000 0.790000  8.560000 0.960000 ;
      RECT  7.235000 1.130000  8.900000 1.300000 ;
      RECT  7.235000 1.300000  7.415000 1.470000 ;
      RECT  7.785000 2.190000  8.125000 2.705000 ;
      RECT  8.225000 1.470000  8.490000 1.970000 ;
      RECT  8.390000 0.360000  9.240000 0.530000 ;
      RECT  8.390000 0.530000  8.560000 0.790000 ;
      RECT  8.730000 0.700000  8.900000 1.130000 ;
      RECT  8.730000 1.300000  8.900000 1.970000 ;
      RECT  8.730000 1.970000  9.495000 2.165000 ;
      RECT  8.795000 2.165000  9.495000 2.980000 ;
      RECT  9.070000 0.530000  9.240000 1.030000 ;
      RECT  9.070000 1.030000  9.825000 1.200000 ;
      RECT  9.070000 1.370000 10.395000 1.540000 ;
      RECT  9.070000 1.540000  9.350000 1.800000 ;
      RECT  9.410000 0.530000 10.475000 0.860000 ;
      RECT  9.735000 1.710000 11.025000 1.880000 ;
      RECT  9.735000 1.880000 10.065000 2.980000 ;
      RECT 10.065000 1.290000 10.395000 1.370000 ;
      RECT 10.305000 0.860000 10.475000 0.870000 ;
      RECT 10.305000 0.870000 11.895000 1.040000 ;
      RECT 10.435000 2.050000 10.685000 2.290000 ;
      RECT 10.435000 2.290000 12.235000 2.460000 ;
      RECT 10.855000 1.880000 11.025000 1.950000 ;
      RECT 10.855000 1.950000 11.895000 2.120000 ;
      RECT 11.380000 2.460000 11.710000 2.980000 ;
      RECT 11.565000 1.040000 11.895000 1.950000 ;
      RECT 11.690000 0.450000 12.235000 0.700000 ;
      RECT 12.065000 0.700000 12.235000 2.290000 ;
      RECT 12.440000 0.350000 12.795000 1.355000 ;
      RECT 12.440000 1.355000 12.810000 1.685000 ;
      RECT 12.440000 1.685000 12.795000 2.980000 ;
  END
END sky130_fd_sc_ms__sdfrtn_1

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__o31ai_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__o31ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.315000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.350000 2.275000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.350000 3.445000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.685000 1.350000 4.695000 1.680000 ;
        RECT 4.365000 1.180000 4.695000 1.350000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.229800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.820000 2.835000 1.950000 ;
        RECT 2.505000 1.950000 4.685000 2.020000 ;
        RECT 2.505000 2.020000 3.785000 2.120000 ;
        RECT 2.505000 2.120000 2.755000 2.735000 ;
        RECT 2.665000 1.010000 4.180000 1.180000 ;
        RECT 2.665000 1.180000 2.835000 1.820000 ;
        RECT 3.455000 2.120000 3.785000 2.980000 ;
        RECT 3.615000 1.850000 4.685000 1.950000 ;
        RECT 3.850000 0.610000 4.180000 1.010000 ;
        RECT 4.355000 2.020000 4.685000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 1.010000 ;
      RECT 0.115000  1.010000 2.445000 1.180000 ;
      RECT 0.120000  1.950000 2.250000 2.120000 ;
      RECT 0.120000  2.120000 0.370000 2.980000 ;
      RECT 0.570000  2.290000 0.820000 3.245000 ;
      RECT 0.615000  0.085000 0.945000 0.825000 ;
      RECT 1.020000  2.120000 1.350000 2.980000 ;
      RECT 1.115000  0.350000 1.445000 1.010000 ;
      RECT 1.550000  2.290000 1.720000 2.905000 ;
      RECT 1.550000  2.905000 3.285000 3.075000 ;
      RECT 1.615000  0.085000 1.945000 0.825000 ;
      RECT 1.920000  2.120000 2.250000 2.735000 ;
      RECT 2.115000  0.350000 2.445000 0.670000 ;
      RECT 2.115000  0.670000 3.670000 0.840000 ;
      RECT 2.115000  0.840000 2.445000 1.010000 ;
      RECT 2.625000  0.085000 3.240000 0.500000 ;
      RECT 2.955000  2.290000 3.285000 2.905000 ;
      RECT 3.420000  0.255000 4.680000 0.425000 ;
      RECT 3.420000  0.425000 3.670000 0.670000 ;
      RECT 3.985000  2.190000 4.155000 3.245000 ;
      RECT 4.350000  0.425000 4.680000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_ms__o31ai_2

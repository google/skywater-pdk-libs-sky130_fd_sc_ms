* NGSPICE file created from sky130_fd_sc_ms__ha_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__ha_1 A B VGND VNB VPB VPWR COUT SUM
M1000 VPWR A a_239_294# VPB pshort w=840000u l=180000u
+  ad=1.6456e+12p pd=9.84e+06u as=2.268e+11p ps=2.22e+06u
M1001 a_695_119# B a_239_294# VNB nlowvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=1.824e+11p ps=1.85e+06u
M1002 VPWR A a_389_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.9e+11p ps=2.78e+06u
M1003 a_389_392# B a_83_260# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.13e+11p ps=2.65e+06u
M1004 COUT a_239_294# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=6.95225e+11p ps=6.36e+06u
M1005 VPWR a_83_260# SUM VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1006 a_83_260# a_239_294# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_305_130# a_239_294# a_83_260# VNB nlowvt w=640000u l=150000u
+  ad=3.616e+11p pd=3.69e+06u as=1.726e+11p ps=1.85e+06u
M1008 COUT a_239_294# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1009 VGND B a_305_130# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A a_695_119# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_83_260# SUM VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1012 a_239_294# B VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_305_130# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


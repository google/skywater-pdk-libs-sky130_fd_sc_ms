* File: sky130_fd_sc_ms__or3_2.spice
* Created: Fri Aug 28 18:07:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__or3_2.pex.spice"
.subckt sky130_fd_sc_ms__or3_2  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_C_M1009_g N_A_27_74#_M1009_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1616 AS=0.1824 PD=1.145 PS=1.85 NRD=20.616 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.6 A=0.096 P=1.58 MULT=1
MM1008 N_A_27_74#_M1008_d N_B_M1008_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.1616 PD=0.99 PS=1.145 NRD=0 NRS=21.552 M=1 R=4.26667 SA=75000.9
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1005 N_VGND_M1005_d N_A_M1005_g N_A_27_74#_M1008_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.179293 AS=0.112 PD=1.21043 PS=0.99 NRD=19.68 NRS=13.116 M=1 R=4.26667
+ SA=75001.4 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1005_d N_A_27_74#_M1000_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.207307 AS=0.1036 PD=1.39957 PS=1.02 NRD=29.184 NRS=0 M=1 R=4.93333
+ SA=75001.8 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_27_74#_M1007_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1003 A_153_392# N_C_M1003_g N_A_27_74#_M1003_s VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.28 PD=1.24 PS=2.56 NRD=12.7853 NRS=0 M=1 R=5.55556 SA=90000.2 SB=90002.3
+ A=0.18 P=2.36 MULT=1
MM1002 A_237_392# N_B_M1002_g A_153_392# VPB PSHORT L=0.18 W=1 AD=0.195 AS=0.12
+ PD=1.39 PS=1.24 NRD=27.5603 NRS=12.7853 M=1 R=5.55556 SA=90000.6 SB=90001.9
+ A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g A_237_392# VPB PSHORT L=0.18 W=1 AD=0.216981
+ AS=0.195 PD=1.46226 PS=1.39 NRD=0 NRS=27.5603 M=1 R=5.55556 SA=90001.2
+ SB=90001.3 A=0.18 P=2.36 MULT=1
MM1004 N_X_M1004_d N_A_27_74#_M1004_g N_VPWR_M1001_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.243019 PD=1.39 PS=1.63774 NRD=0 NRS=27.2451 M=1 R=6.22222
+ SA=90001.6 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1006 N_X_M1004_d N_A_27_74#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__or3_2.pxi.spice"
*
.ends
*
*

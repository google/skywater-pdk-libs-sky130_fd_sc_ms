* File: sky130_fd_sc_ms__dfbbp_1.pex.spice
* Created: Wed Sep  2 12:02:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DFBBP_1%CLK 3 6 8 11 13
r37 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=1.385
+ $X2=0.52 $Y2=1.55
r38 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=1.385
+ $X2=0.52 $Y2=1.22
r39 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.52
+ $Y=1.385 $X2=0.52 $Y2=1.385
r40 8 12 6.22942 $w=3.68e-07 $l=2e-07 $layer=LI1_cond $X=0.72 $Y=1.365 $X2=0.52
+ $Y2=1.365
r41 6 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.595 $Y=2.4
+ $X2=0.595 $Y2=1.55
r42 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=0.74
+ $X2=0.495 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBP_1%D 3 7 9 13
r35 11 13 18 $w=2.41e-07 $l=9e-08 $layer=POLY_cond $X=2.035 $Y=1.99 $X2=2.125
+ $Y2=1.99
r36 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.125
+ $Y=1.99 $X2=2.125 $Y2=1.99
r37 5 13 79 $w=2.41e-07 $l=4.70319e-07 $layer=POLY_cond $X=2.52 $Y=2.155
+ $X2=2.125 $Y2=1.99
r38 5 7 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=2.52 $Y=2.155 $X2=2.52
+ $Y2=2.525
r39 1 11 13.8727 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.035 $Y=1.825
+ $X2=2.035 $Y2=1.99
r40 1 3 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=2.035 $Y=1.825
+ $X2=2.035 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBP_1%A_671_93# 1 2 7 9 12 16 18 20 22 25 26 28 29
+ 32 34 35 36 37 41 45 47 52
c156 37 0 9.9441e-20 $X=5.335 $Y=0.925
c157 29 0 5.24889e-20 $X=3.72 $Y=0.815
c158 25 0 1.13254e-19 $X=3.59 $Y=1.29
c159 7 0 1.68855e-19 $X=3.43 $Y=1.125
r160 46 55 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.015 $Y=1.42
+ $X2=6.015 $Y2=1.585
r161 46 52 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=6.015 $Y=1.42
+ $X2=6.015 $Y2=1.295
r162 45 48 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.015 $Y=1.42
+ $X2=6.015 $Y2=1.585
r163 45 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.015 $Y=1.42
+ $X2=6.015 $Y2=1.255
r164 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.015
+ $Y=1.42 $X2=6.015 $Y2=1.42
r165 41 48 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.935 $Y=1.825
+ $X2=5.935 $Y2=1.585
r166 38 47 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.935 $Y=1.01
+ $X2=5.935 $Y2=1.255
r167 37 43 9.11221 $w=3.9e-07 $l=2.17991e-07 $layer=LI1_cond $X=5.335 $Y=0.925
+ $X2=5.17 $Y2=0.802
r168 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.85 $Y=0.925
+ $X2=5.935 $Y2=1.01
r169 36 37 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=5.85 $Y=0.925
+ $X2=5.335 $Y2=0.925
r170 34 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.85 $Y=1.91
+ $X2=5.935 $Y2=1.825
r171 34 35 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=5.85 $Y=1.91 $X2=4.95
+ $Y2=1.91
r172 30 35 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.825 $Y=1.995
+ $X2=4.95 $Y2=1.91
r173 30 32 2.0744 $w=2.48e-07 $l=4.5e-08 $layer=LI1_cond $X=4.825 $Y=1.995
+ $X2=4.825 $Y2=2.04
r174 28 43 8.79939 $w=3.9e-07 $l=1.61369e-07 $layer=LI1_cond $X=5.015 $Y=0.815
+ $X2=5.17 $Y2=0.802
r175 28 29 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=5.015 $Y=0.815
+ $X2=3.72 $Y2=0.815
r176 26 49 28.8839 $w=2.67e-07 $l=1.6e-07 $layer=POLY_cond $X=3.59 $Y=1.29
+ $X2=3.43 $Y2=1.29
r177 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.59
+ $Y=1.29 $X2=3.59 $Y2=1.29
r178 23 29 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=3.592 $Y=0.9
+ $X2=3.72 $Y2=0.815
r179 23 25 17.6256 $w=2.53e-07 $l=3.9e-07 $layer=LI1_cond $X=3.592 $Y=0.9
+ $X2=3.592 $Y2=1.29
r180 20 22 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.515 $Y=1.22
+ $X2=6.515 $Y2=0.87
r181 19 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.18 $Y=1.295
+ $X2=6.015 $Y2=1.295
r182 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.44 $Y=1.295
+ $X2=6.515 $Y2=1.22
r183 18 19 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=6.44 $Y=1.295
+ $X2=6.18 $Y2=1.295
r184 16 55 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=5.94 $Y=2.315
+ $X2=5.94 $Y2=1.585
r185 10 26 52.3521 $w=2.67e-07 $l=3.63249e-07 $layer=POLY_cond $X=3.88 $Y=1.455
+ $X2=3.59 $Y2=1.29
r186 10 12 252.661 $w=1.8e-07 $l=6.5e-07 $layer=POLY_cond $X=3.88 $Y=1.455
+ $X2=3.88 $Y2=2.105
r187 7 49 16.2448 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.125
+ $X2=3.43 $Y2=1.29
r188 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.43 $Y=1.125
+ $X2=3.43 $Y2=0.805
r189 2 32 300 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_PDIFF $count=2 $X=4.56
+ $Y=1.895 $X2=4.785 $Y2=2.04
r190 1 43 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=5.03
+ $Y=0.595 $X2=5.17 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBP_1%SET_B 3 7 11 15 18 19 20 22 23 24 26 27 28
+ 30 31 32 37 39 44 47
c163 47 0 1.01328e-19 $X=8.405 $Y=1.635
r164 47 50 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.405 $Y=1.635
+ $X2=8.405 $Y2=1.8
r165 47 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.405 $Y=1.635
+ $X2=8.405 $Y2=1.47
r166 39 53 7.33544 $w=3.16e-07 $l=1.9e-07 $layer=LI1_cond $X=8.405 $Y=1.635
+ $X2=8.405 $Y2=1.825
r167 39 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.405
+ $Y=1.635 $X2=8.405 $Y2=1.635
r168 35 44 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.395 $Y=1.53
+ $X2=4.47 $Y2=1.53
r169 35 41 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=4.395 $Y=1.53
+ $X2=4.285 $Y2=1.53
r170 34 37 2.35192 $w=2.43e-07 $l=5e-08 $layer=LI1_cond $X=4.395 $Y=1.532
+ $X2=4.445 $Y2=1.532
r171 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.395
+ $Y=1.53 $X2=4.395 $Y2=1.53
r172 31 53 4.36715 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.24 $Y=1.825
+ $X2=8.405 $Y2=1.825
r173 31 32 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=8.24 $Y=1.825
+ $X2=7.45 $Y2=1.825
r174 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.365 $Y=1.91
+ $X2=7.45 $Y2=1.825
r175 29 30 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=7.365 $Y=1.91
+ $X2=7.365 $Y2=2.905
r176 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.28 $Y=2.99
+ $X2=7.365 $Y2=2.905
r177 27 28 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=7.28 $Y=2.99
+ $X2=6.21 $Y2=2.99
r178 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.125 $Y=2.905
+ $X2=6.21 $Y2=2.99
r179 25 26 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=6.125 $Y=2.335
+ $X2=6.125 $Y2=2.905
r180 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.04 $Y=2.25
+ $X2=6.125 $Y2=2.335
r181 23 24 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=6.04 $Y=2.25
+ $X2=5.33 $Y2=2.25
r182 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.245 $Y=2.335
+ $X2=5.33 $Y2=2.25
r183 21 22 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.245 $Y=2.335
+ $X2=5.245 $Y2=2.905
r184 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.16 $Y=2.99
+ $X2=5.245 $Y2=2.905
r185 19 20 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=5.16 $Y=2.99
+ $X2=4.53 $Y2=2.99
r186 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.445 $Y=2.905
+ $X2=4.53 $Y2=2.99
r187 17 37 2.87745 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=4.445 $Y=1.655
+ $X2=4.445 $Y2=1.532
r188 17 18 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=4.445 $Y=1.655
+ $X2=4.445 $Y2=2.905
r189 15 50 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=8.48 $Y=2.46
+ $X2=8.48 $Y2=1.8
r190 11 49 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=8.465 $Y=0.74
+ $X2=8.465 $Y2=1.47
r191 5 44 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.47 $Y=1.695
+ $X2=4.47 $Y2=1.53
r192 5 7 241 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=4.47 $Y=1.695 $X2=4.47
+ $Y2=2.315
r193 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.285 $Y=1.365
+ $X2=4.285 $Y2=1.53
r194 1 3 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=4.285 $Y=1.365
+ $X2=4.285 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBP_1%A_520_87# 1 2 9 12 14 19 22 24 27 28 29 30
+ 34 36
c102 34 0 9.9441e-20 $X=4.935 $Y=1.42
c103 29 0 1.68855e-19 $X=4.06 $Y=1.155
r104 34 37 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.935 $Y=1.42
+ $X2=4.935 $Y2=1.585
r105 34 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.935 $Y=1.42
+ $X2=4.935 $Y2=1.255
r106 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.935
+ $Y=1.42 $X2=4.935 $Y2=1.42
r107 28 33 11.2257 $w=2.88e-07 $l=3.42243e-07 $layer=LI1_cond $X=4.745 $Y=1.155
+ $X2=4.922 $Y2=1.42
r108 28 29 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=4.745 $Y=1.155
+ $X2=4.06 $Y2=1.155
r109 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.975 $Y=1.24
+ $X2=4.06 $Y2=1.155
r110 26 27 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.975 $Y=1.24
+ $X2=3.975 $Y2=1.625
r111 25 30 2.57001 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.43 $Y=1.71
+ $X2=3.277 $Y2=1.71
r112 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.89 $Y=1.71
+ $X2=3.975 $Y2=1.625
r113 24 25 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.89 $Y=1.71
+ $X2=3.43 $Y2=1.71
r114 20 30 3.87901 $w=2.37e-07 $l=8.5e-08 $layer=LI1_cond $X=3.277 $Y=1.795
+ $X2=3.277 $Y2=1.71
r115 20 22 14.1694 $w=3.03e-07 $l=3.75e-07 $layer=LI1_cond $X=3.277 $Y=1.795
+ $X2=3.277 $Y2=2.17
r116 19 30 3.87901 $w=2.37e-07 $l=1.13666e-07 $layer=LI1_cond $X=3.21 $Y=1.625
+ $X2=3.277 $Y2=1.71
r117 18 19 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=3.21 $Y=0.745
+ $X2=3.21 $Y2=1.625
r118 14 18 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.125 $Y=0.58
+ $X2=3.21 $Y2=0.745
r119 14 16 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=3.125 $Y=0.58
+ $X2=2.74 $Y2=0.58
r120 12 37 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=5.01 $Y=2.315
+ $X2=5.01 $Y2=1.585
r121 9 36 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=4.955 $Y=0.87
+ $X2=4.955 $Y2=1.255
r122 2 22 600 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=1 $X=3.06
+ $Y=2.315 $X2=3.265 $Y2=2.17
r123 1 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.6
+ $Y=0.435 $X2=2.74 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBP_1%A_1062_93# 1 2 9 12 16 18 20 21 23 27 31 33
+ 38 40 41 44 47 48 51 53 55 63
c145 55 0 9.47353e-20 $X=9.875 $Y=1.295
r146 51 54 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.475 $Y=1.42
+ $X2=5.475 $Y2=1.585
r147 51 53 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.475 $Y=1.42
+ $X2=5.475 $Y2=1.255
r148 48 63 6.55126 $w=3.53e-07 $l=1.05e-07 $layer=LI1_cond $X=9.887 $Y=1.295
+ $X2=9.887 $Y2=1.19
r149 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=1.295
+ $X2=9.84 $Y2=1.295
r150 44 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.475
+ $Y=1.42 $X2=5.475 $Y2=1.42
r151 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.295
+ $X2=5.52 $Y2=1.295
r152 41 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=1.295
+ $X2=5.52 $Y2=1.295
r153 40 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.695 $Y=1.295
+ $X2=9.84 $Y2=1.295
r154 40 41 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=9.695 $Y=1.295
+ $X2=5.665 $Y2=1.295
r155 35 38 6.24041 $w=4.58e-07 $l=2.4e-07 $layer=LI1_cond $X=9.98 $Y=0.58
+ $X2=10.22 $Y2=0.58
r156 31 33 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=10.065 $Y=1.945
+ $X2=10.24 $Y2=1.945
r157 29 35 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=9.98 $Y=0.81 $X2=9.98
+ $Y2=0.58
r158 29 63 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.98 $Y=0.81
+ $X2=9.98 $Y2=1.19
r159 28 55 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.875 $Y=1.385
+ $X2=9.875 $Y2=1.295
r160 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.875
+ $Y=1.385 $X2=9.875 $Y2=1.385
r161 25 31 7.08698 $w=2.5e-07 $l=2.32237e-07 $layer=LI1_cond $X=9.887 $Y=1.82
+ $X2=10.065 $Y2=1.945
r162 25 27 14.1215 $w=3.53e-07 $l=4.35e-07 $layer=LI1_cond $X=9.887 $Y=1.82
+ $X2=9.887 $Y2=1.385
r163 24 48 2.33735 $w=3.53e-07 $l=7.2e-08 $layer=LI1_cond $X=9.887 $Y=1.367
+ $X2=9.887 $Y2=1.295
r164 24 27 0.584337 $w=3.53e-07 $l=1.8e-08 $layer=LI1_cond $X=9.887 $Y=1.367
+ $X2=9.887 $Y2=1.385
r165 22 23 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.5 $Y=1.295 $X2=9.41
+ $Y2=1.295
r166 21 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.71 $Y=1.295
+ $X2=9.875 $Y2=1.295
r167 21 22 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=9.71 $Y=1.295
+ $X2=9.5 $Y2=1.295
r168 18 23 18.8402 $w=1.65e-07 $l=7.98436e-08 $layer=POLY_cond $X=9.4 $Y=1.22
+ $X2=9.41 $Y2=1.295
r169 18 20 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.4 $Y=1.22 $X2=9.4
+ $Y2=0.74
r170 14 23 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=9.41 $Y=1.37
+ $X2=9.41 $Y2=1.295
r171 14 16 423.694 $w=1.8e-07 $l=1.09e-06 $layer=POLY_cond $X=9.41 $Y=1.37
+ $X2=9.41 $Y2=2.46
r172 12 54 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=5.43 $Y=2.315
+ $X2=5.43 $Y2=1.585
r173 9 53 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=5.385 $Y=0.87
+ $X2=5.385 $Y2=1.255
r174 2 33 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=10.115
+ $Y=1.84 $X2=10.24 $Y2=1.985
r175 1 38 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=10.075
+ $Y=0.37 $X2=10.22 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBP_1%A_27_74# 1 2 9 13 15 18 19 20 22 23 24 27 31
+ 33 38 41 43 45 48 51 54 58 62 67 68 71 72 74 75 77 78 79 85 91
c219 71 0 1.41865e-20 $X=7.505 $Y=1.065
c220 31 0 1.13254e-19 $X=3.49 $Y=2.105
c221 27 0 1.57784e-19 $X=2.525 $Y=0.645
c222 18 0 9.68576e-20 $X=1.525 $Y=1.3
c223 13 0 7.43587e-20 $X=1.175 $Y=2.4
c224 9 0 6.93165e-20 $X=0.995 $Y=0.74
r225 84 85 33.0969 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.175 $Y=1.465
+ $X2=1.265 $Y2=1.465
r226 78 86 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=6.605 $Y=1.775
+ $X2=6.48 $Y2=1.775
r227 77 79 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.605 $Y=1.775
+ $X2=6.605 $Y2=1.61
r228 77 78 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.605
+ $Y=1.775 $X2=6.605 $Y2=1.775
r229 72 91 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.505 $Y=1.065
+ $X2=7.505 $Y2=0.9
r230 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.505
+ $Y=1.065 $X2=7.505 $Y2=1.065
r231 69 71 22.6943 $w=3.23e-07 $l=6.4e-07 $layer=LI1_cond $X=7.507 $Y=0.425
+ $X2=7.507 $Y2=1.065
r232 67 69 7.72402 $w=1.7e-07 $l=2.00035e-07 $layer=LI1_cond $X=7.345 $Y=0.34
+ $X2=7.507 $Y2=0.425
r233 67 68 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=7.345 $Y=0.34
+ $X2=6.77 $Y2=0.34
r234 65 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.685 $Y=0.425
+ $X2=6.77 $Y2=0.34
r235 65 79 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=6.685 $Y=0.425
+ $X2=6.685 $Y2=1.61
r236 63 84 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=1.06 $Y=1.465
+ $X2=1.175 $Y2=1.465
r237 63 81 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=1.06 $Y=1.465
+ $X2=0.995 $Y2=1.465
r238 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.06
+ $Y=1.465 $X2=1.06 $Y2=1.465
r239 60 62 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.06 $Y=1.72
+ $X2=1.06 $Y2=1.465
r240 59 75 3.57226 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.535 $Y=1.805
+ $X2=0.31 $Y2=1.805
r241 58 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.975 $Y=1.805
+ $X2=1.06 $Y2=1.72
r242 58 59 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=0.975 $Y=1.805
+ $X2=0.535 $Y2=1.805
r243 54 56 22.061 $w=4.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.31 $Y=1.985
+ $X2=0.31 $Y2=2.815
r244 52 75 3.05675 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.31 $Y=1.89
+ $X2=0.31 $Y2=1.805
r245 52 54 2.52505 $w=4.48e-07 $l=9.5e-08 $layer=LI1_cond $X=0.31 $Y=1.89
+ $X2=0.31 $Y2=1.985
r246 51 75 3.05675 $w=3.1e-07 $l=1.77482e-07 $layer=LI1_cond $X=0.17 $Y=1.72
+ $X2=0.31 $Y2=1.805
r247 51 74 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.17 $Y=1.72
+ $X2=0.17 $Y2=1.01
r248 46 74 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.265 $Y=0.83
+ $X2=0.265 $Y2=1.01
r249 46 48 10.0839 $w=3.58e-07 $l=3.15e-07 $layer=LI1_cond $X=0.265 $Y=0.83
+ $X2=0.265 $Y2=0.515
r250 42 43 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.525 $Y=1.375
+ $X2=1.675 $Y2=1.375
r251 41 91 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.415 $Y=0.58
+ $X2=7.415 $Y2=0.9
r252 36 38 207.96 $w=1.8e-07 $l=5.35e-07 $layer=POLY_cond $X=6.48 $Y=3.075
+ $X2=6.48 $Y2=2.54
r253 35 86 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.48 $Y=1.94
+ $X2=6.48 $Y2=1.775
r254 35 38 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=6.48 $Y=1.94 $X2=6.48
+ $Y2=2.54
r255 34 45 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.58 $Y=3.15 $X2=3.49
+ $Y2=3.15
r256 33 36 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.39 $Y=3.15
+ $X2=6.48 $Y2=3.075
r257 33 34 1440.87 $w=1.5e-07 $l=2.81e-06 $layer=POLY_cond $X=6.39 $Y=3.15
+ $X2=3.58 $Y2=3.15
r258 29 45 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.49 $Y=3.075
+ $X2=3.49 $Y2=3.15
r259 29 31 377.048 $w=1.8e-07 $l=9.7e-07 $layer=POLY_cond $X=3.49 $Y=3.075
+ $X2=3.49 $Y2=2.105
r260 25 27 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.525 $Y=0.255
+ $X2=2.525 $Y2=0.645
r261 23 45 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.4 $Y=3.15 $X2=3.49
+ $Y2=3.15
r262 23 24 846.064 $w=1.5e-07 $l=1.65e-06 $layer=POLY_cond $X=3.4 $Y=3.15
+ $X2=1.75 $Y2=3.15
r263 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.675 $Y=3.075
+ $X2=1.75 $Y2=3.15
r264 21 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.675 $Y=1.45
+ $X2=1.675 $Y2=1.375
r265 21 22 833.245 $w=1.5e-07 $l=1.625e-06 $layer=POLY_cond $X=1.675 $Y=1.45
+ $X2=1.675 $Y2=3.075
r266 19 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.45 $Y=0.18
+ $X2=2.525 $Y2=0.255
r267 19 20 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=2.45 $Y=0.18
+ $X2=1.6 $Y2=0.18
r268 18 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.525 $Y=1.3
+ $X2=1.525 $Y2=1.375
r269 17 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.525 $Y=0.255
+ $X2=1.6 $Y2=0.18
r270 17 18 535.84 $w=1.5e-07 $l=1.045e-06 $layer=POLY_cond $X=1.525 $Y=0.255
+ $X2=1.525 $Y2=1.3
r271 15 42 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.45 $Y=1.375
+ $X2=1.525 $Y2=1.375
r272 15 85 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=1.45 $Y=1.375
+ $X2=1.265 $Y2=1.375
r273 11 84 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.175 $Y=1.63
+ $X2=1.175 $Y2=1.465
r274 11 13 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.175 $Y=1.63
+ $X2=1.175 $Y2=2.4
r275 7 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.3
+ $X2=0.995 $Y2=1.465
r276 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.995 $Y=1.3
+ $X2=0.995 $Y2=0.74
r277 2 56 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.225
+ $Y=1.84 $X2=0.37 $Y2=2.815
r278 2 54 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.225
+ $Y=1.84 $X2=0.37 $Y2=1.985
r279 1 48 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBP_1%A_214_74# 1 2 7 12 15 17 18 22 25 29 32 34
+ 35 38 40 42 48 52
c137 48 0 1.57784e-19 $X=2.485 $Y=1.42
c138 32 0 1.41865e-20 $X=7.055 $Y=1.295
c139 12 0 5.24889e-20 $X=2.955 $Y=0.645
r140 49 52 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.485 $Y=1.42
+ $X2=2.485 $Y2=1.33
r141 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.485
+ $Y=1.42 $X2=2.485 $Y2=1.42
r142 46 48 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=1.565 $Y=1.42
+ $X2=2.485 $Y2=1.42
r143 42 44 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=1.44 $Y=1.985
+ $X2=1.44 $Y2=2.815
r144 40 46 7.64946 $w=2.65e-07 $l=2.07123e-07 $layer=LI1_cond $X=1.44 $Y=1.585
+ $X2=1.345 $Y2=1.42
r145 40 42 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=1.44 $Y=1.585
+ $X2=1.44 $Y2=1.985
r146 36 46 16.8014 $w=3.6e-07 $l=4.89592e-07 $layer=LI1_cond $X=1.305 $Y=0.95
+ $X2=1.345 $Y2=1.42
r147 36 38 13.9254 $w=3.58e-07 $l=4.35e-07 $layer=LI1_cond $X=1.305 $Y=0.95
+ $X2=1.305 $Y2=0.515
r148 34 35 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=7.027 $Y=2.18
+ $X2=7.027 $Y2=2.33
r149 30 32 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.875 $Y=1.295
+ $X2=7.055 $Y2=1.295
r150 27 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.055 $Y=1.37
+ $X2=7.055 $Y2=1.295
r151 27 34 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=7.055 $Y=1.37
+ $X2=7.055 $Y2=2.18
r152 25 35 163.258 $w=1.8e-07 $l=4.2e-07 $layer=POLY_cond $X=7.015 $Y=2.75
+ $X2=7.015 $Y2=2.33
r153 20 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.875 $Y=1.22
+ $X2=6.875 $Y2=1.295
r154 20 22 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.875 $Y=1.22
+ $X2=6.875 $Y2=0.87
r155 19 22 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=6.875 $Y=0.255
+ $X2=6.875 $Y2=0.87
r156 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.8 $Y=0.18
+ $X2=6.875 $Y2=0.255
r157 17 18 1933.13 $w=1.5e-07 $l=3.77e-06 $layer=POLY_cond $X=6.8 $Y=0.18
+ $X2=3.03 $Y2=0.18
r158 13 29 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=2.97 $Y=1.405
+ $X2=2.97 $Y2=1.33
r159 13 15 435.355 $w=1.8e-07 $l=1.12e-06 $layer=POLY_cond $X=2.97 $Y=1.405
+ $X2=2.97 $Y2=2.525
r160 10 29 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=2.955 $Y=1.255
+ $X2=2.97 $Y2=1.33
r161 10 12 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.955 $Y=1.255
+ $X2=2.955 $Y2=0.645
r162 9 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.955 $Y=0.255
+ $X2=3.03 $Y2=0.18
r163 9 12 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.955 $Y=0.255
+ $X2=2.955 $Y2=0.645
r164 8 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.65 $Y=1.33
+ $X2=2.485 $Y2=1.33
r165 7 29 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.88 $Y=1.33 $X2=2.97
+ $Y2=1.33
r166 7 8 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.88 $Y=1.33 $X2=2.65
+ $Y2=1.33
r167 2 44 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.265
+ $Y=1.84 $X2=1.4 $Y2=2.815
r168 2 42 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.265
+ $Y=1.84 $X2=1.4 $Y2=1.985
r169 1 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.21 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBP_1%A_1474_446# 1 2 9 12 15 19 23 25 28 30 31 33
+ 34 36 39 43 45 53 57 60 61 64 67 70 74 79 80
c180 64 0 1.25678e-19 $X=10.865 $Y=2.24
c181 53 0 4.99671e-20 $X=7.785 $Y=2.215
c182 39 0 1.35822e-19 $X=7.955 $Y=1.81
c183 12 0 2.35385e-20 $X=7.875 $Y=2.05
r184 79 80 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.955
+ $Y=1.485 $X2=10.955 $Y2=1.485
r185 76 79 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=10.865 $Y=1.485
+ $X2=10.955 $Y2=1.485
r186 72 74 3.63098 $w=3.63e-07 $l=1.15e-07 $layer=LI1_cond $X=9.185 $Y=0.777
+ $X2=9.3 $Y2=0.777
r187 69 70 6.73996 $w=4.38e-07 $l=8.5e-08 $layer=LI1_cond $X=9.3 $Y=2.19
+ $X2=9.385 $Y2=2.19
r188 68 69 12.834 $w=4.38e-07 $l=4.9e-07 $layer=LI1_cond $X=8.81 $Y=2.19 $X2=9.3
+ $Y2=2.19
r189 66 68 1.04768 $w=4.38e-07 $l=4e-08 $layer=LI1_cond $X=8.77 $Y=2.19 $X2=8.81
+ $Y2=2.19
r190 66 67 3.40064 $w=4.38e-07 $l=8.5e-08 $layer=LI1_cond $X=8.77 $Y=2.19
+ $X2=8.685 $Y2=2.19
r191 63 76 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.865 $Y=1.65
+ $X2=10.865 $Y2=1.485
r192 63 64 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=10.865 $Y=1.65
+ $X2=10.865 $Y2=2.24
r193 61 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.78 $Y=2.325
+ $X2=10.865 $Y2=2.24
r194 61 70 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=10.78 $Y=2.325
+ $X2=9.385 $Y2=2.325
r195 60 69 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=9.3 $Y=1.97 $X2=9.3
+ $Y2=2.19
r196 59 74 5.2253 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=9.3 $Y=0.96 $X2=9.3
+ $Y2=0.777
r197 59 60 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=9.3 $Y=0.96
+ $X2=9.3 $Y2=1.97
r198 55 68 4.04531 $w=2.5e-07 $l=2.2e-07 $layer=LI1_cond $X=8.81 $Y=2.41
+ $X2=8.81 $Y2=2.19
r199 55 57 2.99635 $w=2.48e-07 $l=6.5e-08 $layer=LI1_cond $X=8.81 $Y=2.41
+ $X2=8.81 $Y2=2.475
r200 53 84 17.2143 $w=2.52e-07 $l=9e-08 $layer=POLY_cond $X=7.785 $Y=2.215
+ $X2=7.875 $Y2=2.215
r201 52 67 34.5733 $w=2.98e-07 $l=9e-07 $layer=LI1_cond $X=7.785 $Y=2.23
+ $X2=8.685 $Y2=2.23
r202 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.785
+ $Y=2.215 $X2=7.785 $Y2=2.215
r203 41 43 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=11.71 $Y=0.94
+ $X2=12.005 $Y2=0.94
r204 37 39 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=7.875 $Y=1.81
+ $X2=7.955 $Y2=1.81
r205 34 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.005 $Y=0.865
+ $X2=12.005 $Y2=0.94
r206 34 36 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=12.005 $Y=0.865
+ $X2=12.005 $Y2=0.58
r207 31 46 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=11.95 $Y=1.9
+ $X2=11.71 $Y2=1.9
r208 31 33 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=11.95 $Y=1.975
+ $X2=11.95 $Y2=2.47
r209 30 46 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.71 $Y=1.825
+ $X2=11.71 $Y2=1.9
r210 29 45 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.71 $Y=1.65
+ $X2=11.71 $Y2=1.485
r211 29 30 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=11.71 $Y=1.65
+ $X2=11.71 $Y2=1.825
r212 28 45 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.71 $Y=1.32
+ $X2=11.71 $Y2=1.485
r213 27 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.71 $Y=1.015
+ $X2=11.71 $Y2=0.94
r214 27 28 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=11.71 $Y=1.015
+ $X2=11.71 $Y2=1.32
r215 26 80 3.90195 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=11.09 $Y=1.485
+ $X2=10.94 $Y2=1.485
r216 25 45 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=11.635 $Y=1.485
+ $X2=11.71 $Y2=1.485
r217 25 26 95.2994 $w=3.3e-07 $l=5.45e-07 $layer=POLY_cond $X=11.635 $Y=1.485
+ $X2=11.09 $Y2=1.485
r218 21 80 34.7346 $w=1.65e-07 $l=1.98997e-07 $layer=POLY_cond $X=11.015 $Y=1.32
+ $X2=10.94 $Y2=1.485
r219 21 23 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=11.015 $Y=1.32
+ $X2=11.015 $Y2=0.74
r220 17 80 34.7346 $w=1.65e-07 $l=1.83916e-07 $layer=POLY_cond $X=10.98 $Y=1.65
+ $X2=10.94 $Y2=1.485
r221 17 19 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=10.98 $Y=1.65
+ $X2=10.98 $Y2=2.4
r222 13 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.955 $Y=1.735
+ $X2=7.955 $Y2=1.81
r223 13 15 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=7.955 $Y=1.735
+ $X2=7.955 $Y2=0.58
r224 12 84 14.904 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.875 $Y=2.05
+ $X2=7.875 $Y2=2.215
r225 11 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.875 $Y=1.885
+ $X2=7.875 $Y2=1.81
r226 11 12 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.875 $Y=1.885
+ $X2=7.875 $Y2=2.05
r227 7 53 62.1627 $w=2.52e-07 $l=3.99061e-07 $layer=POLY_cond $X=7.46 $Y=2.38
+ $X2=7.785 $Y2=2.215
r228 7 9 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=7.46 $Y=2.38 $X2=7.46
+ $Y2=2.75
r229 2 66 600 $w=1.7e-07 $l=2.73861e-07 $layer=licon1_PDIFF $count=1 $X=8.57
+ $Y=1.96 $X2=8.77 $Y2=2.135
r230 2 57 300 $w=1.7e-07 $l=6.06815e-07 $layer=licon1_PDIFF $count=2 $X=8.57
+ $Y=1.96 $X2=8.77 $Y2=2.475
r231 1 72 182 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_NDIFF $count=1 $X=9.04
+ $Y=0.37 $X2=9.185 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBP_1%A_1314_424# 1 2 9 12 16 20 23 24 26 31 33 34
+ 42 45
c104 31 0 4.99671e-20 $X=7.025 $Y=2.195
c105 26 0 1.01328e-19 $X=8.78 $Y=1.215
c106 23 0 1.59361e-19 $X=7.025 $Y=2.11
r107 42 46 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.945 $Y=1.385
+ $X2=8.945 $Y2=1.55
r108 42 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.945 $Y=1.385
+ $X2=8.945 $Y2=1.22
r109 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.945
+ $Y=1.385 $X2=8.945 $Y2=1.385
r110 34 36 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.985 $Y=1.215
+ $X2=7.985 $Y2=1.485
r111 29 31 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.705 $Y=2.195
+ $X2=7.025 $Y2=2.195
r112 27 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.07 $Y=1.215
+ $X2=7.985 $Y2=1.215
r113 26 41 7.39303 $w=2.63e-07 $l=1.7e-07 $layer=LI1_cond $X=8.912 $Y=1.215
+ $X2=8.912 $Y2=1.385
r114 26 27 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=8.78 $Y=1.215
+ $X2=8.07 $Y2=1.215
r115 25 33 1.97946 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=7.175 $Y=1.485
+ $X2=7.057 $Y2=1.485
r116 24 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=1.485
+ $X2=7.985 $Y2=1.485
r117 24 25 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=7.9 $Y=1.485
+ $X2=7.175 $Y2=1.485
r118 23 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.025 $Y=2.11
+ $X2=7.025 $Y2=2.195
r119 22 33 4.45556 $w=2.02e-07 $l=9.97246e-08 $layer=LI1_cond $X=7.025 $Y=1.57
+ $X2=7.057 $Y2=1.485
r120 22 23 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=7.025 $Y=1.57
+ $X2=7.025 $Y2=2.11
r121 18 33 4.45556 $w=2.02e-07 $l=8.5e-08 $layer=LI1_cond $X=7.057 $Y=1.4
+ $X2=7.057 $Y2=1.485
r122 18 20 31.3857 $w=2.33e-07 $l=6.4e-07 $layer=LI1_cond $X=7.057 $Y=1.4
+ $X2=7.057 $Y2=0.76
r123 16 29 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.705 $Y=2.65
+ $X2=6.705 $Y2=2.28
r124 12 46 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=8.995 $Y=2.46
+ $X2=8.995 $Y2=1.55
r125 9 45 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.965 $Y=0.74
+ $X2=8.965 $Y2=1.22
r126 2 29 600 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=1 $X=6.57
+ $Y=2.12 $X2=6.705 $Y2=2.27
r127 2 16 600 $w=1.7e-07 $l=5.93675e-07 $layer=licon1_PDIFF $count=1 $X=6.57
+ $Y=2.12 $X2=6.705 $Y2=2.65
r128 1 20 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=6.95
+ $Y=0.595 $X2=7.09 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBP_1%RESET_B 3 7 11 12 13 16 17
c46 16 0 1.55842e-19 $X=10.415 $Y=1.145
r47 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.415
+ $Y=1.145 $X2=10.415 $Y2=1.145
r48 13 17 1.69593 $w=6.68e-07 $l=9.5e-08 $layer=LI1_cond $X=10.32 $Y=1.315
+ $X2=10.415 $Y2=1.315
r49 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=10.415 $Y=1.485
+ $X2=10.415 $Y2=1.145
r50 11 12 37.7308 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.415 $Y=1.485
+ $X2=10.415 $Y2=1.65
r51 10 16 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.415 $Y=0.98
+ $X2=10.415 $Y2=1.145
r52 7 12 198.242 $w=1.8e-07 $l=5.1e-07 $layer=POLY_cond $X=10.465 $Y=2.16
+ $X2=10.465 $Y2=1.65
r53 3 10 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=10.435 $Y=0.58
+ $X2=10.435 $Y2=0.98
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBP_1%A_2320_410# 1 2 9 13 15 16 19 23 25 29 32 33
c61 15 0 1.21275e-19 $X=12.375 $Y=1.42
r62 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.19
+ $Y=1.42 $X2=12.19 $Y2=1.42
r63 27 32 0.341012 $w=3.3e-07 $l=1.18e-07 $layer=LI1_cond $X=11.875 $Y=1.42
+ $X2=11.757 $Y2=1.42
r64 27 29 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=11.875 $Y=1.42
+ $X2=12.19 $Y2=1.42
r65 23 33 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=11.765 $Y=2.155
+ $X2=11.765 $Y2=2.03
r66 23 25 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=11.765 $Y=2.155
+ $X2=11.765 $Y2=2.195
r67 21 32 7.59124 $w=2.02e-07 $l=1.80291e-07 $layer=LI1_cond $X=11.725 $Y=1.585
+ $X2=11.757 $Y2=1.42
r68 21 33 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=11.725 $Y=1.585
+ $X2=11.725 $Y2=2.03
r69 17 32 7.59124 $w=2.02e-07 $l=1.65e-07 $layer=LI1_cond $X=11.757 $Y=1.255
+ $X2=11.757 $Y2=1.42
r70 17 19 33.1021 $w=2.33e-07 $l=6.75e-07 $layer=LI1_cond $X=11.757 $Y=1.255
+ $X2=11.757 $Y2=0.58
r71 15 30 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=12.375 $Y=1.42
+ $X2=12.19 $Y2=1.42
r72 15 16 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=12.375 $Y=1.42
+ $X2=12.465 $Y2=1.42
r73 11 16 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=12.48 $Y=1.255
+ $X2=12.465 $Y2=1.42
r74 11 13 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=12.48 $Y=1.255
+ $X2=12.48 $Y2=0.74
r75 7 16 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=12.465 $Y=1.585
+ $X2=12.465 $Y2=1.42
r76 7 9 316.798 $w=1.8e-07 $l=8.15e-07 $layer=POLY_cond $X=12.465 $Y=1.585
+ $X2=12.465 $Y2=2.4
r77 2 25 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=11.6
+ $Y=2.05 $X2=11.725 $Y2=2.195
r78 1 19 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=11.645
+ $Y=0.37 $X2=11.79 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBP_1%VPWR 1 2 3 4 5 6 7 8 29 35 39 43 47 51 55 60
+ 61 62 64 69 77 94 98 105 106 109 112 115 118 123 129 131 134
c146 35 0 7.43587e-20 $X=2.29 $Y=2.59
r147 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r148 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r149 127 129 8.95 $w=7.63e-07 $l=2e-08 $layer=LI1_cond $X=8.4 $Y=3.032 $X2=8.42
+ $Y2=3.032
r150 127 128 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r151 125 127 2.26708 $w=7.63e-07 $l=1.45e-07 $layer=LI1_cond $X=8.255 $Y=3.032
+ $X2=8.4 $Y2=3.032
r152 122 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r153 121 125 5.23773 $w=7.63e-07 $l=3.35e-07 $layer=LI1_cond $X=7.92 $Y=3.032
+ $X2=8.255 $Y2=3.032
r154 121 123 13.3278 $w=7.63e-07 $l=3e-07 $layer=LI1_cond $X=7.92 $Y=3.032
+ $X2=7.62 $Y2=3.032
r155 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r156 118 119 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r157 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r158 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r159 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r160 106 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=12.24 $Y2=3.33
r161 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r162 103 134 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.325 $Y=3.33
+ $X2=12.2 $Y2=3.33
r163 103 105 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=12.325 $Y=3.33
+ $X2=12.72 $Y2=3.33
r164 102 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r165 102 132 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=10.8 $Y2=3.33
r166 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r167 99 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.92 $Y=3.33
+ $X2=10.755 $Y2=3.33
r168 99 101 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=10.92 $Y=3.33
+ $X2=11.76 $Y2=3.33
r169 98 134 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.075 $Y=3.33
+ $X2=12.2 $Y2=3.33
r170 98 101 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.075 $Y=3.33
+ $X2=11.76 $Y2=3.33
r171 97 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r172 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r173 94 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.59 $Y=3.33
+ $X2=10.755 $Y2=3.33
r174 94 96 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=10.59 $Y=3.33
+ $X2=10.32 $Y2=3.33
r175 93 97 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r176 93 128 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.4 $Y2=3.33
r177 92 129 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=9.36 $Y=3.33
+ $X2=8.42 $Y2=3.33
r178 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r179 89 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r180 88 123 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.44 $Y=3.33
+ $X2=7.62 $Y2=3.33
r181 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r182 86 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r183 85 88 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=7.44
+ $Y2=3.33
r184 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r185 83 118 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.87 $Y=3.33
+ $X2=5.685 $Y2=3.33
r186 83 85 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=5.87 $Y=3.33 $X2=6
+ $Y2=3.33
r187 81 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r188 81 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r189 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r190 78 115 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.19 $Y=3.33
+ $X2=4.065 $Y2=3.33
r191 78 80 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.19 $Y=3.33
+ $X2=4.56 $Y2=3.33
r192 77 118 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.5 $Y=3.33
+ $X2=5.685 $Y2=3.33
r193 77 80 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=5.5 $Y=3.33
+ $X2=4.56 $Y2=3.33
r194 76 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r195 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r196 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r197 73 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r198 72 75 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r199 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r200 70 112 12.6176 $w=1.7e-07 $l=3.03e-07 $layer=LI1_cond $X=2.41 $Y=3.33
+ $X2=2.107 $Y2=3.33
r201 70 72 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.41 $Y=3.33
+ $X2=2.64 $Y2=3.33
r202 69 115 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.94 $Y=3.33
+ $X2=4.065 $Y2=3.33
r203 69 75 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.94 $Y=3.33
+ $X2=3.6 $Y2=3.33
r204 68 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r205 68 110 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r206 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r207 65 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=0.87 $Y2=3.33
r208 65 67 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.035 $Y=3.33
+ $X2=1.68 $Y2=3.33
r209 64 112 12.6176 $w=1.7e-07 $l=3.02e-07 $layer=LI1_cond $X=1.805 $Y=3.33
+ $X2=2.107 $Y2=3.33
r210 64 67 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.805 $Y=3.33
+ $X2=1.68 $Y2=3.33
r211 62 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r212 62 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r213 60 92 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=9.47 $Y=3.33
+ $X2=9.36 $Y2=3.33
r214 60 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.47 $Y=3.33
+ $X2=9.635 $Y2=3.33
r215 59 96 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=9.8 $Y=3.33
+ $X2=10.32 $Y2=3.33
r216 59 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.8 $Y=3.33
+ $X2=9.635 $Y2=3.33
r217 55 58 19.1306 $w=2.48e-07 $l=4.15e-07 $layer=LI1_cond $X=12.2 $Y=1.985
+ $X2=12.2 $Y2=2.4
r218 53 134 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.2 $Y=3.245
+ $X2=12.2 $Y2=3.33
r219 53 58 38.9526 $w=2.48e-07 $l=8.45e-07 $layer=LI1_cond $X=12.2 $Y=3.245
+ $X2=12.2 $Y2=2.4
r220 49 131 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.755 $Y=3.245
+ $X2=10.755 $Y2=3.33
r221 49 51 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=10.755 $Y=3.245
+ $X2=10.755 $Y2=2.745
r222 45 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.635 $Y=3.245
+ $X2=9.635 $Y2=3.33
r223 45 47 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=9.635 $Y=3.245
+ $X2=9.635 $Y2=2.78
r224 41 118 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.685 $Y=3.245
+ $X2=5.685 $Y2=3.33
r225 41 43 20.4014 $w=3.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.685 $Y=3.245
+ $X2=5.685 $Y2=2.59
r226 37 115 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.065 $Y=3.245
+ $X2=4.065 $Y2=3.33
r227 37 39 50.477 $w=2.48e-07 $l=1.095e-06 $layer=LI1_cond $X=4.065 $Y=3.245
+ $X2=4.065 $Y2=2.15
r228 33 112 2.53987 $w=6.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.107 $Y=3.245
+ $X2=2.107 $Y2=3.33
r229 33 35 12.9493 $w=6.03e-07 $l=6.55e-07 $layer=LI1_cond $X=2.107 $Y=3.245
+ $X2=2.107 $Y2=2.59
r230 29 32 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.87 $Y=2.145
+ $X2=0.87 $Y2=2.825
r231 27 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=3.245
+ $X2=0.87 $Y2=3.33
r232 27 32 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=0.87 $Y=3.245
+ $X2=0.87 $Y2=2.825
r233 8 58 300 $w=1.7e-07 $l=4.38748e-07 $layer=licon1_PDIFF $count=2 $X=12.04
+ $Y=2.05 $X2=12.24 $Y2=2.4
r234 8 55 600 $w=1.7e-07 $l=2.30217e-07 $layer=licon1_PDIFF $count=1 $X=12.04
+ $Y=2.05 $X2=12.24 $Y2=1.985
r235 7 51 600 $w=1.7e-07 $l=1.00001e-06 $layer=licon1_PDIFF $count=1 $X=10.555
+ $Y=1.84 $X2=10.755 $Y2=2.745
r236 6 47 600 $w=1.7e-07 $l=8.84929e-07 $layer=licon1_PDIFF $count=1 $X=9.5
+ $Y=1.96 $X2=9.635 $Y2=2.78
r237 5 125 300 $w=1.7e-07 $l=8.31204e-07 $layer=licon1_PDIFF $count=2 $X=7.55
+ $Y=2.54 $X2=8.255 $Y2=2.815
r238 4 43 600 $w=1.7e-07 $l=7.73111e-07 $layer=licon1_PDIFF $count=1 $X=5.52
+ $Y=1.895 $X2=5.685 $Y2=2.59
r239 3 39 600 $w=1.7e-07 $l=3.15357e-07 $layer=licon1_PDIFF $count=1 $X=3.97
+ $Y=1.895 $X2=4.105 $Y2=2.15
r240 2 35 300 $w=1.7e-07 $l=5.866e-07 $layer=licon1_PDIFF $count=2 $X=1.825
+ $Y=2.315 $X2=2.29 $Y2=2.59
r241 1 32 400 $w=1.7e-07 $l=1.07352e-06 $layer=licon1_PDIFF $count=1 $X=0.685
+ $Y=1.84 $X2=0.87 $Y2=2.825
r242 1 29 400 $w=1.7e-07 $l=3.86588e-07 $layer=licon1_PDIFF $count=1 $X=0.685
+ $Y=1.84 $X2=0.87 $Y2=2.145
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBP_1%A_422_125# 1 2 9 11 12 16 17
c45 12 0 9.68576e-20 $X=2.335 $Y=1
r46 16 17 10.552 $w=3.73e-07 $l=2.3e-07 $layer=LI1_cond $X=2.767 $Y=2.525
+ $X2=2.767 $Y2=2.295
r47 13 17 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=2.87 $Y=1.085
+ $X2=2.87 $Y2=2.295
r48 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.785 $Y=1
+ $X2=2.87 $Y2=1.085
r49 11 12 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.785 $Y=1 $X2=2.335
+ $Y2=1
r50 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.21 $Y=0.915
+ $X2=2.335 $Y2=1
r51 7 9 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=2.21 $Y=0.915 $X2=2.21
+ $Y2=0.835
r52 2 16 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=2.61
+ $Y=2.315 $X2=2.745 $Y2=2.525
r53 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.11
+ $Y=0.625 $X2=2.25 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBP_1%Q_N 1 2 9 13 14 15 16 23 32
c37 32 0 1.21275e-19 $X=11.29 $Y=1.82
c38 13 0 1.55842e-19 $X=11.262 $Y=1.13
r39 21 23 1.52529 $w=3.38e-07 $l=4.5e-08 $layer=LI1_cond $X=11.29 $Y=1.99
+ $X2=11.29 $Y2=2.035
r40 15 16 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=11.29 $Y=2.405
+ $X2=11.29 $Y2=2.775
r41 14 21 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=11.29 $Y=1.97
+ $X2=11.29 $Y2=1.99
r42 14 32 7.96349 $w=3.38e-07 $l=1.5e-07 $layer=LI1_cond $X=11.29 $Y=1.97
+ $X2=11.29 $Y2=1.82
r43 14 15 11.8634 $w=3.38e-07 $l=3.5e-07 $layer=LI1_cond $X=11.29 $Y=2.055
+ $X2=11.29 $Y2=2.405
r44 14 23 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=11.29 $Y=2.055
+ $X2=11.29 $Y2=2.035
r45 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=11.375 $Y=1.13
+ $X2=11.375 $Y2=1.82
r46 7 13 9.56083 $w=3.93e-07 $l=1.97e-07 $layer=LI1_cond $X=11.262 $Y=0.933
+ $X2=11.262 $Y2=1.13
r47 7 9 12.1955 $w=3.93e-07 $l=4.18e-07 $layer=LI1_cond $X=11.262 $Y=0.933
+ $X2=11.262 $Y2=0.515
r48 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=11.07
+ $Y=1.84 $X2=11.205 $Y2=1.985
r49 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=11.07
+ $Y=1.84 $X2=11.205 $Y2=2.815
r50 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.09
+ $Y=0.37 $X2=11.23 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBP_1%Q 1 2 7 8 9 10 11 12 13
r14 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=12.692 $Y=2.405
+ $X2=12.692 $Y2=2.775
r15 11 12 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=12.692 $Y=1.985
+ $X2=12.692 $Y2=2.405
r16 10 11 11.0084 $w=3.33e-07 $l=3.2e-07 $layer=LI1_cond $X=12.692 $Y=1.665
+ $X2=12.692 $Y2=1.985
r17 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=12.692 $Y=1.295
+ $X2=12.692 $Y2=1.665
r18 8 9 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=12.692 $Y=0.925
+ $X2=12.692 $Y2=1.295
r19 7 8 14.1045 $w=3.33e-07 $l=4.1e-07 $layer=LI1_cond $X=12.692 $Y=0.515
+ $X2=12.692 $Y2=0.925
r20 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=12.555
+ $Y=1.84 $X2=12.69 $Y2=2.815
r21 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=12.555
+ $Y=1.84 $X2=12.69 $Y2=1.985
r22 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.555
+ $Y=0.37 $X2=12.695 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBP_1%VGND 1 2 3 4 5 6 7 24 26 30 33 36 40 44 48
+ 51 52 54 57 58 59 61 66 75 82 92 93 96 99 111 114
c159 30 0 6.93165e-20 $X=1.82 $Y=0.835
r160 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r161 111 112 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r162 104 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0
+ $X2=4.08 $Y2=0
r163 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r164 97 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=1.68 $Y2=0
r165 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r166 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r167 90 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.72 $Y2=0
r168 90 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=10.8 $Y2=0
r169 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r170 87 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.895 $Y=0
+ $X2=10.73 $Y2=0
r171 87 89 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=10.895 $Y=0
+ $X2=11.76 $Y2=0
r172 86 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r173 86 112 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=8.4 $Y2=0
r174 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r175 83 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.415 $Y=0
+ $X2=8.25 $Y2=0
r176 83 85 124.283 $w=1.68e-07 $l=1.905e-06 $layer=LI1_cond $X=8.415 $Y=0
+ $X2=10.32 $Y2=0
r177 82 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.565 $Y=0
+ $X2=10.73 $Y2=0
r178 82 85 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=10.565 $Y=0
+ $X2=10.32 $Y2=0
r179 81 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r180 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r181 77 80 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.48 $Y=0 $X2=7.92
+ $Y2=0
r182 75 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.085 $Y=0
+ $X2=8.25 $Y2=0
r183 75 80 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=8.085 $Y=0
+ $X2=7.92 $Y2=0
r184 74 106 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6 $Y=0 $X2=4.08
+ $Y2=0
r185 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r186 71 73 120.369 $w=1.68e-07 $l=1.845e-06 $layer=LI1_cond $X=4.155 $Y=0 $X2=6
+ $Y2=0
r187 70 104 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=3.6 $Y2=0
r188 70 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r189 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r190 67 99 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.905 $Y=0 $X2=1.78
+ $Y2=0
r191 67 69 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.905 $Y=0
+ $X2=2.16 $Y2=0
r192 66 108 9.54852 $w=5.93e-07 $l=4.75e-07 $layer=LI1_cond $X=3.857 $Y=0
+ $X2=3.857 $Y2=0.475
r193 66 71 8.26286 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=3.857 $Y=0
+ $X2=4.155 $Y2=0
r194 66 106 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r195 66 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r196 66 69 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=3.56 $Y=0 $X2=2.16
+ $Y2=0
r197 64 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r198 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r199 61 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r200 61 63 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r201 59 81 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=7.92 $Y2=0
r202 59 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r203 59 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r204 57 89 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.055 $Y=0
+ $X2=11.76 $Y2=0
r205 57 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.055 $Y=0
+ $X2=12.18 $Y2=0
r206 56 92 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=12.305 $Y=0
+ $X2=12.72 $Y2=0
r207 56 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.305 $Y=0
+ $X2=12.18 $Y2=0
r208 54 55 6.55957 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.245 $Y=0.505
+ $X2=6.245 $Y2=0.67
r209 51 73 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=6.06 $Y=0 $X2=6 $Y2=0
r210 51 52 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.06 $Y=0 $X2=6.245
+ $Y2=0
r211 50 77 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=6.43 $Y=0 $X2=6.48
+ $Y2=0
r212 50 52 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.43 $Y=0 $X2=6.245
+ $Y2=0
r213 46 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.18 $Y=0.085
+ $X2=12.18 $Y2=0
r214 46 48 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=12.18 $Y=0.085
+ $X2=12.18 $Y2=0.58
r215 42 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.73 $Y=0.085
+ $X2=10.73 $Y2=0
r216 42 44 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.73 $Y=0.085
+ $X2=10.73 $Y2=0.58
r217 38 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.25 $Y=0.085
+ $X2=8.25 $Y2=0
r218 38 40 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=8.25 $Y=0.085
+ $X2=8.25 $Y2=0.495
r219 36 55 12.0046 $w=2.38e-07 $l=2.5e-07 $layer=LI1_cond $X=6.31 $Y=0.92
+ $X2=6.31 $Y2=0.67
r220 33 54 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=6.245 $Y=0.485
+ $X2=6.245 $Y2=0.505
r221 32 52 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.245 $Y=0.085
+ $X2=6.245 $Y2=0
r222 32 33 12.4588 $w=3.68e-07 $l=4e-07 $layer=LI1_cond $X=6.245 $Y=0.085
+ $X2=6.245 $Y2=0.485
r223 28 99 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0
r224 28 30 34.5733 $w=2.48e-07 $l=7.5e-07 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0.835
r225 27 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r226 26 99 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.655 $Y=0 $X2=1.78
+ $Y2=0
r227 26 27 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.655 $Y=0
+ $X2=0.945 $Y2=0
r228 22 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r229 22 24 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.515
r230 7 48 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.08
+ $Y=0.37 $X2=12.22 $Y2=0.58
r231 6 44 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=10.51
+ $Y=0.37 $X2=10.73 $Y2=0.58
r232 5 40 91 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=2 $X=8.03
+ $Y=0.37 $X2=8.25 $Y2=0.495
r233 4 54 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.085
+ $Y=0.36 $X2=6.225 $Y2=0.505
r234 4 36 182 $w=1.7e-07 $l=6.58787e-07 $layer=licon1_NDIFF $count=1 $X=6.085
+ $Y=0.36 $X2=6.3 $Y2=0.92
r235 3 108 182 $w=1.7e-07 $l=4.05586e-07 $layer=licon1_NDIFF $count=1 $X=3.505
+ $Y=0.595 $X2=3.855 $Y2=0.475
r236 2 30 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.675
+ $Y=0.625 $X2=1.82 $Y2=0.835
r237 1 24 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBP_1%A_872_119# 1 2 7 9 14
r27 14 17 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=5.675 $Y=0.34
+ $X2=5.675 $Y2=0.5
r28 9 12 3.79463 $w=4.08e-07 $l=1.35e-07 $layer=LI1_cond $X=4.62 $Y=0.34
+ $X2=4.62 $Y2=0.475
r29 8 9 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=4.825 $Y=0.34 $X2=4.62
+ $Y2=0.34
r30 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.51 $Y=0.34
+ $X2=5.675 $Y2=0.34
r31 7 8 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=5.51 $Y=0.34
+ $X2=4.825 $Y2=0.34
r32 2 17 182 $w=1.7e-07 $l=2.58167e-07 $layer=licon1_NDIFF $count=1 $X=5.46
+ $Y=0.595 $X2=5.675 $Y2=0.5
r33 1 12 182 $w=1.7e-07 $l=3.14325e-07 $layer=licon1_NDIFF $count=1 $X=4.36
+ $Y=0.595 $X2=4.62 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_MS__DFBBP_1%A_1708_74# 1 2 9 11 12 15
c29 15 0 9.47353e-20 $X=9.64 $Y=0.515
r30 13 15 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=9.64 $Y=0.425 $X2=9.64
+ $Y2=0.515
r31 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.555 $Y=0.34
+ $X2=9.64 $Y2=0.425
r32 11 12 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=9.555 $Y=0.34
+ $X2=8.915 $Y2=0.34
r33 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.75 $Y=0.425
+ $X2=8.915 $Y2=0.34
r34 7 9 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=8.75 $Y=0.425 $X2=8.75
+ $Y2=0.495
r35 2 15 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=9.475
+ $Y=0.37 $X2=9.64 $Y2=0.515
r36 1 9 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=8.54
+ $Y=0.37 $X2=8.75 $Y2=0.495
.ends


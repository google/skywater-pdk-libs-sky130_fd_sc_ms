* File: sky130_fd_sc_ms__o41a_2.pex.spice
* Created: Wed Sep  2 12:26:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O41A_2%A1 3 7 9 12 13
r29 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.43 $Y=1.515
+ $X2=0.43 $Y2=1.68
r30 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.43 $Y=1.515
+ $X2=0.43 $Y2=1.35
r31 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.43
+ $Y=1.515 $X2=0.43 $Y2=1.515
r32 9 13 5.09219 $w=4.28e-07 $l=1.9e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.43 $Y2=1.565
r33 7 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=0.74
+ $X2=0.495 $Y2=1.35
r34 3 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.505 $Y=2.4
+ $X2=0.505 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_2%A2 3 7 11 12 14 15 16
c42 12 0 1.89954e-19 $X=1 $Y=1.515
r43 15 16 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.075 $Y=2.405
+ $X2=1.075 $Y2=2.775
r44 15 23 6.10498 $w=4.78e-07 $l=2.45e-07 $layer=LI1_cond $X=1.075 $Y=2.405
+ $X2=1.075 $Y2=2.16
r45 14 23 3.11479 $w=4.78e-07 $l=1.25e-07 $layer=LI1_cond $X=1.075 $Y=2.035
+ $X2=1.075 $Y2=2.16
r46 14 30 4.04332 $w=4.78e-07 $l=1.15e-07 $layer=LI1_cond $X=1.075 $Y=2.035
+ $X2=1.075 $Y2=1.92
r47 12 22 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.515 $X2=1
+ $Y2=1.68
r48 12 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.515 $X2=1
+ $Y2=1.35
r49 11 30 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=1 $Y=1.515 $X2=1
+ $Y2=1.92
r50 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.515
+ $X2=1 $Y2=1.515
r51 7 21 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.065 $Y=0.74
+ $X2=1.065 $Y2=1.35
r52 3 22 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.925 $Y=2.4
+ $X2=0.925 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_2%A3 3 7 9 10 11 12 19
c41 3 0 2.29616e-19 $X=1.495 $Y=2.4
r42 19 22 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.57 $Y=1.515
+ $X2=1.57 $Y2=1.68
r43 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.57 $Y=1.515
+ $X2=1.57 $Y2=1.35
r44 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.57
+ $Y=1.515 $X2=1.57 $Y2=1.515
r45 11 12 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=2.405
+ $X2=1.68 $Y2=2.775
r46 10 11 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=2.035
+ $X2=1.68 $Y2=2.405
r47 9 23 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=1.515
+ $X2=1.68 $Y2=1.68
r48 9 20 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=1.68 $Y=1.515
+ $X2=1.57 $Y2=1.515
r49 9 10 16.034 $w=2.28e-07 $l=3.2e-07 $layer=LI1_cond $X=1.68 $Y=1.715 $X2=1.68
+ $Y2=2.035
r50 9 23 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=1.68 $Y=1.715
+ $X2=1.68 $Y2=1.68
r51 7 21 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.495 $Y=0.74
+ $X2=1.495 $Y2=1.35
r52 3 22 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.495 $Y=2.4
+ $X2=1.495 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_2%A4 3 7 9 12 13
c35 13 0 9.34971e-20 $X=2.14 $Y=1.515
r36 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.14 $Y=1.515
+ $X2=2.14 $Y2=1.68
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.14 $Y=1.515
+ $X2=2.14 $Y2=1.35
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.515 $X2=2.14 $Y2=1.515
r39 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.14 $Y=1.665
+ $X2=2.14 $Y2=1.515
r40 7 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.23 $Y=0.74 $X2=2.23
+ $Y2=1.35
r41 3 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.065 $Y=2.4
+ $X2=2.065 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_2%B1 3 7 9 10 14
c41 14 0 8.8899e-20 $X=2.71 $Y=1.515
r42 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.515
+ $X2=2.71 $Y2=1.68
r43 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.515
+ $X2=2.71 $Y2=1.35
r44 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.71
+ $Y=1.515 $X2=2.71 $Y2=1.515
r45 10 15 10.9884 $w=4.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=2.71 $Y2=1.565
r46 9 15 1.87607 $w=4.28e-07 $l=7e-08 $layer=LI1_cond $X=2.64 $Y=1.565 $X2=2.71
+ $Y2=1.565
r47 7 16 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.675 $Y=0.74
+ $X2=2.675 $Y2=1.35
r48 3 17 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.635 $Y=2.34
+ $X2=2.635 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_2%A_431_368# 1 2 9 13 17 21 23 25 27 31 33 34
+ 36 38 46
c81 38 0 8.8899e-20 $X=3.57 $Y=1.465
c82 23 0 1.36119e-19 $X=2.29 $Y=2.12
r83 46 47 9.1519 $w=3.16e-07 $l=6e-08 $layer=POLY_cond $X=4.235 $Y=1.465
+ $X2=4.295 $Y2=1.465
r84 45 46 59.4873 $w=3.16e-07 $l=3.9e-07 $layer=POLY_cond $X=3.845 $Y=1.465
+ $X2=4.235 $Y2=1.465
r85 44 45 6.10127 $w=3.16e-07 $l=4e-08 $layer=POLY_cond $X=3.805 $Y=1.465
+ $X2=3.845 $Y2=1.465
r86 39 44 35.8449 $w=3.16e-07 $l=2.35e-07 $layer=POLY_cond $X=3.57 $Y=1.465
+ $X2=3.805 $Y2=1.465
r87 38 42 14.8553 $w=3.3e-07 $l=3.7e-07 $layer=LI1_cond $X=3.57 $Y=1.465
+ $X2=3.57 $Y2=1.095
r88 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.465 $X2=3.57 $Y2=1.465
r89 36 38 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=3.57 $Y=1.95
+ $X2=3.57 $Y2=1.465
r90 33 42 2.45823 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=1.095
+ $X2=3.57 $Y2=1.095
r91 33 34 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.405 $Y=1.095
+ $X2=3.125 $Y2=1.095
r92 29 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.96 $Y=1.01
+ $X2=3.125 $Y2=1.095
r93 29 31 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.96 $Y=1.01
+ $X2=2.96 $Y2=0.515
r94 28 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.455 $Y=2.035
+ $X2=2.29 $Y2=2.035
r95 27 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.405 $Y=2.035
+ $X2=3.57 $Y2=1.95
r96 27 28 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=3.405 $Y=2.035
+ $X2=2.455 $Y2=2.035
r97 23 41 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=2.12 $X2=2.29
+ $Y2=2.035
r98 23 25 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.29 $Y=2.12
+ $X2=2.29 $Y2=2.815
r99 19 47 15.9236 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.295 $Y=1.63
+ $X2=4.295 $Y2=1.465
r100 19 21 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.295 $Y=1.63
+ $X2=4.295 $Y2=2.4
r101 15 46 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.235 $Y=1.3
+ $X2=4.235 $Y2=1.465
r102 15 17 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.235 $Y=1.3
+ $X2=4.235 $Y2=0.74
r103 11 45 15.9236 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.845 $Y=1.63
+ $X2=3.845 $Y2=1.465
r104 11 13 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=3.845 $Y=1.63
+ $X2=3.845 $Y2=2.4
r105 7 44 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.805 $Y=1.3
+ $X2=3.805 $Y2=1.465
r106 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.805 $Y=1.3
+ $X2=3.805 $Y2=0.74
r107 2 41 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=2.155
+ $Y=1.84 $X2=2.29 $Y2=2.115
r108 2 25 600 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.155
+ $Y=1.84 $X2=2.29 $Y2=2.815
r109 1 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.75
+ $Y=0.37 $X2=2.89 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_2%VPWR 1 2 3 10 12 16 18 22 24 32 41 50
r49 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r50 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 36 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r52 36 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r53 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r54 33 35 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.78 $Y=3.33 $X2=4.08
+ $Y2=3.33
r55 32 49 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=4.355 $Y=3.33
+ $X2=4.577 $Y2=3.33
r56 32 35 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.355 $Y=3.33
+ $X2=4.08 $Y2=3.33
r57 31 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r58 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r60 27 30 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 25 38 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r63 25 27 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 24 33 12.2881 $w=1.7e-07 $l=5.43e-07 $layer=LI1_cond $X=3.237 $Y=3.33
+ $X2=3.78 $Y2=3.33
r65 24 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r66 24 41 10.7382 $w=1.083e-06 $l=9.55e-07 $layer=LI1_cond $X=3.237 $Y=3.33
+ $X2=3.237 $Y2=2.375
r67 24 30 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.695 $Y=3.33
+ $X2=2.64 $Y2=3.33
r68 22 31 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r69 22 28 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=0.72 $Y2=3.33
r70 18 21 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.52 $Y=1.985
+ $X2=4.52 $Y2=2.815
r71 16 49 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.52 $Y=3.245
+ $X2=4.577 $Y2=3.33
r72 16 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.52 $Y=3.245
+ $X2=4.52 $Y2=2.815
r73 12 15 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.28 $Y=2.115 $X2=0.28
+ $Y2=2.815
r74 10 38 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r75 10 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r76 3 21 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.385
+ $Y=1.84 $X2=4.52 $Y2=2.815
r77 3 18 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.385
+ $Y=1.84 $X2=4.52 $Y2=1.985
r78 2 41 300 $w=1.7e-07 $l=1.12617e-06 $layer=licon1_PDIFF $count=2 $X=2.725
+ $Y=1.84 $X2=3.615 $Y2=2.375
r79 2 41 150 $w=1.7e-07 $l=7.40523e-07 $layer=licon1_PDIFF $count=4 $X=2.725
+ $Y=1.84 $X2=3.215 $Y2=2.375
r80 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r81 1 12 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_2%X 1 2 9 11 13 17
r23 13 15 44.9047 $w=2.03e-07 $l=8.3e-07 $layer=LI1_cond $X=4.052 $Y=1.985
+ $X2=4.052 $Y2=2.815
r24 11 17 5.91863 $w=2.75e-07 $l=1.27789e-07 $layer=LI1_cond $X=4.052 $Y=1.41
+ $X2=4.025 $Y2=1.295
r25 11 13 31.1086 $w=2.03e-07 $l=5.75e-07 $layer=LI1_cond $X=4.052 $Y=1.41
+ $X2=4.052 $Y2=1.985
r26 7 17 12.5749 $w=3.3e-07 $l=3.32491e-07 $layer=LI1_cond $X=4.02 $Y=0.965
+ $X2=4.025 $Y2=1.295
r27 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.02 $Y=0.965 $X2=4.02
+ $Y2=0.515
r28 2 15 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.935
+ $Y=1.84 $X2=4.07 $Y2=2.815
r29 2 13 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.935
+ $Y=1.84 $X2=4.07 $Y2=1.985
r30 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.88
+ $Y=0.37 $X2=4.02 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_2%A_27_74# 1 2 3 12 14 15 18 20 24 26
c53 26 0 1.89954e-19 $X=1.28 $Y=1.095
r54 22 24 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.46 $Y=1.01
+ $X2=2.46 $Y2=0.515
r55 21 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=1.095
+ $X2=1.28 $Y2=1.095
r56 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.295 $Y=1.095
+ $X2=2.46 $Y2=1.01
r57 20 21 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=2.295 $Y=1.095
+ $X2=1.445 $Y2=1.095
r58 16 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=1.01 $X2=1.28
+ $Y2=1.095
r59 16 18 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.28 $Y=1.01
+ $X2=1.28 $Y2=0.515
r60 14 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=1.095
+ $X2=1.28 $Y2=1.095
r61 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=1.095
+ $X2=0.445 $Y2=1.095
r62 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.445 $Y2=1.095
r63 10 12 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.28 $Y2=0.515
r64 3 24 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=2.305
+ $Y=0.37 $X2=2.46 $Y2=0.515
r65 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.14
+ $Y=0.37 $X2=1.28 $Y2=0.515
r66 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_2%VGND 1 2 3 4 15 17 21 25 27 29 31 33 38 46 52
+ 55 58 62
r61 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r62 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r63 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r64 53 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r65 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r66 50 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r67 50 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r68 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r69 47 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.52
+ $Y2=0
r70 47 49 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.685 $Y=0 $X2=4.08
+ $Y2=0
r71 46 61 4.01281 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.577
+ $Y2=0
r72 46 49 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.08
+ $Y2=0
r73 45 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r74 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r75 42 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r76 41 44 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r77 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r78 39 55 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=1.87
+ $Y2=0
r79 39 41 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.125 $Y=0 $X2=2.16
+ $Y2=0
r80 38 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.355 $Y=0 $X2=3.52
+ $Y2=0
r81 38 44 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.355 $Y=0 $X2=3.12
+ $Y2=0
r82 36 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r83 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r84 33 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r85 33 35 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r86 31 45 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r87 31 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r88 27 61 3.19941 $w=2.6e-07 $l=1.27609e-07 $layer=LI1_cond $X=4.485 $Y=0.085
+ $X2=4.577 $Y2=0
r89 27 29 18.1731 $w=2.58e-07 $l=4.1e-07 $layer=LI1_cond $X=4.485 $Y=0.085
+ $X2=4.485 $Y2=0.495
r90 23 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.52 $Y=0.085
+ $X2=3.52 $Y2=0
r91 23 25 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=3.52 $Y=0.085
+ $X2=3.52 $Y2=0.655
r92 19 55 2.12513 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.87 $Y=0.085
+ $X2=1.87 $Y2=0
r93 19 21 12.4298 $w=5.08e-07 $l=5.3e-07 $layer=LI1_cond $X=1.87 $Y=0.085
+ $X2=1.87 $Y2=0.615
r94 18 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r95 17 55 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.615 $Y=0 $X2=1.87
+ $Y2=0
r96 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=0 $X2=0.945
+ $Y2=0
r97 13 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r98 13 15 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.595
r99 4 29 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.31
+ $Y=0.37 $X2=4.45 $Y2=0.495
r100 3 25 182 $w=1.7e-07 $l=3.77492e-07 $layer=licon1_NDIFF $count=1 $X=3.375
+ $Y=0.37 $X2=3.59 $Y2=0.655
r101 2 21 182 $w=1.7e-07 $l=4.04351e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.37 $X2=1.87 $Y2=0.615
r102 1 15 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.595
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__and4b_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__and4b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.233700 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.300000 0.455000 1.780000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.350000 3.405000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.505000 1.350000 2.835000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 1.350000 2.295000 1.780000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055000 0.350000 1.385000 1.130000 ;
        RECT 1.055000 1.130000 1.225000 1.820000 ;
        RECT 1.055000 1.820000 1.440000 2.200000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.320000 0.085000 ;
        RECT 0.625000  0.085000 0.875000 0.790000 ;
        RECT 1.555000  0.085000 2.165000 0.790000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 4.320000 3.415000 ;
        RECT 0.650000 2.710000 0.980000 3.245000 ;
        RECT 1.645000 2.710000 1.975000 3.245000 ;
        RECT 2.740000 2.710000 3.070000 3.245000 ;
        RECT 3.850000 2.710000 4.205000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 0.540000 0.445000 0.960000 ;
      RECT 0.115000 0.960000 0.795000 1.130000 ;
      RECT 0.115000 1.950000 0.795000 2.370000 ;
      RECT 0.115000 2.370000 3.985000 2.540000 ;
      RECT 0.115000 2.540000 0.445000 2.700000 ;
      RECT 0.625000 1.130000 0.795000 1.950000 ;
      RECT 1.395000 1.300000 1.780000 1.630000 ;
      RECT 1.610000 0.960000 4.070000 1.130000 ;
      RECT 1.610000 1.130000 1.780000 1.300000 ;
      RECT 1.610000 1.630000 1.780000 1.950000 ;
      RECT 1.610000 1.950000 3.645000 2.200000 ;
      RECT 3.615000 1.350000 3.985000 1.680000 ;
      RECT 3.740000 0.350000 4.070000 0.960000 ;
      RECT 3.815000 1.680000 3.985000 2.370000 ;
  END
END sky130_fd_sc_ms__and4b_2

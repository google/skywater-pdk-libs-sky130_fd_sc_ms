* File: sky130_fd_sc_ms__fa_1.spice
* Created: Wed Sep  2 12:09:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__fa_1.pex.spice"
.subckt sky130_fd_sc_ms__fa_1  VNB VPB A CIN B SUM VPWR COUT VGND
* 
* VGND	VGND
* COUT	COUT
* VPWR	VPWR
* SUM	SUM
* B	B
* CIN	CIN
* A	A
* VPB	VPB
* VNB	VNB
MM1026 N_VGND_M1026_d N_A_69_260#_M1026_g N_SUM_M1026_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.205457 AS=0.2109 PD=1.49609 PS=2.05 NRD=36.096 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75006 A=0.111 P=1.78 MULT=1
MM1011 A_237_75# N_A_M1011_g N_VGND_M1026_d VNB NLOWVT L=0.15 W=0.64 AD=0.0768
+ AS=0.177693 PD=0.88 PS=1.29391 NRD=12.18 NRS=18.744 M=1 R=4.26667 SA=75000.8
+ SB=75006.3 A=0.096 P=1.58 MULT=1
MM1000 A_315_75# N_B_M1000_g A_237_75# VNB NLOWVT L=0.15 W=0.64 AD=0.0768
+ AS=0.0768 PD=0.88 PS=0.88 NRD=12.18 NRS=12.18 M=1 R=4.26667 SA=75001.2
+ SB=75005.9 A=0.096 P=1.58 MULT=1
MM1001 N_A_69_260#_M1001_d N_CIN_M1001_g A_315_75# VNB NLOWVT L=0.15 W=0.64
+ AD=0.1248 AS=0.0768 PD=1.03 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75001.6
+ SB=75005.5 A=0.096 P=1.58 MULT=1
MM1010 N_A_501_75#_M1010_d N_A_465_249#_M1010_g N_A_69_260#_M1001_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1152 AS=0.1248 PD=1 PS=1.03 NRD=7.488 NRS=20.616 M=1
+ R=4.26667 SA=75002.1 SB=75005 A=0.096 P=1.58 MULT=1
MM1014 N_VGND_M1014_d N_B_M1014_g N_A_501_75#_M1010_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.169075 AS=0.1152 PD=1.275 PS=1 NRD=39.216 NRS=0 M=1 R=4.26667 SA=75002.7
+ SB=75004.5 A=0.096 P=1.58 MULT=1
MM1016 N_A_501_75#_M1016_d N_A_M1016_g N_VGND_M1014_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.169075 PD=0.92 PS=1.275 NRD=0 NRS=39.216 M=1 R=4.26667
+ SA=75003.2 SB=75003.9 A=0.096 P=1.58 MULT=1
MM1008 N_VGND_M1008_d N_CIN_M1008_g N_A_501_75#_M1016_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1584 AS=0.0896 PD=1.135 PS=0.92 NRD=26.244 NRS=0 M=1 R=4.26667 SA=75003.7
+ SB=75003.4 A=0.096 P=1.58 MULT=1
MM1002 A_936_75# N_A_M1002_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.64 AD=0.0768
+ AS=0.1584 PD=0.88 PS=1.135 NRD=12.18 NRS=14.052 M=1 R=4.26667 SA=75004.3
+ SB=75002.8 A=0.096 P=1.58 MULT=1
MM1017 N_A_465_249#_M1017_d N_B_M1017_g A_936_75# VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0768 PD=0.92 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75004.7
+ SB=75002.4 A=0.096 P=1.58 MULT=1
MM1024 N_A_1100_75#_M1024_d N_CIN_M1024_g N_A_465_249#_M1017_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.3596 AS=0.0896 PD=1.73 PS=0.92 NRD=95.028 NRS=0 M=1 R=4.26667
+ SA=75005.1 SB=75002 A=0.096 P=1.58 MULT=1
MM1023 N_VGND_M1023_d N_A_M1023_g N_A_1100_75#_M1024_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.212275 AS=0.3596 PD=1.41 PS=1.73 NRD=51.876 NRS=2.808 M=1 R=4.26667
+ SA=75006.2 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1015 N_A_1100_75#_M1015_d N_B_M1015_g N_VGND_M1023_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1696 AS=0.212275 PD=1.81 PS=1.41 NRD=0 NRS=51.876 M=1 R=4.26667
+ SA=75006.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1018 N_COUT_M1018_d N_A_465_249#_M1018_g N_VGND_M1018_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1998 AS=0.1961 PD=2.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1021 N_VPWR_M1021_d N_A_69_260#_M1021_g N_SUM_M1021_s VPB PSHORT L=0.18 W=1.12
+ AD=0.193464 AS=0.3024 PD=1.53736 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90004.9 A=0.2016 P=2.6 MULT=1
MM1027 A_220_368# N_A_M1027_g N_VPWR_M1021_d VPB PSHORT L=0.18 W=1 AD=0.171687
+ AS=0.172736 PD=1.43 PS=1.37264 NRD=22.9702 NRS=12.1352 M=1 R=5.55556
+ SA=90000.7 SB=90004.9 A=0.18 P=2.36 MULT=1
MM1003 A_321_389# N_B_M1003_g A_220_368# VPB PSHORT L=0.18 W=1 AD=0.180875
+ AS=0.171687 PD=1.535 PS=1.43 NRD=24.7826 NRS=22.9702 M=1 R=5.55556 SA=90001.1
+ SB=90004.5 A=0.18 P=2.36 MULT=1
MM1004 N_A_69_260#_M1004_d N_CIN_M1004_g A_321_389# VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.180875 PD=1.27 PS=1.535 NRD=0 NRS=24.7826 M=1 R=5.55556
+ SA=90001.4 SB=90005 A=0.18 P=2.36 MULT=1
MM1006 N_A_512_347#_M1006_d N_A_465_249#_M1006_g N_A_69_260#_M1004_d VPB PSHORT
+ L=0.18 W=1 AD=0.1525 AS=0.135 PD=1.305 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90001.8 SB=90004.6 A=0.18 P=2.36 MULT=1
MM1025 N_VPWR_M1025_d N_B_M1025_g N_A_512_347#_M1006_d VPB PSHORT L=0.18 W=1
+ AD=0.228637 AS=0.1525 PD=1.61 PS=1.305 NRD=34.1992 NRS=0.3152 M=1 R=5.55556
+ SA=90002.3 SB=90004.1 A=0.18 P=2.36 MULT=1
MM1012 N_A_512_347#_M1012_d N_A_M1012_g N_VPWR_M1025_d VPB PSHORT L=0.18 W=1
+ AD=0.1625 AS=0.228637 PD=1.325 PS=1.61 NRD=0 NRS=34.1992 M=1 R=5.55556
+ SA=90002.9 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_CIN_M1005_g N_A_512_347#_M1012_d VPB PSHORT L=0.18 W=1
+ AD=0.14 AS=0.1625 PD=1.28 PS=1.325 NRD=0 NRS=9.8303 M=1 R=5.55556 SA=90003.4
+ SB=90003 A=0.18 P=2.36 MULT=1
MM1019 A_919_347# N_A_M1019_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=1 AD=0.1625
+ AS=0.14 PD=1.325 PS=1.28 NRD=21.1578 NRS=0.9653 M=1 R=5.55556 SA=90003.9
+ SB=90002.5 A=0.18 P=2.36 MULT=1
MM1013 N_A_465_249#_M1013_d N_B_M1013_g A_919_347# VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.1625 PD=1.27 PS=1.325 NRD=0 NRS=21.1578 M=1 R=5.55556 SA=90004.4
+ SB=90002 A=0.18 P=2.36 MULT=1
MM1020 N_A_1110_347#_M1020_d N_CIN_M1020_g N_A_465_249#_M1013_d VPB PSHORT
+ L=0.18 W=1 AD=0.2075 AS=0.135 PD=1.415 PS=1.27 NRD=27.5603 NRS=0 M=1 R=5.55556
+ SA=90004.8 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1022 N_VPWR_M1022_d N_A_M1022_g N_A_1110_347#_M1020_d VPB PSHORT L=0.18 W=1
+ AD=0.334062 AS=0.2075 PD=1.73 PS=1.415 NRD=0 NRS=0 M=1 R=5.55556 SA=90005.4
+ SB=90001 A=0.18 P=2.36 MULT=1
MM1009 N_A_1110_347#_M1009_d N_B_M1009_g N_VPWR_M1022_d VPB PSHORT L=0.18 W=1
+ AD=0.32 AS=0.334062 PD=2.64 PS=1.73 NRD=6.8753 NRS=0 M=1 R=5.55556 SA=90005.9
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1007 N_COUT_M1007_d N_A_465_249#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18
+ W=1.12 AD=0.3024 AS=0.3136 PD=2.78 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX28_noxref VNB VPB NWDIODE A=17.4051 P=21.97
c_83 VNB 0 1.97438e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__fa_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__o2111a_4.pxi.spice
* Created: Fri Aug 28 17:51:48 2020
* 
x_PM_SKY130_FD_SC_MS__O2111A_4%D1 N_D1_M1000_g N_D1_M1010_g N_D1_c_150_n
+ N_D1_M1011_g N_D1_M1023_g N_D1_c_152_n D1 N_D1_c_153_n N_D1_c_154_n
+ PM_SKY130_FD_SC_MS__O2111A_4%D1
x_PM_SKY130_FD_SC_MS__O2111A_4%C1 N_C1_c_207_n N_C1_M1001_g N_C1_M1024_g
+ N_C1_c_208_n N_C1_M1008_g N_C1_M1025_g C1 C1 N_C1_c_210_n
+ PM_SKY130_FD_SC_MS__O2111A_4%C1
x_PM_SKY130_FD_SC_MS__O2111A_4%B1 N_B1_M1013_g N_B1_M1004_g N_B1_M1020_g
+ N_B1_M1026_g B1 N_B1_c_261_n PM_SKY130_FD_SC_MS__O2111A_4%B1
x_PM_SKY130_FD_SC_MS__O2111A_4%A2 N_A2_M1002_g N_A2_M1007_g N_A2_M1003_g
+ N_A2_M1027_g A2 A2 A2 A2 N_A2_c_311_n PM_SKY130_FD_SC_MS__O2111A_4%A2
x_PM_SKY130_FD_SC_MS__O2111A_4%A1 N_A1_M1005_g N_A1_M1018_g N_A1_M1014_g
+ N_A1_c_364_n N_A1_M1022_g A1 N_A1_c_362_n PM_SKY130_FD_SC_MS__O2111A_4%A1
x_PM_SKY130_FD_SC_MS__O2111A_4%A_27_392# N_A_27_392#_M1010_d N_A_27_392#_M1000_s
+ N_A_27_392#_M1023_s N_A_27_392#_M1025_d N_A_27_392#_M1020_s
+ N_A_27_392#_M1003_d N_A_27_392#_M1006_g N_A_27_392#_M1015_g
+ N_A_27_392#_M1009_g N_A_27_392#_M1016_g N_A_27_392#_M1012_g
+ N_A_27_392#_M1017_g N_A_27_392#_c_410_n N_A_27_392#_c_411_n
+ N_A_27_392#_M1019_g N_A_27_392#_M1021_g N_A_27_392#_c_414_n
+ N_A_27_392#_c_423_n N_A_27_392#_c_415_n N_A_27_392#_c_425_n
+ N_A_27_392#_c_426_n N_A_27_392#_c_427_n N_A_27_392#_c_428_n
+ N_A_27_392#_c_429_n N_A_27_392#_c_430_n N_A_27_392#_c_431_n
+ N_A_27_392#_c_432_n N_A_27_392#_c_416_n N_A_27_392#_c_565_p
+ N_A_27_392#_c_433_n N_A_27_392#_c_417_n N_A_27_392#_c_504_p
+ N_A_27_392#_c_434_n N_A_27_392#_c_435_n N_A_27_392#_c_436_n
+ N_A_27_392#_c_437_n PM_SKY130_FD_SC_MS__O2111A_4%A_27_392#
x_PM_SKY130_FD_SC_MS__O2111A_4%VPWR N_VPWR_M1000_d N_VPWR_M1024_s N_VPWR_M1013_d
+ N_VPWR_M1018_s N_VPWR_M1022_s N_VPWR_M1016_d N_VPWR_M1021_d N_VPWR_c_626_n
+ N_VPWR_c_627_n N_VPWR_c_628_n N_VPWR_c_629_n N_VPWR_c_630_n N_VPWR_c_631_n
+ N_VPWR_c_632_n N_VPWR_c_633_n N_VPWR_c_634_n N_VPWR_c_635_n N_VPWR_c_636_n
+ N_VPWR_c_637_n N_VPWR_c_638_n VPWR N_VPWR_c_639_n N_VPWR_c_640_n
+ N_VPWR_c_641_n N_VPWR_c_642_n N_VPWR_c_643_n N_VPWR_c_644_n N_VPWR_c_645_n
+ N_VPWR_c_646_n N_VPWR_c_625_n PM_SKY130_FD_SC_MS__O2111A_4%VPWR
x_PM_SKY130_FD_SC_MS__O2111A_4%A_750_392# N_A_750_392#_M1002_s
+ N_A_750_392#_M1018_d N_A_750_392#_c_747_n N_A_750_392#_c_750_n
+ N_A_750_392#_c_748_n PM_SKY130_FD_SC_MS__O2111A_4%A_750_392#
x_PM_SKY130_FD_SC_MS__O2111A_4%X N_X_M1006_d N_X_M1012_d N_X_M1015_s N_X_M1017_s
+ N_X_c_770_n N_X_c_785_n N_X_c_779_n N_X_c_771_n N_X_c_772_n N_X_c_797_n
+ N_X_c_773_n N_X_c_780_n N_X_c_781_n N_X_c_774_n N_X_c_775_n N_X_c_776_n
+ N_X_c_777_n N_X_c_821_n X PM_SKY130_FD_SC_MS__O2111A_4%X
x_PM_SKY130_FD_SC_MS__O2111A_4%A_27_74# N_A_27_74#_M1010_s N_A_27_74#_M1011_s
+ N_A_27_74#_M1008_s N_A_27_74#_c_850_n N_A_27_74#_c_851_n N_A_27_74#_c_852_n
+ N_A_27_74#_c_853_n N_A_27_74#_c_854_n N_A_27_74#_c_855_n N_A_27_74#_c_856_n
+ PM_SKY130_FD_SC_MS__O2111A_4%A_27_74#
x_PM_SKY130_FD_SC_MS__O2111A_4%A_287_74# N_A_287_74#_M1001_d N_A_287_74#_M1004_d
+ N_A_287_74#_c_889_n N_A_287_74#_c_890_n N_A_287_74#_c_891_n
+ PM_SKY130_FD_SC_MS__O2111A_4%A_287_74#
x_PM_SKY130_FD_SC_MS__O2111A_4%A_477_198# N_A_477_198#_M1004_s
+ N_A_477_198#_M1026_s N_A_477_198#_M1027_d N_A_477_198#_M1005_d
+ N_A_477_198#_c_918_n N_A_477_198#_c_928_n N_A_477_198#_c_919_n
+ N_A_477_198#_c_938_n N_A_477_198#_c_920_n N_A_477_198#_c_921_n
+ N_A_477_198#_c_922_n N_A_477_198#_c_923_n N_A_477_198#_c_924_n
+ N_A_477_198#_c_925_n PM_SKY130_FD_SC_MS__O2111A_4%A_477_198#
x_PM_SKY130_FD_SC_MS__O2111A_4%VGND N_VGND_M1007_s N_VGND_M1005_s N_VGND_M1014_s
+ N_VGND_M1009_s N_VGND_M1019_s N_VGND_c_982_n N_VGND_c_983_n N_VGND_c_984_n
+ N_VGND_c_985_n N_VGND_c_986_n N_VGND_c_987_n N_VGND_c_988_n N_VGND_c_989_n
+ N_VGND_c_990_n N_VGND_c_991_n N_VGND_c_992_n N_VGND_c_993_n VGND
+ N_VGND_c_994_n N_VGND_c_995_n N_VGND_c_996_n N_VGND_c_997_n
+ PM_SKY130_FD_SC_MS__O2111A_4%VGND
cc_1 VNB N_D1_M1010_g 0.0398087f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.74
cc_2 VNB N_D1_c_150_n 0.00856567f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.705
cc_3 VNB N_D1_M1011_g 0.0367314f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.74
cc_4 VNB N_D1_c_152_n 0.00691234f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.705
cc_5 VNB N_D1_c_153_n 0.0245373f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_6 VNB N_D1_c_154_n 0.00919084f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_7 VNB N_C1_c_207_n 0.014489f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.78
cc_8 VNB N_C1_c_208_n 0.0173034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB C1 0.00620616f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.38
cc_10 VNB N_C1_c_210_n 0.0712778f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_11 VNB N_B1_M1004_g 0.0254353f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.74
cc_12 VNB N_B1_M1026_g 0.0198802f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.78
cc_13 VNB B1 9.27509e-19 $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.38
cc_14 VNB N_B1_c_261_n 0.0330379f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_15 VNB N_A2_M1007_g 0.0201199f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.74
cc_16 VNB N_A2_M1027_g 0.026686f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.78
cc_17 VNB A2 0.0142547f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_18 VNB N_A2_c_311_n 0.0285134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_M1005_g 0.0363489f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.38
cc_20 VNB N_A1_M1014_g 0.0297668f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.63
cc_21 VNB A1 9.25683e-19 $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.38
cc_22 VNB N_A1_c_362_n 0.0276117f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_23 VNB N_A_27_392#_M1006_g 0.024894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_392#_M1009_g 0.024924f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_392#_M1012_g 0.0249207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_392#_c_410_n 0.00880736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_392#_c_411_n 0.0560835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_392#_M1019_g 0.0255042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_392#_M1021_g 0.00983424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_392#_c_414_n 0.00854837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_392#_c_415_n 0.00406729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_392#_c_416_n 0.00516444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_392#_c_417_n 0.00199603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_625_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_X_c_770_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.78
cc_36 VNB N_X_c_771_n 0.00323083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_X_c_772_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.615
cc_38 VNB N_X_c_773_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.78
cc_39 VNB N_X_c_774_n 0.00997592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_X_c_775_n 0.0126045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_776_n 8.8527e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_X_c_777_n 0.00273044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB X 0.0155405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_27_74#_c_850_n 0.0167032f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.705
cc_45 VNB N_A_27_74#_c_851_n 0.0219399f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.74
cc_46 VNB N_A_27_74#_c_852_n 0.00272448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_27_74#_c_853_n 0.00226074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_27_74#_c_854_n 0.00123754f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.45
cc_49 VNB N_A_27_74#_c_855_n 0.00987713f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.78
cc_50 VNB N_A_27_74#_c_856_n 0.0027795f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_51 VNB N_A_287_74#_c_889_n 0.0168718f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.74
cc_52 VNB N_A_287_74#_c_890_n 0.00289336f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.74
cc_53 VNB N_A_287_74#_c_891_n 0.00264166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_477_198#_c_918_n 0.0080669f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=0.74
cc_55 VNB N_A_477_198#_c_919_n 0.00267457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_477_198#_c_920_n 0.0101622f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.78
cc_57 VNB N_A_477_198#_c_921_n 0.0252068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_477_198#_c_922_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_477_198#_c_923_n 0.00108544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_477_198#_c_924_n 0.00230918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_477_198#_c_925_n 0.0025485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_982_n 0.0206912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_983_n 0.0166086f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.615
cc_64 VNB N_VGND_c_984_n 0.0151155f $X=-0.19 $Y=-0.245 $X2=0.407 $Y2=1.705
cc_65 VNB N_VGND_c_985_n 0.00830803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_986_n 0.0131737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_987_n 0.029666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_988_n 0.0952344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_989_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_990_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_991_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_992_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_993_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_994_n 0.0222872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_995_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_996_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_997_n 0.456094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VPB N_D1_M1000_g 0.0315139f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.38
cc_79 VPB N_D1_c_150_n 0.00787515f $X=-0.19 $Y=1.66 $X2=0.855 $Y2=1.705
cc_80 VPB N_D1_M1023_g 0.0229449f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.38
cc_81 VPB N_D1_c_152_n 0.00579753f $X=-0.19 $Y=1.66 $X2=1 $Y2=1.705
cc_82 VPB N_D1_c_153_n 0.0128818f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_83 VPB N_D1_c_154_n 0.0054581f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_84 VPB N_C1_M1024_g 0.0224695f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=0.74
cc_85 VPB N_C1_M1025_g 0.0238628f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=0.74
cc_86 VPB C1 0.00250401f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.38
cc_87 VPB N_C1_c_210_n 0.0169586f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_88 VPB N_B1_M1013_g 0.023242f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.38
cc_89 VPB N_B1_M1020_g 0.0228467f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.63
cc_90 VPB B1 0.00138027f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.38
cc_91 VPB N_B1_c_261_n 0.0224208f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_92 VPB N_A2_M1002_g 0.0252218f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.38
cc_93 VPB N_A2_M1003_g 0.0294273f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=1.63
cc_94 VPB A2 0.0119806f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_95 VPB N_A2_c_311_n 0.0168375f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A1_M1018_g 0.0283315f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=0.74
cc_97 VPB N_A1_c_364_n 0.0184525f $X=-0.19 $Y=1.66 $X2=0.93 $Y2=0.74
cc_98 VPB A1 8.34758e-19 $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.38
cc_99 VPB N_A1_c_362_n 0.0227254f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_100 VPB N_A_27_392#_M1015_g 0.0216544f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.45
cc_101 VPB N_A_27_392#_M1016_g 0.0212802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_27_392#_M1017_g 0.0206688f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_27_392#_c_411_n 0.00889192f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_27_392#_M1021_g 0.0273926f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_27_392#_c_423_n 0.00341815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_27_392#_c_415_n 0.00312231f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_27_392#_c_425_n 0.00254216f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_27_392#_c_426_n 0.0067225f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_27_392#_c_427_n 0.00511584f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_27_392#_c_428_n 7.12025e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_27_392#_c_429_n 0.0208772f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_27_392#_c_430_n 0.00241371f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_27_392#_c_431_n 0.00477769f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_27_392#_c_432_n 0.00136086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_27_392#_c_433_n 0.039485f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_27_392#_c_434_n 0.00532065f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_27_392#_c_435_n 0.0150875f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_27_392#_c_436_n 0.00403686f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_27_392#_c_437_n 0.00677628f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_626_n 0.0191643f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.615
cc_121 VPB N_VPWR_c_627_n 0.0193866f $X=-0.19 $Y=1.66 $X2=0.407 $Y2=1.705
cc_122 VPB N_VPWR_c_628_n 0.0156403f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_629_n 0.0127777f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_630_n 0.0127782f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_631_n 0.00582228f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_632_n 0.00274649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_633_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_634_n 0.0594105f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_635_n 0.0216142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_636_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_637_n 0.0432862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_638_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_639_n 0.0198433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_640_n 0.0198086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_641_n 0.0172173f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_642_n 0.0175706f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_643_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_644_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_645_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_646_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_625_n 0.110461f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_750_392#_c_747_n 0.0124765f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=0.74
cc_143 VPB N_A_750_392#_c_748_n 0.00231675f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.38
cc_144 VPB N_X_c_779_n 0.00275545f $X=-0.19 $Y=1.66 $X2=1 $Y2=1.705
cc_145 VPB N_X_c_780_n 0.0016227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_X_c_781_n 0.00202354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 N_D1_M1011_g N_C1_c_207_n 0.0187348f $X=0.93 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_148 N_D1_M1023_g N_C1_M1024_g 0.0145327f $X=1.055 $Y=2.38 $X2=0 $Y2=0
cc_149 N_D1_M1011_g C1 0.00173097f $X=0.93 $Y=0.74 $X2=0 $Y2=0
cc_150 N_D1_c_152_n C1 0.00681629f $X=1 $Y=1.705 $X2=0 $Y2=0
cc_151 N_D1_M1011_g N_C1_c_210_n 0.00802884f $X=0.93 $Y=0.74 $X2=0 $Y2=0
cc_152 N_D1_c_152_n N_C1_c_210_n 0.0145327f $X=1 $Y=1.705 $X2=0 $Y2=0
cc_153 N_D1_M1000_g N_A_27_392#_c_423_n 0.0148113f $X=0.505 $Y=2.38 $X2=0 $Y2=0
cc_154 N_D1_c_150_n N_A_27_392#_c_423_n 0.00118094f $X=0.855 $Y=1.705 $X2=0
+ $Y2=0
cc_155 N_D1_c_154_n N_A_27_392#_c_423_n 0.00746443f $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_156 N_D1_M1000_g N_A_27_392#_c_415_n 0.00389722f $X=0.505 $Y=2.38 $X2=0 $Y2=0
cc_157 N_D1_M1010_g N_A_27_392#_c_415_n 0.00680216f $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_158 N_D1_c_150_n N_A_27_392#_c_415_n 0.00987117f $X=0.855 $Y=1.705 $X2=0
+ $Y2=0
cc_159 N_D1_M1011_g N_A_27_392#_c_415_n 0.0114191f $X=0.93 $Y=0.74 $X2=0 $Y2=0
cc_160 N_D1_M1023_g N_A_27_392#_c_415_n 0.0041557f $X=1.055 $Y=2.38 $X2=0 $Y2=0
cc_161 N_D1_c_152_n N_A_27_392#_c_415_n 0.00297968f $X=1 $Y=1.705 $X2=0 $Y2=0
cc_162 N_D1_c_153_n N_A_27_392#_c_415_n 0.00120381f $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_163 N_D1_c_154_n N_A_27_392#_c_415_n 0.0247006f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_164 N_D1_M1023_g N_A_27_392#_c_425_n 0.016832f $X=1.055 $Y=2.38 $X2=0 $Y2=0
cc_165 N_D1_M1000_g N_A_27_392#_c_433_n 0.0147368f $X=0.505 $Y=2.38 $X2=0 $Y2=0
cc_166 N_D1_M1023_g N_A_27_392#_c_433_n 6.38451e-19 $X=1.055 $Y=2.38 $X2=0 $Y2=0
cc_167 N_D1_c_153_n N_A_27_392#_c_433_n 0.00454265f $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_168 N_D1_c_154_n N_A_27_392#_c_433_n 0.0272436f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_169 N_D1_M1010_g N_A_27_392#_c_417_n 0.00603749f $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_170 N_D1_c_150_n N_A_27_392#_c_417_n 0.00376859f $X=0.855 $Y=1.705 $X2=0
+ $Y2=0
cc_171 N_D1_M1011_g N_A_27_392#_c_417_n 0.00453298f $X=0.93 $Y=0.74 $X2=0 $Y2=0
cc_172 N_D1_c_153_n N_A_27_392#_c_417_n 7.64322e-19 $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_173 N_D1_M1000_g N_A_27_392#_c_434_n 6.38451e-19 $X=0.505 $Y=2.38 $X2=0 $Y2=0
cc_174 N_D1_M1023_g N_A_27_392#_c_434_n 0.0131758f $X=1.055 $Y=2.38 $X2=0 $Y2=0
cc_175 N_D1_M1000_g N_VPWR_c_626_n 0.00421336f $X=0.505 $Y=2.38 $X2=0 $Y2=0
cc_176 N_D1_c_150_n N_VPWR_c_626_n 6.81301e-19 $X=0.855 $Y=1.705 $X2=0 $Y2=0
cc_177 N_D1_M1023_g N_VPWR_c_626_n 0.00280405f $X=1.055 $Y=2.38 $X2=0 $Y2=0
cc_178 N_D1_M1023_g N_VPWR_c_627_n 0.00540023f $X=1.055 $Y=2.38 $X2=0 $Y2=0
cc_179 N_D1_M1000_g N_VPWR_c_639_n 0.00540023f $X=0.505 $Y=2.38 $X2=0 $Y2=0
cc_180 N_D1_M1000_g N_VPWR_c_625_n 0.00595788f $X=0.505 $Y=2.38 $X2=0 $Y2=0
cc_181 N_D1_M1023_g N_VPWR_c_625_n 0.00595788f $X=1.055 $Y=2.38 $X2=0 $Y2=0
cc_182 N_D1_M1010_g N_A_27_74#_c_851_n 9.80934e-19 $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_183 N_D1_c_153_n N_A_27_74#_c_851_n 0.00335778f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_184 N_D1_c_154_n N_A_27_74#_c_851_n 0.0133432f $X=0.385 $Y=1.615 $X2=0 $Y2=0
cc_185 N_D1_M1010_g N_A_27_74#_c_852_n 0.0182491f $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_186 N_D1_M1011_g N_A_27_74#_c_852_n 0.0169848f $X=0.93 $Y=0.74 $X2=0 $Y2=0
cc_187 N_D1_M1011_g N_A_27_74#_c_853_n 3.89484e-19 $X=0.93 $Y=0.74 $X2=0 $Y2=0
cc_188 N_D1_c_152_n N_A_27_74#_c_853_n 0.00113443f $X=1 $Y=1.705 $X2=0 $Y2=0
cc_189 N_D1_M1010_g N_VGND_c_988_n 0.00278271f $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_190 N_D1_M1011_g N_VGND_c_988_n 0.00278271f $X=0.93 $Y=0.74 $X2=0 $Y2=0
cc_191 N_D1_M1010_g N_VGND_c_997_n 0.00357103f $X=0.5 $Y=0.74 $X2=0 $Y2=0
cc_192 N_D1_M1011_g N_VGND_c_997_n 0.00353526f $X=0.93 $Y=0.74 $X2=0 $Y2=0
cc_193 N_C1_M1025_g N_B1_M1013_g 0.0157865f $X=2.005 $Y=2.38 $X2=0 $Y2=0
cc_194 N_C1_c_210_n N_B1_c_261_n 0.0209634f $X=1.79 $Y=1.482 $X2=0 $Y2=0
cc_195 C1 N_A_27_392#_c_415_n 0.0232485f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_196 N_C1_c_210_n N_A_27_392#_c_415_n 0.00145788f $X=1.79 $Y=1.482 $X2=0 $Y2=0
cc_197 C1 N_A_27_392#_c_425_n 0.00210849f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_198 N_C1_M1024_g N_A_27_392#_c_426_n 0.0132272f $X=1.505 $Y=2.38 $X2=0 $Y2=0
cc_199 N_C1_M1025_g N_A_27_392#_c_426_n 0.0224537f $X=2.005 $Y=2.38 $X2=0 $Y2=0
cc_200 C1 N_A_27_392#_c_426_n 0.0257108f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_201 N_C1_c_210_n N_A_27_392#_c_426_n 0.00414484f $X=1.79 $Y=1.482 $X2=0 $Y2=0
cc_202 N_C1_c_207_n N_A_27_392#_c_417_n 6.23466e-19 $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_203 N_C1_M1024_g N_A_27_392#_c_434_n 0.0128698f $X=1.505 $Y=2.38 $X2=0 $Y2=0
cc_204 N_C1_M1025_g N_A_27_392#_c_434_n 0.00102447f $X=2.005 $Y=2.38 $X2=0 $Y2=0
cc_205 C1 N_A_27_392#_c_434_n 0.0286741f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_206 N_C1_M1025_g N_A_27_392#_c_435_n 0.00487985f $X=2.005 $Y=2.38 $X2=0 $Y2=0
cc_207 N_C1_M1024_g N_VPWR_c_627_n 0.00540023f $X=1.505 $Y=2.38 $X2=0 $Y2=0
cc_208 N_C1_M1024_g N_VPWR_c_628_n 0.00262659f $X=1.505 $Y=2.38 $X2=0 $Y2=0
cc_209 N_C1_M1025_g N_VPWR_c_628_n 0.0125741f $X=2.005 $Y=2.38 $X2=0 $Y2=0
cc_210 N_C1_M1025_g N_VPWR_c_629_n 5.95894e-19 $X=2.005 $Y=2.38 $X2=0 $Y2=0
cc_211 N_C1_M1025_g N_VPWR_c_635_n 0.00468007f $X=2.005 $Y=2.38 $X2=0 $Y2=0
cc_212 N_C1_M1024_g N_VPWR_c_625_n 0.00595788f $X=1.505 $Y=2.38 $X2=0 $Y2=0
cc_213 N_C1_M1025_g N_VPWR_c_625_n 0.004998f $X=2.005 $Y=2.38 $X2=0 $Y2=0
cc_214 N_C1_c_207_n N_A_27_74#_c_853_n 4.08775e-19 $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_215 C1 N_A_27_74#_c_853_n 0.00820373f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_216 N_C1_c_207_n N_A_27_74#_c_856_n 0.0122675f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_217 N_C1_c_208_n N_A_27_74#_c_856_n 0.0113109f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_218 N_C1_c_208_n N_A_287_74#_c_889_n 0.0127544f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_219 C1 N_A_287_74#_c_889_n 0.00143794f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_220 N_C1_c_210_n N_A_287_74#_c_889_n 0.00564282f $X=1.79 $Y=1.482 $X2=0 $Y2=0
cc_221 N_C1_c_207_n N_A_287_74#_c_890_n 0.00805309f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_222 N_C1_c_208_n N_A_287_74#_c_890_n 0.0169798f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_223 C1 N_A_287_74#_c_890_n 0.0167849f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_224 N_C1_c_210_n N_A_287_74#_c_890_n 0.00337453f $X=1.79 $Y=1.482 $X2=0 $Y2=0
cc_225 N_C1_c_208_n N_A_477_198#_c_918_n 0.00673386f $X=1.79 $Y=1.185 $X2=0
+ $Y2=0
cc_226 N_C1_c_207_n N_VGND_c_988_n 0.00278271f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_227 N_C1_c_208_n N_VGND_c_988_n 0.00278271f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_228 N_C1_c_207_n N_VGND_c_997_n 0.00353526f $X=1.36 $Y=1.185 $X2=0 $Y2=0
cc_229 N_C1_c_208_n N_VGND_c_997_n 0.00358427f $X=1.79 $Y=1.185 $X2=0 $Y2=0
cc_230 N_B1_M1020_g N_A2_M1002_g 0.0171533f $X=3.075 $Y=2.38 $X2=0 $Y2=0
cc_231 N_B1_M1026_g N_A2_M1007_g 0.0159516f $X=3.255 $Y=0.91 $X2=0 $Y2=0
cc_232 B1 A2 0.0276607f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_233 N_B1_c_261_n A2 0.00240023f $X=3.15 $Y=1.615 $X2=0 $Y2=0
cc_234 B1 N_A2_c_311_n 3.40273e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_235 N_B1_c_261_n N_A2_c_311_n 0.0183165f $X=3.15 $Y=1.615 $X2=0 $Y2=0
cc_236 N_B1_M1013_g N_A_27_392#_c_427_n 0.0188596f $X=2.625 $Y=2.38 $X2=0 $Y2=0
cc_237 N_B1_M1020_g N_A_27_392#_c_427_n 0.0169379f $X=3.075 $Y=2.38 $X2=0 $Y2=0
cc_238 B1 N_A_27_392#_c_427_n 0.016966f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_239 N_B1_c_261_n N_A_27_392#_c_427_n 0.003196f $X=3.15 $Y=1.615 $X2=0 $Y2=0
cc_240 N_B1_M1020_g N_A_27_392#_c_428_n 0.00512167f $X=3.075 $Y=2.38 $X2=0 $Y2=0
cc_241 N_B1_M1020_g N_A_27_392#_c_431_n 2.65336e-19 $X=3.075 $Y=2.38 $X2=0 $Y2=0
cc_242 N_B1_M1013_g N_A_27_392#_c_435_n 0.00487985f $X=2.625 $Y=2.38 $X2=0 $Y2=0
cc_243 B1 N_A_27_392#_c_436_n 0.00796601f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_244 N_B1_c_261_n N_A_27_392#_c_436_n 0.00128085f $X=3.15 $Y=1.615 $X2=0 $Y2=0
cc_245 N_B1_M1013_g N_VPWR_c_628_n 5.95894e-19 $X=2.625 $Y=2.38 $X2=0 $Y2=0
cc_246 N_B1_M1013_g N_VPWR_c_629_n 0.0126452f $X=2.625 $Y=2.38 $X2=0 $Y2=0
cc_247 N_B1_M1020_g N_VPWR_c_629_n 0.0115733f $X=3.075 $Y=2.38 $X2=0 $Y2=0
cc_248 N_B1_M1013_g N_VPWR_c_635_n 0.00468007f $X=2.625 $Y=2.38 $X2=0 $Y2=0
cc_249 N_B1_M1020_g N_VPWR_c_637_n 0.00468007f $X=3.075 $Y=2.38 $X2=0 $Y2=0
cc_250 N_B1_M1013_g N_VPWR_c_625_n 0.004998f $X=2.625 $Y=2.38 $X2=0 $Y2=0
cc_251 N_B1_M1020_g N_VPWR_c_625_n 0.004998f $X=3.075 $Y=2.38 $X2=0 $Y2=0
cc_252 N_B1_M1004_g N_A_27_74#_c_855_n 0.00324596f $X=2.825 $Y=0.91 $X2=0 $Y2=0
cc_253 N_B1_M1004_g N_A_287_74#_c_889_n 0.0109615f $X=2.825 $Y=0.91 $X2=0 $Y2=0
cc_254 N_B1_M1004_g N_A_287_74#_c_891_n 0.00936405f $X=2.825 $Y=0.91 $X2=0 $Y2=0
cc_255 N_B1_c_261_n N_A_477_198#_c_918_n 0.00560629f $X=3.15 $Y=1.615 $X2=0
+ $Y2=0
cc_256 N_B1_M1004_g N_A_477_198#_c_928_n 0.0104018f $X=2.825 $Y=0.91 $X2=0 $Y2=0
cc_257 N_B1_M1026_g N_A_477_198#_c_928_n 0.0125752f $X=3.255 $Y=0.91 $X2=0 $Y2=0
cc_258 B1 N_A_477_198#_c_928_n 0.0216895f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_259 N_B1_c_261_n N_A_477_198#_c_928_n 7.11275e-19 $X=3.15 $Y=1.615 $X2=0
+ $Y2=0
cc_260 N_B1_M1004_g N_A_477_198#_c_919_n 9.14331e-19 $X=2.825 $Y=0.91 $X2=0
+ $Y2=0
cc_261 N_B1_M1026_g N_A_477_198#_c_919_n 0.00758705f $X=3.255 $Y=0.91 $X2=0
+ $Y2=0
cc_262 N_B1_M1004_g N_A_477_198#_c_923_n 0.0023175f $X=2.825 $Y=0.91 $X2=0 $Y2=0
cc_263 N_B1_M1026_g N_A_477_198#_c_924_n 0.00103783f $X=3.255 $Y=0.91 $X2=0
+ $Y2=0
cc_264 B1 N_A_477_198#_c_924_n 7.22171e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_265 N_B1_M1026_g N_VGND_c_982_n 6.8897e-19 $X=3.255 $Y=0.91 $X2=0 $Y2=0
cc_266 N_B1_M1004_g N_VGND_c_988_n 0.00359961f $X=2.825 $Y=0.91 $X2=0 $Y2=0
cc_267 N_B1_M1026_g N_VGND_c_988_n 0.00444543f $X=3.255 $Y=0.91 $X2=0 $Y2=0
cc_268 N_B1_M1004_g N_VGND_c_997_n 0.00493565f $X=2.825 $Y=0.91 $X2=0 $Y2=0
cc_269 N_B1_M1026_g N_VGND_c_997_n 0.00493565f $X=3.255 $Y=0.91 $X2=0 $Y2=0
cc_270 A2 A1 0.0261825f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_271 A2 N_A1_c_362_n 0.0144217f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_272 N_A2_M1002_g N_A_27_392#_c_429_n 0.0146907f $X=3.66 $Y=2.46 $X2=0 $Y2=0
cc_273 N_A2_M1003_g N_A_27_392#_c_429_n 0.0140828f $X=4.16 $Y=2.46 $X2=0 $Y2=0
cc_274 A2 N_A_27_392#_c_429_n 0.122866f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_275 N_A2_c_311_n N_A_27_392#_c_429_n 0.00317828f $X=4.175 $Y=1.615 $X2=0
+ $Y2=0
cc_276 N_A2_M1002_g N_A_27_392#_c_430_n 0.0153671f $X=3.66 $Y=2.46 $X2=0 $Y2=0
cc_277 N_A2_M1003_g N_A_27_392#_c_430_n 0.00937508f $X=4.16 $Y=2.46 $X2=0 $Y2=0
cc_278 A2 N_A_27_392#_c_436_n 0.00575f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_279 N_A2_M1002_g N_A_27_392#_c_437_n 6.38845e-19 $X=3.66 $Y=2.46 $X2=0 $Y2=0
cc_280 N_A2_M1003_g N_A_27_392#_c_437_n 0.00854437f $X=4.16 $Y=2.46 $X2=0 $Y2=0
cc_281 N_A2_M1002_g N_VPWR_c_629_n 7.95254e-19 $X=3.66 $Y=2.46 $X2=0 $Y2=0
cc_282 N_A2_M1003_g N_VPWR_c_630_n 0.00136693f $X=4.16 $Y=2.46 $X2=0 $Y2=0
cc_283 N_A2_M1002_g N_VPWR_c_637_n 0.00333926f $X=3.66 $Y=2.46 $X2=0 $Y2=0
cc_284 N_A2_M1003_g N_VPWR_c_637_n 0.00335119f $X=4.16 $Y=2.46 $X2=0 $Y2=0
cc_285 N_A2_M1002_g N_VPWR_c_625_n 0.00428309f $X=3.66 $Y=2.46 $X2=0 $Y2=0
cc_286 N_A2_M1003_g N_VPWR_c_625_n 0.00427398f $X=4.16 $Y=2.46 $X2=0 $Y2=0
cc_287 N_A2_M1003_g N_A_750_392#_c_747_n 0.0133282f $X=4.16 $Y=2.46 $X2=0 $Y2=0
cc_288 N_A2_M1002_g N_A_750_392#_c_750_n 0.00650386f $X=3.66 $Y=2.46 $X2=0 $Y2=0
cc_289 N_A2_M1007_g N_A_477_198#_c_919_n 3.13308e-19 $X=3.685 $Y=0.91 $X2=0
+ $Y2=0
cc_290 N_A2_M1007_g N_A_477_198#_c_938_n 0.012601f $X=3.685 $Y=0.91 $X2=0 $Y2=0
cc_291 N_A2_M1027_g N_A_477_198#_c_938_n 0.0122289f $X=4.175 $Y=0.91 $X2=0 $Y2=0
cc_292 A2 N_A_477_198#_c_938_n 0.0433751f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_293 N_A2_c_311_n N_A_477_198#_c_938_n 0.00370549f $X=4.175 $Y=1.615 $X2=0
+ $Y2=0
cc_294 N_A2_M1007_g N_A_477_198#_c_920_n 9.05595e-19 $X=3.685 $Y=0.91 $X2=0
+ $Y2=0
cc_295 N_A2_M1027_g N_A_477_198#_c_920_n 0.00850927f $X=4.175 $Y=0.91 $X2=0
+ $Y2=0
cc_296 A2 N_A_477_198#_c_921_n 0.0465439f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_297 A2 N_A_477_198#_c_924_n 0.00597859f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_298 N_A2_M1027_g N_A_477_198#_c_925_n 4.27055e-19 $X=4.175 $Y=0.91 $X2=0
+ $Y2=0
cc_299 A2 N_A_477_198#_c_925_n 0.02594f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_300 N_A2_M1007_g N_VGND_c_982_n 0.00895009f $X=3.685 $Y=0.91 $X2=0 $Y2=0
cc_301 N_A2_M1027_g N_VGND_c_982_n 0.00539056f $X=4.175 $Y=0.91 $X2=0 $Y2=0
cc_302 N_A2_M1027_g N_VGND_c_983_n 0.00356388f $X=4.175 $Y=0.91 $X2=0 $Y2=0
cc_303 N_A2_M1007_g N_VGND_c_988_n 0.00384833f $X=3.685 $Y=0.91 $X2=0 $Y2=0
cc_304 N_A2_M1027_g N_VGND_c_994_n 0.00452252f $X=4.175 $Y=0.91 $X2=0 $Y2=0
cc_305 N_A2_M1007_g N_VGND_c_997_n 0.00414594f $X=3.685 $Y=0.91 $X2=0 $Y2=0
cc_306 N_A2_M1027_g N_VGND_c_997_n 0.00493565f $X=4.175 $Y=0.91 $X2=0 $Y2=0
cc_307 N_A1_M1014_g N_A_27_392#_M1006_g 0.0259675f $X=5.635 $Y=0.74 $X2=0 $Y2=0
cc_308 N_A1_c_362_n N_A_27_392#_M1015_g 0.0287084f $X=5.635 $Y=1.66 $X2=0 $Y2=0
cc_309 A1 N_A_27_392#_c_411_n 3.15573e-19 $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_310 N_A1_c_362_n N_A_27_392#_c_411_n 0.0100415f $X=5.635 $Y=1.66 $X2=0 $Y2=0
cc_311 N_A1_M1018_g N_A_27_392#_c_429_n 0.0161399f $X=5.22 $Y=2.46 $X2=0 $Y2=0
cc_312 N_A1_c_364_n N_A_27_392#_c_429_n 0.0196876f $X=5.67 $Y=1.87 $X2=0 $Y2=0
cc_313 A1 N_A_27_392#_c_429_n 0.0244987f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_314 N_A1_c_362_n N_A_27_392#_c_429_n 6.3257e-19 $X=5.635 $Y=1.66 $X2=0 $Y2=0
cc_315 A1 N_A_27_392#_c_432_n 0.00466348f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_316 N_A1_c_362_n N_A_27_392#_c_432_n 0.00431602f $X=5.635 $Y=1.66 $X2=0 $Y2=0
cc_317 N_A1_M1014_g N_A_27_392#_c_416_n 0.00252208f $X=5.635 $Y=0.74 $X2=0 $Y2=0
cc_318 A1 N_A_27_392#_c_416_n 0.0121153f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_319 N_A1_c_362_n N_A_27_392#_c_416_n 0.0022552f $X=5.635 $Y=1.66 $X2=0 $Y2=0
cc_320 N_A1_M1018_g N_VPWR_c_630_n 0.00534567f $X=5.22 $Y=2.46 $X2=0 $Y2=0
cc_321 N_A1_c_364_n N_VPWR_c_631_n 0.00687499f $X=5.67 $Y=1.87 $X2=0 $Y2=0
cc_322 N_A1_M1018_g N_VPWR_c_640_n 0.005209f $X=5.22 $Y=2.46 $X2=0 $Y2=0
cc_323 N_A1_c_364_n N_VPWR_c_640_n 0.005209f $X=5.67 $Y=1.87 $X2=0 $Y2=0
cc_324 N_A1_M1018_g N_VPWR_c_625_n 0.00986727f $X=5.22 $Y=2.46 $X2=0 $Y2=0
cc_325 N_A1_c_364_n N_VPWR_c_625_n 0.00983239f $X=5.67 $Y=1.87 $X2=0 $Y2=0
cc_326 N_A1_M1018_g N_A_750_392#_c_747_n 0.014819f $X=5.22 $Y=2.46 $X2=0 $Y2=0
cc_327 N_A1_M1018_g N_A_750_392#_c_748_n 0.0129461f $X=5.22 $Y=2.46 $X2=0 $Y2=0
cc_328 N_A1_c_364_n N_A_750_392#_c_748_n 0.00929437f $X=5.67 $Y=1.87 $X2=0 $Y2=0
cc_329 N_A1_M1005_g N_A_477_198#_c_920_n 0.00293386f $X=5.205 $Y=0.74 $X2=0
+ $Y2=0
cc_330 N_A1_M1005_g N_A_477_198#_c_921_n 0.0177833f $X=5.205 $Y=0.74 $X2=0 $Y2=0
cc_331 N_A1_M1014_g N_A_477_198#_c_921_n 0.00415797f $X=5.635 $Y=0.74 $X2=0
+ $Y2=0
cc_332 A1 N_A_477_198#_c_921_n 0.0150501f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_333 N_A1_c_362_n N_A_477_198#_c_921_n 7.88639e-19 $X=5.635 $Y=1.66 $X2=0
+ $Y2=0
cc_334 N_A1_M1005_g N_A_477_198#_c_922_n 3.92313e-19 $X=5.205 $Y=0.74 $X2=0
+ $Y2=0
cc_335 N_A1_M1014_g N_A_477_198#_c_922_n 3.92313e-19 $X=5.635 $Y=0.74 $X2=0
+ $Y2=0
cc_336 N_A1_M1005_g N_VGND_c_983_n 0.0114363f $X=5.205 $Y=0.74 $X2=0 $Y2=0
cc_337 N_A1_M1014_g N_VGND_c_983_n 5.01478e-19 $X=5.635 $Y=0.74 $X2=0 $Y2=0
cc_338 N_A1_M1005_g N_VGND_c_984_n 5.68935e-19 $X=5.205 $Y=0.74 $X2=0 $Y2=0
cc_339 N_A1_M1014_g N_VGND_c_984_n 0.0142039f $X=5.635 $Y=0.74 $X2=0 $Y2=0
cc_340 N_A1_c_362_n N_VGND_c_984_n 0.00170878f $X=5.635 $Y=1.66 $X2=0 $Y2=0
cc_341 N_A1_M1005_g N_VGND_c_990_n 0.00383152f $X=5.205 $Y=0.74 $X2=0 $Y2=0
cc_342 N_A1_M1014_g N_VGND_c_990_n 0.00383152f $X=5.635 $Y=0.74 $X2=0 $Y2=0
cc_343 N_A1_M1005_g N_VGND_c_997_n 0.0075754f $X=5.205 $Y=0.74 $X2=0 $Y2=0
cc_344 N_A1_M1014_g N_VGND_c_997_n 0.0075754f $X=5.635 $Y=0.74 $X2=0 $Y2=0
cc_345 N_A_27_392#_c_423_n N_VPWR_M1000_d 7.5517e-19 $X=0.72 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_346 N_A_27_392#_c_504_p N_VPWR_M1000_d 0.00208437f $X=0.805 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_347 N_A_27_392#_c_426_n N_VPWR_M1024_s 0.00232187f $X=2.15 $Y=2.035 $X2=0
+ $Y2=0
cc_348 N_A_27_392#_c_427_n N_VPWR_M1013_d 0.00175831f $X=3.22 $Y=2.035 $X2=0
+ $Y2=0
cc_349 N_A_27_392#_c_429_n N_VPWR_M1018_s 0.00422922f $X=5.975 $Y=2.035 $X2=0
+ $Y2=0
cc_350 N_A_27_392#_c_429_n N_VPWR_M1022_s 0.00673533f $X=5.975 $Y=2.035 $X2=0
+ $Y2=0
cc_351 N_A_27_392#_c_432_n N_VPWR_M1022_s 0.00130575f $X=6.06 $Y=1.95 $X2=0
+ $Y2=0
cc_352 N_A_27_392#_c_423_n N_VPWR_c_626_n 0.00496126f $X=0.72 $Y=2.035 $X2=0
+ $Y2=0
cc_353 N_A_27_392#_c_425_n N_VPWR_c_626_n 0.00128906f $X=1.115 $Y=2.035 $X2=0
+ $Y2=0
cc_354 N_A_27_392#_c_433_n N_VPWR_c_626_n 0.0197393f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_355 N_A_27_392#_c_504_p N_VPWR_c_626_n 0.0138281f $X=0.805 $Y=2.035 $X2=0
+ $Y2=0
cc_356 N_A_27_392#_c_434_n N_VPWR_c_626_n 0.0197393f $X=1.28 $Y=2.115 $X2=0
+ $Y2=0
cc_357 N_A_27_392#_c_434_n N_VPWR_c_627_n 0.00869594f $X=1.28 $Y=2.115 $X2=0
+ $Y2=0
cc_358 N_A_27_392#_c_426_n N_VPWR_c_628_n 0.0170697f $X=2.15 $Y=2.035 $X2=0
+ $Y2=0
cc_359 N_A_27_392#_c_434_n N_VPWR_c_628_n 0.0197393f $X=1.28 $Y=2.115 $X2=0
+ $Y2=0
cc_360 N_A_27_392#_c_435_n N_VPWR_c_628_n 0.0170056f $X=2.315 $Y=2.105 $X2=0
+ $Y2=0
cc_361 N_A_27_392#_c_427_n N_VPWR_c_629_n 0.0153378f $X=3.22 $Y=2.035 $X2=0
+ $Y2=0
cc_362 N_A_27_392#_c_428_n N_VPWR_c_629_n 0.0228151f $X=3.385 $Y=2.815 $X2=0
+ $Y2=0
cc_363 N_A_27_392#_c_431_n N_VPWR_c_629_n 0.0130717f $X=3.55 $Y=2.99 $X2=0 $Y2=0
cc_364 N_A_27_392#_c_435_n N_VPWR_c_629_n 0.0170056f $X=2.315 $Y=2.105 $X2=0
+ $Y2=0
cc_365 N_A_27_392#_c_437_n N_VPWR_c_630_n 0.0300014f $X=4.385 $Y=2.805 $X2=0
+ $Y2=0
cc_366 N_A_27_392#_M1015_g N_VPWR_c_631_n 0.0125355f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_367 N_A_27_392#_M1016_g N_VPWR_c_631_n 4.98789e-19 $X=6.705 $Y=2.4 $X2=0
+ $Y2=0
cc_368 N_A_27_392#_c_429_n N_VPWR_c_631_n 0.0226691f $X=5.975 $Y=2.035 $X2=0
+ $Y2=0
cc_369 N_A_27_392#_M1015_g N_VPWR_c_632_n 4.88604e-19 $X=6.205 $Y=2.4 $X2=0
+ $Y2=0
cc_370 N_A_27_392#_M1016_g N_VPWR_c_632_n 0.0118758f $X=6.705 $Y=2.4 $X2=0 $Y2=0
cc_371 N_A_27_392#_M1017_g N_VPWR_c_632_n 0.0121532f $X=7.155 $Y=2.4 $X2=0 $Y2=0
cc_372 N_A_27_392#_M1021_g N_VPWR_c_632_n 5.47803e-19 $X=7.605 $Y=2.4 $X2=0
+ $Y2=0
cc_373 N_A_27_392#_M1021_g N_VPWR_c_634_n 0.00540173f $X=7.605 $Y=2.4 $X2=0
+ $Y2=0
cc_374 N_A_27_392#_c_435_n N_VPWR_c_635_n 0.00884037f $X=2.315 $Y=2.105 $X2=0
+ $Y2=0
cc_375 N_A_27_392#_c_430_n N_VPWR_c_637_n 0.0421705f $X=4.22 $Y=2.99 $X2=0 $Y2=0
cc_376 N_A_27_392#_c_431_n N_VPWR_c_637_n 0.0236566f $X=3.55 $Y=2.99 $X2=0 $Y2=0
cc_377 N_A_27_392#_c_437_n N_VPWR_c_637_n 0.0226835f $X=4.385 $Y=2.805 $X2=0
+ $Y2=0
cc_378 N_A_27_392#_c_433_n N_VPWR_c_639_n 0.00876816f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_379 N_A_27_392#_M1015_g N_VPWR_c_641_n 0.00460063f $X=6.205 $Y=2.4 $X2=0
+ $Y2=0
cc_380 N_A_27_392#_M1016_g N_VPWR_c_641_n 0.00460063f $X=6.705 $Y=2.4 $X2=0
+ $Y2=0
cc_381 N_A_27_392#_M1017_g N_VPWR_c_642_n 0.00460063f $X=7.155 $Y=2.4 $X2=0
+ $Y2=0
cc_382 N_A_27_392#_M1021_g N_VPWR_c_642_n 0.005209f $X=7.605 $Y=2.4 $X2=0 $Y2=0
cc_383 N_A_27_392#_M1015_g N_VPWR_c_625_n 0.00909043f $X=6.205 $Y=2.4 $X2=0
+ $Y2=0
cc_384 N_A_27_392#_M1016_g N_VPWR_c_625_n 0.00909043f $X=6.705 $Y=2.4 $X2=0
+ $Y2=0
cc_385 N_A_27_392#_M1017_g N_VPWR_c_625_n 0.00908554f $X=7.155 $Y=2.4 $X2=0
+ $Y2=0
cc_386 N_A_27_392#_M1021_g N_VPWR_c_625_n 0.00985497f $X=7.605 $Y=2.4 $X2=0
+ $Y2=0
cc_387 N_A_27_392#_c_430_n N_VPWR_c_625_n 0.0236848f $X=4.22 $Y=2.99 $X2=0 $Y2=0
cc_388 N_A_27_392#_c_431_n N_VPWR_c_625_n 0.0128296f $X=3.55 $Y=2.99 $X2=0 $Y2=0
cc_389 N_A_27_392#_c_433_n N_VPWR_c_625_n 0.0108652f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_390 N_A_27_392#_c_434_n N_VPWR_c_625_n 0.010834f $X=1.28 $Y=2.115 $X2=0 $Y2=0
cc_391 N_A_27_392#_c_435_n N_VPWR_c_625_n 0.0108964f $X=2.315 $Y=2.105 $X2=0
+ $Y2=0
cc_392 N_A_27_392#_c_437_n N_VPWR_c_625_n 0.0124822f $X=4.385 $Y=2.805 $X2=0
+ $Y2=0
cc_393 N_A_27_392#_c_429_n N_A_750_392#_M1002_s 0.00218982f $X=5.975 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_394 N_A_27_392#_c_430_n N_A_750_392#_M1002_s 0.00218982f $X=4.22 $Y=2.99
+ $X2=-0.19 $Y2=-0.245
cc_395 N_A_27_392#_c_429_n N_A_750_392#_M1018_d 0.00165831f $X=5.975 $Y=2.035
+ $X2=0 $Y2=0
cc_396 N_A_27_392#_M1003_d N_A_750_392#_c_747_n 0.00567673f $X=4.25 $Y=1.96
+ $X2=0 $Y2=0
cc_397 N_A_27_392#_c_429_n N_A_750_392#_c_747_n 0.078691f $X=5.975 $Y=2.035
+ $X2=0 $Y2=0
cc_398 N_A_27_392#_c_430_n N_A_750_392#_c_747_n 0.00464895f $X=4.22 $Y=2.99
+ $X2=0 $Y2=0
cc_399 N_A_27_392#_c_437_n N_A_750_392#_c_747_n 0.0211762f $X=4.385 $Y=2.805
+ $X2=0 $Y2=0
cc_400 N_A_27_392#_c_429_n N_A_750_392#_c_750_n 0.0183291f $X=5.975 $Y=2.035
+ $X2=0 $Y2=0
cc_401 N_A_27_392#_c_430_n N_A_750_392#_c_750_n 0.0171805f $X=4.22 $Y=2.99 $X2=0
+ $Y2=0
cc_402 N_A_27_392#_c_429_n N_A_750_392#_c_748_n 0.0171986f $X=5.975 $Y=2.035
+ $X2=0 $Y2=0
cc_403 N_A_27_392#_M1006_g N_X_c_770_n 0.00792144f $X=6.135 $Y=0.74 $X2=0 $Y2=0
cc_404 N_A_27_392#_M1009_g N_X_c_770_n 0.00993385f $X=6.565 $Y=0.74 $X2=0 $Y2=0
cc_405 N_A_27_392#_M1012_g N_X_c_770_n 7.02145e-19 $X=7.135 $Y=0.74 $X2=0 $Y2=0
cc_406 N_A_27_392#_c_411_n N_X_c_785_n 0.00375441f $X=7.245 $Y=1.425 $X2=0 $Y2=0
cc_407 N_A_27_392#_c_565_p N_X_c_785_n 0.0196131f $X=6.96 $Y=1.515 $X2=0 $Y2=0
cc_408 N_A_27_392#_M1015_g N_X_c_779_n 3.02096e-19 $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_409 N_A_27_392#_M1016_g N_X_c_779_n 3.0062e-19 $X=6.705 $Y=2.4 $X2=0 $Y2=0
cc_410 N_A_27_392#_M1009_g N_X_c_771_n 0.0118691f $X=6.565 $Y=0.74 $X2=0 $Y2=0
cc_411 N_A_27_392#_M1012_g N_X_c_771_n 0.0127389f $X=7.135 $Y=0.74 $X2=0 $Y2=0
cc_412 N_A_27_392#_c_411_n N_X_c_771_n 0.00599162f $X=7.245 $Y=1.425 $X2=0 $Y2=0
cc_413 N_A_27_392#_c_565_p N_X_c_771_n 0.0451032f $X=6.96 $Y=1.515 $X2=0 $Y2=0
cc_414 N_A_27_392#_M1006_g N_X_c_772_n 0.00343246f $X=6.135 $Y=0.74 $X2=0 $Y2=0
cc_415 N_A_27_392#_M1009_g N_X_c_772_n 0.00157732f $X=6.565 $Y=0.74 $X2=0 $Y2=0
cc_416 N_A_27_392#_c_411_n N_X_c_772_n 0.00266482f $X=7.245 $Y=1.425 $X2=0 $Y2=0
cc_417 N_A_27_392#_c_565_p N_X_c_772_n 0.0276081f $X=6.96 $Y=1.515 $X2=0 $Y2=0
cc_418 N_A_27_392#_M1016_g N_X_c_797_n 0.0194167f $X=6.705 $Y=2.4 $X2=0 $Y2=0
cc_419 N_A_27_392#_M1017_g N_X_c_797_n 0.0211218f $X=7.155 $Y=2.4 $X2=0 $Y2=0
cc_420 N_A_27_392#_c_411_n N_X_c_797_n 0.00207011f $X=7.245 $Y=1.425 $X2=0 $Y2=0
cc_421 N_A_27_392#_c_565_p N_X_c_797_n 0.0352986f $X=6.96 $Y=1.515 $X2=0 $Y2=0
cc_422 N_A_27_392#_M1009_g N_X_c_773_n 7.02145e-19 $X=6.565 $Y=0.74 $X2=0 $Y2=0
cc_423 N_A_27_392#_M1012_g N_X_c_773_n 0.00993385f $X=7.135 $Y=0.74 $X2=0 $Y2=0
cc_424 N_A_27_392#_M1019_g N_X_c_773_n 0.0145491f $X=7.565 $Y=0.74 $X2=0 $Y2=0
cc_425 N_A_27_392#_c_411_n N_X_c_780_n 0.00440103f $X=7.245 $Y=1.425 $X2=0 $Y2=0
cc_426 N_A_27_392#_M1021_g N_X_c_780_n 0.00922316f $X=7.605 $Y=2.4 $X2=0 $Y2=0
cc_427 N_A_27_392#_c_565_p N_X_c_780_n 0.00234327f $X=6.96 $Y=1.515 $X2=0 $Y2=0
cc_428 N_A_27_392#_M1017_g N_X_c_781_n 3.63823e-19 $X=7.155 $Y=2.4 $X2=0 $Y2=0
cc_429 N_A_27_392#_M1021_g N_X_c_781_n 0.0102677f $X=7.605 $Y=2.4 $X2=0 $Y2=0
cc_430 N_A_27_392#_M1019_g N_X_c_774_n 0.0131828f $X=7.565 $Y=0.74 $X2=0 $Y2=0
cc_431 N_A_27_392#_c_414_n N_X_c_774_n 0.00153079f $X=7.592 $Y=1.425 $X2=0 $Y2=0
cc_432 N_A_27_392#_M1021_g N_X_c_775_n 0.0117327f $X=7.605 $Y=2.4 $X2=0 $Y2=0
cc_433 N_A_27_392#_c_414_n N_X_c_775_n 0.00293976f $X=7.592 $Y=1.425 $X2=0 $Y2=0
cc_434 N_A_27_392#_c_410_n N_X_c_776_n 0.00565298f $X=7.49 $Y=1.425 $X2=0 $Y2=0
cc_435 N_A_27_392#_c_411_n N_X_c_776_n 0.00146733f $X=7.245 $Y=1.425 $X2=0 $Y2=0
cc_436 N_A_27_392#_M1021_g N_X_c_776_n 0.00172267f $X=7.605 $Y=2.4 $X2=0 $Y2=0
cc_437 N_A_27_392#_c_414_n N_X_c_776_n 0.0010485f $X=7.592 $Y=1.425 $X2=0 $Y2=0
cc_438 N_A_27_392#_c_565_p N_X_c_776_n 0.0150643f $X=6.96 $Y=1.515 $X2=0 $Y2=0
cc_439 N_A_27_392#_M1012_g N_X_c_777_n 0.00192507f $X=7.135 $Y=0.74 $X2=0 $Y2=0
cc_440 N_A_27_392#_c_410_n N_X_c_777_n 0.00245515f $X=7.49 $Y=1.425 $X2=0 $Y2=0
cc_441 N_A_27_392#_M1019_g N_X_c_777_n 0.00164391f $X=7.565 $Y=0.74 $X2=0 $Y2=0
cc_442 N_A_27_392#_M1021_g N_X_c_821_n 0.00388982f $X=7.605 $Y=2.4 $X2=0 $Y2=0
cc_443 N_A_27_392#_M1019_g X 0.00602992f $X=7.565 $Y=0.74 $X2=0 $Y2=0
cc_444 N_A_27_392#_c_414_n X 0.0059128f $X=7.592 $Y=1.425 $X2=0 $Y2=0
cc_445 N_A_27_392#_c_417_n N_A_27_74#_c_851_n 0.0131655f $X=0.715 $Y=0.95 $X2=0
+ $Y2=0
cc_446 N_A_27_392#_M1010_d N_A_27_74#_c_852_n 0.00180346f $X=0.575 $Y=0.37 $X2=0
+ $Y2=0
cc_447 N_A_27_392#_c_417_n N_A_27_74#_c_852_n 0.0176997f $X=0.715 $Y=0.95 $X2=0
+ $Y2=0
cc_448 N_A_27_392#_c_417_n N_A_27_74#_c_853_n 0.0142848f $X=0.715 $Y=0.95 $X2=0
+ $Y2=0
cc_449 N_A_27_392#_c_427_n N_A_477_198#_c_918_n 0.00816198f $X=3.22 $Y=2.035
+ $X2=0 $Y2=0
cc_450 N_A_27_392#_c_435_n N_A_477_198#_c_918_n 0.00394735f $X=2.315 $Y=2.105
+ $X2=0 $Y2=0
cc_451 N_A_27_392#_c_427_n N_A_477_198#_c_928_n 0.00481362f $X=3.22 $Y=2.035
+ $X2=0 $Y2=0
cc_452 N_A_27_392#_c_429_n N_A_477_198#_c_921_n 0.0039109f $X=5.975 $Y=2.035
+ $X2=0 $Y2=0
cc_453 N_A_27_392#_c_436_n N_A_477_198#_c_924_n 0.00481287f $X=3.385 $Y=2.115
+ $X2=0 $Y2=0
cc_454 N_A_27_392#_M1006_g N_VGND_c_984_n 0.00590268f $X=6.135 $Y=0.74 $X2=0
+ $Y2=0
cc_455 N_A_27_392#_c_416_n N_VGND_c_984_n 0.00304495f $X=6.145 $Y=1.515 $X2=0
+ $Y2=0
cc_456 N_A_27_392#_M1009_g N_VGND_c_985_n 0.00469226f $X=6.565 $Y=0.74 $X2=0
+ $Y2=0
cc_457 N_A_27_392#_M1012_g N_VGND_c_985_n 0.00469226f $X=7.135 $Y=0.74 $X2=0
+ $Y2=0
cc_458 N_A_27_392#_M1019_g N_VGND_c_987_n 0.0123273f $X=7.565 $Y=0.74 $X2=0
+ $Y2=0
cc_459 N_A_27_392#_M1006_g N_VGND_c_992_n 0.00434272f $X=6.135 $Y=0.74 $X2=0
+ $Y2=0
cc_460 N_A_27_392#_M1009_g N_VGND_c_992_n 0.00434272f $X=6.565 $Y=0.74 $X2=0
+ $Y2=0
cc_461 N_A_27_392#_M1012_g N_VGND_c_995_n 0.00434272f $X=7.135 $Y=0.74 $X2=0
+ $Y2=0
cc_462 N_A_27_392#_M1019_g N_VGND_c_995_n 0.00434272f $X=7.565 $Y=0.74 $X2=0
+ $Y2=0
cc_463 N_A_27_392#_M1006_g N_VGND_c_997_n 0.00820772f $X=6.135 $Y=0.74 $X2=0
+ $Y2=0
cc_464 N_A_27_392#_M1009_g N_VGND_c_997_n 0.00821294f $X=6.565 $Y=0.74 $X2=0
+ $Y2=0
cc_465 N_A_27_392#_M1012_g N_VGND_c_997_n 0.00821294f $X=7.135 $Y=0.74 $X2=0
+ $Y2=0
cc_466 N_A_27_392#_M1019_g N_VGND_c_997_n 0.00824014f $X=7.565 $Y=0.74 $X2=0
+ $Y2=0
cc_467 N_VPWR_M1018_s N_A_750_392#_c_747_n 0.00720599f $X=4.8 $Y=1.96 $X2=0
+ $Y2=0
cc_468 N_VPWR_c_630_n N_A_750_392#_c_747_n 0.0238156f $X=4.945 $Y=2.805 $X2=0
+ $Y2=0
cc_469 N_VPWR_c_630_n N_A_750_392#_c_748_n 0.0139233f $X=4.945 $Y=2.805 $X2=0
+ $Y2=0
cc_470 N_VPWR_c_631_n N_A_750_392#_c_748_n 0.0174579f $X=5.98 $Y=2.455 $X2=0
+ $Y2=0
cc_471 N_VPWR_c_640_n N_A_750_392#_c_748_n 0.0144776f $X=5.815 $Y=3.33 $X2=0
+ $Y2=0
cc_472 N_VPWR_c_625_n N_A_750_392#_c_748_n 0.0118404f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_473 N_VPWR_c_631_n N_X_c_779_n 0.0266594f $X=5.98 $Y=2.455 $X2=0 $Y2=0
cc_474 N_VPWR_c_632_n N_X_c_779_n 0.023849f $X=6.93 $Y=2.435 $X2=0 $Y2=0
cc_475 N_VPWR_c_641_n N_X_c_779_n 0.0121815f $X=6.765 $Y=3.33 $X2=0 $Y2=0
cc_476 N_VPWR_c_625_n N_X_c_779_n 0.0100828f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_477 N_VPWR_M1016_d N_X_c_797_n 0.00317908f $X=6.795 $Y=1.84 $X2=0 $Y2=0
cc_478 N_VPWR_c_632_n N_X_c_797_n 0.0178311f $X=6.93 $Y=2.435 $X2=0 $Y2=0
cc_479 N_VPWR_c_634_n N_X_c_780_n 0.0018333f $X=7.88 $Y=1.985 $X2=0 $Y2=0
cc_480 N_VPWR_c_632_n N_X_c_781_n 0.0214316f $X=6.93 $Y=2.435 $X2=0 $Y2=0
cc_481 N_VPWR_c_634_n N_X_c_781_n 0.0295221f $X=7.88 $Y=1.985 $X2=0 $Y2=0
cc_482 N_VPWR_c_642_n N_X_c_781_n 0.0109793f $X=7.715 $Y=3.33 $X2=0 $Y2=0
cc_483 N_VPWR_c_625_n N_X_c_781_n 0.00901959f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_484 N_VPWR_c_634_n N_X_c_775_n 0.0289318f $X=7.88 $Y=1.985 $X2=0 $Y2=0
cc_485 N_X_c_772_n N_A_477_198#_c_921_n 0.00152173f $X=6.515 $Y=1.095 $X2=0
+ $Y2=0
cc_486 N_X_c_771_n N_VGND_M1009_s 0.00377777f $X=7.185 $Y=1.095 $X2=0 $Y2=0
cc_487 N_X_c_774_n N_VGND_M1019_s 0.0044011f $X=7.805 $Y=1.095 $X2=0 $Y2=0
cc_488 N_X_c_770_n N_VGND_c_984_n 0.0255177f $X=6.35 $Y=0.515 $X2=0 $Y2=0
cc_489 N_X_c_772_n N_VGND_c_984_n 0.00584871f $X=6.515 $Y=1.095 $X2=0 $Y2=0
cc_490 N_X_c_770_n N_VGND_c_985_n 0.0182384f $X=6.35 $Y=0.515 $X2=0 $Y2=0
cc_491 N_X_c_771_n N_VGND_c_985_n 0.0224739f $X=7.185 $Y=1.095 $X2=0 $Y2=0
cc_492 N_X_c_773_n N_VGND_c_985_n 0.0182384f $X=7.35 $Y=0.515 $X2=0 $Y2=0
cc_493 N_X_c_773_n N_VGND_c_987_n 0.0182384f $X=7.35 $Y=0.515 $X2=0 $Y2=0
cc_494 N_X_c_774_n N_VGND_c_987_n 0.0248922f $X=7.805 $Y=1.095 $X2=0 $Y2=0
cc_495 N_X_c_770_n N_VGND_c_992_n 0.0144922f $X=6.35 $Y=0.515 $X2=0 $Y2=0
cc_496 N_X_c_773_n N_VGND_c_995_n 0.0144922f $X=7.35 $Y=0.515 $X2=0 $Y2=0
cc_497 N_X_c_770_n N_VGND_c_997_n 0.0118826f $X=6.35 $Y=0.515 $X2=0 $Y2=0
cc_498 N_X_c_773_n N_VGND_c_997_n 0.0118826f $X=7.35 $Y=0.515 $X2=0 $Y2=0
cc_499 N_A_27_74#_c_856_n N_A_287_74#_M1001_d 0.00176891f $X=1.92 $Y=0.397
+ $X2=-0.19 $Y2=-0.245
cc_500 N_A_27_74#_M1008_s N_A_287_74#_c_889_n 0.00624487f $X=1.865 $Y=0.37 $X2=0
+ $Y2=0
cc_501 N_A_27_74#_c_855_n N_A_287_74#_c_889_n 0.024192f $X=2.085 $Y=0.375 $X2=0
+ $Y2=0
cc_502 N_A_27_74#_c_856_n N_A_287_74#_c_889_n 0.00497069f $X=1.92 $Y=0.397 $X2=0
+ $Y2=0
cc_503 N_A_27_74#_c_853_n N_A_287_74#_c_890_n 0.0204279f $X=1.145 $Y=0.965 $X2=0
+ $Y2=0
cc_504 N_A_27_74#_c_856_n N_A_287_74#_c_890_n 0.0158153f $X=1.92 $Y=0.397 $X2=0
+ $Y2=0
cc_505 N_A_27_74#_c_855_n N_A_287_74#_c_891_n 5.51636e-19 $X=2.085 $Y=0.375
+ $X2=0 $Y2=0
cc_506 N_A_27_74#_c_850_n N_VGND_c_988_n 0.018997f $X=0.247 $Y=0.6 $X2=0 $Y2=0
cc_507 N_A_27_74#_c_852_n N_VGND_c_988_n 0.0450241f $X=1.06 $Y=0.427 $X2=0 $Y2=0
cc_508 N_A_27_74#_c_854_n N_VGND_c_988_n 0.0121867f $X=1.145 $Y=0.515 $X2=0
+ $Y2=0
cc_509 N_A_27_74#_c_856_n N_VGND_c_988_n 0.0658946f $X=1.92 $Y=0.397 $X2=0 $Y2=0
cc_510 N_A_27_74#_M1008_s N_VGND_c_997_n 0.00242558f $X=1.865 $Y=0.37 $X2=0
+ $Y2=0
cc_511 N_A_27_74#_c_850_n N_VGND_c_997_n 0.0103026f $X=0.247 $Y=0.6 $X2=0 $Y2=0
cc_512 N_A_27_74#_c_852_n N_VGND_c_997_n 0.0245954f $X=1.06 $Y=0.427 $X2=0 $Y2=0
cc_513 N_A_27_74#_c_854_n N_VGND_c_997_n 0.00660921f $X=1.145 $Y=0.515 $X2=0
+ $Y2=0
cc_514 N_A_27_74#_c_856_n N_VGND_c_997_n 0.0372424f $X=1.92 $Y=0.397 $X2=0 $Y2=0
cc_515 N_A_287_74#_c_889_n N_A_477_198#_M1004_s 0.00635284f $X=2.875 $Y=0.795
+ $X2=-0.19 $Y2=-0.245
cc_516 N_A_287_74#_c_889_n N_A_477_198#_c_918_n 0.0333166f $X=2.875 $Y=0.795
+ $X2=0 $Y2=0
cc_517 N_A_287_74#_c_890_n N_A_477_198#_c_918_n 0.00246079f $X=1.74 $Y=0.862
+ $X2=0 $Y2=0
cc_518 N_A_287_74#_M1004_d N_A_477_198#_c_928_n 0.00359685f $X=2.9 $Y=0.54 $X2=0
+ $Y2=0
cc_519 N_A_287_74#_c_891_n N_A_477_198#_c_928_n 0.014851f $X=3.04 $Y=0.7 $X2=0
+ $Y2=0
cc_520 N_A_287_74#_c_891_n N_A_477_198#_c_919_n 0.0130934f $X=3.04 $Y=0.7 $X2=0
+ $Y2=0
cc_521 N_A_287_74#_c_889_n N_VGND_c_988_n 0.0089723f $X=2.875 $Y=0.795 $X2=0
+ $Y2=0
cc_522 N_A_287_74#_c_891_n N_VGND_c_988_n 0.00617201f $X=3.04 $Y=0.7 $X2=0 $Y2=0
cc_523 N_A_287_74#_c_889_n N_VGND_c_997_n 0.0178492f $X=2.875 $Y=0.795 $X2=0
+ $Y2=0
cc_524 N_A_287_74#_c_891_n N_VGND_c_997_n 0.00794446f $X=3.04 $Y=0.7 $X2=0 $Y2=0
cc_525 N_A_477_198#_c_938_n N_VGND_M1007_s 0.00444479f $X=4.235 $Y=1.195
+ $X2=-0.19 $Y2=-0.245
cc_526 N_A_477_198#_c_919_n N_VGND_c_982_n 0.0157813f $X=3.47 $Y=0.685 $X2=0
+ $Y2=0
cc_527 N_A_477_198#_c_938_n N_VGND_c_982_n 0.0202152f $X=4.235 $Y=1.195 $X2=0
+ $Y2=0
cc_528 N_A_477_198#_c_920_n N_VGND_c_982_n 0.0165499f $X=4.4 $Y=0.685 $X2=0
+ $Y2=0
cc_529 N_A_477_198#_c_920_n N_VGND_c_983_n 0.0260211f $X=4.4 $Y=0.685 $X2=0
+ $Y2=0
cc_530 N_A_477_198#_c_921_n N_VGND_c_983_n 0.0243991f $X=5.335 $Y=1.195 $X2=0
+ $Y2=0
cc_531 N_A_477_198#_c_922_n N_VGND_c_983_n 0.0218329f $X=5.42 $Y=0.515 $X2=0
+ $Y2=0
cc_532 N_A_477_198#_c_921_n N_VGND_c_984_n 0.00157055f $X=5.335 $Y=1.195 $X2=0
+ $Y2=0
cc_533 N_A_477_198#_c_922_n N_VGND_c_984_n 0.027926f $X=5.42 $Y=0.515 $X2=0
+ $Y2=0
cc_534 N_A_477_198#_c_919_n N_VGND_c_988_n 0.00645818f $X=3.47 $Y=0.685 $X2=0
+ $Y2=0
cc_535 N_A_477_198#_c_922_n N_VGND_c_990_n 0.00749631f $X=5.42 $Y=0.515 $X2=0
+ $Y2=0
cc_536 N_A_477_198#_c_920_n N_VGND_c_994_n 0.00858533f $X=4.4 $Y=0.685 $X2=0
+ $Y2=0
cc_537 N_A_477_198#_c_919_n N_VGND_c_997_n 0.00815448f $X=3.47 $Y=0.685 $X2=0
+ $Y2=0
cc_538 N_A_477_198#_c_920_n N_VGND_c_997_n 0.0108043f $X=4.4 $Y=0.685 $X2=0
+ $Y2=0
cc_539 N_A_477_198#_c_922_n N_VGND_c_997_n 0.0062048f $X=5.42 $Y=0.515 $X2=0
+ $Y2=0

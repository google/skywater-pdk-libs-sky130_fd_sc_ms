* File: sky130_fd_sc_ms__or4bb_1.pex.spice
* Created: Fri Aug 28 18:10:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__OR4BB_1%C_N 3 7 9 13 16
r28 15 16 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.505 $Y=1.465
+ $X2=0.52 $Y2=1.465
r29 12 15 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.29 $Y=1.465
+ $X2=0.505 $Y2=1.465
r30 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.465 $X2=0.29 $Y2=1.465
r31 9 13 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.29 $Y=1.665 $X2=0.29
+ $Y2=1.465
r32 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=1.3 $X2=0.52
+ $Y2=1.465
r33 5 7 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.52 $Y=1.3 $X2=0.52
+ $Y2=0.645
r34 1 15 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=1.465
r35 1 3 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_MS__OR4BB_1%D_N 2 5 9 11 12 15
r48 15 17 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.105 $Y=1.215
+ $X2=1.105 $Y2=1.05
r49 12 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.13
+ $Y=1.215 $X2=1.13 $Y2=1.215
r50 9 17 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=1.09 $Y=0.645
+ $X2=1.09 $Y2=1.05
r51 5 11 318.742 $w=1.8e-07 $l=8.2e-07 $layer=POLY_cond $X=1.005 $Y=2.54
+ $X2=1.005 $Y2=1.72
r52 2 11 43.2981 $w=3.8e-07 $l=1.9e-07 $layer=POLY_cond $X=1.105 $Y=1.53
+ $X2=1.105 $Y2=1.72
r53 1 15 3.65891 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.105 $Y=1.24
+ $X2=1.105 $Y2=1.215
r54 1 2 42.4433 $w=3.8e-07 $l=2.9e-07 $layer=POLY_cond $X=1.105 $Y=1.24
+ $X2=1.105 $Y2=1.53
.ends

.subckt PM_SKY130_FD_SC_MS__OR4BB_1%A_219_424# 1 2 7 9 10 12 14 21 23 27 30 32
+ 33
r66 30 32 8.7366 $w=4.18e-07 $l=1.65e-07 $layer=LI1_cond $X=1.695 $Y=1.195
+ $X2=1.695 $Y2=1.03
r67 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.74
+ $Y=1.195 $X2=1.74 $Y2=1.195
r68 25 27 5.98039 $w=5.28e-07 $l=2.65e-07 $layer=LI1_cond $X=1.305 $Y=0.615
+ $X2=1.57 $Y2=0.615
r69 23 33 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.57 $Y=1.89
+ $X2=1.57 $Y2=1.7
r70 21 33 9.97136 $w=4.18e-07 $l=2.1e-07 $layer=LI1_cond $X=1.695 $Y=1.49
+ $X2=1.695 $Y2=1.7
r71 20 30 1.23476 $w=4.18e-07 $l=4.5e-08 $layer=LI1_cond $X=1.695 $Y=1.24
+ $X2=1.695 $Y2=1.195
r72 20 21 6.85978 $w=4.18e-07 $l=2.5e-07 $layer=LI1_cond $X=1.695 $Y=1.24
+ $X2=1.695 $Y2=1.49
r73 18 27 7.52407 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=1.57 $Y=0.88
+ $X2=1.57 $Y2=0.615
r74 18 32 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.57 $Y=0.88 $X2=1.57
+ $Y2=1.03
r75 14 23 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.485 $Y=2.015
+ $X2=1.57 $Y2=1.89
r76 14 16 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=1.485 $Y=2.015
+ $X2=1.34 $Y2=2.015
r77 10 31 65.9053 $w=6.41e-07 $l=6.15427e-07 $layer=POLY_cond $X=2.155 $Y=1.7
+ $X2=1.91 $Y2=1.195
r78 10 12 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=2.155 $Y=1.7
+ $X2=2.155 $Y2=2.39
r79 7 31 45.6838 $w=6.41e-07 $l=3.01413e-07 $layer=POLY_cond $X=2.14 $Y=1.03
+ $X2=1.91 $Y2=1.195
r80 7 9 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=2.14 $Y=1.03 $X2=2.14
+ $Y2=0.645
r81 2 16 600 $w=1.7e-07 $l=2.7559e-07 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=2.12 $X2=1.34 $Y2=2.055
r82 1 25 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=1.165
+ $Y=0.37 $X2=1.305 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__OR4BB_1%A_27_424# 1 2 9 13 19 22 23 26 27 28 31 32
+ 35 38 41
r97 37 38 6.145 $w=3.78e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=2.29 $X2=0.795
+ $Y2=2.29
r98 35 37 13.0408 $w=3.78e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=2.29
+ $X2=0.71 $Y2=2.29
r99 32 45 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=1.355
+ $X2=2.59 $Y2=1.52
r100 32 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=1.355
+ $X2=2.59 $Y2=1.19
r101 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.59
+ $Y=1.355 $X2=2.59 $Y2=1.355
r102 29 31 54.1299 $w=3.28e-07 $l=1.55e-06 $layer=LI1_cond $X=2.59 $Y=2.905
+ $X2=2.59 $Y2=1.355
r103 27 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.425 $Y=2.99
+ $X2=2.59 $Y2=2.905
r104 27 28 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=2.425 $Y=2.99
+ $X2=1.285 $Y2=2.99
r105 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.2 $Y=2.905
+ $X2=1.285 $Y2=2.99
r106 25 26 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.2 $Y=2.48
+ $X2=1.2 $Y2=2.905
r107 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.115 $Y=2.395
+ $X2=1.2 $Y2=2.48
r108 23 38 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.115 $Y=2.395
+ $X2=0.795 $Y2=2.395
r109 22 37 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.71 $Y=2.1 $X2=0.71
+ $Y2=2.29
r110 21 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=1.13
+ $X2=0.71 $Y2=1.045
r111 21 22 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=0.71 $Y=1.13
+ $X2=0.71 $Y2=2.1
r112 17 41 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.305 $Y=1.045
+ $X2=0.71 $Y2=1.045
r113 17 19 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.305 $Y=0.96
+ $X2=0.305 $Y2=0.645
r114 13 44 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.625 $Y=0.645
+ $X2=2.625 $Y2=1.19
r115 9 45 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=2.575 $Y=2.39
+ $X2=2.575 $Y2=1.52
r116 2 35 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.265
r117 1 19 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.37 $X2=0.305 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__OR4BB_1%B 3 7 9 10 11 12 18 19
r38 18 21 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.13 $Y=1.515
+ $X2=3.13 $Y2=1.68
r39 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.13 $Y=1.515
+ $X2=3.13 $Y2=1.35
r40 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.13
+ $Y=1.515 $X2=3.13 $Y2=1.515
r41 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.13 $Y=2.405
+ $X2=3.13 $Y2=2.775
r42 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.13 $Y=2.035
+ $X2=3.13 $Y2=2.405
r43 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.13 $Y=1.665
+ $X2=3.13 $Y2=2.035
r44 9 19 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.13 $Y=1.665
+ $X2=3.13 $Y2=1.515
r45 7 20 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=3.19 $Y=0.645 $X2=3.19
+ $Y2=1.35
r46 3 21 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=3.055 $Y=2.39
+ $X2=3.055 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__OR4BB_1%A 3 7 9 12 13
c39 7 0 2.01992e-19 $X=3.69 $Y=0.645
r40 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.515
+ $X2=3.67 $Y2=1.68
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.515
+ $X2=3.67 $Y2=1.35
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.67
+ $Y=1.515 $X2=3.67 $Y2=1.515
r43 9 13 4.93904 $w=3.48e-07 $l=1.5e-07 $layer=LI1_cond $X=3.66 $Y=1.665
+ $X2=3.66 $Y2=1.515
r44 7 14 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=3.69 $Y=0.645 $X2=3.69
+ $Y2=1.35
r45 3 15 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=3.595 $Y=2.39
+ $X2=3.595 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__OR4BB_1%A_357_378# 1 2 3 12 16 24 26 30 32 35 36 37
+ 38 44
c94 44 0 3.95737e-20 $X=4.21 $Y=1.465
c95 26 0 1.25867e-19 $X=3.31 $Y=0.935
r96 44 47 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.21 $Y=1.465
+ $X2=4.21 $Y2=1.63
r97 44 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.21 $Y=1.465
+ $X2=4.21 $Y2=1.3
r98 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.21
+ $Y=1.465 $X2=4.21 $Y2=1.465
r99 38 39 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=3.475 $Y=0.935
+ $X2=3.475 $Y2=1.095
r100 35 36 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=2.045 $Y=2.035
+ $X2=2.045 $Y2=1.87
r101 33 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.64 $Y=1.095
+ $X2=3.475 $Y2=1.095
r102 32 43 16.3551 $w=2.76e-07 $l=4.53156e-07 $layer=LI1_cond $X=4.005 $Y=1.095
+ $X2=4.19 $Y2=1.465
r103 32 33 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.005 $Y=1.095
+ $X2=3.64 $Y2=1.095
r104 28 38 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.475 $Y=0.85
+ $X2=3.475 $Y2=0.935
r105 28 30 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=3.475 $Y=0.85
+ $X2=3.475 $Y2=0.645
r106 27 37 2.76166 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=2.575 $Y=0.935
+ $X2=2.325 $Y2=0.935
r107 26 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.31 $Y=0.935
+ $X2=3.475 $Y2=0.935
r108 26 27 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=3.31 $Y=0.935
+ $X2=2.575 $Y2=0.935
r109 22 37 3.70735 $w=2.5e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.41 $Y=0.85
+ $X2=2.325 $Y2=0.935
r110 22 24 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=2.41 $Y=0.85
+ $X2=2.41 $Y2=0.645
r111 20 37 3.70735 $w=2.5e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.16 $Y=1.02
+ $X2=2.325 $Y2=0.935
r112 20 36 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=2.16 $Y=1.02
+ $X2=2.16 $Y2=1.87
r113 16 46 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.295 $Y=0.74
+ $X2=4.295 $Y2=1.3
r114 12 47 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.18 $Y=2.4
+ $X2=4.18 $Y2=1.63
r115 3 35 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.785
+ $Y=1.89 $X2=1.93 $Y2=2.035
r116 2 30 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=3.265
+ $Y=0.37 $X2=3.475 $Y2=0.645
r117 1 24 182 $w=1.7e-07 $l=3.59514e-07 $layer=licon1_NDIFF $count=1 $X=2.215
+ $Y=0.37 $X2=2.41 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__OR4BB_1%VPWR 1 2 9 13 18 19 20 22 35 36 39
r46 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r48 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r49 32 33 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r50 30 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 29 32 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=3.6
+ $Y2=3.33
r52 29 30 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r53 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r54 27 29 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r57 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r58 22 24 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r59 20 33 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=3.6
+ $Y2=3.33
r60 20 30 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r61 18 32 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.74 $Y=3.33 $X2=3.6
+ $Y2=3.33
r62 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.74 $Y=3.33
+ $X2=3.905 $Y2=3.33
r63 17 35 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=4.07 $Y=3.33
+ $X2=4.56 $Y2=3.33
r64 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.07 $Y=3.33
+ $X2=3.905 $Y2=3.33
r65 13 16 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=3.905 $Y=2.115
+ $X2=3.905 $Y2=2.815
r66 11 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.905 $Y=3.245
+ $X2=3.905 $Y2=3.33
r67 11 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.905 $Y=3.245
+ $X2=3.905 $Y2=2.815
r68 7 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245 $X2=0.78
+ $Y2=3.33
r69 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.78 $Y=3.245 $X2=0.78
+ $Y2=2.815
r70 2 16 600 $w=1.7e-07 $l=1.02914e-06 $layer=licon1_PDIFF $count=1 $X=3.685
+ $Y=1.89 $X2=3.905 $Y2=2.815
r71 2 13 300 $w=1.7e-07 $l=3.16425e-07 $layer=licon1_PDIFF $count=2 $X=3.685
+ $Y=1.89 $X2=3.905 $Y2=2.115
r72 1 9 600 $w=1.7e-07 $l=7.82049e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=2.12 $X2=0.78 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__OR4BB_1%X 1 2 9 14 15 16 17 28
c25 17 0 1.15698e-19 $X=4.475 $Y=0.84
r26 21 28 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=4.53 $Y=0.945
+ $X2=4.53 $Y2=0.925
r27 17 30 8.16504 $w=3.68e-07 $l=1.53e-07 $layer=LI1_cond $X=4.53 $Y=0.977
+ $X2=4.53 $Y2=1.13
r28 17 21 0.996707 $w=3.68e-07 $l=3.2e-08 $layer=LI1_cond $X=4.53 $Y=0.977
+ $X2=4.53 $Y2=0.945
r29 17 28 1.02785 $w=3.68e-07 $l=3.3e-08 $layer=LI1_cond $X=4.53 $Y=0.892
+ $X2=4.53 $Y2=0.925
r30 16 17 11.7425 $w=3.68e-07 $l=3.77e-07 $layer=LI1_cond $X=4.53 $Y=0.515
+ $X2=4.53 $Y2=0.892
r31 15 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.63 $Y=1.82 $X2=4.63
+ $Y2=1.13
r32 14 15 9.3668 $w=4.73e-07 $l=1.65e-07 $layer=LI1_cond $X=4.477 $Y=1.985
+ $X2=4.477 $Y2=1.82
r33 7 14 1.813 $w=4.73e-07 $l=7.2e-08 $layer=LI1_cond $X=4.477 $Y=2.057
+ $X2=4.477 $Y2=1.985
r34 7 9 19.0869 $w=4.73e-07 $l=7.58e-07 $layer=LI1_cond $X=4.477 $Y=2.057
+ $X2=4.477 $Y2=2.815
r35 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.27
+ $Y=1.84 $X2=4.405 $Y2=1.985
r36 2 9 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.27
+ $Y=1.84 $X2=4.405 $Y2=2.815
r37 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.37
+ $Y=0.37 $X2=4.51 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR4BB_1%VGND 1 2 3 4 17 21 25 29 32 33 35 36 38 39
+ 40 53 54 57
r66 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r67 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r68 51 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r69 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r70 48 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r71 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r72 45 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r73 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r74 42 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=0 $X2=0.805
+ $Y2=0
r75 42 44 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.97 $Y=0 $X2=1.68
+ $Y2=0
r76 40 48 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r77 40 45 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.68
+ $Y2=0
r78 38 50 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.81 $Y=0 $X2=3.6
+ $Y2=0
r79 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.81 $Y=0 $X2=3.975
+ $Y2=0
r80 37 53 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=4.14 $Y=0 $X2=4.56
+ $Y2=0
r81 37 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.14 $Y=0 $X2=3.975
+ $Y2=0
r82 35 47 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.64
+ $Y2=0
r83 35 36 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.942
+ $Y2=0
r84 34 50 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.14 $Y=0 $X2=3.6
+ $Y2=0
r85 34 36 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=3.14 $Y=0 $X2=2.942
+ $Y2=0
r86 32 44 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.825 $Y=0 $X2=1.68
+ $Y2=0
r87 32 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.825 $Y=0 $X2=1.95
+ $Y2=0
r88 31 47 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.64
+ $Y2=0
r89 31 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.075 $Y=0 $X2=1.95
+ $Y2=0
r90 27 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.975 $Y=0.085
+ $X2=3.975 $Y2=0
r91 27 29 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=3.975 $Y=0.085
+ $X2=3.975 $Y2=0.595
r92 23 36 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.942 $Y=0.085
+ $X2=2.942 $Y2=0
r93 23 25 12.5456 $w=3.93e-07 $l=4.3e-07 $layer=LI1_cond $X=2.942 $Y=0.085
+ $X2=2.942 $Y2=0.515
r94 19 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.95 $Y=0.085
+ $X2=1.95 $Y2=0
r95 19 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=1.95 $Y=0.085
+ $X2=1.95 $Y2=0.515
r96 15 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=0.085
+ $X2=0.805 $Y2=0
r97 15 17 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=0.805 $Y=0.085
+ $X2=0.805 $Y2=0.57
r98 4 29 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=3.765
+ $Y=0.37 $X2=3.975 $Y2=0.595
r99 3 25 182 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.37 $X2=2.94 $Y2=0.515
r100 2 21 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=1.765
+ $Y=0.37 $X2=1.91 $Y2=0.515
r101 1 17 182 $w=1.7e-07 $l=2.93428e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.37 $X2=0.805 $Y2=0.57
.ends


* File: sky130_fd_sc_ms__sdfxtp_4.pex.spice
* Created: Wed Sep  2 12:31:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SDFXTP_4%A_36_74# 1 2 9 13 15 17 19 22 24 28 29 34
+ 42
c94 42 0 1.57125e-19 $X=0.915 $Y=1.825
c95 15 0 1.95114e-19 $X=0.965 $Y=1.69
c96 13 0 5.7257e-20 $X=1.985 $Y=2.64
r97 40 42 10.1561 $w=5.98e-07 $l=1.65e-07 $layer=LI1_cond $X=0.75 $Y=1.825
+ $X2=0.915 $Y2=1.825
r98 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.69 $X2=0.75 $Y2=1.69
r99 38 40 8.5719 $w=5.98e-07 $l=4.3e-07 $layer=LI1_cond $X=0.32 $Y=1.825
+ $X2=0.75 $Y2=1.825
r100 36 38 2.9902 $w=5.98e-07 $l=1.5e-07 $layer=LI1_cond $X=0.17 $Y=1.825
+ $X2=0.32 $Y2=1.825
r101 31 34 4.10641 $w=4.33e-07 $l=1.55e-07 $layer=LI1_cond $X=0.17 $Y=0.567
+ $X2=0.325 $Y2=0.567
r102 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.03
+ $Y=1.635 $X2=2.03 $Y2=1.635
r103 26 28 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=2.03 $Y=1.955
+ $X2=2.03 $Y2=1.635
r104 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.865 $Y=2.04
+ $X2=2.03 $Y2=1.955
r105 24 42 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=1.865 $Y=2.04
+ $X2=0.915 $Y2=2.04
r106 20 38 2.16985 $w=4.7e-07 $l=3e-07 $layer=LI1_cond $X=0.32 $Y=2.125 $X2=0.32
+ $Y2=1.825
r107 20 22 8.65248 $w=4.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.32 $Y=2.125
+ $X2=0.32 $Y2=2.465
r108 19 36 8.31678 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=0.17 $Y=1.525 $X2=0.17
+ $Y2=1.825
r109 18 31 6.29128 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.17 $Y=0.785
+ $X2=0.17 $Y2=0.567
r110 18 19 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.17 $Y=0.785
+ $X2=0.17 $Y2=1.525
r111 16 29 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.03 $Y=1.975
+ $X2=2.03 $Y2=1.635
r112 16 17 37.308 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.03 $Y=1.975
+ $X2=2.03 $Y2=2.14
r113 15 41 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.965 $Y=1.69
+ $X2=0.75 $Y2=1.69
r114 13 17 194.355 $w=1.8e-07 $l=5e-07 $layer=POLY_cond $X=1.985 $Y=2.64
+ $X2=1.985 $Y2=2.14
r115 7 15 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.04 $Y=1.525
+ $X2=0.965 $Y2=1.69
r116 7 9 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=1.04 $Y=1.525
+ $X2=1.04 $Y2=0.58
r117 2 22 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.245
+ $Y=2.32 $X2=0.39 $Y2=2.465
r118 1 34 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=0.18
+ $Y=0.37 $X2=0.325 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_4%SCE 2 3 4 7 9 11 12 14 16 17 19 20 26 29 33
+ 35 38
r80 32 35 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=2.03 $Y=1.065
+ $X2=2.185 $Y2=1.065
r81 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.03
+ $Y=1.065 $X2=2.03 $Y2=1.065
r82 26 33 8.81321 $w=4.73e-07 $l=3.5e-07 $layer=LI1_cond $X=1.68 $Y=1.047
+ $X2=2.03 $Y2=1.047
r83 26 38 4.02225 $w=4.73e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=1.047
+ $X2=1.565 $Y2=1.047
r84 24 29 9.41406 $w=2.56e-07 $l=5e-08 $layer=POLY_cond $X=0.59 $Y=1.12 $X2=0.54
+ $Y2=1.12
r85 23 38 34.0495 $w=3.28e-07 $l=9.75e-07 $layer=LI1_cond $X=0.59 $Y=1.12
+ $X2=1.565 $Y2=1.12
r86 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.12 $X2=0.59 $Y2=1.12
r87 17 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.185 $Y=0.9
+ $X2=2.185 $Y2=1.065
r88 17 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.185 $Y=0.9
+ $X2=2.185 $Y2=0.58
r89 14 16 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.115 $Y=2.245
+ $X2=1.115 $Y2=2.64
r90 13 20 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.705 $Y=2.17
+ $X2=0.615 $Y2=2.17
r91 12 14 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.025 $Y=2.17
+ $X2=1.115 $Y2=2.245
r92 12 13 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.025 $Y=2.17
+ $X2=0.705 $Y2=2.17
r93 9 20 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=0.615 $Y=2.245
+ $X2=0.615 $Y2=2.17
r94 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.615 $Y=2.245
+ $X2=0.615 $Y2=2.64
r95 5 29 15.2686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=0.955
+ $X2=0.54 $Y2=1.12
r96 5 7 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=0.54 $Y=0.955
+ $X2=0.54 $Y2=0.58
r97 3 20 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.525 $Y=2.17 $X2=0.615
+ $Y2=2.17
r98 3 4 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.525 $Y=2.17
+ $X2=0.345 $Y2=2.17
r99 2 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.27 $Y=2.095
+ $X2=0.345 $Y2=2.17
r100 1 29 50.8359 $w=2.56e-07 $l=3.4271e-07 $layer=POLY_cond $X=0.27 $Y=1.285
+ $X2=0.54 $Y2=1.12
r101 1 2 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.27 $Y=1.285 $X2=0.27
+ $Y2=2.095
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_4%D 3 7 9 12 13
c39 12 0 1.57125e-19 $X=1.49 $Y=1.62
r40 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.49 $Y=1.62
+ $X2=1.49 $Y2=1.785
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.49 $Y=1.62
+ $X2=1.49 $Y2=1.455
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.49
+ $Y=1.62 $X2=1.49 $Y2=1.62
r43 9 13 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.2 $Y=1.62 $X2=1.49
+ $Y2=1.62
r44 7 15 332.347 $w=1.8e-07 $l=8.55e-07 $layer=POLY_cond $X=1.535 $Y=2.64
+ $X2=1.535 $Y2=1.785
r45 3 14 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=1.43 $Y=0.58 $X2=1.43
+ $Y2=1.455
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_4%SCD 3 7 9 10 14
c45 9 0 5.7257e-20 $X=2.64 $Y=1.665
c46 7 0 2.97692e-19 $X=2.575 $Y=0.58
r47 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.6 $Y=1.775
+ $X2=2.6 $Y2=1.94
r48 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.6 $Y=1.775
+ $X2=2.6 $Y2=1.61
r49 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.6
+ $Y=1.775 $X2=2.6 $Y2=1.775
r50 10 15 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.6 $Y=2.035 $X2=2.6
+ $Y2=1.775
r51 9 15 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=2.6 $Y=1.665 $X2=2.6
+ $Y2=1.775
r52 7 16 528.149 $w=1.5e-07 $l=1.03e-06 $layer=POLY_cond $X=2.575 $Y=0.58
+ $X2=2.575 $Y2=1.61
r53 3 17 272.097 $w=1.8e-07 $l=7e-07 $layer=POLY_cond $X=2.525 $Y=2.64 $X2=2.525
+ $Y2=1.94
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_4%CLK 1 3 6 8 11
c43 8 0 9.81103e-20 $X=3.6 $Y=1.295
c44 6 0 6.78871e-20 $X=3.265 $Y=2.4
r45 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.44
+ $Y=1.385 $X2=3.44 $Y2=1.385
r46 11 13 30.4513 $w=2.77e-07 $l=1.75e-07 $layer=POLY_cond $X=3.265 $Y=1.385
+ $X2=3.44 $Y2=1.385
r47 8 14 4.98354 $w=3.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.6 $Y=1.365 $X2=3.44
+ $Y2=1.365
r48 4 11 12.8788 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.265 $Y=1.55
+ $X2=3.265 $Y2=1.385
r49 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.265 $Y=1.55
+ $X2=3.265 $Y2=2.4
r50 1 11 33.0614 $w=2.77e-07 $l=2.59711e-07 $layer=POLY_cond $X=3.075 $Y=1.22
+ $X2=3.265 $Y2=1.385
r51 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.075 $Y=1.22 $X2=3.075
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_4%A_828_74# 1 2 9 11 13 16 20 24 26 27 29 30
+ 33 36 37 39 42 43 44 46 47 54 55 56 59 62 63 67
c191 67 0 7.63119e-20 $X=8.7 $Y=1.55
c192 59 0 1.06925e-20 $X=7.8 $Y=1.22
c193 54 0 6.02966e-20 $X=5.24 $Y=2.205
c194 33 0 1.815e-19 $X=5.86 $Y=0.77
r195 67 80 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.7 $Y=1.55
+ $X2=8.7 $Y2=1.715
r196 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.7
+ $Y=1.55 $X2=8.7 $Y2=1.55
r197 63 66 8.36451 $w=3.08e-07 $l=2.25e-07 $layer=LI1_cond $X=8.69 $Y=1.325
+ $X2=8.69 $Y2=1.55
r198 59 76 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.8 $Y=1.22
+ $X2=7.8 $Y2=1.055
r199 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.8
+ $Y=1.22 $X2=7.8 $Y2=1.22
r200 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.24
+ $Y=2.205 $X2=5.24 $Y2=2.205
r201 47 63 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=8.535 $Y=1.325
+ $X2=8.69 $Y2=1.325
r202 47 62 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=8.535 $Y=1.325
+ $X2=8.125 $Y2=1.325
r203 46 62 5.902 $w=3.53e-07 $l=8.5e-08 $layer=LI1_cond $X=8.04 $Y=1.232
+ $X2=8.125 $Y2=1.232
r204 46 58 7.79116 $w=3.53e-07 $l=2.4e-07 $layer=LI1_cond $X=8.04 $Y=1.232
+ $X2=7.8 $Y2=1.232
r205 45 46 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.04 $Y=0.465
+ $X2=8.04 $Y2=1.055
r206 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.955 $Y=0.38
+ $X2=8.04 $Y2=0.465
r207 43 44 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=7.955 $Y=0.38
+ $X2=7.16 $Y2=0.38
r208 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.075 $Y=0.465
+ $X2=7.16 $Y2=0.38
r209 41 42 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.075 $Y=0.465
+ $X2=7.075 $Y2=0.77
r210 40 56 2.53056 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.075 $Y=0.855
+ $X2=5.925 $Y2=0.855
r211 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.99 $Y=0.855
+ $X2=7.075 $Y2=0.77
r212 39 40 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=6.99 $Y=0.855
+ $X2=6.075 $Y2=0.855
r213 37 71 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=5.91 $Y=1.195
+ $X2=5.735 $Y2=1.195
r214 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.91
+ $Y=1.195 $X2=5.91 $Y2=1.195
r215 34 56 3.91525 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=5.925 $Y=0.94
+ $X2=5.925 $Y2=0.855
r216 34 36 9.79577 $w=2.98e-07 $l=2.55e-07 $layer=LI1_cond $X=5.925 $Y=0.94
+ $X2=5.925 $Y2=1.195
r217 33 56 3.91525 $w=2.35e-07 $l=1.12916e-07 $layer=LI1_cond $X=5.86 $Y=0.77
+ $X2=5.925 $Y2=0.855
r218 32 33 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.86 $Y=0.425
+ $X2=5.86 $Y2=0.77
r219 31 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.265 $Y=0.34
+ $X2=5.18 $Y2=0.34
r220 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.775 $Y=0.34
+ $X2=5.86 $Y2=0.425
r221 30 31 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.775 $Y=0.34
+ $X2=5.265 $Y2=0.34
r222 29 53 2.26625 $w=3.23e-07 $l=6e-08 $layer=LI1_cond $X=5.18 $Y=2.095
+ $X2=5.24 $Y2=2.095
r223 29 50 15.8638 $w=3.23e-07 $l=4.2e-07 $layer=LI1_cond $X=5.18 $Y=2.095
+ $X2=4.76 $Y2=2.095
r224 28 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.18 $Y=0.425
+ $X2=5.18 $Y2=0.34
r225 28 29 105.364 $w=1.68e-07 $l=1.615e-06 $layer=LI1_cond $X=5.18 $Y=0.425
+ $X2=5.18 $Y2=2.04
r226 26 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.095 $Y=0.34
+ $X2=5.18 $Y2=0.34
r227 26 27 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.095 $Y=0.34
+ $X2=4.445 $Y2=0.34
r228 22 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.32 $Y=0.425
+ $X2=4.445 $Y2=0.34
r229 22 24 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.32 $Y=0.425
+ $X2=4.32 $Y2=0.515
r230 20 80 340.121 $w=1.8e-07 $l=8.75e-07 $layer=POLY_cond $X=8.745 $Y=2.59
+ $X2=8.745 $Y2=1.715
r231 16 76 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=7.86 $Y=0.645
+ $X2=7.86 $Y2=1.055
r232 11 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.735 $Y=1.03
+ $X2=5.735 $Y2=1.195
r233 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.735 $Y=1.03
+ $X2=5.735 $Y2=0.71
r234 7 54 57.4258 $w=2.56e-07 $l=3.78616e-07 $layer=POLY_cond $X=5.545 $Y=2.37
+ $X2=5.24 $Y2=2.205
r235 7 9 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=5.545 $Y=2.37
+ $X2=5.545 $Y2=2.74
r236 2 50 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=4.625
+ $Y=1.84 $X2=4.76 $Y2=2.02
r237 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.14
+ $Y=0.37 $X2=4.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_4%A_630_74# 1 2 9 11 15 17 21 23 29 33 36 37
+ 38 41 43 44 47 48 51 53 54 55 59 62 63 65 66 67 69 70 75 78 80 83 94
c206 80 0 6.02966e-20 $X=6.19 $Y=2.115
c207 67 0 1.65237e-19 $X=6.275 $Y=2.6
c208 55 0 6.78871e-20 $X=3.855 $Y=1.905
c209 51 0 1.99582e-19 $X=3.29 $Y=0.515
c210 44 0 1.68504e-19 $X=5.055 $Y=1.555
c211 41 0 8.3449e-20 $X=8.755 $Y=0.58
c212 37 0 1.81826e-20 $X=8.68 $Y=1.07
c213 21 0 1.815e-19 $X=5.055 $Y=0.71
r214 83 86 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.935 $Y=1.79
+ $X2=7.935 $Y2=1.955
r215 83 84 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.935
+ $Y=1.79 $X2=7.935 $Y2=1.79
r216 78 94 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.07 $Y=2.115
+ $X2=6.07 $Y2=2.28
r217 77 80 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=6.07 $Y=2.115
+ $X2=6.19 $Y2=2.115
r218 77 78 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.07
+ $Y=2.115 $X2=6.07 $Y2=2.115
r219 70 73 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.49 $Y=1.905
+ $X2=3.49 $Y2=2.02
r220 69 86 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.015 $Y=2.515
+ $X2=8.015 $Y2=1.955
r221 66 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.93 $Y=2.6
+ $X2=8.015 $Y2=2.515
r222 66 67 107.973 $w=1.68e-07 $l=1.655e-06 $layer=LI1_cond $X=7.93 $Y=2.6
+ $X2=6.275 $Y2=2.6
r223 65 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.19 $Y=2.515
+ $X2=6.275 $Y2=2.6
r224 64 80 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.19 $Y=2.28
+ $X2=6.19 $Y2=2.115
r225 64 65 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.19 $Y=2.28
+ $X2=6.19 $Y2=2.515
r226 63 91 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.01 $Y=1.465
+ $X2=4.01 $Y2=1.555
r227 63 90 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.01 $Y=1.465
+ $X2=4.01 $Y2=1.3
r228 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.01
+ $Y=1.465 $X2=4.01 $Y2=1.465
r229 60 62 13.1973 $w=3.08e-07 $l=3.55e-07 $layer=LI1_cond $X=4.01 $Y=1.82
+ $X2=4.01 $Y2=1.465
r230 59 75 8.09553 $w=3.08e-07 $l=1.55e-07 $layer=LI1_cond $X=4.01 $Y=1.455
+ $X2=4.01 $Y2=1.3
r231 59 62 0.371756 $w=3.08e-07 $l=1e-08 $layer=LI1_cond $X=4.01 $Y=1.455
+ $X2=4.01 $Y2=1.465
r232 57 75 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.94 $Y=1.01
+ $X2=3.94 $Y2=1.3
r233 56 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.655 $Y=1.905
+ $X2=3.49 $Y2=1.905
r234 55 60 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=3.855 $Y=1.905
+ $X2=4.01 $Y2=1.82
r235 55 56 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.855 $Y=1.905
+ $X2=3.655 $Y2=1.905
r236 53 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.855 $Y=0.925
+ $X2=3.94 $Y2=1.01
r237 53 54 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.855 $Y=0.925
+ $X2=3.455 $Y2=0.925
r238 49 54 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.29 $Y=0.84
+ $X2=3.455 $Y2=0.925
r239 49 51 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.29 $Y=0.84
+ $X2=3.29 $Y2=0.515
r240 47 84 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=8.115 $Y=1.79
+ $X2=7.935 $Y2=1.79
r241 47 48 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.115 $Y=1.79
+ $X2=8.115 $Y2=1.625
r242 44 45 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=5.055 $Y=1.555
+ $X2=5.055 $Y2=1.755
r243 39 41 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=8.755 $Y=0.995
+ $X2=8.755 $Y2=0.58
r244 37 39 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.68 $Y=1.07
+ $X2=8.755 $Y2=0.995
r245 37 38 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=8.68 $Y=1.07
+ $X2=8.325 $Y2=1.07
r246 36 48 34.7346 $w=1.65e-07 $l=1.35e-07 $layer=POLY_cond $X=8.25 $Y=1.625
+ $X2=8.115 $Y2=1.625
r247 35 38 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.25 $Y=1.145
+ $X2=8.325 $Y2=1.07
r248 35 36 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.25 $Y=1.145
+ $X2=8.25 $Y2=1.625
r249 31 48 34.7346 $w=1.65e-07 $l=3.7229e-07 $layer=POLY_cond $X=8.205 $Y=1.955
+ $X2=8.115 $Y2=1.625
r250 31 33 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=8.205 $Y=1.955
+ $X2=8.205 $Y2=2.535
r251 29 94 178.806 $w=1.8e-07 $l=4.6e-07 $layer=POLY_cond $X=5.995 $Y=2.74
+ $X2=5.995 $Y2=2.28
r252 25 78 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=6.07 $Y=1.83
+ $X2=6.07 $Y2=2.115
r253 24 45 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.13 $Y=1.755
+ $X2=5.055 $Y2=1.755
r254 23 25 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.905 $Y=1.755
+ $X2=6.07 $Y2=1.83
r255 23 24 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=5.905 $Y=1.755
+ $X2=5.13 $Y2=1.755
r256 19 44 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.055 $Y=1.48
+ $X2=5.055 $Y2=1.555
r257 19 21 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=5.055 $Y=1.48
+ $X2=5.055 $Y2=0.71
r258 18 43 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.625 $Y=1.555
+ $X2=4.535 $Y2=1.555
r259 17 44 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.98 $Y=1.555
+ $X2=5.055 $Y2=1.555
r260 17 18 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=4.98 $Y=1.555
+ $X2=4.625 $Y2=1.555
r261 13 43 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.535 $Y=1.63
+ $X2=4.535 $Y2=1.555
r262 13 15 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.535 $Y=1.63
+ $X2=4.535 $Y2=2.4
r263 12 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.175 $Y=1.555
+ $X2=4.01 $Y2=1.555
r264 11 43 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.445 $Y=1.555
+ $X2=4.535 $Y2=1.555
r265 11 12 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.445 $Y=1.555
+ $X2=4.175 $Y2=1.555
r266 9 90 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.065 $Y=0.74
+ $X2=4.065 $Y2=1.3
r267 2 73 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=3.355
+ $Y=1.84 $X2=3.49 $Y2=2.02
r268 1 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.15
+ $Y=0.37 $X2=3.29 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_4%A_1257_74# 1 2 9 13 15 21 23 25 29 31 35
r72 26 29 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=7.415 $Y=0.76
+ $X2=7.555 $Y2=0.76
r73 23 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.415 $Y=2.175
+ $X2=7.415 $Y2=2.26
r74 22 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.415 $Y=1.44
+ $X2=7.415 $Y2=1.275
r75 22 23 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=7.415 $Y=1.44
+ $X2=7.415 $Y2=2.175
r76 21 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.415 $Y=1.11
+ $X2=7.415 $Y2=1.275
r77 20 26 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.415 $Y=0.885
+ $X2=7.415 $Y2=0.76
r78 20 21 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.415 $Y=0.885
+ $X2=7.415 $Y2=1.11
r79 18 35 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.46 $Y=1.275
+ $X2=6.535 $Y2=1.275
r80 18 32 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=6.46 $Y=1.275 $X2=6.36
+ $Y2=1.275
r81 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.46
+ $Y=1.275 $X2=6.46 $Y2=1.275
r82 15 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.33 $Y=1.275
+ $X2=7.415 $Y2=1.275
r83 15 17 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=7.33 $Y=1.275
+ $X2=6.46 $Y2=1.275
r84 11 35 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.535 $Y=1.44
+ $X2=6.535 $Y2=1.275
r85 11 13 505.323 $w=1.8e-07 $l=1.3e-06 $layer=POLY_cond $X=6.535 $Y=1.44
+ $X2=6.535 $Y2=2.74
r86 7 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.36 $Y=1.11
+ $X2=6.36 $Y2=1.275
r87 7 9 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=6.36 $Y=1.11 $X2=6.36
+ $Y2=0.71
r88 2 25 600 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_PDIFF $count=1 $X=7.245
+ $Y=2.115 $X2=7.485 $Y2=2.26
r89 1 29 182 $w=1.7e-07 $l=4.38748e-07 $layer=licon1_NDIFF $count=1 $X=7.355
+ $Y=0.37 $X2=7.555 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_4%A_1026_100# 1 2 9 13 17 21 22 27 28 39
c81 22 0 1.3178e-19 $X=5.745 $Y=1.695
r82 38 39 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=7.155 $Y=1.775
+ $X2=7.28 $Y2=1.775
r83 34 38 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=7 $Y=1.775
+ $X2=7.155 $Y2=1.775
r84 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7 $Y=1.775
+ $X2=7 $Y2=1.775
r85 27 28 10.5918 $w=3.58e-07 $l=2.3e-07 $layer=LI1_cond $X=5.755 $Y=2.74
+ $X2=5.755 $Y2=2.51
r86 23 25 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.52 $Y=1.695
+ $X2=5.66 $Y2=1.695
r87 22 25 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.745 $Y=1.695
+ $X2=5.66 $Y2=1.695
r88 21 33 2.83678 $w=3.23e-07 $l=8e-08 $layer=LI1_cond $X=6.997 $Y=1.695
+ $X2=6.997 $Y2=1.775
r89 21 22 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=6.835 $Y=1.695
+ $X2=5.745 $Y2=1.695
r90 19 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.66 $Y=1.78
+ $X2=5.66 $Y2=1.695
r91 19 28 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.66 $Y=1.78
+ $X2=5.66 $Y2=2.51
r92 15 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.52 $Y=1.61
+ $X2=5.52 $Y2=1.695
r93 15 17 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=5.52 $Y=1.61
+ $X2=5.52 $Y2=0.765
r94 11 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.28 $Y=1.61
+ $X2=7.28 $Y2=1.775
r95 11 13 494.819 $w=1.5e-07 $l=9.65e-07 $layer=POLY_cond $X=7.28 $Y=1.61
+ $X2=7.28 $Y2=0.645
r96 7 38 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.155 $Y=1.94
+ $X2=7.155 $Y2=1.775
r97 7 9 231.282 $w=1.8e-07 $l=5.95e-07 $layer=POLY_cond $X=7.155 $Y=1.94
+ $X2=7.155 $Y2=2.535
r98 2 27 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=5.635
+ $Y=2.53 $X2=5.77 $Y2=2.74
r99 1 17 182 $w=1.7e-07 $l=5.05421e-07 $layer=licon1_NDIFF $count=1 $X=5.13
+ $Y=0.5 $X2=5.52 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_4%A_1814_48# 1 2 7 9 10 12 18 22 26 30 34 38
+ 42 46 49 50 55 59 64 69 73 74 87
c152 74 0 1.73925e-19 $X=9.932 $Y=1.97
c153 59 0 2.26236e-19 $X=10.135 $Y=1.465
c154 10 0 6.75189e-20 $X=9.165 $Y=1.475
r155 86 87 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=11.975 $Y=1.465
+ $X2=11.985 $Y2=1.465
r156 85 86 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=11.555 $Y=1.465
+ $X2=11.975 $Y2=1.465
r157 84 85 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=11.525 $Y=1.465
+ $X2=11.555 $Y2=1.465
r158 81 82 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=11.075 $Y=1.465
+ $X2=11.125 $Y2=1.465
r159 77 79 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=10.61 $Y=1.465
+ $X2=10.625 $Y2=1.465
r160 73 74 8.6688 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=9.932 $Y=2.135
+ $X2=9.932 $Y2=1.97
r161 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.5
+ $Y=1.065 $X2=9.5 $Y2=1.065
r162 65 84 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=11.38 $Y=1.465
+ $X2=11.525 $Y2=1.465
r163 65 82 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=11.38 $Y=1.465
+ $X2=11.125 $Y2=1.465
r164 64 65 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=11.38
+ $Y=1.465 $X2=11.38 $Y2=1.465
r165 62 81 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=10.7 $Y=1.465
+ $X2=11.075 $Y2=1.465
r166 62 79 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=10.7 $Y=1.465
+ $X2=10.625 $Y2=1.465
r167 61 64 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=10.7 $Y=1.465
+ $X2=11.38 $Y2=1.465
r168 61 62 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=10.7
+ $Y=1.465 $X2=10.7 $Y2=1.465
r169 59 71 3.11411 $w=3.33e-07 $l=2.38747e-07 $layer=LI1_cond $X=10.135 $Y=1.465
+ $X2=10.05 $Y2=1.265
r170 59 61 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=10.135 $Y=1.465
+ $X2=10.7 $Y2=1.465
r171 57 71 4.67747 $w=1.7e-07 $l=3.65e-07 $layer=LI1_cond $X=10.05 $Y=1.63
+ $X2=10.05 $Y2=1.265
r172 57 74 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=10.05 $Y=1.63
+ $X2=10.05 $Y2=1.97
r173 53 71 4.76276 $w=3.33e-07 $l=1.3e-07 $layer=LI1_cond $X=9.92 $Y=1.265
+ $X2=10.05 $Y2=1.265
r174 53 68 15.3874 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=9.92 $Y=1.265
+ $X2=9.5 $Y2=1.265
r175 53 55 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=9.92 $Y=1.13
+ $X2=9.92 $Y2=0.515
r176 48 69 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=9.255 $Y=1.065
+ $X2=9.5 $Y2=1.065
r177 48 49 5.03009 $w=3.3e-07 $l=2.5446e-07 $layer=POLY_cond $X=9.255 $Y=1.065
+ $X2=9.07 $Y2=0.9
r178 44 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.985 $Y=1.3
+ $X2=11.985 $Y2=1.465
r179 44 46 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.985 $Y=1.3
+ $X2=11.985 $Y2=0.74
r180 40 86 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=11.975 $Y=1.63
+ $X2=11.975 $Y2=1.465
r181 40 42 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=11.975 $Y=1.63
+ $X2=11.975 $Y2=2.4
r182 36 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.555 $Y=1.3
+ $X2=11.555 $Y2=1.465
r183 36 38 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.555 $Y=1.3
+ $X2=11.555 $Y2=0.74
r184 32 84 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=11.525 $Y=1.63
+ $X2=11.525 $Y2=1.465
r185 32 34 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=11.525 $Y=1.63
+ $X2=11.525 $Y2=2.4
r186 28 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.125 $Y=1.3
+ $X2=11.125 $Y2=1.465
r187 28 30 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.125 $Y=1.3
+ $X2=11.125 $Y2=0.74
r188 24 81 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=11.075 $Y=1.63
+ $X2=11.075 $Y2=1.465
r189 24 26 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=11.075 $Y=1.63
+ $X2=11.075 $Y2=2.4
r190 20 79 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.625 $Y=1.63
+ $X2=10.625 $Y2=1.465
r191 20 22 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=10.625 $Y=1.63
+ $X2=10.625 $Y2=2.4
r192 16 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.61 $Y=1.3
+ $X2=10.61 $Y2=1.465
r193 16 18 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=10.61 $Y=1.3
+ $X2=10.61 $Y2=0.74
r194 14 49 37.0704 $w=1.5e-07 $l=3.81051e-07 $layer=POLY_cond $X=9.18 $Y=1.23
+ $X2=9.07 $Y2=0.9
r195 14 50 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=9.18 $Y=1.23
+ $X2=9.18 $Y2=1.385
r196 10 50 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=9.165 $Y=1.475
+ $X2=9.165 $Y2=1.385
r197 10 12 433.411 $w=1.8e-07 $l=1.115e-06 $layer=POLY_cond $X=9.165 $Y=1.475
+ $X2=9.165 $Y2=2.59
r198 7 49 37.0704 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.145 $Y=0.9
+ $X2=9.07 $Y2=0.9
r199 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.145 $Y=0.9
+ $X2=9.145 $Y2=0.58
r200 2 73 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=9.76
+ $Y=1.96 $X2=9.895 $Y2=2.135
r201 1 55 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=9.775
+ $Y=0.37 $X2=9.92 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_4%A_1587_74# 1 2 9 11 15 19 21 24 28 30 31 32
+ 33 35 37 40 43 44
c112 43 0 6.75189e-20 $X=9.1 $Y=1.635
c113 33 0 8.70044e-20 $X=8.625 $Y=0.985
c114 15 0 1.24604e-19 $X=10.12 $Y=2.38
r115 41 47 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.63 $Y=1.635
+ $X2=9.63 $Y2=1.8
r116 41 44 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.63 $Y=1.635
+ $X2=9.63 $Y2=1.545
r117 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.63
+ $Y=1.635 $X2=9.63 $Y2=1.635
r118 38 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.185 $Y=1.635
+ $X2=9.1 $Y2=1.635
r119 38 40 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=9.185 $Y=1.635
+ $X2=9.63 $Y2=1.635
r120 36 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.1 $Y=1.8 $X2=9.1
+ $Y2=1.635
r121 36 37 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=9.1 $Y=1.8 $X2=9.1
+ $Y2=2.02
r122 35 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.1 $Y=1.47 $X2=9.1
+ $Y2=1.635
r123 34 35 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=9.1 $Y=1.07 $X2=9.1
+ $Y2=1.47
r124 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.015 $Y=0.985
+ $X2=9.1 $Y2=1.07
r125 32 33 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=9.015 $Y=0.985
+ $X2=8.625 $Y2=0.985
r126 30 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.015 $Y=2.105
+ $X2=9.1 $Y2=2.02
r127 30 31 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=9.015 $Y=2.105
+ $X2=8.6 $Y2=2.105
r128 26 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.46 $Y=0.9
+ $X2=8.625 $Y2=0.985
r129 26 28 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=8.46 $Y=0.9
+ $X2=8.46 $Y2=0.615
r130 22 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.435 $Y=2.19
+ $X2=8.6 $Y2=2.105
r131 22 24 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=8.435 $Y=2.19
+ $X2=8.435 $Y2=2.26
r132 17 21 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=10.135 $Y=1.47
+ $X2=10.12 $Y2=1.545
r133 17 19 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=10.135 $Y=1.47
+ $X2=10.135 $Y2=0.74
r134 13 21 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=10.12 $Y=1.62
+ $X2=10.12 $Y2=1.545
r135 13 15 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=10.12 $Y=1.62
+ $X2=10.12 $Y2=2.38
r136 12 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.795 $Y=1.545
+ $X2=9.63 $Y2=1.545
r137 11 21 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=10.03 $Y=1.545
+ $X2=10.12 $Y2=1.545
r138 11 12 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=10.03 $Y=1.545
+ $X2=9.795 $Y2=1.545
r139 9 47 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=9.67 $Y=2.38
+ $X2=9.67 $Y2=1.8
r140 2 24 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=8.295
+ $Y=2.115 $X2=8.435 $Y2=2.26
r141 1 28 182 $w=1.7e-07 $l=6.35807e-07 $layer=licon1_NDIFF $count=1 $X=7.935
+ $Y=0.37 $X2=8.46 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_4%VPWR 1 2 3 4 5 6 7 8 27 31 35 37 41 43 47
+ 49 51 54 55 56 62 66 71 79 84 90 99 106 109 112 115 119
c147 27 0 1.95114e-19 $X=0.89 $Y=2.465
r148 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r149 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r150 113 116 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r151 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r152 110 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r153 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r154 106 107 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r155 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r156 99 102 10.4403 $w=5.88e-07 $l=5.15e-07 $layer=LI1_cond $X=4.18 $Y=2.815
+ $X2=4.18 $Y2=3.33
r157 94 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r158 93 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r159 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r160 90 93 9.93517 $w=6.18e-07 $l=5.15e-07 $layer=LI1_cond $X=2.895 $Y=2.815
+ $X2=2.895 $Y2=3.33
r161 88 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r162 88 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=11.28 $Y2=3.33
r163 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r164 85 115 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.465 $Y=3.33
+ $X2=11.34 $Y2=3.33
r165 85 87 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=11.465 $Y=3.33
+ $X2=11.76 $Y2=3.33
r166 84 118 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=12.035 $Y=3.33
+ $X2=12.257 $Y2=3.33
r167 84 87 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=12.035 $Y=3.33
+ $X2=11.76 $Y2=3.33
r168 83 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r169 83 107 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=6.96 $Y2=3.33
r170 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r171 80 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.01 $Y=3.33
+ $X2=6.845 $Y2=3.33
r172 80 82 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=7.01 $Y=3.33 $X2=8.88
+ $Y2=3.33
r173 79 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.225 $Y=3.33
+ $X2=9.39 $Y2=3.33
r174 79 82 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.225 $Y=3.33
+ $X2=8.88 $Y2=3.33
r175 78 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r176 77 78 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r177 75 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r178 74 77 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r179 74 75 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r180 72 102 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=4.475 $Y=3.33
+ $X2=4.18 $Y2=3.33
r181 72 74 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.475 $Y=3.33
+ $X2=4.56 $Y2=3.33
r182 71 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.68 $Y=3.33
+ $X2=6.845 $Y2=3.33
r183 71 77 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=6.68 $Y=3.33 $X2=6.48
+ $Y2=3.33
r184 70 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r185 70 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r186 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r187 67 93 8.52869 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=3.205 $Y=3.33
+ $X2=2.895 $Y2=3.33
r188 67 69 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.205 $Y=3.33
+ $X2=3.6 $Y2=3.33
r189 66 102 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=3.885 $Y=3.33
+ $X2=4.18 $Y2=3.33
r190 66 69 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.885 $Y=3.33
+ $X2=3.6 $Y2=3.33
r191 65 94 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r192 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r193 62 93 8.52869 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=2.585 $Y=3.33
+ $X2=2.895 $Y2=3.33
r194 62 64 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=2.585 $Y=3.33
+ $X2=1.2 $Y2=3.33
r195 60 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r196 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r197 56 78 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.24 $Y=3.33
+ $X2=6.48 $Y2=3.33
r198 56 75 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.24 $Y=3.33
+ $X2=4.56 $Y2=3.33
r199 54 59 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.72 $Y2=3.33
r200 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.89 $Y2=3.33
r201 53 64 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.2 $Y2=3.33
r202 53 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.89 $Y2=3.33
r203 49 118 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=12.2 $Y=3.245
+ $X2=12.257 $Y2=3.33
r204 49 51 34.0495 $w=3.28e-07 $l=9.75e-07 $layer=LI1_cond $X=12.2 $Y=3.245
+ $X2=12.2 $Y2=2.27
r205 45 115 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.34 $Y=3.245
+ $X2=11.34 $Y2=3.33
r206 45 47 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=11.34 $Y=3.245
+ $X2=11.34 $Y2=2.305
r207 44 112 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.475 $Y=3.33
+ $X2=10.39 $Y2=3.33
r208 43 115 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.215 $Y=3.33
+ $X2=11.34 $Y2=3.33
r209 43 44 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=11.215 $Y=3.33
+ $X2=10.475 $Y2=3.33
r210 39 112 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.39 $Y=3.245
+ $X2=10.39 $Y2=3.33
r211 39 41 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=10.39 $Y=3.245
+ $X2=10.39 $Y2=2.105
r212 38 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.555 $Y=3.33
+ $X2=9.39 $Y2=3.33
r213 37 112 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.305 $Y=3.33
+ $X2=10.39 $Y2=3.33
r214 37 38 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=10.305 $Y=3.33
+ $X2=9.555 $Y2=3.33
r215 33 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.39 $Y=3.245
+ $X2=9.39 $Y2=3.33
r216 33 35 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=9.39 $Y=3.245
+ $X2=9.39 $Y2=2.59
r217 29 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.845 $Y=3.245
+ $X2=6.845 $Y2=3.33
r218 29 31 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=6.845 $Y=3.245
+ $X2=6.845 $Y2=3.02
r219 25 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=3.245
+ $X2=0.89 $Y2=3.33
r220 25 27 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=0.89 $Y=3.245
+ $X2=0.89 $Y2=2.465
r221 8 51 300 $w=1.7e-07 $l=4.929e-07 $layer=licon1_PDIFF $count=2 $X=12.065
+ $Y=1.84 $X2=12.2 $Y2=2.27
r222 7 47 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=11.165
+ $Y=1.84 $X2=11.3 $Y2=2.305
r223 6 41 300 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=2 $X=10.21
+ $Y=1.96 $X2=10.39 $Y2=2.105
r224 5 35 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=9.255
+ $Y=2.38 $X2=9.39 $Y2=2.59
r225 4 31 600 $w=1.7e-07 $l=5.89831e-07 $layer=licon1_PDIFF $count=1 $X=6.625
+ $Y=2.53 $X2=6.845 $Y2=3.02
r226 3 99 600 $w=1.7e-07 $l=1.10397e-06 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=1.84 $X2=4.18 $Y2=2.815
r227 2 90 600 $w=1.7e-07 $l=6.19375e-07 $layer=licon1_PDIFF $count=1 $X=2.615
+ $Y=2.32 $X2=2.895 $Y2=2.815
r228 1 27 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=0.705
+ $Y=2.32 $X2=0.89 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_4%A_301_74# 1 2 3 4 13 19 22 23 24 26 27 30
+ 31 33 35 36 38 39 45
c128 31 0 1.68504e-19 $X=4.8 $Y=1.48
r129 45 48 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=5.28 $Y=2.625
+ $X2=5.28 $Y2=2.755
r130 36 44 22.3289 $w=2.23e-07 $l=4.30871e-07 $layer=LI1_cond $X=4.815 $Y=2.625
+ $X2=4.42 $Y2=2.55
r131 35 45 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.155 $Y=2.625
+ $X2=5.28 $Y2=2.625
r132 35 36 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.155 $Y=2.625
+ $X2=4.815 $Y2=2.625
r133 31 40 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.8 $Y=1.565
+ $X2=4.42 $Y2=1.565
r134 31 33 32.9599 $w=2.48e-07 $l=7.15e-07 $layer=LI1_cond $X=4.8 $Y=1.48
+ $X2=4.8 $Y2=0.765
r135 30 44 2.32876 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=4.42 $Y=2.39
+ $X2=4.42 $Y2=2.55
r136 29 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.42 $Y=1.65
+ $X2=4.42 $Y2=1.565
r137 29 30 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=4.42 $Y=1.65
+ $X2=4.42 $Y2=2.39
r138 28 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.105 $Y=2.475
+ $X2=3.02 $Y2=2.475
r139 27 44 5.36928 $w=2.23e-07 $l=1.16619e-07 $layer=LI1_cond $X=4.335 $Y=2.475
+ $X2=4.42 $Y2=2.55
r140 27 28 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=4.335 $Y=2.475
+ $X2=3.105 $Y2=2.475
r141 26 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.02 $Y=2.39
+ $X2=3.02 $Y2=2.475
r142 25 26 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=3.02 $Y=1.35
+ $X2=3.02 $Y2=2.39
r143 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.935 $Y=1.265
+ $X2=3.02 $Y2=1.35
r144 23 24 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.935 $Y=1.265
+ $X2=2.535 $Y2=1.265
r145 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.45 $Y=1.18
+ $X2=2.535 $Y2=1.265
r146 21 22 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.45 $Y=0.64
+ $X2=2.45 $Y2=1.18
r147 20 38 4.82444 $w=1.7e-07 $l=1.83916e-07 $layer=LI1_cond $X=1.925 $Y=2.475
+ $X2=1.76 $Y2=2.435
r148 19 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.935 $Y=2.475
+ $X2=3.02 $Y2=2.475
r149 19 20 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=2.935 $Y=2.475
+ $X2=1.925 $Y2=2.475
r150 13 21 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.365 $Y=0.515
+ $X2=2.45 $Y2=0.64
r151 13 15 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=2.365 $Y=0.515
+ $X2=1.805 $Y2=0.515
r152 4 48 600 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_PDIFF $count=1 $X=5.175
+ $Y=2.53 $X2=5.32 $Y2=2.755
r153 3 38 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=1.625
+ $Y=2.32 $X2=1.76 $Y2=2.475
r154 2 33 182 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_NDIFF $count=1 $X=4.695
+ $Y=0.5 $X2=4.84 $Y2=0.765
r155 1 15 182 $w=1.7e-07 $l=3.81445e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.37 $X2=1.805 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_4%Q 1 2 3 4 15 19 21 23 25 26 29 33 39 42 43
r73 40 43 3.31686 $w=5.93e-07 $l=1.65e-07 $layer=LI1_cond $X=12.057 $Y=1.13
+ $X2=12.057 $Y2=1.295
r74 40 42 3.49788 $w=3.92e-07 $l=1.44482e-07 $layer=LI1_cond $X=12.057 $Y=1.13
+ $X2=12.015 $Y2=1.005
r75 37 43 10.1516 $w=5.93e-07 $l=5.05e-07 $layer=LI1_cond $X=12.057 $Y=1.8
+ $X2=12.057 $Y2=1.295
r76 37 39 2.46131 $w=3.92e-07 $l=1.28367e-07 $layer=LI1_cond $X=12.057 $Y=1.8
+ $X2=12.01 $Y2=1.907
r77 31 42 3.49788 $w=3.92e-07 $l=3.01081e-07 $layer=LI1_cond $X=11.77 $Y=0.88
+ $X2=12.015 $Y2=1.005
r78 31 33 21.3062 $w=1.88e-07 $l=3.65e-07 $layer=LI1_cond $X=11.77 $Y=0.88
+ $X2=11.77 $Y2=0.515
r79 27 39 2.46131 $w=3.92e-07 $l=2.99165e-07 $layer=LI1_cond $X=11.76 $Y=2.015
+ $X2=12.01 $Y2=1.907
r80 27 29 46.6986 $w=1.88e-07 $l=8e-07 $layer=LI1_cond $X=11.76 $Y=2.015
+ $X2=11.76 $Y2=2.815
r81 25 39 4.47094 $w=1.7e-07 $l=3.5583e-07 $layer=LI1_cond $X=11.665 $Y=1.885
+ $X2=12.01 $Y2=1.907
r82 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=11.665 $Y=1.885
+ $X2=11.015 $Y2=1.885
r83 24 36 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=10.995 $Y=1.005
+ $X2=10.87 $Y2=1.005
r84 23 42 3.00706 $w=2.5e-07 $l=3.4e-07 $layer=LI1_cond $X=11.675 $Y=1.005
+ $X2=12.015 $Y2=1.005
r85 23 24 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=11.675 $Y=1.005
+ $X2=10.995 $Y2=1.005
r86 19 36 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=10.87 $Y=0.88
+ $X2=10.87 $Y2=1.005
r87 19 21 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=10.87 $Y=0.88
+ $X2=10.87 $Y2=0.515
r88 15 17 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=10.85 $Y=1.985
+ $X2=10.85 $Y2=2.815
r89 13 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.85 $Y=1.97
+ $X2=11.015 $Y2=1.885
r90 13 15 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=10.85 $Y=1.97
+ $X2=10.85 $Y2=1.985
r91 4 39 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=11.615
+ $Y=1.84 $X2=11.75 $Y2=1.985
r92 4 29 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=11.615
+ $Y=1.84 $X2=11.75 $Y2=2.815
r93 3 17 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.715
+ $Y=1.84 $X2=10.85 $Y2=2.815
r94 3 15 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.715
+ $Y=1.84 $X2=10.85 $Y2=1.985
r95 2 42 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=11.63
+ $Y=0.37 $X2=11.77 $Y2=0.965
r96 2 33 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=11.63
+ $Y=0.37 $X2=11.77 $Y2=0.515
r97 1 36 182 $w=1.7e-07 $l=6.98498e-07 $layer=licon1_NDIFF $count=1 $X=10.685
+ $Y=0.37 $X2=10.91 $Y2=0.965
r98 1 21 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=10.685
+ $Y=0.37 $X2=10.91 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXTP_4%VGND 1 2 3 4 5 6 7 8 29 33 37 41 45 49 53
+ 55 57 60 61 63 64 66 67 68 86 93 98 103 109 112 115 118 122
r145 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r146 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r147 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r148 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r149 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r150 107 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r151 107 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r152 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r153 104 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.505 $Y=0
+ $X2=11.34 $Y2=0
r154 104 106 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.505 $Y=0
+ $X2=11.76 $Y2=0
r155 103 121 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=12.035 $Y=0
+ $X2=12.257 $Y2=0
r156 103 106 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=12.035 $Y=0
+ $X2=11.76 $Y2=0
r157 102 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r158 102 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r159 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r160 99 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.515 $Y=0
+ $X2=10.35 $Y2=0
r161 99 101 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=10.515 $Y=0
+ $X2=10.8 $Y2=0
r162 98 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.175 $Y=0
+ $X2=11.34 $Y2=0
r163 98 101 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.175 $Y=0
+ $X2=10.8 $Y2=0
r164 97 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r165 97 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=9.36 $Y2=0
r166 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r167 94 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.525 $Y=0
+ $X2=9.36 $Y2=0
r168 94 96 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.525 $Y=0
+ $X2=9.84 $Y2=0
r169 93 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.185 $Y=0
+ $X2=10.35 $Y2=0
r170 93 96 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=10.185 $Y=0
+ $X2=9.84 $Y2=0
r171 92 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r172 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r173 89 92 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=8.88 $Y2=0
r174 88 91 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.96 $Y=0 $X2=8.88
+ $Y2=0
r175 88 89 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r176 86 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.195 $Y=0
+ $X2=9.36 $Y2=0
r177 86 91 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.195 $Y=0
+ $X2=8.88 $Y2=0
r178 85 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r179 84 85 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r180 81 84 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6.48
+ $Y2=0
r181 81 82 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r182 79 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r183 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r184 76 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r185 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r186 73 76 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r187 73 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r188 72 75 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r189 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r190 70 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=0
+ $X2=0.825 $Y2=0
r191 70 72 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.2
+ $Y2=0
r192 68 85 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.24 $Y=0
+ $X2=6.48 $Y2=0
r193 68 82 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=6.24 $Y=0
+ $X2=4.08 $Y2=0
r194 66 84 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=6.49 $Y=0 $X2=6.48
+ $Y2=0
r195 66 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.49 $Y=0 $X2=6.655
+ $Y2=0
r196 65 88 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.82 $Y=0 $X2=6.96
+ $Y2=0
r197 65 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.82 $Y=0 $X2=6.655
+ $Y2=0
r198 63 78 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.6
+ $Y2=0
r199 63 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.85
+ $Y2=0
r200 62 81 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.015 $Y=0 $X2=4.08
+ $Y2=0
r201 62 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.015 $Y=0 $X2=3.85
+ $Y2=0
r202 60 75 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.705 $Y=0 $X2=2.64
+ $Y2=0
r203 60 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.705 $Y=0 $X2=2.83
+ $Y2=0
r204 59 78 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=2.955 $Y=0 $X2=3.6
+ $Y2=0
r205 59 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.955 $Y=0 $X2=2.83
+ $Y2=0
r206 55 121 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=12.2 $Y=0.085
+ $X2=12.257 $Y2=0
r207 55 57 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=12.2 $Y=0.085
+ $X2=12.2 $Y2=0.57
r208 51 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.34 $Y=0.085
+ $X2=11.34 $Y2=0
r209 51 53 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=11.34 $Y=0.085
+ $X2=11.34 $Y2=0.53
r210 47 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.35 $Y=0.085
+ $X2=10.35 $Y2=0
r211 47 49 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=10.35 $Y=0.085
+ $X2=10.35 $Y2=0.495
r212 43 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.36 $Y=0.085
+ $X2=9.36 $Y2=0
r213 43 45 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=9.36 $Y=0.085
+ $X2=9.36 $Y2=0.54
r214 39 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.655 $Y=0.085
+ $X2=6.655 $Y2=0
r215 39 41 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.655 $Y=0.085
+ $X2=6.655 $Y2=0.515
r216 35 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=0.085
+ $X2=3.85 $Y2=0
r217 35 37 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.85 $Y=0.085
+ $X2=3.85 $Y2=0.55
r218 31 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.83 $Y=0.085
+ $X2=2.83 $Y2=0
r219 31 33 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=2.83 $Y=0.085
+ $X2=2.83 $Y2=0.58
r220 27 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0
r221 27 29 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0.565
r222 8 57 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=12.06
+ $Y=0.37 $X2=12.2 $Y2=0.57
r223 7 53 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=11.2
+ $Y=0.37 $X2=11.34 $Y2=0.53
r224 6 49 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=10.21
+ $Y=0.37 $X2=10.35 $Y2=0.495
r225 5 45 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=9.22
+ $Y=0.37 $X2=9.36 $Y2=0.54
r226 4 41 182 $w=1.7e-07 $l=2.27376e-07 $layer=licon1_NDIFF $count=1 $X=6.435
+ $Y=0.5 $X2=6.655 $Y2=0.515
r227 3 37 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=3.705
+ $Y=0.37 $X2=3.85 $Y2=0.55
r228 2 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.65
+ $Y=0.37 $X2=2.79 $Y2=0.58
r229 1 29 182 $w=1.7e-07 $l=2.91633e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.37 $X2=0.825 $Y2=0.565
.ends


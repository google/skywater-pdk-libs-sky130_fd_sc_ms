* NGSPICE file created from sky130_fd_sc_ms__a41oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__a41oi_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 VPWR A2 a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=1.1648e+12p pd=6.56e+06u as=9.744e+11p ps=8.46e+06u
M1001 Y A1 a_469_74# VNB nlowvt w=740000u l=150000u
+  ad=4.218e+11p pd=4.1e+06u as=3.108e+11p ps=2.32e+06u
M1002 VPWR A4 a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_119_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1004 a_119_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_277_74# A4 VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=4.921e+11p ps=2.81e+06u
M1006 a_355_74# A3 a_277_74# VNB nlowvt w=740000u l=150000u
+  ad=3.108e+11p pd=2.32e+06u as=0p ps=0u
M1007 VGND B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_469_74# A2 a_355_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_119_368# A3 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


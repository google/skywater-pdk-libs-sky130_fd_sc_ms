* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__ha_2 A B VGND VNB VPB VPWR COUT SUM
X0 a_278_74# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_394_388# a_27_74# a_278_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 VGND a_27_74# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VPWR B a_27_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X4 SUM a_394_388# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 COUT a_27_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_394_388# a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X7 VPWR A a_310_388# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X8 a_27_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X9 VPWR a_394_388# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X10 a_310_388# B a_394_388# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X11 SUM a_394_388# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VGND A a_278_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 VPWR a_27_74# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X14 VGND a_394_388# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 a_27_74# B a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 a_114_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 COUT a_27_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
.ends

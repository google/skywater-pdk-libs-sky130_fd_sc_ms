* File: sky130_fd_sc_ms__o21ai_4.spice
* Created: Fri Aug 28 17:55:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o21ai_4.pex.spice"
.subckt sky130_fd_sc_ms__o21ai_4  VNB VPB A1 B1 A2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2	A2
* B1	B1
* A1	A1
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A1_M1009_g N_A_27_74#_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75005 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1009_d N_A1_M1018_g N_A_27_74#_M1018_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75004.5 A=0.111 P=1.78 MULT=1
MM1019 N_VGND_M1019_d N_A1_M1019_g N_A_27_74#_M1018_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10915 AS=0.1036 PD=1.035 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75004.1 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1019_d N_A1_M1021_g N_A_27_74#_M1021_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10915 AS=0.1036 PD=1.035 PS=1.02 NRD=2.424 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75003.7 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_B1_M1002_g N_A_27_74#_M1021_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1002_d N_B1_M1003_g N_A_27_74#_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.4
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1010 N_Y_M1010_d N_B1_M1010_g N_A_27_74#_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1017 N_Y_M1010_d N_B1_M1017_g N_A_27_74#_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.11285 PD=1.02 PS=1.045 NRD=0 NRS=4.044 M=1 R=4.93333 SA=75003.2
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_27_74#_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.11285 PD=1.02 PS=1.045 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.7
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1000_d N_A2_M1001_g N_A_27_74#_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.1
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_A2_M1008_g N_A_27_74#_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.5
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1008_d N_A2_M1016_g N_A_27_74#_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75005
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_A_119_368#_M1004_d N_A1_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90002.5 A=0.2016 P=2.6 MULT=1
MM1005 N_A_119_368#_M1004_d N_A1_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90002.1 A=0.2016 P=2.6 MULT=1
MM1006 N_A_119_368#_M1006_d N_A1_M1006_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1007 N_A_119_368#_M1006_d N_A1_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1011 N_Y_M1011_d N_B1_M1011_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1012 N_Y_M1011_d N_B1_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.4088 PD=1.39 PS=2.97 NRD=0 NRS=14.0658 M=1 R=6.22222 SA=90002.4
+ SB=90000.3 A=0.2016 P=2.6 MULT=1
MM1013 N_A_119_368#_M1013_d N_A2_M1013_g N_Y_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1792 PD=2.8 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.2
+ SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1014 N_A_119_368#_M1014_d N_A2_M1014_g N_Y_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.7
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1015 N_A_119_368#_M1014_d N_A2_M1015_g N_Y_M1015_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1020 N_A_119_368#_M1020_d N_A2_M1020_g N_Y_M1015_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX22_noxref VNB VPB NWDIODE A=11.4204 P=16
c_57 VNB 0 1.07857e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__o21ai_4.pxi.spice"
*
.ends
*
*

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__sdfbbn_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__sdfbbn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  16.80000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.480000 1.815000 1.810000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.524500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.335000 0.350000 16.715000 1.050000 ;
        RECT 16.355000 1.820000 16.715000 2.980000 ;
        RECT 16.545000 1.050000 16.715000 1.820000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.524500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.890000 1.820000 15.275000 2.980000 ;
        RECT 14.915000 0.350000 15.275000 1.130000 ;
        RECT 15.105000 1.130000 15.275000 1.820000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.075000 1.190000 14.380000 1.550000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.205000 0.550000 1.875000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.805000 1.205000 1.315000 1.875000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.524700 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  8.285000 1.790000  8.990000 1.960000 ;
        RECT  8.285000 1.960000  8.490000 2.140000 ;
        RECT  8.660000 1.630000  8.990000 1.790000 ;
        RECT 11.630000 1.470000 11.960000 2.120000 ;
      LAYER mcon ;
        RECT  8.315000 1.950000  8.485000 2.120000 ;
        RECT 11.675000 1.950000 11.845000 2.120000 ;
      LAYER met1 ;
        RECT  8.255000 1.920000  8.545000 1.965000 ;
        RECT  8.255000 1.965000 11.905000 2.105000 ;
        RECT  8.255000 2.105000  8.545000 2.150000 ;
        RECT 11.615000 1.920000 11.905000 1.965000 ;
        RECT 11.615000 2.105000 11.905000 2.150000 ;
    END
  END SET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.470000 1.350000 3.800000 1.780000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 16.800000 0.085000 ;
        RECT  0.140000  0.085000  0.470000 1.035000 ;
        RECT  1.890000  0.085000  2.220000 0.970000 ;
        RECT  3.800000  0.085000  4.130000 0.410000 ;
        RECT  5.300000  0.085000  5.630000 1.035000 ;
        RECT  8.795000  0.085000  9.125000 1.080000 ;
        RECT 11.415000  0.085000 11.755000 0.410000 ;
        RECT 14.415000  0.085000 14.735000 0.680000 ;
        RECT 15.905000  0.085000 16.155000 1.050000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
        RECT 15.035000 -0.085000 15.205000 0.085000 ;
        RECT 15.515000 -0.085000 15.685000 0.085000 ;
        RECT 15.995000 -0.085000 16.165000 0.085000 ;
        RECT 16.475000 -0.085000 16.645000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 16.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 16.800000 3.415000 ;
        RECT  0.565000 2.385000  0.895000 3.245000 ;
        RECT  2.470000 2.300000  2.720000 3.245000 ;
        RECT  3.930000 2.290000  4.180000 3.245000 ;
        RECT  5.020000 2.465000  5.270000 3.245000 ;
        RECT  8.125000 2.650000  8.295000 3.245000 ;
        RECT  9.050000 2.470000  9.380000 3.245000 ;
        RECT 10.900000 2.970000 11.230000 3.245000 ;
        RECT 11.995000 2.970000 12.325000 3.245000 ;
        RECT 14.000000 2.550000 14.690000 3.245000 ;
        RECT 15.905000 1.900000 16.155000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
        RECT 14.555000 3.245000 14.725000 3.415000 ;
        RECT 15.035000 3.245000 15.205000 3.415000 ;
        RECT 15.515000 3.245000 15.685000 3.415000 ;
        RECT 15.995000 3.245000 16.165000 3.415000 ;
        RECT 16.475000 3.245000 16.645000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 16.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.115000 2.045000  1.235000 2.215000 ;
      RECT  0.115000 2.215000  0.395000 2.980000 ;
      RECT  0.960000 0.575000  1.290000 0.865000 ;
      RECT  0.960000 0.865000  1.655000 1.035000 ;
      RECT  1.065000 2.215000  1.235000 2.905000 ;
      RECT  1.065000 2.905000  2.245000 3.075000 ;
      RECT  1.465000 2.300000  1.715000 2.735000 ;
      RECT  1.485000 1.035000  1.655000 1.140000 ;
      RECT  1.485000 1.140000  2.560000 1.310000 ;
      RECT  1.545000 1.980000  2.155000 2.150000 ;
      RECT  1.545000 2.150000  1.715000 2.300000 ;
      RECT  1.915000 2.320000  2.245000 2.905000 ;
      RECT  1.985000 1.310000  2.155000 1.980000 ;
      RECT  2.390000 0.255000  3.400000 0.425000 ;
      RECT  2.390000 0.425000  2.560000 1.140000 ;
      RECT  2.510000 1.480000  3.060000 1.810000 ;
      RECT  2.730000 0.595000  3.060000 1.480000 ;
      RECT  2.890000 1.810000  3.060000 2.300000 ;
      RECT  2.890000 2.300000  3.250000 2.980000 ;
      RECT  3.230000 0.425000  3.400000 0.580000 ;
      RECT  3.230000 0.580000  5.130000 0.750000 ;
      RECT  3.290000 0.920000  4.140000 1.170000 ;
      RECT  3.480000 1.950000  4.140000 2.120000 ;
      RECT  3.480000 2.120000  3.730000 2.980000 ;
      RECT  3.970000 1.170000  4.140000 1.340000 ;
      RECT  3.970000 1.340000  4.440000 1.670000 ;
      RECT  3.970000 1.670000  4.140000 1.950000 ;
      RECT  4.310000 0.920000  4.790000 1.170000 ;
      RECT  4.380000 1.840000  4.780000 2.980000 ;
      RECT  4.610000 1.170000  4.790000 1.550000 ;
      RECT  4.610000 1.550000  6.710000 1.720000 ;
      RECT  4.610000 1.720000  4.780000 1.840000 ;
      RECT  4.950000 1.965000  5.215000 2.125000 ;
      RECT  4.950000 2.125000  5.610000 2.295000 ;
      RECT  4.960000 0.750000  5.130000 1.205000 ;
      RECT  4.960000 1.205000  5.970000 1.375000 ;
      RECT  5.405000 1.720000  6.710000 1.800000 ;
      RECT  5.405000 1.800000  5.755000 1.905000 ;
      RECT  5.440000 2.295000  5.610000 2.905000 ;
      RECT  5.440000 2.905000  7.505000 3.075000 ;
      RECT  5.800000 0.255000  6.925000 0.425000 ;
      RECT  5.800000 0.425000  5.970000 1.205000 ;
      RECT  5.865000 2.245000  6.195000 2.735000 ;
      RECT  6.025000 1.970000  7.250000 2.140000 ;
      RECT  6.025000 2.140000  6.195000 2.245000 ;
      RECT  6.170000 0.595000  6.420000 1.130000 ;
      RECT  6.170000 1.130000  7.250000 1.300000 ;
      RECT  6.365000 2.310000  7.590000 2.480000 ;
      RECT  6.365000 2.480000  6.695000 2.735000 ;
      RECT  6.380000 1.470000  6.710000 1.550000 ;
      RECT  6.595000 0.425000  6.925000 0.790000 ;
      RECT  6.595000 0.790000  7.590000 0.960000 ;
      RECT  6.920000 1.300000  7.250000 1.970000 ;
      RECT  6.925000 2.650000  7.930000 2.820000 ;
      RECT  6.925000 2.820000  7.505000 2.905000 ;
      RECT  7.150000 0.255000  8.590000 0.425000 ;
      RECT  7.150000 0.425000  7.480000 0.620000 ;
      RECT  7.420000 0.960000  7.590000 2.310000 ;
      RECT  7.760000 0.595000  8.090000 1.080000 ;
      RECT  7.760000 1.080000  7.930000 2.310000 ;
      RECT  7.760000 2.310000  8.830000 2.480000 ;
      RECT  7.760000 2.480000  7.930000 2.650000 ;
      RECT  8.100000 1.290000  9.555000 1.460000 ;
      RECT  8.100000 1.460000  8.430000 1.620000 ;
      RECT  8.260000 0.425000  8.590000 1.080000 ;
      RECT  8.495000 2.480000  8.830000 2.980000 ;
      RECT  8.660000 2.130000  9.530000 2.300000 ;
      RECT  8.660000 2.300000  8.830000 2.310000 ;
      RECT  9.200000 1.630000  9.530000 2.130000 ;
      RECT  9.385000 0.365000 10.920000 0.535000 ;
      RECT  9.385000 0.535000  9.555000 1.290000 ;
      RECT  9.725000 1.260000 11.000000 1.555000 ;
      RECT  9.725000 1.555000 10.070000 1.940000 ;
      RECT  9.745000 0.705000 10.580000 0.920000 ;
      RECT  9.745000 0.920000 11.340000 1.090000 ;
      RECT  9.890000 2.110000 10.410000 2.280000 ;
      RECT  9.890000 2.280000 10.220000 2.980000 ;
      RECT 10.240000 1.725000 11.340000 1.895000 ;
      RECT 10.240000 1.895000 10.410000 2.110000 ;
      RECT 10.665000 2.065000 10.995000 2.630000 ;
      RECT 10.665000 2.630000 13.280000 2.800000 ;
      RECT 10.750000 0.535000 10.920000 0.580000 ;
      RECT 10.750000 0.580000 11.680000 0.750000 ;
      RECT 11.170000 1.090000 11.340000 1.725000 ;
      RECT 11.170000 1.895000 11.340000 2.290000 ;
      RECT 11.170000 2.290000 12.780000 2.460000 ;
      RECT 11.460000 2.800000 11.790000 2.980000 ;
      RECT 11.510000 0.750000 11.680000 1.130000 ;
      RECT 11.510000 1.130000 13.905000 1.300000 ;
      RECT 11.935000 0.255000 13.225000 0.425000 ;
      RECT 11.935000 0.425000 12.265000 0.960000 ;
      RECT 12.200000 1.300000 12.530000 1.550000 ;
      RECT 12.465000 0.595000 12.795000 0.790000 ;
      RECT 12.465000 0.790000 13.565000 0.960000 ;
      RECT 12.610000 1.720000 13.440000 1.890000 ;
      RECT 12.610000 1.890000 12.780000 2.290000 ;
      RECT 12.770000 1.470000 13.440000 1.720000 ;
      RECT 12.950000 2.060000 13.280000 2.210000 ;
      RECT 12.950000 2.210000 14.720000 2.380000 ;
      RECT 12.950000 2.380000 13.280000 2.630000 ;
      RECT 12.950000 2.800000 13.280000 2.980000 ;
      RECT 12.975000 0.425000 13.225000 0.620000 ;
      RECT 13.395000 0.330000 14.245000 0.500000 ;
      RECT 13.395000 0.500000 13.565000 0.790000 ;
      RECT 13.610000 1.300000 13.780000 1.790000 ;
      RECT 13.610000 1.790000 14.130000 2.040000 ;
      RECT 13.735000 0.670000 13.905000 1.130000 ;
      RECT 14.075000 0.500000 14.245000 0.850000 ;
      RECT 14.075000 0.850000 14.720000 1.020000 ;
      RECT 14.550000 1.020000 14.720000 1.300000 ;
      RECT 14.550000 1.300000 14.935000 1.630000 ;
      RECT 14.550000 1.630000 14.720000 2.210000 ;
      RECT 15.450000 0.350000 15.725000 1.220000 ;
      RECT 15.450000 1.220000 16.375000 1.550000 ;
      RECT 15.450000 1.550000 15.700000 2.780000 ;
    LAYER mcon ;
      RECT 5.435000 1.580000 5.605000 1.750000 ;
      RECT 9.755000 1.580000 9.925000 1.750000 ;
    LAYER met1 ;
      RECT 5.375000 1.550000 5.665000 1.595000 ;
      RECT 5.375000 1.595000 9.985000 1.735000 ;
      RECT 5.375000 1.735000 5.665000 1.780000 ;
      RECT 9.695000 1.550000 9.985000 1.595000 ;
      RECT 9.695000 1.735000 9.985000 1.780000 ;
  END
END sky130_fd_sc_ms__sdfbbn_1

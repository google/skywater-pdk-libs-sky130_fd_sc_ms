* NGSPICE file created from sky130_fd_sc_ms__xnor3_4.ext - technology: sky130A

.subckt sky130_fd_sc_ms__xnor3_4 A B C VGND VNB VPB VPWR X
M1000 a_75_227# a_386_23# a_321_77# VPB pshort w=840000u l=180000u
+  ad=7.2195e+11p pd=5.6e+06u as=4.964e+11p ps=4.58e+06u
M1001 X a_1057_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=2.35215e+12p ps=1.359e+07u
M1002 X a_1057_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=2.2864e+12p ps=1.53e+07u
M1003 a_75_227# A VGND VNB nlowvt w=640000u l=150000u
+  ad=5.611e+11p pd=4.74e+06u as=0p ps=0u
M1004 X a_1057_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_327_373# B a_27_373# VNB nlowvt w=640000u l=150000u
+  ad=3.84e+11p pd=3.76e+06u as=4.635e+11p ps=4.06e+06u
M1006 a_27_373# a_386_23# a_321_77# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=3.739e+11p ps=3.78e+06u
M1007 VPWR B a_386_23# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1008 VPWR a_1057_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_75_227# a_386_23# a_327_373# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_327_373# C a_1057_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.592e+11p ps=2.09e+06u
M1011 VGND a_1057_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR C a_1024_300# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1013 VGND a_1057_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_373# a_386_23# a_327_373# VPB pshort w=640000u l=180000u
+  ad=4.528e+11p pd=4.38e+06u as=6.18e+11p ps=4.96e+06u
M1015 a_321_77# B a_27_373# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_75_227# a_27_373# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND C a_1024_300# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1018 a_75_227# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_321_77# C a_1057_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=4.305e+11p ps=2.98e+06u
M1020 VPWR a_75_227# a_27_373# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1057_74# a_1024_300# a_327_373# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND B a_386_23# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1023 X a_1057_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_321_77# B a_75_227# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_327_373# B a_75_227# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_1057_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1057_74# a_1024_300# a_321_77# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__xnor3_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__xnor3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.845000 1.425000 7.205000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.771000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.705000 1.350000 4.375000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.425400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 1.350000 1.325000 1.780000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.513300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.440000 0.445000 1.170000 ;
        RECT 0.085000 1.170000 0.255000 1.840000 ;
        RECT 0.085000 1.840000 0.355000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.160000 0.085000 ;
        RECT 0.625000  0.085000 0.955000 0.490000 ;
        RECT 3.395000  0.085000 3.725000 0.500000 ;
        RECT 7.205000  0.085000 7.615000 0.915000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 8.160000 3.415000 ;
        RECT 0.555000 2.290000 0.805000 3.245000 ;
        RECT 3.395000 2.710000 3.725000 3.245000 ;
        RECT 7.260000 2.290000 7.590000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.425000 1.340000 0.785000 1.670000 ;
      RECT 0.615000 0.660000 1.665000 0.830000 ;
      RECT 0.615000 0.830000 0.785000 1.340000 ;
      RECT 0.615000 1.670000 0.785000 1.950000 ;
      RECT 0.615000 1.950000 1.145000 2.120000 ;
      RECT 0.975000 2.120000 1.145000 2.905000 ;
      RECT 0.975000 2.905000 2.655000 3.075000 ;
      RECT 1.135000 1.000000 1.665000 1.170000 ;
      RECT 1.315000 1.950000 1.665000 2.500000 ;
      RECT 1.495000 0.255000 2.665000 0.425000 ;
      RECT 1.495000 0.425000 1.665000 0.660000 ;
      RECT 1.495000 1.170000 1.665000 1.580000 ;
      RECT 1.495000 1.580000 2.845000 1.750000 ;
      RECT 1.495000 1.750000 1.665000 1.950000 ;
      RECT 1.835000 0.595000 2.165000 1.140000 ;
      RECT 1.835000 1.140000 3.185000 1.310000 ;
      RECT 1.835000 1.310000 2.275000 1.410000 ;
      RECT 1.875000 1.950000 2.125000 2.370000 ;
      RECT 1.875000 2.370000 5.265000 2.540000 ;
      RECT 1.875000 2.540000 2.125000 2.735000 ;
      RECT 2.325000 2.710000 2.655000 2.905000 ;
      RECT 2.335000 0.425000 2.665000 0.970000 ;
      RECT 2.515000 1.480000 2.845000 1.580000 ;
      RECT 2.515000 1.750000 2.845000 1.810000 ;
      RECT 2.835000 0.350000 3.165000 0.670000 ;
      RECT 2.835000 0.670000 6.535000 0.765000 ;
      RECT 2.835000 0.765000 5.180000 0.840000 ;
      RECT 2.835000 0.840000 3.525000 0.970000 ;
      RECT 2.850000 2.030000 3.185000 2.200000 ;
      RECT 3.015000 1.310000 3.185000 2.030000 ;
      RECT 3.355000 0.970000 3.525000 2.370000 ;
      RECT 3.905000 1.010000 4.715000 1.180000 ;
      RECT 3.920000 1.950000 4.715000 2.200000 ;
      RECT 4.465000 0.255000 7.035000 0.425000 ;
      RECT 4.465000 0.425000 4.840000 0.500000 ;
      RECT 4.490000 2.710000 4.820000 2.905000 ;
      RECT 4.490000 2.905000 7.090000 3.075000 ;
      RECT 4.545000 1.180000 4.715000 1.355000 ;
      RECT 4.545000 1.355000 5.045000 1.685000 ;
      RECT 4.545000 1.685000 4.715000 1.950000 ;
      RECT 5.010000 0.595000 6.535000 0.670000 ;
      RECT 5.015000 1.855000 5.265000 2.370000 ;
      RECT 5.015000 2.540000 5.265000 2.575000 ;
      RECT 5.020000 1.015000 5.485000 1.180000 ;
      RECT 5.020000 1.180000 5.605000 1.185000 ;
      RECT 5.315000 1.185000 5.605000 1.410000 ;
      RECT 5.435000 1.410000 5.605000 1.765000 ;
      RECT 5.435000 1.765000 6.250000 1.935000 ;
      RECT 5.550000 2.105000 5.880000 2.565000 ;
      RECT 5.550000 2.565000 6.590000 2.735000 ;
      RECT 5.775000 0.935000 6.085000 1.425000 ;
      RECT 5.775000 1.425000 6.590000 1.595000 ;
      RECT 6.080000 1.935000 6.250000 2.395000 ;
      RECT 6.255000 0.765000 6.535000 1.210000 ;
      RECT 6.420000 1.595000 6.590000 2.565000 ;
      RECT 6.705000 0.425000 7.035000 1.085000 ;
      RECT 6.705000 1.085000 7.620000 1.255000 ;
      RECT 6.760000 1.950000 7.620000 2.120000 ;
      RECT 6.760000 2.120000 7.090000 2.905000 ;
      RECT 7.415000 1.255000 7.620000 1.425000 ;
      RECT 7.415000 1.425000 7.665000 1.755000 ;
      RECT 7.415000 1.755000 7.620000 1.950000 ;
      RECT 7.790000 2.190000 8.075000 2.930000 ;
      RECT 7.795000 0.585000 8.075000 1.255000 ;
      RECT 7.835000 1.255000 8.075000 2.190000 ;
    LAYER mcon ;
      RECT 2.075000 1.210000 2.245000 1.380000 ;
      RECT 5.435000 1.210000 5.605000 1.380000 ;
      RECT 5.915000 1.210000 6.085000 1.380000 ;
      RECT 7.835000 1.210000 8.005000 1.380000 ;
    LAYER met1 ;
      RECT 2.015000 1.180000 2.305000 1.225000 ;
      RECT 2.015000 1.225000 5.665000 1.365000 ;
      RECT 2.015000 1.365000 2.305000 1.410000 ;
      RECT 5.375000 1.180000 5.665000 1.225000 ;
      RECT 5.375000 1.365000 5.665000 1.410000 ;
      RECT 5.855000 1.180000 6.145000 1.225000 ;
      RECT 5.855000 1.225000 8.065000 1.365000 ;
      RECT 5.855000 1.365000 6.145000 1.410000 ;
      RECT 7.775000 1.180000 8.065000 1.225000 ;
      RECT 7.775000 1.365000 8.065000 1.410000 ;
  END
END sky130_fd_sc_ms__xnor3_1

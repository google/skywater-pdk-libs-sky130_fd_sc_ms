# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__o2111ai_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__o2111ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.350000 5.635000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.350000 4.675000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.350000 3.715000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.345000 1.300000 2.015000 1.630000 ;
        RECT 1.565000 1.180000 1.795000 1.300000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.550000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  1.416800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.180000 0.935000 1.800000 ;
        RECT 0.605000 1.800000 1.885000 1.950000 ;
        RECT 0.605000 1.950000 4.245000 1.970000 ;
        RECT 0.605000 1.970000 0.935000 2.980000 ;
        RECT 0.690000 0.595000 0.940000 1.130000 ;
        RECT 0.690000 1.130000 0.935000 1.180000 ;
        RECT 1.555000 1.970000 4.245000 2.120000 ;
        RECT 1.555000 2.120000 1.885000 2.980000 ;
        RECT 2.455000 2.120000 2.785000 2.980000 ;
        RECT 3.915000 2.120000 4.245000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.155000  1.820000 0.405000 3.245000 ;
      RECT 0.180000  0.255000 1.290000 0.425000 ;
      RECT 0.180000  0.425000 0.510000 1.010000 ;
      RECT 1.105000  2.140000 1.355000 3.245000 ;
      RECT 1.120000  0.425000 1.290000 0.840000 ;
      RECT 1.120000  0.840000 2.300000 1.010000 ;
      RECT 1.120000  1.010000 1.290000 1.130000 ;
      RECT 1.470000  0.255000 3.360000 0.425000 ;
      RECT 1.470000  0.425000 1.800000 0.670000 ;
      RECT 1.970000  0.595000 2.300000 0.840000 ;
      RECT 1.970000  1.010000 2.300000 1.130000 ;
      RECT 2.085000  2.290000 2.255000 3.245000 ;
      RECT 2.530000  0.595000 2.860000 1.010000 ;
      RECT 2.530000  1.010000 5.600000 1.180000 ;
      RECT 2.985000  2.290000 3.235000 3.245000 ;
      RECT 3.030000  0.425000 3.360000 0.840000 ;
      RECT 3.465000  2.290000 3.715000 2.905000 ;
      RECT 3.465000  2.905000 4.615000 3.075000 ;
      RECT 3.540000  0.350000 3.710000 1.010000 ;
      RECT 3.890000  0.085000 4.220000 0.840000 ;
      RECT 4.420000  0.350000 4.670000 1.010000 ;
      RECT 4.445000  1.950000 5.645000 2.120000 ;
      RECT 4.445000  2.120000 4.615000 2.905000 ;
      RECT 4.815000  2.290000 5.145000 3.245000 ;
      RECT 4.840000  0.085000 5.170000 0.840000 ;
      RECT 5.315000  2.120000 5.645000 2.980000 ;
      RECT 5.350000  0.350000 5.600000 1.010000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_ms__o2111ai_2

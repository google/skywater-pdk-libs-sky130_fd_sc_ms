* File: sky130_fd_sc_ms__a211oi_1.spice
* Created: Fri Aug 28 16:57:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a211oi_1.pex.spice"
.subckt sky130_fd_sc_ms__a211oi_1  VNB VPB A2 A1 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1003 A_159_74# N_A2_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74 AD=0.0777
+ AS=0.1961 PD=0.95 PS=2.01 NRD=8.1 NRS=0 M=1 R=4.93333 SA=75000.2 SB=75001.6
+ A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_A1_M1001_g A_159_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1443
+ AS=0.0777 PD=1.13 PS=0.95 NRD=3.24 NRS=8.1 M=1 R=4.93333 SA=75000.6 SB=75001.3
+ A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_B1_M1004_g N_Y_M1001_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.1443 PD=1.13 PS=1.13 NRD=3.24 NRS=14.592 M=1 R=4.93333
+ SA=75001.1 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1007 N_Y_M1007_d N_C1_M1007_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1443 PD=2.01 PS=1.13 NRD=0 NRS=14.592 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_A2_M1005_g N_A_71_368#_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2016 AS=0.2912 PD=1.48 PS=2.76 NRD=2.6201 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1000 N_A_71_368#_M1000_d N_A1_M1000_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2016 PD=1.39 PS=1.48 NRD=0 NRS=11.426 M=1 R=6.22222 SA=90000.7
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1002 A_357_368# N_B1_M1002_g N_A_71_368#_M1000_d VPB PSHORT L=0.18 W=1.12
+ AD=0.168 AS=0.1512 PD=1.42 PS=1.39 NRD=16.7056 NRS=0 M=1 R=6.22222 SA=90001.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1006 N_Y_M1006_d N_C1_M1006_g A_357_368# VPB PSHORT L=0.18 W=1.12 AD=0.2912
+ AS=0.168 PD=2.76 PS=1.42 NRD=0 NRS=16.7056 M=1 R=6.22222 SA=90001.6 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ms__a211oi_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__a21o_4.spice
* Created: Wed Sep  2 11:51:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a21o_4.pex.spice"
.subckt sky130_fd_sc_ms__a21o_4  VNB VPB B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1001 N_X_M1001_d N_A_91_48#_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1004 N_X_M1001_d N_A_91_48#_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1010 N_X_M1010_d N_A_91_48#_M1010_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75001.4 A=0.111 P=1.78 MULT=1
MM1012 N_X_M1010_d N_A_91_48#_M1012_g N_VGND_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.130894 PD=1.02 PS=1.15826 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001 A=0.111 P=1.78 MULT=1
MM1005 N_A_91_48#_M1005_d N_B1_M1005_g N_VGND_M1012_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.113206 PD=0.92 PS=1.00174 NRD=0 NRS=11.244 M=1 R=4.26667
+ SA=75002 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1019 N_A_91_48#_M1005_d N_B1_M1019_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.4
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1003 N_A_700_74#_M1003_d N_A1_M1003_g N_A_91_48#_M1003_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1017 N_A_700_74#_M1017_d N_A1_M1017_g N_A_91_48#_M1003_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1000 N_A_700_74#_M1017_d N_A2_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1015 N_A_700_74#_M1015_d N_A2_M1015_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_X_M1007_d N_A_91_48#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1008 N_X_M1007_d N_A_91_48#_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1011 N_X_M1011_d N_A_91_48#_M1011_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1014 N_X_M1011_d N_A_91_48#_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1006 N_A_91_48#_M1006_d N_B1_M1006_g N_A_503_392#_M1006_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90002.4 A=0.18 P=2.36 MULT=1
MM1009 N_A_91_48#_M1006_d N_B1_M1009_g N_A_503_392#_M1009_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.6
+ SB=90002 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1013_d N_A1_M1013_g N_A_503_392#_M1009_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.1
+ SB=90001.5 A=0.18 P=2.36 MULT=1
MM1016 N_VPWR_M1013_d N_A1_M1016_g N_A_503_392#_M1016_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.5
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1002 N_A_503_392#_M1016_s N_A2_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90002
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1018 N_A_503_392#_M1018_d N_A2_M1018_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1
+ AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90002.4
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ms__a21o_4.pxi.spice"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlrtn_4 D GATE_N RESET_B VGND VNB VPB VPWR Q
M1000 a_750_504# a_232_98# a_642_392# VPB pshort w=420000u l=180000u
+  ad=2.898e+11p pd=2.22e+06u as=3.158e+11p ps=2.72e+06u
M1001 VGND a_888_406# Q VNB nlowvt w=740000u l=150000u
+  ad=2.1144e+12p pd=1.632e+07u as=4.144e+11p ps=4.08e+06u
M1002 a_1035_74# RESET_B VGND VNB nlowvt w=640000u l=150000u
+  ad=5.44e+11p pd=5.54e+06u as=0p ps=0u
M1003 a_232_98# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=0p ps=0u
M1004 VGND a_888_406# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_564_392# a_27_136# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.1e+11p pd=2.42e+06u as=2.5597e+12p ps=1.989e+07u
M1006 a_839_74# a_348_392# a_642_392# VNB nlowvt w=420000u l=150000u
+  ad=1.155e+11p pd=1.39e+06u as=1.915e+11p ps=1.93e+06u
M1007 a_232_98# GATE_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1008 VPWR a_232_98# a_348_392# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1009 a_1035_74# a_642_392# a_888_406# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1010 VPWR a_888_406# a_750_504# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Q a_888_406# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_888_406# a_642_392# VPWR VPB pshort w=840000u l=180000u
+  ad=5.124e+11p pd=4.58e+06u as=0p ps=0u
M1013 VPWR D a_27_136# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1014 a_888_406# RESET_B VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_888_406# a_839_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_642_392# a_888_406# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_642_392# a_232_98# a_666_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1018 a_666_74# a_27_136# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_888_406# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=7.168e+11p ps=5.76e+06u
M1020 VGND a_232_98# a_348_392# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1021 VGND RESET_B a_1035_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Q a_888_406# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q a_888_406# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND D a_27_136# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1025 Q a_888_406# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_888_406# a_642_392# a_1035_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR a_888_406# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_642_392# a_348_392# a_564_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR RESET_B a_888_406# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

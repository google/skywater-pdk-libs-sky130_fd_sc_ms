* File: sky130_fd_sc_ms__mux2_4.pxi.spice
* Created: Fri Aug 28 17:39:53 2020
* 
x_PM_SKY130_FD_SC_MS__MUX2_4%S N_S_M1009_g N_S_M1002_g N_S_M1001_g N_S_M1010_g
+ N_S_M1024_g N_S_M1013_g N_S_c_166_n N_S_c_176_p N_S_c_177_p N_S_c_182_p
+ N_S_c_167_n N_S_c_158_n N_S_c_159_n N_S_c_183_p S N_S_c_160_n N_S_c_161_n
+ N_S_c_162_n PM_SKY130_FD_SC_MS__MUX2_4%S
x_PM_SKY130_FD_SC_MS__MUX2_4%A_27_368# N_A_27_368#_M1002_s N_A_27_368#_M1009_s
+ N_A_27_368#_M1015_g N_A_27_368#_M1003_g N_A_27_368#_M1007_g
+ N_A_27_368#_M1018_g N_A_27_368#_c_300_n N_A_27_368#_c_312_n
+ N_A_27_368#_c_301_n N_A_27_368#_c_317_n N_A_27_368#_c_321_n
+ N_A_27_368#_c_302_n N_A_27_368#_c_303_n N_A_27_368#_c_304_n
+ N_A_27_368#_c_293_n N_A_27_368#_c_294_n N_A_27_368#_c_295_n
+ N_A_27_368#_c_306_n N_A_27_368#_c_296_n N_A_27_368#_c_348_n
+ N_A_27_368#_c_297_n PM_SKY130_FD_SC_MS__MUX2_4%A_27_368#
x_PM_SKY130_FD_SC_MS__MUX2_4%A_193_241# N_A_193_241#_M1017_s
+ N_A_193_241#_M1022_s N_A_193_241#_M1025_d N_A_193_241#_M1011_s
+ N_A_193_241#_M1016_s N_A_193_241#_M1008_s N_A_193_241#_M1000_g
+ N_A_193_241#_M1006_g N_A_193_241#_c_429_n N_A_193_241#_c_430_n
+ N_A_193_241#_c_431_n N_A_193_241#_M1004_g N_A_193_241#_M1012_g
+ N_A_193_241#_c_434_n N_A_193_241#_M1021_g N_A_193_241#_c_436_n
+ N_A_193_241#_M1019_g N_A_193_241#_c_438_n N_A_193_241#_M1023_g
+ N_A_193_241#_c_440_n N_A_193_241#_c_441_n N_A_193_241#_M1020_g
+ N_A_193_241#_c_443_n N_A_193_241#_c_444_n N_A_193_241#_c_445_n
+ N_A_193_241#_c_446_n N_A_193_241#_c_447_n N_A_193_241#_c_448_n
+ N_A_193_241#_c_449_n N_A_193_241#_c_465_n N_A_193_241#_c_466_n
+ N_A_193_241#_c_467_n N_A_193_241#_c_450_n N_A_193_241#_c_526_p
+ N_A_193_241#_c_451_n N_A_193_241#_c_452_n N_A_193_241#_c_468_n
+ N_A_193_241#_c_453_n N_A_193_241#_c_454_n N_A_193_241#_c_455_n
+ N_A_193_241#_c_456_n N_A_193_241#_c_457_n N_A_193_241#_c_470_n
+ N_A_193_241#_c_458_n PM_SKY130_FD_SC_MS__MUX2_4%A_193_241#
x_PM_SKY130_FD_SC_MS__MUX2_4%A0 N_A0_M1017_g N_A0_M1011_g N_A0_M1022_g
+ N_A0_M1016_g A0 N_A0_c_648_n PM_SKY130_FD_SC_MS__MUX2_4%A0
x_PM_SKY130_FD_SC_MS__MUX2_4%A1 N_A1_M1005_g N_A1_M1014_g N_A1_M1008_g
+ N_A1_M1025_g A1 A1 N_A1_c_692_n N_A1_c_693_n PM_SKY130_FD_SC_MS__MUX2_4%A1
x_PM_SKY130_FD_SC_MS__MUX2_4%VPWR N_VPWR_M1009_d N_VPWR_M1004_s N_VPWR_M1020_s
+ N_VPWR_M1013_s N_VPWR_M1018_s N_VPWR_c_737_n N_VPWR_c_738_n N_VPWR_c_739_n
+ N_VPWR_c_740_n N_VPWR_c_741_n N_VPWR_c_742_n N_VPWR_c_743_n N_VPWR_c_744_n
+ N_VPWR_c_745_n N_VPWR_c_746_n N_VPWR_c_747_n VPWR N_VPWR_c_748_n
+ N_VPWR_c_749_n N_VPWR_c_736_n N_VPWR_c_751_n N_VPWR_c_752_n
+ PM_SKY130_FD_SC_MS__MUX2_4%VPWR
x_PM_SKY130_FD_SC_MS__MUX2_4%X N_X_M1006_d N_X_M1021_d N_X_M1000_d N_X_M1019_d
+ N_X_c_837_n N_X_c_838_n N_X_c_839_n N_X_c_840_n X X X N_X_c_841_n X
+ PM_SKY130_FD_SC_MS__MUX2_4%X
x_PM_SKY130_FD_SC_MS__MUX2_4%A_725_391# N_A_725_391#_M1010_d
+ N_A_725_391#_M1011_d N_A_725_391#_c_895_n N_A_725_391#_c_896_n
+ N_A_725_391#_c_897_n N_A_725_391#_c_898_n
+ PM_SKY130_FD_SC_MS__MUX2_4%A_725_391#
x_PM_SKY130_FD_SC_MS__MUX2_4%A_939_391# N_A_939_391#_M1015_d
+ N_A_939_391#_M1005_d N_A_939_391#_c_941_n N_A_939_391#_c_942_n
+ N_A_939_391#_c_943_n N_A_939_391#_c_944_n N_A_939_391#_c_945_n
+ PM_SKY130_FD_SC_MS__MUX2_4%A_939_391#
x_PM_SKY130_FD_SC_MS__MUX2_4%VGND N_VGND_M1002_d N_VGND_M1012_s N_VGND_M1023_s
+ N_VGND_M1024_s N_VGND_M1007_s N_VGND_c_988_n N_VGND_c_989_n N_VGND_c_990_n
+ N_VGND_c_991_n N_VGND_c_992_n N_VGND_c_993_n N_VGND_c_994_n N_VGND_c_995_n
+ N_VGND_c_996_n N_VGND_c_997_n VGND N_VGND_c_998_n N_VGND_c_999_n
+ N_VGND_c_1000_n N_VGND_c_1001_n N_VGND_c_1002_n N_VGND_c_1003_n
+ N_VGND_c_1004_n PM_SKY130_FD_SC_MS__MUX2_4%VGND
x_PM_SKY130_FD_SC_MS__MUX2_4%A_709_119# N_A_709_119#_M1001_d
+ N_A_709_119#_M1014_s N_A_709_119#_c_1094_n N_A_709_119#_c_1095_n
+ N_A_709_119#_c_1096_n N_A_709_119#_c_1097_n N_A_709_119#_c_1098_n
+ N_A_709_119#_c_1099_n PM_SKY130_FD_SC_MS__MUX2_4%A_709_119#
x_PM_SKY130_FD_SC_MS__MUX2_4%A_937_119# N_A_937_119#_M1003_d
+ N_A_937_119#_M1017_d N_A_937_119#_c_1154_n N_A_937_119#_c_1155_n
+ N_A_937_119#_c_1160_n N_A_937_119#_c_1156_n N_A_937_119#_c_1171_n
+ PM_SKY130_FD_SC_MS__MUX2_4%A_937_119#
cc_1 VNB N_S_M1002_g 0.0294058f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.81
cc_2 VNB N_S_M1001_g 0.0228248f $X=-0.19 $Y=-0.245 $X2=3.47 $Y2=0.915
cc_3 VNB N_S_M1024_g 0.0216899f $X=-0.19 $Y=-0.245 $X2=3.97 $Y2=0.915
cc_4 VNB N_S_c_158_n 0.00152914f $X=-0.19 $Y=-0.245 $X2=3.165 $Y2=1.6
cc_5 VNB N_S_c_159_n 0.00633555f $X=-0.19 $Y=-0.245 $X2=3.58 $Y2=1.6
cc_6 VNB N_S_c_160_n 0.0272156f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.515
cc_7 VNB N_S_c_161_n 0.00610825f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.515
cc_8 VNB N_S_c_162_n 0.0278221f $X=-0.19 $Y=-0.245 $X2=3.985 $Y2=1.6
cc_9 VNB N_A_27_368#_M1003_g 0.0215488f $X=-0.19 $Y=-0.245 $X2=3.535 $Y2=1.765
cc_10 VNB N_A_27_368#_M1007_g 0.0232446f $X=-0.19 $Y=-0.245 $X2=3.97 $Y2=1.435
cc_11 VNB N_A_27_368#_c_293_n 3.75525e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_368#_c_294_n 0.00212795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_368#_c_295_n 0.0447788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_368#_c_296_n 0.0242993f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.68
cc_15 VNB N_A_27_368#_c_297_n 0.0356331f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.665
cc_16 VNB N_A_193_241#_M1000_g 0.00622475f $X=-0.19 $Y=-0.245 $X2=3.985
+ $Y2=1.765
cc_17 VNB N_A_193_241#_M1006_g 0.0119056f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=2.05
cc_18 VNB N_A_193_241#_c_429_n 0.0188836f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=2.135
cc_19 VNB N_A_193_241#_c_430_n 0.0125025f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=2.135
cc_20 VNB N_A_193_241#_c_431_n 0.0059089f $X=-0.19 $Y=-0.245 $X2=2.995 $Y2=2.24
cc_21 VNB N_A_193_241#_M1004_g 0.0126506f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=1.765
cc_22 VNB N_A_193_241#_M1012_g 0.011601f $X=-0.19 $Y=-0.245 $X2=3.58 $Y2=1.6
cc_23 VNB N_A_193_241#_c_434_n 0.0274798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_193_241#_M1021_g 0.0112763f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_25 VNB N_A_193_241#_c_436_n 0.00575367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_193_241#_M1019_g 0.0149832f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.515
cc_27 VNB N_A_193_241#_c_438_n 0.016028f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.35
cc_28 VNB N_A_193_241#_M1023_g 0.0129289f $X=-0.19 $Y=-0.245 $X2=3.58 $Y2=1.6
cc_29 VNB N_A_193_241#_c_440_n 0.219476f $X=-0.19 $Y=-0.245 $X2=3.97 $Y2=1.6
cc_30 VNB N_A_193_241#_c_441_n 0.0261863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_193_241#_M1020_g 0.00887312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_193_241#_c_443_n 0.0853864f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.78
cc_33 VNB N_A_193_241#_c_444_n 0.0201879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_193_241#_c_445_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_193_241#_c_446_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_193_241#_c_447_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_193_241#_c_448_n 0.00467671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_193_241#_c_449_n 0.0313614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_193_241#_c_450_n 0.0026202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_193_241#_c_451_n 0.012433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_193_241#_c_452_n 0.0165854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_193_241#_c_453_n 0.0302575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_193_241#_c_454_n 0.00938153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_193_241#_c_455_n 0.00139572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_193_241#_c_456_n 0.0022133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_193_241#_c_457_n 0.0133735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_193_241#_c_458_n 0.0171429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A0_M1017_g 0.0448307f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.34
cc_49 VNB N_A0_M1022_g 0.0336114f $X=-0.19 $Y=-0.245 $X2=3.47 $Y2=0.915
cc_50 VNB N_A0_c_648_n 0.0251436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A1_M1014_g 0.0337961f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.81
cc_52 VNB N_A1_M1025_g 0.0391319f $X=-0.19 $Y=-0.245 $X2=3.535 $Y2=2.455
cc_53 VNB N_A1_c_692_n 0.00508237f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=2.05
cc_54 VNB N_A1_c_693_n 0.0282231f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=2.135
cc_55 VNB N_VPWR_c_736_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_X_c_837_n 0.00243486f $X=-0.19 $Y=-0.245 $X2=3.535 $Y2=1.765
cc_57 VNB N_X_c_838_n 0.00541625f $X=-0.19 $Y=-0.245 $X2=3.535 $Y2=2.455
cc_58 VNB N_X_c_839_n 7.61737e-19 $X=-0.19 $Y=-0.245 $X2=3.97 $Y2=1.435
cc_59 VNB N_X_c_840_n 0.00215099f $X=-0.19 $Y=-0.245 $X2=3.97 $Y2=0.915
cc_60 VNB N_X_c_841_n 0.00882506f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=2.24
cc_61 VNB N_VGND_c_988_n 0.0228137f $X=-0.19 $Y=-0.245 $X2=3.97 $Y2=0.915
cc_62 VNB N_VGND_c_989_n 0.00298812f $X=-0.19 $Y=-0.245 $X2=3.985 $Y2=2.455
cc_63 VNB N_VGND_c_990_n 0.0157969f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=2.05
cc_64 VNB N_VGND_c_991_n 0.0205418f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=2.24
cc_65 VNB N_VGND_c_992_n 0.0195912f $X=-0.19 $Y=-0.245 $X2=3.58 $Y2=1.6
cc_66 VNB N_VGND_c_993_n 0.0128294f $X=-0.19 $Y=-0.245 $X2=1.59 $Y2=2.135
cc_67 VNB N_VGND_c_994_n 0.0234806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_995_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_69 VNB N_VGND_c_996_n 0.0190194f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_70 VNB N_VGND_c_997_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.515
cc_71 VNB N_VGND_c_998_n 0.0196457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_999_n 0.0171982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1000_n 0.0724602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1001_n 0.434755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1002_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1003_n 0.00625894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1004_n 0.00536684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_709_119#_c_1094_n 0.00267057f $X=-0.19 $Y=-0.245 $X2=3.47
+ $Y2=1.435
cc_79 VNB N_A_709_119#_c_1095_n 0.00289807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_709_119#_c_1096_n 0.0407711f $X=-0.19 $Y=-0.245 $X2=3.535
+ $Y2=1.765
cc_81 VNB N_A_709_119#_c_1097_n 0.00218005f $X=-0.19 $Y=-0.245 $X2=3.97
+ $Y2=1.435
cc_82 VNB N_A_709_119#_c_1098_n 0.00740417f $X=-0.19 $Y=-0.245 $X2=3.97
+ $Y2=0.915
cc_83 VNB N_A_709_119#_c_1099_n 0.00609138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_937_119#_c_1154_n 0.00160098f $X=-0.19 $Y=-0.245 $X2=3.47
+ $Y2=1.435
cc_85 VNB N_A_937_119#_c_1155_n 0.00224578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_937_119#_c_1156_n 0.00151525f $X=-0.19 $Y=-0.245 $X2=3.97
+ $Y2=1.435
cc_87 VPB N_S_M1009_g 0.0257961f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.34
cc_88 VPB N_S_M1010_g 0.0250865f $X=-0.19 $Y=1.66 $X2=3.535 $Y2=2.455
cc_89 VPB N_S_M1013_g 0.0240397f $X=-0.19 $Y=1.66 $X2=3.985 $Y2=2.455
cc_90 VPB N_S_c_166_n 8.59789e-19 $X=-0.19 $Y=1.66 $X2=0.75 $Y2=2.05
cc_91 VPB N_S_c_167_n 7.75131e-19 $X=-0.19 $Y=1.66 $X2=3.08 $Y2=2.155
cc_92 VPB N_S_c_159_n 0.00697023f $X=-0.19 $Y=1.66 $X2=3.58 $Y2=1.6
cc_93 VPB N_S_c_160_n 0.005975f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.515
cc_94 VPB N_S_c_161_n 0.00195922f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.515
cc_95 VPB N_S_c_162_n 0.0140668f $X=-0.19 $Y=1.66 $X2=3.985 $Y2=1.6
cc_96 VPB N_A_27_368#_M1015_g 0.0253068f $X=-0.19 $Y=1.66 $X2=3.47 $Y2=1.435
cc_97 VPB N_A_27_368#_M1018_g 0.0289604f $X=-0.19 $Y=1.66 $X2=3.985 $Y2=1.765
cc_98 VPB N_A_27_368#_c_300_n 0.0101859f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=2.05
cc_99 VPB N_A_27_368#_c_301_n 0.0226151f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=2.135
cc_100 VPB N_A_27_368#_c_302_n 0.00331455f $X=-0.19 $Y=1.66 $X2=3.165 $Y2=1.6
cc_101 VPB N_A_27_368#_c_303_n 0.00100408f $X=-0.19 $Y=1.66 $X2=3.58 $Y2=1.6
cc_102 VPB N_A_27_368#_c_304_n 0.00202119f $X=-0.19 $Y=1.66 $X2=3.58 $Y2=1.6
cc_103 VPB N_A_27_368#_c_294_n 0.00390775f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_27_368#_c_306_n 0.00710642f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.35
cc_105 VPB N_A_27_368#_c_296_n 0.0126837f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.68
cc_106 VPB N_A_27_368#_c_297_n 0.0213701f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.665
cc_107 VPB N_A_193_241#_M1000_g 0.0359259f $X=-0.19 $Y=1.66 $X2=3.985 $Y2=1.765
cc_108 VPB N_A_193_241#_M1004_g 0.0326126f $X=-0.19 $Y=1.66 $X2=3.08 $Y2=1.765
cc_109 VPB N_A_193_241#_M1019_g 0.0294803f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.515
cc_110 VPB N_A_193_241#_M1020_g 0.0283526f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_193_241#_c_448_n 0.00179237f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_193_241#_c_449_n 0.0266663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_193_241#_c_465_n 0.00737845f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_193_241#_c_466_n 0.0108831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_193_241#_c_467_n 0.00724744f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_193_241#_c_468_n 0.0327257f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_193_241#_c_453_n 0.0139254f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_193_241#_c_470_n 0.0169387f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_193_241#_c_458_n 0.017241f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A0_M1011_g 0.0269203f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=0.81
cc_121 VPB N_A0_M1016_g 0.0229491f $X=-0.19 $Y=1.66 $X2=3.535 $Y2=2.455
cc_122 VPB N_A0_c_648_n 0.0145222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A1_M1005_g 0.022963f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.34
cc_124 VPB N_A1_M1008_g 0.0281372f $X=-0.19 $Y=1.66 $X2=3.47 $Y2=0.915
cc_125 VPB N_A1_c_692_n 0.00361007f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=2.05
cc_126 VPB N_A1_c_693_n 0.0164486f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=2.135
cc_127 VPB N_VPWR_c_737_n 0.0110391f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_738_n 0.00799777f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_739_n 0.00799536f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=2.135
cc_130 VPB N_VPWR_c_740_n 0.00867756f $X=-0.19 $Y=1.66 $X2=3.08 $Y2=2.155
cc_131 VPB N_VPWR_c_741_n 0.00686253f $X=-0.19 $Y=1.66 $X2=3.58 $Y2=1.6
cc_132 VPB N_VPWR_c_742_n 0.0232884f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_743_n 0.00631622f $X=-0.19 $Y=1.66 $X2=1.59 $Y2=2.24
cc_134 VPB N_VPWR_c_744_n 0.0203178f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_135 VPB N_VPWR_c_745_n 0.00631953f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_746_n 0.0207444f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.515
cc_137 VPB N_VPWR_c_747_n 0.00478125f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.515
cc_138 VPB N_VPWR_c_748_n 0.025094f $X=-0.19 $Y=1.66 $X2=3.97 $Y2=1.6
cc_139 VPB N_VPWR_c_749_n 0.0862348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_736_n 0.0941944f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_751_n 0.0270156f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_752_n 0.00631622f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_X_c_837_n 5.32607e-19 $X=-0.19 $Y=1.66 $X2=3.535 $Y2=1.765
cc_144 VPB N_X_c_839_n 0.00278012f $X=-0.19 $Y=1.66 $X2=3.97 $Y2=1.435
cc_145 VPB N_X_c_841_n 7.84116e-19 $X=-0.19 $Y=1.66 $X2=1.675 $Y2=2.24
cc_146 VPB N_A_725_391#_c_895_n 0.00357339f $X=-0.19 $Y=1.66 $X2=3.47 $Y2=1.435
cc_147 VPB N_A_725_391#_c_896_n 0.0210801f $X=-0.19 $Y=1.66 $X2=3.535 $Y2=1.765
cc_148 VPB N_A_725_391#_c_897_n 0.00205552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_725_391#_c_898_n 0.0177038f $X=-0.19 $Y=1.66 $X2=3.97 $Y2=1.435
cc_150 VPB N_A_939_391#_c_941_n 0.0116868f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=0.81
cc_151 VPB N_A_939_391#_c_942_n 0.00548534f $X=-0.19 $Y=1.66 $X2=3.47 $Y2=1.435
cc_152 VPB N_A_939_391#_c_943_n 0.00221956f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_939_391#_c_944_n 0.0162501f $X=-0.19 $Y=1.66 $X2=3.97 $Y2=1.435
cc_154 VPB N_A_939_391#_c_945_n 0.00231152f $X=-0.19 $Y=1.66 $X2=3.985 $Y2=2.455
cc_155 N_S_M1013_g N_A_27_368#_M1015_g 0.0324544f $X=3.985 $Y=2.455 $X2=0 $Y2=0
cc_156 N_S_M1024_g N_A_27_368#_M1003_g 0.0210679f $X=3.97 $Y=0.915 $X2=0 $Y2=0
cc_157 N_S_M1009_g N_A_27_368#_c_300_n 0.00624542f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_158 N_S_M1009_g N_A_27_368#_c_312_n 0.0120277f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_159 N_S_c_176_p N_A_27_368#_c_312_n 0.0174664f $X=1.505 $Y=2.135 $X2=0 $Y2=0
cc_160 N_S_c_177_p N_A_27_368#_c_312_n 0.0137412f $X=0.835 $Y=2.135 $X2=0 $Y2=0
cc_161 N_S_c_161_n N_A_27_368#_c_312_n 0.00522503f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_162 N_S_M1009_g N_A_27_368#_c_301_n 0.0086473f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_163 N_S_M1010_g N_A_27_368#_c_317_n 0.00638734f $X=3.535 $Y=2.455 $X2=0 $Y2=0
cc_164 N_S_c_176_p N_A_27_368#_c_317_n 0.00866703f $X=1.505 $Y=2.135 $X2=0 $Y2=0
cc_165 N_S_c_182_p N_A_27_368#_c_317_n 0.0862432f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_166 N_S_c_183_p N_A_27_368#_c_317_n 0.00796293f $X=1.59 $Y=2.135 $X2=0 $Y2=0
cc_167 N_S_M1010_g N_A_27_368#_c_321_n 0.0100402f $X=3.535 $Y=2.455 $X2=0 $Y2=0
cc_168 N_S_M1013_g N_A_27_368#_c_321_n 7.93935e-19 $X=3.985 $Y=2.455 $X2=0 $Y2=0
cc_169 N_S_c_182_p N_A_27_368#_c_321_n 0.0138308f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_170 N_S_c_167_n N_A_27_368#_c_321_n 0.00355899f $X=3.08 $Y=2.155 $X2=0 $Y2=0
cc_171 N_S_M1010_g N_A_27_368#_c_302_n 0.0106802f $X=3.535 $Y=2.455 $X2=0 $Y2=0
cc_172 N_S_M1013_g N_A_27_368#_c_302_n 0.00992587f $X=3.985 $Y=2.455 $X2=0 $Y2=0
cc_173 N_S_c_159_n N_A_27_368#_c_302_n 0.0175559f $X=3.58 $Y=1.6 $X2=0 $Y2=0
cc_174 N_S_c_162_n N_A_27_368#_c_302_n 0.00231283f $X=3.985 $Y=1.6 $X2=0 $Y2=0
cc_175 N_S_M1010_g N_A_27_368#_c_303_n 0.00345703f $X=3.535 $Y=2.455 $X2=0 $Y2=0
cc_176 N_S_c_167_n N_A_27_368#_c_303_n 0.0138661f $X=3.08 $Y=2.155 $X2=0 $Y2=0
cc_177 N_S_c_159_n N_A_27_368#_c_303_n 0.0143138f $X=3.58 $Y=1.6 $X2=0 $Y2=0
cc_178 N_S_c_162_n N_A_27_368#_c_303_n 0.00136199f $X=3.985 $Y=1.6 $X2=0 $Y2=0
cc_179 N_S_M1010_g N_A_27_368#_c_304_n 0.00104675f $X=3.535 $Y=2.455 $X2=0 $Y2=0
cc_180 N_S_M1013_g N_A_27_368#_c_304_n 0.00576f $X=3.985 $Y=2.455 $X2=0 $Y2=0
cc_181 N_S_c_159_n N_A_27_368#_c_293_n 0.0277655f $X=3.58 $Y=1.6 $X2=0 $Y2=0
cc_182 N_S_c_162_n N_A_27_368#_c_293_n 0.0150349f $X=3.985 $Y=1.6 $X2=0 $Y2=0
cc_183 N_S_M1002_g N_A_27_368#_c_295_n 0.00855288f $X=0.65 $Y=0.81 $X2=0 $Y2=0
cc_184 N_S_c_160_n N_A_27_368#_c_295_n 0.00164811f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_185 N_S_c_161_n N_A_27_368#_c_295_n 0.013094f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_186 N_S_M1009_g N_A_27_368#_c_306_n 0.00299985f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_187 N_S_c_166_n N_A_27_368#_c_306_n 0.00606514f $X=0.75 $Y=2.05 $X2=0 $Y2=0
cc_188 N_S_c_177_p N_A_27_368#_c_306_n 0.0115465f $X=0.835 $Y=2.135 $X2=0 $Y2=0
cc_189 N_S_c_161_n N_A_27_368#_c_306_n 0.00147239f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_190 N_S_M1002_g N_A_27_368#_c_296_n 0.00436189f $X=0.65 $Y=0.81 $X2=0 $Y2=0
cc_191 N_S_c_166_n N_A_27_368#_c_296_n 0.00470078f $X=0.75 $Y=2.05 $X2=0 $Y2=0
cc_192 N_S_c_160_n N_A_27_368#_c_296_n 0.0122425f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_193 N_S_c_161_n N_A_27_368#_c_296_n 0.032823f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_194 N_S_c_176_p N_A_27_368#_c_348_n 0.00999494f $X=1.505 $Y=2.135 $X2=0 $Y2=0
cc_195 N_S_c_162_n N_A_27_368#_c_297_n 0.0183107f $X=3.985 $Y=1.6 $X2=0 $Y2=0
cc_196 N_S_M1009_g N_A_193_241#_M1000_g 0.0321131f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_197 N_S_c_166_n N_A_193_241#_M1000_g 0.0039804f $X=0.75 $Y=2.05 $X2=0 $Y2=0
cc_198 N_S_c_176_p N_A_193_241#_M1000_g 0.0159432f $X=1.505 $Y=2.135 $X2=0 $Y2=0
cc_199 N_S_c_183_p N_A_193_241#_M1000_g 0.00201814f $X=1.59 $Y=2.135 $X2=0 $Y2=0
cc_200 N_S_M1002_g N_A_193_241#_M1006_g 0.0166337f $X=0.65 $Y=0.81 $X2=0 $Y2=0
cc_201 N_S_c_176_p N_A_193_241#_M1004_g 3.99741e-19 $X=1.505 $Y=2.135 $X2=0
+ $Y2=0
cc_202 N_S_c_182_p N_A_193_241#_M1004_g 0.00757545f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_203 N_S_c_183_p N_A_193_241#_M1004_g 0.00940567f $X=1.59 $Y=2.135 $X2=0 $Y2=0
cc_204 N_S_c_182_p N_A_193_241#_M1019_g 0.0140996f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_205 N_S_c_167_n N_A_193_241#_M1019_g 8.30962e-19 $X=3.08 $Y=2.155 $X2=0 $Y2=0
cc_206 N_S_c_158_n N_A_193_241#_M1019_g 2.07883e-19 $X=3.165 $Y=1.6 $X2=0 $Y2=0
cc_207 N_S_c_183_p N_A_193_241#_M1019_g 6.06311e-19 $X=1.59 $Y=2.135 $X2=0 $Y2=0
cc_208 N_S_M1001_g N_A_193_241#_M1023_g 0.00801147f $X=3.47 $Y=0.915 $X2=0 $Y2=0
cc_209 N_S_M1001_g N_A_193_241#_c_440_n 0.0103003f $X=3.47 $Y=0.915 $X2=0 $Y2=0
cc_210 N_S_M1024_g N_A_193_241#_c_440_n 0.0103107f $X=3.97 $Y=0.915 $X2=0 $Y2=0
cc_211 N_S_M1001_g N_A_193_241#_c_441_n 0.00703294f $X=3.47 $Y=0.915 $X2=0 $Y2=0
cc_212 N_S_c_182_p N_A_193_241#_c_441_n 9.15503e-19 $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_213 N_S_c_158_n N_A_193_241#_c_441_n 9.10335e-19 $X=3.165 $Y=1.6 $X2=0 $Y2=0
cc_214 N_S_M1010_g N_A_193_241#_M1020_g 0.0306142f $X=3.535 $Y=2.455 $X2=0 $Y2=0
cc_215 N_S_c_182_p N_A_193_241#_M1020_g 0.0174187f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_216 N_S_c_167_n N_A_193_241#_M1020_g 0.00988809f $X=3.08 $Y=2.155 $X2=0 $Y2=0
cc_217 N_S_c_158_n N_A_193_241#_M1020_g 0.00816553f $X=3.165 $Y=1.6 $X2=0 $Y2=0
cc_218 N_S_c_162_n N_A_193_241#_M1020_g 0.00703294f $X=3.985 $Y=1.6 $X2=0 $Y2=0
cc_219 N_S_M1002_g N_A_193_241#_c_444_n 0.00854554f $X=0.65 $Y=0.81 $X2=0 $Y2=0
cc_220 N_S_c_160_n N_A_193_241#_c_444_n 0.0196459f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_221 N_S_c_161_n N_A_193_241#_c_444_n 0.0039804f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_222 N_S_c_166_n N_VPWR_M1009_d 0.00511674f $X=0.75 $Y=2.05 $X2=-0.19
+ $Y2=-0.245
cc_223 N_S_c_176_p N_VPWR_M1009_d 0.00351444f $X=1.505 $Y=2.135 $X2=-0.19
+ $Y2=-0.245
cc_224 N_S_c_177_p N_VPWR_M1009_d 0.00453484f $X=0.835 $Y=2.135 $X2=-0.19
+ $Y2=-0.245
cc_225 N_S_c_182_p N_VPWR_M1004_s 0.00853823f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_226 N_S_c_182_p N_VPWR_M1020_s 0.00267546f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_227 N_S_c_167_n N_VPWR_M1020_s 0.00310809f $X=3.08 $Y=2.155 $X2=0 $Y2=0
cc_228 N_S_M1009_g N_VPWR_c_737_n 0.0039575f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_229 N_S_M1010_g N_VPWR_c_739_n 0.00422816f $X=3.535 $Y=2.455 $X2=0 $Y2=0
cc_230 N_S_M1013_g N_VPWR_c_740_n 0.00459019f $X=3.985 $Y=2.455 $X2=0 $Y2=0
cc_231 N_S_M1010_g N_VPWR_c_744_n 0.00496376f $X=3.535 $Y=2.455 $X2=0 $Y2=0
cc_232 N_S_M1013_g N_VPWR_c_744_n 0.00391326f $X=3.985 $Y=2.455 $X2=0 $Y2=0
cc_233 N_S_M1009_g N_VPWR_c_736_n 0.00610055f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_234 N_S_M1010_g N_VPWR_c_736_n 0.00653145f $X=3.535 $Y=2.455 $X2=0 $Y2=0
cc_235 N_S_M1013_g N_VPWR_c_736_n 0.00653145f $X=3.985 $Y=2.455 $X2=0 $Y2=0
cc_236 N_S_M1009_g N_VPWR_c_751_n 0.00567028f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_237 N_S_c_176_p N_X_M1000_d 0.0079533f $X=1.505 $Y=2.135 $X2=0 $Y2=0
cc_238 N_S_c_183_p N_X_M1000_d 0.00234678f $X=1.59 $Y=2.135 $X2=0 $Y2=0
cc_239 N_S_c_182_p N_X_M1019_d 0.00759035f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_240 N_S_c_176_p N_X_c_837_n 0.0289114f $X=1.505 $Y=2.135 $X2=0 $Y2=0
cc_241 N_S_c_183_p N_X_c_837_n 0.00617282f $X=1.59 $Y=2.135 $X2=0 $Y2=0
cc_242 N_S_c_160_n N_X_c_837_n 2.82822e-19 $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_243 N_S_c_161_n N_X_c_837_n 0.0320616f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_244 N_S_c_161_n N_X_c_838_n 8.05573e-19 $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_245 N_S_M1001_g N_X_c_839_n 2.44849e-19 $X=3.47 $Y=0.915 $X2=0 $Y2=0
cc_246 N_S_c_182_p N_X_c_839_n 0.0292685f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_247 N_S_c_167_n N_X_c_839_n 0.00878443f $X=3.08 $Y=2.155 $X2=0 $Y2=0
cc_248 N_S_c_158_n N_X_c_839_n 0.0227181f $X=3.165 $Y=1.6 $X2=0 $Y2=0
cc_249 N_S_M1001_g N_X_c_840_n 0.00101895f $X=3.47 $Y=0.915 $X2=0 $Y2=0
cc_250 N_S_c_182_p N_X_c_841_n 0.0289077f $X=2.995 $Y=2.24 $X2=0 $Y2=0
cc_251 N_S_c_183_p N_X_c_841_n 0.00257766f $X=1.59 $Y=2.135 $X2=0 $Y2=0
cc_252 N_S_M1013_g N_A_725_391#_c_895_n 0.0116375f $X=3.985 $Y=2.455 $X2=0 $Y2=0
cc_253 N_S_M1013_g N_A_725_391#_c_897_n 0.0107236f $X=3.985 $Y=2.455 $X2=0 $Y2=0
cc_254 N_S_M1013_g N_A_939_391#_c_943_n 8.64576e-19 $X=3.985 $Y=2.455 $X2=0
+ $Y2=0
cc_255 N_S_M1002_g N_VGND_c_988_n 0.0074703f $X=0.65 $Y=0.81 $X2=0 $Y2=0
cc_256 N_S_c_161_n N_VGND_c_988_n 0.00525943f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_257 N_S_M1001_g N_VGND_c_990_n 0.0108034f $X=3.47 $Y=0.915 $X2=0 $Y2=0
cc_258 N_S_c_158_n N_VGND_c_990_n 0.0152459f $X=3.165 $Y=1.6 $X2=0 $Y2=0
cc_259 N_S_c_159_n N_VGND_c_990_n 0.00752017f $X=3.58 $Y=1.6 $X2=0 $Y2=0
cc_260 N_S_M1001_g N_VGND_c_992_n 6.03908e-19 $X=3.47 $Y=0.915 $X2=0 $Y2=0
cc_261 N_S_M1024_g N_VGND_c_992_n 0.0133679f $X=3.97 $Y=0.915 $X2=0 $Y2=0
cc_262 N_S_M1002_g N_VGND_c_994_n 0.00473385f $X=0.65 $Y=0.81 $X2=0 $Y2=0
cc_263 N_S_M1002_g N_VGND_c_1001_n 0.00508379f $X=0.65 $Y=0.81 $X2=0 $Y2=0
cc_264 N_S_M1001_g N_VGND_c_1001_n 9.39239e-19 $X=3.47 $Y=0.915 $X2=0 $Y2=0
cc_265 N_S_M1024_g N_VGND_c_1001_n 7.88961e-19 $X=3.97 $Y=0.915 $X2=0 $Y2=0
cc_266 N_S_M1001_g N_A_709_119#_c_1094_n 0.00735844f $X=3.47 $Y=0.915 $X2=0
+ $Y2=0
cc_267 N_S_M1024_g N_A_709_119#_c_1094_n 0.00277359f $X=3.97 $Y=0.915 $X2=0
+ $Y2=0
cc_268 N_S_M1001_g N_A_709_119#_c_1095_n 0.00334323f $X=3.47 $Y=0.915 $X2=0
+ $Y2=0
cc_269 N_S_c_159_n N_A_709_119#_c_1095_n 0.0188868f $X=3.58 $Y=1.6 $X2=0 $Y2=0
cc_270 N_S_c_162_n N_A_709_119#_c_1095_n 0.00467964f $X=3.985 $Y=1.6 $X2=0 $Y2=0
cc_271 N_S_M1024_g N_A_709_119#_c_1098_n 0.0157636f $X=3.97 $Y=0.915 $X2=0 $Y2=0
cc_272 N_S_c_162_n N_A_709_119#_c_1098_n 2.0866e-19 $X=3.985 $Y=1.6 $X2=0 $Y2=0
cc_273 N_S_M1024_g N_A_937_119#_c_1155_n 2.92953e-19 $X=3.97 $Y=0.915 $X2=0
+ $Y2=0
cc_274 N_A_27_368#_c_300_n N_A_193_241#_M1000_g 7.78621e-19 $X=0.265 $Y=2.39
+ $X2=0 $Y2=0
cc_275 N_A_27_368#_c_312_n N_A_193_241#_M1000_g 0.0125257f $X=1.165 $Y=2.475
+ $X2=0 $Y2=0
cc_276 N_A_27_368#_c_301_n N_A_193_241#_M1000_g 5.17124e-19 $X=0.445 $Y=2.475
+ $X2=0 $Y2=0
cc_277 N_A_27_368#_c_317_n N_A_193_241#_M1004_g 0.0142782f $X=3.335 $Y=2.58
+ $X2=0 $Y2=0
cc_278 N_A_27_368#_c_348_n N_A_193_241#_M1004_g 0.0023389f $X=1.25 $Y=2.475
+ $X2=0 $Y2=0
cc_279 N_A_27_368#_c_317_n N_A_193_241#_M1019_g 0.0149641f $X=3.335 $Y=2.58
+ $X2=0 $Y2=0
cc_280 N_A_27_368#_M1003_g N_A_193_241#_c_440_n 0.0103003f $X=4.61 $Y=0.915
+ $X2=0 $Y2=0
cc_281 N_A_27_368#_M1007_g N_A_193_241#_c_440_n 0.00991298f $X=5.04 $Y=0.915
+ $X2=0 $Y2=0
cc_282 N_A_27_368#_c_317_n N_A_193_241#_M1020_g 0.0149124f $X=3.335 $Y=2.58
+ $X2=0 $Y2=0
cc_283 N_A_27_368#_c_321_n N_A_193_241#_M1020_g 0.00366232f $X=3.42 $Y=2.495
+ $X2=0 $Y2=0
cc_284 N_A_27_368#_c_303_n N_A_193_241#_M1020_g 5.23016e-19 $X=3.505 $Y=2.02
+ $X2=0 $Y2=0
cc_285 N_A_27_368#_M1007_g N_A_193_241#_c_443_n 0.0193743f $X=5.04 $Y=0.915
+ $X2=0 $Y2=0
cc_286 N_A_27_368#_c_294_n N_A_193_241#_c_448_n 0.0132241f $X=4.82 $Y=1.6 $X2=0
+ $Y2=0
cc_287 N_A_27_368#_c_297_n N_A_193_241#_c_448_n 0.00154423f $X=5.055 $Y=1.6
+ $X2=0 $Y2=0
cc_288 N_A_27_368#_c_294_n N_A_193_241#_c_458_n 3.11698e-19 $X=4.82 $Y=1.6 $X2=0
+ $Y2=0
cc_289 N_A_27_368#_c_297_n N_A_193_241#_c_458_n 0.0186824f $X=5.055 $Y=1.6 $X2=0
+ $Y2=0
cc_290 N_A_27_368#_c_312_n N_VPWR_M1009_d 0.00558527f $X=1.165 $Y=2.475
+ $X2=-0.19 $Y2=-0.245
cc_291 N_A_27_368#_c_317_n N_VPWR_M1004_s 0.00756667f $X=3.335 $Y=2.58 $X2=0
+ $Y2=0
cc_292 N_A_27_368#_c_317_n N_VPWR_M1020_s 0.0116374f $X=3.335 $Y=2.58 $X2=0
+ $Y2=0
cc_293 N_A_27_368#_c_321_n N_VPWR_M1020_s 0.00417874f $X=3.42 $Y=2.495 $X2=0
+ $Y2=0
cc_294 N_A_27_368#_c_303_n N_VPWR_M1020_s 0.00138996f $X=3.505 $Y=2.02 $X2=0
+ $Y2=0
cc_295 N_A_27_368#_c_312_n N_VPWR_c_737_n 0.022352f $X=1.165 $Y=2.475 $X2=0
+ $Y2=0
cc_296 N_A_27_368#_c_301_n N_VPWR_c_737_n 0.00497591f $X=0.445 $Y=2.475 $X2=0
+ $Y2=0
cc_297 N_A_27_368#_c_317_n N_VPWR_c_738_n 0.0250819f $X=3.335 $Y=2.58 $X2=0
+ $Y2=0
cc_298 N_A_27_368#_c_317_n N_VPWR_c_739_n 0.0254753f $X=3.335 $Y=2.58 $X2=0
+ $Y2=0
cc_299 N_A_27_368#_M1015_g N_VPWR_c_740_n 0.00495234f $X=4.605 $Y=2.455 $X2=0
+ $Y2=0
cc_300 N_A_27_368#_M1018_g N_VPWR_c_741_n 0.00896155f $X=5.055 $Y=2.455 $X2=0
+ $Y2=0
cc_301 N_A_27_368#_c_317_n N_VPWR_c_742_n 0.00690659f $X=3.335 $Y=2.58 $X2=0
+ $Y2=0
cc_302 N_A_27_368#_c_348_n N_VPWR_c_742_n 0.0025644f $X=1.25 $Y=2.475 $X2=0
+ $Y2=0
cc_303 N_A_27_368#_c_317_n N_VPWR_c_744_n 0.00149501f $X=3.335 $Y=2.58 $X2=0
+ $Y2=0
cc_304 N_A_27_368#_M1015_g N_VPWR_c_746_n 0.0039878f $X=4.605 $Y=2.455 $X2=0
+ $Y2=0
cc_305 N_A_27_368#_M1018_g N_VPWR_c_746_n 0.0039878f $X=5.055 $Y=2.455 $X2=0
+ $Y2=0
cc_306 N_A_27_368#_c_317_n N_VPWR_c_748_n 0.0128314f $X=3.335 $Y=2.58 $X2=0
+ $Y2=0
cc_307 N_A_27_368#_M1015_g N_VPWR_c_736_n 0.00653145f $X=4.605 $Y=2.455 $X2=0
+ $Y2=0
cc_308 N_A_27_368#_M1018_g N_VPWR_c_736_n 0.00653145f $X=5.055 $Y=2.455 $X2=0
+ $Y2=0
cc_309 N_A_27_368#_c_312_n N_VPWR_c_736_n 0.0134442f $X=1.165 $Y=2.475 $X2=0
+ $Y2=0
cc_310 N_A_27_368#_c_301_n N_VPWR_c_736_n 0.0122603f $X=0.445 $Y=2.475 $X2=0
+ $Y2=0
cc_311 N_A_27_368#_c_317_n N_VPWR_c_736_n 0.0423238f $X=3.335 $Y=2.58 $X2=0
+ $Y2=0
cc_312 N_A_27_368#_c_348_n N_VPWR_c_736_n 0.00478779f $X=1.25 $Y=2.475 $X2=0
+ $Y2=0
cc_313 N_A_27_368#_c_301_n N_VPWR_c_751_n 0.010702f $X=0.445 $Y=2.475 $X2=0
+ $Y2=0
cc_314 N_A_27_368#_c_317_n N_X_M1000_d 0.00702265f $X=3.335 $Y=2.58 $X2=0 $Y2=0
cc_315 N_A_27_368#_c_348_n N_X_M1000_d 0.00570046f $X=1.25 $Y=2.475 $X2=0 $Y2=0
cc_316 N_A_27_368#_c_317_n N_X_M1019_d 0.0100898f $X=3.335 $Y=2.58 $X2=0 $Y2=0
cc_317 N_A_27_368#_c_302_n N_A_725_391#_M1010_d 0.00165831f $X=3.915 $Y=2.02
+ $X2=-0.19 $Y2=-0.245
cc_318 N_A_27_368#_M1015_g N_A_725_391#_c_895_n 0.016645f $X=4.605 $Y=2.455
+ $X2=0 $Y2=0
cc_319 N_A_27_368#_M1018_g N_A_725_391#_c_895_n 0.0153685f $X=5.055 $Y=2.455
+ $X2=0 $Y2=0
cc_320 N_A_27_368#_c_302_n N_A_725_391#_c_895_n 0.00667344f $X=3.915 $Y=2.02
+ $X2=0 $Y2=0
cc_321 N_A_27_368#_c_294_n N_A_725_391#_c_895_n 0.0136596f $X=4.82 $Y=1.6 $X2=0
+ $Y2=0
cc_322 N_A_27_368#_c_297_n N_A_725_391#_c_895_n 0.00285921f $X=5.055 $Y=1.6
+ $X2=0 $Y2=0
cc_323 N_A_27_368#_M1015_g N_A_725_391#_c_897_n 0.00151074f $X=4.605 $Y=2.455
+ $X2=0 $Y2=0
cc_324 N_A_27_368#_c_302_n N_A_725_391#_c_897_n 0.0150202f $X=3.915 $Y=2.02
+ $X2=0 $Y2=0
cc_325 N_A_27_368#_M1018_g N_A_725_391#_c_898_n 0.00500066f $X=5.055 $Y=2.455
+ $X2=0 $Y2=0
cc_326 N_A_27_368#_M1018_g N_A_939_391#_c_941_n 0.00413049f $X=5.055 $Y=2.455
+ $X2=0 $Y2=0
cc_327 N_A_27_368#_M1015_g N_A_939_391#_c_943_n 0.00817393f $X=4.605 $Y=2.455
+ $X2=0 $Y2=0
cc_328 N_A_27_368#_M1018_g N_A_939_391#_c_943_n 0.0193943f $X=5.055 $Y=2.455
+ $X2=0 $Y2=0
cc_329 N_A_27_368#_c_302_n N_A_939_391#_c_943_n 0.00281074f $X=3.915 $Y=2.02
+ $X2=0 $Y2=0
cc_330 N_A_27_368#_c_294_n N_A_939_391#_c_943_n 0.0251231f $X=4.82 $Y=1.6 $X2=0
+ $Y2=0
cc_331 N_A_27_368#_c_297_n N_A_939_391#_c_943_n 0.00205041f $X=5.055 $Y=1.6
+ $X2=0 $Y2=0
cc_332 N_A_27_368#_c_295_n N_VGND_c_988_n 0.0288933f $X=0.435 $Y=0.635 $X2=0
+ $Y2=0
cc_333 N_A_27_368#_M1003_g N_VGND_c_992_n 0.00585775f $X=4.61 $Y=0.915 $X2=0
+ $Y2=0
cc_334 N_A_27_368#_M1007_g N_VGND_c_993_n 0.00351782f $X=5.04 $Y=0.915 $X2=0
+ $Y2=0
cc_335 N_A_27_368#_c_295_n N_VGND_c_994_n 0.0153192f $X=0.435 $Y=0.635 $X2=0
+ $Y2=0
cc_336 N_A_27_368#_M1003_g N_VGND_c_1001_n 9.39239e-19 $X=4.61 $Y=0.915 $X2=0
+ $Y2=0
cc_337 N_A_27_368#_M1007_g N_VGND_c_1001_n 9.39239e-19 $X=5.04 $Y=0.915 $X2=0
+ $Y2=0
cc_338 N_A_27_368#_c_295_n N_VGND_c_1001_n 0.0175003f $X=0.435 $Y=0.635 $X2=0
+ $Y2=0
cc_339 N_A_27_368#_c_302_n N_A_709_119#_c_1095_n 0.00336384f $X=3.915 $Y=2.02
+ $X2=0 $Y2=0
cc_340 N_A_27_368#_M1003_g N_A_709_119#_c_1098_n 0.0150485f $X=4.61 $Y=0.915
+ $X2=0 $Y2=0
cc_341 N_A_27_368#_M1007_g N_A_709_119#_c_1098_n 0.0133803f $X=5.04 $Y=0.915
+ $X2=0 $Y2=0
cc_342 N_A_27_368#_c_302_n N_A_709_119#_c_1098_n 0.00170556f $X=3.915 $Y=2.02
+ $X2=0 $Y2=0
cc_343 N_A_27_368#_c_293_n N_A_709_119#_c_1098_n 0.0131287f $X=4.085 $Y=1.6
+ $X2=0 $Y2=0
cc_344 N_A_27_368#_c_294_n N_A_709_119#_c_1098_n 0.0679154f $X=4.82 $Y=1.6 $X2=0
+ $Y2=0
cc_345 N_A_27_368#_c_297_n N_A_709_119#_c_1098_n 0.00828243f $X=5.055 $Y=1.6
+ $X2=0 $Y2=0
cc_346 N_A_27_368#_M1007_g N_A_709_119#_c_1099_n 4.91777e-19 $X=5.04 $Y=0.915
+ $X2=0 $Y2=0
cc_347 N_A_27_368#_M1003_g N_A_937_119#_c_1155_n 0.00472551f $X=4.61 $Y=0.915
+ $X2=0 $Y2=0
cc_348 N_A_27_368#_M1007_g N_A_937_119#_c_1155_n 0.00553184f $X=5.04 $Y=0.915
+ $X2=0 $Y2=0
cc_349 N_A_27_368#_M1007_g N_A_937_119#_c_1160_n 0.0101743f $X=5.04 $Y=0.915
+ $X2=0 $Y2=0
cc_350 N_A_27_368#_M1007_g N_A_937_119#_c_1156_n 3.25189e-19 $X=5.04 $Y=0.915
+ $X2=0 $Y2=0
cc_351 N_A_193_241#_c_450_n N_A0_M1017_g 0.0121398f $X=7.26 $Y=0.34 $X2=0 $Y2=0
cc_352 N_A_193_241#_c_465_n N_A0_M1011_g 0.00592185f $X=6.385 $Y=1.95 $X2=0
+ $Y2=0
cc_353 N_A_193_241#_c_466_n N_A0_M1011_g 0.0122909f $X=8.195 $Y=2.075 $X2=0
+ $Y2=0
cc_354 N_A_193_241#_c_450_n N_A0_M1022_g 0.013161f $X=7.26 $Y=0.34 $X2=0 $Y2=0
cc_355 N_A_193_241#_c_466_n N_A0_M1016_g 0.0147743f $X=8.195 $Y=2.075 $X2=0
+ $Y2=0
cc_356 N_A_193_241#_c_448_n A0 0.02833f $X=6.3 $Y=1.615 $X2=0 $Y2=0
cc_357 N_A_193_241#_c_449_n A0 3.51297e-19 $X=6.23 $Y=1.615 $X2=0 $Y2=0
cc_358 N_A_193_241#_c_466_n A0 0.0329931f $X=8.195 $Y=2.075 $X2=0 $Y2=0
cc_359 N_A_193_241#_c_448_n N_A0_c_648_n 0.00239229f $X=6.3 $Y=1.615 $X2=0 $Y2=0
cc_360 N_A_193_241#_c_449_n N_A0_c_648_n 0.0182643f $X=6.23 $Y=1.615 $X2=0 $Y2=0
cc_361 N_A_193_241#_c_466_n N_A0_c_648_n 0.00203619f $X=8.195 $Y=2.075 $X2=0
+ $Y2=0
cc_362 N_A_193_241#_c_466_n N_A1_M1005_g 0.0121406f $X=8.195 $Y=2.075 $X2=0
+ $Y2=0
cc_363 N_A_193_241#_c_526_p N_A1_M1014_g 0.00708055f $X=7.425 $Y=0.495 $X2=0
+ $Y2=0
cc_364 N_A_193_241#_c_451_n N_A1_M1014_g 0.0102487f $X=8.19 $Y=0.34 $X2=0 $Y2=0
cc_365 N_A_193_241#_c_456_n N_A1_M1014_g 0.00203192f $X=7.425 $Y=0.34 $X2=0
+ $Y2=0
cc_366 N_A_193_241#_c_466_n N_A1_M1008_g 0.0170307f $X=8.195 $Y=2.075 $X2=0
+ $Y2=0
cc_367 N_A_193_241#_c_468_n N_A1_M1008_g 4.8138e-19 $X=8.36 $Y=2.465 $X2=0 $Y2=0
cc_368 N_A_193_241#_c_526_p N_A1_M1025_g 6.1326e-19 $X=7.425 $Y=0.495 $X2=0
+ $Y2=0
cc_369 N_A_193_241#_c_451_n N_A1_M1025_g 0.0142468f $X=8.19 $Y=0.34 $X2=0 $Y2=0
cc_370 N_A_193_241#_c_453_n N_A1_M1025_g 0.00991507f $X=8.44 $Y=1.95 $X2=0 $Y2=0
cc_371 N_A_193_241#_c_457_n N_A1_M1025_g 4.67633e-19 $X=8.357 $Y=1.03 $X2=0
+ $Y2=0
cc_372 N_A_193_241#_c_466_n N_A1_c_692_n 0.0651388f $X=8.195 $Y=2.075 $X2=0
+ $Y2=0
cc_373 N_A_193_241#_c_453_n N_A1_c_692_n 0.025097f $X=8.44 $Y=1.95 $X2=0 $Y2=0
cc_374 N_A_193_241#_c_466_n N_A1_c_693_n 0.00294117f $X=8.195 $Y=2.075 $X2=0
+ $Y2=0
cc_375 N_A_193_241#_c_453_n N_A1_c_693_n 0.00642921f $X=8.44 $Y=1.95 $X2=0 $Y2=0
cc_376 N_A_193_241#_M1000_g N_VPWR_c_737_n 0.0114012f $X=1.055 $Y=2.4 $X2=0
+ $Y2=0
cc_377 N_A_193_241#_M1004_g N_VPWR_c_737_n 0.001604f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_378 N_A_193_241#_M1004_g N_VPWR_c_738_n 0.00456895f $X=1.675 $Y=2.4 $X2=0
+ $Y2=0
cc_379 N_A_193_241#_M1019_g N_VPWR_c_738_n 0.00456895f $X=2.295 $Y=2.4 $X2=0
+ $Y2=0
cc_380 N_A_193_241#_M1020_g N_VPWR_c_739_n 0.00462601f $X=2.915 $Y=2.4 $X2=0
+ $Y2=0
cc_381 N_A_193_241#_M1000_g N_VPWR_c_742_n 0.00460063f $X=1.055 $Y=2.4 $X2=0
+ $Y2=0
cc_382 N_A_193_241#_M1004_g N_VPWR_c_742_n 0.0039528f $X=1.675 $Y=2.4 $X2=0
+ $Y2=0
cc_383 N_A_193_241#_M1019_g N_VPWR_c_748_n 0.0039528f $X=2.295 $Y=2.4 $X2=0
+ $Y2=0
cc_384 N_A_193_241#_M1020_g N_VPWR_c_748_n 0.0039528f $X=2.915 $Y=2.4 $X2=0
+ $Y2=0
cc_385 N_A_193_241#_c_468_n N_VPWR_c_749_n 0.0146357f $X=8.36 $Y=2.465 $X2=0
+ $Y2=0
cc_386 N_A_193_241#_M1000_g N_VPWR_c_736_n 0.00444732f $X=1.055 $Y=2.4 $X2=0
+ $Y2=0
cc_387 N_A_193_241#_M1004_g N_VPWR_c_736_n 0.00505754f $X=1.675 $Y=2.4 $X2=0
+ $Y2=0
cc_388 N_A_193_241#_M1019_g N_VPWR_c_736_n 0.00505754f $X=2.295 $Y=2.4 $X2=0
+ $Y2=0
cc_389 N_A_193_241#_M1020_g N_VPWR_c_736_n 0.00509401f $X=2.915 $Y=2.4 $X2=0
+ $Y2=0
cc_390 N_A_193_241#_c_468_n N_VPWR_c_736_n 0.0121141f $X=8.36 $Y=2.465 $X2=0
+ $Y2=0
cc_391 N_A_193_241#_M1000_g N_X_c_837_n 0.0193092f $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_392 N_A_193_241#_M1004_g N_X_c_837_n 0.0119463f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_393 N_A_193_241#_c_444_n N_X_c_837_n 0.00827407f $X=1.22 $Y=1.28 $X2=0 $Y2=0
cc_394 N_A_193_241#_M1006_g N_X_c_838_n 0.00662985f $X=1.22 $Y=0.76 $X2=0 $Y2=0
cc_395 N_A_193_241#_c_429_n N_X_c_838_n 0.00327521f $X=1.615 $Y=0.18 $X2=0 $Y2=0
cc_396 N_A_193_241#_c_431_n N_X_c_838_n 0.00379483f $X=1.675 $Y=1.295 $X2=0
+ $Y2=0
cc_397 N_A_193_241#_M1004_g N_X_c_838_n 0.00250774f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_398 N_A_193_241#_M1012_g N_X_c_838_n 0.0120726f $X=1.69 $Y=0.76 $X2=0 $Y2=0
cc_399 N_A_193_241#_M1021_g N_X_c_838_n 0.00149354f $X=2.28 $Y=0.76 $X2=0 $Y2=0
cc_400 N_A_193_241#_M1019_g N_X_c_839_n 0.0108f $X=2.295 $Y=2.4 $X2=0 $Y2=0
cc_401 N_A_193_241#_c_441_n N_X_c_839_n 0.00715706f $X=2.915 $Y=1.46 $X2=0 $Y2=0
cc_402 N_A_193_241#_M1020_g N_X_c_839_n 0.00525344f $X=2.915 $Y=2.4 $X2=0 $Y2=0
cc_403 N_A_193_241#_M1012_g N_X_c_840_n 0.00150338f $X=1.69 $Y=0.76 $X2=0 $Y2=0
cc_404 N_A_193_241#_M1021_g N_X_c_840_n 0.0125712f $X=2.28 $Y=0.76 $X2=0 $Y2=0
cc_405 N_A_193_241#_c_436_n N_X_c_840_n 0.00389807f $X=2.295 $Y=1.295 $X2=0
+ $Y2=0
cc_406 N_A_193_241#_M1019_g N_X_c_840_n 0.00255008f $X=2.295 $Y=2.4 $X2=0 $Y2=0
cc_407 N_A_193_241#_c_438_n N_X_c_840_n 0.00233944f $X=2.635 $Y=0.18 $X2=0 $Y2=0
cc_408 N_A_193_241#_M1023_g N_X_c_840_n 0.021545f $X=2.71 $Y=0.76 $X2=0 $Y2=0
cc_409 N_A_193_241#_c_441_n N_X_c_840_n 0.00253386f $X=2.915 $Y=1.46 $X2=0 $Y2=0
cc_410 N_A_193_241#_M1004_g N_X_c_841_n 0.0227963f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_411 N_A_193_241#_M1019_g N_X_c_841_n 0.0229567f $X=2.295 $Y=2.4 $X2=0 $Y2=0
cc_412 N_A_193_241#_c_466_n N_A_725_391#_M1011_d 0.00168223f $X=8.195 $Y=2.075
+ $X2=0 $Y2=0
cc_413 N_A_193_241#_M1011_s N_A_725_391#_c_896_n 0.00464935f $X=6.32 $Y=1.96
+ $X2=0 $Y2=0
cc_414 N_A_193_241#_c_466_n N_A_939_391#_M1005_d 0.00167813f $X=8.195 $Y=2.075
+ $X2=0 $Y2=0
cc_415 N_A_193_241#_c_448_n N_A_939_391#_c_941_n 0.0270752f $X=6.3 $Y=1.615
+ $X2=0 $Y2=0
cc_416 N_A_193_241#_c_458_n N_A_939_391#_c_941_n 0.0121277f $X=5.78 $Y=1.615
+ $X2=0 $Y2=0
cc_417 N_A_193_241#_M1011_s N_A_939_391#_c_942_n 0.00663104f $X=6.32 $Y=1.96
+ $X2=0 $Y2=0
cc_418 N_A_193_241#_M1016_s N_A_939_391#_c_942_n 0.00493062f $X=7.265 $Y=1.96
+ $X2=0 $Y2=0
cc_419 N_A_193_241#_c_448_n N_A_939_391#_c_942_n 0.00496304f $X=6.3 $Y=1.615
+ $X2=0 $Y2=0
cc_420 N_A_193_241#_c_449_n N_A_939_391#_c_942_n 0.00303812f $X=6.23 $Y=1.615
+ $X2=0 $Y2=0
cc_421 N_A_193_241#_c_466_n N_A_939_391#_c_942_n 0.067604f $X=8.195 $Y=2.075
+ $X2=0 $Y2=0
cc_422 N_A_193_241#_c_467_n N_A_939_391#_c_942_n 0.013893f $X=6.47 $Y=2.075
+ $X2=0 $Y2=0
cc_423 N_A_193_241#_c_448_n N_A_939_391#_c_944_n 0.00864147f $X=6.3 $Y=1.615
+ $X2=0 $Y2=0
cc_424 N_A_193_241#_c_449_n N_A_939_391#_c_944_n 0.00352482f $X=6.23 $Y=1.615
+ $X2=0 $Y2=0
cc_425 N_A_193_241#_c_467_n N_A_939_391#_c_944_n 0.00886829f $X=6.47 $Y=2.075
+ $X2=0 $Y2=0
cc_426 N_A_193_241#_c_466_n N_A_939_391#_c_945_n 0.0174907f $X=8.195 $Y=2.075
+ $X2=0 $Y2=0
cc_427 N_A_193_241#_c_468_n N_A_939_391#_c_945_n 0.0172628f $X=8.36 $Y=2.465
+ $X2=0 $Y2=0
cc_428 N_A_193_241#_c_430_n N_VGND_c_988_n 0.0155675f $X=1.295 $Y=0.18 $X2=0
+ $Y2=0
cc_429 N_A_193_241#_c_444_n N_VGND_c_988_n 0.00703432f $X=1.22 $Y=1.28 $X2=0
+ $Y2=0
cc_430 N_A_193_241#_M1012_g N_VGND_c_989_n 0.00786117f $X=1.69 $Y=0.76 $X2=0
+ $Y2=0
cc_431 N_A_193_241#_c_434_n N_VGND_c_989_n 0.0244461f $X=2.205 $Y=0.18 $X2=0
+ $Y2=0
cc_432 N_A_193_241#_M1021_g N_VGND_c_989_n 0.00999417f $X=2.28 $Y=0.76 $X2=0
+ $Y2=0
cc_433 N_A_193_241#_M1021_g N_VGND_c_990_n 0.00138461f $X=2.28 $Y=0.76 $X2=0
+ $Y2=0
cc_434 N_A_193_241#_M1023_g N_VGND_c_990_n 0.0100627f $X=2.71 $Y=0.76 $X2=0
+ $Y2=0
cc_435 N_A_193_241#_c_440_n N_VGND_c_990_n 0.0261591f $X=5.63 $Y=0.18 $X2=0
+ $Y2=0
cc_436 N_A_193_241#_c_441_n N_VGND_c_990_n 0.00409955f $X=2.915 $Y=1.46 $X2=0
+ $Y2=0
cc_437 N_A_193_241#_c_440_n N_VGND_c_991_n 0.0232603f $X=5.63 $Y=0.18 $X2=0
+ $Y2=0
cc_438 N_A_193_241#_c_440_n N_VGND_c_992_n 0.0334796f $X=5.63 $Y=0.18 $X2=0
+ $Y2=0
cc_439 N_A_193_241#_c_440_n N_VGND_c_993_n 0.0277529f $X=5.63 $Y=0.18 $X2=0
+ $Y2=0
cc_440 N_A_193_241#_c_443_n N_VGND_c_993_n 0.00432999f $X=5.705 $Y=1.45 $X2=0
+ $Y2=0
cc_441 N_A_193_241#_c_454_n N_VGND_c_993_n 0.021907f $X=6.425 $Y=0.515 $X2=0
+ $Y2=0
cc_442 N_A_193_241#_c_430_n N_VGND_c_996_n 0.0208701f $X=1.295 $Y=0.18 $X2=0
+ $Y2=0
cc_443 N_A_193_241#_c_434_n N_VGND_c_998_n 0.0241797f $X=2.205 $Y=0.18 $X2=0
+ $Y2=0
cc_444 N_A_193_241#_c_440_n N_VGND_c_999_n 0.0185474f $X=5.63 $Y=0.18 $X2=0
+ $Y2=0
cc_445 N_A_193_241#_c_440_n N_VGND_c_1000_n 0.00710974f $X=5.63 $Y=0.18 $X2=0
+ $Y2=0
cc_446 N_A_193_241#_c_451_n N_VGND_c_1000_n 0.0618101f $X=8.19 $Y=0.34 $X2=0
+ $Y2=0
cc_447 N_A_193_241#_c_454_n N_VGND_c_1000_n 0.0933251f $X=6.425 $Y=0.515 $X2=0
+ $Y2=0
cc_448 N_A_193_241#_c_456_n N_VGND_c_1000_n 0.0235818f $X=7.425 $Y=0.34 $X2=0
+ $Y2=0
cc_449 N_A_193_241#_c_429_n N_VGND_c_1001_n 0.00836613f $X=1.615 $Y=0.18 $X2=0
+ $Y2=0
cc_450 N_A_193_241#_c_430_n N_VGND_c_1001_n 0.0114564f $X=1.295 $Y=0.18 $X2=0
+ $Y2=0
cc_451 N_A_193_241#_c_434_n N_VGND_c_1001_n 0.00646961f $X=2.205 $Y=0.18 $X2=0
+ $Y2=0
cc_452 N_A_193_241#_c_438_n N_VGND_c_1001_n 0.00686833f $X=2.635 $Y=0.18 $X2=0
+ $Y2=0
cc_453 N_A_193_241#_c_440_n N_VGND_c_1001_n 0.0624474f $X=5.63 $Y=0.18 $X2=0
+ $Y2=0
cc_454 N_A_193_241#_c_445_n N_VGND_c_1001_n 0.00824287f $X=1.69 $Y=0.18 $X2=0
+ $Y2=0
cc_455 N_A_193_241#_c_446_n N_VGND_c_1001_n 0.00829753f $X=2.28 $Y=0.18 $X2=0
+ $Y2=0
cc_456 N_A_193_241#_c_447_n N_VGND_c_1001_n 0.00491962f $X=2.71 $Y=0.18 $X2=0
+ $Y2=0
cc_457 N_A_193_241#_c_451_n N_VGND_c_1001_n 0.0343238f $X=8.19 $Y=0.34 $X2=0
+ $Y2=0
cc_458 N_A_193_241#_c_454_n N_VGND_c_1001_n 0.052653f $X=6.425 $Y=0.515 $X2=0
+ $Y2=0
cc_459 N_A_193_241#_c_456_n N_VGND_c_1001_n 0.0127177f $X=7.425 $Y=0.34 $X2=0
+ $Y2=0
cc_460 N_A_193_241#_c_451_n N_A_709_119#_M1014_s 0.00208352f $X=8.19 $Y=0.34
+ $X2=0 $Y2=0
cc_461 N_A_193_241#_c_440_n N_A_709_119#_c_1094_n 0.00622628f $X=5.63 $Y=0.18
+ $X2=0 $Y2=0
cc_462 N_A_193_241#_c_443_n N_A_709_119#_c_1096_n 0.0135146f $X=5.705 $Y=1.45
+ $X2=0 $Y2=0
cc_463 N_A_193_241#_c_448_n N_A_709_119#_c_1096_n 0.0820582f $X=6.3 $Y=1.615
+ $X2=0 $Y2=0
cc_464 N_A_193_241#_c_449_n N_A_709_119#_c_1096_n 0.0123082f $X=6.23 $Y=1.615
+ $X2=0 $Y2=0
cc_465 N_A_193_241#_c_466_n N_A_709_119#_c_1096_n 0.0111911f $X=8.195 $Y=2.075
+ $X2=0 $Y2=0
cc_466 N_A_193_241#_c_526_p N_A_709_119#_c_1096_n 0.0229858f $X=7.425 $Y=0.495
+ $X2=0 $Y2=0
cc_467 N_A_193_241#_c_453_n N_A_709_119#_c_1096_n 0.00893256f $X=8.44 $Y=1.95
+ $X2=0 $Y2=0
cc_468 N_A_193_241#_c_458_n N_A_709_119#_c_1096_n 0.00549303f $X=5.78 $Y=1.615
+ $X2=0 $Y2=0
cc_469 N_A_193_241#_c_451_n N_A_709_119#_c_1097_n 0.0149266f $X=8.19 $Y=0.34
+ $X2=0 $Y2=0
cc_470 N_A_193_241#_c_453_n N_A_709_119#_c_1097_n 0.00142601f $X=8.44 $Y=1.95
+ $X2=0 $Y2=0
cc_471 N_A_193_241#_c_457_n N_A_709_119#_c_1097_n 0.00155021f $X=8.357 $Y=1.03
+ $X2=0 $Y2=0
cc_472 N_A_193_241#_c_443_n N_A_709_119#_c_1099_n 3.54931e-19 $X=5.705 $Y=1.45
+ $X2=0 $Y2=0
cc_473 N_A_193_241#_c_450_n N_A_937_119#_M1017_d 0.00197722f $X=7.26 $Y=0.34
+ $X2=0 $Y2=0
cc_474 N_A_193_241#_M1017_s N_A_937_119#_c_1154_n 0.019235f $X=5.855 $Y=0.37
+ $X2=0 $Y2=0
cc_475 N_A_193_241#_c_443_n N_A_937_119#_c_1154_n 0.009911f $X=5.705 $Y=1.45
+ $X2=0 $Y2=0
cc_476 N_A_193_241#_c_450_n N_A_937_119#_c_1154_n 0.00418581f $X=7.26 $Y=0.34
+ $X2=0 $Y2=0
cc_477 N_A_193_241#_c_454_n N_A_937_119#_c_1154_n 0.0552517f $X=6.425 $Y=0.515
+ $X2=0 $Y2=0
cc_478 N_A_193_241#_c_440_n N_A_937_119#_c_1155_n 0.00557458f $X=5.63 $Y=0.18
+ $X2=0 $Y2=0
cc_479 N_A_193_241#_c_443_n N_A_937_119#_c_1155_n 8.19579e-19 $X=5.705 $Y=1.45
+ $X2=0 $Y2=0
cc_480 N_A_193_241#_c_440_n N_A_937_119#_c_1160_n 0.00156495f $X=5.63 $Y=0.18
+ $X2=0 $Y2=0
cc_481 N_A_193_241#_c_443_n N_A_937_119#_c_1156_n 0.0057997f $X=5.705 $Y=1.45
+ $X2=0 $Y2=0
cc_482 N_A_193_241#_c_450_n N_A_937_119#_c_1171_n 0.0152769f $X=7.26 $Y=0.34
+ $X2=0 $Y2=0
cc_483 N_A0_M1016_g N_A1_M1005_g 0.0452083f $X=7.175 $Y=2.46 $X2=0 $Y2=0
cc_484 N_A0_M1022_g N_A1_M1014_g 0.022348f $X=7.16 $Y=0.69 $X2=0 $Y2=0
cc_485 A0 N_A1_c_692_n 0.0211953f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_486 N_A0_c_648_n N_A1_c_692_n 0.0034029f $X=7.16 $Y=1.615 $X2=0 $Y2=0
cc_487 A0 N_A1_c_693_n 2.45568e-19 $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_488 N_A0_c_648_n N_A1_c_693_n 0.0168961f $X=7.16 $Y=1.615 $X2=0 $Y2=0
cc_489 N_A0_M1011_g N_VPWR_c_749_n 0.00349978f $X=6.725 $Y=2.46 $X2=0 $Y2=0
cc_490 N_A0_M1016_g N_VPWR_c_749_n 0.00519794f $X=7.175 $Y=2.46 $X2=0 $Y2=0
cc_491 N_A0_M1011_g N_VPWR_c_736_n 0.00434652f $X=6.725 $Y=2.46 $X2=0 $Y2=0
cc_492 N_A0_M1016_g N_VPWR_c_736_n 0.00522701f $X=7.175 $Y=2.46 $X2=0 $Y2=0
cc_493 N_A0_M1011_g N_A_725_391#_c_896_n 0.015498f $X=6.725 $Y=2.46 $X2=0 $Y2=0
cc_494 N_A0_M1016_g N_A_725_391#_c_896_n 0.00611637f $X=7.175 $Y=2.46 $X2=0
+ $Y2=0
cc_495 N_A0_M1011_g N_A_939_391#_c_942_n 0.0135003f $X=6.725 $Y=2.46 $X2=0 $Y2=0
cc_496 N_A0_M1016_g N_A_939_391#_c_942_n 0.0129227f $X=7.175 $Y=2.46 $X2=0 $Y2=0
cc_497 N_A0_M1011_g N_A_939_391#_c_944_n 0.00323126f $X=6.725 $Y=2.46 $X2=0
+ $Y2=0
cc_498 N_A0_M1016_g N_A_939_391#_c_945_n 0.00160299f $X=7.175 $Y=2.46 $X2=0
+ $Y2=0
cc_499 N_A0_M1017_g N_VGND_c_1000_n 0.00278271f $X=6.71 $Y=0.69 $X2=0 $Y2=0
cc_500 N_A0_M1022_g N_VGND_c_1000_n 0.00278271f $X=7.16 $Y=0.69 $X2=0 $Y2=0
cc_501 N_A0_M1017_g N_VGND_c_1001_n 0.00357715f $X=6.71 $Y=0.69 $X2=0 $Y2=0
cc_502 N_A0_M1022_g N_VGND_c_1001_n 0.00350534f $X=7.16 $Y=0.69 $X2=0 $Y2=0
cc_503 N_A0_M1017_g N_A_709_119#_c_1096_n 0.0127144f $X=6.71 $Y=0.69 $X2=0 $Y2=0
cc_504 N_A0_M1022_g N_A_709_119#_c_1096_n 0.0175267f $X=7.16 $Y=0.69 $X2=0 $Y2=0
cc_505 A0 N_A_709_119#_c_1096_n 0.032153f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_506 N_A0_c_648_n N_A_709_119#_c_1096_n 0.00359019f $X=7.16 $Y=1.615 $X2=0
+ $Y2=0
cc_507 N_A0_M1017_g N_A_937_119#_c_1154_n 0.0112042f $X=6.71 $Y=0.69 $X2=0 $Y2=0
cc_508 N_A0_M1017_g N_A_937_119#_c_1171_n 0.00916617f $X=6.71 $Y=0.69 $X2=0
+ $Y2=0
cc_509 N_A0_M1022_g N_A_937_119#_c_1171_n 0.0030388f $X=7.16 $Y=0.69 $X2=0 $Y2=0
cc_510 N_A1_M1005_g N_VPWR_c_749_n 0.005209f $X=7.635 $Y=2.46 $X2=0 $Y2=0
cc_511 N_A1_M1008_g N_VPWR_c_749_n 0.005209f $X=8.085 $Y=2.46 $X2=0 $Y2=0
cc_512 N_A1_M1005_g N_VPWR_c_736_n 0.00521734f $X=7.635 $Y=2.46 $X2=0 $Y2=0
cc_513 N_A1_M1008_g N_VPWR_c_736_n 0.00987267f $X=8.085 $Y=2.46 $X2=0 $Y2=0
cc_514 N_A1_M1005_g N_A_725_391#_c_896_n 7.86993e-19 $X=7.635 $Y=2.46 $X2=0
+ $Y2=0
cc_515 N_A1_M1005_g N_A_939_391#_c_942_n 0.00963291f $X=7.635 $Y=2.46 $X2=0
+ $Y2=0
cc_516 N_A1_M1005_g N_A_939_391#_c_945_n 0.00983358f $X=7.635 $Y=2.46 $X2=0
+ $Y2=0
cc_517 N_A1_M1008_g N_A_939_391#_c_945_n 0.00807054f $X=8.085 $Y=2.46 $X2=0
+ $Y2=0
cc_518 N_A1_M1014_g N_VGND_c_1000_n 0.00278247f $X=7.64 $Y=0.69 $X2=0 $Y2=0
cc_519 N_A1_M1025_g N_VGND_c_1000_n 0.00278271f $X=8.1 $Y=0.69 $X2=0 $Y2=0
cc_520 N_A1_M1014_g N_VGND_c_1001_n 0.00354264f $X=7.64 $Y=0.69 $X2=0 $Y2=0
cc_521 N_A1_M1025_g N_VGND_c_1001_n 0.00357524f $X=8.1 $Y=0.69 $X2=0 $Y2=0
cc_522 N_A1_M1014_g N_A_709_119#_c_1096_n 0.0144407f $X=7.64 $Y=0.69 $X2=0 $Y2=0
cc_523 N_A1_M1025_g N_A_709_119#_c_1096_n 0.00220281f $X=8.1 $Y=0.69 $X2=0 $Y2=0
cc_524 N_A1_c_692_n N_A_709_119#_c_1096_n 0.054688f $X=8.01 $Y=1.615 $X2=0 $Y2=0
cc_525 N_A1_c_693_n N_A_709_119#_c_1096_n 0.00460576f $X=8.1 $Y=1.615 $X2=0
+ $Y2=0
cc_526 N_A1_M1014_g N_A_709_119#_c_1097_n 0.00268042f $X=7.64 $Y=0.69 $X2=0
+ $Y2=0
cc_527 N_A1_M1025_g N_A_709_119#_c_1097_n 0.00201605f $X=8.1 $Y=0.69 $X2=0 $Y2=0
cc_528 N_VPWR_M1004_s N_X_c_841_n 0.00464694f $X=1.765 $Y=1.84 $X2=0 $Y2=0
cc_529 N_VPWR_M1013_s N_A_725_391#_c_895_n 0.0106235f $X=4.075 $Y=1.955 $X2=0
+ $Y2=0
cc_530 N_VPWR_M1018_s N_A_725_391#_c_895_n 0.00861488f $X=5.145 $Y=1.955 $X2=0
+ $Y2=0
cc_531 N_VPWR_c_740_n N_A_725_391#_c_895_n 0.025501f $X=4.295 $Y=2.94 $X2=0
+ $Y2=0
cc_532 N_VPWR_c_741_n N_A_725_391#_c_895_n 0.0193213f $X=5.365 $Y=2.94 $X2=0
+ $Y2=0
cc_533 N_VPWR_c_744_n N_A_725_391#_c_895_n 0.00241745f $X=4.13 $Y=3.33 $X2=0
+ $Y2=0
cc_534 N_VPWR_c_746_n N_A_725_391#_c_895_n 0.00878572f $X=5.2 $Y=3.33 $X2=0
+ $Y2=0
cc_535 N_VPWR_c_749_n N_A_725_391#_c_895_n 0.00253166f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_536 N_VPWR_c_736_n N_A_725_391#_c_895_n 0.0295184f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_537 N_VPWR_c_749_n N_A_725_391#_c_896_n 0.0545953f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_538 N_VPWR_c_736_n N_A_725_391#_c_896_n 0.0464727f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_539 N_VPWR_c_739_n N_A_725_391#_c_897_n 0.00107993f $X=3.225 $Y=3 $X2=0 $Y2=0
cc_540 N_VPWR_c_740_n N_A_725_391#_c_897_n 0.00688434f $X=4.295 $Y=2.94 $X2=0
+ $Y2=0
cc_541 N_VPWR_c_744_n N_A_725_391#_c_897_n 0.010785f $X=4.13 $Y=3.33 $X2=0 $Y2=0
cc_542 N_VPWR_c_736_n N_A_725_391#_c_897_n 0.00900085f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_543 N_VPWR_c_741_n N_A_725_391#_c_898_n 0.0156058f $X=5.365 $Y=2.94 $X2=0
+ $Y2=0
cc_544 N_VPWR_c_749_n N_A_725_391#_c_898_n 0.00737699f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_545 N_VPWR_c_736_n N_A_725_391#_c_898_n 0.0061588f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_546 N_VPWR_M1018_s N_A_939_391#_c_941_n 0.0134142f $X=5.145 $Y=1.955 $X2=0
+ $Y2=0
cc_547 N_VPWR_c_736_n N_A_939_391#_c_942_n 0.0201929f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_548 N_VPWR_c_749_n N_A_939_391#_c_945_n 0.0143496f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_549 N_VPWR_c_736_n N_A_939_391#_c_945_n 0.01179f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_550 N_X_c_837_n N_VGND_c_988_n 0.00100635f $X=1.475 $Y=1.37 $X2=0 $Y2=0
cc_551 N_X_c_838_n N_VGND_c_988_n 0.00272557f $X=1.475 $Y=0.535 $X2=0 $Y2=0
cc_552 N_X_c_838_n N_VGND_c_989_n 0.0270562f $X=1.475 $Y=0.535 $X2=0 $Y2=0
cc_553 N_X_c_840_n N_VGND_c_989_n 0.0508519f $X=2.495 $Y=0.535 $X2=0 $Y2=0
cc_554 N_X_c_841_n N_VGND_c_989_n 0.0192123f $X=2.33 $Y=1.625 $X2=0 $Y2=0
cc_555 N_X_c_840_n N_VGND_c_990_n 0.0702289f $X=2.495 $Y=0.535 $X2=0 $Y2=0
cc_556 N_X_c_838_n N_VGND_c_996_n 0.0134715f $X=1.475 $Y=0.535 $X2=0 $Y2=0
cc_557 N_X_c_840_n N_VGND_c_998_n 0.017052f $X=2.495 $Y=0.535 $X2=0 $Y2=0
cc_558 N_X_c_838_n N_VGND_c_1001_n 0.0106052f $X=1.475 $Y=0.535 $X2=0 $Y2=0
cc_559 N_X_c_840_n N_VGND_c_1001_n 0.0135629f $X=2.495 $Y=0.535 $X2=0 $Y2=0
cc_560 N_A_725_391#_c_895_n N_A_939_391#_M1015_d 0.00458554f $X=5.62 $Y=2.52
+ $X2=-0.19 $Y2=1.66
cc_561 N_A_725_391#_c_896_n N_A_939_391#_c_941_n 0.00682381f $X=6.95 $Y=2.805
+ $X2=0 $Y2=0
cc_562 N_A_725_391#_c_898_n N_A_939_391#_c_941_n 0.0139328f $X=5.705 $Y=2.52
+ $X2=0 $Y2=0
cc_563 N_A_725_391#_M1011_d N_A_939_391#_c_942_n 0.00321075f $X=6.815 $Y=1.96
+ $X2=0 $Y2=0
cc_564 N_A_725_391#_c_896_n N_A_939_391#_c_942_n 0.0589027f $X=6.95 $Y=2.805
+ $X2=0 $Y2=0
cc_565 N_A_725_391#_c_895_n N_A_939_391#_c_943_n 0.0574455f $X=5.62 $Y=2.52
+ $X2=0 $Y2=0
cc_566 N_A_725_391#_c_896_n N_A_939_391#_c_944_n 0.0137316f $X=6.95 $Y=2.805
+ $X2=0 $Y2=0
cc_567 N_A_725_391#_c_898_n N_A_939_391#_c_944_n 0.0079066f $X=5.705 $Y=2.52
+ $X2=0 $Y2=0
cc_568 N_A_725_391#_c_896_n N_A_939_391#_c_945_n 0.00774758f $X=6.95 $Y=2.805
+ $X2=0 $Y2=0
cc_569 N_A_939_391#_c_943_n N_A_709_119#_c_1098_n 0.00360319f $X=5.14 $Y=2.1
+ $X2=0 $Y2=0
cc_570 N_VGND_c_990_n N_A_709_119#_c_1094_n 0.0287269f $X=3.09 $Y=0.535 $X2=0
+ $Y2=0
cc_571 N_VGND_c_991_n N_A_709_119#_c_1094_n 0.0075028f $X=4.02 $Y=0 $X2=0 $Y2=0
cc_572 N_VGND_c_992_n N_A_709_119#_c_1094_n 0.0138611f $X=4.255 $Y=0.74 $X2=0
+ $Y2=0
cc_573 N_VGND_c_1001_n N_A_709_119#_c_1094_n 0.00907938f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_574 N_VGND_c_990_n N_A_709_119#_c_1095_n 0.00939066f $X=3.09 $Y=0.535 $X2=0
+ $Y2=0
cc_575 N_VGND_M1007_s N_A_709_119#_c_1096_n 0.00335654f $X=5.115 $Y=0.595 $X2=0
+ $Y2=0
cc_576 N_VGND_M1024_s N_A_709_119#_c_1098_n 0.00519037f $X=4.045 $Y=0.595 $X2=0
+ $Y2=0
cc_577 N_VGND_c_992_n N_A_709_119#_c_1098_n 0.0298247f $X=4.255 $Y=0.74 $X2=0
+ $Y2=0
cc_578 N_VGND_M1007_s N_A_709_119#_c_1099_n 0.00207907f $X=5.115 $Y=0.595 $X2=0
+ $Y2=0
cc_579 N_VGND_c_1001_n N_A_937_119#_c_1154_n 0.00702266f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_580 N_VGND_c_992_n N_A_937_119#_c_1155_n 0.0132163f $X=4.255 $Y=0.74 $X2=0
+ $Y2=0
cc_581 N_VGND_c_993_n N_A_937_119#_c_1155_n 7.70571e-19 $X=5.37 $Y=0.5 $X2=0
+ $Y2=0
cc_582 N_VGND_c_999_n N_A_937_119#_c_1155_n 0.0070895f $X=5.17 $Y=0 $X2=0 $Y2=0
cc_583 N_VGND_c_1001_n N_A_937_119#_c_1155_n 0.00875466f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_584 N_VGND_M1007_s N_A_937_119#_c_1160_n 0.00778741f $X=5.115 $Y=0.595 $X2=0
+ $Y2=0
cc_585 N_VGND_c_993_n N_A_937_119#_c_1160_n 0.0318174f $X=5.37 $Y=0.5 $X2=0
+ $Y2=0
cc_586 N_VGND_c_999_n N_A_937_119#_c_1160_n 0.00195503f $X=5.17 $Y=0 $X2=0 $Y2=0
cc_587 N_VGND_c_1001_n N_A_937_119#_c_1160_n 0.005356f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_588 N_VGND_M1007_s N_A_937_119#_c_1156_n 0.00137378f $X=5.115 $Y=0.595 $X2=0
+ $Y2=0
cc_589 N_VGND_c_1000_n N_A_937_119#_c_1156_n 0.00122935f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_590 N_VGND_c_1001_n N_A_937_119#_c_1156_n 0.00198148f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_591 N_A_709_119#_c_1098_n N_A_937_119#_M1003_d 0.00176461f $X=5.155 $Y=1.187
+ $X2=-0.19 $Y2=-0.245
cc_592 N_A_709_119#_c_1098_n N_A_937_119#_c_1155_n 0.0161925f $X=5.155 $Y=1.187
+ $X2=0 $Y2=0
cc_593 N_A_709_119#_c_1096_n N_A_937_119#_c_1160_n 0.0115278f $X=7.77 $Y=1.195
+ $X2=0 $Y2=0
cc_594 N_A_709_119#_c_1098_n N_A_937_119#_c_1160_n 0.0196564f $X=5.155 $Y=1.187
+ $X2=0 $Y2=0
cc_595 N_A_709_119#_c_1096_n N_A_937_119#_c_1156_n 0.089963f $X=7.77 $Y=1.195
+ $X2=0 $Y2=0
cc_596 N_A_709_119#_c_1096_n N_A_937_119#_c_1171_n 0.0208323f $X=7.77 $Y=1.195
+ $X2=0 $Y2=0

* NGSPICE file created from sky130_fd_sc_ms__o41a_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 VPWR a_83_270# X VPB pshort w=1.12e+06u l=180000u
+  ad=1.3554e+12p pd=7.11e+06u as=3.136e+11p ps=2.8e+06u
M1001 VGND A4 a_326_74# VNB nlowvt w=640000u l=150000u
+  ad=8.899e+11p pd=6.71e+06u as=6.24e+11p ps=5.79e+06u
M1002 a_83_270# B1 VPWR VPB pshort w=840000u l=180000u
+  ad=3.7225e+11p pd=2.95e+06u as=0p ps=0u
M1003 a_446_368# A4 a_83_270# VPB pshort w=1.12e+06u l=180000u
+  ad=2.688e+11p pd=2.72e+06u as=0p ps=0u
M1004 a_326_74# B1 a_83_270# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1005 a_644_368# A2 a_530_368# VPB pshort w=1.12e+06u l=180000u
+  ad=4.368e+11p pd=3.02e+06u as=4.368e+11p ps=3.02e+06u
M1006 VGND A2 a_326_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_530_368# A3 a_446_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_326_74# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_644_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_83_270# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1011 a_326_74# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_ms__nor2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__nor2b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.028400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.790000 1.010000 3.975000 1.180000 ;
        RECT 0.790000 1.180000 1.795000 1.340000 ;
        RECT 1.085000 1.340000 1.795000 1.410000 ;
        RECT 3.645000 1.180000 3.975000 1.550000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.413400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.750000 1.180000 5.155000 1.825000 ;
    END
  END B_N
  PIN Y
    ANTENNADIFFAREA  1.019200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.670000 3.810000 0.840000 ;
        RECT 0.125000 0.840000 0.355000 1.410000 ;
        RECT 0.185000 1.410000 0.355000 1.510000 ;
        RECT 0.185000 1.510000 0.705000 1.580000 ;
        RECT 0.185000 1.580000 2.055000 1.680000 ;
        RECT 0.535000 1.680000 2.055000 1.750000 ;
        RECT 1.885000 1.750000 2.055000 1.850000 ;
        RECT 1.885000 1.850000 2.165000 2.060000 ;
        RECT 1.885000 2.060000 3.145000 2.230000 ;
        RECT 1.885000 2.230000 2.165000 2.735000 ;
        RECT 2.060000 0.530000 2.390000 0.670000 ;
        RECT 2.895000 2.230000 3.145000 2.735000 ;
        RECT 3.560000 0.510000 3.810000 0.670000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 5.280000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.660000 5.470000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.115000  1.850000 0.365000 3.245000 ;
      RECT 0.565000  1.920000 1.715000 2.090000 ;
      RECT 0.565000  2.090000 0.895000 2.980000 ;
      RECT 1.095000  2.260000 1.265000 3.245000 ;
      RECT 1.465000  2.090000 1.715000 2.905000 ;
      RECT 1.465000  2.905000 3.645000 3.075000 ;
      RECT 1.550000  0.085000 1.880000 0.500000 ;
      RECT 2.225000  1.350000 3.225000 1.680000 ;
      RECT 2.365000  2.400000 2.695000 2.905000 ;
      RECT 2.570000  0.085000 3.380000 0.500000 ;
      RECT 3.055000  1.680000 3.225000 1.720000 ;
      RECT 3.055000  1.720000 4.580000 1.890000 ;
      RECT 3.315000  2.060000 3.645000 2.905000 ;
      RECT 3.815000  2.060000 4.145000 3.245000 ;
      RECT 3.990000  0.085000 4.240000 0.840000 ;
      RECT 4.350000  1.890000 4.580000 1.995000 ;
      RECT 4.350000  1.995000 4.680000 2.875000 ;
      RECT 4.410000  0.345000 5.165000 1.010000 ;
      RECT 4.410000  1.010000 4.580000 1.720000 ;
      RECT 4.880000  1.995000 5.130000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_ms__nor2b_4
END LIBRARY

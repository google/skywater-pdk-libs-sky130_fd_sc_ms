* File: sky130_fd_sc_ms__a311oi_2.pex.spice
* Created: Wed Sep  2 11:54:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A311OI_2%A3 3 5 7 8 10 13 15 22
r41 22 23 2.12647 $w=3.4e-07 $l=1.5e-08 $layer=POLY_cond $X=0.995 $Y=1.43
+ $X2=1.01 $Y2=1.43
r42 20 22 51.0353 $w=3.4e-07 $l=3.6e-07 $layer=POLY_cond $X=0.635 $Y=1.43
+ $X2=0.995 $Y2=1.43
r43 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.635
+ $Y=1.385 $X2=0.635 $Y2=1.385
r44 18 20 9.92353 $w=3.4e-07 $l=7e-08 $layer=POLY_cond $X=0.565 $Y=1.43
+ $X2=0.635 $Y2=1.43
r45 15 21 3.13714 $w=3.5e-07 $l=9e-08 $layer=LI1_cond $X=0.652 $Y=1.295
+ $X2=0.652 $Y2=1.385
r46 11 23 17.6285 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=1.01 $Y=1.64
+ $X2=1.01 $Y2=1.43
r47 11 13 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=1.01 $Y=1.64
+ $X2=1.01 $Y2=2.4
r48 8 22 21.9347 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.995 $Y=1.22
+ $X2=0.995 $Y2=1.43
r49 8 10 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.995 $Y=1.22
+ $X2=0.995 $Y2=0.74
r50 5 18 21.9347 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.565 $Y=1.22
+ $X2=0.565 $Y2=1.43
r51 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.565 $Y=1.22 $X2=0.565
+ $Y2=0.74
r52 1 18 0.708824 $w=3.4e-07 $l=5e-09 $layer=POLY_cond $X=0.56 $Y=1.43 $X2=0.565
+ $Y2=1.43
r53 1 3 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.56 $Y=1.55 $X2=0.56
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_2%A2 1 3 6 8 10 13 20 23 29 34
c56 29 0 9.06755e-20 $X=1.91 $Y=1.385
c57 1 0 1.90514e-19 $X=1.425 $Y=1.22
r58 28 29 8.15692 $w=3.25e-07 $l=5.5e-08 $layer=POLY_cond $X=1.855 $Y=1.385
+ $X2=1.91 $Y2=1.385
r59 25 26 5.19077 $w=3.25e-07 $l=3.5e-08 $layer=POLY_cond $X=1.425 $Y=1.385
+ $X2=1.46 $Y2=1.385
r60 23 34 3.7435 $w=3.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.365
+ $X2=1.315 $Y2=1.365
r61 21 29 2.22462 $w=3.25e-07 $l=1.5e-08 $layer=POLY_cond $X=1.925 $Y=1.385
+ $X2=1.91 $Y2=1.385
r62 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.925
+ $Y=1.385 $X2=1.925 $Y2=1.385
r63 18 28 47.4585 $w=3.25e-07 $l=3.2e-07 $layer=POLY_cond $X=1.535 $Y=1.385
+ $X2=1.855 $Y2=1.385
r64 18 26 11.1231 $w=3.25e-07 $l=7.5e-08 $layer=POLY_cond $X=1.535 $Y=1.385
+ $X2=1.46 $Y2=1.385
r65 17 20 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=1.535 $Y=1.385
+ $X2=1.925 $Y2=1.385
r66 17 34 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.535 $Y=1.385
+ $X2=1.315 $Y2=1.385
r67 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.535
+ $Y=1.385 $X2=1.535 $Y2=1.385
r68 11 29 16.5763 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.91 $Y=1.55
+ $X2=1.91 $Y2=1.385
r69 11 13 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.91 $Y=1.55
+ $X2=1.91 $Y2=2.4
r70 8 28 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.22
+ $X2=1.855 $Y2=1.385
r71 8 10 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.855 $Y=1.22
+ $X2=1.855 $Y2=0.74
r72 4 26 16.5763 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.46 $Y=1.55
+ $X2=1.46 $Y2=1.385
r73 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.46 $Y=1.55 $X2=1.46
+ $Y2=2.4
r74 1 25 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.22
+ $X2=1.425 $Y2=1.385
r75 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.425 $Y=1.22 $X2=1.425
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_2%A1 3 7 11 15 17 22 29
r54 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.035
+ $Y=1.515 $X2=3.035 $Y2=1.515
r55 27 29 14.9226 $w=3.23e-07 $l=1e-07 $layer=POLY_cond $X=2.935 $Y=1.49
+ $X2=3.035 $Y2=1.49
r56 26 27 14.1765 $w=3.23e-07 $l=9.5e-08 $layer=POLY_cond $X=2.84 $Y=1.49
+ $X2=2.935 $Y2=1.49
r57 22 30 4.73607 $w=3.63e-07 $l=1.5e-07 $layer=LI1_cond $X=3.052 $Y=1.665
+ $X2=3.052 $Y2=1.515
r58 20 26 55.9598 $w=3.23e-07 $l=3.75e-07 $layer=POLY_cond $X=2.465 $Y=1.49
+ $X2=2.84 $Y2=1.49
r59 20 24 11.192 $w=3.23e-07 $l=7.5e-08 $layer=POLY_cond $X=2.465 $Y=1.49
+ $X2=2.39 $Y2=1.49
r60 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.465
+ $Y=1.465 $X2=2.465 $Y2=1.465
r61 17 30 2.0523 $w=3.63e-07 $l=6.5e-08 $layer=LI1_cond $X=3.052 $Y=1.45
+ $X2=3.052 $Y2=1.515
r62 17 19 22.4591 $w=1.98e-07 $l=4.05e-07 $layer=LI1_cond $X=2.87 $Y=1.45
+ $X2=2.465 $Y2=1.45
r63 13 29 49.2446 $w=3.23e-07 $l=3.3e-07 $layer=POLY_cond $X=3.365 $Y=1.49
+ $X2=3.035 $Y2=1.49
r64 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.365 $Y=1.35
+ $X2=3.365 $Y2=0.74
r65 9 27 20.7134 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.935 $Y=1.3
+ $X2=2.935 $Y2=1.49
r66 9 11 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.935 $Y=1.3
+ $X2=2.935 $Y2=0.74
r67 5 26 16.4327 $w=1.8e-07 $l=1.9e-07 $layer=POLY_cond $X=2.84 $Y=1.68 $X2=2.84
+ $Y2=1.49
r68 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.84 $Y=1.68 $X2=2.84
+ $Y2=2.4
r69 1 24 16.4327 $w=1.8e-07 $l=1.9e-07 $layer=POLY_cond $X=2.39 $Y=1.68 $X2=2.39
+ $Y2=1.49
r70 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.39 $Y=1.68 $X2=2.39
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_2%B1 3 7 11 13 14 15 25
c49 25 0 1.60946e-19 $X=4.26 $Y=1.515
c50 15 0 7.19971e-20 $X=4.56 $Y=1.665
c51 3 0 1.0484e-19 $X=3.795 $Y=0.74
r52 23 25 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.185 $Y=1.515
+ $X2=4.26 $Y2=1.515
r53 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.185
+ $Y=1.515 $X2=4.185 $Y2=1.515
r54 21 23 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=3.81 $Y=1.515
+ $X2=4.185 $Y2=1.515
r55 19 21 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.795 $Y=1.515
+ $X2=3.81 $Y2=1.515
r56 15 24 10.0504 $w=4.28e-07 $l=3.75e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.185 $Y2=1.565
r57 14 24 2.81411 $w=4.28e-07 $l=1.05e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=4.185 $Y2=1.565
r58 13 14 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=4.08 $Y2=1.565
r59 9 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.26 $Y=1.68
+ $X2=4.26 $Y2=1.515
r60 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.26 $Y=1.68 $X2=4.26
+ $Y2=2.4
r61 5 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.81 $Y=1.68
+ $X2=3.81 $Y2=1.515
r62 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.81 $Y=1.68 $X2=3.81
+ $Y2=2.4
r63 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.795 $Y=1.35
+ $X2=3.795 $Y2=1.515
r64 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.795 $Y=1.35
+ $X2=3.795 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_2%C1 3 7 11 13 20 21
c39 20 0 1.60946e-19 $X=5.01 $Y=1.515
c40 11 0 7.19971e-20 $X=5.16 $Y=2.4
r41 19 21 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=5.01 $Y=1.515
+ $X2=5.16 $Y2=1.515
r42 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.01
+ $Y=1.515 $X2=5.01 $Y2=1.515
r43 17 19 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=4.71 $Y=1.515 $X2=5.01
+ $Y2=1.515
r44 15 17 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.635 $Y=1.515
+ $X2=4.71 $Y2=1.515
r45 13 20 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=5.01 $Y=1.665
+ $X2=5.01 $Y2=1.515
r46 9 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.16 $Y=1.68
+ $X2=5.16 $Y2=1.515
r47 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.16 $Y=1.68 $X2=5.16
+ $Y2=2.4
r48 5 17 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.71 $Y=1.68
+ $X2=4.71 $Y2=1.515
r49 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.71 $Y=1.68 $X2=4.71
+ $Y2=2.4
r50 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.635 $Y=1.35
+ $X2=4.635 $Y2=1.515
r51 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.635 $Y=1.35
+ $X2=4.635 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_2%VPWR 1 2 3 4 13 15 19 23 27 31 33 35 40 50
+ 51 57 60 63
r72 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r73 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r74 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r75 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r76 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r77 50 51 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r78 48 51 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r79 48 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r80 47 50 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r81 47 48 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r82 45 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.23 $Y=3.33
+ $X2=3.065 $Y2=3.33
r83 45 47 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.23 $Y=3.33 $X2=3.6
+ $Y2=3.33
r84 44 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r85 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r86 41 60 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.33 $Y=3.33 $X2=2.19
+ $Y2=3.33
r87 41 43 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.33 $Y=3.33
+ $X2=2.64 $Y2=3.33
r88 40 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.9 $Y=3.33
+ $X2=3.065 $Y2=3.33
r89 40 43 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.9 $Y=3.33 $X2=2.64
+ $Y2=3.33
r90 39 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r91 39 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r92 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r93 36 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.32 $Y=3.33
+ $X2=1.235 $Y2=3.33
r94 36 38 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.32 $Y=3.33
+ $X2=1.68 $Y2=3.33
r95 35 60 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.05 $Y=3.33 $X2=2.19
+ $Y2=3.33
r96 35 38 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.05 $Y=3.33 $X2=1.68
+ $Y2=3.33
r97 33 64 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r98 33 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r99 29 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=3.245
+ $X2=3.065 $Y2=3.33
r100 29 31 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=3.065 $Y=3.245
+ $X2=3.065 $Y2=2.405
r101 25 60 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=3.33
r102 25 27 41.9819 $w=2.78e-07 $l=1.02e-06 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=2.225
r103 21 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=3.245
+ $X2=1.235 $Y2=3.33
r104 21 23 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.235 $Y=3.245
+ $X2=1.235 $Y2=2.225
r105 20 54 3.94754 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=0.42 $Y=3.33
+ $X2=0.21 $Y2=3.33
r106 19 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=3.33
+ $X2=1.235 $Y2=3.33
r107 19 20 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.15 $Y=3.33
+ $X2=0.42 $Y2=3.33
r108 15 18 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.295 $Y=1.985
+ $X2=0.295 $Y2=2.815
r109 13 54 3.19563 $w=2.5e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.21 $Y2=3.33
r110 13 18 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.295 $Y2=2.815
r111 4 31 300 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=2 $X=2.93
+ $Y=1.84 $X2=3.065 $Y2=2.405
r112 3 27 300 $w=1.7e-07 $l=4.53845e-07 $layer=licon1_PDIFF $count=2 $X=2
+ $Y=1.84 $X2=2.15 $Y2=2.225
r113 2 23 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=1.1
+ $Y=1.84 $X2=1.235 $Y2=2.225
r114 1 18 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.21
+ $Y=1.84 $X2=0.335 $Y2=2.815
r115 1 15 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.21
+ $Y=1.84 $X2=0.335 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_2%A_130_368# 1 2 3 4 15 19 20 23 27 31 33 37
+ 38 43
c69 19 0 9.06755e-20 $X=1.52 $Y=1.805
r70 38 41 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.615 $Y=1.805
+ $X2=2.615 $Y2=1.985
r71 34 41 0.716491 $w=1.7e-07 $l=1.07121e-07 $layer=LI1_cond $X=2.7 $Y=2.035
+ $X2=2.615 $Y2=1.985
r72 33 43 3.65518 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=3.925 $Y=2.035
+ $X2=4.022 $Y2=2.035
r73 33 34 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=3.925 $Y=2.035
+ $X2=2.7 $Y2=2.035
r74 29 41 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.615 $Y=2.12
+ $X2=2.615 $Y2=1.985
r75 29 31 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.615 $Y=2.12
+ $X2=2.615 $Y2=2.4
r76 28 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.85 $Y=1.805
+ $X2=1.685 $Y2=1.805
r77 27 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=1.805
+ $X2=2.615 $Y2=1.805
r78 27 28 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.53 $Y=1.805
+ $X2=1.85 $Y2=1.805
r79 23 25 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.685 $Y=1.985
+ $X2=1.685 $Y2=2.815
r80 21 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.685 $Y=1.89
+ $X2=1.685 $Y2=1.805
r81 21 23 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.685 $Y=1.89
+ $X2=1.685 $Y2=1.985
r82 19 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=1.805
+ $X2=1.685 $Y2=1.805
r83 19 20 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.52 $Y=1.805
+ $X2=0.95 $Y2=1.805
r84 15 17 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.785 $Y=1.985
+ $X2=0.785 $Y2=2.815
r85 13 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.785 $Y=1.89
+ $X2=0.95 $Y2=1.805
r86 13 15 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.785 $Y=1.89
+ $X2=0.785 $Y2=1.985
r87 4 43 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=3.9
+ $Y=1.84 $X2=4.035 $Y2=2.115
r88 3 41 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.84 $X2=2.615 $Y2=1.985
r89 3 31 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=2.48
+ $Y=1.84 $X2=2.615 $Y2=2.4
r90 2 25 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.55
+ $Y=1.84 $X2=1.685 $Y2=2.815
r91 2 23 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.55
+ $Y=1.84 $X2=1.685 $Y2=1.985
r92 1 17 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.84 $X2=0.785 $Y2=2.815
r93 1 15 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.84 $X2=0.785 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_2%A_692_368# 1 2 3 12 14 15 18 22 26 28
r44 24 26 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.385 $Y=2.905
+ $X2=5.385 $Y2=2.425
r45 23 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.65 $Y=2.99
+ $X2=4.485 $Y2=2.99
r46 22 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.22 $Y=2.99
+ $X2=5.385 $Y2=2.905
r47 22 23 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.22 $Y=2.99
+ $X2=4.65 $Y2=2.99
r48 18 21 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=4.485 $Y=2.07
+ $X2=4.485 $Y2=2.815
r49 16 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.485 $Y=2.905
+ $X2=4.485 $Y2=2.99
r50 16 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.485 $Y=2.905
+ $X2=4.485 $Y2=2.815
r51 14 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=2.99
+ $X2=4.485 $Y2=2.99
r52 14 15 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=4.32 $Y=2.99
+ $X2=3.755 $Y2=2.99
r53 10 15 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=3.587 $Y=2.905
+ $X2=3.755 $Y2=2.99
r54 10 12 17.3726 $w=3.33e-07 $l=5.05e-07 $layer=LI1_cond $X=3.587 $Y=2.905
+ $X2=3.587 $Y2=2.4
r55 3 26 300 $w=1.7e-07 $l=6.48999e-07 $layer=licon1_PDIFF $count=2 $X=5.25
+ $Y=1.84 $X2=5.385 $Y2=2.425
r56 2 21 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.35
+ $Y=1.84 $X2=4.485 $Y2=2.815
r57 2 18 400 $w=1.7e-07 $l=2.89741e-07 $layer=licon1_PDIFF $count=1 $X=4.35
+ $Y=1.84 $X2=4.485 $Y2=2.07
r58 1 12 300 $w=1.7e-07 $l=6.19354e-07 $layer=licon1_PDIFF $count=2 $X=3.46
+ $Y=1.84 $X2=3.585 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_2%Y 1 2 3 4 13 19 25 28 30 32 34 35 47
r53 46 47 11.617 $w=8.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.85 $Y=0.765
+ $X2=4.685 $Y2=0.765
r54 34 35 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=5.52 $Y=1.295
+ $X2=5.52 $Y2=1.665
r55 34 40 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=5.52 $Y=1.295
+ $X2=5.52 $Y2=1.18
r56 32 40 8.46024 $w=2.3e-07 $l=4.15e-07 $layer=LI1_cond $X=5.52 $Y=0.765
+ $X2=5.52 $Y2=1.18
r57 32 46 9.65509 $w=8.28e-07 $l=6.7e-07 $layer=LI1_cond $X=5.52 $Y=0.765
+ $X2=4.85 $Y2=0.765
r58 31 35 14.2803 $w=2.28e-07 $l=2.85e-07 $layer=LI1_cond $X=5.52 $Y=1.95
+ $X2=5.52 $Y2=1.665
r59 26 30 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.02 $Y=2.035
+ $X2=4.935 $Y2=2.035
r60 25 31 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=5.405 $Y=2.035
+ $X2=5.52 $Y2=1.95
r61 25 26 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=5.405 $Y=2.035
+ $X2=5.02 $Y2=2.035
r62 22 28 5.16603 $w=2.5e-07 $l=1.60078e-07 $layer=LI1_cond $X=3.745 $Y=1.095
+ $X2=3.62 $Y2=1.015
r63 22 47 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.745 $Y=1.095
+ $X2=4.685 $Y2=1.095
r64 17 28 1.34256 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=3.62 $Y=0.85
+ $X2=3.62 $Y2=1.015
r65 17 19 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.62 $Y=0.85
+ $X2=3.62 $Y2=0.515
r66 13 28 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=3.495 $Y=1.015
+ $X2=3.62 $Y2=1.015
r67 13 15 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=3.495 $Y=1.015
+ $X2=2.72 $Y2=1.015
r68 4 30 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=4.8
+ $Y=1.84 $X2=4.935 $Y2=2.115
r69 3 46 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.71
+ $Y=0.37 $X2=4.85 $Y2=0.515
r70 2 28 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=3.44
+ $Y=0.37 $X2=3.58 $Y2=0.965
r71 2 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.44
+ $Y=0.37 $X2=3.58 $Y2=0.515
r72 1 15 182 $w=1.7e-07 $l=6.39453e-07 $layer=licon1_NDIFF $count=1 $X=2.595
+ $Y=0.37 $X2=2.72 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_2%A_45_74# 1 2 3 12 14 15 18 22 24 25
c35 24 0 1.90514e-19 $X=2.07 $Y=0.87
r36 24 25 7.05875 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=2.07 $Y=0.91
+ $X2=1.905 $Y2=0.91
r37 21 22 4.40882 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.295 $Y=0.89
+ $X2=1.21 $Y2=0.89
r38 21 25 29.2913 $w=2.38e-07 $l=6.1e-07 $layer=LI1_cond $X=1.295 $Y=0.89
+ $X2=1.905 $Y2=0.89
r39 16 22 2.0246 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.21 $Y=0.77 $X2=1.21
+ $Y2=0.89
r40 16 18 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.21 $Y=0.77
+ $X2=1.21 $Y2=0.495
r41 14 22 4.40882 $w=2.05e-07 $l=1.00995e-07 $layer=LI1_cond $X=1.125 $Y=0.925
+ $X2=1.21 $Y2=0.89
r42 14 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.125 $Y=0.925
+ $X2=0.435 $Y2=0.925
r43 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.31 $Y=0.84
+ $X2=0.435 $Y2=0.925
r44 10 12 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=0.31 $Y=0.84
+ $X2=0.31 $Y2=0.515
r45 3 24 182 $w=1.7e-07 $l=5.65685e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.37 $X2=2.07 $Y2=0.87
r46 2 18 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.21 $Y2=0.495
r47 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.225
+ $Y=0.37 $X2=0.35 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_2%VGND 1 2 9 13 15 17 22 35 36 39 42
r50 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r51 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r52 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r53 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r54 33 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r55 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r56 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r57 30 42 12.559 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=4.515 $Y=0 $X2=4.215
+ $Y2=0
r58 30 32 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.515 $Y=0 $X2=4.56
+ $Y2=0
r59 29 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r60 28 29 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r61 26 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r62 25 28 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r63 25 26 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r64 23 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r65 23 25 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r66 22 42 12.559 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=3.915 $Y=0 $X2=4.215
+ $Y2=0
r67 22 28 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.915 $Y=0 $X2=3.6
+ $Y2=0
r68 20 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r69 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r70 17 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r71 17 19 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r72 15 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.6
+ $Y2=0
r73 15 26 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=1.2
+ $Y2=0
r74 11 42 2.52064 $w=6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.215 $Y=0.085
+ $X2=4.215 $Y2=0
r75 11 13 11.7614 $w=5.98e-07 $l=5.9e-07 $layer=LI1_cond $X=4.215 $Y=0.085
+ $X2=4.215 $Y2=0.675
r76 7 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0
r77 7 9 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0.55
r78 2 13 91 $w=1.7e-07 $l=6.85748e-07 $layer=licon1_NDIFF $count=2 $X=3.87
+ $Y=0.37 $X2=4.42 $Y2=0.675
r79 1 9 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.64 $Y=0.37
+ $X2=0.78 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_2%A_300_74# 1 2 12 13
c18 12 0 1.0484e-19 $X=3.15 $Y=0.515
r19 12 13 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.15 $Y=0.515
+ $X2=2.985 $Y2=0.515
r20 9 13 62.0014 $w=2.48e-07 $l=1.345e-06 $layer=LI1_cond $X=1.64 $Y=0.475
+ $X2=2.985 $Y2=0.475
r21 2 12 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.01
+ $Y=0.37 $X2=3.15 $Y2=0.515
r22 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.64 $Y2=0.515
.ends


* NGSPICE file created from sky130_fd_sc_ms__a32o_4.ext - technology: sky130A

.subckt sky130_fd_sc_ms__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 a_587_110# B2 VGND VNB nlowvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=1.47252e+12p ps=1.141e+07u
M1001 a_83_283# B1 a_587_110# VNB nlowvt w=640000u l=150000u
+  ad=4.34975e+11p pd=4.13e+06u as=0p ps=0u
M1002 a_992_122# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=5.568e+11p pd=5.58e+06u as=0p ps=0u
M1003 X a_83_283# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=2.0706e+12p ps=1.665e+07u
M1004 X a_83_283# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_83_283# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_83_283# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_83_283# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.255e+11p pd=4.11e+06u as=0p ps=0u
M1008 X a_83_283# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_992_122# A2 a_1079_122# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.096e+11p ps=3.84e+06u
M1010 VPWR A2 a_509_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=1.955e+12p ps=1.591e+07u
M1011 a_509_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A3 a_992_122# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_509_392# A3 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_83_283# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_509_392# B2 a_83_283# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=6.4e+11p ps=5.28e+06u
M1016 a_509_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A3 a_509_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_509_392# B1 a_83_283# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_83_283# B1 a_509_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_83_283# B2 a_509_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_587_110# B1 a_83_283# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND B2 a_587_110# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND a_83_283# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1079_122# A2 a_992_122# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_83_283# A1 a_1079_122# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1079_122# A1 a_83_283# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR A1 a_509_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__and4_2.pxi.spice
* Created: Fri Aug 28 17:13:19 2020
* 
x_PM_SKY130_FD_SC_MS__AND4_2%A N_A_M1001_g N_A_M1005_g N_A_c_69_n N_A_c_70_n A
+ N_A_c_71_n PM_SKY130_FD_SC_MS__AND4_2%A
x_PM_SKY130_FD_SC_MS__AND4_2%B N_B_M1000_g N_B_M1003_g B B B N_B_c_98_n
+ N_B_c_99_n PM_SKY130_FD_SC_MS__AND4_2%B
x_PM_SKY130_FD_SC_MS__AND4_2%C N_C_M1011_g N_C_M1006_g C C C N_C_c_135_n
+ N_C_c_136_n PM_SKY130_FD_SC_MS__AND4_2%C
x_PM_SKY130_FD_SC_MS__AND4_2%D N_D_c_172_n N_D_M1007_g N_D_M1004_g N_D_c_168_n D
+ N_D_c_169_n N_D_c_170_n N_D_c_171_n PM_SKY130_FD_SC_MS__AND4_2%D
x_PM_SKY130_FD_SC_MS__AND4_2%A_56_74# N_A_56_74#_M1005_s N_A_56_74#_M1001_d
+ N_A_56_74#_M1006_d N_A_56_74#_M1002_g N_A_56_74#_M1009_g N_A_56_74#_M1008_g
+ N_A_56_74#_M1010_g N_A_56_74#_c_210_n N_A_56_74#_c_211_n N_A_56_74#_c_212_n
+ N_A_56_74#_c_219_n N_A_56_74#_c_220_n N_A_56_74#_c_244_n N_A_56_74#_c_221_n
+ N_A_56_74#_c_222_n N_A_56_74#_c_213_n N_A_56_74#_c_214_n N_A_56_74#_c_215_n
+ N_A_56_74#_c_224_n N_A_56_74#_c_255_n PM_SKY130_FD_SC_MS__AND4_2%A_56_74#
x_PM_SKY130_FD_SC_MS__AND4_2%VPWR N_VPWR_M1001_s N_VPWR_M1003_d N_VPWR_M1007_d
+ N_VPWR_M1010_s N_VPWR_c_317_n N_VPWR_c_318_n N_VPWR_c_319_n N_VPWR_c_320_n
+ N_VPWR_c_321_n N_VPWR_c_322_n N_VPWR_c_323_n N_VPWR_c_324_n N_VPWR_c_325_n
+ N_VPWR_c_326_n VPWR N_VPWR_c_327_n N_VPWR_c_316_n
+ PM_SKY130_FD_SC_MS__AND4_2%VPWR
x_PM_SKY130_FD_SC_MS__AND4_2%X N_X_M1002_s N_X_M1009_d X X X X N_X_c_367_n
+ PM_SKY130_FD_SC_MS__AND4_2%X
x_PM_SKY130_FD_SC_MS__AND4_2%VGND N_VGND_M1004_d N_VGND_M1008_d N_VGND_c_389_n
+ N_VGND_c_390_n N_VGND_c_391_n N_VGND_c_392_n N_VGND_c_393_n N_VGND_c_394_n
+ N_VGND_c_395_n VGND N_VGND_c_396_n N_VGND_c_397_n
+ PM_SKY130_FD_SC_MS__AND4_2%VGND
cc_1 VNB N_A_M1001_g 0.00155843f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.46
cc_2 VNB N_A_M1005_g 0.0287743f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.74
cc_3 VNB N_A_c_69_n 0.0547136f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_4 VNB N_A_c_70_n 0.013266f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.3
cc_5 VNB N_A_c_71_n 0.0086234f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.465
cc_6 VNB N_B_M1003_g 0.00695258f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.74
cc_7 VNB B 0.00459753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B_c_98_n 0.0308071f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.465
cc_9 VNB N_B_c_99_n 0.0180773f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.465
cc_10 VNB N_C_M1006_g 0.00710459f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.74
cc_11 VNB C 0.00242177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_C_c_135_n 0.0326376f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.465
cc_13 VNB N_C_c_136_n 0.0195889f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.465
cc_14 VNB N_D_c_168_n 0.00655899f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_15 VNB N_D_c_169_n 0.033522f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.465
cc_16 VNB N_D_c_170_n 0.0100678f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.465
cc_17 VNB N_D_c_171_n 0.0197696f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.465
cc_18 VNB N_A_56_74#_M1002_g 0.0225826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_56_74#_M1009_g 0.00335088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_56_74#_M1008_g 0.0273222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_56_74#_M1010_g 0.00156177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_56_74#_c_210_n 0.0366222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_56_74#_c_211_n 0.0258829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_56_74#_c_212_n 0.00377606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_56_74#_c_213_n 0.00710428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_56_74#_c_214_n 0.0577987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_56_74#_c_215_n 0.0094188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_316_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB X 0.00144878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_X_c_367_n 7.53866e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_389_n 0.0091706f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_32 VNB N_VGND_c_390_n 0.016267f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_33 VNB N_VGND_c_391_n 0.0111347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_392_n 0.0182112f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.465
cc_35 VNB N_VGND_c_393_n 0.0671414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_394_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.665
cc_37 VNB N_VGND_c_395_n 0.00867839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_396_n 0.0196671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_397_n 0.258397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VPB N_A_M1001_g 0.0343146f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=2.46
cc_41 VPB N_A_c_71_n 0.00823058f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.465
cc_42 VPB N_B_M1003_g 0.0307765f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=0.74
cc_43 VPB N_C_M1006_g 0.0309436f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=0.74
cc_44 VPB N_D_c_172_n 0.0244118f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.63
cc_45 VPB N_D_c_168_n 0.00740068f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_46 VPB N_A_56_74#_M1009_g 0.0240885f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_56_74#_M1010_g 0.0233476f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_56_74#_c_212_n 5.66269e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_56_74#_c_219_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_56_74#_c_220_n 0.0265271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A_56_74#_c_221_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_56_74#_c_222_n 0.00748573f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_56_74#_c_213_n 0.026491f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_56_74#_c_224_n 0.00692367f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_317_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.465
cc_56 VPB N_VPWR_c_318_n 0.0539876f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.465
cc_57 VPB N_VPWR_c_319_n 0.00987717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_320_n 0.00991277f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_321_n 0.0126718f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_322_n 0.0254067f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_323_n 0.0215645f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_324_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_325_n 0.0213997f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_326_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_327_n 0.0234846f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_316_n 0.0629723f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 N_A_M1001_g N_B_M1003_g 0.0146007f $X=0.595 $Y=2.46 $X2=0 $Y2=0
cc_68 N_A_M1005_g B 0.00235149f $X=0.64 $Y=0.74 $X2=0 $Y2=0
cc_69 N_A_c_70_n N_B_c_98_n 0.0449896f $X=0.505 $Y=1.3 $X2=0 $Y2=0
cc_70 N_A_M1005_g N_B_c_99_n 0.0303889f $X=0.64 $Y=0.74 $X2=0 $Y2=0
cc_71 N_A_M1005_g N_A_56_74#_c_211_n 0.0109243f $X=0.64 $Y=0.74 $X2=0 $Y2=0
cc_72 N_A_M1001_g N_A_56_74#_c_212_n 0.00179792f $X=0.595 $Y=2.46 $X2=0 $Y2=0
cc_73 N_A_M1005_g N_A_56_74#_c_212_n 0.00887397f $X=0.64 $Y=0.74 $X2=0 $Y2=0
cc_74 N_A_c_70_n N_A_56_74#_c_212_n 0.00952112f $X=0.505 $Y=1.3 $X2=0 $Y2=0
cc_75 N_A_c_71_n N_A_56_74#_c_212_n 0.030293f $X=0.28 $Y=1.465 $X2=0 $Y2=0
cc_76 N_A_M1001_g N_A_56_74#_c_219_n 0.019438f $X=0.595 $Y=2.46 $X2=0 $Y2=0
cc_77 N_A_M1005_g N_A_56_74#_c_215_n 0.0116482f $X=0.64 $Y=0.74 $X2=0 $Y2=0
cc_78 N_A_c_69_n N_A_56_74#_c_215_n 0.00605879f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_79 N_A_c_71_n N_A_56_74#_c_215_n 0.0143044f $X=0.28 $Y=1.465 $X2=0 $Y2=0
cc_80 N_A_M1001_g N_A_56_74#_c_224_n 0.00843804f $X=0.595 $Y=2.46 $X2=0 $Y2=0
cc_81 N_A_c_71_n N_A_56_74#_c_224_n 0.00503427f $X=0.28 $Y=1.465 $X2=0 $Y2=0
cc_82 N_A_M1001_g N_VPWR_c_318_n 0.0284032f $X=0.595 $Y=2.46 $X2=0 $Y2=0
cc_83 N_A_c_69_n N_VPWR_c_318_n 0.00181048f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_84 N_A_c_71_n N_VPWR_c_318_n 0.0299469f $X=0.28 $Y=1.465 $X2=0 $Y2=0
cc_85 N_A_M1001_g N_VPWR_c_323_n 0.0047558f $X=0.595 $Y=2.46 $X2=0 $Y2=0
cc_86 N_A_M1001_g N_VPWR_c_316_n 0.00839869f $X=0.595 $Y=2.46 $X2=0 $Y2=0
cc_87 N_A_M1005_g N_VGND_c_393_n 0.00434272f $X=0.64 $Y=0.74 $X2=0 $Y2=0
cc_88 N_A_M1005_g N_VGND_c_397_n 0.0082504f $X=0.64 $Y=0.74 $X2=0 $Y2=0
cc_89 N_B_M1003_g N_C_M1006_g 0.0291116f $X=1.045 $Y=2.46 $X2=0 $Y2=0
cc_90 B C 0.0744187f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_91 N_B_c_98_n C 3.9854e-19 $X=1.12 $Y=1.385 $X2=0 $Y2=0
cc_92 N_B_c_99_n C 7.46328e-19 $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_93 N_B_c_98_n N_C_c_135_n 0.0175135f $X=1.12 $Y=1.385 $X2=0 $Y2=0
cc_94 B N_C_c_136_n 0.00774327f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_95 N_B_c_99_n N_C_c_136_n 0.024906f $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_96 B N_A_56_74#_c_211_n 0.0212655f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_97 N_B_c_99_n N_A_56_74#_c_211_n 0.00182282f $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_98 B N_A_56_74#_c_212_n 0.031739f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_99 N_B_c_99_n N_A_56_74#_c_212_n 0.00586721f $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_100 N_B_M1003_g N_A_56_74#_c_219_n 0.016996f $X=1.045 $Y=2.46 $X2=0 $Y2=0
cc_101 N_B_M1003_g N_A_56_74#_c_220_n 0.0138724f $X=1.045 $Y=2.46 $X2=0 $Y2=0
cc_102 B N_A_56_74#_c_220_n 0.025829f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_103 N_B_c_98_n N_A_56_74#_c_220_n 0.00105742f $X=1.12 $Y=1.385 $X2=0 $Y2=0
cc_104 N_B_M1003_g N_A_56_74#_c_244_n 7.91299e-19 $X=1.045 $Y=2.46 $X2=0 $Y2=0
cc_105 B N_A_56_74#_c_215_n 0.0137062f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_106 N_B_c_99_n N_A_56_74#_c_215_n 9.65577e-19 $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_107 N_B_M1003_g N_A_56_74#_c_224_n 0.00282746f $X=1.045 $Y=2.46 $X2=0 $Y2=0
cc_108 B N_A_56_74#_c_224_n 0.00245488f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_109 N_B_M1003_g N_VPWR_c_319_n 0.0129189f $X=1.045 $Y=2.46 $X2=0 $Y2=0
cc_110 N_B_M1003_g N_VPWR_c_323_n 0.005209f $X=1.045 $Y=2.46 $X2=0 $Y2=0
cc_111 N_B_M1003_g N_VPWR_c_316_n 0.00984824f $X=1.045 $Y=2.46 $X2=0 $Y2=0
cc_112 B A_221_74# 0.00939544f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_113 B N_VGND_c_393_n 0.0102495f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_114 N_B_c_99_n N_VGND_c_393_n 0.00304348f $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_115 B N_VGND_c_397_n 0.0117398f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_116 N_B_c_99_n N_VGND_c_397_n 0.00371612f $X=1.12 $Y=1.22 $X2=0 $Y2=0
cc_117 N_C_M1006_g N_D_c_172_n 0.0140074f $X=1.705 $Y=2.46 $X2=-0.19 $Y2=-0.245
cc_118 N_C_M1006_g N_D_c_168_n 0.0110466f $X=1.705 $Y=2.46 $X2=0 $Y2=0
cc_119 C N_D_c_169_n 3.80049e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_120 N_C_c_135_n N_D_c_169_n 0.0174582f $X=1.69 $Y=1.385 $X2=0 $Y2=0
cc_121 C N_D_c_170_n 0.0273797f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_122 N_C_c_135_n N_D_c_170_n 0.00202602f $X=1.69 $Y=1.385 $X2=0 $Y2=0
cc_123 C N_D_c_171_n 0.00922273f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_124 N_C_c_136_n N_D_c_171_n 0.0242189f $X=1.69 $Y=1.22 $X2=0 $Y2=0
cc_125 N_C_M1006_g N_A_56_74#_c_219_n 9.35852e-19 $X=1.705 $Y=2.46 $X2=0 $Y2=0
cc_126 N_C_M1006_g N_A_56_74#_c_220_n 0.0167877f $X=1.705 $Y=2.46 $X2=0 $Y2=0
cc_127 C N_A_56_74#_c_220_n 0.0263044f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_128 N_C_c_135_n N_A_56_74#_c_220_n 0.00108599f $X=1.69 $Y=1.385 $X2=0 $Y2=0
cc_129 N_C_M1006_g N_A_56_74#_c_244_n 0.00782968f $X=1.705 $Y=2.46 $X2=0 $Y2=0
cc_130 N_C_M1006_g N_A_56_74#_c_221_n 0.0067134f $X=1.705 $Y=2.46 $X2=0 $Y2=0
cc_131 N_C_M1006_g N_A_56_74#_c_255_n 0.00216667f $X=1.705 $Y=2.46 $X2=0 $Y2=0
cc_132 N_C_M1006_g N_VPWR_c_319_n 0.0130077f $X=1.705 $Y=2.46 $X2=0 $Y2=0
cc_133 N_C_M1006_g N_VPWR_c_325_n 0.005209f $X=1.705 $Y=2.46 $X2=0 $Y2=0
cc_134 N_C_M1006_g N_VPWR_c_316_n 0.009846f $X=1.705 $Y=2.46 $X2=0 $Y2=0
cc_135 C A_335_74# 0.0102591f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_136 C N_VGND_c_393_n 0.00930091f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_137 N_C_c_136_n N_VGND_c_393_n 0.00304348f $X=1.69 $Y=1.22 $X2=0 $Y2=0
cc_138 C N_VGND_c_397_n 0.0106938f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_139 N_C_c_136_n N_VGND_c_397_n 0.00373154f $X=1.69 $Y=1.22 $X2=0 $Y2=0
cc_140 N_D_c_169_n N_A_56_74#_M1002_g 0.0181812f $X=2.26 $Y=1.385 $X2=0 $Y2=0
cc_141 N_D_c_170_n N_A_56_74#_M1002_g 0.00180549f $X=2.26 $Y=1.385 $X2=0 $Y2=0
cc_142 N_D_c_171_n N_A_56_74#_M1002_g 0.0138101f $X=2.26 $Y=1.22 $X2=0 $Y2=0
cc_143 N_D_c_168_n N_A_56_74#_M1009_g 0.0361195f $X=2.155 $Y=1.79 $X2=0 $Y2=0
cc_144 N_D_c_168_n N_A_56_74#_c_210_n 0.00174393f $X=2.155 $Y=1.79 $X2=0 $Y2=0
cc_145 N_D_c_172_n N_A_56_74#_c_220_n 0.00391559f $X=2.155 $Y=1.88 $X2=0 $Y2=0
cc_146 N_D_c_168_n N_A_56_74#_c_220_n 0.00235788f $X=2.155 $Y=1.79 $X2=0 $Y2=0
cc_147 N_D_c_170_n N_A_56_74#_c_220_n 0.00445923f $X=2.26 $Y=1.385 $X2=0 $Y2=0
cc_148 N_D_c_172_n N_A_56_74#_c_244_n 0.0100464f $X=2.155 $Y=1.88 $X2=0 $Y2=0
cc_149 N_D_c_172_n N_A_56_74#_c_221_n 0.00809344f $X=2.155 $Y=1.88 $X2=0 $Y2=0
cc_150 N_D_c_172_n N_A_56_74#_c_222_n 0.0151322f $X=2.155 $Y=1.88 $X2=0 $Y2=0
cc_151 N_D_c_172_n N_A_56_74#_c_255_n 4.64231e-19 $X=2.155 $Y=1.88 $X2=0 $Y2=0
cc_152 N_D_c_172_n N_VPWR_c_320_n 0.005335f $X=2.155 $Y=1.88 $X2=0 $Y2=0
cc_153 N_D_c_172_n N_VPWR_c_325_n 0.005209f $X=2.155 $Y=1.88 $X2=0 $Y2=0
cc_154 N_D_c_172_n N_VPWR_c_316_n 0.00534649f $X=2.155 $Y=1.88 $X2=0 $Y2=0
cc_155 N_D_c_168_n X 0.00261816f $X=2.155 $Y=1.79 $X2=0 $Y2=0
cc_156 N_D_c_169_n X 2.48447e-19 $X=2.26 $Y=1.385 $X2=0 $Y2=0
cc_157 N_D_c_170_n X 0.0146227f $X=2.26 $Y=1.385 $X2=0 $Y2=0
cc_158 N_D_c_171_n N_X_c_367_n 3.54267e-19 $X=2.26 $Y=1.22 $X2=0 $Y2=0
cc_159 N_D_c_169_n N_VGND_c_389_n 0.00103009f $X=2.26 $Y=1.385 $X2=0 $Y2=0
cc_160 N_D_c_170_n N_VGND_c_389_n 0.0122839f $X=2.26 $Y=1.385 $X2=0 $Y2=0
cc_161 N_D_c_171_n N_VGND_c_389_n 0.00413006f $X=2.26 $Y=1.22 $X2=0 $Y2=0
cc_162 N_D_c_171_n N_VGND_c_393_n 0.00461464f $X=2.26 $Y=1.22 $X2=0 $Y2=0
cc_163 N_D_c_171_n N_VGND_c_397_n 0.00910053f $X=2.26 $Y=1.22 $X2=0 $Y2=0
cc_164 N_A_56_74#_c_222_n N_VPWR_M1007_d 0.0166011f $X=3.405 $Y=2.405 $X2=0
+ $Y2=0
cc_165 N_A_56_74#_c_222_n N_VPWR_M1010_s 0.00615092f $X=3.405 $Y=2.405 $X2=0
+ $Y2=0
cc_166 N_A_56_74#_c_213_n N_VPWR_M1010_s 0.0115413f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_167 N_A_56_74#_c_219_n N_VPWR_c_318_n 0.080681f $X=0.82 $Y=2.105 $X2=0 $Y2=0
cc_168 N_A_56_74#_c_219_n N_VPWR_c_319_n 0.0571321f $X=0.82 $Y=2.105 $X2=0 $Y2=0
cc_169 N_A_56_74#_c_220_n N_VPWR_c_319_n 0.0271222f $X=1.765 $Y=1.805 $X2=0
+ $Y2=0
cc_170 N_A_56_74#_c_244_n N_VPWR_c_319_n 0.0165244f $X=1.93 $Y=2.105 $X2=0 $Y2=0
cc_171 N_A_56_74#_c_221_n N_VPWR_c_319_n 0.0312007f $X=1.93 $Y=2.815 $X2=0 $Y2=0
cc_172 N_A_56_74#_c_255_n N_VPWR_c_319_n 0.0114734f $X=1.93 $Y=2.405 $X2=0 $Y2=0
cc_173 N_A_56_74#_M1009_g N_VPWR_c_320_n 0.00569715f $X=2.775 $Y=2.4 $X2=0 $Y2=0
cc_174 N_A_56_74#_c_221_n N_VPWR_c_320_n 0.0110297f $X=1.93 $Y=2.815 $X2=0 $Y2=0
cc_175 N_A_56_74#_c_222_n N_VPWR_c_320_n 0.0259418f $X=3.405 $Y=2.405 $X2=0
+ $Y2=0
cc_176 N_A_56_74#_M1010_g N_VPWR_c_322_n 0.0115497f $X=3.225 $Y=2.4 $X2=0 $Y2=0
cc_177 N_A_56_74#_c_222_n N_VPWR_c_322_n 0.0306825f $X=3.405 $Y=2.405 $X2=0
+ $Y2=0
cc_178 N_A_56_74#_c_219_n N_VPWR_c_323_n 0.0161276f $X=0.82 $Y=2.105 $X2=0 $Y2=0
cc_179 N_A_56_74#_c_221_n N_VPWR_c_325_n 0.0144623f $X=1.93 $Y=2.815 $X2=0 $Y2=0
cc_180 N_A_56_74#_M1009_g N_VPWR_c_327_n 0.00553757f $X=2.775 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A_56_74#_M1010_g N_VPWR_c_327_n 0.00553757f $X=3.225 $Y=2.4 $X2=0 $Y2=0
cc_182 N_A_56_74#_M1009_g N_VPWR_c_316_n 0.00556599f $X=2.775 $Y=2.4 $X2=0 $Y2=0
cc_183 N_A_56_74#_M1010_g N_VPWR_c_316_n 0.00559162f $X=3.225 $Y=2.4 $X2=0 $Y2=0
cc_184 N_A_56_74#_c_219_n N_VPWR_c_316_n 0.0131188f $X=0.82 $Y=2.105 $X2=0 $Y2=0
cc_185 N_A_56_74#_c_221_n N_VPWR_c_316_n 0.0118344f $X=1.93 $Y=2.815 $X2=0 $Y2=0
cc_186 N_A_56_74#_c_222_n N_VPWR_c_316_n 0.0318244f $X=3.405 $Y=2.405 $X2=0
+ $Y2=0
cc_187 N_A_56_74#_c_222_n N_X_M1009_d 0.00479467f $X=3.405 $Y=2.405 $X2=0 $Y2=0
cc_188 N_A_56_74#_M1002_g X 0.00294214f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A_56_74#_M1009_g X 0.0153087f $X=2.775 $Y=2.4 $X2=0 $Y2=0
cc_190 N_A_56_74#_M1008_g X 0.0106301f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_191 N_A_56_74#_M1010_g X 0.0124113f $X=3.225 $Y=2.4 $X2=0 $Y2=0
cc_192 N_A_56_74#_c_210_n X 0.025387f $X=3.315 $Y=1.465 $X2=0 $Y2=0
cc_193 N_A_56_74#_c_222_n X 0.0223581f $X=3.405 $Y=2.405 $X2=0 $Y2=0
cc_194 N_A_56_74#_c_213_n X 0.0663601f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_195 N_A_56_74#_M1002_g N_X_c_367_n 0.00713606f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A_56_74#_M1008_g N_X_c_367_n 0.0119323f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A_56_74#_c_215_n A_143_74# 0.00178387f $X=0.7 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_198 N_A_56_74#_M1002_g N_VGND_c_389_n 0.0125291f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A_56_74#_M1002_g N_VGND_c_391_n 0.00110029f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A_56_74#_M1008_g N_VGND_c_391_n 0.00595376f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A_56_74#_M1008_g N_VGND_c_392_n 0.0103157f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A_56_74#_c_213_n N_VGND_c_392_n 0.0178142f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_203 N_A_56_74#_c_214_n N_VGND_c_392_n 0.00190129f $X=3.57 $Y=1.465 $X2=0
+ $Y2=0
cc_204 N_A_56_74#_c_211_n N_VGND_c_393_n 0.0144497f $X=0.425 $Y=0.515 $X2=0
+ $Y2=0
cc_205 N_A_56_74#_M1008_g N_VGND_c_395_n 0.00481221f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A_56_74#_c_210_n N_VGND_c_395_n 0.00345718f $X=3.315 $Y=1.465 $X2=0
+ $Y2=0
cc_207 N_A_56_74#_M1002_g N_VGND_c_396_n 0.00461464f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A_56_74#_M1008_g N_VGND_c_396_n 0.00383152f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A_56_74#_M1002_g N_VGND_c_397_n 0.00835925f $X=2.74 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A_56_74#_M1008_g N_VGND_c_397_n 0.0036906f $X=3.17 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A_56_74#_c_211_n N_VGND_c_397_n 0.0119539f $X=0.425 $Y=0.515 $X2=0
+ $Y2=0
cc_212 N_X_c_367_n N_VGND_c_389_n 0.017139f $X=2.955 $Y=0.91 $X2=0 $Y2=0
cc_213 N_X_c_367_n N_VGND_c_392_n 0.0241034f $X=2.955 $Y=0.91 $X2=0 $Y2=0
cc_214 N_X_c_367_n N_VGND_c_395_n 0.00106652f $X=2.955 $Y=0.91 $X2=0 $Y2=0
cc_215 N_X_c_367_n N_VGND_c_397_n 0.0167375f $X=2.955 $Y=0.91 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__mux2_4.pex.spice
* Created: Wed Sep  2 12:11:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__MUX2_4%S 3 7 11 15 19 23 26 27 28 29 32 33 35 38 42
+ 45 46 54
c136 54 0 1.32825e-20 $X=3.985 $Y=1.6
c137 35 0 1.42621e-19 $X=3.58 $Y=1.6
c138 15 0 1.78467e-19 $X=3.535 $Y=2.455
c139 3 0 7.82978e-20 $X=0.505 $Y=2.34
r140 53 54 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.97 $Y=1.6
+ $X2=3.985 $Y2=1.6
r141 49 51 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=3.47 $Y=1.6
+ $X2=3.535 $Y2=1.6
r142 45 48 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.515
+ $X2=0.585 $Y2=1.68
r143 45 47 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.515
+ $X2=0.585 $Y2=1.35
r144 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.515 $X2=0.59 $Y2=1.515
r145 42 60 7.28531 $w=4.08e-07 $l=1.15e-07 $layer=LI1_cond $X=0.63 $Y=1.665
+ $X2=0.63 $Y2=1.78
r146 42 46 4.21625 $w=4.08e-07 $l=1.5e-07 $layer=LI1_cond $X=0.63 $Y=1.665
+ $X2=0.63 $Y2=1.515
r147 38 40 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.59 $Y=2.135
+ $X2=1.59 $Y2=2.24
r148 36 53 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=3.58 $Y=1.6
+ $X2=3.97 $Y2=1.6
r149 36 51 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=3.58 $Y=1.6
+ $X2=3.535 $Y2=1.6
r150 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.58
+ $Y=1.6 $X2=3.58 $Y2=1.6
r151 33 35 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=3.165 $Y=1.6
+ $X2=3.58 $Y2=1.6
r152 31 33 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.08 $Y=1.765
+ $X2=3.165 $Y2=1.6
r153 31 32 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.08 $Y=1.765
+ $X2=3.08 $Y2=2.155
r154 30 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.675 $Y=2.24
+ $X2=1.59 $Y2=2.24
r155 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.995 $Y=2.24
+ $X2=3.08 $Y2=2.155
r156 29 30 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=2.995 $Y=2.24
+ $X2=1.675 $Y2=2.24
r157 27 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.505 $Y=2.135
+ $X2=1.59 $Y2=2.135
r158 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.505 $Y=2.135
+ $X2=0.835 $Y2=2.135
r159 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.75 $Y=2.05
+ $X2=0.835 $Y2=2.135
r160 26 60 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.75 $Y=2.05
+ $X2=0.75 $Y2=1.78
r161 21 54 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.985 $Y=1.765
+ $X2=3.985 $Y2=1.6
r162 21 23 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=3.985 $Y=1.765
+ $X2=3.985 $Y2=2.455
r163 17 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.97 $Y=1.435
+ $X2=3.97 $Y2=1.6
r164 17 19 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=3.97 $Y=1.435
+ $X2=3.97 $Y2=0.915
r165 13 51 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.535 $Y=1.765
+ $X2=3.535 $Y2=1.6
r166 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=3.535 $Y=1.765
+ $X2=3.535 $Y2=2.455
r167 9 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.47 $Y=1.435
+ $X2=3.47 $Y2=1.6
r168 9 11 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=3.47 $Y=1.435
+ $X2=3.47 $Y2=0.915
r169 7 47 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=0.65 $Y=0.81
+ $X2=0.65 $Y2=1.35
r170 3 48 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=0.505 $Y=2.34
+ $X2=0.505 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2_4%A_27_368# 1 2 9 13 17 21 26 27 28 29 32 33 34
+ 36 37 39 43 47 48 49 58
c136 58 0 1.42621e-19 $X=5.055 $Y=1.6
c137 47 0 1.47206e-19 $X=0.28 $Y=2.115
c138 29 0 5.64602e-20 $X=3.335 $Y=2.58
r139 57 58 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.04 $Y=1.6
+ $X2=5.055 $Y2=1.6
r140 53 55 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=4.605 $Y=1.6
+ $X2=4.61 $Y2=1.6
r141 49 51 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.25 $Y=2.475
+ $X2=1.25 $Y2=2.58
r142 47 48 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.265 $Y=2.115
+ $X2=0.265 $Y2=1.95
r143 45 48 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=0.17 $Y=1.15 $X2=0.17
+ $Y2=1.95
r144 43 45 17.7387 $w=5.13e-07 $l=5.15e-07 $layer=LI1_cond $X=0.342 $Y=0.635
+ $X2=0.342 $Y2=1.15
r145 40 57 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=4.82 $Y=1.6
+ $X2=5.04 $Y2=1.6
r146 40 55 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.82 $Y=1.6
+ $X2=4.61 $Y2=1.6
r147 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.82
+ $Y=1.6 $X2=4.82 $Y2=1.6
r148 37 39 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=4.085 $Y=1.6
+ $X2=4.82 $Y2=1.6
r149 35 37 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=4 $Y=1.765
+ $X2=4.085 $Y2=1.6
r150 35 36 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4 $Y=1.765 $X2=4
+ $Y2=1.935
r151 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.915 $Y=2.02
+ $X2=4 $Y2=1.935
r152 33 34 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.915 $Y=2.02
+ $X2=3.505 $Y2=2.02
r153 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.42 $Y=2.105
+ $X2=3.505 $Y2=2.02
r154 31 32 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.42 $Y=2.105
+ $X2=3.42 $Y2=2.495
r155 30 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.335 $Y=2.58
+ $X2=1.25 $Y2=2.58
r156 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.335 $Y=2.58
+ $X2=3.42 $Y2=2.495
r157 29 30 130.481 $w=1.68e-07 $l=2e-06 $layer=LI1_cond $X=3.335 $Y=2.58
+ $X2=1.335 $Y2=2.58
r158 27 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.165 $Y=2.475
+ $X2=1.25 $Y2=2.475
r159 27 28 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.165 $Y=2.475
+ $X2=0.445 $Y2=2.475
r160 26 28 8.02311 $w=1.7e-07 $l=2.18403e-07 $layer=LI1_cond $X=0.265 $Y=2.39
+ $X2=0.445 $Y2=2.475
r161 25 47 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=0.265 $Y=2.13
+ $X2=0.265 $Y2=2.115
r162 25 26 8.3232 $w=3.58e-07 $l=2.6e-07 $layer=LI1_cond $X=0.265 $Y=2.13
+ $X2=0.265 $Y2=2.39
r163 19 58 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.055 $Y=1.765
+ $X2=5.055 $Y2=1.6
r164 19 21 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=5.055 $Y=1.765
+ $X2=5.055 $Y2=2.455
r165 15 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.04 $Y=1.435
+ $X2=5.04 $Y2=1.6
r166 15 17 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=5.04 $Y=1.435
+ $X2=5.04 $Y2=0.915
r167 11 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.61 $Y=1.435
+ $X2=4.61 $Y2=1.6
r168 11 13 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=4.61 $Y=1.435
+ $X2=4.61 $Y2=0.915
r169 7 53 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.605 $Y=1.765
+ $X2=4.605 $Y2=1.6
r170 7 9 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=4.605 $Y=1.765
+ $X2=4.605 $Y2=2.455
r171 2 47 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r172 1 43 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.29
+ $Y=0.49 $X2=0.435 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2_4%A_193_241# 1 2 3 4 5 6 21 26 27 28 29 31 36
+ 37 42 43 45 47 52 53 55 57 60 63 66 67 69 74 81 85 86 87 92 96 98 103 106 109
+ 111 112 113 114 116 117
c219 43 0 5.9954e-20 $X=2.295 $Y=1.295
c220 21 0 3.09329e-19 $X=1.055 $Y=2.4
r221 117 122 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.78 $Y=1.615
+ $X2=5.705 $Y2=1.615
r222 111 112 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=6.425 $Y=0.427
+ $X2=6.59 $Y2=0.427
r223 109 116 5.16603 $w=2.5e-07 $l=1.60078e-07 $layer=LI1_cond $X=8.44 $Y=1.95
+ $X2=8.36 $Y2=2.075
r224 109 114 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.44 $Y=1.95
+ $X2=8.44 $Y2=1.03
r225 104 116 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=8.36 $Y=2.2
+ $X2=8.36 $Y2=2.075
r226 104 106 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=8.36 $Y=2.2
+ $X2=8.36 $Y2=2.465
r227 101 114 8.53494 $w=3.33e-07 $l=1.67e-07 $layer=LI1_cond $X=8.357 $Y=0.863
+ $X2=8.357 $Y2=1.03
r228 101 103 11.9716 $w=3.33e-07 $l=3.48e-07 $layer=LI1_cond $X=8.357 $Y=0.863
+ $X2=8.357 $Y2=0.515
r229 100 103 3.09612 $w=3.33e-07 $l=9e-08 $layer=LI1_cond $X=8.357 $Y=0.425
+ $X2=8.357 $Y2=0.515
r230 99 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.59 $Y=0.34
+ $X2=7.425 $Y2=0.34
r231 98 100 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=8.19 $Y=0.34
+ $X2=8.357 $Y2=0.425
r232 98 99 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=8.19 $Y=0.34 $X2=7.59
+ $Y2=0.34
r233 94 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.425 $Y=0.425
+ $X2=7.425 $Y2=0.34
r234 94 96 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=7.425 $Y=0.425
+ $X2=7.425 $Y2=0.495
r235 92 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.26 $Y=0.34
+ $X2=7.425 $Y2=0.34
r236 92 112 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.26 $Y=0.34
+ $X2=6.59 $Y2=0.34
r237 89 91 42.6404 $w=2.48e-07 $l=9.25e-07 $layer=LI1_cond $X=6.48 $Y=2.075
+ $X2=7.405 $Y2=2.075
r238 87 89 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=6.47 $Y=2.075
+ $X2=6.48 $Y2=2.075
r239 86 116 1.34256 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=8.195 $Y=2.075
+ $X2=8.36 $Y2=2.075
r240 86 91 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=8.195 $Y=2.075
+ $X2=7.405 $Y2=2.075
r241 85 87 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.385 $Y=1.95
+ $X2=6.47 $Y2=2.075
r242 84 85 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.385 $Y=1.78
+ $X2=6.385 $Y2=1.95
r243 81 117 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=6.23 $Y=1.615
+ $X2=5.78 $Y2=1.615
r244 80 81 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.23
+ $Y=1.615 $X2=6.23 $Y2=1.615
r245 77 122 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=5.55 $Y=1.615
+ $X2=5.705 $Y2=1.615
r246 76 80 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.55 $Y=1.615
+ $X2=6.23 $Y2=1.615
r247 76 77 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.55
+ $Y=1.615 $X2=5.55 $Y2=1.615
r248 74 84 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.3 $Y=1.615
+ $X2=6.385 $Y2=1.78
r249 74 80 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=6.3 $Y=1.615 $X2=6.23
+ $Y2=1.615
r250 60 122 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.705 $Y=1.45
+ $X2=5.705 $Y2=1.615
r251 59 60 612.755 $w=1.5e-07 $l=1.195e-06 $layer=POLY_cond $X=5.705 $Y=0.255
+ $X2=5.705 $Y2=1.45
r252 55 70 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.915 $Y=1.385
+ $X2=2.71 $Y2=1.385
r253 55 57 365.387 $w=1.8e-07 $l=9.4e-07 $layer=POLY_cond $X=2.915 $Y=1.46
+ $X2=2.915 $Y2=2.4
r254 54 69 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.785 $Y=0.18
+ $X2=2.71 $Y2=0.18
r255 53 59 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.63 $Y=0.18
+ $X2=5.705 $Y2=0.255
r256 53 54 1458.82 $w=1.5e-07 $l=2.845e-06 $layer=POLY_cond $X=5.63 $Y=0.18
+ $X2=2.785 $Y2=0.18
r257 50 70 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.71 $Y=1.31
+ $X2=2.71 $Y2=1.385
r258 50 52 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.71 $Y=1.31
+ $X2=2.71 $Y2=0.76
r259 49 69 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.71 $Y=0.255
+ $X2=2.71 $Y2=0.18
r260 49 52 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.71 $Y=0.255
+ $X2=2.71 $Y2=0.76
r261 48 67 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.355 $Y=0.18
+ $X2=2.28 $Y2=0.18
r262 47 69 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.635 $Y=0.18
+ $X2=2.71 $Y2=0.18
r263 47 48 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.635 $Y=0.18
+ $X2=2.355 $Y2=0.18
r264 43 68 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.295 $Y=1.295
+ $X2=2.295 $Y2=1.205
r265 43 45 429.524 $w=1.8e-07 $l=1.105e-06 $layer=POLY_cond $X=2.295 $Y=1.295
+ $X2=2.295 $Y2=2.4
r266 42 68 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.28 $Y=0.76
+ $X2=2.28 $Y2=1.205
r267 39 67 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.28 $Y=0.255
+ $X2=2.28 $Y2=0.18
r268 39 42 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.28 $Y=0.255
+ $X2=2.28 $Y2=0.76
r269 38 66 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=0.18
+ $X2=1.69 $Y2=0.18
r270 37 67 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.205 $Y=0.18
+ $X2=2.28 $Y2=0.18
r271 37 38 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=2.205 $Y=0.18
+ $X2=1.765 $Y2=0.18
r272 36 65 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.69 $Y=0.76
+ $X2=1.69 $Y2=1.205
r273 33 66 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=0.255
+ $X2=1.69 $Y2=0.18
r274 33 36 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.69 $Y=0.255
+ $X2=1.69 $Y2=0.76
r275 29 65 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.675 $Y=1.295
+ $X2=1.675 $Y2=1.205
r276 29 31 429.524 $w=1.8e-07 $l=1.105e-06 $layer=POLY_cond $X=1.675 $Y=1.295
+ $X2=1.675 $Y2=2.4
r277 27 66 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.615 $Y=0.18
+ $X2=1.69 $Y2=0.18
r278 27 28 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.615 $Y=0.18
+ $X2=1.295 $Y2=0.18
r279 24 63 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.22 $Y=1.205
+ $X2=1.22 $Y2=1.28
r280 24 26 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.22 $Y=1.205
+ $X2=1.22 $Y2=0.76
r281 23 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.22 $Y=0.255
+ $X2=1.295 $Y2=0.18
r282 23 26 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.22 $Y=0.255
+ $X2=1.22 $Y2=0.76
r283 19 63 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.28
+ $X2=1.22 $Y2=1.28
r284 19 21 406.202 $w=1.8e-07 $l=1.045e-06 $layer=POLY_cond $X=1.055 $Y=1.355
+ $X2=1.055 $Y2=2.4
r285 6 116 600 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_PDIFF $count=1 $X=8.175
+ $Y=1.96 $X2=8.36 $Y2=2.115
r286 6 106 300 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_PDIFF $count=2 $X=8.175
+ $Y=1.96 $X2=8.36 $Y2=2.465
r287 5 91 600 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=7.265
+ $Y=1.96 $X2=7.405 $Y2=2.115
r288 4 89 600 $w=1.7e-07 $l=2.24499e-07 $layer=licon1_PDIFF $count=1 $X=6.32
+ $Y=1.96 $X2=6.48 $Y2=2.115
r289 3 103 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=8.175
+ $Y=0.37 $X2=8.355 $Y2=0.515
r290 2 96 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=7.235
+ $Y=0.37 $X2=7.425 $Y2=0.495
r291 1 111 91 $w=1.7e-07 $l=6.38396e-07 $layer=licon1_NDIFF $count=2 $X=5.855
+ $Y=0.37 $X2=6.425 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2_4%A0 3 7 11 15 17 24
r44 24 25 2.24534 $w=3.22e-07 $l=1.5e-08 $layer=POLY_cond $X=7.16 $Y=1.615
+ $X2=7.175 $Y2=1.615
r45 22 24 53.1398 $w=3.22e-07 $l=3.55e-07 $layer=POLY_cond $X=6.805 $Y=1.615
+ $X2=7.16 $Y2=1.615
r46 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.805
+ $Y=1.615 $X2=6.805 $Y2=1.615
r47 20 22 11.9752 $w=3.22e-07 $l=8e-08 $layer=POLY_cond $X=6.725 $Y=1.615
+ $X2=6.805 $Y2=1.615
r48 19 20 2.24534 $w=3.22e-07 $l=1.5e-08 $layer=POLY_cond $X=6.71 $Y=1.615
+ $X2=6.725 $Y2=1.615
r49 17 23 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=6.96 $Y=1.615
+ $X2=6.805 $Y2=1.615
r50 13 25 16.3606 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.175 $Y=1.78
+ $X2=7.175 $Y2=1.615
r51 13 15 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=7.175 $Y=1.78
+ $X2=7.175 $Y2=2.46
r52 9 24 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.16 $Y=1.45
+ $X2=7.16 $Y2=1.615
r53 9 11 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=7.16 $Y=1.45 $X2=7.16
+ $Y2=0.69
r54 5 20 16.3606 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.725 $Y=1.78
+ $X2=6.725 $Y2=1.615
r55 5 7 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=6.725 $Y=1.78
+ $X2=6.725 $Y2=2.46
r56 1 19 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.71 $Y=1.45
+ $X2=6.71 $Y2=1.615
r57 1 3 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=6.71 $Y=1.45 $X2=6.71
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2_4%A1 3 7 11 15 17 18 26 28
r46 27 28 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=8.085 $Y=1.615
+ $X2=8.1 $Y2=1.615
r47 25 27 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.01 $Y=1.615
+ $X2=8.085 $Y2=1.615
r48 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.01
+ $Y=1.615 $X2=8.01 $Y2=1.615
r49 23 25 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=7.64 $Y=1.615
+ $X2=8.01 $Y2=1.615
r50 21 23 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=7.635 $Y=1.615
+ $X2=7.64 $Y2=1.615
r51 18 26 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=7.92 $Y=1.615 $X2=8.01
+ $Y2=1.615
r52 17 18 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.615
+ $X2=7.92 $Y2=1.615
r53 13 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.1 $Y=1.45 $X2=8.1
+ $Y2=1.615
r54 13 15 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=8.1 $Y=1.45 $X2=8.1
+ $Y2=0.69
r55 9 27 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.085 $Y=1.78
+ $X2=8.085 $Y2=1.615
r56 9 11 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=8.085 $Y=1.78
+ $X2=8.085 $Y2=2.46
r57 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.64 $Y=1.45
+ $X2=7.64 $Y2=1.615
r58 5 7 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=7.64 $Y=1.45 $X2=7.64
+ $Y2=0.69
r59 1 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.635 $Y=1.78
+ $X2=7.635 $Y2=1.615
r60 1 3 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=7.635 $Y=1.78
+ $X2=7.635 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2_4%VPWR 1 2 3 4 5 20 24 28 32 36 39 40 42 43 45
+ 46 47 53 68 69 72 75
r101 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r102 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r103 68 69 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r104 66 69 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=8.4 $Y2=3.33
r105 65 68 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=8.4 $Y2=3.33
r106 65 66 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r107 63 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r108 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r109 60 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r110 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r111 57 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.39 $Y=3.33
+ $X2=3.225 $Y2=3.33
r112 57 59 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.39 $Y=3.33
+ $X2=4.08 $Y2=3.33
r113 56 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r114 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r115 53 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.06 $Y=3.33
+ $X2=3.225 $Y2=3.33
r116 53 55 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=3.06 $Y=3.33 $X2=2.16
+ $Y2=3.33
r117 52 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r118 52 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r119 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r120 49 72 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=0.822 $Y2=3.33
r121 49 51 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=1.68 $Y2=3.33
r122 47 63 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=5.04 $Y2=3.33
r123 47 60 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r124 45 62 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.2 $Y=3.33
+ $X2=5.04 $Y2=3.33
r125 45 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.2 $Y=3.33
+ $X2=5.325 $Y2=3.33
r126 44 65 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=5.45 $Y=3.33 $X2=5.52
+ $Y2=3.33
r127 44 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.45 $Y=3.33
+ $X2=5.325 $Y2=3.33
r128 42 59 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=4.13 $Y=3.33 $X2=4.08
+ $Y2=3.33
r129 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.13 $Y=3.33
+ $X2=4.295 $Y2=3.33
r130 41 62 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.46 $Y=3.33
+ $X2=5.04 $Y2=3.33
r131 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.46 $Y=3.33
+ $X2=4.295 $Y2=3.33
r132 39 51 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.82 $Y=3.33
+ $X2=1.68 $Y2=3.33
r133 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.82 $Y=3.33
+ $X2=1.985 $Y2=3.33
r134 38 55 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=2.15 $Y=3.33
+ $X2=2.16 $Y2=3.33
r135 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.15 $Y=3.33
+ $X2=1.985 $Y2=3.33
r136 34 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.325 $Y=3.245
+ $X2=5.325 $Y2=3.33
r137 34 36 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=5.325 $Y=3.245
+ $X2=5.325 $Y2=2.94
r138 30 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.295 $Y=3.245
+ $X2=4.295 $Y2=3.33
r139 30 32 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.295 $Y=3.245
+ $X2=4.295 $Y2=2.94
r140 26 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.225 $Y=3.245
+ $X2=3.225 $Y2=3.33
r141 26 28 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=3.225 $Y=3.245
+ $X2=3.225 $Y2=3
r142 22 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=3.245
+ $X2=1.985 $Y2=3.33
r143 22 24 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=1.985 $Y=3.245
+ $X2=1.985 $Y2=3
r144 18 72 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=0.822 $Y=3.245
+ $X2=0.822 $Y2=3.33
r145 18 20 14.3638 $w=3.43e-07 $l=4.3e-07 $layer=LI1_cond $X=0.822 $Y=3.245
+ $X2=0.822 $Y2=2.815
r146 5 36 600 $w=1.7e-07 $l=1.08946e-06 $layer=licon1_PDIFF $count=1 $X=5.145
+ $Y=1.955 $X2=5.365 $Y2=2.94
r147 4 32 600 $w=1.7e-07 $l=1.08946e-06 $layer=licon1_PDIFF $count=1 $X=4.075
+ $Y=1.955 $X2=4.295 $Y2=2.94
r148 3 28 600 $w=1.7e-07 $l=1.26523e-06 $layer=licon1_PDIFF $count=1 $X=3.005
+ $Y=1.84 $X2=3.225 $Y2=3
r149 2 24 600 $w=1.7e-07 $l=1.26523e-06 $layer=licon1_PDIFF $count=1 $X=1.765
+ $Y=1.84 $X2=1.985 $Y2=3
r150 1 20 600 $w=1.7e-07 $l=1.08167e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.82 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2_4%X 1 2 3 4 13 15 17 19 21 23 24 30 33
c58 30 0 2.54869e-20 $X=2.33 $Y=1.625
c59 17 0 1.32825e-20 $X=2.542 $Y=1.37
c60 15 0 1.62123e-19 $X=1.475 $Y=0.535
c61 13 0 1.09271e-19 $X=1.475 $Y=1.37
r62 31 33 0.938101 $w=5.08e-07 $l=4e-08 $layer=LI1_cond $X=1.64 $Y=1.625
+ $X2=1.68 $Y2=1.625
r63 24 30 3.19265 $w=5.1e-07 $l=2.44622e-07 $layer=LI1_cond $X=2.55 $Y=1.677
+ $X2=2.33 $Y2=1.625
r64 23 30 3.98693 $w=5.08e-07 $l=1.7e-07 $layer=LI1_cond $X=2.16 $Y=1.625
+ $X2=2.33 $Y2=1.625
r65 21 31 3.11208 $w=5.1e-07 $l=2.78e-07 $layer=LI1_cond $X=1.362 $Y=1.625
+ $X2=1.64 $Y2=1.625
r66 21 23 10.7413 $w=5.08e-07 $l=4.58e-07 $layer=LI1_cond $X=1.702 $Y=1.625
+ $X2=2.16 $Y2=1.625
r67 21 33 0.515955 $w=5.08e-07 $l=2.2e-08 $layer=LI1_cond $X=1.702 $Y=1.625
+ $X2=1.68 $Y2=1.625
r68 17 24 3.69737 $w=4.25e-07 $l=3.10974e-07 $layer=LI1_cond $X=2.542 $Y=1.37
+ $X2=2.55 $Y2=1.677
r69 17 19 22.6421 $w=4.23e-07 $l=8.35e-07 $layer=LI1_cond $X=2.542 $Y=1.37
+ $X2=2.542 $Y2=0.535
r70 13 21 4.11959 $w=3.3e-07 $l=3.06333e-07 $layer=LI1_cond $X=1.475 $Y=1.37
+ $X2=1.362 $Y2=1.625
r71 13 15 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=1.475 $Y=1.37
+ $X2=1.475 $Y2=0.535
r72 4 24 600 $w=1.7e-07 $l=2.48193e-07 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=1.84 $X2=2.605 $Y2=1.9
r73 3 21 600 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.84 $X2=1.365 $Y2=1.795
r74 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.355
+ $Y=0.39 $X2=2.495 $Y2=0.535
r75 1 15 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=1.295
+ $Y=0.39 $X2=1.475 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2_4%A_725_391# 1 2 9 13 16 17
c46 16 0 1.78467e-19 $X=3.76 $Y=2.44
r47 11 17 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.705 $Y=2.845
+ $X2=5.705 $Y2=2.52
r48 11 13 49.5124 $w=2.68e-07 $l=1.16e-06 $layer=LI1_cond $X=5.79 $Y=2.845
+ $X2=6.95 $Y2=2.845
r49 10 16 3.9577 $w=1.7e-07 $l=1.60078e-07 $layer=LI1_cond $X=3.925 $Y=2.52
+ $X2=3.8 $Y2=2.44
r50 9 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.62 $Y=2.52
+ $X2=5.705 $Y2=2.52
r51 9 10 110.583 $w=1.68e-07 $l=1.695e-06 $layer=LI1_cond $X=5.62 $Y=2.52
+ $X2=3.925 $Y2=2.52
r52 2 13 600 $w=1.7e-07 $l=9.1e-07 $layer=licon1_PDIFF $count=1 $X=6.815 $Y=1.96
+ $X2=6.95 $Y2=2.805
r53 1 16 300 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=2 $X=3.625
+ $Y=1.955 $X2=3.76 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2_4%A_939_391# 1 2 7 9 16 17 22
r47 17 19 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.045 $Y=2.18
+ $X2=6.045 $Y2=2.455
r48 14 16 13.5259 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=4.83 $Y=2.1 $X2=5.14
+ $Y2=2.1
r49 10 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.13 $Y=2.455
+ $X2=6.045 $Y2=2.455
r50 9 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.695 $Y=2.455
+ $X2=7.86 $Y2=2.455
r51 9 10 102.102 $w=1.68e-07 $l=1.565e-06 $layer=LI1_cond $X=7.695 $Y=2.455
+ $X2=6.13 $Y2=2.455
r52 7 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.96 $Y=2.18
+ $X2=6.045 $Y2=2.18
r53 7 16 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=5.96 $Y=2.18 $X2=5.14
+ $Y2=2.18
r54 2 22 300 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=2 $X=7.725
+ $Y=1.96 $X2=7.86 $Y2=2.455
r55 1 14 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.695
+ $Y=1.955 $X2=4.83 $Y2=2.1
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2_4%VGND 1 2 3 4 5 18 22 26 30 34 38 41 42 44 45
+ 46 55 59 66 67 70 73 76
c106 26 0 5.9954e-20 $X=3.09 $Y=0.535
r107 76 77 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r108 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r109 71 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r110 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r111 67 77 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=8.4 $Y=0 $X2=5.52
+ $Y2=0
r112 66 67 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r113 64 76 9.89127 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=5.575 $Y=0
+ $X2=5.372 $Y2=0
r114 64 66 184.305 $w=1.68e-07 $l=2.825e-06 $layer=LI1_cond $X=5.575 $Y=0
+ $X2=8.4 $Y2=0
r115 63 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r116 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r117 60 73 10.873 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=4.49 $Y=0 $X2=4.255
+ $Y2=0
r118 60 62 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=4.49 $Y=0 $X2=5.04
+ $Y2=0
r119 59 76 9.89127 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=5.17 $Y=0 $X2=5.372
+ $Y2=0
r120 59 62 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=5.17 $Y=0 $X2=5.04
+ $Y2=0
r121 58 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r122 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r123 55 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.925 $Y=0 $X2=3.09
+ $Y2=0
r124 55 57 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.925 $Y=0
+ $X2=2.64 $Y2=0
r125 54 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r126 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r127 50 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r128 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r129 46 63 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.32 $Y=0 $X2=5.04
+ $Y2=0
r130 46 74 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.08 $Y2=0
r131 44 53 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.81 $Y=0 $X2=1.68
+ $Y2=0
r132 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.81 $Y=0 $X2=1.975
+ $Y2=0
r133 43 57 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.14 $Y=0 $X2=2.64
+ $Y2=0
r134 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.14 $Y=0 $X2=1.975
+ $Y2=0
r135 41 49 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=0.77 $Y=0 $X2=0.72
+ $Y2=0
r136 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=0 $X2=0.935
+ $Y2=0
r137 40 53 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=1.1 $Y=0 $X2=1.68
+ $Y2=0
r138 40 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.1 $Y=0 $X2=0.935
+ $Y2=0
r139 36 76 1.50354 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.372 $Y=0.085
+ $X2=5.372 $Y2=0
r140 36 38 11.809 $w=4.03e-07 $l=4.15e-07 $layer=LI1_cond $X=5.372 $Y=0.085
+ $X2=5.372 $Y2=0.5
r141 32 73 1.91284 $w=4.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.255 $Y=0.085
+ $X2=4.255 $Y2=0
r142 32 34 16.6688 $w=4.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.255 $Y=0.085
+ $X2=4.255 $Y2=0.74
r143 31 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.09
+ $Y2=0
r144 30 73 10.873 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=4.02 $Y=0 $X2=4.255
+ $Y2=0
r145 30 31 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=4.02 $Y=0
+ $X2=3.255 $Y2=0
r146 26 28 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=3.09 $Y=0.535
+ $X2=3.09 $Y2=1.09
r147 24 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.09 $Y=0.085
+ $X2=3.09 $Y2=0
r148 24 26 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.09 $Y=0.085
+ $X2=3.09 $Y2=0.535
r149 20 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.975 $Y=0.085
+ $X2=1.975 $Y2=0
r150 20 22 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.975 $Y=0.085
+ $X2=1.975 $Y2=0.535
r151 16 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.935 $Y=0.085
+ $X2=0.935 $Y2=0
r152 16 18 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=0.935 $Y=0.085
+ $X2=0.935 $Y2=0.635
r153 5 38 182 $w=1.7e-07 $l=2.98747e-07 $layer=licon1_NDIFF $count=1 $X=5.115
+ $Y=0.595 $X2=5.37 $Y2=0.5
r154 4 34 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=4.045
+ $Y=0.595 $X2=4.255 $Y2=0.74
r155 3 28 182 $w=1.7e-07 $l=8.38749e-07 $layer=licon1_NDIFF $count=1 $X=2.785
+ $Y=0.39 $X2=3.09 $Y2=1.09
r156 3 26 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=2.785
+ $Y=0.39 $X2=3.09 $Y2=0.535
r157 2 22 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.765
+ $Y=0.39 $X2=1.975 $Y2=0.535
r158 1 18 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=0.725
+ $Y=0.49 $X2=0.935 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2_4%A_709_119# 1 2 9 12 13 17 19 20
r60 19 20 10.1916 $w=1.83e-07 $l=1.7e-07 $layer=LI1_cond $X=5.155 $Y=1.187
+ $X2=5.325 $Y2=1.187
r61 15 17 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=7.895 $Y=1.11
+ $X2=7.895 $Y2=0.81
r62 13 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.77 $Y=1.195
+ $X2=7.895 $Y2=1.11
r63 13 20 159.513 $w=1.68e-07 $l=2.445e-06 $layer=LI1_cond $X=7.77 $Y=1.195
+ $X2=5.325 $Y2=1.195
r64 12 19 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=3.85 $Y=1.18
+ $X2=5.155 $Y2=1.18
r65 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.685 $Y=1.095
+ $X2=3.85 $Y2=1.18
r66 7 9 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.685 $Y=1.095
+ $X2=3.685 $Y2=0.74
r67 2 17 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=7.715
+ $Y=0.37 $X2=7.855 $Y2=0.81
r68 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.545
+ $Y=0.595 $X2=3.685 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2_4%A_937_119# 1 2 9 12 16 17 19
r39 19 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.925 $Y=0.765
+ $X2=6.925 $Y2=0.855
r40 16 17 10.1916 $w=1.83e-07 $l=1.7e-07 $layer=LI1_cond $X=5.495 $Y=0.847
+ $X2=5.665 $Y2=0.847
r41 12 14 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.825 $Y=0.75
+ $X2=4.825 $Y2=0.84
r42 9 21 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.76 $Y=0.855
+ $X2=6.925 $Y2=0.855
r43 9 17 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=6.76 $Y=0.855
+ $X2=5.665 $Y2=0.855
r44 8 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.99 $Y=0.84
+ $X2=4.825 $Y2=0.84
r45 8 16 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=4.99 $Y=0.84
+ $X2=5.495 $Y2=0.84
r46 2 19 182 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_NDIFF $count=1 $X=6.785
+ $Y=0.37 $X2=6.925 $Y2=0.765
r47 1 12 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=4.685
+ $Y=0.595 $X2=4.825 $Y2=0.75
.ends


* File: sky130_fd_sc_ms__edfxbp_1.pex.spice
* Created: Wed Sep  2 12:07:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__EDFXBP_1%D 2 5 9 11 12 16 17 20
c40 20 0 4.29314e-20 $X=0.59 $Y=1.825
r41 20 22 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.825
+ $X2=0.585 $Y2=1.99
r42 20 21 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.825 $X2=0.59 $Y2=1.825
r43 16 18 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.145
+ $X2=0.585 $Y2=0.98
r44 16 17 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.145 $X2=0.59 $Y2=1.145
r45 12 21 4.49734 $w=4.08e-07 $l=1.6e-07 $layer=LI1_cond $X=0.63 $Y=1.665
+ $X2=0.63 $Y2=1.825
r46 11 12 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.63 $Y=1.295
+ $X2=0.63 $Y2=1.665
r47 11 17 4.21625 $w=4.08e-07 $l=1.5e-07 $layer=LI1_cond $X=0.63 $Y=1.295
+ $X2=0.63 $Y2=1.145
r48 9 18 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.65 $Y=0.58 $X2=0.65
+ $Y2=0.98
r49 5 22 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=0.505 $Y=2.75
+ $X2=0.505 $Y2=1.99
r50 2 20 0.848592 $w=3.4e-07 $l=5e-09 $layer=POLY_cond $X=0.585 $Y=1.82
+ $X2=0.585 $Y2=1.825
r51 1 16 0.848592 $w=3.4e-07 $l=5e-09 $layer=POLY_cond $X=0.585 $Y=1.15
+ $X2=0.585 $Y2=1.145
r52 1 2 113.711 $w=3.4e-07 $l=6.7e-07 $layer=POLY_cond $X=0.585 $Y=1.15
+ $X2=0.585 $Y2=1.82
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXBP_1%A_161_446# 1 2 7 9 13 23 24 25 26 27 28 31
+ 35 37 41 42 44
c109 41 0 1.52853e-19 $X=2.5 $Y=1.145
c110 28 0 4.29314e-20 $X=1.335 $Y=2.035
r111 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.5
+ $Y=1.145 $X2=2.5 $Y2=1.145
r112 39 41 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=2.5 $Y=1.95
+ $X2=2.5 $Y2=1.145
r113 38 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.885 $Y=2.035
+ $X2=1.8 $Y2=2.035
r114 37 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.335 $Y=2.035
+ $X2=2.5 $Y2=1.95
r115 37 38 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.335 $Y=2.035
+ $X2=1.885 $Y2=2.035
r116 33 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.8 $Y=2.12 $X2=1.8
+ $Y2=2.035
r117 33 35 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.8 $Y=2.12
+ $X2=1.8 $Y2=2.505
r118 29 31 15.311 $w=3.48e-07 $l=4.65e-07 $layer=LI1_cond $X=1.825 $Y=1.11
+ $X2=1.825 $Y2=0.645
r119 27 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.715 $Y=2.035
+ $X2=1.8 $Y2=2.035
r120 27 28 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.715 $Y=2.035
+ $X2=1.335 $Y2=2.035
r121 25 29 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=1.65 $Y=1.195
+ $X2=1.825 $Y2=1.11
r122 25 26 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.65 $Y=1.195
+ $X2=1.335 $Y2=1.195
r123 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.17
+ $Y=1.615 $X2=1.17 $Y2=1.615
r124 21 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.17 $Y=1.95
+ $X2=1.335 $Y2=2.035
r125 21 23 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.17 $Y=1.95
+ $X2=1.17 $Y2=1.615
r126 20 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.17 $Y=1.28
+ $X2=1.335 $Y2=1.195
r127 20 23 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.17 $Y=1.28
+ $X2=1.17 $Y2=1.615
r128 19 42 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.5 $Y=0.98
+ $X2=2.5 $Y2=1.145
r129 17 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.17 $Y=1.955
+ $X2=1.17 $Y2=1.615
r130 13 19 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.56 $Y=0.58 $X2=2.56
+ $Y2=0.98
r131 7 17 57.1336 $w=2.32e-07 $l=5.45436e-07 $layer=POLY_cond $X=0.895 $Y=2.38
+ $X2=1.17 $Y2=1.955
r132 7 9 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=0.895 $Y=2.38
+ $X2=0.895 $Y2=2.75
r133 2 35 600 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=1 $X=1.655
+ $Y=2.3 $X2=1.8 $Y2=2.505
r134 1 31 182 $w=1.7e-07 $l=3.43875e-07 $layer=licon1_NDIFF $count=1 $X=1.67
+ $Y=0.37 $X2=1.825 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXBP_1%DE 1 3 4 5 8 12 14 16 17 20 21 23 25 30 33
+ 35
c87 23 0 9.594e-20 $X=2.705 $Y=2.73
c88 17 0 2.45649e-19 $X=2.44 $Y=1.965
c89 8 0 1.52853e-19 $X=1.975 $Y=0.94
r90 36 37 32.9693 $w=5.4e-07 $l=7.5e-08 $layer=POLY_cond $X=1.845 $Y=1.965
+ $X2=1.845 $Y2=2.04
r91 33 36 34.6778 $w=5.4e-07 $l=3.5e-07 $layer=POLY_cond $X=1.845 $Y=1.615
+ $X2=1.845 $Y2=1.965
r92 33 35 47.7034 $w=5.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.615
+ $X2=1.845 $Y2=1.45
r93 30 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.74
+ $Y=1.615 $X2=1.74 $Y2=1.615
r94 21 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.705 $Y=2.305
+ $X2=2.515 $Y2=2.305
r95 21 23 136.048 $w=1.8e-07 $l=3.5e-07 $layer=POLY_cond $X=2.705 $Y=2.38
+ $X2=2.705 $Y2=2.73
r96 20 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.515 $Y=2.23
+ $X2=2.515 $Y2=2.305
r97 19 20 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.515 $Y=2.04
+ $X2=2.515 $Y2=2.23
r98 18 36 33.3633 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.115 $Y=1.965
+ $X2=1.845 $Y2=1.965
r99 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.44 $Y=1.965
+ $X2=2.515 $Y2=2.04
r100 17 18 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=2.44 $Y=1.965
+ $X2=2.115 $Y2=1.965
r101 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.05 $Y=0.865
+ $X2=2.05 $Y2=0.58
r102 12 37 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=2.025 $Y=2.62
+ $X2=2.025 $Y2=2.04
r103 9 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.725 $Y=0.94
+ $X2=1.65 $Y2=0.94
r104 8 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.975 $Y=0.94
+ $X2=2.05 $Y2=0.865
r105 8 9 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.975 $Y=0.94
+ $X2=1.725 $Y2=0.94
r106 6 25 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.65 $Y=1.015
+ $X2=1.65 $Y2=0.94
r107 6 35 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.65 $Y=1.015
+ $X2=1.65 $Y2=1.45
r108 4 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.575 $Y=0.94
+ $X2=1.65 $Y2=0.94
r109 4 5 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=1.575 $Y=0.94
+ $X2=1.115 $Y2=0.94
r110 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.04 $Y=0.865
+ $X2=1.115 $Y2=0.94
r111 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.04 $Y=0.865 $X2=1.04
+ $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXBP_1%A_575_48# 1 2 9 13 17 21 25 29 33 40 42 43
+ 45 46 48 49 54 55 56 62 67 68 70 72 74 84
c230 72 0 1.37757e-19 $X=3.04 $Y=1.99
c231 68 0 1.15042e-19 $X=3.04 $Y=1.145
c232 55 0 2.25169e-19 $X=12.095 $Y=1.665
c233 49 0 7.45843e-20 $X=13.865 $Y=1.485
c234 33 0 7.24209e-20 $X=12.155 $Y=1.922
r235 73 74 2.31731 $w=3.12e-07 $l=1.5e-08 $layer=POLY_cond $X=11.435 $Y=1.89
+ $X2=11.45 $Y2=1.89
r236 70 72 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.04 $Y=1.825
+ $X2=3.04 $Y2=1.99
r237 67 70 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=3.04 $Y=1.145
+ $X2=3.04 $Y2=1.825
r238 67 68 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.04
+ $Y=1.145 $X2=3.04 $Y2=1.145
r239 63 84 40.1609 $w=3.28e-07 $l=1.15e-06 $layer=LI1_cond $X=12.32 $Y=1.665
+ $X2=12.32 $Y2=0.515
r240 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=1.665
+ $X2=12.24 $Y2=1.665
r241 59 68 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=3.04 $Y=1.665
+ $X2=3.04 $Y2=1.145
r242 59 70 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.04
+ $Y=1.825 $X2=3.04 $Y2=1.825
r243 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.665
+ $X2=3.12 $Y2=1.665
r244 56 58 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=1.665
+ $X2=3.12 $Y2=1.665
r245 55 62 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.095 $Y=1.665
+ $X2=12.24 $Y2=1.665
r246 55 56 10.9282 $w=1.4e-07 $l=8.83e-06 $layer=MET1_cond $X=12.095 $Y=1.665
+ $X2=3.265 $Y2=1.665
r247 52 63 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=12.32 $Y=1.725
+ $X2=12.32 $Y2=1.665
r248 52 54 6.62588 $w=2.9e-07 $l=1.65e-07 $layer=LI1_cond $X=12.32 $Y=1.725
+ $X2=12.155 $Y2=1.725
r249 51 84 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=12.32 $Y=0.425
+ $X2=12.32 $Y2=0.515
r250 49 78 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.865 $Y=1.485
+ $X2=13.865 $Y2=1.65
r251 49 77 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.865 $Y=1.485
+ $X2=13.865 $Y2=1.32
r252 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.865
+ $Y=1.485 $X2=13.865 $Y2=1.485
r253 46 48 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.435 $Y=1.485
+ $X2=13.865 $Y2=1.485
r254 45 46 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=13.35 $Y=1.32
+ $X2=13.435 $Y2=1.485
r255 44 45 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=13.35 $Y=0.425
+ $X2=13.35 $Y2=1.32
r256 43 51 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.485 $Y=0.34
+ $X2=12.32 $Y2=0.425
r257 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.265 $Y=0.34
+ $X2=13.35 $Y2=0.425
r258 42 43 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=13.265 $Y=0.34
+ $X2=12.485 $Y2=0.34
r259 38 54 6.62588 $w=2.9e-07 $l=5.85064e-07 $layer=LI1_cond $X=12.575 $Y=2.12
+ $X2=12.155 $Y2=1.725
r260 38 40 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=12.575 $Y=2.12
+ $X2=12.575 $Y2=2.68
r261 36 74 42.484 $w=3.12e-07 $l=2.75e-07 $layer=POLY_cond $X=11.725 $Y=1.89
+ $X2=11.45 $Y2=1.89
r262 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.725
+ $Y=1.89 $X2=11.725 $Y2=1.89
r263 33 54 0.257366 $w=3.95e-07 $l=1.97e-07 $layer=LI1_cond $X=12.155 $Y=1.922
+ $X2=12.155 $Y2=1.725
r264 33 35 12.5456 $w=3.93e-07 $l=4.3e-07 $layer=LI1_cond $X=12.155 $Y=1.922
+ $X2=11.725 $Y2=1.922
r265 32 67 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.04 $Y=0.98
+ $X2=3.04 $Y2=1.145
r266 29 77 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.905 $Y=0.76
+ $X2=13.905 $Y2=1.32
r267 25 78 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=13.85 $Y=2.4
+ $X2=13.85 $Y2=1.65
r268 19 74 19.893 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.45 $Y=1.725
+ $X2=11.45 $Y2=1.89
r269 19 21 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=11.45 $Y=1.725
+ $X2=11.45 $Y2=0.8
r270 15 73 15.628 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=11.435 $Y=2.055
+ $X2=11.435 $Y2=1.89
r271 15 17 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=11.435 $Y=2.055
+ $X2=11.435 $Y2=2.425
r272 13 72 287.645 $w=1.8e-07 $l=7.4e-07 $layer=POLY_cond $X=3.095 $Y=2.73
+ $X2=3.095 $Y2=1.99
r273 9 32 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.95 $Y=0.58 $X2=2.95
+ $Y2=0.98
r274 2 54 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=12.48
+ $Y=1.825 $X2=12.615 $Y2=1.97
r275 2 40 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=12.48
+ $Y=1.825 $X2=12.615 $Y2=2.68
r276 1 84 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.18
+ $Y=0.37 $X2=12.32 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXBP_1%CLK 1 3 6 8 14
c38 14 0 5.19822e-20 $X=4.22 $Y=1.385
r39 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.22
+ $Y=1.385 $X2=4.22 $Y2=1.385
r40 12 14 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=4.105 $Y=1.385
+ $X2=4.22 $Y2=1.385
r41 10 12 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.015 $Y=1.385
+ $X2=4.105 $Y2=1.385
r42 8 15 1.60667 $w=6.68e-07 $l=9e-08 $layer=LI1_cond $X=4.05 $Y=1.295 $X2=4.05
+ $Y2=1.385
r43 4 12 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.105 $Y=1.55
+ $X2=4.105 $Y2=1.385
r44 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=4.105 $Y=1.55
+ $X2=4.105 $Y2=2.4
r45 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.015 $Y=1.22
+ $X2=4.015 $Y2=1.385
r46 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.015 $Y=1.22 $X2=4.015
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXBP_1%A_1008_74# 1 2 9 11 13 14 16 18 21 25 27 28
+ 29 34 35 38 39 42 43 44 46 48 51 55 56 58 59 62 63 66 68 69 71 72 73 81
c221 66 0 1.31135e-19 $X=6.72 $Y=1.18
c222 62 0 1.41465e-19 $X=6.19 $Y=2.215
c223 56 0 2.75085e-19 $X=11 $Y=1.635
c224 55 0 5.74077e-20 $X=11 $Y=1.635
c225 44 0 1.9677e-19 $X=7.81 $Y=0.34
c226 21 0 7.24209e-20 $X=10.955 $Y=2.425
c227 18 0 3.32586e-20 $X=9.395 $Y=1.26
r228 72 81 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.92 $Y=1.285
+ $X2=9.755 $Y2=1.285
r229 71 73 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.92 $Y=1.285
+ $X2=10.085 $Y2=1.285
r230 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.92
+ $Y=1.285 $X2=9.92 $Y2=1.285
r231 69 71 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=9.37 $Y=1.285
+ $X2=9.92 $Y2=1.285
r232 68 69 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=9.2 $Y=1.207
+ $X2=9.37 $Y2=1.207
r233 66 76 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=6.72 $Y=1.18
+ $X2=6.595 $Y2=1.18
r234 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.72
+ $Y=1.18 $X2=6.72 $Y2=1.18
r235 63 65 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=6.76 $Y=1.05
+ $X2=6.76 $Y2=1.18
r236 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.19
+ $Y=2.215 $X2=6.19 $Y2=2.215
r237 59 61 8.7403 $w=3.35e-07 $l=2.4e-07 $layer=LI1_cond $X=6.155 $Y=1.975
+ $X2=6.155 $Y2=2.215
r238 56 85 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11 $Y=1.635 $X2=11
+ $Y2=1.8
r239 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11
+ $Y=1.635 $X2=11 $Y2=1.635
r240 53 55 14.7257 $w=2.68e-07 $l=3.45e-07 $layer=LI1_cond $X=10.97 $Y=1.29
+ $X2=10.97 $Y2=1.635
r241 51 53 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=10.835 $Y=1.205
+ $X2=10.97 $Y2=1.29
r242 51 73 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=10.835 $Y=1.205
+ $X2=10.085 $Y2=1.205
r243 48 68 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=8.49 $Y=1.05
+ $X2=9.2 $Y2=1.05
r244 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.405 $Y=0.965
+ $X2=8.49 $Y2=1.05
r245 45 46 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=8.405 $Y=0.425
+ $X2=8.405 $Y2=0.965
r246 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.32 $Y=0.34
+ $X2=8.405 $Y2=0.425
r247 43 44 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.32 $Y=0.34
+ $X2=7.81 $Y2=0.34
r248 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.725 $Y=0.425
+ $X2=7.81 $Y2=0.34
r249 41 42 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=7.725 $Y=0.425
+ $X2=7.725 $Y2=0.965
r250 40 63 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.885 $Y=1.05
+ $X2=6.76 $Y2=1.05
r251 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.64 $Y=1.05
+ $X2=7.725 $Y2=0.965
r252 39 40 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=7.64 $Y=1.05
+ $X2=6.885 $Y2=1.05
r253 38 63 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=6.76 $Y=0.965
+ $X2=6.76 $Y2=1.05
r254 37 38 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=6.76 $Y=0.425
+ $X2=6.76 $Y2=0.965
r255 36 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.125 $Y=0.34
+ $X2=6.04 $Y2=0.34
r256 35 37 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.635 $Y=0.34
+ $X2=6.76 $Y2=0.425
r257 35 36 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.635 $Y=0.34
+ $X2=6.125 $Y2=0.34
r258 34 59 8.96243 $w=3.35e-07 $l=2.14942e-07 $layer=LI1_cond $X=6.04 $Y=1.81
+ $X2=6.155 $Y2=1.975
r259 33 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.04 $Y=0.425
+ $X2=6.04 $Y2=0.34
r260 33 34 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=6.04 $Y=0.425
+ $X2=6.04 $Y2=1.81
r261 29 59 0.808037 $w=3.3e-07 $l=2e-07 $layer=LI1_cond $X=5.955 $Y=1.975
+ $X2=6.155 $Y2=1.975
r262 29 31 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=5.955 $Y=1.975
+ $X2=5.72 $Y2=1.975
r263 27 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.955 $Y=0.34
+ $X2=6.04 $Y2=0.34
r264 27 28 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.955 $Y=0.34
+ $X2=5.345 $Y2=0.34
r265 23 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.22 $Y=0.425
+ $X2=5.345 $Y2=0.34
r266 23 25 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=5.22 $Y=0.425
+ $X2=5.22 $Y2=0.515
r267 21 85 242.944 $w=1.8e-07 $l=6.25e-07 $layer=POLY_cond $X=10.955 $Y=2.425
+ $X2=10.955 $Y2=1.8
r268 18 81 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=9.395 $Y=1.26
+ $X2=9.755 $Y2=1.26
r269 14 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.32 $Y=1.185
+ $X2=9.395 $Y2=1.26
r270 14 16 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=9.32 $Y=1.185
+ $X2=9.32 $Y2=0.74
r271 11 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.595 $Y=1.015
+ $X2=6.595 $Y2=1.18
r272 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.595 $Y=1.015
+ $X2=6.595 $Y2=0.695
r273 7 62 76.2055 $w=2.53e-07 $l=4.80833e-07 $layer=POLY_cond $X=6.59 $Y=2.405
+ $X2=6.19 $Y2=2.227
r274 7 9 134.105 $w=1.8e-07 $l=3.45e-07 $layer=POLY_cond $X=6.59 $Y=2.405
+ $X2=6.59 $Y2=2.75
r275 2 31 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.585
+ $Y=1.83 $X2=5.72 $Y2=1.975
r276 1 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.04
+ $Y=0.37 $X2=5.18 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXBP_1%A_818_74# 1 2 9 11 13 15 16 20 22 28 32 36
+ 37 38 40 41 42 46 48 53 55 56 57 58 61 62 63 66 70 75 77 79 84 85 89 94 96
c227 84 0 3.39525e-20 $X=10.46 $Y=1.625
c228 79 0 1.50728e-19 $X=8.28 $Y=2.63
c229 77 0 1.41465e-19 $X=7.235 $Y=2.23
c230 36 0 1.59075e-19 $X=10.985 $Y=1.185
c231 32 0 5.74077e-20 $X=10.385 $Y=2.46
c232 22 0 1.37651e-20 $X=6.595 $Y=1.68
r233 89 90 33.431 $w=4.05e-07 $l=7.5e-08 $layer=POLY_cond $X=4.837 $Y=1.68
+ $X2=4.837 $Y2=1.605
r234 85 97 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.46 $Y=1.625
+ $X2=10.46 $Y2=1.79
r235 85 96 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.46 $Y=1.625
+ $X2=10.46 $Y2=1.46
r236 84 87 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=10.46 $Y=1.625
+ $X2=10.46 $Y2=1.705
r237 84 85 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.46
+ $Y=1.625 $X2=10.46 $Y2=1.625
r238 79 81 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=8.28 $Y=2.63
+ $X2=8.28 $Y2=2.84
r239 75 94 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.055 $Y=2.215
+ $X2=7.055 $Y2=2.38
r240 74 77 6.91466 $w=2.98e-07 $l=1.8e-07 $layer=LI1_cond $X=7.055 $Y=2.23
+ $X2=7.235 $Y2=2.23
r241 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.055
+ $Y=2.215 $X2=7.055 $Y2=2.215
r242 71 89 40.51 $w=4.05e-07 $l=2.95e-07 $layer=POLY_cond $X=4.837 $Y=1.975
+ $X2=4.837 $Y2=1.68
r243 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.8
+ $Y=1.975 $X2=4.8 $Y2=1.975
r244 68 70 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.64 $Y=1.975
+ $X2=4.8 $Y2=1.975
r245 62 87 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.295 $Y=1.705
+ $X2=10.46 $Y2=1.705
r246 62 63 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=10.295 $Y=1.705
+ $X2=9.405 $Y2=1.705
r247 60 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.32 $Y=1.79
+ $X2=9.405 $Y2=1.705
r248 60 61 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=9.32 $Y=1.79
+ $X2=9.32 $Y2=2.755
r249 59 81 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.365 $Y=2.84
+ $X2=8.28 $Y2=2.84
r250 58 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.235 $Y=2.84
+ $X2=9.32 $Y2=2.755
r251 58 59 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=9.235 $Y=2.84
+ $X2=8.365 $Y2=2.84
r252 56 79 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.195 $Y=2.63
+ $X2=8.28 $Y2=2.63
r253 56 57 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=8.195 $Y=2.63
+ $X2=7.32 $Y2=2.63
r254 55 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.235 $Y=2.545
+ $X2=7.32 $Y2=2.63
r255 54 77 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=7.235 $Y=2.38
+ $X2=7.235 $Y2=2.23
r256 54 55 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.235 $Y=2.38
+ $X2=7.235 $Y2=2.545
r257 53 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.64 $Y=1.81
+ $X2=4.64 $Y2=1.975
r258 52 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.64 $Y=1.01
+ $X2=4.64 $Y2=0.925
r259 52 53 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=4.64 $Y=1.01 $X2=4.64
+ $Y2=1.81
r260 48 68 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.555 $Y=1.975
+ $X2=4.64 $Y2=1.975
r261 48 50 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=4.555 $Y=1.975
+ $X2=4.33 $Y2=1.975
r262 44 66 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=4.23 $Y=0.925
+ $X2=4.64 $Y2=0.925
r263 44 46 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.23 $Y=0.84
+ $X2=4.23 $Y2=0.515
r264 38 40 99.6133 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=11.06 $Y=1.11
+ $X2=11.06 $Y2=0.8
r265 36 38 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.985 $Y=1.185
+ $X2=11.06 $Y2=1.11
r266 36 37 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=10.985 $Y=1.185
+ $X2=10.625 $Y2=1.185
r267 34 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.55 $Y=1.26
+ $X2=10.625 $Y2=1.185
r268 34 96 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=10.55 $Y=1.26
+ $X2=10.55 $Y2=1.46
r269 32 97 260.435 $w=1.8e-07 $l=6.7e-07 $layer=POLY_cond $X=10.385 $Y=2.46
+ $X2=10.385 $Y2=1.79
r270 28 94 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=7.04 $Y=2.75
+ $X2=7.04 $Y2=2.38
r271 24 75 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=7.055 $Y=2.015
+ $X2=7.055 $Y2=2.215
r272 23 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.99 $Y=1.68
+ $X2=5.915 $Y2=1.68
r273 22 24 108.771 $w=2.12e-07 $l=5.44702e-07 $layer=POLY_cond $X=6.595 $Y=1.68
+ $X2=7.055 $Y2=1.865
r274 22 23 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=6.595 $Y=1.68
+ $X2=5.99 $Y2=1.68
r275 18 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.915 $Y=1.605
+ $X2=5.915 $Y2=1.68
r276 18 20 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=5.915 $Y=1.605
+ $X2=5.915 $Y2=0.695
r277 17 41 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.585 $Y=1.68
+ $X2=5.495 $Y2=1.68
r278 16 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.84 $Y=1.68
+ $X2=5.915 $Y2=1.68
r279 16 17 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=5.84 $Y=1.68
+ $X2=5.585 $Y2=1.68
r280 13 41 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=5.495 $Y=1.755
+ $X2=5.495 $Y2=1.68
r281 13 15 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=5.495 $Y=1.755
+ $X2=5.495 $Y2=2.39
r282 12 89 26.1659 $w=1.5e-07 $l=2.03e-07 $layer=POLY_cond $X=5.04 $Y=1.68
+ $X2=4.837 $Y2=1.68
r283 11 41 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.405 $Y=1.68
+ $X2=5.495 $Y2=1.68
r284 11 12 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=5.405 $Y=1.68
+ $X2=5.04 $Y2=1.68
r285 9 90 443.543 $w=1.5e-07 $l=8.65e-07 $layer=POLY_cond $X=4.965 $Y=0.74
+ $X2=4.965 $Y2=1.605
r286 2 50 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=4.195
+ $Y=1.84 $X2=4.33 $Y2=2.02
r287 1 46 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.09
+ $Y=0.37 $X2=4.23 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXBP_1%A_1419_71# 1 2 9 13 17 19 21 23 24 28 30 32
+ 37 39 40 43 45 46 49
c135 49 0 1.50728e-19 $X=8.865 $Y=2.42
c136 45 0 1.30788e-19 $X=7.535 $Y=1.437
c137 30 0 3.32586e-20 $X=8.7 $Y=1.39
c138 19 0 3.39525e-20 $X=9.875 $Y=1.81
c139 9 0 1.9677e-19 $X=7.17 $Y=0.695
r140 50 58 12.9189 $w=3.35e-07 $l=7.5e-08 $layer=POLY_cond $X=8.867 $Y=1.885
+ $X2=8.867 $Y2=1.81
r141 49 50 92.1545 $w=3.35e-07 $l=5.35e-07 $layer=POLY_cond $X=8.867 $Y=2.42
+ $X2=8.867 $Y2=1.885
r142 48 49 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.865
+ $Y=2.42 $X2=8.865 $Y2=2.42
r143 42 45 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=7.37 $Y=1.437
+ $X2=7.535 $Y2=1.437
r144 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.37
+ $Y=1.435 $X2=7.37 $Y2=1.435
r145 40 58 12.0576 $w=3.35e-07 $l=7e-08 $layer=POLY_cond $X=8.867 $Y=1.74
+ $X2=8.867 $Y2=1.81
r146 40 57 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=8.867 $Y=1.74
+ $X2=8.867 $Y2=1.575
r147 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.865
+ $Y=1.74 $X2=8.865 $Y2=1.74
r148 37 48 3.2138 $w=3.3e-07 $l=2.3e-07 $layer=LI1_cond $X=8.865 $Y=2.125
+ $X2=8.865 $Y2=2.355
r149 37 39 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=8.865 $Y=2.125
+ $X2=8.865 $Y2=1.74
r150 36 39 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=8.865 $Y=1.475
+ $X2=8.865 $Y2=1.74
r151 32 48 3.77273 $w=2.5e-07 $l=2.11069e-07 $layer=LI1_cond $X=8.7 $Y=2.25
+ $X2=8.865 $Y2=2.355
r152 32 34 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=8.7 $Y=2.25
+ $X2=8.395 $Y2=2.25
r153 31 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.15 $Y=1.39
+ $X2=8.065 $Y2=1.39
r154 30 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.7 $Y=1.39
+ $X2=8.865 $Y2=1.475
r155 30 31 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=8.7 $Y=1.39
+ $X2=8.15 $Y2=1.39
r156 26 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.065 $Y=1.305
+ $X2=8.065 $Y2=1.39
r157 26 28 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=8.065 $Y=1.305
+ $X2=8.065 $Y2=0.81
r158 24 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.98 $Y=1.39
+ $X2=8.065 $Y2=1.39
r159 24 45 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=7.98 $Y=1.39
+ $X2=7.535 $Y2=1.39
r160 21 23 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.965 $Y=1.885
+ $X2=9.965 $Y2=2.46
r161 20 58 21.5811 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=9.035 $Y=1.81
+ $X2=8.867 $Y2=1.81
r162 19 21 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=9.875 $Y=1.81
+ $X2=9.965 $Y2=1.885
r163 19 20 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=9.875 $Y=1.81
+ $X2=9.035 $Y2=1.81
r164 17 57 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=8.96 $Y=0.74
+ $X2=8.96 $Y2=1.575
r165 11 43 30.0208 $w=2.89e-07 $l=2.80936e-07 $layer=POLY_cond $X=7.55 $Y=1.625
+ $X2=7.37 $Y2=1.42
r166 11 13 437.298 $w=1.8e-07 $l=1.125e-06 $layer=POLY_cond $X=7.55 $Y=1.625
+ $X2=7.55 $Y2=2.75
r167 7 43 33.3564 $w=2.89e-07 $l=2.88141e-07 $layer=POLY_cond $X=7.17 $Y=1.215
+ $X2=7.37 $Y2=1.42
r168 7 9 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=7.17 $Y=1.215
+ $X2=7.17 $Y2=0.695
r169 2 34 600 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=8.26
+ $Y=2.12 $X2=8.395 $Y2=2.29
r170 1 28 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=7.925
+ $Y=0.37 $X2=8.065 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXBP_1%A_1198_97# 1 2 7 9 14 18 22 25 27 34 35 36
+ 39
r105 35 40 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.095 $Y=1.79
+ $X2=8.095 $Y2=1.955
r106 35 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.095 $Y=1.79
+ $X2=8.095 $Y2=1.625
r107 34 36 8.46729 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=8.095 $Y=1.8
+ $X2=7.93 $Y2=1.8
r108 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.095
+ $Y=1.79 $X2=8.095 $Y2=1.79
r109 28 29 11.9654 $w=2.6e-07 $l=2.55e-07 $layer=LI1_cond $X=6.38 $Y=1.685
+ $X2=6.635 $Y2=1.685
r110 27 29 5.4494 $w=2.6e-07 $l=1.77482e-07 $layer=LI1_cond $X=6.72 $Y=1.825
+ $X2=6.635 $Y2=1.685
r111 27 36 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=6.72 $Y=1.825
+ $X2=7.93 $Y2=1.825
r112 25 32 5.95122 $w=3.69e-07 $l=2.91419e-07 $layer=LI1_cond $X=6.635 $Y=2.55
+ $X2=6.815 $Y2=2.765
r113 24 29 3.22376 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=6.635 $Y=1.91
+ $X2=6.635 $Y2=1.685
r114 24 25 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=6.635 $Y=1.91
+ $X2=6.635 $Y2=2.55
r115 20 28 3.22376 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.38 $Y=1.515
+ $X2=6.38 $Y2=1.685
r116 20 22 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=6.38 $Y=1.515
+ $X2=6.38 $Y2=0.76
r117 16 18 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=7.85 $Y=1.16
+ $X2=8.005 $Y2=1.16
r118 14 40 227.395 $w=1.8e-07 $l=5.85e-07 $layer=POLY_cond $X=8.17 $Y=2.54
+ $X2=8.17 $Y2=1.955
r119 10 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.005 $Y=1.235
+ $X2=8.005 $Y2=1.16
r120 10 39 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=8.005 $Y=1.235
+ $X2=8.005 $Y2=1.625
r121 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.85 $Y=1.085
+ $X2=7.85 $Y2=1.16
r122 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=7.85 $Y=1.085
+ $X2=7.85 $Y2=0.69
r123 2 32 600 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_PDIFF $count=1 $X=6.68
+ $Y=2.54 $X2=6.815 $Y2=2.765
r124 1 22 182 $w=1.7e-07 $l=5.09264e-07 $layer=licon1_NDIFF $count=1 $X=5.99
+ $Y=0.485 $X2=6.38 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXBP_1%A_1879_74# 1 2 9 11 13 14 15 16 18 21 24 26
+ 32 34 36 39 41 44 49
c126 49 0 1.03676e-19 $X=11.36 $Y=1.32
c127 26 0 1.71408e-19 $X=11.275 $Y=0.785
r128 51 52 31.363 $w=4.38e-07 $l=2.85e-07 $layer=POLY_cond $X=12.105 $Y=1.45
+ $X2=12.39 $Y2=1.45
r129 45 51 22.5594 $w=4.38e-07 $l=2.05e-07 $layer=POLY_cond $X=11.9 $Y=1.45
+ $X2=12.105 $Y2=1.45
r130 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.9
+ $Y=1.32 $X2=11.9 $Y2=1.32
r131 42 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.445 $Y=1.32
+ $X2=11.36 $Y2=1.32
r132 42 44 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=11.445 $Y=1.32
+ $X2=11.9 $Y2=1.32
r133 40 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.36 $Y=1.485
+ $X2=11.36 $Y2=1.32
r134 40 41 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=11.36 $Y=1.485
+ $X2=11.36 $Y2=1.985
r135 39 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.36 $Y=1.155
+ $X2=11.36 $Y2=1.32
r136 38 39 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=11.36 $Y=0.95
+ $X2=11.36 $Y2=1.155
r137 37 48 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.775 $Y=2.07
+ $X2=10.61 $Y2=2.07
r138 36 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.275 $Y=2.07
+ $X2=11.36 $Y2=1.985
r139 36 37 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=11.275 $Y=2.07
+ $X2=10.775 $Y2=2.07
r140 32 48 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.61 $Y=2.155
+ $X2=10.61 $Y2=2.07
r141 32 34 23.0489 $w=3.28e-07 $l=6.6e-07 $layer=LI1_cond $X=10.61 $Y=2.155
+ $X2=10.61 $Y2=2.815
r142 28 31 42.6055 $w=3.28e-07 $l=1.22e-06 $layer=LI1_cond $X=9.625 $Y=0.785
+ $X2=10.845 $Y2=0.785
r143 26 38 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.275 $Y=0.785
+ $X2=11.36 $Y2=0.95
r144 26 31 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.275 $Y=0.785
+ $X2=10.845 $Y2=0.785
r145 23 24 47.4664 $w=3.1e-07 $l=2.55e-07 $layer=POLY_cond $X=13.145 $Y=1.36
+ $X2=13.4 $Y2=1.36
r146 19 24 15.4789 $w=1.8e-07 $l=1.55e-07 $layer=POLY_cond $X=13.4 $Y=1.515
+ $X2=13.4 $Y2=1.36
r147 19 21 344.008 $w=1.8e-07 $l=8.85e-07 $layer=POLY_cond $X=13.4 $Y=1.515
+ $X2=13.4 $Y2=2.4
r148 16 23 19.7411 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=13.145 $Y=1.205
+ $X2=13.145 $Y2=1.36
r149 16 18 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=13.145 $Y=1.205
+ $X2=13.145 $Y2=0.76
r150 15 52 14.0844 $w=4.38e-07 $l=1.27279e-07 $layer=POLY_cond $X=12.48 $Y=1.36
+ $X2=12.39 $Y2=1.45
r151 14 23 13.9607 $w=3.1e-07 $l=7.5e-08 $layer=POLY_cond $X=13.07 $Y=1.36
+ $X2=13.145 $Y2=1.36
r152 14 15 109.824 $w=3.1e-07 $l=5.9e-07 $layer=POLY_cond $X=13.07 $Y=1.36
+ $X2=12.48 $Y2=1.36
r153 11 52 23.6381 $w=1.8e-07 $l=2.95e-07 $layer=POLY_cond $X=12.39 $Y=1.745
+ $X2=12.39 $Y2=1.45
r154 11 13 155.311 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=12.39 $Y=1.745
+ $X2=12.39 $Y2=2.325
r155 7 51 28.0956 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=12.105 $Y=1.155
+ $X2=12.105 $Y2=1.45
r156 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=12.105 $Y=1.155
+ $X2=12.105 $Y2=0.69
r157 2 48 300 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=2 $X=10.475
+ $Y=1.96 $X2=10.61 $Y2=2.125
r158 2 34 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=10.475
+ $Y=1.96 $X2=10.61 $Y2=2.815
r159 1 31 91 $w=1.7e-07 $l=1.64446e-06 $layer=licon1_NDIFF $count=2 $X=9.395
+ $Y=0.37 $X2=10.845 $Y2=0.785
r160 1 28 91 $w=1.7e-07 $l=5.17373e-07 $layer=licon1_NDIFF $count=2 $X=9.395
+ $Y=0.37 $X2=9.625 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXBP_1%A_27_74# 1 2 3 4 5 6 20 23 25 28 29 30 32
+ 33 34 37 40 41 44 45 47 49 52 53 55 60 62 66 68 73
c175 68 0 2.33697e-19 $X=3.35 $Y=2.385
c176 34 0 1.30607e-19 $X=2.225 $Y=2.375
r177 64 66 7.6705 $w=4.58e-07 $l=2.95e-07 $layer=LI1_cond $X=3.165 $Y=0.58
+ $X2=3.46 $Y2=0.58
r178 57 60 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.17 $Y=0.585
+ $X2=0.435 $Y2=0.585
r179 53 55 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=5.775 $Y=2.975
+ $X2=6.28 $Y2=2.975
r180 52 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.69 $Y=2.89
+ $X2=5.775 $Y2=2.975
r181 51 52 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=5.69 $Y=2.48
+ $X2=5.69 $Y2=2.89
r182 47 69 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=5.66 $Y=1.385
+ $X2=5.3 $Y2=1.385
r183 47 49 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=5.66 $Y=1.3
+ $X2=5.66 $Y2=0.76
r184 46 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.385 $Y=2.395
+ $X2=5.3 $Y2=2.395
r185 45 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.605 $Y=2.395
+ $X2=5.69 $Y2=2.48
r186 45 46 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.605 $Y=2.395
+ $X2=5.385 $Y2=2.395
r187 44 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=2.31 $X2=5.3
+ $Y2=2.395
r188 43 69 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=1.47 $X2=5.3
+ $Y2=1.385
r189 43 44 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=5.3 $Y=1.47 $X2=5.3
+ $Y2=2.31
r190 42 68 4.69131 $w=1.7e-07 $l=1.99937e-07 $layer=LI1_cond $X=3.545 $Y=2.395
+ $X2=3.35 $Y2=2.385
r191 41 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.215 $Y=2.395
+ $X2=5.3 $Y2=2.395
r192 41 42 108.952 $w=1.68e-07 $l=1.67e-06 $layer=LI1_cond $X=5.215 $Y=2.395
+ $X2=3.545 $Y2=2.395
r193 40 68 1.68048 $w=1.7e-07 $l=1.50167e-07 $layer=LI1_cond $X=3.46 $Y=2.29
+ $X2=3.35 $Y2=2.385
r194 39 66 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.46 $Y=0.81 $X2=3.46
+ $Y2=0.58
r195 39 40 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=3.46 $Y=0.81
+ $X2=3.46 $Y2=2.29
r196 35 68 1.68048 $w=3.9e-07 $l=9.5e-08 $layer=LI1_cond $X=3.35 $Y=2.48
+ $X2=3.35 $Y2=2.385
r197 35 37 7.38745 $w=3.88e-07 $l=2.5e-07 $layer=LI1_cond $X=3.35 $Y=2.48
+ $X2=3.35 $Y2=2.73
r198 33 68 4.69131 $w=1.7e-07 $l=1.99937e-07 $layer=LI1_cond $X=3.155 $Y=2.375
+ $X2=3.35 $Y2=2.385
r199 33 34 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.155 $Y=2.375
+ $X2=2.225 $Y2=2.375
r200 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.14 $Y=2.46
+ $X2=2.225 $Y2=2.375
r201 31 32 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.14 $Y=2.46
+ $X2=2.14 $Y2=2.905
r202 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.055 $Y=2.99
+ $X2=2.14 $Y2=2.905
r203 29 30 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.055 $Y=2.99
+ $X2=1.545 $Y2=2.99
r204 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.46 $Y=2.905
+ $X2=1.545 $Y2=2.99
r205 27 28 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.46 $Y=2.46
+ $X2=1.46 $Y2=2.905
r206 26 62 2.98021 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.445 $Y=2.375
+ $X2=0.265 $Y2=2.375
r207 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.375 $Y=2.375
+ $X2=1.46 $Y2=2.46
r208 25 26 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=1.375 $Y=2.375
+ $X2=0.445 $Y2=2.375
r209 21 62 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=2.46
+ $X2=0.265 $Y2=2.375
r210 21 23 9.28357 $w=3.58e-07 $l=2.9e-07 $layer=LI1_cond $X=0.265 $Y=2.46
+ $X2=0.265 $Y2=2.75
r211 20 62 3.52026 $w=2.65e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.17 $Y=2.29
+ $X2=0.265 $Y2=2.375
r212 19 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=0.75
+ $X2=0.17 $Y2=0.585
r213 19 20 100.471 $w=1.68e-07 $l=1.54e-06 $layer=LI1_cond $X=0.17 $Y=0.75
+ $X2=0.17 $Y2=2.29
r214 6 55 600 $w=1.7e-07 $l=5.02295e-07 $layer=licon1_PDIFF $count=1 $X=6.135
+ $Y=2.54 $X2=6.28 $Y2=2.975
r215 5 37 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=3.185
+ $Y=2.52 $X2=3.32 $Y2=2.73
r216 4 23 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.28 $Y2=2.75
r217 3 49 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=5.575
+ $Y=0.485 $X2=5.7 $Y2=0.76
r218 2 64 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.025
+ $Y=0.37 $X2=3.165 $Y2=0.58
r219 1 60 182 $w=1.7e-07 $l=3.93065e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.435 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXBP_1%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 47 53
+ 57 62 63 65 66 67 69 74 89 96 104 109 116 117 120 123 126 129 132 137
r160 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r161 133 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r162 132 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r163 132 133 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r164 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r165 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r166 123 124 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r167 120 121 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r168 117 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.68 $Y2=3.33
r169 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r170 114 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.79 $Y=3.33
+ $X2=13.665 $Y2=3.33
r171 114 116 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=13.79 $Y=3.33
+ $X2=14.16 $Y2=3.33
r172 113 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r173 113 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.24 $Y2=3.33
r174 112 113 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r175 110 132 14.4958 $w=1.7e-07 $l=3.93e-07 $layer=LI1_cond $X=12.28 $Y=3.33
+ $X2=11.887 $Y2=3.33
r176 110 112 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=12.28 $Y=3.33
+ $X2=13.2 $Y2=3.33
r177 109 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.54 $Y=3.33
+ $X2=13.665 $Y2=3.33
r178 109 112 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=13.54 $Y=3.33
+ $X2=13.2 $Y2=3.33
r179 108 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r180 108 130 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=9.84 $Y2=3.33
r181 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r182 105 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.905 $Y=3.33
+ $X2=9.74 $Y2=3.33
r183 105 107 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=9.905 $Y=3.33
+ $X2=11.28 $Y2=3.33
r184 104 132 14.4958 $w=1.7e-07 $l=3.92e-07 $layer=LI1_cond $X=11.495 $Y=3.33
+ $X2=11.887 $Y2=3.33
r185 104 107 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=11.495 $Y=3.33
+ $X2=11.28 $Y2=3.33
r186 103 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r187 102 103 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r188 100 103 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r189 100 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r190 99 102 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r191 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r192 97 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=7.86 $Y2=3.33
r193 97 99 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=8.4 $Y2=3.33
r194 96 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.575 $Y=3.33
+ $X2=9.74 $Y2=3.33
r195 96 102 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=9.575 $Y=3.33
+ $X2=9.36 $Y2=3.33
r196 95 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r197 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r198 91 94 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=7.44 $Y2=3.33
r199 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r200 89 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.695 $Y=3.33
+ $X2=7.86 $Y2=3.33
r201 89 94 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.695 $Y=3.33
+ $X2=7.44 $Y2=3.33
r202 88 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r203 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r204 85 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r205 84 87 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r206 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r207 82 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r208 82 124 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r209 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r210 79 123 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.645 $Y=3.33
+ $X2=2.52 $Y2=3.33
r211 79 81 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=2.645 $Y=3.33
+ $X2=3.6 $Y2=3.33
r212 78 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r213 78 121 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r214 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r215 75 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.205 $Y=3.33
+ $X2=1.08 $Y2=3.33
r216 75 77 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.205 $Y=3.33
+ $X2=2.16 $Y2=3.33
r217 74 123 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.52 $Y2=3.33
r218 74 77 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.395 $Y=3.33
+ $X2=2.16 $Y2=3.33
r219 72 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r220 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r221 69 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=1.08 $Y2=3.33
r222 69 71 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=0.72 $Y2=3.33
r223 67 95 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=7.44 $Y2=3.33
r224 67 92 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=5.52 $Y2=3.33
r225 65 87 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.105 $Y=3.33
+ $X2=5.04 $Y2=3.33
r226 65 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.105 $Y=3.33
+ $X2=5.27 $Y2=3.33
r227 64 91 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.435 $Y=3.33
+ $X2=5.52 $Y2=3.33
r228 64 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.435 $Y=3.33
+ $X2=5.27 $Y2=3.33
r229 62 81 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.715 $Y=3.33
+ $X2=3.6 $Y2=3.33
r230 62 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.715 $Y=3.33
+ $X2=3.88 $Y2=3.33
r231 61 84 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=4.08 $Y2=3.33
r232 61 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=3.88 $Y2=3.33
r233 57 60 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=13.665 $Y=1.985
+ $X2=13.665 $Y2=2.815
r234 55 137 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.665 $Y=3.245
+ $X2=13.665 $Y2=3.33
r235 55 60 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=13.665 $Y=3.245
+ $X2=13.665 $Y2=2.815
r236 51 132 3.09511 $w=7.85e-07 $l=8.5e-08 $layer=LI1_cond $X=11.887 $Y=3.245
+ $X2=11.887 $Y2=3.33
r237 51 53 11.5037 $w=7.83e-07 $l=7.55e-07 $layer=LI1_cond $X=11.887 $Y=3.245
+ $X2=11.887 $Y2=2.49
r238 47 50 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=9.74 $Y=2.125
+ $X2=9.74 $Y2=2.815
r239 45 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.74 $Y=3.245
+ $X2=9.74 $Y2=3.33
r240 45 50 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=9.74 $Y=3.245
+ $X2=9.74 $Y2=2.815
r241 41 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.86 $Y=3.245
+ $X2=7.86 $Y2=3.33
r242 41 43 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=7.86 $Y=3.245
+ $X2=7.86 $Y2=3.05
r243 37 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.27 $Y=3.245
+ $X2=5.27 $Y2=3.33
r244 37 39 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=5.27 $Y=3.245
+ $X2=5.27 $Y2=2.77
r245 33 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.88 $Y=3.245
+ $X2=3.88 $Y2=3.33
r246 33 35 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.88 $Y=3.245
+ $X2=3.88 $Y2=2.815
r247 29 123 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=3.245
+ $X2=2.52 $Y2=3.33
r248 29 31 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=2.52 $Y=3.245
+ $X2=2.52 $Y2=2.795
r249 25 120 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.08 $Y=3.245
+ $X2=1.08 $Y2=3.33
r250 25 27 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=1.08 $Y=3.245
+ $X2=1.08 $Y2=2.805
r251 8 60 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=13.49
+ $Y=1.84 $X2=13.625 $Y2=2.815
r252 8 57 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=13.49
+ $Y=1.84 $X2=13.625 $Y2=1.985
r253 7 53 300 $w=1.7e-07 $l=7.14388e-07 $layer=licon1_PDIFF $count=2 $X=11.525
+ $Y=2.215 $X2=12.115 $Y2=2.49
r254 6 50 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=9.595
+ $Y=1.96 $X2=9.74 $Y2=2.815
r255 6 47 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=9.595
+ $Y=1.96 $X2=9.74 $Y2=2.125
r256 5 43 600 $w=1.7e-07 $l=6.10164e-07 $layer=licon1_PDIFF $count=1 $X=7.64
+ $Y=2.54 $X2=7.86 $Y2=3.05
r257 4 39 600 $w=1.7e-07 $l=1.0099e-06 $layer=licon1_PDIFF $count=1 $X=5.125
+ $Y=1.83 $X2=5.27 $Y2=2.77
r258 3 35 600 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=3.735
+ $Y=1.84 $X2=3.88 $Y2=2.815
r259 2 31 600 $w=1.7e-07 $l=6.52457e-07 $layer=licon1_PDIFF $count=1 $X=2.115
+ $Y=2.3 $X2=2.48 $Y2=2.795
r260 1 27 600 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=2.54 $X2=1.12 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXBP_1%Q 1 2 10 13 14 15 22 32
c32 32 0 7.45843e-20 $X=13.132 $Y=1.82
r33 20 22 0.222158 $w=4.13e-07 $l=8e-09 $layer=LI1_cond $X=13.132 $Y=2.027
+ $X2=13.132 $Y2=2.035
r34 14 15 10.2748 $w=4.13e-07 $l=3.7e-07 $layer=LI1_cond $X=13.132 $Y=2.405
+ $X2=13.132 $Y2=2.775
r35 13 20 1.16633 $w=4.13e-07 $l=4.2e-08 $layer=LI1_cond $X=13.132 $Y=1.985
+ $X2=13.132 $Y2=2.027
r36 13 32 8.71334 $w=4.13e-07 $l=1.65e-07 $layer=LI1_cond $X=13.132 $Y=1.985
+ $X2=13.132 $Y2=1.82
r37 13 14 9.21954 $w=4.13e-07 $l=3.32e-07 $layer=LI1_cond $X=13.132 $Y=2.073
+ $X2=13.132 $Y2=2.405
r38 13 22 1.05525 $w=4.13e-07 $l=3.8e-08 $layer=LI1_cond $X=13.132 $Y=2.073
+ $X2=13.132 $Y2=2.035
r39 12 32 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=13.01 $Y=1 $X2=13.01
+ $Y2=1.82
r40 10 12 9.33524 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=12.93 $Y=0.81
+ $X2=12.93 $Y2=1
r41 2 13 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=13.03
+ $Y=1.84 $X2=13.175 $Y2=1.985
r42 2 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=13.03
+ $Y=1.84 $X2=13.175 $Y2=2.815
r43 1 10 182 $w=1.7e-07 $l=4.87134e-07 $layer=licon1_NDIFF $count=1 $X=12.785
+ $Y=0.39 $X2=12.93 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXBP_1%Q_N 1 2 7 9 15 16 17 28
r22 21 28 1.44055 $w=3.58e-07 $l=4.5e-08 $layer=LI1_cond $X=14.135 $Y=0.97
+ $X2=14.135 $Y2=0.925
r23 17 30 8.35096 $w=3.58e-07 $l=1.6e-07 $layer=LI1_cond $X=14.135 $Y=0.99
+ $X2=14.135 $Y2=1.15
r24 17 21 0.640246 $w=3.58e-07 $l=2e-08 $layer=LI1_cond $X=14.135 $Y=0.99
+ $X2=14.135 $Y2=0.97
r25 17 28 0.640246 $w=3.58e-07 $l=2e-08 $layer=LI1_cond $X=14.135 $Y=0.905
+ $X2=14.135 $Y2=0.925
r26 16 17 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=14.135 $Y=0.535
+ $X2=14.135 $Y2=0.905
r27 15 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=14.23 $Y=1.82
+ $X2=14.23 $Y2=1.15
r28 9 11 29.4316 $w=3.23e-07 $l=8.3e-07 $layer=LI1_cond $X=14.152 $Y=1.985
+ $X2=14.152 $Y2=2.815
r29 7 15 8.35379 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=14.152 $Y=1.982
+ $X2=14.152 $Y2=1.82
r30 7 9 0.106379 $w=3.23e-07 $l=3e-09 $layer=LI1_cond $X=14.152 $Y=1.982
+ $X2=14.152 $Y2=1.985
r31 2 11 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=13.94
+ $Y=1.84 $X2=14.075 $Y2=2.815
r32 2 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=13.94
+ $Y=1.84 $X2=14.075 $Y2=1.985
r33 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.98
+ $Y=0.39 $X2=14.12 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_MS__EDFXBP_1%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 51
+ 55 58 59 61 62 64 65 66 68 86 93 98 103 110 111 114 117 120 123 126
r153 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r154 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r155 120 121 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r156 117 118 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r157 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r158 111 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=13.68 $Y2=0
r159 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r160 108 126 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.775 $Y=0
+ $X2=13.69 $Y2=0
r161 108 110 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=13.775 $Y=0
+ $X2=14.16 $Y2=0
r162 107 127 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=13.68 $Y2=0
r163 107 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r164 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r165 104 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.985 $Y=0
+ $X2=11.82 $Y2=0
r166 104 106 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.985 $Y=0
+ $X2=12.24 $Y2=0
r167 103 126 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.605 $Y=0
+ $X2=13.69 $Y2=0
r168 103 106 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=13.605 $Y=0
+ $X2=12.24 $Y2=0
r169 102 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r170 102 121 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=8.88 $Y2=0
r171 101 102 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r172 99 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.91 $Y=0
+ $X2=8.785 $Y2=0
r173 99 101 154.62 $w=1.68e-07 $l=2.37e-06 $layer=LI1_cond $X=8.91 $Y=0
+ $X2=11.28 $Y2=0
r174 98 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.655 $Y=0
+ $X2=11.82 $Y2=0
r175 98 101 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.655 $Y=0
+ $X2=11.28 $Y2=0
r176 97 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r177 97 118 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.44
+ $Y2=0
r178 96 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r179 94 117 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.47 $Y=0
+ $X2=7.345 $Y2=0
r180 94 96 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=7.47 $Y=0 $X2=8.4
+ $Y2=0
r181 93 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.66 $Y=0
+ $X2=8.785 $Y2=0
r182 93 96 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=8.66 $Y=0 $X2=8.4
+ $Y2=0
r183 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r184 89 92 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.96 $Y2=0
r185 88 91 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=6.96
+ $Y2=0
r186 88 89 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r187 86 117 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.22 $Y=0
+ $X2=7.345 $Y2=0
r188 86 91 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.22 $Y=0 $X2=6.96
+ $Y2=0
r189 85 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r190 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r191 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r192 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r193 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r194 78 81 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r195 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r196 76 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r197 76 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r198 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r199 73 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.42 $Y=0
+ $X2=1.255 $Y2=0
r200 73 75 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.42 $Y=0 $X2=2.16
+ $Y2=0
r201 71 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r202 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r203 68 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.09 $Y=0
+ $X2=1.255 $Y2=0
r204 68 70 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.09 $Y=0 $X2=0.72
+ $Y2=0
r205 66 118 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=0
+ $X2=7.44 $Y2=0
r206 66 92 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=0 $X2=6.96
+ $Y2=0
r207 64 84 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.585 $Y=0 $X2=4.56
+ $Y2=0
r208 64 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.585 $Y=0 $X2=4.75
+ $Y2=0
r209 63 88 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.915 $Y=0
+ $X2=5.04 $Y2=0
r210 63 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.915 $Y=0 $X2=4.75
+ $Y2=0
r211 61 81 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.6
+ $Y2=0
r212 61 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.8
+ $Y2=0
r213 60 84 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=3.885 $Y=0
+ $X2=4.56 $Y2=0
r214 60 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.885 $Y=0 $X2=3.8
+ $Y2=0
r215 58 75 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=2.17 $Y=0 $X2=2.16
+ $Y2=0
r216 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.17 $Y=0 $X2=2.335
+ $Y2=0
r217 57 78 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.5 $Y=0 $X2=2.64
+ $Y2=0
r218 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.5 $Y=0 $X2=2.335
+ $Y2=0
r219 53 126 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.69 $Y=0.085
+ $X2=13.69 $Y2=0
r220 53 55 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=13.69 $Y=0.085
+ $X2=13.69 $Y2=0.535
r221 49 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.82 $Y=0.085
+ $X2=11.82 $Y2=0
r222 49 51 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.82 $Y=0.085
+ $X2=11.82 $Y2=0.515
r223 45 120 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.785 $Y=0.085
+ $X2=8.785 $Y2=0
r224 45 47 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=8.785 $Y=0.085
+ $X2=8.785 $Y2=0.595
r225 41 117 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.345 $Y=0.085
+ $X2=7.345 $Y2=0
r226 41 43 25.1233 $w=2.48e-07 $l=5.45e-07 $layer=LI1_cond $X=7.345 $Y=0.085
+ $X2=7.345 $Y2=0.63
r227 37 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.75 $Y=0.085
+ $X2=4.75 $Y2=0
r228 37 39 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.75 $Y=0.085
+ $X2=4.75 $Y2=0.55
r229 33 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.8 $Y=0.085 $X2=3.8
+ $Y2=0
r230 33 35 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.8 $Y=0.085
+ $X2=3.8 $Y2=0.505
r231 29 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.335 $Y=0.085
+ $X2=2.335 $Y2=0
r232 29 31 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.335 $Y=0.085
+ $X2=2.335 $Y2=0.58
r233 25 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.255 $Y=0.085
+ $X2=1.255 $Y2=0
r234 25 27 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.255 $Y=0.085
+ $X2=1.255 $Y2=0.58
r235 8 55 91 $w=1.7e-07 $l=5.37634e-07 $layer=licon1_NDIFF $count=2 $X=13.22
+ $Y=0.39 $X2=13.69 $Y2=0.535
r236 7 51 91 $w=1.7e-07 $l=3.30379e-07 $layer=licon1_NDIFF $count=2 $X=11.525
+ $Y=0.59 $X2=11.82 $Y2=0.515
r237 6 47 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=8.6
+ $Y=0.37 $X2=8.745 $Y2=0.595
r238 5 43 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.245
+ $Y=0.485 $X2=7.385 $Y2=0.63
r239 4 39 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=4.625
+ $Y=0.37 $X2=4.75 $Y2=0.55
r240 3 35 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.655
+ $Y=0.37 $X2=3.8 $Y2=0.505
r241 2 31 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=2.125
+ $Y=0.37 $X2=2.335 $Y2=0.58
r242 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.115
+ $Y=0.37 $X2=1.255 $Y2=0.58
.ends


* File: sky130_fd_sc_ms__dfrbp_2.pex.spice
* Created: Fri Aug 28 17:22:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DFRBP_2%D 3 7 9 10 12 13 14 18
c31 9 0 8.70277e-20 $X=0.5 $Y=0.9
r32 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.065 $X2=0.385 $Y2=1.065
r33 14 19 6.79646 $w=3.88e-07 $l=2.3e-07 $layer=LI1_cond $X=0.32 $Y=1.295
+ $X2=0.32 $Y2=1.065
r34 13 19 4.13697 $w=3.88e-07 $l=1.4e-07 $layer=LI1_cond $X=0.32 $Y=0.925
+ $X2=0.32 $Y2=1.065
r35 11 18 28.3893 $w=4.9e-07 $l=2.6e-07 $layer=POLY_cond $X=0.465 $Y=1.325
+ $X2=0.465 $Y2=1.065
r36 11 12 49.2579 $w=4.9e-07 $l=2.45e-07 $layer=POLY_cond $X=0.465 $Y=1.325
+ $X2=0.465 $Y2=1.57
r37 10 18 1.63785 $w=4.9e-07 $l=1.5e-08 $layer=POLY_cond $X=0.465 $Y=1.05
+ $X2=0.465 $Y2=1.065
r38 9 10 44.6155 $w=4.9e-07 $l=1.5e-07 $layer=POLY_cond $X=0.5 $Y=0.9 $X2=0.5
+ $Y2=1.05
r39 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.705 $Y=0.58
+ $X2=0.705 $Y2=0.9
r40 3 12 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=0.62 $Y=2.17 $X2=0.62
+ $Y2=1.57
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_2%A_298_294# 1 2 3 12 16 19 22 23 27 29 30 33
+ 36 40 42
c106 42 0 1.97119e-19 $X=4.05 $Y=1.44
c107 30 0 4.31709e-20 $X=2.435 $Y=2.03
c108 23 0 3.04161e-20 $X=1.99 $Y=1.635
c109 16 0 5.72834e-20 $X=1.595 $Y=0.965
r110 42 44 7.89247 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=4.01 $Y=1.44
+ $X2=4.01 $Y2=1.61
r111 36 40 3.32435 $w=2.82e-07 $l=1.05924e-07 $layer=LI1_cond $X=4.002 $Y=1.945
+ $X2=3.955 $Y2=2.03
r112 36 44 16.4284 $w=2.33e-07 $l=3.35e-07 $layer=LI1_cond $X=4.002 $Y=1.945
+ $X2=4.002 $Y2=1.61
r113 31 40 3.32435 $w=2.82e-07 $l=8.5e-08 $layer=LI1_cond $X=3.955 $Y=2.115
+ $X2=3.955 $Y2=2.03
r114 31 33 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=3.955 $Y=2.115
+ $X2=3.955 $Y2=2.57
r115 29 40 3.22099 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.79 $Y=2.03
+ $X2=3.955 $Y2=2.03
r116 29 30 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=3.79 $Y=2.03
+ $X2=2.435 $Y2=2.03
r117 25 30 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.31 $Y=2.03
+ $X2=2.435 $Y2=2.03
r118 25 27 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=2.31 $Y=2.115
+ $X2=2.31 $Y2=2.57
r119 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.99
+ $Y=1.635 $X2=1.99 $Y2=1.635
r120 20 25 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.99 $Y=2.03
+ $X2=2.31 $Y2=2.03
r121 20 22 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.99 $Y=1.945
+ $X2=1.99 $Y2=1.635
r122 18 23 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=1.67 $Y=1.635
+ $X2=1.99 $Y2=1.635
r123 18 19 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.67 $Y=1.635
+ $X2=1.58 $Y2=1.635
r124 14 19 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=1.595 $Y=1.47
+ $X2=1.58 $Y2=1.635
r125 14 16 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.595 $Y=1.47
+ $X2=1.595 $Y2=0.965
r126 10 19 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.58 $Y=1.8
+ $X2=1.58 $Y2=1.635
r127 10 12 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.58 $Y=1.8
+ $X2=1.58 $Y2=2.46
r128 3 33 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.82
+ $Y=2.425 $X2=3.955 $Y2=2.57
r129 2 27 600 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=2.22
+ $Y=2.425 $X2=2.35 $Y2=2.57
r130 1 42 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=3.91
+ $Y=1.16 $X2=4.05 $Y2=1.44
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_2%RESET_B 3 8 9 10 13 18 21 25 27 28 29 30 36
+ 39 42 43 47 48 52 53
c205 53 0 1.1019e-19 $X=9.705 $Y=1.615
c206 52 0 1.06861e-19 $X=9.705 $Y=1.615
c207 43 0 5.72834e-20 $X=1.115 $Y=1.615
c208 30 0 3.6858e-19 $X=2.785 $Y=1.665
c209 21 0 1.76421e-19 $X=9.77 $Y=2.155
r210 52 55 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.705 $Y=1.615
+ $X2=9.705 $Y2=1.78
r211 52 54 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.705 $Y=1.615
+ $X2=9.705 $Y2=1.45
r212 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.705
+ $Y=1.615 $X2=9.705 $Y2=1.615
r213 47 50 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.55 $Y=1.61
+ $X2=2.55 $Y2=1.775
r214 47 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.55 $Y=1.61
+ $X2=2.55 $Y2=1.445
r215 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.55
+ $Y=1.61 $X2=2.55 $Y2=1.61
r216 42 45 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.115 $Y=1.615
+ $X2=1.115 $Y2=1.78
r217 42 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.115 $Y=1.615
+ $X2=1.115 $Y2=1.45
r218 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.115
+ $Y=1.615 $X2=1.115 $Y2=1.615
r219 39 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=1.665
r220 36 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=1.665
+ $X2=9.84 $Y2=1.665
r221 32 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=1.665
+ $X2=1.2 $Y2=1.665
r222 30 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=1.665
+ $X2=2.64 $Y2=1.665
r223 29 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.695 $Y=1.665
+ $X2=9.84 $Y2=1.665
r224 29 30 8.55196 $w=1.4e-07 $l=6.91e-06 $layer=MET1_cond $X=9.695 $Y=1.665
+ $X2=2.785 $Y2=1.665
r225 28 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=1.665
+ $X2=1.2 $Y2=1.665
r226 27 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.495 $Y=1.665
+ $X2=2.64 $Y2=1.665
r227 27 28 1.42326 $w=1.4e-07 $l=1.15e-06 $layer=MET1_cond $X=2.495 $Y=1.665
+ $X2=1.345 $Y2=1.665
r228 25 54 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=9.795 $Y=0.58
+ $X2=9.795 $Y2=1.45
r229 21 55 145.766 $w=1.8e-07 $l=3.75e-07 $layer=POLY_cond $X=9.77 $Y=2.155
+ $X2=9.77 $Y2=1.78
r230 18 49 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=2.605 $Y=0.615
+ $X2=2.605 $Y2=1.445
r231 15 18 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=2.605 $Y=0.255
+ $X2=2.605 $Y2=0.615
r232 13 50 334.29 $w=1.8e-07 $l=8.6e-07 $layer=POLY_cond $X=2.575 $Y=2.635
+ $X2=2.575 $Y2=1.775
r233 9 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.53 $Y=0.18
+ $X2=2.605 $Y2=0.255
r234 9 10 712.745 $w=1.5e-07 $l=1.39e-06 $layer=POLY_cond $X=2.53 $Y=0.18
+ $X2=1.14 $Y2=0.18
r235 8 44 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=1.065 $Y=0.58
+ $X2=1.065 $Y2=1.45
r236 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.065 $Y=0.255
+ $X2=1.14 $Y2=0.18
r237 5 8 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=1.065 $Y=0.255
+ $X2=1.065 $Y2=0.58
r238 3 45 151.597 $w=1.8e-07 $l=3.9e-07 $layer=POLY_cond $X=1.07 $Y=2.17
+ $X2=1.07 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_2%A_334_119# 1 2 3 4 15 17 20 22 23 25 28 30
+ 32 34 35 37 38 39 41 43 44 45 47 48 49 51 54 56 57 60 65 70 73 77
c222 77 0 1.92736e-19 $X=3.34 $Y=1.68
c223 60 0 6.79844e-20 $X=7.795 $Y=2.09
c224 56 0 1.4118e-19 $X=7.71 $Y=1.44
c225 51 0 8.33581e-20 $X=7.3 $Y=1.355
c226 41 0 1.45428e-19 $X=3.01 $Y=1.555
c227 35 0 4.31709e-20 $X=2.155 $Y=1.1
r228 71 77 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.09 $Y=1.68
+ $X2=3.34 $Y2=1.68
r229 71 74 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=3.09 $Y=1.68 $X2=3.03
+ $Y2=1.68
r230 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.68 $X2=3.09 $Y2=1.68
r231 67 70 4.1907 $w=2.18e-07 $l=8e-08 $layer=LI1_cond $X=3.01 $Y=1.665 $X2=3.09
+ $Y2=1.665
r232 64 65 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.79 $Y=1.1
+ $X2=3.01 $Y2=1.1
r233 58 60 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=7.795 $Y=1.525
+ $X2=7.795 $Y2=2.09
r234 56 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.71 $Y=1.44
+ $X2=7.795 $Y2=1.525
r235 56 57 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.71 $Y=1.44
+ $X2=7.385 $Y2=1.44
r236 52 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.385 $Y=0.34
+ $X2=7.3 $Y2=0.34
r237 52 54 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=7.385 $Y=0.34
+ $X2=8.615 $Y2=0.34
r238 51 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.3 $Y=1.355
+ $X2=7.385 $Y2=1.44
r239 50 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.3 $Y=0.425 $X2=7.3
+ $Y2=0.34
r240 50 51 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=7.3 $Y=0.425
+ $X2=7.3 $Y2=1.355
r241 48 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.215 $Y=0.34
+ $X2=7.3 $Y2=0.34
r242 48 49 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=7.215 $Y=0.34
+ $X2=6.195 $Y2=0.34
r243 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.11 $Y=0.425
+ $X2=6.195 $Y2=0.34
r244 46 47 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.11 $Y=0.425
+ $X2=6.11 $Y2=0.66
r245 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.025 $Y=0.745
+ $X2=6.11 $Y2=0.66
r246 44 45 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=6.025 $Y=0.745
+ $X2=5.235 $Y2=0.745
r247 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.15 $Y=0.66
+ $X2=5.235 $Y2=0.745
r248 42 43 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.15 $Y=0.425
+ $X2=5.15 $Y2=0.66
r249 41 67 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.01 $Y=1.555
+ $X2=3.01 $Y2=1.665
r250 40 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.01 $Y=1.185
+ $X2=3.01 $Y2=1.1
r251 40 41 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.01 $Y=1.185
+ $X2=3.01 $Y2=1.555
r252 38 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.065 $Y=0.34
+ $X2=5.15 $Y2=0.425
r253 38 39 142.877 $w=1.68e-07 $l=2.19e-06 $layer=LI1_cond $X=5.065 $Y=0.34
+ $X2=2.875 $Y2=0.34
r254 37 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.79 $Y=1.015
+ $X2=2.79 $Y2=1.1
r255 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.79 $Y=0.425
+ $X2=2.875 $Y2=0.34
r256 36 37 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.79 $Y=0.425
+ $X2=2.79 $Y2=1.015
r257 34 64 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=1.1
+ $X2=2.79 $Y2=1.1
r258 34 35 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.705 $Y=1.1
+ $X2=2.155 $Y2=1.1
r259 30 32 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.655 $Y=2.37
+ $X2=1.805 $Y2=2.37
r260 26 35 17.2543 $w=2.7e-07 $l=3.72411e-07 $layer=LI1_cond $X=1.81 $Y=1.157
+ $X2=2.155 $Y2=1.1
r261 26 62 10.8444 $w=2.7e-07 $l=2.4e-07 $layer=LI1_cond $X=1.81 $Y=1.157
+ $X2=1.57 $Y2=1.157
r262 26 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.81 $Y=1.015
+ $X2=1.81 $Y2=0.74
r263 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.57 $Y=2.285
+ $X2=1.655 $Y2=2.37
r264 24 62 3.44395 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.57 $Y=1.3
+ $X2=1.57 $Y2=1.157
r265 24 25 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=1.57 $Y=1.3
+ $X2=1.57 $Y2=2.285
r266 22 23 55.4135 $w=1.85e-07 $l=1.5e-07 $layer=POLY_cond $X=3.012 $Y=0.9
+ $X2=3.012 $Y2=1.05
r267 18 77 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.34 $Y=1.845
+ $X2=3.34 $Y2=1.68
r268 18 20 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=3.34 $Y=1.845
+ $X2=3.34 $Y2=2.635
r269 17 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.03 $Y=1.515
+ $X2=3.03 $Y2=1.68
r270 17 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.03 $Y=1.515
+ $X2=3.03 $Y2=1.05
r271 15 22 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.995 $Y=0.615
+ $X2=2.995 $Y2=0.9
r272 4 60 300 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=2 $X=7.665
+ $Y=1.945 $X2=7.795 $Y2=2.09
r273 3 32 600 $w=1.7e-07 $l=4.72705e-07 $layer=licon1_PDIFF $count=1 $X=1.67
+ $Y=1.96 $X2=1.805 $Y2=2.37
r274 2 54 182 $w=1.7e-07 $l=2.48898e-07 $layer=licon1_NDIFF $count=1 $X=8.405
+ $Y=0.425 $X2=8.615 $Y2=0.34
r275 1 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.67
+ $Y=0.595 $X2=1.81 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_2%A_818_418# 1 2 9 13 17 19 22 24 25 26 31 34
+ 37 39 42 43 44 46 48 49 54 56 60 61
c157 61 0 2.09165e-19 $X=8.455 $Y=1.44
c158 22 0 2.33767e-20 $X=8.7 $Y=2.155
c159 13 0 1.97119e-19 $X=4.265 $Y=1.37
c160 9 0 7.64129e-20 $X=4.18 $Y=2.635
r161 61 67 37.1352 $w=3.18e-07 $l=2.45e-07 $layer=POLY_cond $X=8.455 $Y=1.44
+ $X2=8.7 $Y2=1.44
r162 61 65 18.9465 $w=3.18e-07 $l=1.25e-07 $layer=POLY_cond $X=8.455 $Y=1.44
+ $X2=8.33 $Y2=1.44
r163 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.455
+ $Y=1.44 $X2=8.455 $Y2=1.44
r164 57 60 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=8.135 $Y=1.44
+ $X2=8.455 $Y2=1.44
r165 52 54 0.432166 $w=3.98e-07 $l=1.5e-08 $layer=LI1_cond $X=5.605 $Y=2.04
+ $X2=5.62 $Y2=2.04
r166 51 52 9.93982 $w=3.98e-07 $l=3.45e-07 $layer=LI1_cond $X=5.26 $Y=2.04
+ $X2=5.605 $Y2=2.04
r167 48 51 3.16922 $w=3.98e-07 $l=1.1e-07 $layer=LI1_cond $X=5.15 $Y=2.04
+ $X2=5.26 $Y2=2.04
r168 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.15
+ $Y=2.075 $X2=5.15 $Y2=2.075
r169 45 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.135 $Y=1.605
+ $X2=8.135 $Y2=1.44
r170 45 46 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=8.135 $Y=1.605
+ $X2=8.135 $Y2=2.905
r171 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.05 $Y=2.99
+ $X2=8.135 $Y2=2.905
r172 43 44 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=8.05 $Y=2.99
+ $X2=7.505 $Y2=2.99
r173 42 44 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=7.41 $Y=2.905
+ $X2=7.505 $Y2=2.99
r174 41 42 18.0957 $w=1.88e-07 $l=3.1e-07 $layer=LI1_cond $X=7.41 $Y=2.595
+ $X2=7.41 $Y2=2.905
r175 40 56 4.14084 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=5.785 $Y=2.51
+ $X2=5.605 $Y2=2.51
r176 39 41 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=7.315 $Y=2.51
+ $X2=7.41 $Y2=2.595
r177 39 40 99.8182 $w=1.68e-07 $l=1.53e-06 $layer=LI1_cond $X=7.315 $Y=2.51
+ $X2=5.785 $Y2=2.51
r178 35 56 2.66603 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.605 $Y=2.595
+ $X2=5.605 $Y2=2.51
r179 35 37 7.04271 $w=3.58e-07 $l=2.2e-07 $layer=LI1_cond $X=5.605 $Y=2.595
+ $X2=5.605 $Y2=2.815
r180 34 56 2.66603 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.605 $Y=2.425
+ $X2=5.605 $Y2=2.51
r181 33 52 1.35108 $w=3.6e-07 $l=2e-07 $layer=LI1_cond $X=5.605 $Y=2.24
+ $X2=5.605 $Y2=2.04
r182 33 34 5.92228 $w=3.58e-07 $l=1.85e-07 $layer=LI1_cond $X=5.605 $Y=2.24
+ $X2=5.605 $Y2=2.425
r183 29 51 1.86583 $w=3.3e-07 $l=2e-07 $layer=LI1_cond $X=5.26 $Y=1.84 $X2=5.26
+ $Y2=2.04
r184 29 31 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=5.26 $Y=1.84
+ $X2=5.26 $Y2=1.085
r185 25 49 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.81 $Y=2.075
+ $X2=5.15 $Y2=2.075
r186 25 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.81 $Y=2.075
+ $X2=4.645 $Y2=2.075
r187 20 67 16.0701 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.7 $Y=1.605
+ $X2=8.7 $Y2=1.44
r188 20 22 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=8.7 $Y=1.605 $X2=8.7
+ $Y2=2.155
r189 17 65 20.3436 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.33 $Y=1.275
+ $X2=8.33 $Y2=1.44
r190 17 19 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.33 $Y=1.275
+ $X2=8.33 $Y2=0.795
r191 16 24 6.66866 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=4.34 $Y=2.165
+ $X2=4.215 $Y2=2.165
r192 16 26 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=4.34 $Y=2.165
+ $X2=4.645 $Y2=2.165
r193 11 24 18.8402 $w=1.65e-07 $l=9.68246e-08 $layer=POLY_cond $X=4.265 $Y=2.09
+ $X2=4.215 $Y2=2.165
r194 11 13 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=4.265 $Y=2.09
+ $X2=4.265 $Y2=1.37
r195 7 24 18.8402 $w=1.65e-07 $l=9.08295e-08 $layer=POLY_cond $X=4.18 $Y=2.24
+ $X2=4.215 $Y2=2.165
r196 7 9 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=4.18 $Y=2.24 $X2=4.18
+ $Y2=2.635
r197 2 54 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=5.475
+ $Y=1.84 $X2=5.62 $Y2=2.005
r198 2 37 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=5.475
+ $Y=1.84 $X2=5.62 $Y2=2.815
r199 1 31 182 $w=1.7e-07 $l=6.56791e-07 $layer=licon1_NDIFF $count=1 $X=5.13
+ $Y=0.49 $X2=5.26 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_2%A_728_331# 1 2 9 14 15 16 20 23 25 29 31 33
+ 35 42 44 46 49 53 54 56 61 65 66 72
c163 46 0 9.04021e-20 $X=6.45 $Y=1.34
c164 31 0 1.9418e-19 $X=8.02 $Y=1.87
c165 9 0 1.97872e-19 $X=3.73 $Y=2.635
r166 67 69 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=5.475 $Y=1.505
+ $X2=5.845 $Y2=1.505
r167 64 66 5.09823 $w=4.13e-07 $l=1.65e-07 $layer=LI1_cond $X=6.87 $Y=2.047
+ $X2=7.035 $Y2=2.047
r168 64 65 5.09823 $w=4.13e-07 $l=1.65e-07 $layer=LI1_cond $X=6.87 $Y=2.047
+ $X2=6.705 $Y2=2.047
r169 58 61 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=6.45 $Y=0.8
+ $X2=6.795 $Y2=0.8
r170 55 56 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=6.18 $Y=1.505
+ $X2=6.45 $Y2=1.505
r171 54 69 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=6.1 $Y=1.505
+ $X2=5.845 $Y2=1.505
r172 53 55 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=6.1 $Y=1.505 $X2=6.18
+ $Y2=1.505
r173 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.1
+ $Y=1.505 $X2=6.1 $Y2=1.505
r174 50 72 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=7.34 $Y=2.005
+ $X2=7.34 $Y2=1.795
r175 49 66 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=7.34 $Y=2.005
+ $X2=7.035 $Y2=2.005
r176 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.34
+ $Y=2.005 $X2=7.34 $Y2=2.005
r177 46 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.45 $Y=1.34
+ $X2=6.45 $Y2=1.505
r178 45 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.45 $Y=0.965
+ $X2=6.45 $Y2=0.8
r179 45 46 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.45 $Y=0.965
+ $X2=6.45 $Y2=1.34
r180 44 65 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=6.265 $Y=2.005
+ $X2=6.705 $Y2=2.005
r181 42 44 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.18 $Y=1.84
+ $X2=6.265 $Y2=2.005
r182 41 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.18 $Y=1.67
+ $X2=6.18 $Y2=1.505
r183 41 42 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.18 $Y=1.67
+ $X2=6.18 $Y2=1.84
r184 34 35 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.775 $Y=1.655
+ $X2=3.775 $Y2=1.805
r185 31 36 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.02 $Y=1.795
+ $X2=7.855 $Y2=1.795
r186 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.02 $Y=1.87
+ $X2=8.02 $Y2=2.445
r187 27 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.855 $Y=1.72
+ $X2=7.855 $Y2=1.795
r188 27 29 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=7.855 $Y=1.72
+ $X2=7.855 $Y2=0.955
r189 26 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.505 $Y=1.795
+ $X2=7.34 $Y2=1.795
r190 25 36 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.78 $Y=1.795
+ $X2=7.855 $Y2=1.795
r191 25 26 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=7.78 $Y=1.795
+ $X2=7.505 $Y2=1.795
r192 21 69 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.845 $Y=1.67
+ $X2=5.845 $Y2=1.505
r193 21 23 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=5.845 $Y=1.67
+ $X2=5.845 $Y2=2.4
r194 18 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.475 $Y=1.34
+ $X2=5.475 $Y2=1.505
r195 18 20 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.475 $Y=1.34
+ $X2=5.475 $Y2=0.86
r196 17 20 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.475 $Y=0.415
+ $X2=5.475 $Y2=0.86
r197 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.4 $Y=0.34
+ $X2=5.475 $Y2=0.415
r198 15 16 764.021 $w=1.5e-07 $l=1.49e-06 $layer=POLY_cond $X=5.4 $Y=0.34
+ $X2=3.91 $Y2=0.34
r199 14 34 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.835 $Y=1.37
+ $X2=3.835 $Y2=1.655
r200 11 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.835 $Y=0.415
+ $X2=3.91 $Y2=0.34
r201 11 14 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=3.835 $Y=0.415
+ $X2=3.835 $Y2=1.37
r202 9 35 322.629 $w=1.8e-07 $l=8.3e-07 $layer=POLY_cond $X=3.73 $Y=2.635
+ $X2=3.73 $Y2=1.805
r203 2 64 600 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_PDIFF $count=1 $X=6.735
+ $Y=1.84 $X2=6.87 $Y2=2.045
r204 1 61 182 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_NDIFF $count=1 $X=6.655
+ $Y=0.49 $X2=6.795 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_2%CLK 1 3 6 8 11
c42 11 0 1.7376e-19 $X=6.645 $Y=1.505
r43 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.8
+ $Y=1.505 $X2=6.8 $Y2=1.505
r44 11 13 24.1 $w=3.1e-07 $l=1.55e-07 $layer=POLY_cond $X=6.645 $Y=1.505 $X2=6.8
+ $Y2=1.505
r45 10 11 10.1065 $w=3.1e-07 $l=6.5e-08 $layer=POLY_cond $X=6.58 $Y=1.505
+ $X2=6.645 $Y2=1.505
r46 8 14 7.11803 $w=3.38e-07 $l=2.1e-07 $layer=LI1_cond $X=6.875 $Y=1.295
+ $X2=6.875 $Y2=1.505
r47 4 11 15.4789 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.645 $Y=1.67
+ $X2=6.645 $Y2=1.505
r48 4 6 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=6.645 $Y=1.67
+ $X2=6.645 $Y2=2.4
r49 1 10 19.7411 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.58 $Y=1.34
+ $X2=6.58 $Y2=1.505
r50 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.58 $Y=1.34 $X2=6.58
+ $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_2%A_1800_291# 1 2 9 13 15 18 22 23 26 27 30 33
+ 34 38 41
c92 30 0 1.06861e-19 $X=10.59 $Y=1.95
c93 23 0 1.76421e-19 $X=9.165 $Y=1.62
c94 22 0 2.33767e-20 $X=9.165 $Y=1.62
r95 36 38 6.10934 $w=4.13e-07 $l=2.2e-07 $layer=LI1_cond $X=10.37 $Y=0.557
+ $X2=10.59 $Y2=0.557
r96 32 34 8.80985 $w=4.33e-07 $l=1.65e-07 $layer=LI1_cond $X=9.995 $Y=2.167
+ $X2=10.16 $Y2=2.167
r97 32 33 8.80985 $w=4.33e-07 $l=1.65e-07 $layer=LI1_cond $X=9.995 $Y=2.167
+ $X2=9.83 $Y2=2.167
r98 29 38 6.00275 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=10.59 $Y=0.765
+ $X2=10.59 $Y2=0.557
r99 29 30 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=10.59 $Y=0.765
+ $X2=10.59 $Y2=1.95
r100 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.505 $Y=2.035
+ $X2=10.59 $Y2=1.95
r101 27 34 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=10.505 $Y=2.035
+ $X2=10.16 $Y2=2.035
r102 26 33 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=9.33 $Y=2.035
+ $X2=9.83 $Y2=2.035
r103 23 42 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.165 $Y=1.62
+ $X2=9.165 $Y2=1.785
r104 23 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.165 $Y=1.62
+ $X2=9.165 $Y2=1.455
r105 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.165
+ $Y=1.62 $X2=9.165 $Y2=1.62
r106 20 26 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=9.197 $Y=1.95
+ $X2=9.33 $Y2=2.035
r107 20 22 14.3512 $w=2.63e-07 $l=3.3e-07 $layer=LI1_cond $X=9.197 $Y=1.95
+ $X2=9.197 $Y2=1.62
r108 16 18 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=9.225 $Y=0.94
+ $X2=9.365 $Y2=0.94
r109 13 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.365 $Y=0.865
+ $X2=9.365 $Y2=0.94
r110 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.365 $Y=0.865
+ $X2=9.365 $Y2=0.58
r111 11 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.225 $Y=1.015
+ $X2=9.225 $Y2=0.94
r112 11 41 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=9.225 $Y=1.015
+ $X2=9.225 $Y2=1.455
r113 9 42 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=9.12 $Y=2.155
+ $X2=9.12 $Y2=1.785
r114 2 32 600 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_PDIFF $count=1 $X=9.86
+ $Y=1.945 $X2=9.995 $Y2=2.165
r115 1 36 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=10.23
+ $Y=0.37 $X2=10.37 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_2%A_1586_149# 1 2 9 13 17 19 21 24 26 28 31 35
+ 37 43 46 49 54 56 64
c136 46 0 3.0437e-19 $X=8.81 $Y=1.925
r137 57 58 6.9933 $w=4.48e-07 $l=6.5e-08 $layer=POLY_cond $X=10.155 $Y=1.267
+ $X2=10.22 $Y2=1.267
r138 50 60 54.8705 $w=4.48e-07 $l=5.1e-07 $layer=POLY_cond $X=10.245 $Y=1.267
+ $X2=10.755 $Y2=1.267
r139 50 58 2.68973 $w=4.48e-07 $l=2.5e-08 $layer=POLY_cond $X=10.245 $Y=1.267
+ $X2=10.22 $Y2=1.267
r140 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.245
+ $Y=1.1 $X2=10.245 $Y2=1.1
r141 47 56 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.895 $Y=1.1
+ $X2=8.81 $Y2=1.1
r142 47 49 47.1454 $w=3.28e-07 $l=1.35e-06 $layer=LI1_cond $X=8.895 $Y=1.1
+ $X2=10.245 $Y2=1.1
r143 46 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.81 $Y=1.925
+ $X2=8.81 $Y2=2.01
r144 45 56 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.81 $Y=1.265
+ $X2=8.81 $Y2=1.1
r145 45 46 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=8.81 $Y=1.265
+ $X2=8.81 $Y2=1.925
r146 41 54 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.515 $Y=2.01
+ $X2=8.81 $Y2=2.01
r147 41 43 2.76586 $w=2.48e-07 $l=6e-08 $layer=LI1_cond $X=8.515 $Y=2.095
+ $X2=8.515 $Y2=2.155
r148 37 56 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=8.725 $Y=1.02
+ $X2=8.81 $Y2=1.1
r149 37 39 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.725 $Y=1.02
+ $X2=8.09 $Y2=1.02
r150 33 64 33.3527 $w=4.48e-07 $l=3.1e-07 $layer=POLY_cond $X=12.05 $Y=1.267
+ $X2=11.74 $Y2=1.267
r151 33 35 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=12.05 $Y=1.185
+ $X2=12.05 $Y2=0.69
r152 29 64 24.1837 $w=1.8e-07 $l=3.33e-07 $layer=POLY_cond $X=11.74 $Y=1.6
+ $X2=11.74 $Y2=1.267
r153 29 31 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=11.74 $Y=1.6
+ $X2=11.74 $Y2=2.26
r154 26 64 17.7522 $w=4.48e-07 $l=1.65e-07 $layer=POLY_cond $X=11.575 $Y=1.267
+ $X2=11.74 $Y2=1.267
r155 26 62 39.808 $w=4.48e-07 $l=3.7e-07 $layer=POLY_cond $X=11.575 $Y=1.267
+ $X2=11.205 $Y2=1.267
r156 26 28 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=11.575 $Y=1.185
+ $X2=11.575 $Y2=0.74
r157 22 62 24.1837 $w=1.8e-07 $l=3.33e-07 $layer=POLY_cond $X=11.205 $Y=1.6
+ $X2=11.205 $Y2=1.267
r158 22 24 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=11.205 $Y=1.6
+ $X2=11.205 $Y2=2.32
r159 19 62 6.45536 $w=4.48e-07 $l=6e-08 $layer=POLY_cond $X=11.145 $Y=1.267
+ $X2=11.205 $Y2=1.267
r160 19 60 41.9598 $w=4.48e-07 $l=3.9e-07 $layer=POLY_cond $X=11.145 $Y=1.267
+ $X2=10.755 $Y2=1.267
r161 19 21 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=11.145 $Y=1.185
+ $X2=11.145 $Y2=0.74
r162 15 60 24.1837 $w=1.8e-07 $l=3.33e-07 $layer=POLY_cond $X=10.755 $Y=1.6
+ $X2=10.755 $Y2=1.267
r163 15 17 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=10.755 $Y=1.6
+ $X2=10.755 $Y2=2.32
r164 11 58 24.1837 $w=1.8e-07 $l=3.33e-07 $layer=POLY_cond $X=10.22 $Y=1.6
+ $X2=10.22 $Y2=1.267
r165 11 13 215.734 $w=1.8e-07 $l=5.55e-07 $layer=POLY_cond $X=10.22 $Y=1.6
+ $X2=10.22 $Y2=2.155
r166 7 57 28.6558 $w=1.5e-07 $l=3.32e-07 $layer=POLY_cond $X=10.155 $Y=0.935
+ $X2=10.155 $Y2=1.267
r167 7 9 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=10.155 $Y=0.935
+ $X2=10.155 $Y2=0.58
r168 2 43 600 $w=1.7e-07 $l=4.58121e-07 $layer=licon1_PDIFF $count=1 $X=8.11
+ $Y=1.945 $X2=8.475 $Y2=2.155
r169 1 39 182 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_NDIFF $count=1 $X=7.93
+ $Y=0.745 $X2=8.09 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_2%A_2366_352# 1 2 9 13 17 21 23 25 29 33 42
r61 42 43 11.4038 $w=3.17e-07 $l=7.5e-08 $layer=POLY_cond $X=13.365 $Y=1.465
+ $X2=13.44 $Y2=1.465
r62 41 42 53.9779 $w=3.17e-07 $l=3.55e-07 $layer=POLY_cond $X=13.01 $Y=1.465
+ $X2=13.365 $Y2=1.465
r63 40 41 14.4448 $w=3.17e-07 $l=9.5e-08 $layer=POLY_cond $X=12.915 $Y=1.465
+ $X2=13.01 $Y2=1.465
r64 36 38 17.3161 $w=3.1e-07 $l=4.4e-07 $layer=LI1_cond $X=12.162 $Y=1.465
+ $X2=12.162 $Y2=1.905
r65 34 40 17.4858 $w=3.17e-07 $l=1.15e-07 $layer=POLY_cond $X=12.8 $Y=1.465
+ $X2=12.915 $Y2=1.465
r66 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.8
+ $Y=1.465 $X2=12.8 $Y2=1.465
r67 31 36 0.331605 $w=3.3e-07 $l=2.68e-07 $layer=LI1_cond $X=12.43 $Y=1.465
+ $X2=12.162 $Y2=1.465
r68 31 33 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.43 $Y=1.465
+ $X2=12.8 $Y2=1.465
r69 27 36 6.53365 $w=3.1e-07 $l=2.16852e-07 $layer=LI1_cond $X=12.282 $Y=1.3
+ $X2=12.162 $Y2=1.465
r70 27 29 30.6667 $w=2.93e-07 $l=7.85e-07 $layer=LI1_cond $X=12.282 $Y=1.3
+ $X2=12.282 $Y2=0.515
r71 23 38 1.94469 $w=4.1e-07 $l=7.95236e-08 $layer=LI1_cond $X=12.1 $Y=1.945
+ $X2=12.162 $Y2=1.905
r72 23 25 18.8326 $w=4.08e-07 $l=6.7e-07 $layer=LI1_cond $X=12.1 $Y=1.945
+ $X2=12.1 $Y2=2.615
r73 19 43 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.44 $Y=1.3
+ $X2=13.44 $Y2=1.465
r74 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.44 $Y=1.3
+ $X2=13.44 $Y2=0.74
r75 15 42 15.9969 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=13.365 $Y=1.63
+ $X2=13.365 $Y2=1.465
r76 15 17 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=13.365 $Y=1.63
+ $X2=13.365 $Y2=2.4
r77 11 41 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.01 $Y=1.3
+ $X2=13.01 $Y2=1.465
r78 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.01 $Y=1.3
+ $X2=13.01 $Y2=0.74
r79 7 40 15.9969 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=12.915 $Y=1.63
+ $X2=12.915 $Y2=1.465
r80 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=12.915 $Y=1.63
+ $X2=12.915 $Y2=2.4
r81 2 38 400 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_PDIFF $count=1 $X=11.83
+ $Y=1.76 $X2=12.06 $Y2=1.905
r82 2 25 400 $w=1.7e-07 $l=9.63159e-07 $layer=licon1_PDIFF $count=1 $X=11.83
+ $Y=1.76 $X2=12.06 $Y2=2.615
r83 1 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.125
+ $Y=0.37 $X2=12.265 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_2%VPWR 1 2 3 4 5 6 7 8 9 28 30 34 36 40 44 46
+ 50 56 60 62 67 70 71 72 73 79 86 95 100 110 113 122 125 128 132
r149 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r150 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r151 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r152 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r153 117 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r154 116 119 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r155 116 117 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6 $Y=3.33
+ $X2=6 $Y2=3.33
r156 113 116 11.2572 $w=5.08e-07 $l=4.8e-07 $layer=LI1_cond $X=6.245 $Y=2.85
+ $X2=6.245 $Y2=3.33
r157 111 117 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=6 $Y2=3.33
r158 110 111 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r159 106 107 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r160 104 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r161 104 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.72 $Y2=3.33
r162 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r163 101 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.805 $Y=3.33
+ $X2=12.64 $Y2=3.33
r164 101 103 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=12.805 $Y=3.33
+ $X2=13.2 $Y2=3.33
r165 100 131 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=13.475 $Y=3.33
+ $X2=13.697 $Y2=3.33
r166 100 103 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=13.475 $Y=3.33
+ $X2=13.2 $Y2=3.33
r167 99 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r168 99 126 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.28 $Y2=3.33
r169 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r170 96 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.595 $Y=3.33
+ $X2=11.43 $Y2=3.33
r171 96 98 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=11.595 $Y=3.33
+ $X2=12.24 $Y2=3.33
r172 95 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.475 $Y=3.33
+ $X2=12.64 $Y2=3.33
r173 95 98 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=12.475 $Y=3.33
+ $X2=12.24 $Y2=3.33
r174 94 126 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r175 94 123 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.36 $Y2=3.33
r176 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r177 91 122 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=9.625 $Y=3.33
+ $X2=9.445 $Y2=3.33
r178 91 93 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=9.625 $Y=3.33
+ $X2=10.32 $Y2=3.33
r179 90 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r180 89 90 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r181 87 116 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=6.5 $Y=3.33
+ $X2=6.245 $Y2=3.33
r182 87 89 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=6.5 $Y=3.33
+ $X2=8.88 $Y2=3.33
r183 86 122 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=9.265 $Y=3.33
+ $X2=9.445 $Y2=3.33
r184 86 89 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=9.265 $Y=3.33
+ $X2=8.88 $Y2=3.33
r185 85 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r186 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r187 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r188 81 84 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r189 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r190 79 110 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=3.07 $Y2=3.33
r191 79 84 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=2.64 $Y2=3.33
r192 78 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r193 78 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r194 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r195 75 106 3.25475 $w=4.5e-07 $l=2.55e-07 $layer=LI1_cond $X=0.51 $Y=3.19
+ $X2=0.255 $Y2=3.19
r196 75 77 18.3399 $w=4.48e-07 $l=6.9e-07 $layer=LI1_cond $X=0.51 $Y=3.19
+ $X2=1.2 $Y2=3.19
r197 73 90 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.88 $Y2=3.33
r198 73 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r199 71 93 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=10.365 $Y=3.33
+ $X2=10.32 $Y2=3.33
r200 71 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.365 $Y=3.33
+ $X2=10.53 $Y2=3.33
r201 70 81 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.435 $Y=3.33
+ $X2=1.68 $Y2=3.33
r202 69 70 9.22412 $w=4.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.27 $Y=3.19
+ $X2=1.435 $Y2=3.19
r203 67 77 0.265795 $w=4.48e-07 $l=1e-08 $layer=LI1_cond $X=1.21 $Y=3.19 $X2=1.2
+ $Y2=3.19
r204 67 69 1.59477 $w=4.48e-07 $l=6e-08 $layer=LI1_cond $X=1.21 $Y=3.19 $X2=1.27
+ $Y2=3.19
r205 62 65 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=13.64 $Y=1.985
+ $X2=13.64 $Y2=2.815
r206 60 131 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=13.64 $Y=3.245
+ $X2=13.697 $Y2=3.33
r207 60 65 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.64 $Y=3.245
+ $X2=13.64 $Y2=2.815
r208 56 59 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=12.64 $Y=1.985
+ $X2=12.64 $Y2=2.815
r209 54 128 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.64 $Y=3.245
+ $X2=12.64 $Y2=3.33
r210 54 59 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=12.64 $Y=3.245
+ $X2=12.64 $Y2=2.815
r211 50 53 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=11.43 $Y=1.905
+ $X2=11.43 $Y2=2.735
r212 48 125 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.43 $Y=3.245
+ $X2=11.43 $Y2=3.33
r213 48 53 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=11.43 $Y=3.245
+ $X2=11.43 $Y2=2.735
r214 47 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.695 $Y=3.33
+ $X2=10.53 $Y2=3.33
r215 46 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.265 $Y=3.33
+ $X2=11.43 $Y2=3.33
r216 46 47 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=11.265 $Y=3.33
+ $X2=10.695 $Y2=3.33
r217 42 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.53 $Y=3.245
+ $X2=10.53 $Y2=3.33
r218 42 44 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=10.53 $Y=3.245
+ $X2=10.53 $Y2=2.375
r219 38 122 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.445 $Y=3.245
+ $X2=9.445 $Y2=3.33
r220 38 40 25.2897 $w=3.58e-07 $l=7.9e-07 $layer=LI1_cond $X=9.445 $Y=3.245
+ $X2=9.445 $Y2=2.455
r221 37 110 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.195 $Y=3.33
+ $X2=3.07 $Y2=3.33
r222 36 116 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=5.99 $Y=3.33
+ $X2=6.245 $Y2=3.33
r223 36 37 182.348 $w=1.68e-07 $l=2.795e-06 $layer=LI1_cond $X=5.99 $Y=3.33
+ $X2=3.195 $Y2=3.33
r224 32 110 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.07 $Y=3.245
+ $X2=3.07 $Y2=3.33
r225 32 34 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=3.07 $Y=3.245
+ $X2=3.07 $Y2=2.79
r226 28 106 3.59937 $w=3.95e-07 $l=2.51893e-07 $layer=LI1_cond $X=0.312 $Y=2.965
+ $X2=0.255 $Y2=3.19
r227 28 30 23.1947 $w=3.93e-07 $l=7.95e-07 $layer=LI1_cond $X=0.312 $Y=2.965
+ $X2=0.312 $Y2=2.17
r228 9 65 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=13.455
+ $Y=1.84 $X2=13.64 $Y2=2.815
r229 9 62 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=13.455
+ $Y=1.84 $X2=13.64 $Y2=1.985
r230 8 59 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=12.495
+ $Y=1.84 $X2=12.64 $Y2=2.815
r231 8 56 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=12.495
+ $Y=1.84 $X2=12.64 $Y2=1.985
r232 7 53 600 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=11.295
+ $Y=1.76 $X2=11.43 $Y2=2.735
r233 7 50 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=11.295
+ $Y=1.76 $X2=11.43 $Y2=1.905
r234 6 44 300 $w=1.7e-07 $l=5.28678e-07 $layer=licon1_PDIFF $count=2 $X=10.31
+ $Y=1.945 $X2=10.53 $Y2=2.375
r235 5 40 600 $w=1.7e-07 $l=6.16401e-07 $layer=licon1_PDIFF $count=1 $X=9.21
+ $Y=1.945 $X2=9.445 $Y2=2.455
r236 4 113 600 $w=1.7e-07 $l=1.15464e-06 $layer=licon1_PDIFF $count=1 $X=5.935
+ $Y=1.84 $X2=6.245 $Y2=2.85
r237 3 34 600 $w=1.7e-07 $l=5.16188e-07 $layer=licon1_PDIFF $count=1 $X=2.665
+ $Y=2.425 $X2=3.03 $Y2=2.79
r238 2 106 600 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.81 $X2=0.28 $Y2=3.05
r239 2 69 300 $w=1.7e-07 $l=1.24925e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.81 $X2=1.27 $Y2=3.05
r240 1 30 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.2
+ $Y=1.96 $X2=0.345 $Y2=2.17
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_2%A_70_74# 1 2 3 4 13 17 20 23 24 25 28 29 30
+ 32 33 34 35 38 39 41 43 44 48
c151 38 0 1.97872e-19 $X=4.39 $Y=2.41
r152 48 51 8.72119 $w=3.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.53 $Y=1.02
+ $X2=3.53 $Y2=1.3
r153 44 46 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.69 $Y=2.71
+ $X2=1.69 $Y2=2.99
r154 39 54 23.1732 $w=1.79e-07 $l=3.4e-07 $layer=LI1_cond $X=4.382 $Y=2.65
+ $X2=4.382 $Y2=2.99
r155 39 41 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=4.475 $Y=2.65
+ $X2=4.795 $Y2=2.65
r156 38 39 16.4005 $w=1.79e-07 $l=2.43967e-07 $layer=LI1_cond $X=4.39 $Y=2.41
+ $X2=4.382 $Y2=2.65
r157 37 38 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=4.39 $Y=1.105
+ $X2=4.39 $Y2=2.41
r158 36 48 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.715 $Y=1.02
+ $X2=3.53 $Y2=1.02
r159 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.305 $Y=1.02
+ $X2=4.39 $Y2=1.105
r160 35 36 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.305 $Y=1.02
+ $X2=3.715 $Y2=1.02
r161 33 54 1.02909 $w=1.7e-07 $l=9.2e-08 $layer=LI1_cond $X=4.29 $Y=2.99
+ $X2=4.382 $Y2=2.99
r162 33 34 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4.29 $Y=2.99
+ $X2=3.535 $Y2=2.99
r163 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.45 $Y=2.905
+ $X2=3.535 $Y2=2.99
r164 31 32 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.45 $Y=2.455
+ $X2=3.45 $Y2=2.905
r165 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.365 $Y=2.37
+ $X2=3.45 $Y2=2.455
r166 29 30 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.365 $Y=2.37
+ $X2=2.775 $Y2=2.37
r167 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.69 $Y=2.455
+ $X2=2.775 $Y2=2.37
r168 27 28 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.69 $Y=2.455
+ $X2=2.69 $Y2=2.905
r169 26 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.775 $Y=2.99
+ $X2=1.69 $Y2=2.99
r170 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.605 $Y=2.99
+ $X2=2.69 $Y2=2.905
r171 25 26 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.605 $Y=2.99
+ $X2=1.775 $Y2=2.99
r172 23 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=2.71
+ $X2=1.69 $Y2=2.71
r173 23 24 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=1.605 $Y=2.71
+ $X2=1.01 $Y2=2.71
r174 21 43 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=0.77 $Y=0.64
+ $X2=0.77 $Y2=1.95
r175 18 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.845 $Y=2.625
+ $X2=1.01 $Y2=2.71
r176 18 20 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.845 $Y=2.625
+ $X2=0.845 $Y2=2.175
r177 17 43 8.30336 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=2.115
+ $X2=0.845 $Y2=1.95
r178 17 20 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=0.845 $Y=2.115
+ $X2=0.845 $Y2=2.175
r179 13 21 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.685 $Y=0.515
+ $X2=0.77 $Y2=0.64
r180 13 15 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=0.685 $Y=0.515
+ $X2=0.49 $Y2=0.515
r181 4 41 300 $w=1.7e-07 $l=6.27495e-07 $layer=licon1_PDIFF $count=2 $X=4.27
+ $Y=2.425 $X2=4.795 $Y2=2.65
r182 3 20 600 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=0.71
+ $Y=1.96 $X2=0.845 $Y2=2.175
r183 2 51 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=1.16 $X2=3.53 $Y2=1.3
r184 1 15 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=0.35
+ $Y=0.37 $X2=0.49 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_2%Q_N 1 2 9 15 17
r29 22 24 0.73494 $w=5.81e-07 $l=3.5e-08 $layer=LI1_cond $X=11.325 $Y=1.155
+ $X2=11.36 $Y2=1.155
r30 17 24 8.39931 $w=5.81e-07 $l=4e-07 $layer=LI1_cond $X=11.76 $Y=1.155
+ $X2=11.36 $Y2=1.155
r31 13 22 5.46591 $w=2.6e-07 $l=3.85e-07 $layer=LI1_cond $X=11.325 $Y=0.77
+ $X2=11.325 $Y2=1.155
r32 13 15 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=11.325 $Y=0.77
+ $X2=11.325 $Y2=0.515
r33 9 11 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=10.98 $Y=1.935
+ $X2=10.98 $Y2=2.735
r34 7 22 7.24441 $w=5.81e-07 $l=5.30141e-07 $layer=LI1_cond $X=10.98 $Y=1.54
+ $X2=11.325 $Y2=1.155
r35 7 9 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.98 $Y=1.54
+ $X2=10.98 $Y2=1.935
r36 2 11 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.845
+ $Y=1.76 $X2=10.98 $Y2=2.735
r37 2 9 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=10.845
+ $Y=1.76 $X2=10.98 $Y2=1.935
r38 1 24 182 $w=1.7e-07 $l=6.3113e-07 $layer=licon1_NDIFF $count=1 $X=11.22
+ $Y=0.37 $X2=11.36 $Y2=0.935
r39 1 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=11.22
+ $Y=0.37 $X2=11.36 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_2%Q 1 2 9 11 15 16 21 25
r29 19 25 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=13.225 $Y=0.965
+ $X2=13.225 $Y2=0.925
r30 16 27 7.69388 $w=3.28e-07 $l=1.43e-07 $layer=LI1_cond $X=13.225 $Y=0.987
+ $X2=13.225 $Y2=1.13
r31 16 19 0.768295 $w=3.28e-07 $l=2.2e-08 $layer=LI1_cond $X=13.225 $Y=0.987
+ $X2=13.225 $Y2=0.965
r32 16 25 0.803218 $w=3.28e-07 $l=2.3e-08 $layer=LI1_cond $X=13.225 $Y=0.902
+ $X2=13.225 $Y2=0.925
r33 16 21 14.2135 $w=3.28e-07 $l=4.07e-07 $layer=LI1_cond $X=13.225 $Y=0.902
+ $X2=13.225 $Y2=0.495
r34 15 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=13.22 $Y=1.82
+ $X2=13.22 $Y2=1.13
r35 9 15 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=13.14 $Y=1.985
+ $X2=13.14 $Y2=1.82
r36 9 11 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=13.14 $Y=1.985
+ $X2=13.14 $Y2=2.815
r37 2 11 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=13.005
+ $Y=1.84 $X2=13.14 $Y2=2.815
r38 2 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=13.005
+ $Y=1.84 $X2=13.14 $Y2=1.985
r39 1 21 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=13.085
+ $Y=0.37 $X2=13.225 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_2%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 51 53
+ 55 58 59 61 62 64 65 67 68 69 71 98 102 107 113 116 119 123
c145 27 0 8.70277e-20 $X=1.31 $Y=0.645
r146 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r147 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r148 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r149 113 114 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r150 111 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=13.68 $Y2=0
r151 111 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=12.72 $Y2=0
r152 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r153 108 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.88 $Y=0
+ $X2=12.755 $Y2=0
r154 108 110 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=12.88 $Y=0
+ $X2=13.2 $Y2=0
r155 107 122 4.12127 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=13.56 $Y=0
+ $X2=13.74 $Y2=0
r156 107 110 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=13.56 $Y=0
+ $X2=13.2 $Y2=0
r157 106 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r158 106 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r159 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r160 103 116 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=11.965 $Y=0
+ $X2=11.795 $Y2=0
r161 103 105 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.965 $Y=0
+ $X2=12.24 $Y2=0
r162 102 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.63 $Y=0
+ $X2=12.755 $Y2=0
r163 102 105 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=12.63 $Y=0
+ $X2=12.24 $Y2=0
r164 101 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r165 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r166 98 116 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=11.625 $Y=0
+ $X2=11.795 $Y2=0
r167 98 100 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=11.625 $Y=0
+ $X2=11.28 $Y2=0
r168 97 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r169 96 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r170 94 97 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=10.8
+ $Y2=0
r171 93 96 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=9.84 $Y=0 $X2=10.8
+ $Y2=0
r172 93 94 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r173 91 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=9.84
+ $Y2=0
r174 90 91 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r175 87 90 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=6 $Y=0 $X2=9.36
+ $Y2=0
r176 87 88 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=6 $Y=0 $X2=6
+ $Y2=0
r177 85 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r178 84 85 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r179 82 85 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=5.52 $Y2=0
r180 81 84 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=5.52
+ $Y2=0
r181 81 82 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r182 79 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r183 79 114 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r184 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r185 76 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.475 $Y=0
+ $X2=1.31 $Y2=0
r186 76 78 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.475 $Y=0
+ $X2=2.16 $Y2=0
r187 74 114 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r188 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r189 71 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.145 $Y=0
+ $X2=1.31 $Y2=0
r190 71 73 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=1.145 $Y=0
+ $X2=0.24 $Y2=0
r191 69 91 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=6.96 $Y=0 $X2=9.36
+ $Y2=0
r192 69 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6
+ $Y2=0
r193 67 96 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=10.845 $Y=0
+ $X2=10.8 $Y2=0
r194 67 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.845 $Y=0
+ $X2=10.93 $Y2=0
r195 66 100 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=11.015 $Y=0
+ $X2=11.28 $Y2=0
r196 66 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.015 $Y=0
+ $X2=10.93 $Y2=0
r197 64 90 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=9.415 $Y=0 $X2=9.36
+ $Y2=0
r198 64 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.415 $Y=0 $X2=9.58
+ $Y2=0
r199 63 93 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=9.745 $Y=0 $X2=9.84
+ $Y2=0
r200 63 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.745 $Y=0 $X2=9.58
+ $Y2=0
r201 61 84 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.605 $Y=0 $X2=5.52
+ $Y2=0
r202 61 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.605 $Y=0 $X2=5.73
+ $Y2=0
r203 60 87 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=5.855 $Y=0 $X2=6
+ $Y2=0
r204 60 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.855 $Y=0 $X2=5.73
+ $Y2=0
r205 58 78 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.16
+ $Y2=0
r206 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.37
+ $Y2=0
r207 57 81 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.535 $Y=0
+ $X2=2.64 $Y2=0
r208 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.535 $Y=0 $X2=2.37
+ $Y2=0
r209 53 122 3.09095 $w=2.6e-07 $l=1.07121e-07 $layer=LI1_cond $X=13.69 $Y=0.085
+ $X2=13.74 $Y2=0
r210 53 55 19.0596 $w=2.58e-07 $l=4.3e-07 $layer=LI1_cond $X=13.69 $Y=0.085
+ $X2=13.69 $Y2=0.515
r211 49 119 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.755 $Y=0.085
+ $X2=12.755 $Y2=0
r212 49 51 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=12.755 $Y=0.085
+ $X2=12.755 $Y2=0.515
r213 45 116 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=11.795 $Y=0.085
+ $X2=11.795 $Y2=0
r214 45 47 14.575 $w=3.38e-07 $l=4.3e-07 $layer=LI1_cond $X=11.795 $Y=0.085
+ $X2=11.795 $Y2=0.515
r215 41 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.93 $Y=0.085
+ $X2=10.93 $Y2=0
r216 41 43 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=10.93 $Y=0.085
+ $X2=10.93 $Y2=0.515
r217 37 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.58 $Y=0.085
+ $X2=9.58 $Y2=0
r218 37 39 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=9.58 $Y=0.085
+ $X2=9.58 $Y2=0.555
r219 33 62 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.73 $Y=0.085
+ $X2=5.73 $Y2=0
r220 33 35 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=5.73 $Y=0.085
+ $X2=5.73 $Y2=0.325
r221 29 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.37 $Y=0.085
+ $X2=2.37 $Y2=0
r222 29 31 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=2.37 $Y=0.085
+ $X2=2.37 $Y2=0.615
r223 25 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.31 $Y=0.085
+ $X2=1.31 $Y2=0
r224 25 27 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=1.31 $Y=0.085
+ $X2=1.31 $Y2=0.645
r225 8 55 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.515
+ $Y=0.37 $X2=13.655 $Y2=0.515
r226 7 51 91 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_NDIFF $count=2 $X=12.665
+ $Y=0.37 $X2=12.795 $Y2=0.515
r227 6 47 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=11.65
+ $Y=0.37 $X2=11.795 $Y2=0.515
r228 5 43 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=10.785
+ $Y=0.37 $X2=10.93 $Y2=0.515
r229 4 39 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=9.44
+ $Y=0.37 $X2=9.58 $Y2=0.555
r230 3 35 182 $w=1.7e-07 $l=2.91033e-07 $layer=licon1_NDIFF $count=1 $X=5.55
+ $Y=0.49 $X2=5.77 $Y2=0.325
r231 2 31 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.405 $X2=2.37 $Y2=0.615
r232 1 27 182 $w=1.7e-07 $l=3.49821e-07 $layer=licon1_NDIFF $count=1 $X=1.14
+ $Y=0.37 $X2=1.31 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_2%A_614_81# 1 2 7 13
r24 11 13 27.8891 $w=2.48e-07 $l=6.05e-07 $layer=LI1_cond $X=4.77 $Y=0.765
+ $X2=4.77 $Y2=1.37
r25 7 11 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.645 $Y=0.68
+ $X2=4.77 $Y2=0.765
r26 7 9 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=4.645 $Y=0.68
+ $X2=3.21 $Y2=0.68
r27 2 13 182 $w=1.7e-07 $l=4.83735e-07 $layer=licon1_NDIFF $count=1 $X=4.34
+ $Y=1.16 $X2=4.73 $Y2=1.37
r28 1 9 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.07
+ $Y=0.405 $X2=3.21 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_2%A_1499_149# 1 2 9 11 12 14
r31 14 16 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=9.11 $Y=0.555
+ $X2=9.11 $Y2=0.68
r32 11 16 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.985 $Y=0.68
+ $X2=9.11 $Y2=0.68
r33 11 12 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=8.985 $Y=0.68
+ $X2=7.725 $Y2=0.68
r34 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.64 $Y=0.765
+ $X2=7.725 $Y2=0.68
r35 7 9 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=7.64 $Y=0.765 $X2=7.64
+ $Y2=0.955
r36 2 14 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=9.015
+ $Y=0.37 $X2=9.15 $Y2=0.555
r37 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=7.495
+ $Y=0.745 $X2=7.64 $Y2=0.955
.ends


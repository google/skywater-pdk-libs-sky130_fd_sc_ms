* File: sky130_fd_sc_ms__ha_2.spice
* Created: Wed Sep  2 12:10:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__ha_2.pex.spice"
.subckt sky130_fd_sc_ms__ha_2  VNB VPB B A VPWR SUM COUT VGND
* 
* VGND	VGND
* COUT	COUT
* SUM	SUM
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1016 A_114_74# N_B_M1016_g N_A_27_74#_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.4 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_M1009_g A_114_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.0888 PD=1.02 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75000.6 SB=75001
+ A=0.111 P=1.78 MULT=1
MM1001 N_A_278_74#_M1001_d N_A_M1001_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_B_M1007_g N_A_278_74#_M1001_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.19515 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1017 N_A_278_74#_M1017_d N_A_27_74#_M1017_g N_A_394_388#_M1017_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2011 AS=0.201625 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_SUM_M1004_d N_A_394_388#_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1221 AS=0.1962 PD=1.07 PS=2.05 NRD=4.044 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1012 N_SUM_M1004_d N_A_394_388#_M1012_g N_VGND_M1012_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1221 AS=0.1036 PD=1.07 PS=1.02 NRD=4.044 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1000 N_COUT_M1000_d N_A_27_74#_M1000_g N_VGND_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1008 N_COUT_M1000_d N_A_27_74#_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1014 N_A_27_74#_M1014_d N_B_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90004.9 A=0.18 P=2.36 MULT=1
MM1015 N_VPWR_M1015_d N_A_M1015_g N_A_27_74#_M1014_d VPB PSHORT L=0.18 W=1
+ AD=0.16425 AS=0.135 PD=1.345 PS=1.27 NRD=3.9203 NRS=0 M=1 R=5.55556 SA=90000.6
+ SB=90004.4 A=0.18 P=2.36 MULT=1
MM1005 A_310_388# N_A_M1005_g N_VPWR_M1015_d VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.16425 PD=1.24 PS=1.345 NRD=12.7853 NRS=4.9053 M=1 R=5.55556 SA=90001.1
+ SB=90004 A=0.18 P=2.36 MULT=1
MM1010 N_A_394_388#_M1010_d N_B_M1010_g A_310_388# VPB PSHORT L=0.18 W=1 AD=0.48
+ AS=0.12 PD=1.96 PS=1.24 NRD=134.925 NRS=12.7853 M=1 R=5.55556 SA=90001.5
+ SB=90003.6 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1013_d N_A_27_74#_M1013_g N_A_394_388#_M1010_d VPB PSHORT L=0.18
+ W=1 AD=0.349953 AS=0.48 PD=1.7217 PS=1.96 NRD=0 NRS=0 M=1 R=5.55556 SA=90002.7
+ SB=90002.4 A=0.18 P=2.36 MULT=1
MM1002 N_SUM_M1002_d N_A_394_388#_M1002_g N_VPWR_M1013_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.391947 PD=1.39 PS=1.9283 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90003.2 SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1003 N_SUM_M1002_d N_A_394_388#_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90003.7 SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1006 N_COUT_M1006_d N_A_27_74#_M1006_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.1
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1011 N_COUT_M1006_d N_A_27_74#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX18_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ms__ha_2.pxi.spice"
*
.ends
*
*

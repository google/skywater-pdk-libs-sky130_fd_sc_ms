* File: sky130_fd_sc_ms__o311a_2.pxi.spice
* Created: Fri Aug 28 18:00:54 2020
* 
x_PM_SKY130_FD_SC_MS__O311A_2%C1 N_C1_c_75_n N_C1_M1001_g N_C1_M1007_g
+ N_C1_c_77_n N_C1_c_78_n C1 PM_SKY130_FD_SC_MS__O311A_2%C1
x_PM_SKY130_FD_SC_MS__O311A_2%B1 N_B1_M1013_g N_B1_M1006_g B1 N_B1_c_105_n
+ N_B1_c_106_n PM_SKY130_FD_SC_MS__O311A_2%B1
x_PM_SKY130_FD_SC_MS__O311A_2%A3 N_A3_M1002_g N_A3_M1010_g A3 N_A3_c_143_n
+ N_A3_c_144_n PM_SKY130_FD_SC_MS__O311A_2%A3
x_PM_SKY130_FD_SC_MS__O311A_2%A2 N_A2_M1003_g N_A2_M1000_g A2 A2 A2 A2
+ N_A2_c_180_n N_A2_c_181_n PM_SKY130_FD_SC_MS__O311A_2%A2
x_PM_SKY130_FD_SC_MS__O311A_2%A1 N_A1_M1004_g N_A1_M1008_g A1 N_A1_c_218_n
+ N_A1_c_219_n PM_SKY130_FD_SC_MS__O311A_2%A1
x_PM_SKY130_FD_SC_MS__O311A_2%A_32_74# N_A_32_74#_M1001_s N_A_32_74#_M1007_s
+ N_A_32_74#_M1006_d N_A_32_74#_M1011_g N_A_32_74#_c_253_n N_A_32_74#_M1005_g
+ N_A_32_74#_M1012_g N_A_32_74#_c_255_n N_A_32_74#_M1009_g N_A_32_74#_c_262_n
+ N_A_32_74#_c_256_n N_A_32_74#_c_257_n N_A_32_74#_c_270_n N_A_32_74#_c_293_n
+ N_A_32_74#_c_263_n N_A_32_74#_c_264_n N_A_32_74#_c_258_n N_A_32_74#_c_259_n
+ PM_SKY130_FD_SC_MS__O311A_2%A_32_74#
x_PM_SKY130_FD_SC_MS__O311A_2%VPWR N_VPWR_M1007_d N_VPWR_M1004_d N_VPWR_M1012_s
+ N_VPWR_c_359_n N_VPWR_c_360_n N_VPWR_c_361_n N_VPWR_c_362_n N_VPWR_c_363_n
+ N_VPWR_c_364_n N_VPWR_c_365_n N_VPWR_c_366_n VPWR N_VPWR_c_367_n
+ N_VPWR_c_358_n PM_SKY130_FD_SC_MS__O311A_2%VPWR
x_PM_SKY130_FD_SC_MS__O311A_2%X N_X_M1005_d N_X_M1011_d N_X_c_416_n N_X_c_413_n
+ N_X_c_417_n N_X_c_418_n N_X_c_432_n N_X_c_433_n X X X N_X_c_415_n N_X_c_420_n
+ X PM_SKY130_FD_SC_MS__O311A_2%X
x_PM_SKY130_FD_SC_MS__O311A_2%A_219_74# N_A_219_74#_M1013_d N_A_219_74#_M1000_d
+ N_A_219_74#_c_462_n N_A_219_74#_c_459_n N_A_219_74#_c_460_n
+ PM_SKY130_FD_SC_MS__O311A_2%A_219_74#
x_PM_SKY130_FD_SC_MS__O311A_2%VGND N_VGND_M1002_d N_VGND_M1008_d N_VGND_M1009_s
+ N_VGND_c_487_n N_VGND_c_488_n N_VGND_c_489_n N_VGND_c_490_n N_VGND_c_491_n
+ N_VGND_c_492_n N_VGND_c_493_n VGND N_VGND_c_494_n N_VGND_c_495_n
+ PM_SKY130_FD_SC_MS__O311A_2%VGND
cc_1 VNB N_C1_c_75_n 0.0223455f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.22
cc_2 VNB N_C1_M1007_g 0.00857766f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.34
cc_3 VNB N_C1_c_77_n 0.0558804f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.385
cc_4 VNB N_C1_c_78_n 0.0109812f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.385
cc_5 VNB C1 0.0144311f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_B1_M1013_g 0.0252948f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.74
cc_7 VNB N_B1_c_105_n 0.0246651f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_8 VNB N_B1_c_106_n 0.00392806f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_9 VNB N_A3_M1002_g 0.0286878f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.74
cc_10 VNB N_A3_c_143_n 0.0262505f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_11 VNB N_A3_c_144_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_12 VNB N_A2_M1000_g 0.027243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_c_180_n 0.02663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_181_n 0.0016809f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_15 VNB N_A1_M1008_g 0.0257689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A1_c_218_n 0.0252921f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_17 VNB N_A1_c_219_n 0.00420079f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_18 VNB N_A_32_74#_M1011_g 0.00591612f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_19 VNB N_A_32_74#_c_253_n 0.0181781f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_20 VNB N_A_32_74#_M1012_g 0.00639648f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_21 VNB N_A_32_74#_c_255_n 0.0181832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_32_74#_c_256_n 0.00466883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_32_74#_c_257_n 0.0440786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_32_74#_c_258_n 0.00348446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_32_74#_c_259_n 0.0417409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_358_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_X_c_413_n 0.00208471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB X 0.0311383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_X_c_415_n 0.00995846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_219_74#_c_459_n 0.00284354f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_31 VNB N_A_219_74#_c_460_n 0.00238751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_487_n 0.00979921f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_33 VNB N_VGND_c_488_n 0.0125758f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_34 VNB N_VGND_c_489_n 0.0227978f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_35 VNB N_VGND_c_490_n 0.0173724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_491_n 0.0481805f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_37 VNB N_VGND_c_492_n 0.0182861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_493_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_494_n 0.0201153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_495_n 0.260862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VPB N_C1_M1007_g 0.0308788f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=2.34
cc_42 VPB N_B1_M1006_g 0.0216192f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_B1_c_105_n 0.00551218f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_44 VPB N_B1_c_106_n 0.00316297f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_45 VPB N_A3_M1010_g 0.023332f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A3_c_143_n 0.00561631f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_47 VPB N_A3_c_144_n 0.00200497f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_48 VPB N_A2_M1003_g 0.0211582f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=0.74
cc_49 VPB N_A2_c_180_n 0.0056136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A2_c_181_n 0.00258229f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_51 VPB N_A1_M1004_g 0.0226927f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=0.74
cc_52 VPB N_A1_c_218_n 0.00556387f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_53 VPB N_A1_c_219_n 0.00578906f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_54 VPB N_A_32_74#_M1011_g 0.0237717f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_55 VPB N_A_32_74#_M1012_g 0.0242679f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_56 VPB N_A_32_74#_c_262_n 0.0317411f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_32_74#_c_263_n 0.00367939f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_32_74#_c_264_n 0.0151235f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_32_74#_c_258_n 0.001194f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_359_n 0.0138424f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_61 VPB N_VPWR_c_360_n 0.00646754f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_62 VPB N_VPWR_c_361_n 0.0136263f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_362_n 0.0476283f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_363_n 0.0244728f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_364_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_365_n 0.0472569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_366_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_367_n 0.0213997f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_358_n 0.0941341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_X_c_416_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.385
cc_71 VPB N_X_c_417_n 0.00234139f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_X_c_418_n 0.00284528f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB X 0.00313078f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_X_c_420_n 0.00953878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 N_C1_c_75_n N_B1_M1013_g 0.0435734f $X=0.6 $Y=1.22 $X2=0 $Y2=0
cc_76 N_C1_c_78_n N_B1_M1013_g 0.0119264f $X=0.615 $Y=1.385 $X2=0 $Y2=0
cc_77 N_C1_M1007_g N_B1_M1006_g 0.0250444f $X=0.615 $Y=2.34 $X2=0 $Y2=0
cc_78 N_C1_M1007_g N_B1_c_105_n 0.0119264f $X=0.615 $Y=2.34 $X2=0 $Y2=0
cc_79 N_C1_M1007_g N_B1_c_106_n 3.28591e-19 $X=0.615 $Y=2.34 $X2=0 $Y2=0
cc_80 N_C1_c_78_n N_B1_c_106_n 3.63567e-19 $X=0.615 $Y=1.385 $X2=0 $Y2=0
cc_81 N_C1_M1007_g N_A_32_74#_c_262_n 0.0140228f $X=0.615 $Y=2.34 $X2=0 $Y2=0
cc_82 N_C1_c_75_n N_A_32_74#_c_256_n 0.0296397f $X=0.6 $Y=1.22 $X2=0 $Y2=0
cc_83 N_C1_c_77_n N_A_32_74#_c_256_n 0.00413135f $X=0.525 $Y=1.385 $X2=0 $Y2=0
cc_84 C1 N_A_32_74#_c_256_n 0.0200679f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_85 N_C1_M1007_g N_A_32_74#_c_270_n 3.90346e-19 $X=0.615 $Y=2.34 $X2=0 $Y2=0
cc_86 N_C1_M1007_g N_A_32_74#_c_264_n 0.0169706f $X=0.615 $Y=2.34 $X2=0 $Y2=0
cc_87 N_C1_c_77_n N_A_32_74#_c_264_n 0.00517127f $X=0.525 $Y=1.385 $X2=0 $Y2=0
cc_88 C1 N_A_32_74#_c_264_n 0.0125623f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_89 N_C1_c_75_n N_A_32_74#_c_258_n 7.45067e-19 $X=0.6 $Y=1.22 $X2=0 $Y2=0
cc_90 N_C1_M1007_g N_A_32_74#_c_258_n 0.0141394f $X=0.615 $Y=2.34 $X2=0 $Y2=0
cc_91 N_C1_c_78_n N_A_32_74#_c_258_n 0.00973665f $X=0.615 $Y=1.385 $X2=0 $Y2=0
cc_92 C1 N_A_32_74#_c_258_n 0.0265183f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_93 N_C1_M1007_g N_VPWR_c_359_n 0.00811426f $X=0.615 $Y=2.34 $X2=0 $Y2=0
cc_94 N_C1_M1007_g N_VPWR_c_363_n 0.00524835f $X=0.615 $Y=2.34 $X2=0 $Y2=0
cc_95 N_C1_M1007_g N_VPWR_c_358_n 0.00610055f $X=0.615 $Y=2.34 $X2=0 $Y2=0
cc_96 N_C1_c_75_n N_VGND_c_491_n 0.00291513f $X=0.6 $Y=1.22 $X2=0 $Y2=0
cc_97 N_C1_c_75_n N_VGND_c_495_n 0.00362985f $X=0.6 $Y=1.22 $X2=0 $Y2=0
cc_98 N_B1_M1013_g N_A3_M1002_g 0.028005f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_99 N_B1_M1006_g N_A3_M1010_g 0.02311f $X=1.185 $Y=2.34 $X2=0 $Y2=0
cc_100 N_B1_c_106_n N_A3_M1010_g 2.6794e-19 $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_101 N_B1_c_105_n N_A3_c_143_n 0.0206294f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_102 N_B1_c_106_n N_A3_c_143_n 0.00188197f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_103 N_B1_M1006_g N_A3_c_144_n 3.38956e-19 $X=1.185 $Y=2.34 $X2=0 $Y2=0
cc_104 N_B1_c_105_n N_A3_c_144_n 3.80681e-19 $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_105 N_B1_c_106_n N_A3_c_144_n 0.0347534f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_106 N_B1_M1006_g N_A_32_74#_c_262_n 6.86853e-19 $X=1.185 $Y=2.34 $X2=0 $Y2=0
cc_107 N_B1_M1013_g N_A_32_74#_c_256_n 0.00911188f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_108 N_B1_M1013_g N_A_32_74#_c_257_n 0.0154674f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_109 N_B1_c_105_n N_A_32_74#_c_257_n 0.00125196f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_110 N_B1_c_106_n N_A_32_74#_c_257_n 0.0279742f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_111 N_B1_M1006_g N_A_32_74#_c_270_n 0.0175737f $X=1.185 $Y=2.34 $X2=0 $Y2=0
cc_112 N_B1_c_105_n N_A_32_74#_c_270_n 6.98124e-19 $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_113 N_B1_c_106_n N_A_32_74#_c_270_n 0.0247432f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_114 N_B1_M1006_g N_A_32_74#_c_263_n 0.0113003f $X=1.185 $Y=2.34 $X2=0 $Y2=0
cc_115 N_B1_M1013_g N_A_32_74#_c_258_n 0.00530675f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_116 N_B1_M1006_g N_A_32_74#_c_258_n 0.0039546f $X=1.185 $Y=2.34 $X2=0 $Y2=0
cc_117 N_B1_c_106_n N_A_32_74#_c_258_n 0.03302f $X=1.11 $Y=1.515 $X2=0 $Y2=0
cc_118 N_B1_M1006_g N_VPWR_c_359_n 0.00972401f $X=1.185 $Y=2.34 $X2=0 $Y2=0
cc_119 N_B1_M1006_g N_VPWR_c_365_n 0.0055879f $X=1.185 $Y=2.34 $X2=0 $Y2=0
cc_120 N_B1_M1006_g N_VPWR_c_358_n 0.00579552f $X=1.185 $Y=2.34 $X2=0 $Y2=0
cc_121 N_B1_M1013_g N_A_219_74#_c_459_n 0.00577459f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_122 N_B1_M1013_g N_VGND_c_491_n 0.00461464f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_123 N_B1_M1013_g N_VGND_c_495_n 0.0091035f $X=1.02 $Y=0.74 $X2=0 $Y2=0
cc_124 N_A3_M1010_g N_A2_M1003_g 0.0728203f $X=1.725 $Y=2.4 $X2=0 $Y2=0
cc_125 N_A3_M1002_g N_A2_M1000_g 0.0201424f $X=1.56 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A3_c_143_n N_A2_c_180_n 0.0201104f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_127 N_A3_c_144_n N_A2_c_180_n 0.00114936f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_128 N_A3_M1010_g N_A2_c_181_n 0.00481666f $X=1.725 $Y=2.4 $X2=0 $Y2=0
cc_129 N_A3_c_143_n N_A2_c_181_n 0.00114936f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_130 N_A3_c_144_n N_A2_c_181_n 0.0276387f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_131 N_A3_M1002_g N_A_32_74#_c_257_n 0.0121365f $X=1.56 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A3_c_143_n N_A_32_74#_c_257_n 0.001245f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_133 N_A3_c_144_n N_A_32_74#_c_257_n 0.0247243f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_134 N_A3_M1010_g N_A_32_74#_c_293_n 0.00302493f $X=1.725 $Y=2.4 $X2=0 $Y2=0
cc_135 N_A3_c_143_n N_A_32_74#_c_293_n 7.63688e-19 $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_136 N_A3_c_144_n N_A_32_74#_c_293_n 0.0130747f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_137 N_A3_M1010_g N_A_32_74#_c_263_n 0.014026f $X=1.725 $Y=2.4 $X2=0 $Y2=0
cc_138 N_A3_M1010_g N_VPWR_c_359_n 0.00303034f $X=1.725 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A3_M1010_g N_VPWR_c_365_n 0.005209f $X=1.725 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A3_M1010_g N_VPWR_c_358_n 0.00988313f $X=1.725 $Y=2.4 $X2=0 $Y2=0
cc_141 N_A3_M1002_g N_A_219_74#_c_462_n 0.0101937f $X=1.56 $Y=0.74 $X2=0 $Y2=0
cc_142 N_A3_M1002_g N_A_219_74#_c_459_n 0.00821463f $X=1.56 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A3_M1002_g N_A_219_74#_c_460_n 8.12228e-19 $X=1.56 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A3_M1002_g N_VGND_c_490_n 0.00472847f $X=1.56 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A3_M1002_g N_VGND_c_491_n 0.00324657f $X=1.56 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A3_M1002_g N_VGND_c_495_n 0.00412987f $X=1.56 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A2_M1003_g N_A1_M1004_g 0.0432723f $X=2.145 $Y=2.4 $X2=0 $Y2=0
cc_148 N_A2_c_181_n N_A1_M1004_g 0.0121366f $X=2.19 $Y=1.515 $X2=0 $Y2=0
cc_149 N_A2_M1000_g N_A1_M1008_g 0.0340316f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A2_c_180_n N_A1_c_218_n 0.0173872f $X=2.19 $Y=1.515 $X2=0 $Y2=0
cc_151 N_A2_c_181_n N_A1_c_218_n 3.65288e-19 $X=2.19 $Y=1.515 $X2=0 $Y2=0
cc_152 N_A2_M1003_g N_A1_c_219_n 2.89892e-19 $X=2.145 $Y=2.4 $X2=0 $Y2=0
cc_153 N_A2_c_180_n N_A1_c_219_n 0.00202953f $X=2.19 $Y=1.515 $X2=0 $Y2=0
cc_154 N_A2_c_181_n N_A1_c_219_n 0.0349694f $X=2.19 $Y=1.515 $X2=0 $Y2=0
cc_155 N_A2_M1000_g N_A_32_74#_c_257_n 0.0115698f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A2_c_180_n N_A_32_74#_c_257_n 0.00124773f $X=2.19 $Y=1.515 $X2=0 $Y2=0
cc_157 N_A2_c_181_n N_A_32_74#_c_257_n 0.0256551f $X=2.19 $Y=1.515 $X2=0 $Y2=0
cc_158 N_A2_M1003_g N_A_32_74#_c_263_n 0.0011964f $X=2.145 $Y=2.4 $X2=0 $Y2=0
cc_159 N_A2_M1003_g N_VPWR_c_360_n 0.00177473f $X=2.145 $Y=2.4 $X2=0 $Y2=0
cc_160 N_A2_c_181_n N_VPWR_c_360_n 0.0385262f $X=2.19 $Y=1.515 $X2=0 $Y2=0
cc_161 N_A2_M1003_g N_VPWR_c_365_n 0.00363952f $X=2.145 $Y=2.4 $X2=0 $Y2=0
cc_162 N_A2_c_181_n N_VPWR_c_365_n 0.00882659f $X=2.19 $Y=1.515 $X2=0 $Y2=0
cc_163 N_A2_M1003_g N_VPWR_c_358_n 0.00445309f $X=2.145 $Y=2.4 $X2=0 $Y2=0
cc_164 N_A2_c_181_n N_VPWR_c_358_n 0.0105393f $X=2.19 $Y=1.515 $X2=0 $Y2=0
cc_165 N_A2_c_181_n A_447_368# 0.0139977f $X=2.19 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_166 N_A2_M1000_g N_A_219_74#_c_462_n 0.0101837f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A2_M1000_g N_A_219_74#_c_459_n 8.12228e-19 $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A2_M1000_g N_A_219_74#_c_460_n 0.00810322f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A2_M1000_g N_VGND_c_490_n 0.00472847f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A2_M1000_g N_VGND_c_492_n 0.00324657f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A2_M1000_g N_VGND_c_495_n 0.00412056f $X=2.28 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A1_M1004_g N_A_32_74#_M1011_g 0.021306f $X=2.685 $Y=2.4 $X2=0 $Y2=0
cc_173 N_A1_c_219_n N_A_32_74#_M1011_g 0.00231652f $X=2.76 $Y=1.515 $X2=0 $Y2=0
cc_174 N_A1_M1008_g N_A_32_74#_c_253_n 0.0202161f $X=2.71 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A1_M1008_g N_A_32_74#_c_257_n 0.0186271f $X=2.71 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A1_c_218_n N_A_32_74#_c_257_n 0.0025321f $X=2.76 $Y=1.515 $X2=0 $Y2=0
cc_177 N_A1_c_219_n N_A_32_74#_c_257_n 0.0468355f $X=2.76 $Y=1.515 $X2=0 $Y2=0
cc_178 N_A1_M1008_g N_A_32_74#_c_259_n 0.00338438f $X=2.71 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A1_c_218_n N_A_32_74#_c_259_n 0.0166495f $X=2.76 $Y=1.515 $X2=0 $Y2=0
cc_180 N_A1_c_219_n N_A_32_74#_c_259_n 2.14068e-19 $X=2.76 $Y=1.515 $X2=0 $Y2=0
cc_181 N_A1_M1004_g N_VPWR_c_360_n 0.0221038f $X=2.685 $Y=2.4 $X2=0 $Y2=0
cc_182 N_A1_c_218_n N_VPWR_c_360_n 7.73517e-19 $X=2.76 $Y=1.515 $X2=0 $Y2=0
cc_183 N_A1_c_219_n N_VPWR_c_360_n 0.0129929f $X=2.76 $Y=1.515 $X2=0 $Y2=0
cc_184 N_A1_M1004_g N_VPWR_c_365_n 0.00460063f $X=2.685 $Y=2.4 $X2=0 $Y2=0
cc_185 N_A1_M1004_g N_VPWR_c_358_n 0.00909457f $X=2.685 $Y=2.4 $X2=0 $Y2=0
cc_186 N_A1_M1004_g N_X_c_416_n 4.96188e-19 $X=2.685 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A1_M1004_g N_X_c_418_n 5.44109e-19 $X=2.685 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A1_c_219_n N_X_c_418_n 0.00266255f $X=2.76 $Y=1.515 $X2=0 $Y2=0
cc_189 N_A1_M1008_g N_A_219_74#_c_460_n 0.00681223f $X=2.71 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A1_M1008_g N_VGND_c_487_n 0.00640249f $X=2.71 $Y=0.74 $X2=0 $Y2=0
cc_191 N_A1_M1008_g N_VGND_c_492_n 0.00434272f $X=2.71 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A1_M1008_g N_VGND_c_495_n 0.00821587f $X=2.71 $Y=0.74 $X2=0 $Y2=0
cc_193 N_A_32_74#_c_270_n N_VPWR_M1007_d 0.010783f $X=1.335 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_194 N_A_32_74#_c_264_n N_VPWR_M1007_d 0.00264313f $X=0.39 $Y=1.985 $X2=-0.19
+ $Y2=-0.245
cc_195 N_A_32_74#_c_262_n N_VPWR_c_359_n 0.0447429f $X=0.39 $Y=2.695 $X2=0 $Y2=0
cc_196 N_A_32_74#_c_270_n N_VPWR_c_359_n 0.0219594f $X=1.335 $Y=2.035 $X2=0
+ $Y2=0
cc_197 N_A_32_74#_c_263_n N_VPWR_c_359_n 0.0427309f $X=1.5 $Y=2.815 $X2=0 $Y2=0
cc_198 N_A_32_74#_M1011_g N_VPWR_c_360_n 0.0129017f $X=3.27 $Y=2.4 $X2=0 $Y2=0
cc_199 N_A_32_74#_M1012_g N_VPWR_c_362_n 0.00534567f $X=3.72 $Y=2.4 $X2=0 $Y2=0
cc_200 N_A_32_74#_c_262_n N_VPWR_c_363_n 0.0111301f $X=0.39 $Y=2.695 $X2=0 $Y2=0
cc_201 N_A_32_74#_c_263_n N_VPWR_c_365_n 0.014549f $X=1.5 $Y=2.815 $X2=0 $Y2=0
cc_202 N_A_32_74#_M1011_g N_VPWR_c_367_n 0.005209f $X=3.27 $Y=2.4 $X2=0 $Y2=0
cc_203 N_A_32_74#_M1012_g N_VPWR_c_367_n 0.005209f $X=3.72 $Y=2.4 $X2=0 $Y2=0
cc_204 N_A_32_74#_M1011_g N_VPWR_c_358_n 0.00984616f $X=3.27 $Y=2.4 $X2=0 $Y2=0
cc_205 N_A_32_74#_M1012_g N_VPWR_c_358_n 0.00985623f $X=3.72 $Y=2.4 $X2=0 $Y2=0
cc_206 N_A_32_74#_c_262_n N_VPWR_c_358_n 0.0128323f $X=0.39 $Y=2.695 $X2=0 $Y2=0
cc_207 N_A_32_74#_c_263_n N_VPWR_c_358_n 0.0119743f $X=1.5 $Y=2.815 $X2=0 $Y2=0
cc_208 N_A_32_74#_M1011_g N_X_c_416_n 0.0161638f $X=3.27 $Y=2.4 $X2=0 $Y2=0
cc_209 N_A_32_74#_M1012_g N_X_c_416_n 0.0193526f $X=3.72 $Y=2.4 $X2=0 $Y2=0
cc_210 N_A_32_74#_c_255_n N_X_c_413_n 0.0118569f $X=3.735 $Y=1.22 $X2=0 $Y2=0
cc_211 N_A_32_74#_M1012_g N_X_c_417_n 0.0167628f $X=3.72 $Y=2.4 $X2=0 $Y2=0
cc_212 N_A_32_74#_M1011_g N_X_c_418_n 0.0053409f $X=3.27 $Y=2.4 $X2=0 $Y2=0
cc_213 N_A_32_74#_M1012_g N_X_c_418_n 0.0027041f $X=3.72 $Y=2.4 $X2=0 $Y2=0
cc_214 N_A_32_74#_c_257_n N_X_c_418_n 0.0151207f $X=3.095 $Y=1.095 $X2=0 $Y2=0
cc_215 N_A_32_74#_c_259_n N_X_c_418_n 0.00137795f $X=3.735 $Y=1.385 $X2=0 $Y2=0
cc_216 N_A_32_74#_c_255_n N_X_c_432_n 0.0142632f $X=3.735 $Y=1.22 $X2=0 $Y2=0
cc_217 N_A_32_74#_c_255_n N_X_c_433_n 0.00119573f $X=3.735 $Y=1.22 $X2=0 $Y2=0
cc_218 N_A_32_74#_c_257_n N_X_c_433_n 0.00614869f $X=3.095 $Y=1.095 $X2=0 $Y2=0
cc_219 N_A_32_74#_c_259_n N_X_c_433_n 0.00224023f $X=3.735 $Y=1.385 $X2=0 $Y2=0
cc_220 N_A_32_74#_c_255_n X 0.0220789f $X=3.735 $Y=1.22 $X2=0 $Y2=0
cc_221 N_A_32_74#_c_257_n X 0.0123458f $X=3.095 $Y=1.095 $X2=0 $Y2=0
cc_222 N_A_32_74#_c_256_n A_135_74# 0.00814767f $X=0.69 $Y=1.18 $X2=-0.19
+ $Y2=-0.245
cc_223 N_A_32_74#_c_257_n A_135_74# 0.00427342f $X=3.095 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_224 N_A_32_74#_c_257_n N_A_219_74#_M1013_d 0.00389656f $X=3.095 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_225 N_A_32_74#_c_257_n N_A_219_74#_M1000_d 0.00176461f $X=3.095 $Y=1.095
+ $X2=0 $Y2=0
cc_226 N_A_32_74#_c_257_n N_A_219_74#_c_462_n 0.0500659f $X=3.095 $Y=1.095 $X2=0
+ $Y2=0
cc_227 N_A_32_74#_c_256_n N_A_219_74#_c_459_n 0.0216996f $X=0.69 $Y=1.18 $X2=0
+ $Y2=0
cc_228 N_A_32_74#_c_257_n N_A_219_74#_c_459_n 0.0213487f $X=3.095 $Y=1.095 $X2=0
+ $Y2=0
cc_229 N_A_32_74#_c_257_n N_A_219_74#_c_460_n 0.0167101f $X=3.095 $Y=1.095 $X2=0
+ $Y2=0
cc_230 N_A_32_74#_c_257_n N_VGND_M1002_d 0.00600992f $X=3.095 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_231 N_A_32_74#_c_257_n N_VGND_M1008_d 0.00426848f $X=3.095 $Y=1.095 $X2=0
+ $Y2=0
cc_232 N_A_32_74#_c_253_n N_VGND_c_487_n 0.00845049f $X=3.305 $Y=1.22 $X2=0
+ $Y2=0
cc_233 N_A_32_74#_c_257_n N_VGND_c_487_n 0.0262206f $X=3.095 $Y=1.095 $X2=0
+ $Y2=0
cc_234 N_A_32_74#_c_255_n N_VGND_c_489_n 0.00957981f $X=3.735 $Y=1.22 $X2=0
+ $Y2=0
cc_235 N_A_32_74#_c_256_n N_VGND_c_491_n 0.0249477f $X=0.69 $Y=1.18 $X2=0 $Y2=0
cc_236 N_A_32_74#_c_253_n N_VGND_c_494_n 0.00461464f $X=3.305 $Y=1.22 $X2=0
+ $Y2=0
cc_237 N_A_32_74#_c_255_n N_VGND_c_494_n 0.00434272f $X=3.735 $Y=1.22 $X2=0
+ $Y2=0
cc_238 N_A_32_74#_c_253_n N_VGND_c_495_n 0.00910098f $X=3.305 $Y=1.22 $X2=0
+ $Y2=0
cc_239 N_A_32_74#_c_255_n N_VGND_c_495_n 0.00442526f $X=3.735 $Y=1.22 $X2=0
+ $Y2=0
cc_240 N_A_32_74#_c_256_n N_VGND_c_495_n 0.0203135f $X=0.69 $Y=1.18 $X2=0 $Y2=0
cc_241 N_VPWR_c_360_n N_X_c_416_n 0.0586176f $X=2.91 $Y=2.115 $X2=0 $Y2=0
cc_242 N_VPWR_c_362_n N_X_c_416_n 0.0353111f $X=3.995 $Y=2.145 $X2=0 $Y2=0
cc_243 N_VPWR_c_367_n N_X_c_416_n 0.0144623f $X=3.83 $Y=3.33 $X2=0 $Y2=0
cc_244 N_VPWR_c_358_n N_X_c_416_n 0.0118344f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_245 N_VPWR_M1012_s N_X_c_417_n 0.00103113f $X=3.81 $Y=1.84 $X2=0 $Y2=0
cc_246 N_VPWR_c_362_n N_X_c_417_n 0.00793666f $X=3.995 $Y=2.145 $X2=0 $Y2=0
cc_247 N_VPWR_M1012_s N_X_c_420_n 0.00235172f $X=3.81 $Y=1.84 $X2=0 $Y2=0
cc_248 N_VPWR_c_362_n N_X_c_420_n 0.0175586f $X=3.995 $Y=2.145 $X2=0 $Y2=0
cc_249 N_X_c_432_n N_VGND_M1009_s 0.00306514f $X=3.965 $Y=0.93 $X2=0 $Y2=0
cc_250 X N_VGND_M1009_s 0.0013398f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_251 N_X_c_415_n N_VGND_M1009_s 0.00521203f $X=4.08 $Y=1.05 $X2=0 $Y2=0
cc_252 N_X_c_413_n N_VGND_c_487_n 0.0135169f $X=3.52 $Y=0.515 $X2=0 $Y2=0
cc_253 N_X_c_413_n N_VGND_c_489_n 0.00978743f $X=3.52 $Y=0.515 $X2=0 $Y2=0
cc_254 N_X_c_432_n N_VGND_c_489_n 0.00664376f $X=3.965 $Y=0.93 $X2=0 $Y2=0
cc_255 N_X_c_415_n N_VGND_c_489_n 0.0169147f $X=4.08 $Y=1.05 $X2=0 $Y2=0
cc_256 N_X_c_413_n N_VGND_c_494_n 0.0110175f $X=3.52 $Y=0.515 $X2=0 $Y2=0
cc_257 N_X_c_413_n N_VGND_c_495_n 0.0090528f $X=3.52 $Y=0.515 $X2=0 $Y2=0
cc_258 N_X_c_432_n N_VGND_c_495_n 0.00573789f $X=3.965 $Y=0.93 $X2=0 $Y2=0
cc_259 N_X_c_415_n N_VGND_c_495_n 9.73527e-19 $X=4.08 $Y=1.05 $X2=0 $Y2=0
cc_260 N_A_219_74#_c_462_n N_VGND_M1002_d 0.0112181f $X=2.33 $Y=0.755 $X2=-0.19
+ $Y2=-0.245
cc_261 N_A_219_74#_c_460_n N_VGND_c_487_n 0.0191765f $X=2.495 $Y=0.595 $X2=0
+ $Y2=0
cc_262 N_A_219_74#_c_462_n N_VGND_c_490_n 0.0351355f $X=2.33 $Y=0.755 $X2=0
+ $Y2=0
cc_263 N_A_219_74#_c_459_n N_VGND_c_490_n 0.00617451f $X=1.345 $Y=0.595 $X2=0
+ $Y2=0
cc_264 N_A_219_74#_c_460_n N_VGND_c_490_n 0.00617451f $X=2.495 $Y=0.595 $X2=0
+ $Y2=0
cc_265 N_A_219_74#_c_462_n N_VGND_c_491_n 0.00237563f $X=2.33 $Y=0.755 $X2=0
+ $Y2=0
cc_266 N_A_219_74#_c_459_n N_VGND_c_491_n 0.0142249f $X=1.345 $Y=0.595 $X2=0
+ $Y2=0
cc_267 N_A_219_74#_c_462_n N_VGND_c_492_n 0.00237563f $X=2.33 $Y=0.755 $X2=0
+ $Y2=0
cc_268 N_A_219_74#_c_460_n N_VGND_c_492_n 0.0141563f $X=2.495 $Y=0.595 $X2=0
+ $Y2=0
cc_269 N_A_219_74#_c_462_n N_VGND_c_495_n 0.0107664f $X=2.33 $Y=0.755 $X2=0
+ $Y2=0
cc_270 N_A_219_74#_c_459_n N_VGND_c_495_n 0.011867f $X=1.345 $Y=0.595 $X2=0
+ $Y2=0
cc_271 N_A_219_74#_c_460_n N_VGND_c_495_n 0.0117515f $X=2.495 $Y=0.595 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__o21bai_1.spice
* Created: Wed Sep  2 12:22:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o21bai_1.pex.spice"
.subckt sky130_fd_sc_ms__o21bai_1  VNB VPB B1_N A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_B1_N_M1001_g N_A_27_74#_M1001_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.15125 AS=0.154 PD=1.65 PS=1.66 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1003 N_A_308_74#_M1003_d N_A_27_74#_M1003_g N_Y_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1221 AS=0.2072 PD=1.07 PS=2.04 NRD=8.1 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g N_A_308_74#_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1073 AS=0.1221 PD=1.03 PS=1.07 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1002 N_A_308_74#_M1002_d N_A1_M1002_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1073 PD=2.05 PS=1.03 NRD=0 NRS=0.804 M=1 R=4.93333 SA=75001.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_B1_N_M1005_g N_A_27_74#_M1005_s VPB PSHORT L=0.18 W=0.84
+ AD=0.2982 AS=0.2352 PD=1.59857 PS=2.24 NRD=10.5395 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90002 A=0.1512 P=2.04 MULT=1
MM1006 N_Y_M1006_d N_A_27_74#_M1006_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3976 PD=1.39 PS=2.13143 NRD=0 NRS=14.0658 M=1 R=6.22222
+ SA=90000.9 SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1007 A_398_368# N_A2_M1007_g N_Y_M1006_d VPB PSHORT L=0.18 W=1.12 AD=0.168
+ AS=0.1512 PD=1.42 PS=1.39 NRD=16.7056 NRS=0 M=1 R=6.22222 SA=90001.3
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g A_398_368# VPB PSHORT L=0.18 W=1.12 AD=0.308
+ AS=0.168 PD=2.79 PS=1.42 NRD=0 NRS=16.7056 M=1 R=6.22222 SA=90001.8 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ms__o21bai_1.pxi.spice"
*
.ends
*
*

* NGSPICE file created from sky130_fd_sc_ms__o21ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 VPWR A1 a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=9.296e+11p pd=8.38e+06u as=6.608e+11p ps=5.66e+06u
M1001 a_119_368# A2 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=6.608e+11p ps=5.66e+06u
M1002 a_119_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y A2 a_119_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=2.331e+11p pd=2.11e+06u as=8.806e+11p ps=8.3e+06u
M1006 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=5.069e+11p ps=4.33e+06u
M1008 a_27_74# B1 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


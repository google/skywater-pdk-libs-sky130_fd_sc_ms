# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__or4bb_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__or4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.471000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.525000 1.180000 8.535000 1.550000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.471000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.450000 7.075000 1.780000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.375000 1.350000 3.715000 1.780000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.350000 0.835000 1.780000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  1.610300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.180000 1.450000 2.050000 ;
        RECT 1.085000 2.050000 2.525000 2.220000 ;
        RECT 1.120000 0.350000 1.450000 0.580000 ;
        RECT 1.120000 0.580000 2.775000 0.750000 ;
        RECT 1.120000 0.750000 1.450000 1.180000 ;
        RECT 2.140000 0.420000 2.775000 0.580000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.640000 0.085000 ;
        RECT 0.615000  0.085000 0.915000 1.130000 ;
        RECT 1.630000  0.085000 1.960000 0.410000 ;
        RECT 2.945000  0.085000 3.275000 0.750000 ;
        RECT 4.015000  0.085000 4.605000 0.410000 ;
        RECT 6.450000  0.085000 6.780000 0.920000 ;
        RECT 7.640000  0.085000 8.310000 0.985000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 8.640000 3.415000 ;
        RECT 0.650000 2.730000 0.995000 3.245000 ;
        RECT 1.565000 2.730000 1.990000 3.245000 ;
        RECT 2.840000 2.730000 3.170000 3.245000 ;
        RECT 7.745000 2.410000 8.075000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.450000 0.445000 1.130000 ;
      RECT 0.085000 1.130000 0.255000 1.950000 ;
      RECT 0.085000 1.950000 0.445000 2.390000 ;
      RECT 0.085000 2.390000 2.865000 2.560000 ;
      RECT 0.085000 2.560000 0.445000 2.860000 ;
      RECT 1.620000 0.920000 4.275000 1.090000 ;
      RECT 1.620000 1.090000 1.790000 1.710000 ;
      RECT 1.620000 1.710000 2.865000 1.880000 ;
      RECT 1.960000 1.260000 3.205000 1.540000 ;
      RECT 2.695000 1.880000 2.865000 2.390000 ;
      RECT 3.035000 1.540000 3.205000 2.290000 ;
      RECT 3.035000 2.290000 4.715000 2.460000 ;
      RECT 3.375000 1.950000 4.055000 2.120000 ;
      RECT 3.455000 0.450000 3.785000 0.580000 ;
      RECT 3.455000 0.580000 4.615000 0.750000 ;
      RECT 3.885000 1.420000 5.805000 1.590000 ;
      RECT 3.885000 1.590000 4.055000 1.950000 ;
      RECT 3.935000 2.630000 5.165000 2.905000 ;
      RECT 3.935000 2.905000 6.115000 2.980000 ;
      RECT 3.945000 1.090000 4.275000 1.250000 ;
      RECT 4.385000 1.760000 6.145000 1.930000 ;
      RECT 4.385000 1.930000 4.715000 2.290000 ;
      RECT 4.445000 0.750000 4.615000 1.260000 ;
      RECT 4.445000 1.260000 5.805000 1.420000 ;
      RECT 4.785000 0.350000 6.280000 1.090000 ;
      RECT 4.835000 2.980000 6.115000 3.075000 ;
      RECT 5.335000 2.100000 7.045000 2.270000 ;
      RECT 5.335000 2.270000 5.665000 2.735000 ;
      RECT 5.865000 2.440000 6.115000 2.905000 ;
      RECT 5.975000 1.090000 7.355000 1.260000 ;
      RECT 5.975000 1.260000 6.145000 1.760000 ;
      RECT 6.345000 2.440000 6.675000 2.905000 ;
      RECT 6.345000 2.905000 7.575000 3.075000 ;
      RECT 6.575000 1.950000 7.045000 2.100000 ;
      RECT 6.875000 2.270000 7.045000 2.735000 ;
      RECT 7.025000 0.350000 7.355000 1.090000 ;
      RECT 7.245000 1.950000 8.525000 2.240000 ;
      RECT 7.245000 2.240000 7.575000 2.905000 ;
      RECT 8.195000 1.940000 8.525000 1.950000 ;
      RECT 8.250000 2.240000 8.525000 2.990000 ;
  END
END sky130_fd_sc_ms__or4bb_4

* NGSPICE file created from sky130_fd_sc_ms__nand2b_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__nand2b_1 A_N B VGND VNB VPB VPWR Y
M1000 Y a_27_112# a_269_74# VNB nlowvt w=740000u l=150000u
+  ad=3.182e+11p pd=2.34e+06u as=1.776e+11p ps=1.96e+06u
M1001 a_269_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.4825e+11p ps=2.73e+06u
M1002 VPWR A_N a_27_112# VPB pshort w=840000u l=180000u
+  ad=8.47e+11p pd=6.03e+06u as=2.352e+11p ps=2.24e+06u
M1003 VGND A_N a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1004 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.584e+11p pd=2.88e+06u as=0p ps=0u
M1005 VPWR a_27_112# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__mux4_1.pxi.spice
* Created: Fri Aug 28 17:40:51 2020
* 
x_PM_SKY130_FD_SC_MS__MUX4_1%A0 N_A0_M1020_g N_A0_M1014_g A0 N_A0_c_184_n
+ N_A0_c_185_n PM_SKY130_FD_SC_MS__MUX4_1%A0
x_PM_SKY130_FD_SC_MS__MUX4_1%A_27_74# N_A_27_74#_M1021_s N_A_27_74#_M1009_s
+ N_A_27_74#_M1015_g N_A_27_74#_M1013_g N_A_27_74#_M1022_g N_A_27_74#_M1005_g
+ N_A_27_74#_c_218_n N_A_27_74#_c_241_n N_A_27_74#_c_219_n N_A_27_74#_c_308_p
+ N_A_27_74#_c_220_n N_A_27_74#_c_221_n N_A_27_74#_c_260_p N_A_27_74#_c_222_n
+ N_A_27_74#_c_223_n N_A_27_74#_c_224_n N_A_27_74#_c_225_n N_A_27_74#_c_226_n
+ N_A_27_74#_c_227_n N_A_27_74#_c_228_n N_A_27_74#_c_229_n N_A_27_74#_c_230_n
+ N_A_27_74#_c_231_n N_A_27_74#_c_245_n N_A_27_74#_c_232_n N_A_27_74#_c_342_p
+ N_A_27_74#_c_233_n N_A_27_74#_c_234_n N_A_27_74#_c_235_n N_A_27_74#_c_236_n
+ N_A_27_74#_c_237_n N_A_27_74#_c_238_n PM_SKY130_FD_SC_MS__MUX4_1%A_27_74#
x_PM_SKY130_FD_SC_MS__MUX4_1%A1 N_A1_M1001_g N_A1_M1000_g A1 A1 N_A1_c_401_n
+ N_A1_c_402_n PM_SKY130_FD_SC_MS__MUX4_1%A1
x_PM_SKY130_FD_SC_MS__MUX4_1%A2 N_A2_M1002_g N_A2_M1023_g A2 A2 N_A2_c_441_n
+ N_A2_c_442_n PM_SKY130_FD_SC_MS__MUX4_1%A2
x_PM_SKY130_FD_SC_MS__MUX4_1%S0 N_S0_M1021_g N_S0_M1009_g N_S0_c_488_n
+ N_S0_c_489_n N_S0_c_479_n N_S0_M1010_g N_S0_M1019_g N_S0_c_491_n N_S0_M1008_g
+ N_S0_c_493_n N_S0_c_494_n N_S0_c_481_n N_S0_c_482_n N_S0_M1003_g N_S0_c_483_n
+ N_S0_c_496_n N_S0_c_484_n S0 N_S0_c_485_n N_S0_c_486_n
+ PM_SKY130_FD_SC_MS__MUX4_1%S0
x_PM_SKY130_FD_SC_MS__MUX4_1%A3 N_A3_c_599_n N_A3_M1025_g N_A3_c_600_n
+ N_A3_c_601_n N_A3_c_602_n N_A3_M1012_g A3 PM_SKY130_FD_SC_MS__MUX4_1%A3
x_PM_SKY130_FD_SC_MS__MUX4_1%A_1396_99# N_A_1396_99#_M1011_s
+ N_A_1396_99#_M1016_s N_A_1396_99#_M1024_g N_A_1396_99#_M1006_g
+ N_A_1396_99#_c_643_n N_A_1396_99#_c_644_n N_A_1396_99#_c_650_n
+ N_A_1396_99#_c_645_n N_A_1396_99#_c_646_n N_A_1396_99#_c_652_n
+ N_A_1396_99#_c_647_n N_A_1396_99#_c_648_n
+ PM_SKY130_FD_SC_MS__MUX4_1%A_1396_99#
x_PM_SKY130_FD_SC_MS__MUX4_1%S1 N_S1_M1004_g N_S1_M1007_g N_S1_c_706_n
+ N_S1_c_707_n N_S1_c_708_n N_S1_M1016_g N_S1_M1011_g N_S1_c_710_n S1
+ N_S1_c_711_n PM_SKY130_FD_SC_MS__MUX4_1%S1
x_PM_SKY130_FD_SC_MS__MUX4_1%A_1338_125# N_A_1338_125#_M1004_d
+ N_A_1338_125#_M1007_d N_A_1338_125#_M1017_g N_A_1338_125#_M1018_g
+ N_A_1338_125#_c_782_n N_A_1338_125#_c_783_n N_A_1338_125#_c_788_n
+ N_A_1338_125#_c_789_n N_A_1338_125#_c_808_n N_A_1338_125#_c_809_n
+ N_A_1338_125#_c_810_n N_A_1338_125#_c_790_n N_A_1338_125#_c_784_n
+ N_A_1338_125#_c_785_n PM_SKY130_FD_SC_MS__MUX4_1%A_1338_125#
x_PM_SKY130_FD_SC_MS__MUX4_1%VPWR N_VPWR_M1009_d N_VPWR_M1000_d N_VPWR_M1012_d
+ N_VPWR_M1016_d N_VPWR_c_862_n N_VPWR_c_863_n N_VPWR_c_864_n N_VPWR_c_865_n
+ N_VPWR_c_866_n N_VPWR_c_867_n N_VPWR_c_868_n N_VPWR_c_869_n VPWR
+ N_VPWR_c_870_n N_VPWR_c_871_n N_VPWR_c_872_n N_VPWR_c_861_n N_VPWR_c_874_n
+ N_VPWR_c_875_n PM_SKY130_FD_SC_MS__MUX4_1%VPWR
x_PM_SKY130_FD_SC_MS__MUX4_1%A_342_74# N_A_342_74#_M1015_d N_A_342_74#_M1024_d
+ N_A_342_74#_M1010_d N_A_342_74#_M1007_s N_A_342_74#_c_970_n
+ N_A_342_74#_c_971_n N_A_342_74#_c_958_n N_A_342_74#_c_959_n
+ N_A_342_74#_c_960_n N_A_342_74#_c_1088_p N_A_342_74#_c_961_n
+ N_A_342_74#_c_1072_p N_A_342_74#_c_962_n N_A_342_74#_c_963_n
+ N_A_342_74#_c_964_n N_A_342_74#_c_952_n N_A_342_74#_c_953_n
+ N_A_342_74#_c_965_n N_A_342_74#_c_954_n N_A_342_74#_c_967_n
+ N_A_342_74#_c_955_n N_A_342_74#_c_1035_n N_A_342_74#_c_956_n
+ N_A_342_74#_c_957_n PM_SKY130_FD_SC_MS__MUX4_1%A_342_74#
x_PM_SKY130_FD_SC_MS__MUX4_1%A_846_74# N_A_846_74#_M1022_d N_A_846_74#_M1004_s
+ N_A_846_74#_M1008_d N_A_846_74#_M1006_d N_A_846_74#_c_1110_n
+ N_A_846_74#_c_1094_n N_A_846_74#_c_1095_n N_A_846_74#_c_1096_n
+ N_A_846_74#_c_1119_n N_A_846_74#_c_1097_n N_A_846_74#_c_1098_n
+ N_A_846_74#_c_1099_n N_A_846_74#_c_1100_n N_A_846_74#_c_1206_p
+ N_A_846_74#_c_1101_n N_A_846_74#_c_1107_n N_A_846_74#_c_1102_n
+ N_A_846_74#_c_1122_n N_A_846_74#_c_1146_n N_A_846_74#_c_1103_n
+ N_A_846_74#_c_1104_n N_A_846_74#_c_1105_n PM_SKY130_FD_SC_MS__MUX4_1%A_846_74#
x_PM_SKY130_FD_SC_MS__MUX4_1%X N_X_M1017_d N_X_M1018_d X X X X X X X X
+ PM_SKY130_FD_SC_MS__MUX4_1%X
x_PM_SKY130_FD_SC_MS__MUX4_1%VGND N_VGND_M1021_d N_VGND_M1001_d N_VGND_M1025_d
+ N_VGND_M1011_d N_VGND_c_1239_n N_VGND_c_1240_n N_VGND_c_1241_n N_VGND_c_1242_n
+ N_VGND_c_1243_n N_VGND_c_1244_n VGND N_VGND_c_1245_n N_VGND_c_1246_n
+ N_VGND_c_1247_n N_VGND_c_1248_n N_VGND_c_1249_n N_VGND_c_1250_n
+ N_VGND_c_1251_n PM_SKY130_FD_SC_MS__MUX4_1%VGND
cc_1 VNB N_A0_M1014_g 0.025411f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=0.69
cc_2 VNB N_A0_c_184_n 0.0262565f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.38
cc_3 VNB N_A0_c_185_n 0.00172497f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.38
cc_4 VNB N_A_27_74#_M1015_g 0.0203542f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_5 VNB N_A_27_74#_M1013_g 0.00427099f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.38
cc_6 VNB N_A_27_74#_c_218_n 0.0221849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_74#_c_219_n 0.0160355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_74#_c_220_n 0.00764472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_74#_c_221_n 0.00122403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_74#_c_222_n 0.00549441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_74#_c_223_n 0.0361351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_c_224_n 0.022974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_225_n 0.00637819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_74#_c_226_n 0.0332145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_74#_c_227_n 0.00221525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_74#_c_228_n 0.00857418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_229_n 0.00416738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_74#_c_230_n 0.0189146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_231_n 0.0128604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_74#_c_232_n 0.0293842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_74#_c_233_n 0.00555713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_234_n 0.0272559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_74#_c_235_n 0.00165995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_74#_c_236_n 2.44719e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_74#_c_237_n 0.00316465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_74#_c_238_n 0.0184364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A1_M1001_g 0.0261196f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=2.205
cc_28 VNB N_A1_c_401_n 0.0265401f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.215
cc_29 VNB N_A1_c_402_n 0.0016809f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.545
cc_30 VNB N_A2_M1023_g 0.0239399f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=0.69
cc_31 VNB N_A2_c_441_n 0.0268555f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.215
cc_32 VNB N_A2_c_442_n 0.00393472f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.545
cc_33 VNB N_S0_M1021_g 0.031278f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=2.205
cc_34 VNB N_S0_M1009_g 0.00513885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_S0_c_479_n 0.00575642f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.38
cc_36 VNB N_S0_M1010_g 0.0162592f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.215
cc_37 VNB N_S0_c_481_n 0.0262749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_S0_c_482_n 0.016835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_S0_c_483_n 0.017478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_S0_c_484_n 0.0137658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_S0_c_485_n 0.0324204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_S0_c_486_n 0.00535787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A3_c_599_n 0.018887f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.545
cc_44 VNB N_A3_c_600_n 0.0207701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A3_c_601_n 0.00576594f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=1.215
cc_46 VNB N_A3_c_602_n 0.0818175f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=0.69
cc_47 VNB N_A_1396_99#_M1024_g 0.0192719f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_48 VNB N_A_1396_99#_M1006_g 0.0037316f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.38
cc_49 VNB N_A_1396_99#_c_643_n 0.0201559f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.545
cc_50 VNB N_A_1396_99#_c_644_n 0.0139349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1396_99#_c_645_n 0.00131118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1396_99#_c_646_n 0.0053947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1396_99#_c_647_n 0.0242514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1396_99#_c_648_n 0.0246298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_S1_M1004_g 0.0301207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_S1_M1007_g 0.0101629f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=0.69
cc_57 VNB N_S1_c_706_n 0.133558f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_58 VNB N_S1_c_707_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_S1_c_708_n 0.0272457f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.38
cc_60 VNB N_S1_M1011_g 0.0314088f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.665
cc_61 VNB N_S1_c_710_n 0.0125302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_S1_c_711_n 0.00166449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1338_125#_M1017_g 0.0266178f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_64 VNB N_A_1338_125#_c_782_n 0.00113767f $X=-0.19 $Y=-0.245 $X2=1.155
+ $Y2=1.545
cc_65 VNB N_A_1338_125#_c_783_n 0.00247606f $X=-0.19 $Y=-0.245 $X2=1.155
+ $Y2=1.665
cc_66 VNB N_A_1338_125#_c_784_n 0.00326383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1338_125#_c_785_n 0.0342137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VPWR_c_861_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_342_74#_c_952_n 6.34967e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_342_74#_c_953_n 0.00629701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_342_74#_c_954_n 0.00353895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_342_74#_c_955_n 0.00426504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_342_74#_c_956_n 0.00154297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_342_74#_c_957_n 0.00195188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_846_74#_c_1094_n 0.00145889f $X=-0.19 $Y=-0.245 $X2=1.155
+ $Y2=1.665
cc_76 VNB N_A_846_74#_c_1095_n 0.00881326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_846_74#_c_1096_n 0.00249378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_846_74#_c_1097_n 0.00712355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_846_74#_c_1098_n 0.00336014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_846_74#_c_1099_n 0.00209848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_846_74#_c_1100_n 0.0127993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_846_74#_c_1101_n 0.0219922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_846_74#_c_1102_n 0.0175843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_846_74#_c_1103_n 4.2192e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_846_74#_c_1104_n 0.00737477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_846_74#_c_1105_n 0.00444966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB X 0.0276704f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=0.69
cc_88 VNB X 0.012293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB X 0.0245106f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_90 VNB N_VGND_c_1239_n 0.0104518f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1240_n 0.00587384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1241_n 0.0153613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1242_n 0.0220288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1243_n 0.0761732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1244_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1245_n 0.0538813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1246_n 0.0422501f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1247_n 0.0212465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1248_n 0.521376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1249_n 0.0293189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1250_n 0.0109694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1251_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VPB N_A0_M1020_g 0.0253526f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=2.205
cc_104 VPB N_A0_c_184_n 0.00611024f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=1.38
cc_105 VPB N_A0_c_185_n 0.00695763f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=1.38
cc_106 VPB N_A_27_74#_M1013_g 0.0212724f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=1.38
cc_107 VPB N_A_27_74#_M1005_g 0.0245197f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_27_74#_c_241_n 0.035176f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_27_74#_c_228_n 0.00122182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_27_74#_c_229_n 0.00287633f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_27_74#_c_230_n 0.010399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_27_74#_c_245_n 0.00968222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_27_74#_c_232_n 0.0132382f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_27_74#_c_233_n 0.012813f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_27_74#_c_234_n 0.00971065f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A1_M1000_g 0.0200372f $X=-0.19 $Y=1.66 $X2=1.245 $Y2=0.69
cc_117 VPB N_A1_c_401_n 0.00566934f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=1.215
cc_118 VPB N_A1_c_402_n 0.00284782f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=1.545
cc_119 VPB N_A2_M1002_g 0.0209248f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=2.205
cc_120 VPB N_A2_c_441_n 0.00618392f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=1.215
cc_121 VPB N_A2_c_442_n 0.00680087f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=1.545
cc_122 VPB N_S0_M1009_g 0.0341131f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_S0_c_488_n 0.111725f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_124 VPB N_S0_c_489_n 0.0143041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_S0_M1010_g 0.0497941f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=1.215
cc_126 VPB N_S0_c_491_n 0.149869f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=1.665
cc_127 VPB N_S0_M1008_g 0.0187908f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_S0_c_493_n 0.0290327f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_S0_c_494_n 0.00937629f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_S0_c_481_n 0.00158796f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_S0_c_496_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_S0_c_485_n 0.00255986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_S0_c_486_n 0.00515833f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A3_c_602_n 0.0473878f $X=-0.19 $Y=1.66 $X2=1.245 $Y2=0.69
cc_135 VPB A3 0.00514791f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_136 VPB N_A_1396_99#_M1006_g 0.030987f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=1.38
cc_137 VPB N_A_1396_99#_c_650_n 0.00722388f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_1396_99#_c_645_n 0.0088679f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_1396_99#_c_652_n 0.00287634f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_1396_99#_c_648_n 0.0170937f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_S1_M1007_g 0.0335261f $X=-0.19 $Y=1.66 $X2=1.245 $Y2=0.69
cc_142 VPB N_S1_c_708_n 0.0112636f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=1.38
cc_143 VPB N_S1_M1016_g 0.0264805f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=1.38
cc_144 VPB N_S1_c_711_n 0.00219047f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_1338_125#_M1018_g 0.0285688f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=1.38
cc_146 VPB N_A_1338_125#_c_783_n 0.00268751f $X=-0.19 $Y=1.66 $X2=1.155
+ $Y2=1.665
cc_147 VPB N_A_1338_125#_c_788_n 0.0213298f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_1338_125#_c_789_n 0.00377614f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_1338_125#_c_790_n 0.00254161f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_1338_125#_c_784_n 0.00121771f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_1338_125#_c_785_n 0.00865749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_862_n 0.0135861f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=1.545
cc_153 VPB N_VPWR_c_863_n 0.0136326f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_864_n 0.010261f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_865_n 0.00661086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_866_n 0.0213239f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_867_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_868_n 0.0657218f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_869_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_870_n 0.0501803f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_871_n 0.0646356f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_872_n 0.0187203f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_861_n 0.0925525f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_874_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_875_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_342_74#_c_958_n 6.73981e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_342_74#_c_959_n 0.0129277f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_342_74#_c_960_n 0.00208963f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_342_74#_c_961_n 0.0110072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_342_74#_c_962_n 0.00315704f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_342_74#_c_963_n 0.006983f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_342_74#_c_964_n 0.00786605f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_342_74#_c_965_n 0.00975699f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_342_74#_c_954_n 0.00532049f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_342_74#_c_967_n 0.00393611f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_342_74#_c_955_n 0.00571116f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_846_74#_c_1097_n 0.00222895f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_846_74#_c_1107_n 0.00945754f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_846_74#_c_1105_n 0.00547853f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB X 0.0355463f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_181 VPB X 0.0123936f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=1.38
cc_182 N_A0_M1014_g N_A_27_74#_M1015_g 0.0488224f $X=1.245 $Y=0.69 $X2=0 $Y2=0
cc_183 N_A0_M1014_g N_A_27_74#_c_219_n 0.0129855f $X=1.245 $Y=0.69 $X2=0 $Y2=0
cc_184 N_A0_c_184_n N_A_27_74#_c_219_n 0.00123356f $X=1.155 $Y=1.38 $X2=0 $Y2=0
cc_185 N_A0_c_185_n N_A_27_74#_c_219_n 0.0236578f $X=1.155 $Y=1.38 $X2=0 $Y2=0
cc_186 N_A0_M1014_g N_A_27_74#_c_221_n 0.00120821f $X=1.245 $Y=0.69 $X2=0 $Y2=0
cc_187 N_A0_M1014_g N_A_27_74#_c_233_n 0.00119474f $X=1.245 $Y=0.69 $X2=0 $Y2=0
cc_188 N_A0_c_185_n N_A_27_74#_c_233_n 0.0199626f $X=1.155 $Y=1.38 $X2=0 $Y2=0
cc_189 N_A0_M1014_g N_A_27_74#_c_234_n 0.0201322f $X=1.245 $Y=0.69 $X2=0 $Y2=0
cc_190 N_A0_c_185_n N_A_27_74#_c_234_n 0.00109712f $X=1.155 $Y=1.38 $X2=0 $Y2=0
cc_191 N_A0_M1014_g N_A_27_74#_c_235_n 0.00324727f $X=1.245 $Y=0.69 $X2=0 $Y2=0
cc_192 N_A0_M1014_g N_S0_M1021_g 0.0162779f $X=1.245 $Y=0.69 $X2=0 $Y2=0
cc_193 N_A0_M1020_g N_S0_M1009_g 0.0198108f $X=1.2 $Y=2.205 $X2=0 $Y2=0
cc_194 N_A0_c_185_n N_S0_M1009_g 6.88557e-19 $X=1.155 $Y=1.38 $X2=0 $Y2=0
cc_195 N_A0_M1020_g N_S0_c_488_n 0.0108881f $X=1.2 $Y=2.205 $X2=0 $Y2=0
cc_196 N_A0_c_184_n N_S0_c_485_n 0.020639f $X=1.155 $Y=1.38 $X2=0 $Y2=0
cc_197 N_A0_c_185_n N_S0_c_485_n 3.80229e-19 $X=1.155 $Y=1.38 $X2=0 $Y2=0
cc_198 N_A0_M1020_g N_S0_c_486_n 6.93468e-19 $X=1.2 $Y=2.205 $X2=0 $Y2=0
cc_199 N_A0_c_184_n N_S0_c_486_n 0.00188197f $X=1.155 $Y=1.38 $X2=0 $Y2=0
cc_200 N_A0_c_185_n N_S0_c_486_n 0.0459773f $X=1.155 $Y=1.38 $X2=0 $Y2=0
cc_201 N_A0_c_185_n N_VPWR_M1009_d 0.0013515f $X=1.155 $Y=1.38 $X2=-0.19
+ $Y2=-0.245
cc_202 N_A0_M1020_g N_VPWR_c_862_n 0.00828236f $X=1.2 $Y=2.205 $X2=0 $Y2=0
cc_203 N_A0_c_184_n N_VPWR_c_862_n 2.91996e-19 $X=1.155 $Y=1.38 $X2=0 $Y2=0
cc_204 N_A0_c_185_n N_VPWR_c_862_n 0.00551427f $X=1.155 $Y=1.38 $X2=0 $Y2=0
cc_205 N_A0_M1020_g N_VPWR_c_861_n 0.00113998f $X=1.2 $Y=2.205 $X2=0 $Y2=0
cc_206 N_A0_M1014_g N_VGND_c_1239_n 0.00674196f $X=1.245 $Y=0.69 $X2=0 $Y2=0
cc_207 N_A0_M1014_g N_VGND_c_1245_n 0.00461464f $X=1.245 $Y=0.69 $X2=0 $Y2=0
cc_208 N_A0_M1014_g N_VGND_c_1248_n 0.00471211f $X=1.245 $Y=0.69 $X2=0 $Y2=0
cc_209 N_A_27_74#_c_220_n N_A1_M1001_g 0.00325205f $X=2.46 $Y=0.34 $X2=0 $Y2=0
cc_210 N_A_27_74#_c_260_p N_A1_M1001_g 0.00986281f $X=2.545 $Y=0.875 $X2=0 $Y2=0
cc_211 N_A_27_74#_c_222_n N_A1_M1001_g 0.00409499f $X=2.625 $Y=1.285 $X2=0 $Y2=0
cc_212 N_A_27_74#_c_223_n N_A1_M1001_g 0.0203929f $X=2.625 $Y=1.285 $X2=0 $Y2=0
cc_213 N_A_27_74#_c_224_n N_A1_M1001_g 0.0170535f $X=4.08 $Y=0.96 $X2=0 $Y2=0
cc_214 N_A_27_74#_M1013_g N_A1_M1000_g 0.0470724f $X=2.61 $Y=2.205 $X2=0 $Y2=0
cc_215 N_A_27_74#_M1013_g N_A1_c_401_n 0.00424196f $X=2.61 $Y=2.205 $X2=0 $Y2=0
cc_216 N_A_27_74#_c_224_n N_A1_c_401_n 0.00125621f $X=4.08 $Y=0.96 $X2=0 $Y2=0
cc_217 N_A_27_74#_M1013_g N_A1_c_402_n 0.00505379f $X=2.61 $Y=2.205 $X2=0 $Y2=0
cc_218 N_A_27_74#_c_222_n N_A1_c_402_n 0.0148928f $X=2.625 $Y=1.285 $X2=0 $Y2=0
cc_219 N_A_27_74#_c_223_n N_A1_c_402_n 8.18483e-19 $X=2.625 $Y=1.285 $X2=0 $Y2=0
cc_220 N_A_27_74#_c_224_n N_A1_c_402_n 0.0256551f $X=4.08 $Y=0.96 $X2=0 $Y2=0
cc_221 N_A_27_74#_c_224_n N_A2_M1023_g 0.0149383f $X=4.08 $Y=0.96 $X2=0 $Y2=0
cc_222 N_A_27_74#_c_225_n N_A2_M1023_g 0.00109506f $X=4.245 $Y=1.285 $X2=0 $Y2=0
cc_223 N_A_27_74#_c_238_n N_A2_M1023_g 0.0517658f $X=4.245 $Y=1.12 $X2=0 $Y2=0
cc_224 N_A_27_74#_c_224_n N_A2_c_441_n 0.00125809f $X=4.08 $Y=0.96 $X2=0 $Y2=0
cc_225 N_A_27_74#_c_225_n N_A2_c_441_n 8.18483e-19 $X=4.245 $Y=1.285 $X2=0 $Y2=0
cc_226 N_A_27_74#_c_226_n N_A2_c_441_n 0.014321f $X=4.245 $Y=1.285 $X2=0 $Y2=0
cc_227 N_A_27_74#_c_224_n N_A2_c_442_n 0.0290252f $X=4.08 $Y=0.96 $X2=0 $Y2=0
cc_228 N_A_27_74#_c_225_n N_A2_c_442_n 0.0150243f $X=4.245 $Y=1.285 $X2=0 $Y2=0
cc_229 N_A_27_74#_c_226_n N_A2_c_442_n 8.18053e-19 $X=4.245 $Y=1.285 $X2=0 $Y2=0
cc_230 N_A_27_74#_c_218_n N_S0_M1021_g 0.0126407f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_231 N_A_27_74#_c_219_n N_S0_M1021_g 0.0100334f $X=1.53 $Y=0.945 $X2=0 $Y2=0
cc_232 N_A_27_74#_c_231_n N_S0_M1021_g 0.00194563f $X=0.277 $Y=0.945 $X2=0 $Y2=0
cc_233 N_A_27_74#_c_232_n N_S0_M1021_g 0.0125596f $X=0.332 $Y=1.95 $X2=0 $Y2=0
cc_234 N_A_27_74#_c_241_n N_S0_M1009_g 0.00940135f $X=0.39 $Y=2.715 $X2=0 $Y2=0
cc_235 N_A_27_74#_c_245_n N_S0_M1009_g 0.00293377f $X=0.39 $Y=2.035 $X2=0 $Y2=0
cc_236 N_A_27_74#_c_232_n N_S0_M1009_g 0.00426393f $X=0.332 $Y=1.95 $X2=0 $Y2=0
cc_237 N_A_27_74#_M1015_g N_S0_c_479_n 0.00339648f $X=1.635 $Y=0.69 $X2=0 $Y2=0
cc_238 N_A_27_74#_c_222_n N_S0_c_479_n 0.00107031f $X=2.625 $Y=1.285 $X2=0 $Y2=0
cc_239 N_A_27_74#_c_223_n N_S0_c_479_n 0.0193839f $X=2.625 $Y=1.285 $X2=0 $Y2=0
cc_240 N_A_27_74#_M1013_g N_S0_M1010_g 0.0190645f $X=2.61 $Y=2.205 $X2=0 $Y2=0
cc_241 N_A_27_74#_c_233_n N_S0_M1010_g 3.83861e-19 $X=1.695 $Y=1.365 $X2=0 $Y2=0
cc_242 N_A_27_74#_c_234_n N_S0_M1010_g 0.0205629f $X=1.695 $Y=1.365 $X2=0 $Y2=0
cc_243 N_A_27_74#_M1013_g N_S0_c_491_n 0.0102729f $X=2.61 $Y=2.205 $X2=0 $Y2=0
cc_244 N_A_27_74#_M1005_g N_S0_c_493_n 0.00297154f $X=5.25 $Y=2.435 $X2=0 $Y2=0
cc_245 N_A_27_74#_c_228_n N_S0_c_493_n 0.0084145f $X=4.75 $Y=1.61 $X2=0 $Y2=0
cc_246 N_A_27_74#_c_229_n N_S0_c_493_n 0.0015562f $X=5.175 $Y=1.61 $X2=0 $Y2=0
cc_247 N_A_27_74#_c_237_n N_S0_c_493_n 0.00371216f $X=4.665 $Y=0.96 $X2=0 $Y2=0
cc_248 N_A_27_74#_c_225_n N_S0_c_494_n 0.00156542f $X=4.245 $Y=1.285 $X2=0 $Y2=0
cc_249 N_A_27_74#_c_226_n N_S0_c_494_n 0.0139782f $X=4.245 $Y=1.285 $X2=0 $Y2=0
cc_250 N_A_27_74#_c_227_n N_S0_c_481_n 0.00933773f $X=4.665 $Y=1.445 $X2=0 $Y2=0
cc_251 N_A_27_74#_c_228_n N_S0_c_481_n 0.00602925f $X=4.75 $Y=1.61 $X2=0 $Y2=0
cc_252 N_A_27_74#_c_229_n N_S0_c_481_n 0.00563781f $X=5.175 $Y=1.61 $X2=0 $Y2=0
cc_253 N_A_27_74#_c_230_n N_S0_c_481_n 0.0213539f $X=5.175 $Y=1.61 $X2=0 $Y2=0
cc_254 N_A_27_74#_c_227_n N_S0_c_482_n 7.98674e-19 $X=4.665 $Y=1.445 $X2=0 $Y2=0
cc_255 N_A_27_74#_c_237_n N_S0_c_482_n 0.00454612f $X=4.665 $Y=0.96 $X2=0 $Y2=0
cc_256 N_A_27_74#_c_238_n N_S0_c_482_n 0.017978f $X=4.245 $Y=1.12 $X2=0 $Y2=0
cc_257 N_A_27_74#_M1015_g N_S0_c_483_n 0.017745f $X=1.635 $Y=0.69 $X2=0 $Y2=0
cc_258 N_A_27_74#_c_308_p N_S0_c_483_n 0.00106602f $X=1.615 $Y=0.86 $X2=0 $Y2=0
cc_259 N_A_27_74#_c_220_n N_S0_c_483_n 0.0127838f $X=2.46 $Y=0.34 $X2=0 $Y2=0
cc_260 N_A_27_74#_c_260_p N_S0_c_483_n 0.0109342f $X=2.545 $Y=0.875 $X2=0 $Y2=0
cc_261 N_A_27_74#_c_222_n N_S0_c_483_n 0.00147926f $X=2.625 $Y=1.285 $X2=0 $Y2=0
cc_262 N_A_27_74#_c_236_n N_S0_c_483_n 0.00347791f $X=2.625 $Y=0.96 $X2=0 $Y2=0
cc_263 N_A_27_74#_c_225_n N_S0_c_484_n 4.84738e-19 $X=4.245 $Y=1.285 $X2=0 $Y2=0
cc_264 N_A_27_74#_c_226_n N_S0_c_484_n 0.0172982f $X=4.245 $Y=1.285 $X2=0 $Y2=0
cc_265 N_A_27_74#_c_227_n N_S0_c_484_n 0.00481074f $X=4.665 $Y=1.445 $X2=0 $Y2=0
cc_266 N_A_27_74#_c_229_n N_S0_c_484_n 0.00403701f $X=5.175 $Y=1.61 $X2=0 $Y2=0
cc_267 N_A_27_74#_c_237_n N_S0_c_484_n 9.49459e-19 $X=4.665 $Y=0.96 $X2=0 $Y2=0
cc_268 N_A_27_74#_c_238_n N_S0_c_484_n 8.87846e-19 $X=4.245 $Y=1.12 $X2=0 $Y2=0
cc_269 N_A_27_74#_c_219_n N_S0_c_485_n 0.00144141f $X=1.53 $Y=0.945 $X2=0 $Y2=0
cc_270 N_A_27_74#_c_245_n N_S0_c_485_n 0.00140016f $X=0.39 $Y=2.035 $X2=0 $Y2=0
cc_271 N_A_27_74#_c_219_n N_S0_c_486_n 0.0269006f $X=1.53 $Y=0.945 $X2=0 $Y2=0
cc_272 N_A_27_74#_c_245_n N_S0_c_486_n 0.00651637f $X=0.39 $Y=2.035 $X2=0 $Y2=0
cc_273 N_A_27_74#_c_232_n N_S0_c_486_n 0.0438201f $X=0.332 $Y=1.95 $X2=0 $Y2=0
cc_274 N_A_27_74#_c_229_n N_A3_c_601_n 2.34704e-19 $X=5.175 $Y=1.61 $X2=0 $Y2=0
cc_275 N_A_27_74#_c_230_n N_A3_c_601_n 0.0134856f $X=5.175 $Y=1.61 $X2=0 $Y2=0
cc_276 N_A_27_74#_M1005_g N_A3_c_602_n 0.06388f $X=5.25 $Y=2.435 $X2=0 $Y2=0
cc_277 N_A_27_74#_c_229_n N_A3_c_602_n 3.43922e-19 $X=5.175 $Y=1.61 $X2=0 $Y2=0
cc_278 N_A_27_74#_c_230_n N_A3_c_602_n 0.0157269f $X=5.175 $Y=1.61 $X2=0 $Y2=0
cc_279 N_A_27_74#_c_245_n N_VPWR_c_862_n 0.0381122f $X=0.39 $Y=2.035 $X2=0 $Y2=0
cc_280 N_A_27_74#_c_241_n N_VPWR_c_866_n 0.0139866f $X=0.39 $Y=2.715 $X2=0 $Y2=0
cc_281 N_A_27_74#_M1005_g N_VPWR_c_870_n 0.00113339f $X=5.25 $Y=2.435 $X2=0
+ $Y2=0
cc_282 N_A_27_74#_M1013_g N_VPWR_c_861_n 0.00113998f $X=2.61 $Y=2.205 $X2=0
+ $Y2=0
cc_283 N_A_27_74#_c_241_n N_VPWR_c_861_n 0.015197f $X=0.39 $Y=2.715 $X2=0 $Y2=0
cc_284 N_A_27_74#_c_220_n N_A_342_74#_M1015_d 0.00600069f $X=2.46 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_285 N_A_27_74#_M1013_g N_A_342_74#_c_970_n 0.00739494f $X=2.61 $Y=2.205 $X2=0
+ $Y2=0
cc_286 N_A_27_74#_M1013_g N_A_342_74#_c_971_n 0.0132149f $X=2.61 $Y=2.205 $X2=0
+ $Y2=0
cc_287 N_A_27_74#_M1005_g N_A_342_74#_c_959_n 0.0181045f $X=5.25 $Y=2.435 $X2=0
+ $Y2=0
cc_288 N_A_27_74#_M1015_g N_A_342_74#_c_953_n 0.00309442f $X=1.635 $Y=0.69 $X2=0
+ $Y2=0
cc_289 N_A_27_74#_c_308_p N_A_342_74#_c_953_n 0.0191397f $X=1.615 $Y=0.86 $X2=0
+ $Y2=0
cc_290 N_A_27_74#_c_220_n N_A_342_74#_c_953_n 0.0191354f $X=2.46 $Y=0.34 $X2=0
+ $Y2=0
cc_291 N_A_27_74#_c_260_p N_A_342_74#_c_953_n 0.0148708f $X=2.545 $Y=0.875 $X2=0
+ $Y2=0
cc_292 N_A_27_74#_c_342_p N_A_342_74#_c_953_n 0.0136961f $X=1.615 $Y=0.945 $X2=0
+ $Y2=0
cc_293 N_A_27_74#_c_236_n N_A_342_74#_c_953_n 0.00923031f $X=2.625 $Y=0.96 $X2=0
+ $Y2=0
cc_294 N_A_27_74#_M1013_g N_A_342_74#_c_965_n 0.00523363f $X=2.61 $Y=2.205 $X2=0
+ $Y2=0
cc_295 N_A_27_74#_c_222_n N_A_342_74#_c_965_n 0.00601104f $X=2.625 $Y=1.285
+ $X2=0 $Y2=0
cc_296 N_A_27_74#_c_223_n N_A_342_74#_c_965_n 4.48835e-19 $X=2.625 $Y=1.285
+ $X2=0 $Y2=0
cc_297 N_A_27_74#_M1015_g N_A_342_74#_c_954_n 0.00105664f $X=1.635 $Y=0.69 $X2=0
+ $Y2=0
cc_298 N_A_27_74#_M1013_g N_A_342_74#_c_954_n 0.00136529f $X=2.61 $Y=2.205 $X2=0
+ $Y2=0
cc_299 N_A_27_74#_c_222_n N_A_342_74#_c_954_n 0.0208345f $X=2.625 $Y=1.285 $X2=0
+ $Y2=0
cc_300 N_A_27_74#_c_223_n N_A_342_74#_c_954_n 0.00106957f $X=2.625 $Y=1.285
+ $X2=0 $Y2=0
cc_301 N_A_27_74#_c_233_n N_A_342_74#_c_954_n 0.0248017f $X=1.695 $Y=1.365 $X2=0
+ $Y2=0
cc_302 N_A_27_74#_c_234_n N_A_342_74#_c_954_n 0.00174016f $X=1.695 $Y=1.365
+ $X2=0 $Y2=0
cc_303 N_A_27_74#_c_235_n N_A_342_74#_c_954_n 0.00738764f $X=1.695 $Y=1.2 $X2=0
+ $Y2=0
cc_304 N_A_27_74#_c_236_n N_A_342_74#_c_954_n 8.82522e-19 $X=2.625 $Y=0.96 $X2=0
+ $Y2=0
cc_305 N_A_27_74#_M1013_g N_A_342_74#_c_967_n 0.00620023f $X=2.61 $Y=2.205 $X2=0
+ $Y2=0
cc_306 N_A_27_74#_c_237_n N_A_846_74#_M1022_d 0.00463813f $X=4.665 $Y=0.96
+ $X2=-0.19 $Y2=-0.245
cc_307 N_A_27_74#_c_237_n N_A_846_74#_c_1110_n 0.0324305f $X=4.665 $Y=0.96 $X2=0
+ $Y2=0
cc_308 N_A_27_74#_c_238_n N_A_846_74#_c_1110_n 0.0118221f $X=4.245 $Y=1.12 $X2=0
+ $Y2=0
cc_309 N_A_27_74#_c_227_n N_A_846_74#_c_1094_n 0.00421927f $X=4.665 $Y=1.445
+ $X2=0 $Y2=0
cc_310 N_A_27_74#_c_237_n N_A_846_74#_c_1094_n 0.00832361f $X=4.665 $Y=0.96
+ $X2=0 $Y2=0
cc_311 N_A_27_74#_c_229_n N_A_846_74#_c_1095_n 0.0187515f $X=5.175 $Y=1.61 $X2=0
+ $Y2=0
cc_312 N_A_27_74#_c_230_n N_A_846_74#_c_1095_n 0.00219571f $X=5.175 $Y=1.61
+ $X2=0 $Y2=0
cc_313 N_A_27_74#_c_227_n N_A_846_74#_c_1096_n 0.0136801f $X=4.665 $Y=1.445
+ $X2=0 $Y2=0
cc_314 N_A_27_74#_c_229_n N_A_846_74#_c_1096_n 0.0147082f $X=5.175 $Y=1.61 $X2=0
+ $Y2=0
cc_315 N_A_27_74#_c_230_n N_A_846_74#_c_1096_n 0.00186365f $X=5.175 $Y=1.61
+ $X2=0 $Y2=0
cc_316 N_A_27_74#_M1005_g N_A_846_74#_c_1119_n 0.0148921f $X=5.25 $Y=2.435 $X2=0
+ $Y2=0
cc_317 N_A_27_74#_c_229_n N_A_846_74#_c_1097_n 0.0262124f $X=5.175 $Y=1.61 $X2=0
+ $Y2=0
cc_318 N_A_27_74#_c_230_n N_A_846_74#_c_1097_n 0.00550326f $X=5.175 $Y=1.61
+ $X2=0 $Y2=0
cc_319 N_A_27_74#_M1005_g N_A_846_74#_c_1122_n 0.00947737f $X=5.25 $Y=2.435
+ $X2=0 $Y2=0
cc_320 N_A_27_74#_c_225_n N_A_846_74#_c_1122_n 0.00233591f $X=4.245 $Y=1.285
+ $X2=0 $Y2=0
cc_321 N_A_27_74#_c_228_n N_A_846_74#_c_1122_n 0.0120851f $X=4.75 $Y=1.61 $X2=0
+ $Y2=0
cc_322 N_A_27_74#_c_229_n N_A_846_74#_c_1122_n 0.0368437f $X=5.175 $Y=1.61 $X2=0
+ $Y2=0
cc_323 N_A_27_74#_c_230_n N_A_846_74#_c_1122_n 0.00320169f $X=5.175 $Y=1.61
+ $X2=0 $Y2=0
cc_324 N_A_27_74#_c_219_n N_VGND_M1021_d 0.00815441f $X=1.53 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_325 N_A_27_74#_c_224_n N_VGND_M1001_d 0.00613658f $X=4.08 $Y=0.96 $X2=0 $Y2=0
cc_326 N_A_27_74#_c_218_n N_VGND_c_1239_n 0.0190719f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_327 N_A_27_74#_c_219_n N_VGND_c_1239_n 0.0295177f $X=1.53 $Y=0.945 $X2=0
+ $Y2=0
cc_328 N_A_27_74#_c_221_n N_VGND_c_1239_n 0.00638964f $X=1.7 $Y=0.34 $X2=0 $Y2=0
cc_329 N_A_27_74#_c_220_n N_VGND_c_1240_n 0.00658648f $X=2.46 $Y=0.34 $X2=0
+ $Y2=0
cc_330 N_A_27_74#_c_260_p N_VGND_c_1240_n 0.00855501f $X=2.545 $Y=0.875 $X2=0
+ $Y2=0
cc_331 N_A_27_74#_c_224_n N_VGND_c_1240_n 0.0345611f $X=4.08 $Y=0.96 $X2=0 $Y2=0
cc_332 N_A_27_74#_c_238_n N_VGND_c_1240_n 0.00154479f $X=4.245 $Y=1.12 $X2=0
+ $Y2=0
cc_333 N_A_27_74#_M1015_g N_VGND_c_1245_n 0.00278135f $X=1.635 $Y=0.69 $X2=0
+ $Y2=0
cc_334 N_A_27_74#_c_220_n N_VGND_c_1245_n 0.0606235f $X=2.46 $Y=0.34 $X2=0 $Y2=0
cc_335 N_A_27_74#_c_221_n N_VGND_c_1245_n 0.0116947f $X=1.7 $Y=0.34 $X2=0 $Y2=0
cc_336 N_A_27_74#_c_238_n N_VGND_c_1246_n 0.00439269f $X=4.245 $Y=1.12 $X2=0
+ $Y2=0
cc_337 N_A_27_74#_M1015_g N_VGND_c_1248_n 0.00354157f $X=1.635 $Y=0.69 $X2=0
+ $Y2=0
cc_338 N_A_27_74#_c_218_n N_VGND_c_1248_n 0.012183f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_339 N_A_27_74#_c_219_n N_VGND_c_1248_n 0.0229194f $X=1.53 $Y=0.945 $X2=0
+ $Y2=0
cc_340 N_A_27_74#_c_220_n N_VGND_c_1248_n 0.034448f $X=2.46 $Y=0.34 $X2=0 $Y2=0
cc_341 N_A_27_74#_c_221_n N_VGND_c_1248_n 0.00596862f $X=1.7 $Y=0.34 $X2=0 $Y2=0
cc_342 N_A_27_74#_c_238_n N_VGND_c_1248_n 0.00837941f $X=4.245 $Y=1.12 $X2=0
+ $Y2=0
cc_343 N_A_27_74#_c_218_n N_VGND_c_1249_n 0.014787f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_344 N_A_27_74#_c_219_n A_264_74# 0.00257608f $X=1.53 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_345 N_A_27_74#_c_220_n A_450_74# 0.00722946f $X=2.46 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_346 N_A_27_74#_c_260_p A_450_74# 0.0152875f $X=2.545 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_347 N_A_27_74#_c_224_n A_450_74# 0.00590237f $X=4.08 $Y=0.96 $X2=-0.19
+ $Y2=-0.245
cc_348 N_A_27_74#_c_236_n A_450_74# 0.00963213f $X=2.625 $Y=0.96 $X2=-0.19
+ $Y2=-0.245
cc_349 N_A_27_74#_c_224_n A_768_74# 0.0048076f $X=4.08 $Y=0.96 $X2=-0.19
+ $Y2=-0.245
cc_350 N_A1_M1000_g N_A2_M1002_g 0.0328679f $X=3.12 $Y=2.205 $X2=0 $Y2=0
cc_351 N_A1_c_402_n N_A2_M1002_g 0.00167677f $X=3.165 $Y=1.38 $X2=0 $Y2=0
cc_352 N_A1_M1001_g N_A2_M1023_g 0.0203478f $X=3.075 $Y=0.69 $X2=0 $Y2=0
cc_353 N_A1_c_401_n N_A2_c_441_n 0.0206294f $X=3.165 $Y=1.38 $X2=0 $Y2=0
cc_354 N_A1_c_402_n N_A2_c_441_n 3.80681e-19 $X=3.165 $Y=1.38 $X2=0 $Y2=0
cc_355 N_A1_M1000_g N_A2_c_442_n 0.00182567f $X=3.12 $Y=2.205 $X2=0 $Y2=0
cc_356 N_A1_c_401_n N_A2_c_442_n 0.00188197f $X=3.165 $Y=1.38 $X2=0 $Y2=0
cc_357 N_A1_c_402_n N_A2_c_442_n 0.0757936f $X=3.165 $Y=1.38 $X2=0 $Y2=0
cc_358 N_A1_M1000_g N_S0_c_491_n 0.0103286f $X=3.12 $Y=2.205 $X2=0 $Y2=0
cc_359 N_A1_c_402_n N_VPWR_M1000_d 0.00474029f $X=3.165 $Y=1.38 $X2=0 $Y2=0
cc_360 N_A1_M1000_g N_VPWR_c_863_n 0.00398531f $X=3.12 $Y=2.205 $X2=0 $Y2=0
cc_361 N_A1_M1000_g N_VPWR_c_861_n 0.00113998f $X=3.12 $Y=2.205 $X2=0 $Y2=0
cc_362 N_A1_M1000_g N_A_342_74#_c_970_n 8.59113e-19 $X=3.12 $Y=2.205 $X2=0 $Y2=0
cc_363 N_A1_M1000_g N_A_342_74#_c_971_n 0.0121605f $X=3.12 $Y=2.205 $X2=0 $Y2=0
cc_364 N_A1_c_402_n N_A_342_74#_c_971_n 0.0175433f $X=3.165 $Y=1.38 $X2=0 $Y2=0
cc_365 N_A1_M1000_g N_A_342_74#_c_958_n 7.95693e-19 $X=3.12 $Y=2.205 $X2=0 $Y2=0
cc_366 N_A1_M1000_g N_A_342_74#_c_965_n 4.59945e-19 $X=3.12 $Y=2.205 $X2=0 $Y2=0
cc_367 N_A1_c_402_n N_A_342_74#_c_965_n 0.00888376f $X=3.165 $Y=1.38 $X2=0 $Y2=0
cc_368 N_A1_M1000_g N_A_342_74#_c_967_n 0.00109651f $X=3.12 $Y=2.205 $X2=0 $Y2=0
cc_369 N_A1_M1001_g N_VGND_c_1240_n 0.0174878f $X=3.075 $Y=0.69 $X2=0 $Y2=0
cc_370 N_A1_M1001_g N_VGND_c_1245_n 0.00383152f $X=3.075 $Y=0.69 $X2=0 $Y2=0
cc_371 N_A1_M1001_g N_VGND_c_1248_n 0.00762539f $X=3.075 $Y=0.69 $X2=0 $Y2=0
cc_372 N_A2_M1002_g N_S0_c_491_n 0.0102489f $X=3.74 $Y=2.205 $X2=0 $Y2=0
cc_373 N_A2_M1002_g N_S0_c_494_n 0.0405301f $X=3.74 $Y=2.205 $X2=0 $Y2=0
cc_374 N_A2_c_442_n N_S0_c_494_n 0.00188646f $X=3.705 $Y=1.38 $X2=0 $Y2=0
cc_375 N_A2_c_442_n N_VPWR_M1000_d 0.00505088f $X=3.705 $Y=1.38 $X2=0 $Y2=0
cc_376 N_A2_M1002_g N_VPWR_c_863_n 0.00151557f $X=3.74 $Y=2.205 $X2=0 $Y2=0
cc_377 N_A2_M1002_g N_VPWR_c_861_n 9.20984e-19 $X=3.74 $Y=2.205 $X2=0 $Y2=0
cc_378 N_A2_M1002_g N_A_342_74#_c_971_n 0.0111608f $X=3.74 $Y=2.205 $X2=0 $Y2=0
cc_379 N_A2_c_442_n N_A_342_74#_c_971_n 0.0200788f $X=3.705 $Y=1.38 $X2=0 $Y2=0
cc_380 N_A2_M1002_g N_A_342_74#_c_958_n 0.00903954f $X=3.74 $Y=2.205 $X2=0 $Y2=0
cc_381 N_A2_M1023_g N_A_846_74#_c_1110_n 9.6691e-19 $X=3.765 $Y=0.69 $X2=0 $Y2=0
cc_382 N_A2_M1002_g N_A_846_74#_c_1122_n 0.00133006f $X=3.74 $Y=2.205 $X2=0
+ $Y2=0
cc_383 N_A2_M1023_g N_VGND_c_1240_n 0.0165996f $X=3.765 $Y=0.69 $X2=0 $Y2=0
cc_384 N_A2_M1023_g N_VGND_c_1246_n 0.00383152f $X=3.765 $Y=0.69 $X2=0 $Y2=0
cc_385 N_A2_M1023_g N_VGND_c_1248_n 0.0075725f $X=3.765 $Y=0.69 $X2=0 $Y2=0
cc_386 N_S0_c_482_n N_A3_c_599_n 0.0237287f $X=4.82 $Y=1.085 $X2=-0.19
+ $Y2=-0.245
cc_387 N_S0_c_484_n N_A3_c_601_n 0.0237287f $X=4.82 $Y=1.16 $X2=0 $Y2=0
cc_388 N_S0_M1009_g N_VPWR_c_862_n 0.00963357f $X=0.615 $Y=2.34 $X2=0 $Y2=0
cc_389 N_S0_c_488_n N_VPWR_c_862_n 0.0239494f $X=2.07 $Y=3.15 $X2=0 $Y2=0
cc_390 N_S0_c_486_n N_VPWR_c_862_n 0.00680686f $X=0.615 $Y=1.38 $X2=0 $Y2=0
cc_391 N_S0_c_491_n N_VPWR_c_863_n 0.0253068f $X=4.155 $Y=3.15 $X2=0 $Y2=0
cc_392 N_S0_M1008_g N_VPWR_c_863_n 7.10911e-19 $X=4.245 $Y=2.435 $X2=0 $Y2=0
cc_393 N_S0_c_489_n N_VPWR_c_866_n 0.00739826f $X=0.705 $Y=3.15 $X2=0 $Y2=0
cc_394 N_S0_c_488_n N_VPWR_c_868_n 0.0735781f $X=2.07 $Y=3.15 $X2=0 $Y2=0
cc_395 N_S0_c_491_n N_VPWR_c_870_n 0.0188949f $X=4.155 $Y=3.15 $X2=0 $Y2=0
cc_396 N_S0_c_488_n N_VPWR_c_861_n 0.0517272f $X=2.07 $Y=3.15 $X2=0 $Y2=0
cc_397 N_S0_c_489_n N_VPWR_c_861_n 0.0118361f $X=0.705 $Y=3.15 $X2=0 $Y2=0
cc_398 N_S0_c_491_n N_VPWR_c_861_n 0.0496362f $X=4.155 $Y=3.15 $X2=0 $Y2=0
cc_399 N_S0_c_496_n N_VPWR_c_861_n 0.00508464f $X=2.16 $Y=3.15 $X2=0 $Y2=0
cc_400 N_S0_M1010_g N_A_342_74#_c_970_n 0.0122619f $X=2.16 $Y=2.205 $X2=0 $Y2=0
cc_401 N_S0_c_491_n N_A_342_74#_c_971_n 0.00881413f $X=4.155 $Y=3.15 $X2=0 $Y2=0
cc_402 N_S0_M1008_g N_A_342_74#_c_971_n 0.00161022f $X=4.245 $Y=2.435 $X2=0
+ $Y2=0
cc_403 N_S0_M1008_g N_A_342_74#_c_958_n 0.00686069f $X=4.245 $Y=2.435 $X2=0
+ $Y2=0
cc_404 N_S0_c_491_n N_A_342_74#_c_959_n 0.00105363f $X=4.155 $Y=3.15 $X2=0 $Y2=0
cc_405 N_S0_M1008_g N_A_342_74#_c_959_n 0.019036f $X=4.245 $Y=2.435 $X2=0 $Y2=0
cc_406 N_S0_c_491_n N_A_342_74#_c_960_n 0.00499425f $X=4.155 $Y=3.15 $X2=0 $Y2=0
cc_407 N_S0_c_479_n N_A_342_74#_c_953_n 2.58461e-19 $X=2.16 $Y=1.175 $X2=0 $Y2=0
cc_408 N_S0_c_483_n N_A_342_74#_c_953_n 0.0100031f $X=2.16 $Y=1.085 $X2=0 $Y2=0
cc_409 N_S0_M1010_g N_A_342_74#_c_965_n 0.0110299f $X=2.16 $Y=2.205 $X2=0 $Y2=0
cc_410 N_S0_c_479_n N_A_342_74#_c_954_n 0.00281389f $X=2.16 $Y=1.175 $X2=0 $Y2=0
cc_411 N_S0_M1010_g N_A_342_74#_c_954_n 0.0146683f $X=2.16 $Y=2.205 $X2=0 $Y2=0
cc_412 N_S0_c_483_n N_A_342_74#_c_954_n 0.00169124f $X=2.16 $Y=1.085 $X2=0 $Y2=0
cc_413 N_S0_M1010_g N_A_342_74#_c_967_n 0.0164897f $X=2.16 $Y=2.205 $X2=0 $Y2=0
cc_414 N_S0_c_491_n N_A_342_74#_c_967_n 0.00365848f $X=4.155 $Y=3.15 $X2=0 $Y2=0
cc_415 N_S0_c_482_n N_A_846_74#_c_1110_n 0.021291f $X=4.82 $Y=1.085 $X2=0 $Y2=0
cc_416 N_S0_c_482_n N_A_846_74#_c_1094_n 0.00186119f $X=4.82 $Y=1.085 $X2=0
+ $Y2=0
cc_417 N_S0_c_481_n N_A_846_74#_c_1096_n 8.31322e-19 $X=4.725 $Y=1.69 $X2=0
+ $Y2=0
cc_418 N_S0_c_484_n N_A_846_74#_c_1096_n 0.00110457f $X=4.82 $Y=1.16 $X2=0 $Y2=0
cc_419 N_S0_M1008_g N_A_846_74#_c_1122_n 0.0156011f $X=4.245 $Y=2.435 $X2=0
+ $Y2=0
cc_420 N_S0_c_493_n N_A_846_74#_c_1122_n 0.0142819f $X=4.65 $Y=1.765 $X2=0 $Y2=0
cc_421 N_S0_M1021_g N_VGND_c_1239_n 0.00676114f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_422 N_S0_c_482_n N_VGND_c_1241_n 0.00100982f $X=4.82 $Y=1.085 $X2=0 $Y2=0
cc_423 N_S0_c_483_n N_VGND_c_1245_n 0.00278271f $X=2.16 $Y=1.085 $X2=0 $Y2=0
cc_424 N_S0_c_482_n N_VGND_c_1246_n 0.00295004f $X=4.82 $Y=1.085 $X2=0 $Y2=0
cc_425 N_S0_M1021_g N_VGND_c_1248_n 0.00456213f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_426 N_S0_c_482_n N_VGND_c_1248_n 0.00363625f $X=4.82 $Y=1.085 $X2=0 $Y2=0
cc_427 N_S0_c_483_n N_VGND_c_1248_n 0.00359456f $X=2.16 $Y=1.085 $X2=0 $Y2=0
cc_428 N_S0_M1021_g N_VGND_c_1249_n 0.00434272f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_429 N_A3_c_602_n N_S1_M1004_g 0.0130295f $X=5.67 $Y=1.865 $X2=0 $Y2=0
cc_430 N_A3_c_602_n N_S1_M1007_g 0.00656387f $X=5.67 $Y=1.865 $X2=0 $Y2=0
cc_431 N_A3_c_602_n N_VPWR_c_864_n 0.00803321f $X=5.67 $Y=1.865 $X2=0 $Y2=0
cc_432 N_A3_c_602_n N_VPWR_c_870_n 0.00558361f $X=5.67 $Y=1.865 $X2=0 $Y2=0
cc_433 N_A3_c_602_n N_VPWR_c_861_n 0.00541439f $X=5.67 $Y=1.865 $X2=0 $Y2=0
cc_434 N_A3_c_602_n N_A_342_74#_c_959_n 0.00119995f $X=5.67 $Y=1.865 $X2=0 $Y2=0
cc_435 N_A3_c_602_n N_A_342_74#_c_961_n 0.0205301f $X=5.67 $Y=1.865 $X2=0 $Y2=0
cc_436 A3 N_A_342_74#_c_961_n 0.0111922f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_437 N_A3_c_602_n N_A_342_74#_c_963_n 0.00788538f $X=5.67 $Y=1.865 $X2=0 $Y2=0
cc_438 N_A3_c_602_n N_A_342_74#_c_964_n 0.00388244f $X=5.67 $Y=1.865 $X2=0 $Y2=0
cc_439 N_A3_c_602_n N_A_342_74#_c_955_n 0.0105151f $X=5.67 $Y=1.865 $X2=0 $Y2=0
cc_440 A3 N_A_342_74#_c_955_n 0.0204305f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_441 N_A3_c_599_n N_A_846_74#_c_1094_n 0.00337564f $X=5.21 $Y=1.085 $X2=0
+ $Y2=0
cc_442 N_A3_c_600_n N_A_846_74#_c_1095_n 0.00654084f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_443 N_A3_c_601_n N_A_846_74#_c_1095_n 0.00910877f $X=5.285 $Y=1.16 $X2=0
+ $Y2=0
cc_444 N_A3_c_602_n N_A_846_74#_c_1119_n 0.00780058f $X=5.67 $Y=1.865 $X2=0
+ $Y2=0
cc_445 N_A3_c_602_n N_A_846_74#_c_1097_n 0.0301535f $X=5.67 $Y=1.865 $X2=0 $Y2=0
cc_446 A3 N_A_846_74#_c_1097_n 0.0239436f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_447 N_A3_c_602_n N_A_846_74#_c_1098_n 0.0320376f $X=5.67 $Y=1.865 $X2=0 $Y2=0
cc_448 A3 N_A_846_74#_c_1098_n 0.0251382f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_449 N_A3_c_599_n N_A_846_74#_c_1099_n 6.44102e-19 $X=5.21 $Y=1.085 $X2=0
+ $Y2=0
cc_450 N_A3_c_602_n N_A_846_74#_c_1100_n 0.00621898f $X=5.67 $Y=1.865 $X2=0
+ $Y2=0
cc_451 N_A3_c_602_n N_A_846_74#_c_1122_n 9.56141e-19 $X=5.67 $Y=1.865 $X2=0
+ $Y2=0
cc_452 N_A3_c_600_n N_A_846_74#_c_1146_n 0.00473182f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_453 N_A3_c_602_n N_A_846_74#_c_1146_n 0.00509879f $X=5.67 $Y=1.865 $X2=0
+ $Y2=0
cc_454 N_A3_c_599_n N_VGND_c_1241_n 0.0114303f $X=5.21 $Y=1.085 $X2=0 $Y2=0
cc_455 N_A3_c_600_n N_VGND_c_1241_n 0.00601958f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_456 N_A3_c_599_n N_VGND_c_1246_n 0.00383152f $X=5.21 $Y=1.085 $X2=0 $Y2=0
cc_457 N_A3_c_599_n N_VGND_c_1248_n 0.0075725f $X=5.21 $Y=1.085 $X2=0 $Y2=0
cc_458 N_A_1396_99#_M1024_g N_S1_M1004_g 0.0214569f $X=7.055 $Y=0.945 $X2=0
+ $Y2=0
cc_459 N_A_1396_99#_M1006_g N_S1_M1007_g 0.0170074f $X=7.18 $Y=2.46 $X2=0 $Y2=0
cc_460 N_A_1396_99#_c_644_n N_S1_M1007_g 0.00743862f $X=7.125 $Y=1.515 $X2=0
+ $Y2=0
cc_461 N_A_1396_99#_M1024_g N_S1_c_706_n 0.00737233f $X=7.055 $Y=0.945 $X2=0
+ $Y2=0
cc_462 N_A_1396_99#_c_647_n N_S1_c_706_n 0.00919339f $X=8.245 $Y=0.665 $X2=0
+ $Y2=0
cc_463 N_A_1396_99#_c_645_n N_S1_c_708_n 0.00245034f $X=7.795 $Y=1.61 $X2=0
+ $Y2=0
cc_464 N_A_1396_99#_c_646_n N_S1_c_708_n 0.00350686f $X=7.832 $Y=1.445 $X2=0
+ $Y2=0
cc_465 N_A_1396_99#_c_647_n N_S1_c_708_n 0.00156332f $X=8.245 $Y=0.665 $X2=0
+ $Y2=0
cc_466 N_A_1396_99#_c_648_n N_S1_c_708_n 0.0171154f $X=7.795 $Y=1.515 $X2=0
+ $Y2=0
cc_467 N_A_1396_99#_c_652_n N_S1_M1016_g 0.00245034f $X=8.015 $Y=1.95 $X2=0
+ $Y2=0
cc_468 N_A_1396_99#_c_646_n N_S1_M1011_g 0.00337861f $X=7.832 $Y=1.445 $X2=0
+ $Y2=0
cc_469 N_A_1396_99#_c_647_n N_S1_M1011_g 0.00866907f $X=8.245 $Y=0.665 $X2=0
+ $Y2=0
cc_470 N_A_1396_99#_M1024_g N_S1_c_710_n 0.00743862f $X=7.055 $Y=0.945 $X2=0
+ $Y2=0
cc_471 N_A_1396_99#_c_646_n N_S1_c_711_n 0.0339526f $X=7.832 $Y=1.445 $X2=0
+ $Y2=0
cc_472 N_A_1396_99#_c_647_n N_S1_c_711_n 0.0174115f $X=8.245 $Y=0.665 $X2=0
+ $Y2=0
cc_473 N_A_1396_99#_c_648_n N_S1_c_711_n 3.6795e-19 $X=7.795 $Y=1.515 $X2=0
+ $Y2=0
cc_474 N_A_1396_99#_M1024_g N_A_1338_125#_c_782_n 0.00606704f $X=7.055 $Y=0.945
+ $X2=0 $Y2=0
cc_475 N_A_1396_99#_M1024_g N_A_1338_125#_c_783_n 0.00389469f $X=7.055 $Y=0.945
+ $X2=0 $Y2=0
cc_476 N_A_1396_99#_M1006_g N_A_1338_125#_c_783_n 0.025007f $X=7.18 $Y=2.46
+ $X2=0 $Y2=0
cc_477 N_A_1396_99#_c_644_n N_A_1338_125#_c_783_n 0.00782459f $X=7.125 $Y=1.515
+ $X2=0 $Y2=0
cc_478 N_A_1396_99#_M1016_s N_A_1338_125#_c_788_n 0.00314282f $X=7.87 $Y=1.935
+ $X2=0 $Y2=0
cc_479 N_A_1396_99#_M1006_g N_A_1338_125#_c_788_n 0.0137576f $X=7.18 $Y=2.46
+ $X2=0 $Y2=0
cc_480 N_A_1396_99#_c_650_n N_A_1338_125#_c_788_n 0.02228f $X=8.015 $Y=2.115
+ $X2=0 $Y2=0
cc_481 N_A_1396_99#_M1006_g N_A_1338_125#_c_789_n 0.00190737f $X=7.18 $Y=2.46
+ $X2=0 $Y2=0
cc_482 N_A_1396_99#_M1006_g N_VPWR_c_871_n 0.00333896f $X=7.18 $Y=2.46 $X2=0
+ $Y2=0
cc_483 N_A_1396_99#_M1006_g N_VPWR_c_861_n 0.00428385f $X=7.18 $Y=2.46 $X2=0
+ $Y2=0
cc_484 N_A_1396_99#_M1024_g N_A_342_74#_c_955_n 7.43538e-19 $X=7.055 $Y=0.945
+ $X2=0 $Y2=0
cc_485 N_A_1396_99#_M1024_g N_A_342_74#_c_956_n 0.00433321f $X=7.055 $Y=0.945
+ $X2=0 $Y2=0
cc_486 N_A_1396_99#_c_644_n N_A_342_74#_c_956_n 0.00418768f $X=7.125 $Y=1.515
+ $X2=0 $Y2=0
cc_487 N_A_1396_99#_M1024_g N_A_342_74#_c_957_n 0.00738537f $X=7.055 $Y=0.945
+ $X2=0 $Y2=0
cc_488 N_A_1396_99#_M1024_g N_A_846_74#_c_1101_n 0.00120987f $X=7.055 $Y=0.945
+ $X2=0 $Y2=0
cc_489 N_A_1396_99#_c_643_n N_A_846_74#_c_1107_n 0.00168494f $X=7.63 $Y=1.515
+ $X2=0 $Y2=0
cc_490 N_A_1396_99#_c_650_n N_A_846_74#_c_1107_n 0.0265879f $X=8.015 $Y=2.115
+ $X2=0 $Y2=0
cc_491 N_A_1396_99#_c_652_n N_A_846_74#_c_1107_n 0.0265879f $X=8.015 $Y=1.95
+ $X2=0 $Y2=0
cc_492 N_A_1396_99#_M1024_g N_A_846_74#_c_1102_n 0.00632515f $X=7.055 $Y=0.945
+ $X2=0 $Y2=0
cc_493 N_A_1396_99#_c_647_n N_A_846_74#_c_1102_n 0.0499511f $X=8.245 $Y=0.665
+ $X2=0 $Y2=0
cc_494 N_A_1396_99#_M1024_g N_A_846_74#_c_1104_n 0.00335241f $X=7.055 $Y=0.945
+ $X2=0 $Y2=0
cc_495 N_A_1396_99#_c_643_n N_A_846_74#_c_1104_n 0.00721105f $X=7.63 $Y=1.515
+ $X2=0 $Y2=0
cc_496 N_A_1396_99#_c_645_n N_A_846_74#_c_1104_n 0.00483371f $X=7.795 $Y=1.61
+ $X2=0 $Y2=0
cc_497 N_A_1396_99#_c_647_n N_A_846_74#_c_1104_n 0.0145371f $X=8.245 $Y=0.665
+ $X2=0 $Y2=0
cc_498 N_A_1396_99#_M1024_g N_A_846_74#_c_1105_n 0.00317042f $X=7.055 $Y=0.945
+ $X2=0 $Y2=0
cc_499 N_A_1396_99#_M1006_g N_A_846_74#_c_1105_n 0.00747972f $X=7.18 $Y=2.46
+ $X2=0 $Y2=0
cc_500 N_A_1396_99#_c_643_n N_A_846_74#_c_1105_n 0.0117865f $X=7.63 $Y=1.515
+ $X2=0 $Y2=0
cc_501 N_A_1396_99#_c_645_n N_A_846_74#_c_1105_n 0.024653f $X=7.795 $Y=1.61
+ $X2=0 $Y2=0
cc_502 N_A_1396_99#_c_646_n N_A_846_74#_c_1105_n 0.00697275f $X=7.832 $Y=1.445
+ $X2=0 $Y2=0
cc_503 N_A_1396_99#_c_652_n N_A_846_74#_c_1105_n 0.0074274f $X=8.015 $Y=1.95
+ $X2=0 $Y2=0
cc_504 N_A_1396_99#_c_648_n N_A_846_74#_c_1105_n 0.00132855f $X=7.795 $Y=1.515
+ $X2=0 $Y2=0
cc_505 N_A_1396_99#_c_647_n N_VGND_c_1242_n 0.0291305f $X=8.245 $Y=0.665 $X2=0
+ $Y2=0
cc_506 N_A_1396_99#_c_647_n N_VGND_c_1243_n 0.014939f $X=8.245 $Y=0.665 $X2=0
+ $Y2=0
cc_507 N_A_1396_99#_c_647_n N_VGND_c_1248_n 0.0159507f $X=8.245 $Y=0.665 $X2=0
+ $Y2=0
cc_508 N_S1_M1011_g N_A_1338_125#_M1017_g 0.0228209f $X=8.46 $Y=0.84 $X2=0 $Y2=0
cc_509 N_S1_c_708_n N_A_1338_125#_M1018_g 0.0130484f $X=8.29 $Y=1.77 $X2=0 $Y2=0
cc_510 N_S1_c_710_n N_A_1338_125#_c_782_n 0.00125953f $X=6.655 $Y=1.49 $X2=0
+ $Y2=0
cc_511 N_S1_M1004_g N_A_1338_125#_c_783_n 4.10822e-19 $X=6.615 $Y=0.945 $X2=0
+ $Y2=0
cc_512 N_S1_c_710_n N_A_1338_125#_c_783_n 0.00556483f $X=6.655 $Y=1.49 $X2=0
+ $Y2=0
cc_513 N_S1_M1016_g N_A_1338_125#_c_788_n 0.0176693f $X=8.29 $Y=2.435 $X2=0
+ $Y2=0
cc_514 N_S1_M1007_g N_A_1338_125#_c_789_n 0.003398f $X=6.68 $Y=2.46 $X2=0 $Y2=0
cc_515 N_S1_M1016_g N_A_1338_125#_c_808_n 0.0242179f $X=8.29 $Y=2.435 $X2=0
+ $Y2=0
cc_516 N_S1_c_711_n N_A_1338_125#_c_809_n 0.00108383f $X=8.37 $Y=1.515 $X2=0
+ $Y2=0
cc_517 N_S1_c_708_n N_A_1338_125#_c_810_n 7.09324e-19 $X=8.29 $Y=1.77 $X2=0
+ $Y2=0
cc_518 N_S1_M1016_g N_A_1338_125#_c_810_n 0.00562853f $X=8.29 $Y=2.435 $X2=0
+ $Y2=0
cc_519 N_S1_c_711_n N_A_1338_125#_c_810_n 0.0123177f $X=8.37 $Y=1.515 $X2=0
+ $Y2=0
cc_520 N_S1_c_708_n N_A_1338_125#_c_790_n 2.8046e-19 $X=8.29 $Y=1.77 $X2=0 $Y2=0
cc_521 N_S1_M1016_g N_A_1338_125#_c_790_n 0.00318956f $X=8.29 $Y=2.435 $X2=0
+ $Y2=0
cc_522 N_S1_c_708_n N_A_1338_125#_c_784_n 0.00114936f $X=8.29 $Y=1.77 $X2=0
+ $Y2=0
cc_523 N_S1_c_711_n N_A_1338_125#_c_784_n 0.0277175f $X=8.37 $Y=1.515 $X2=0
+ $Y2=0
cc_524 N_S1_c_708_n N_A_1338_125#_c_785_n 0.0205025f $X=8.29 $Y=1.77 $X2=0 $Y2=0
cc_525 N_S1_c_711_n N_A_1338_125#_c_785_n 0.00120518f $X=8.37 $Y=1.515 $X2=0
+ $Y2=0
cc_526 N_S1_M1007_g N_VPWR_c_864_n 0.00337872f $X=6.68 $Y=2.46 $X2=0 $Y2=0
cc_527 N_S1_M1016_g N_VPWR_c_865_n 0.00241293f $X=8.29 $Y=2.435 $X2=0 $Y2=0
cc_528 N_S1_M1007_g N_VPWR_c_871_n 0.005209f $X=6.68 $Y=2.46 $X2=0 $Y2=0
cc_529 N_S1_M1016_g N_VPWR_c_871_n 0.00115241f $X=8.29 $Y=2.435 $X2=0 $Y2=0
cc_530 N_S1_M1007_g N_VPWR_c_861_n 0.00989063f $X=6.68 $Y=2.46 $X2=0 $Y2=0
cc_531 N_S1_M1007_g N_A_342_74#_c_962_n 0.00245662f $X=6.68 $Y=2.46 $X2=0 $Y2=0
cc_532 N_S1_M1007_g N_A_342_74#_c_963_n 0.00354685f $X=6.68 $Y=2.46 $X2=0 $Y2=0
cc_533 N_S1_c_710_n N_A_342_74#_c_963_n 5.34817e-19 $X=6.655 $Y=1.49 $X2=0 $Y2=0
cc_534 N_S1_M1007_g N_A_342_74#_c_964_n 0.00600945f $X=6.68 $Y=2.46 $X2=0 $Y2=0
cc_535 N_S1_M1004_g N_A_342_74#_c_952_n 0.00397185f $X=6.615 $Y=0.945 $X2=0
+ $Y2=0
cc_536 N_S1_M1004_g N_A_342_74#_c_955_n 0.0146218f $X=6.615 $Y=0.945 $X2=0 $Y2=0
cc_537 N_S1_M1007_g N_A_342_74#_c_955_n 0.00724414f $X=6.68 $Y=2.46 $X2=0 $Y2=0
cc_538 N_S1_c_710_n N_A_342_74#_c_955_n 0.00422159f $X=6.655 $Y=1.49 $X2=0 $Y2=0
cc_539 N_S1_M1007_g N_A_342_74#_c_1035_n 0.00192359f $X=6.68 $Y=2.46 $X2=0 $Y2=0
cc_540 N_S1_M1004_g N_A_342_74#_c_956_n 4.65959e-19 $X=6.615 $Y=0.945 $X2=0
+ $Y2=0
cc_541 N_S1_M1004_g N_A_342_74#_c_957_n 0.0104485f $X=6.615 $Y=0.945 $X2=0 $Y2=0
cc_542 N_S1_c_710_n N_A_342_74#_c_957_n 9.14496e-19 $X=6.655 $Y=1.49 $X2=0 $Y2=0
cc_543 N_S1_M1004_g N_A_846_74#_c_1098_n 5.28281e-19 $X=6.615 $Y=0.945 $X2=0
+ $Y2=0
cc_544 N_S1_M1004_g N_A_846_74#_c_1100_n 0.00779557f $X=6.615 $Y=0.945 $X2=0
+ $Y2=0
cc_545 N_S1_M1004_g N_A_846_74#_c_1101_n 0.0137511f $X=6.615 $Y=0.945 $X2=0
+ $Y2=0
cc_546 N_S1_c_706_n N_A_846_74#_c_1101_n 0.0191695f $X=8.385 $Y=0.18 $X2=0 $Y2=0
cc_547 N_S1_M1011_g N_A_846_74#_c_1101_n 0.00409369f $X=8.46 $Y=0.84 $X2=0 $Y2=0
cc_548 N_S1_M1011_g N_A_846_74#_c_1102_n 0.00185502f $X=8.46 $Y=0.84 $X2=0 $Y2=0
cc_549 N_S1_M1004_g N_A_846_74#_c_1103_n 3.99719e-19 $X=6.615 $Y=0.945 $X2=0
+ $Y2=0
cc_550 N_S1_M1011_g N_A_846_74#_c_1104_n 7.07925e-19 $X=8.46 $Y=0.84 $X2=0 $Y2=0
cc_551 N_S1_c_706_n N_VGND_c_1242_n 0.0178023f $X=8.385 $Y=0.18 $X2=0 $Y2=0
cc_552 N_S1_c_707_n N_VGND_c_1243_n 0.0482304f $X=6.69 $Y=0.18 $X2=0 $Y2=0
cc_553 N_S1_c_706_n N_VGND_c_1248_n 0.0565635f $X=8.385 $Y=0.18 $X2=0 $Y2=0
cc_554 N_S1_c_707_n N_VGND_c_1248_n 0.00604685f $X=6.69 $Y=0.18 $X2=0 $Y2=0
cc_555 N_A_1338_125#_c_788_n N_VPWR_M1016_d 2.9285e-19 $X=8.35 $Y=2.99 $X2=0
+ $Y2=0
cc_556 N_A_1338_125#_c_808_n N_VPWR_M1016_d 0.00829346f $X=8.435 $Y=2.905 $X2=0
+ $Y2=0
cc_557 N_A_1338_125#_c_809_n N_VPWR_M1016_d 0.0219794f $X=8.745 $Y=2.035 $X2=0
+ $Y2=0
cc_558 N_A_1338_125#_c_810_n N_VPWR_M1016_d 7.49093e-19 $X=8.52 $Y=2.035 $X2=0
+ $Y2=0
cc_559 N_A_1338_125#_c_790_n N_VPWR_M1016_d 0.00347934f $X=8.83 $Y=1.95 $X2=0
+ $Y2=0
cc_560 N_A_1338_125#_M1018_g N_VPWR_c_865_n 0.0199952f $X=9.08 $Y=2.4 $X2=0
+ $Y2=0
cc_561 N_A_1338_125#_c_788_n N_VPWR_c_865_n 0.0149386f $X=8.35 $Y=2.99 $X2=0
+ $Y2=0
cc_562 N_A_1338_125#_c_808_n N_VPWR_c_865_n 0.0469629f $X=8.435 $Y=2.905 $X2=0
+ $Y2=0
cc_563 N_A_1338_125#_c_809_n N_VPWR_c_865_n 0.0195942f $X=8.745 $Y=2.035 $X2=0
+ $Y2=0
cc_564 N_A_1338_125#_c_784_n N_VPWR_c_865_n 0.00207826f $X=8.91 $Y=1.515 $X2=0
+ $Y2=0
cc_565 N_A_1338_125#_c_785_n N_VPWR_c_865_n 7.7246e-19 $X=9.08 $Y=1.515 $X2=0
+ $Y2=0
cc_566 N_A_1338_125#_c_788_n N_VPWR_c_871_n 0.0909292f $X=8.35 $Y=2.99 $X2=0
+ $Y2=0
cc_567 N_A_1338_125#_c_789_n N_VPWR_c_871_n 0.0234823f $X=7.12 $Y=2.99 $X2=0
+ $Y2=0
cc_568 N_A_1338_125#_M1018_g N_VPWR_c_872_n 0.00460063f $X=9.08 $Y=2.4 $X2=0
+ $Y2=0
cc_569 N_A_1338_125#_M1018_g N_VPWR_c_861_n 0.00912347f $X=9.08 $Y=2.4 $X2=0
+ $Y2=0
cc_570 N_A_1338_125#_c_788_n N_VPWR_c_861_n 0.0521645f $X=8.35 $Y=2.99 $X2=0
+ $Y2=0
cc_571 N_A_1338_125#_c_789_n N_VPWR_c_861_n 0.0126824f $X=7.12 $Y=2.99 $X2=0
+ $Y2=0
cc_572 N_A_1338_125#_c_783_n N_A_342_74#_c_963_n 0.0147455f $X=6.955 $Y=2.105
+ $X2=0 $Y2=0
cc_573 N_A_1338_125#_c_789_n N_A_342_74#_c_964_n 0.0037133f $X=7.12 $Y=2.99
+ $X2=0 $Y2=0
cc_574 N_A_1338_125#_c_782_n N_A_342_74#_c_955_n 0.0120468f $X=6.955 $Y=1.285
+ $X2=0 $Y2=0
cc_575 N_A_1338_125#_c_783_n N_A_342_74#_c_955_n 0.043798f $X=6.955 $Y=2.105
+ $X2=0 $Y2=0
cc_576 N_A_1338_125#_c_782_n N_A_342_74#_c_956_n 0.00114341f $X=6.955 $Y=1.285
+ $X2=0 $Y2=0
cc_577 N_A_1338_125#_M1004_d N_A_342_74#_c_957_n 0.00184734f $X=6.69 $Y=0.625
+ $X2=0 $Y2=0
cc_578 N_A_1338_125#_c_782_n N_A_342_74#_c_957_n 0.019663f $X=6.955 $Y=1.285
+ $X2=0 $Y2=0
cc_579 N_A_1338_125#_c_788_n N_A_846_74#_M1006_d 0.00335038f $X=8.35 $Y=2.99
+ $X2=0 $Y2=0
cc_580 N_A_1338_125#_c_788_n N_A_846_74#_c_1107_n 0.02228f $X=8.35 $Y=2.99 $X2=0
+ $Y2=0
cc_581 N_A_1338_125#_c_782_n N_A_846_74#_c_1104_n 0.0127985f $X=6.955 $Y=1.285
+ $X2=0 $Y2=0
cc_582 N_A_1338_125#_c_782_n N_A_846_74#_c_1105_n 7.62674e-19 $X=6.955 $Y=1.285
+ $X2=0 $Y2=0
cc_583 N_A_1338_125#_c_783_n N_A_846_74#_c_1105_n 0.0791124f $X=6.955 $Y=2.105
+ $X2=0 $Y2=0
cc_584 N_A_1338_125#_M1017_g X 0.00790145f $X=9.03 $Y=0.79 $X2=0 $Y2=0
cc_585 N_A_1338_125#_M1017_g X 0.00373467f $X=9.03 $Y=0.79 $X2=0 $Y2=0
cc_586 N_A_1338_125#_c_785_n X 0.00314505f $X=9.08 $Y=1.515 $X2=0 $Y2=0
cc_587 N_A_1338_125#_M1017_g X 0.00622745f $X=9.03 $Y=0.79 $X2=0 $Y2=0
cc_588 N_A_1338_125#_c_809_n X 0.00854274f $X=8.745 $Y=2.035 $X2=0 $Y2=0
cc_589 N_A_1338_125#_c_790_n X 0.0127776f $X=8.83 $Y=1.95 $X2=0 $Y2=0
cc_590 N_A_1338_125#_c_784_n X 0.0254663f $X=8.91 $Y=1.515 $X2=0 $Y2=0
cc_591 N_A_1338_125#_c_785_n X 0.0322073f $X=9.08 $Y=1.515 $X2=0 $Y2=0
cc_592 N_A_1338_125#_M1017_g N_VGND_c_1242_n 0.00807764f $X=9.03 $Y=0.79 $X2=0
+ $Y2=0
cc_593 N_A_1338_125#_c_784_n N_VGND_c_1242_n 0.0145322f $X=8.91 $Y=1.515 $X2=0
+ $Y2=0
cc_594 N_A_1338_125#_c_785_n N_VGND_c_1242_n 0.0012901f $X=9.08 $Y=1.515 $X2=0
+ $Y2=0
cc_595 N_A_1338_125#_M1017_g N_VGND_c_1247_n 0.00517302f $X=9.03 $Y=0.79 $X2=0
+ $Y2=0
cc_596 N_A_1338_125#_M1017_g N_VGND_c_1248_n 0.00529924f $X=9.03 $Y=0.79 $X2=0
+ $Y2=0
cc_597 N_VPWR_M1000_d N_A_342_74#_c_971_n 0.0121013f $X=3.21 $Y=1.705 $X2=0
+ $Y2=0
cc_598 N_VPWR_c_863_n N_A_342_74#_c_971_n 0.0259076f $X=3.43 $Y=2.84 $X2=0 $Y2=0
cc_599 N_VPWR_c_861_n N_A_342_74#_c_971_n 0.0280744f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_600 N_VPWR_c_863_n N_A_342_74#_c_958_n 0.0147765f $X=3.43 $Y=2.84 $X2=0 $Y2=0
cc_601 N_VPWR_c_864_n N_A_342_74#_c_959_n 0.0123841f $X=5.895 $Y=2.775 $X2=0
+ $Y2=0
cc_602 N_VPWR_c_870_n N_A_342_74#_c_959_n 0.0994305f $X=5.73 $Y=3.33 $X2=0 $Y2=0
cc_603 N_VPWR_c_861_n N_A_342_74#_c_959_n 0.056386f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_604 N_VPWR_c_863_n N_A_342_74#_c_960_n 0.013408f $X=3.43 $Y=2.84 $X2=0 $Y2=0
cc_605 N_VPWR_c_870_n N_A_342_74#_c_960_n 0.0153388f $X=5.73 $Y=3.33 $X2=0 $Y2=0
cc_606 N_VPWR_c_861_n N_A_342_74#_c_960_n 0.00771797f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_607 N_VPWR_M1012_d N_A_342_74#_c_961_n 0.0069031f $X=5.76 $Y=1.935 $X2=0
+ $Y2=0
cc_608 N_VPWR_c_864_n N_A_342_74#_c_961_n 0.0214055f $X=5.895 $Y=2.775 $X2=0
+ $Y2=0
cc_609 N_VPWR_c_861_n N_A_342_74#_c_961_n 0.0149483f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_610 N_VPWR_c_864_n N_A_342_74#_c_964_n 0.0205626f $X=5.895 $Y=2.775 $X2=0
+ $Y2=0
cc_611 N_VPWR_c_871_n N_A_342_74#_c_964_n 0.014549f $X=8.69 $Y=3.33 $X2=0 $Y2=0
cc_612 N_VPWR_c_861_n N_A_342_74#_c_964_n 0.0119743f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_613 N_VPWR_c_868_n N_A_342_74#_c_967_n 0.0106786f $X=3.265 $Y=3.33 $X2=0
+ $Y2=0
cc_614 N_VPWR_c_861_n N_A_342_74#_c_967_n 0.013737f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_615 N_VPWR_c_865_n X 0.0164587f $X=8.855 $Y=2.455 $X2=0 $Y2=0
cc_616 N_VPWR_c_872_n X 0.0082217f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_617 N_VPWR_c_861_n X 0.0091476f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_618 N_A_342_74#_c_971_n A_540_341# 0.0100794f $X=3.795 $Y=2.42 $X2=-0.19
+ $Y2=-0.245
cc_619 N_A_342_74#_c_971_n A_766_341# 0.00789917f $X=3.795 $Y=2.42 $X2=-0.19
+ $Y2=-0.245
cc_620 N_A_342_74#_c_958_n A_766_341# 0.00444759f $X=3.907 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_621 N_A_342_74#_c_959_n A_766_341# 0.00293798f $X=5.35 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_622 N_A_342_74#_c_952_n N_A_846_74#_M1004_s 0.00252297f $X=6.575 $Y=0.7 $X2=0
+ $Y2=0
cc_623 N_A_342_74#_c_955_n N_A_846_74#_M1004_s 0.00471995f $X=6.455 $Y=1.95
+ $X2=0 $Y2=0
cc_624 N_A_342_74#_c_959_n N_A_846_74#_M1008_d 0.00832289f $X=5.35 $Y=2.99 $X2=0
+ $Y2=0
cc_625 N_A_342_74#_c_961_n N_A_846_74#_c_1119_n 0.0075754f $X=6.29 $Y=2.42 $X2=0
+ $Y2=0
cc_626 N_A_342_74#_c_1072_p N_A_846_74#_c_1119_n 0.0102841f $X=5.55 $Y=2.42
+ $X2=0 $Y2=0
cc_627 N_A_342_74#_c_963_n N_A_846_74#_c_1119_n 0.00536899f $X=6.455 $Y=2.115
+ $X2=0 $Y2=0
cc_628 N_A_342_74#_c_963_n N_A_846_74#_c_1097_n 0.00128656f $X=6.455 $Y=2.115
+ $X2=0 $Y2=0
cc_629 N_A_342_74#_c_955_n N_A_846_74#_c_1098_n 0.0141439f $X=6.455 $Y=1.95
+ $X2=0 $Y2=0
cc_630 N_A_342_74#_c_952_n N_A_846_74#_c_1100_n 0.0141996f $X=6.575 $Y=0.7 $X2=0
+ $Y2=0
cc_631 N_A_342_74#_c_955_n N_A_846_74#_c_1100_n 0.0240517f $X=6.455 $Y=1.95
+ $X2=0 $Y2=0
cc_632 N_A_342_74#_c_952_n N_A_846_74#_c_1101_n 0.00649084f $X=6.575 $Y=0.7
+ $X2=0 $Y2=0
cc_633 N_A_342_74#_c_956_n N_A_846_74#_c_1101_n 0.0185392f $X=7.27 $Y=0.77 $X2=0
+ $Y2=0
cc_634 N_A_342_74#_c_957_n N_A_846_74#_c_1101_n 0.034646f $X=7.105 $Y=0.77 $X2=0
+ $Y2=0
cc_635 N_A_342_74#_c_956_n N_A_846_74#_c_1102_n 0.0261742f $X=7.27 $Y=0.77 $X2=0
+ $Y2=0
cc_636 N_A_342_74#_c_971_n N_A_846_74#_c_1122_n 0.00996195f $X=3.795 $Y=2.42
+ $X2=0 $Y2=0
cc_637 N_A_342_74#_c_958_n N_A_846_74#_c_1122_n 0.0122884f $X=3.907 $Y=2.905
+ $X2=0 $Y2=0
cc_638 N_A_342_74#_c_959_n N_A_846_74#_c_1122_n 0.0562506f $X=5.35 $Y=2.99 $X2=0
+ $Y2=0
cc_639 N_A_342_74#_c_952_n N_A_846_74#_c_1103_n 0.00619865f $X=6.575 $Y=0.7
+ $X2=0 $Y2=0
cc_640 N_A_342_74#_M1024_d N_A_846_74#_c_1104_n 0.00425603f $X=7.13 $Y=0.625
+ $X2=0 $Y2=0
cc_641 N_A_342_74#_c_956_n N_A_846_74#_c_1104_n 0.00496742f $X=7.27 $Y=0.77
+ $X2=0 $Y2=0
cc_642 N_A_342_74#_c_1088_p A_1068_387# 3.52028e-19 $X=5.45 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_643 N_A_342_74#_c_1072_p A_1068_387# 0.00141309f $X=5.55 $Y=2.42 $X2=-0.19
+ $Y2=-0.245
cc_644 N_A_846_74#_c_1119_n A_1068_387# 0.0055968f $X=5.51 $Y=2.08 $X2=-0.19
+ $Y2=-0.245
cc_645 N_A_846_74#_c_1097_n A_1068_387# 6.84302e-19 $X=5.595 $Y=1.995 $X2=-0.19
+ $Y2=-0.245
cc_646 N_A_846_74#_c_1110_n N_VGND_c_1240_n 0.0105681f $X=4.92 $Y=0.54 $X2=0
+ $Y2=0
cc_647 N_A_846_74#_c_1095_n N_VGND_c_1241_n 0.0169193f $X=5.51 $Y=1.19 $X2=0
+ $Y2=0
cc_648 N_A_846_74#_c_1099_n N_VGND_c_1241_n 0.00886151f $X=6.11 $Y=0.445 $X2=0
+ $Y2=0
cc_649 N_A_846_74#_c_1100_n N_VGND_c_1241_n 0.0222988f $X=6.15 $Y=0.82 $X2=0
+ $Y2=0
cc_650 N_A_846_74#_c_1146_n N_VGND_c_1241_n 0.00693814f $X=5.595 $Y=1.19 $X2=0
+ $Y2=0
cc_651 N_A_846_74#_c_1099_n N_VGND_c_1243_n 0.0165298f $X=6.11 $Y=0.445 $X2=0
+ $Y2=0
cc_652 N_A_846_74#_c_1206_p N_VGND_c_1243_n 0.0774851f $X=6.395 $Y=0.355 $X2=0
+ $Y2=0
cc_653 N_A_846_74#_c_1101_n N_VGND_c_1243_n 0.0114574f $X=7.525 $Y=0.35 $X2=0
+ $Y2=0
cc_654 N_A_846_74#_c_1110_n N_VGND_c_1246_n 0.0298469f $X=4.92 $Y=0.54 $X2=0
+ $Y2=0
cc_655 N_A_846_74#_M1004_s N_VGND_c_1248_n 0.00415243f $X=5.995 $Y=0.215 $X2=0
+ $Y2=0
cc_656 N_A_846_74#_c_1110_n N_VGND_c_1248_n 0.0305311f $X=4.92 $Y=0.54 $X2=0
+ $Y2=0
cc_657 N_A_846_74#_c_1099_n N_VGND_c_1248_n 0.00967329f $X=6.11 $Y=0.445 $X2=0
+ $Y2=0
cc_658 N_A_846_74#_c_1206_p N_VGND_c_1248_n 0.0441596f $X=6.395 $Y=0.355 $X2=0
+ $Y2=0
cc_659 N_A_846_74#_c_1101_n N_VGND_c_1248_n 0.00589978f $X=7.525 $Y=0.35 $X2=0
+ $Y2=0
cc_660 N_A_846_74#_c_1110_n A_979_74# 0.00161992f $X=4.92 $Y=0.54 $X2=-0.19
+ $Y2=-0.245
cc_661 N_A_846_74#_c_1094_n A_979_74# 3.36419e-19 $X=5.005 $Y=1.105 $X2=-0.19
+ $Y2=-0.245
cc_662 X N_VGND_c_1242_n 0.0317414f $X=9.275 $Y=0.47 $X2=0 $Y2=0
cc_663 X N_VGND_c_1247_n 0.014899f $X=9.275 $Y=0.47 $X2=0 $Y2=0
cc_664 X N_VGND_c_1248_n 0.014405f $X=9.275 $Y=0.47 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__dfstp_1.spice
* Created: Fri Aug 28 17:24:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dfstp_1.pex.spice"
.subckt sky130_fd_sc_ms__dfstp_1  VNB VPB D CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* D	D
* VPB	VPB
* VNB	VNB
MM1028 N_VGND_M1028_d N_D_M1028_g N_A_27_74#_M1028_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1031 N_VGND_M1031_d N_CLK_M1031_g N_A_224_350#_M1031_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1020 N_A_398_74#_M1020_d N_A_224_350#_M1020_g N_VGND_M1031_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1013 N_A_604_74#_M1013_d N_A_224_350#_M1013_g N_A_27_74#_M1013_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.17595 PD=0.95 PS=1.76 NRD=71.424 NRS=24.276 M=1
+ R=2.8 SA=75000.3 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1024 A_740_74# N_A_398_74#_M1024_g N_A_604_74#_M1013_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.1113 PD=0.66 PS=0.95 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_A_760_395#_M1022_g A_740_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1449 AS=0.0504 PD=1.53 PS=0.66 NRD=8.568 NRS=18.564 M=1 R=2.8 SA=75001.3
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1011 A_1027_118# N_A_604_74#_M1011_g N_A_760_395#_M1011_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1176 PD=0.63 PS=1.4 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_SET_B_M1009_g A_1027_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0964019 AS=0.0441 PD=0.847925 PS=0.63 NRD=43.56 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1003 A_1215_74# N_A_604_74#_M1003_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.12 AS=0.146898 PD=1.015 PS=1.29208 NRD=24.84 NRS=0 M=1 R=4.26667
+ SA=75000.8 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1007 N_A_1301_392#_M1007_d N_A_398_74#_M1007_g A_1215_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.129147 AS=0.12 PD=1.20755 PS=1.015 NRD=0 NRS=24.84 M=1 R=4.26667
+ SA=75001.3 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1018 A_1422_74# N_A_224_350#_M1018_g N_A_1301_392#_M1007_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0847528 PD=0.66 PS=0.792453 NRD=18.564 NRS=24.276 M=1
+ R=2.8 SA=75001.7 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1019 A_1500_74# N_A_1470_48#_M1019_g A_1422_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75002.1
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_SET_B_M1023_g A_1500_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.19215 AS=0.0504 PD=1.335 PS=0.66 NRD=1.428 NRS=18.564 M=1 R=2.8
+ SA=75002.5 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1005 N_A_1470_48#_M1005_d N_A_1301_392#_M1005_g N_VGND_M1023_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1197 AS=0.19215 PD=1.41 PS=1.335 NRD=0 NRS=19.992 M=1 R=2.8
+ SA=75003.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_A_1301_392#_M1026_g N_A_1902_74#_M1026_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.129591 AS=0.15675 PD=0.997674 PS=1.67 NRD=17.988 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1014 N_Q_M1014_d N_A_1902_74#_M1014_g N_VGND_M1026_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VPWR_M1008_d N_D_M1008_g N_A_27_74#_M1008_s VPB PSHORT L=0.18 W=0.42
+ AD=0.1113 AS=0.1134 PD=1.37 PS=1.38 NRD=0 NRS=0 M=1 R=2.33333 SA=90000.2
+ SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1004 N_VPWR_M1004_d N_CLK_M1004_g N_A_224_350#_M1004_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3024 PD=1.39 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1010 N_A_398_74#_M1010_d N_A_224_350#_M1010_g N_VPWR_M1004_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1017 N_A_604_74#_M1017_d N_A_398_74#_M1017_g N_A_27_74#_M1017_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0672 AS=0.1176 PD=0.74 PS=1.4 NRD=21.0987 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90004.2 A=0.0756 P=1.2 MULT=1
MM1015 A_712_463# N_A_224_350#_M1015_g N_A_604_74#_M1017_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0672 PD=0.66 PS=0.74 NRD=30.4759 NRS=0 M=1 R=2.33333
+ SA=90000.7 SB=90003.7 A=0.0756 P=1.2 MULT=1
MM1030 N_VPWR_M1030_d N_A_760_395#_M1030_g A_712_463# VPB PSHORT L=0.18 W=0.42
+ AD=0.13545 AS=0.0504 PD=1.065 PS=0.66 NRD=4.6886 NRS=30.4759 M=1 R=2.33333
+ SA=90001.1 SB=90003.3 A=0.0756 P=1.2 MULT=1
MM1000 N_A_760_395#_M1000_d N_A_604_74#_M1000_g N_VPWR_M1030_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0567 AS=0.13545 PD=0.69 PS=1.065 NRD=0 NRS=166.504 M=1 R=2.33333
+ SA=90001.9 SB=90002.5 A=0.0756 P=1.2 MULT=1
MM1012 N_VPWR_M1012_d N_SET_B_M1012_g N_A_760_395#_M1000_d VPB PSHORT L=0.18
+ W=0.42 AD=0.133394 AS=0.0567 PD=1.08254 PS=0.69 NRD=123.164 NRS=0 M=1
+ R=2.33333 SA=90002.4 SB=90002 A=0.0756 P=1.2 MULT=1
MM1001 A_1200_341# N_A_604_74#_M1001_g N_VPWR_M1012_d VPB PSHORT L=0.18 W=1
+ AD=0.184812 AS=0.317606 PD=1.58 PS=2.57746 NRD=25.5706 NRS=51.7322 M=1
+ R=5.55556 SA=90001.3 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1021 N_A_1301_392#_M1021_d N_A_224_350#_M1021_g A_1200_341# VPB PSHORT L=0.18
+ W=1 AD=0.290141 AS=0.184812 PD=2.27465 PS=1.58 NRD=0 NRS=25.5706 M=1 R=5.55556
+ SA=90001.7 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1027 A_1460_508# N_A_398_74#_M1027_g N_A_1301_392#_M1021_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.121859 PD=0.66 PS=0.955352 NRD=30.4759 NRS=79.7259 M=1
+ R=2.33333 SA=90002.3 SB=90001 A=0.0756 P=1.2 MULT=1
MM1002 N_VPWR_M1002_d N_A_1470_48#_M1002_g A_1460_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.0567 AS=0.0504 PD=0.69 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.33333 SA=90002.7
+ SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1006 N_A_1301_392#_M1006_d N_SET_B_M1006_g N_VPWR_M1002_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90003.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1016 N_A_1470_48#_M1016_d N_A_1301_392#_M1016_g N_VPWR_M1016_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.1092 AS=0.1113 PD=1.36 PS=1.37 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1029 N_VPWR_M1029_d N_A_1301_392#_M1029_g N_A_1902_74#_M1029_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1542 AS=0.2184 PD=1.25143 PS=2.2 NRD=30.4759 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1025 N_Q_M1025_d N_A_1902_74#_M1025_g N_VPWR_M1029_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3024 AS=0.2056 PD=2.78 PS=1.66857 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX32_noxref VNB VPB NWDIODE A=21.7821 P=26.83
c_1633 A_1200_341# 0 1.09525e-19 $X=6 $Y=1.705
*
.include "sky130_fd_sc_ms__dfstp_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__and3b_1.pxi.spice
* Created: Wed Sep  2 11:57:57 2020
* 
x_PM_SKY130_FD_SC_MS__AND3B_1%A_N N_A_N_M1006_g N_A_N_c_75_n N_A_N_M1002_g
+ N_A_N_c_71_n N_A_N_c_72_n N_A_N_c_77_n A_N A_N N_A_N_c_73_n N_A_N_c_74_n
+ PM_SKY130_FD_SC_MS__AND3B_1%A_N
x_PM_SKY130_FD_SC_MS__AND3B_1%A_114_74# N_A_114_74#_M1006_d N_A_114_74#_M1002_d
+ N_A_114_74#_c_101_n N_A_114_74#_M1009_g N_A_114_74#_c_103_n
+ N_A_114_74#_M1004_g N_A_114_74#_c_104_n N_A_114_74#_c_105_n
+ N_A_114_74#_c_111_n N_A_114_74#_c_106_n N_A_114_74#_c_107_n
+ N_A_114_74#_c_108_n N_A_114_74#_c_113_n N_A_114_74#_c_109_n
+ PM_SKY130_FD_SC_MS__AND3B_1%A_114_74#
x_PM_SKY130_FD_SC_MS__AND3B_1%B N_B_M1005_g N_B_M1000_g B N_B_c_168_n
+ N_B_c_171_n PM_SKY130_FD_SC_MS__AND3B_1%B
x_PM_SKY130_FD_SC_MS__AND3B_1%C N_C_M1007_g N_C_M1008_g C N_C_c_204_n
+ N_C_c_205_n PM_SKY130_FD_SC_MS__AND3B_1%C
x_PM_SKY130_FD_SC_MS__AND3B_1%A_266_94# N_A_266_94#_M1004_s N_A_266_94#_M1009_s
+ N_A_266_94#_M1000_d N_A_266_94#_M1001_g N_A_266_94#_M1003_g
+ N_A_266_94#_c_239_n N_A_266_94#_c_240_n N_A_266_94#_c_241_n
+ N_A_266_94#_c_259_n N_A_266_94#_c_242_n N_A_266_94#_c_246_n
+ N_A_266_94#_c_247_n N_A_266_94#_c_243_n PM_SKY130_FD_SC_MS__AND3B_1%A_266_94#
x_PM_SKY130_FD_SC_MS__AND3B_1%VPWR N_VPWR_M1002_s N_VPWR_M1009_d N_VPWR_M1008_d
+ N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_334_n N_VPWR_c_335_n N_VPWR_c_336_n
+ N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n VPWR N_VPWR_c_340_n
+ N_VPWR_c_331_n PM_SKY130_FD_SC_MS__AND3B_1%VPWR
x_PM_SKY130_FD_SC_MS__AND3B_1%X N_X_M1003_d N_X_M1001_d N_X_c_377_n N_X_c_378_n
+ X X X X N_X_c_381_n N_X_c_379_n PM_SKY130_FD_SC_MS__AND3B_1%X
x_PM_SKY130_FD_SC_MS__AND3B_1%VGND N_VGND_M1006_s N_VGND_M1007_d N_VGND_c_402_n
+ N_VGND_c_403_n N_VGND_c_404_n VGND N_VGND_c_405_n N_VGND_c_406_n
+ N_VGND_c_407_n N_VGND_c_408_n PM_SKY130_FD_SC_MS__AND3B_1%VGND
cc_1 VNB N_A_N_M1006_g 0.0315936f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_2 VNB N_A_N_c_71_n 0.0275245f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_3 VNB N_A_N_c_72_n 0.0036645f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.78
cc_4 VNB N_A_N_c_73_n 0.0185743f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.275
cc_5 VNB N_A_N_c_74_n 0.0240162f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.275
cc_6 VNB N_A_114_74#_c_101_n 0.0344902f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.54
cc_7 VNB N_A_114_74#_M1009_g 0.0129028f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.78
cc_8 VNB N_A_114_74#_c_103_n 0.0161108f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_9 VNB N_A_114_74#_c_104_n 0.0107445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_114_74#_c_105_n 0.00839405f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.275
cc_11 VNB N_A_114_74#_c_106_n 0.0205614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_114_74#_c_107_n 0.00199474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_114_74#_c_108_n 0.0493999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_114_74#_c_109_n 9.31753e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_M1005_g 0.0236487f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_16 VNB N_B_c_168_n 0.0258546f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_17 VNB N_C_M1007_g 0.0263528f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_18 VNB N_C_c_204_n 0.023996f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_19 VNB N_C_c_205_n 0.00189186f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.78
cc_20 VNB N_A_266_94#_M1001_g 0.00182608f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.615
cc_21 VNB N_A_266_94#_M1003_g 0.0294556f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_22 VNB N_A_266_94#_c_239_n 0.010932f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.275
cc_23 VNB N_A_266_94#_c_240_n 0.00257034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_266_94#_c_241_n 0.0351178f $X=-0.19 $Y=-0.245 $X2=0.347 $Y2=1.665
cc_25 VNB N_A_266_94#_c_242_n 8.27411e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_266_94#_c_243_n 0.0341041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_331_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_X_c_377_n 0.0267746f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.54
cc_29 VNB N_X_c_378_n 0.0144258f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.78
cc_30 VNB N_X_c_379_n 0.0248166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_402_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.03
cc_32 VNB N_VGND_c_403_n 0.0342445f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.54
cc_33 VNB N_VGND_c_404_n 0.0134281f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.78
cc_34 VNB N_VGND_c_405_n 0.0644827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_406_n 0.0191572f $X=-0.19 $Y=-0.245 $X2=0.347 $Y2=1.295
cc_36 VNB N_VGND_c_407_n 0.267554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_408_n 0.0113485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_A_N_c_75_n 0.0350681f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.03
cc_39 VPB N_A_N_c_72_n 0.0154589f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.78
cc_40 VPB N_A_N_c_77_n 0.0135533f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.94
cc_41 VPB N_A_N_c_74_n 0.00817485f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.275
cc_42 VPB N_A_114_74#_M1009_g 0.0271295f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.78
cc_43 VPB N_A_114_74#_c_111_n 0.0248397f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A_114_74#_c_108_n 0.0122024f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A_114_74#_c_113_n 0.00902376f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_114_74#_c_109_n 0.00814936f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_B_M1000_g 0.0223623f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.03
cc_48 VPB N_B_c_168_n 0.0056223f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_49 VPB N_B_c_171_n 0.00219656f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.78
cc_50 VPB N_C_M1008_g 0.0221631f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.03
cc_51 VPB N_C_c_204_n 0.0055832f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_52 VPB N_C_c_205_n 0.00512011f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.78
cc_53 VPB N_A_266_94#_M1001_g 0.0303296f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_54 VPB N_A_266_94#_c_240_n 0.00419179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_266_94#_c_246_n 0.0140282f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_266_94#_c_247_n 0.00361747f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_332_n 0.0120013f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.275
cc_58 VPB N_VPWR_c_333_n 0.0459907f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.615
cc_59 VPB N_VPWR_c_334_n 0.033688f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_60 VPB N_VPWR_c_335_n 0.0202647f $X=-0.19 $Y=1.66 $X2=0.405 $Y2=1.275
cc_61 VPB N_VPWR_c_336_n 0.0391783f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_337_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.347 $Y2=1.295
cc_63 VPB N_VPWR_c_338_n 0.0208961f $X=-0.19 $Y=1.66 $X2=0.347 $Y2=1.665
cc_64 VPB N_VPWR_c_339_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_340_n 0.0201177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_331_n 0.0857233f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB X 0.0433299f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_X_c_381_n 0.0158501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_X_c_379_n 0.00779946f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 N_A_N_M1006_g N_A_114_74#_c_105_n 0.00829387f $X=0.495 $Y=0.645 $X2=0
+ $Y2=0
cc_71 N_A_N_c_75_n N_A_114_74#_c_111_n 0.00430801f $X=0.51 $Y=2.03 $X2=0 $Y2=0
cc_72 N_A_N_M1006_g N_A_114_74#_c_106_n 0.00867488f $X=0.495 $Y=0.645 $X2=0
+ $Y2=0
cc_73 N_A_N_c_74_n N_A_114_74#_c_106_n 0.00725794f $X=0.405 $Y=1.275 $X2=0 $Y2=0
cc_74 N_A_N_c_73_n N_A_114_74#_c_107_n 0.00332712f $X=0.405 $Y=1.275 $X2=0 $Y2=0
cc_75 N_A_N_c_74_n N_A_114_74#_c_107_n 0.0397534f $X=0.405 $Y=1.275 $X2=0 $Y2=0
cc_76 N_A_N_M1006_g N_A_114_74#_c_108_n 0.0176124f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_77 N_A_N_c_71_n N_A_114_74#_c_108_n 0.0176124f $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_78 N_A_N_c_74_n N_A_114_74#_c_108_n 7.04297e-19 $X=0.405 $Y=1.275 $X2=0 $Y2=0
cc_79 N_A_N_c_75_n N_A_114_74#_c_113_n 0.00552779f $X=0.51 $Y=2.03 $X2=0 $Y2=0
cc_80 N_A_N_c_72_n N_A_114_74#_c_113_n 0.00332712f $X=0.405 $Y=1.78 $X2=0 $Y2=0
cc_81 N_A_N_c_71_n N_A_114_74#_c_109_n 0.00332712f $X=0.405 $Y=1.615 $X2=0 $Y2=0
cc_82 N_A_N_c_75_n N_VPWR_c_333_n 0.0219555f $X=0.51 $Y=2.03 $X2=0 $Y2=0
cc_83 N_A_N_c_72_n N_VPWR_c_333_n 0.00130639f $X=0.405 $Y=1.78 $X2=0 $Y2=0
cc_84 N_A_N_c_74_n N_VPWR_c_333_n 0.0180519f $X=0.405 $Y=1.275 $X2=0 $Y2=0
cc_85 N_A_N_c_75_n N_VPWR_c_336_n 0.00475445f $X=0.51 $Y=2.03 $X2=0 $Y2=0
cc_86 N_A_N_c_75_n N_VPWR_c_331_n 0.00943794f $X=0.51 $Y=2.03 $X2=0 $Y2=0
cc_87 N_A_N_M1006_g N_VGND_c_403_n 0.0180652f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_88 N_A_N_c_73_n N_VGND_c_403_n 0.0014092f $X=0.405 $Y=1.275 $X2=0 $Y2=0
cc_89 N_A_N_c_74_n N_VGND_c_403_n 0.0287296f $X=0.405 $Y=1.275 $X2=0 $Y2=0
cc_90 N_A_N_M1006_g N_VGND_c_405_n 0.00383152f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_91 N_A_N_M1006_g N_VGND_c_407_n 0.00762539f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_92 N_A_114_74#_c_103_n N_B_M1005_g 0.0548083f $X=1.69 $Y=1.185 $X2=0 $Y2=0
cc_93 N_A_114_74#_c_104_n N_B_M1005_g 0.0101789f $X=1.61 $Y=1.185 $X2=0 $Y2=0
cc_94 N_A_114_74#_M1009_g N_B_M1000_g 0.0225583f $X=1.7 $Y=2.26 $X2=0 $Y2=0
cc_95 N_A_114_74#_M1009_g N_B_c_168_n 0.0101789f $X=1.7 $Y=2.26 $X2=0 $Y2=0
cc_96 N_A_114_74#_M1009_g N_B_c_171_n 8.68275e-19 $X=1.7 $Y=2.26 $X2=0 $Y2=0
cc_97 N_A_114_74#_c_104_n N_B_c_171_n 0.00102127f $X=1.61 $Y=1.185 $X2=0 $Y2=0
cc_98 N_A_114_74#_c_103_n N_A_266_94#_c_239_n 0.0112826f $X=1.69 $Y=1.185 $X2=0
+ $Y2=0
cc_99 N_A_114_74#_c_105_n N_A_266_94#_c_239_n 0.0159343f $X=0.78 $Y=0.645 $X2=0
+ $Y2=0
cc_100 N_A_114_74#_c_106_n N_A_266_94#_c_239_n 0.013901f $X=0.957 $Y=1.212 $X2=0
+ $Y2=0
cc_101 N_A_114_74#_c_101_n N_A_266_94#_c_240_n 0.00983996f $X=1.61 $Y=1.26 $X2=0
+ $Y2=0
cc_102 N_A_114_74#_M1009_g N_A_266_94#_c_240_n 0.0156157f $X=1.7 $Y=2.26 $X2=0
+ $Y2=0
cc_103 N_A_114_74#_c_104_n N_A_266_94#_c_240_n 0.00489741f $X=1.61 $Y=1.185
+ $X2=0 $Y2=0
cc_104 N_A_114_74#_c_107_n N_A_266_94#_c_240_n 0.0376823f $X=0.957 $Y=1.518
+ $X2=0 $Y2=0
cc_105 N_A_114_74#_c_108_n N_A_266_94#_c_240_n 0.00320796f $X=0.975 $Y=1.195
+ $X2=0 $Y2=0
cc_106 N_A_114_74#_c_113_n N_A_266_94#_c_240_n 0.0116419f $X=0.78 $Y=2.1 $X2=0
+ $Y2=0
cc_107 N_A_114_74#_c_103_n N_A_266_94#_c_241_n 0.00839128f $X=1.69 $Y=1.185
+ $X2=0 $Y2=0
cc_108 N_A_114_74#_c_104_n N_A_266_94#_c_241_n 0.00733763f $X=1.61 $Y=1.185
+ $X2=0 $Y2=0
cc_109 N_A_114_74#_M1009_g N_A_266_94#_c_259_n 0.0179146f $X=1.7 $Y=2.26 $X2=0
+ $Y2=0
cc_110 N_A_114_74#_c_101_n N_A_266_94#_c_242_n 0.00878777f $X=1.61 $Y=1.26 $X2=0
+ $Y2=0
cc_111 N_A_114_74#_c_103_n N_A_266_94#_c_242_n 0.00134888f $X=1.69 $Y=1.185
+ $X2=0 $Y2=0
cc_112 N_A_114_74#_c_104_n N_A_266_94#_c_242_n 2.24561e-19 $X=1.61 $Y=1.185
+ $X2=0 $Y2=0
cc_113 N_A_114_74#_c_106_n N_A_266_94#_c_242_n 0.013702f $X=0.957 $Y=1.212 $X2=0
+ $Y2=0
cc_114 N_A_114_74#_c_107_n N_A_266_94#_c_242_n 6.05e-19 $X=0.957 $Y=1.518 $X2=0
+ $Y2=0
cc_115 N_A_114_74#_c_108_n N_A_266_94#_c_242_n 6.14826e-19 $X=0.975 $Y=1.195
+ $X2=0 $Y2=0
cc_116 N_A_114_74#_M1009_g N_A_266_94#_c_246_n 0.0127862f $X=1.7 $Y=2.26 $X2=0
+ $Y2=0
cc_117 N_A_114_74#_c_111_n N_A_266_94#_c_246_n 0.0284313f $X=0.78 $Y=2.265 $X2=0
+ $Y2=0
cc_118 N_A_114_74#_c_113_n N_A_266_94#_c_246_n 0.00847258f $X=0.78 $Y=2.1 $X2=0
+ $Y2=0
cc_119 N_A_114_74#_M1009_g N_A_266_94#_c_247_n 5.36924e-19 $X=1.7 $Y=2.26 $X2=0
+ $Y2=0
cc_120 N_A_114_74#_c_111_n N_VPWR_c_333_n 0.0346006f $X=0.78 $Y=2.265 $X2=0
+ $Y2=0
cc_121 N_A_114_74#_M1009_g N_VPWR_c_334_n 0.00363277f $X=1.7 $Y=2.26 $X2=0 $Y2=0
cc_122 N_A_114_74#_M1009_g N_VPWR_c_336_n 0.00465228f $X=1.7 $Y=2.26 $X2=0 $Y2=0
cc_123 N_A_114_74#_c_111_n N_VPWR_c_336_n 0.0146357f $X=0.78 $Y=2.265 $X2=0
+ $Y2=0
cc_124 N_A_114_74#_M1009_g N_VPWR_c_331_n 0.00555093f $X=1.7 $Y=2.26 $X2=0 $Y2=0
cc_125 N_A_114_74#_c_111_n N_VPWR_c_331_n 0.0121141f $X=0.78 $Y=2.265 $X2=0
+ $Y2=0
cc_126 N_A_114_74#_c_105_n N_VGND_c_403_n 0.0167375f $X=0.78 $Y=0.645 $X2=0
+ $Y2=0
cc_127 N_A_114_74#_c_106_n N_VGND_c_403_n 0.00701512f $X=0.957 $Y=1.212 $X2=0
+ $Y2=0
cc_128 N_A_114_74#_c_103_n N_VGND_c_405_n 0.00485498f $X=1.69 $Y=1.185 $X2=0
+ $Y2=0
cc_129 N_A_114_74#_c_105_n N_VGND_c_405_n 0.0145628f $X=0.78 $Y=0.645 $X2=0
+ $Y2=0
cc_130 N_A_114_74#_c_103_n N_VGND_c_407_n 0.00514438f $X=1.69 $Y=1.185 $X2=0
+ $Y2=0
cc_131 N_A_114_74#_c_105_n N_VGND_c_407_n 0.012086f $X=0.78 $Y=0.645 $X2=0 $Y2=0
cc_132 N_B_M1005_g N_C_M1007_g 0.0335091f $X=2.08 $Y=0.79 $X2=0 $Y2=0
cc_133 N_B_M1000_g N_C_M1008_g 0.0187829f $X=2.245 $Y=2.26 $X2=0 $Y2=0
cc_134 N_B_c_168_n N_C_c_204_n 0.0211575f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_135 N_B_c_171_n N_C_c_204_n 3.50941e-19 $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_136 N_B_c_168_n N_C_c_205_n 0.00226045f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_137 N_B_c_171_n N_C_c_205_n 0.0284944f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_138 N_B_M1005_g N_A_266_94#_c_239_n 0.00297121f $X=2.08 $Y=0.79 $X2=0 $Y2=0
cc_139 N_B_M1005_g N_A_266_94#_c_240_n 0.00165598f $X=2.08 $Y=0.79 $X2=0 $Y2=0
cc_140 N_B_M1000_g N_A_266_94#_c_240_n 8.6467e-19 $X=2.245 $Y=2.26 $X2=0 $Y2=0
cc_141 N_B_c_171_n N_A_266_94#_c_240_n 0.0162405f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_142 N_B_M1005_g N_A_266_94#_c_241_n 0.0152776f $X=2.08 $Y=0.79 $X2=0 $Y2=0
cc_143 N_B_c_168_n N_A_266_94#_c_241_n 0.00498422f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_144 N_B_c_171_n N_A_266_94#_c_241_n 0.0245335f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_145 N_B_M1000_g N_A_266_94#_c_259_n 0.013768f $X=2.245 $Y=2.26 $X2=0 $Y2=0
cc_146 N_B_c_168_n N_A_266_94#_c_259_n 6.98124e-19 $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_147 N_B_c_171_n N_A_266_94#_c_259_n 0.0209931f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_148 N_B_M1000_g N_A_266_94#_c_246_n 5.42137e-19 $X=2.245 $Y=2.26 $X2=0 $Y2=0
cc_149 N_B_M1000_g N_A_266_94#_c_247_n 0.00970529f $X=2.245 $Y=2.26 $X2=0 $Y2=0
cc_150 N_B_c_171_n N_A_266_94#_c_247_n 0.00194922f $X=2.17 $Y=1.515 $X2=0 $Y2=0
cc_151 N_B_M1000_g N_VPWR_c_334_n 0.0036579f $X=2.245 $Y=2.26 $X2=0 $Y2=0
cc_152 N_B_M1000_g N_VPWR_c_338_n 0.00468269f $X=2.245 $Y=2.26 $X2=0 $Y2=0
cc_153 N_B_M1000_g N_VPWR_c_331_n 0.00555093f $X=2.245 $Y=2.26 $X2=0 $Y2=0
cc_154 N_B_M1005_g N_VGND_c_404_n 0.00268474f $X=2.08 $Y=0.79 $X2=0 $Y2=0
cc_155 N_B_M1005_g N_VGND_c_405_n 0.00507111f $X=2.08 $Y=0.79 $X2=0 $Y2=0
cc_156 N_B_M1005_g N_VGND_c_407_n 0.00514438f $X=2.08 $Y=0.79 $X2=0 $Y2=0
cc_157 N_C_M1008_g N_A_266_94#_M1001_g 0.0176825f $X=2.7 $Y=2.26 $X2=0 $Y2=0
cc_158 N_C_c_204_n N_A_266_94#_M1001_g 0.00208102f $X=2.71 $Y=1.515 $X2=0 $Y2=0
cc_159 N_C_c_205_n N_A_266_94#_M1001_g 0.00241556f $X=2.71 $Y=1.515 $X2=0 $Y2=0
cc_160 N_C_M1007_g N_A_266_94#_M1003_g 0.00939291f $X=2.62 $Y=0.79 $X2=0 $Y2=0
cc_161 N_C_M1007_g N_A_266_94#_c_241_n 0.0170163f $X=2.62 $Y=0.79 $X2=0 $Y2=0
cc_162 N_C_c_204_n N_A_266_94#_c_241_n 0.00695803f $X=2.71 $Y=1.515 $X2=0 $Y2=0
cc_163 N_C_c_205_n N_A_266_94#_c_241_n 0.0454831f $X=2.71 $Y=1.515 $X2=0 $Y2=0
cc_164 N_C_M1008_g N_A_266_94#_c_247_n 0.0106357f $X=2.7 $Y=2.26 $X2=0 $Y2=0
cc_165 N_C_c_204_n N_A_266_94#_c_247_n 2.52994e-19 $X=2.71 $Y=1.515 $X2=0 $Y2=0
cc_166 N_C_c_205_n N_A_266_94#_c_247_n 0.0072311f $X=2.71 $Y=1.515 $X2=0 $Y2=0
cc_167 N_C_M1007_g N_A_266_94#_c_243_n 0.00132954f $X=2.62 $Y=0.79 $X2=0 $Y2=0
cc_168 N_C_c_204_n N_A_266_94#_c_243_n 0.0175012f $X=2.71 $Y=1.515 $X2=0 $Y2=0
cc_169 N_C_c_205_n N_A_266_94#_c_243_n 2.7599e-19 $X=2.71 $Y=1.515 $X2=0 $Y2=0
cc_170 N_C_M1008_g N_VPWR_c_335_n 0.00776968f $X=2.7 $Y=2.26 $X2=0 $Y2=0
cc_171 N_C_c_205_n N_VPWR_c_335_n 0.00242374f $X=2.71 $Y=1.515 $X2=0 $Y2=0
cc_172 N_C_M1008_g N_VPWR_c_338_n 0.00465228f $X=2.7 $Y=2.26 $X2=0 $Y2=0
cc_173 N_C_M1008_g N_VPWR_c_331_n 0.00555093f $X=2.7 $Y=2.26 $X2=0 $Y2=0
cc_174 N_C_M1007_g N_X_c_377_n 6.21799e-19 $X=2.62 $Y=0.79 $X2=0 $Y2=0
cc_175 N_C_M1008_g N_X_c_381_n 7.50962e-19 $X=2.7 $Y=2.26 $X2=0 $Y2=0
cc_176 N_C_M1007_g N_VGND_c_404_n 0.0203753f $X=2.62 $Y=0.79 $X2=0 $Y2=0
cc_177 N_C_M1007_g N_VGND_c_405_n 0.00269285f $X=2.62 $Y=0.79 $X2=0 $Y2=0
cc_178 N_C_M1007_g N_VGND_c_407_n 0.00277796f $X=2.62 $Y=0.79 $X2=0 $Y2=0
cc_179 N_A_266_94#_c_259_n N_VPWR_M1009_d 0.00957916f $X=2.31 $Y=2.035 $X2=0
+ $Y2=0
cc_180 N_A_266_94#_c_259_n N_VPWR_c_334_n 0.020421f $X=2.31 $Y=2.035 $X2=0 $Y2=0
cc_181 N_A_266_94#_c_246_n N_VPWR_c_334_n 0.0161747f $X=1.475 $Y=1.985 $X2=0
+ $Y2=0
cc_182 N_A_266_94#_c_247_n N_VPWR_c_334_n 0.0161746f $X=2.475 $Y=2.115 $X2=0
+ $Y2=0
cc_183 N_A_266_94#_M1001_g N_VPWR_c_335_n 0.00917005f $X=3.285 $Y=2.4 $X2=0
+ $Y2=0
cc_184 N_A_266_94#_c_241_n N_VPWR_c_335_n 0.00600469f $X=3.045 $Y=1.135 $X2=0
+ $Y2=0
cc_185 N_A_266_94#_c_247_n N_VPWR_c_335_n 0.019396f $X=2.475 $Y=2.115 $X2=0
+ $Y2=0
cc_186 N_A_266_94#_c_243_n N_VPWR_c_335_n 5.04644e-19 $X=3.25 $Y=1.465 $X2=0
+ $Y2=0
cc_187 N_A_266_94#_c_246_n N_VPWR_c_336_n 0.0066444f $X=1.475 $Y=1.985 $X2=0
+ $Y2=0
cc_188 N_A_266_94#_c_247_n N_VPWR_c_338_n 0.00658022f $X=2.475 $Y=2.115 $X2=0
+ $Y2=0
cc_189 N_A_266_94#_M1001_g N_VPWR_c_340_n 0.005209f $X=3.285 $Y=2.4 $X2=0 $Y2=0
cc_190 N_A_266_94#_M1001_g N_VPWR_c_331_n 0.0099063f $X=3.285 $Y=2.4 $X2=0 $Y2=0
cc_191 N_A_266_94#_c_246_n N_VPWR_c_331_n 0.00995531f $X=1.475 $Y=1.985 $X2=0
+ $Y2=0
cc_192 N_A_266_94#_c_247_n N_VPWR_c_331_n 0.00992017f $X=2.475 $Y=2.115 $X2=0
+ $Y2=0
cc_193 N_A_266_94#_M1003_g N_X_c_377_n 0.00888737f $X=3.335 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A_266_94#_M1003_g N_X_c_378_n 0.00396511f $X=3.335 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A_266_94#_c_241_n N_X_c_378_n 0.00630461f $X=3.045 $Y=1.135 $X2=0 $Y2=0
cc_196 N_A_266_94#_M1001_g X 0.0126855f $X=3.285 $Y=2.4 $X2=0 $Y2=0
cc_197 N_A_266_94#_M1001_g N_X_c_381_n 0.0045115f $X=3.285 $Y=2.4 $X2=0 $Y2=0
cc_198 N_A_266_94#_c_241_n N_X_c_381_n 0.00524276f $X=3.045 $Y=1.135 $X2=0 $Y2=0
cc_199 N_A_266_94#_c_243_n N_X_c_381_n 3.09009e-19 $X=3.25 $Y=1.465 $X2=0 $Y2=0
cc_200 N_A_266_94#_M1001_g N_X_c_379_n 0.00467041f $X=3.285 $Y=2.4 $X2=0 $Y2=0
cc_201 N_A_266_94#_M1003_g N_X_c_379_n 0.00252147f $X=3.335 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A_266_94#_c_241_n N_X_c_379_n 0.0306189f $X=3.045 $Y=1.135 $X2=0 $Y2=0
cc_203 N_A_266_94#_c_243_n N_X_c_379_n 0.00232633f $X=3.25 $Y=1.465 $X2=0 $Y2=0
cc_204 N_A_266_94#_c_241_n N_VGND_M1007_d 0.00592064f $X=3.045 $Y=1.135 $X2=0
+ $Y2=0
cc_205 N_A_266_94#_M1003_g N_VGND_c_404_n 0.00656426f $X=3.335 $Y=0.74 $X2=0
+ $Y2=0
cc_206 N_A_266_94#_c_241_n N_VGND_c_404_n 0.043095f $X=3.045 $Y=1.135 $X2=0
+ $Y2=0
cc_207 N_A_266_94#_c_243_n N_VGND_c_404_n 5.6341e-19 $X=3.25 $Y=1.465 $X2=0
+ $Y2=0
cc_208 N_A_266_94#_c_239_n N_VGND_c_405_n 0.0103491f $X=1.475 $Y=0.615 $X2=0
+ $Y2=0
cc_209 N_A_266_94#_M1003_g N_VGND_c_406_n 0.00434272f $X=3.335 $Y=0.74 $X2=0
+ $Y2=0
cc_210 N_A_266_94#_M1003_g N_VGND_c_407_n 0.00828751f $X=3.335 $Y=0.74 $X2=0
+ $Y2=0
cc_211 N_A_266_94#_c_239_n N_VGND_c_407_n 0.0113354f $X=1.475 $Y=0.615 $X2=0
+ $Y2=0
cc_212 N_A_266_94#_c_241_n A_353_94# 0.0048076f $X=3.045 $Y=1.135 $X2=-0.19
+ $Y2=-0.245
cc_213 N_A_266_94#_c_241_n A_431_94# 0.0106289f $X=3.045 $Y=1.135 $X2=-0.19
+ $Y2=-0.245
cc_214 N_VPWR_c_340_n X 0.0181186f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_215 N_VPWR_c_331_n X 0.0149289f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_216 N_VPWR_c_335_n N_X_c_381_n 0.0407049f $X=3.01 $Y=2.115 $X2=0 $Y2=0
cc_217 N_X_c_377_n N_VGND_c_404_n 0.0211012f $X=3.55 $Y=0.515 $X2=0 $Y2=0
cc_218 N_X_c_377_n N_VGND_c_406_n 0.0163488f $X=3.55 $Y=0.515 $X2=0 $Y2=0
cc_219 N_X_c_377_n N_VGND_c_407_n 0.0134757f $X=3.55 $Y=0.515 $X2=0 $Y2=0

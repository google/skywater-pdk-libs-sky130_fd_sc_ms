* File: sky130_fd_sc_ms__or4_4.pxi.spice
* Created: Fri Aug 28 18:09:05 2020
* 
x_PM_SKY130_FD_SC_MS__OR4_4%A_83_264# N_A_83_264#_M1004_d N_A_83_264#_M1015_d
+ N_A_83_264#_M1000_d N_A_83_264#_M1005_g N_A_83_264#_M1001_g
+ N_A_83_264#_M1006_g N_A_83_264#_M1007_g N_A_83_264#_M1008_g
+ N_A_83_264#_M1010_g N_A_83_264#_M1011_g N_A_83_264#_M1012_g
+ N_A_83_264#_c_117_n N_A_83_264#_c_118_n N_A_83_264#_c_134_p
+ N_A_83_264#_c_262_p N_A_83_264#_c_119_n N_A_83_264#_c_141_p
+ N_A_83_264#_c_120_n N_A_83_264#_c_121_n N_A_83_264#_c_129_n
+ N_A_83_264#_c_122_n N_A_83_264#_c_123_n N_A_83_264#_c_140_p
+ N_A_83_264#_c_124_n N_A_83_264#_c_131_n PM_SKY130_FD_SC_MS__OR4_4%A_83_264#
x_PM_SKY130_FD_SC_MS__OR4_4%B N_B_c_273_n N_B_M1014_g N_B_c_275_n N_B_M1004_g
+ N_B_M1018_g N_B_c_277_n N_B_c_278_n N_B_c_279_n N_B_c_280_n B B
+ PM_SKY130_FD_SC_MS__OR4_4%B
x_PM_SKY130_FD_SC_MS__OR4_4%A N_A_M1013_g N_A_M1016_g N_A_M1017_g A N_A_c_358_n
+ PM_SKY130_FD_SC_MS__OR4_4%A
x_PM_SKY130_FD_SC_MS__OR4_4%C N_C_M1015_g N_C_M1003_g N_C_M1019_g C C C
+ N_C_c_404_n N_C_c_405_n N_C_c_406_n N_C_c_407_n PM_SKY130_FD_SC_MS__OR4_4%C
x_PM_SKY130_FD_SC_MS__OR4_4%D N_D_c_470_n N_D_M1009_g N_D_M1000_g N_D_M1002_g
+ N_D_c_473_n N_D_c_474_n N_D_c_475_n N_D_c_476_n D N_D_c_477_n N_D_c_478_n
+ PM_SKY130_FD_SC_MS__OR4_4%D
x_PM_SKY130_FD_SC_MS__OR4_4%VPWR N_VPWR_M1005_s N_VPWR_M1006_s N_VPWR_M1011_s
+ N_VPWR_M1016_d N_VPWR_c_527_n N_VPWR_c_528_n N_VPWR_c_529_n N_VPWR_c_530_n
+ N_VPWR_c_531_n VPWR N_VPWR_c_532_n N_VPWR_c_533_n N_VPWR_c_534_n
+ N_VPWR_c_535_n N_VPWR_c_526_n N_VPWR_c_537_n N_VPWR_c_538_n N_VPWR_c_539_n
+ PM_SKY130_FD_SC_MS__OR4_4%VPWR
x_PM_SKY130_FD_SC_MS__OR4_4%X N_X_M1001_s N_X_M1010_s N_X_M1005_d N_X_M1008_d
+ N_X_c_612_n N_X_c_613_n N_X_c_617_n N_X_c_614_n N_X_c_618_n N_X_c_615_n X X X
+ X N_X_c_621_n PM_SKY130_FD_SC_MS__OR4_4%X
x_PM_SKY130_FD_SC_MS__OR4_4%A_499_392# N_A_499_392#_M1014_s N_A_499_392#_M1018_s
+ N_A_499_392#_M1019_d N_A_499_392#_c_681_n N_A_499_392#_c_682_n
+ N_A_499_392#_c_699_n N_A_499_392#_c_683_n N_A_499_392#_c_690_n
+ N_A_499_392#_c_684_n N_A_499_392#_c_691_n N_A_499_392#_c_722_n
+ N_A_499_392#_c_685_n PM_SKY130_FD_SC_MS__OR4_4%A_499_392#
x_PM_SKY130_FD_SC_MS__OR4_4%A_591_392# N_A_591_392#_M1014_d N_A_591_392#_M1017_s
+ N_A_591_392#_c_753_n N_A_591_392#_c_751_n N_A_591_392#_c_757_n
+ N_A_591_392#_c_755_n N_A_591_392#_c_752_n PM_SKY130_FD_SC_MS__OR4_4%A_591_392#
x_PM_SKY130_FD_SC_MS__OR4_4%A_965_392# N_A_965_392#_M1003_s N_A_965_392#_M1002_s
+ N_A_965_392#_c_779_n PM_SKY130_FD_SC_MS__OR4_4%A_965_392#
x_PM_SKY130_FD_SC_MS__OR4_4%VGND N_VGND_M1001_d N_VGND_M1007_d N_VGND_M1012_d
+ N_VGND_M1013_d N_VGND_M1009_d N_VGND_c_792_n N_VGND_c_793_n N_VGND_c_794_n
+ N_VGND_c_795_n VGND N_VGND_c_796_n N_VGND_c_797_n N_VGND_c_798_n
+ N_VGND_c_799_n N_VGND_c_800_n N_VGND_c_801_n N_VGND_c_802_n N_VGND_c_803_n
+ N_VGND_c_804_n N_VGND_c_805_n PM_SKY130_FD_SC_MS__OR4_4%VGND
cc_1 VNB N_A_83_264#_M1005_g 0.00539279f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A_83_264#_M1001_g 0.0272031f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_3 VNB N_A_83_264#_M1006_g 0.00433407f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_4 VNB N_A_83_264#_M1007_g 0.0219865f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_5 VNB N_A_83_264#_M1008_g 4.7811e-19 $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_6 VNB N_A_83_264#_M1010_g 0.0256793f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=0.74
cc_7 VNB N_A_83_264#_M1011_g 7.57144e-19 $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_8 VNB N_A_83_264#_M1012_g 0.0265883f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=0.74
cc_9 VNB N_A_83_264#_c_117_n 6.71782e-19 $X=-0.19 $Y=-0.245 $X2=2.155 $Y2=1.485
cc_10 VNB N_A_83_264#_c_118_n 0.008967f $X=-0.19 $Y=-0.245 $X2=2.24 $Y2=1.32
cc_11 VNB N_A_83_264#_c_119_n 0.00239713f $X=-0.19 $Y=-0.245 $X2=3.085 $Y2=0.515
cc_12 VNB N_A_83_264#_c_120_n 0.00280366f $X=-0.19 $Y=-0.245 $X2=4.935 $Y2=0.515
cc_13 VNB N_A_83_264#_c_121_n 0.0283703f $X=-0.19 $Y=-0.245 $X2=6.465 $Y2=1.11
cc_14 VNB N_A_83_264#_c_122_n 0.0231448f $X=-0.19 $Y=-0.245 $X2=6.55 $Y2=1.95
cc_15 VNB N_A_83_264#_c_123_n 0.113549f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.485
cc_16 VNB N_A_83_264#_c_124_n 0.00258271f $X=-0.19 $Y=-0.245 $X2=4.935 $Y2=0.875
cc_17 VNB N_B_c_273_n 0.0361513f $X=-0.19 $Y=-0.245 $X2=2.945 $Y2=0.37
cc_18 VNB N_B_M1014_g 0.00142475f $X=-0.19 $Y=-0.245 $X2=5.325 $Y2=1.96
cc_19 VNB N_B_c_275_n 0.0182315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B_M1018_g 0.00629716f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.57
cc_21 VNB N_B_c_277_n 0.0154954f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_22 VNB N_B_c_278_n 0.0151427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B_c_279_n 0.0060756f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.32
cc_24 VNB N_B_c_280_n 0.0397096f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.57
cc_25 VNB N_A_M1013_g 0.0336515f $X=-0.19 $Y=-0.245 $X2=5.325 $Y2=1.96
cc_26 VNB A 0.00304223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_c_358_n 0.032858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_C_M1015_g 0.0306063f $X=-0.19 $Y=-0.245 $X2=5.325 $Y2=1.96
cc_29 VNB N_C_c_404_n 0.0176735f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_30 VNB N_C_c_405_n 0.0286189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_C_c_406_n 0.00148209f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.65
cc_32 VNB N_C_c_407_n 0.00637831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_D_c_470_n 0.0169511f $X=-0.19 $Y=-0.245 $X2=2.945 $Y2=0.37
cc_34 VNB N_D_M1000_g 0.00733563f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_D_M1002_g 0.00733563f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.57
cc_36 VNB N_D_c_473_n 0.0176918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_D_c_474_n 0.054246f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.32
cc_38 VNB N_D_c_475_n 0.00909013f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_39 VNB N_D_c_476_n 0.0403232f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_40 VNB N_D_c_477_n 0.0691165f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.65
cc_41 VNB N_D_c_478_n 0.00238263f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_42 VNB N_VPWR_c_526_n 0.283096f $X=-0.19 $Y=-0.245 $X2=3.085 $Y2=0.515
cc_43 VNB N_X_c_612_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_44 VNB N_X_c_613_n 0.0209897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_X_c_614_n 0.00674496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_X_c_615_n 0.0033365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_792_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_48 VNB N_VGND_c_793_n 0.0449905f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.57
cc_49 VNB N_VGND_c_794_n 0.00571618f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.32
cc_50 VNB N_VGND_c_795_n 0.00950637f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.65
cc_51 VNB N_VGND_c_796_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=1.32
cc_52 VNB N_VGND_c_797_n 0.0269696f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_53 VNB N_VGND_c_798_n 0.018096f $X=-0.19 $Y=-0.245 $X2=3.085 $Y2=0.515
cc_54 VNB N_VGND_c_799_n 0.362172f $X=-0.19 $Y=-0.245 $X2=3.085 $Y2=0.515
cc_55 VNB N_VGND_c_800_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=4.935 $Y2=0.515
cc_56 VNB N_VGND_c_801_n 0.00689995f $X=-0.19 $Y=-0.245 $X2=5.1 $Y2=1.11
cc_57 VNB N_VGND_c_802_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=6.55 $Y2=1.95
cc_58 VNB N_VGND_c_803_n 0.0378507f $X=-0.19 $Y=-0.245 $X2=5.46 $Y2=2.105
cc_59 VNB N_VGND_c_804_n 0.0176133f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.485
cc_60 VNB N_VGND_c_805_n 0.0344666f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=1.485
cc_61 VPB N_A_83_264#_M1005_g 0.0251338f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_62 VPB N_A_83_264#_M1006_g 0.0209526f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_63 VPB N_A_83_264#_M1008_g 0.0216178f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_64 VPB N_A_83_264#_M1011_g 0.0289227f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_65 VPB N_A_83_264#_c_129_n 0.0181071f $X=-0.19 $Y=1.66 $X2=6.465 $Y2=2.035
cc_66 VPB N_A_83_264#_c_122_n 0.0141543f $X=-0.19 $Y=1.66 $X2=6.55 $Y2=1.95
cc_67 VPB N_A_83_264#_c_131_n 0.00230067f $X=-0.19 $Y=1.66 $X2=5.625 $Y2=2.07
cc_68 VPB N_B_M1014_g 0.0376488f $X=-0.19 $Y=1.66 $X2=5.325 $Y2=1.96
cc_69 VPB N_B_M1018_g 0.0312878f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.57
cc_70 VPB N_A_M1016_g 0.0212401f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_M1017_g 0.0214621f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_72 VPB A 8.34758e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_c_358_n 0.0175259f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_C_M1003_g 0.0251301f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_C_M1019_g 0.027499f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_76 VPB N_C_c_404_n 0.0107264f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_77 VPB N_C_c_405_n 0.0119929f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_C_c_406_n 0.0043287f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.65
cc_79 VPB N_C_c_407_n 0.0070921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_D_M1000_g 0.0285359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_D_M1002_g 0.0277964f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.57
cc_82 VPB N_VPWR_c_527_n 0.0119967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_528_n 0.0340261f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_84 VPB N_VPWR_c_529_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_85 VPB N_VPWR_c_530_n 0.0120686f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_86 VPB N_VPWR_c_531_n 0.00396467f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_87 VPB N_VPWR_c_532_n 0.0159778f $X=-0.19 $Y=1.66 $X2=1.495 $Y2=0.74
cc_88 VPB N_VPWR_c_533_n 0.0159778f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_89 VPB N_VPWR_c_534_n 0.0313938f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_535_n 0.0810424f $X=-0.19 $Y=1.66 $X2=3.085 $Y2=0.79
cc_91 VPB N_VPWR_c_526_n 0.0829084f $X=-0.19 $Y=1.66 $X2=3.085 $Y2=0.515
cc_92 VPB N_VPWR_c_537_n 0.00601644f $X=-0.19 $Y=1.66 $X2=4.935 $Y2=0.515
cc_93 VPB N_VPWR_c_538_n 0.0061274f $X=-0.19 $Y=1.66 $X2=6.465 $Y2=1.11
cc_94 VPB N_VPWR_c_539_n 0.00601668f $X=-0.19 $Y=1.66 $X2=5.625 $Y2=2.035
cc_95 VPB N_X_c_613_n 0.0208972f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_X_c_617_n 0.00233077f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_97 VPB N_X_c_618_n 0.00233077f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB X 0.00186725f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.65
cc_99 VPB X 0.00755712f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_100 VPB N_X_c_621_n 0.00375655f $X=-0.19 $Y=1.66 $X2=2.155 $Y2=1.485
cc_101 VPB N_A_499_392#_c_681_n 0.00738124f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.57
cc_102 VPB N_A_499_392#_c_682_n 0.0103883f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_103 VPB N_A_499_392#_c_683_n 0.00948185f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_104 VPB N_A_499_392#_c_684_n 0.00275675f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_105 VPB N_A_499_392#_c_685_n 0.0300793f $X=-0.19 $Y=1.66 $X2=1.495 $Y2=0.74
cc_106 VPB N_A_591_392#_c_751_n 0.00228692f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_591_392#_c_752_n 0.00230033f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_108 VPB N_A_965_392#_c_779_n 0.00728342f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_109 N_A_83_264#_M1012_g N_B_c_273_n 0.0139171f $X=2.25 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_110 N_A_83_264#_c_118_n N_B_c_273_n 9.47471e-19 $X=2.24 $Y=1.32 $X2=-0.19
+ $Y2=-0.245
cc_111 N_A_83_264#_c_134_p N_B_c_273_n 8.96913e-19 $X=2.92 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_112 N_A_83_264#_c_123_n N_B_c_273_n 0.00225496f $X=2.16 $Y=1.485 $X2=-0.19
+ $Y2=-0.245
cc_113 N_A_83_264#_M1012_g N_B_c_275_n 0.0204288f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_114 N_A_83_264#_c_118_n N_B_c_275_n 0.00101364f $X=2.24 $Y=1.32 $X2=0 $Y2=0
cc_115 N_A_83_264#_c_134_p N_B_c_275_n 0.0092233f $X=2.92 $Y=0.875 $X2=0 $Y2=0
cc_116 N_A_83_264#_c_119_n N_B_c_275_n 0.00689388f $X=3.085 $Y=0.515 $X2=0 $Y2=0
cc_117 N_A_83_264#_c_140_p N_B_c_275_n 7.15033e-19 $X=3.085 $Y=0.875 $X2=0 $Y2=0
cc_118 N_A_83_264#_c_141_p N_B_c_277_n 0.0574059f $X=4.77 $Y=0.875 $X2=0 $Y2=0
cc_119 N_A_83_264#_c_140_p N_B_c_277_n 0.00109891f $X=3.085 $Y=0.875 $X2=0 $Y2=0
cc_120 N_A_83_264#_M1012_g N_B_c_278_n 0.00140149f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_121 N_A_83_264#_c_118_n N_B_c_278_n 0.0283182f $X=2.24 $Y=1.32 $X2=0 $Y2=0
cc_122 N_A_83_264#_c_134_p N_B_c_278_n 0.02837f $X=2.92 $Y=0.875 $X2=0 $Y2=0
cc_123 N_A_83_264#_c_123_n N_B_c_278_n 5.52866e-19 $X=2.16 $Y=1.485 $X2=0 $Y2=0
cc_124 N_A_83_264#_c_140_p N_B_c_278_n 0.0223159f $X=3.085 $Y=0.875 $X2=0 $Y2=0
cc_125 N_A_83_264#_c_141_p N_B_c_279_n 0.0261968f $X=4.77 $Y=0.875 $X2=0 $Y2=0
cc_126 N_A_83_264#_c_124_n N_B_c_279_n 0.00285444f $X=4.935 $Y=0.875 $X2=0 $Y2=0
cc_127 N_A_83_264#_c_141_p N_B_c_280_n 0.00181415f $X=4.77 $Y=0.875 $X2=0 $Y2=0
cc_128 N_A_83_264#_c_119_n N_A_M1013_g 0.010756f $X=3.085 $Y=0.515 $X2=0 $Y2=0
cc_129 N_A_83_264#_c_141_p N_A_M1013_g 0.0104279f $X=4.77 $Y=0.875 $X2=0 $Y2=0
cc_130 N_A_83_264#_c_140_p N_A_M1013_g 7.15645e-19 $X=3.085 $Y=0.875 $X2=0 $Y2=0
cc_131 N_A_83_264#_c_141_p N_C_M1015_g 0.0120241f $X=4.77 $Y=0.875 $X2=0 $Y2=0
cc_132 N_A_83_264#_c_120_n N_C_M1015_g 0.0114883f $X=4.935 $Y=0.515 $X2=0 $Y2=0
cc_133 N_A_83_264#_c_124_n N_C_M1015_g 0.0106918f $X=4.935 $Y=0.875 $X2=0 $Y2=0
cc_134 N_A_83_264#_c_131_n N_C_M1003_g 7.19448e-19 $X=5.625 $Y=2.07 $X2=0 $Y2=0
cc_135 N_A_83_264#_c_129_n N_C_M1019_g 0.013807f $X=6.465 $Y=2.035 $X2=0 $Y2=0
cc_136 N_A_83_264#_c_122_n N_C_M1019_g 0.00547941f $X=6.55 $Y=1.95 $X2=0 $Y2=0
cc_137 N_A_83_264#_c_131_n N_C_M1019_g 3.29019e-19 $X=5.625 $Y=2.07 $X2=0 $Y2=0
cc_138 N_A_83_264#_c_124_n N_C_c_404_n 9.09904e-19 $X=4.935 $Y=0.875 $X2=0 $Y2=0
cc_139 N_A_83_264#_c_121_n N_C_c_405_n 0.00338597f $X=6.465 $Y=1.11 $X2=0 $Y2=0
cc_140 N_A_83_264#_c_129_n N_C_c_405_n 0.0039803f $X=6.465 $Y=2.035 $X2=0 $Y2=0
cc_141 N_A_83_264#_c_122_n N_C_c_405_n 0.00960216f $X=6.55 $Y=1.95 $X2=0 $Y2=0
cc_142 N_A_83_264#_c_121_n N_C_c_406_n 0.0715147f $X=6.465 $Y=1.11 $X2=0 $Y2=0
cc_143 N_A_83_264#_c_122_n N_C_c_406_n 0.0315994f $X=6.55 $Y=1.95 $X2=0 $Y2=0
cc_144 N_A_83_264#_c_131_n N_C_c_406_n 0.0734148f $X=5.625 $Y=2.07 $X2=0 $Y2=0
cc_145 N_A_83_264#_c_141_p N_C_c_407_n 0.00546445f $X=4.77 $Y=0.875 $X2=0 $Y2=0
cc_146 N_A_83_264#_c_121_n N_C_c_407_n 0.01791f $X=6.465 $Y=1.11 $X2=0 $Y2=0
cc_147 N_A_83_264#_c_124_n N_C_c_407_n 0.0293972f $X=4.935 $Y=0.875 $X2=0 $Y2=0
cc_148 N_A_83_264#_c_131_n N_C_c_407_n 0.0034967f $X=5.625 $Y=2.07 $X2=0 $Y2=0
cc_149 N_A_83_264#_c_120_n N_D_c_470_n 0.00358648f $X=4.935 $Y=0.515 $X2=-0.19
+ $Y2=-0.245
cc_150 N_A_83_264#_c_121_n N_D_c_470_n 0.0113592f $X=6.465 $Y=1.11 $X2=-0.19
+ $Y2=-0.245
cc_151 N_A_83_264#_c_124_n N_D_c_470_n 4.42511e-19 $X=4.935 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_152 N_A_83_264#_c_131_n N_D_M1000_g 0.00572858f $X=5.625 $Y=2.07 $X2=0 $Y2=0
cc_153 N_A_83_264#_c_129_n N_D_M1002_g 0.00875219f $X=6.465 $Y=2.035 $X2=0 $Y2=0
cc_154 N_A_83_264#_c_131_n N_D_M1002_g 0.00269754f $X=5.625 $Y=2.07 $X2=0 $Y2=0
cc_155 N_A_83_264#_c_121_n N_D_c_473_n 0.0105003f $X=6.465 $Y=1.11 $X2=0 $Y2=0
cc_156 N_A_83_264#_c_121_n N_D_c_474_n 0.0192499f $X=6.465 $Y=1.11 $X2=0 $Y2=0
cc_157 N_A_83_264#_c_121_n N_D_c_476_n 0.0120613f $X=6.465 $Y=1.11 $X2=0 $Y2=0
cc_158 N_A_83_264#_c_122_n N_D_c_476_n 0.00405285f $X=6.55 $Y=1.95 $X2=0 $Y2=0
cc_159 N_A_83_264#_c_131_n N_D_c_476_n 3.42297e-19 $X=5.625 $Y=2.07 $X2=0 $Y2=0
cc_160 N_A_83_264#_c_121_n N_D_c_478_n 0.0272875f $X=6.465 $Y=1.11 $X2=0 $Y2=0
cc_161 N_A_83_264#_M1005_g N_VPWR_c_528_n 0.013475f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_162 N_A_83_264#_M1006_g N_VPWR_c_528_n 5.02386e-19 $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_163 N_A_83_264#_M1005_g N_VPWR_c_529_n 5.02386e-19 $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_164 N_A_83_264#_M1006_g N_VPWR_c_529_n 0.012204f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_165 N_A_83_264#_M1008_g N_VPWR_c_529_n 0.012204f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_166 N_A_83_264#_M1011_g N_VPWR_c_529_n 5.02386e-19 $X=1.855 $Y=2.4 $X2=0
+ $Y2=0
cc_167 N_A_83_264#_M1008_g N_VPWR_c_530_n 5.02386e-19 $X=1.405 $Y=2.4 $X2=0
+ $Y2=0
cc_168 N_A_83_264#_M1011_g N_VPWR_c_530_n 0.0134762f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_169 N_A_83_264#_M1005_g N_VPWR_c_532_n 0.00460063f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_170 N_A_83_264#_M1006_g N_VPWR_c_532_n 0.00460063f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_171 N_A_83_264#_M1008_g N_VPWR_c_533_n 0.00460063f $X=1.405 $Y=2.4 $X2=0
+ $Y2=0
cc_172 N_A_83_264#_M1011_g N_VPWR_c_533_n 0.00460063f $X=1.855 $Y=2.4 $X2=0
+ $Y2=0
cc_173 N_A_83_264#_M1005_g N_VPWR_c_526_n 0.00908554f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_174 N_A_83_264#_M1006_g N_VPWR_c_526_n 0.00908554f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_175 N_A_83_264#_M1008_g N_VPWR_c_526_n 0.00908554f $X=1.405 $Y=2.4 $X2=0
+ $Y2=0
cc_176 N_A_83_264#_M1011_g N_VPWR_c_526_n 0.00908554f $X=1.855 $Y=2.4 $X2=0
+ $Y2=0
cc_177 N_A_83_264#_M1001_g N_X_c_612_n 0.00788812f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A_83_264#_M1007_g N_X_c_612_n 0.00926373f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A_83_264#_M1010_g N_X_c_612_n 6.73969e-19 $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_180 N_A_83_264#_M1005_g N_X_c_613_n 0.0326548f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A_83_264#_M1001_g N_X_c_613_n 0.0189011f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A_83_264#_M1006_g N_X_c_613_n 0.0144752f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_183 N_A_83_264#_M1007_g N_X_c_613_n 0.00535402f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_184 N_A_83_264#_M1010_g N_X_c_613_n 5.67152e-19 $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A_83_264#_c_117_n N_X_c_613_n 0.0147668f $X=2.155 $Y=1.485 $X2=0 $Y2=0
cc_186 N_A_83_264#_c_123_n N_X_c_613_n 0.0295009f $X=2.16 $Y=1.485 $X2=0 $Y2=0
cc_187 N_A_83_264#_M1005_g N_X_c_617_n 3.8104e-19 $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A_83_264#_M1006_g N_X_c_617_n 3.8104e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_189 N_A_83_264#_M1007_g N_X_c_614_n 0.0133712f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A_83_264#_M1010_g N_X_c_614_n 0.0155759f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_191 N_A_83_264#_M1012_g N_X_c_614_n 8.15014e-19 $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A_83_264#_c_117_n N_X_c_614_n 0.0497808f $X=2.155 $Y=1.485 $X2=0 $Y2=0
cc_193 N_A_83_264#_c_118_n N_X_c_614_n 0.00786297f $X=2.24 $Y=1.32 $X2=0 $Y2=0
cc_194 N_A_83_264#_c_123_n N_X_c_614_n 0.012612f $X=2.16 $Y=1.485 $X2=0 $Y2=0
cc_195 N_A_83_264#_M1008_g N_X_c_618_n 3.8104e-19 $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_196 N_A_83_264#_M1011_g N_X_c_618_n 3.8104e-19 $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_197 N_A_83_264#_M1010_g N_X_c_615_n 0.00516826f $X=1.495 $Y=0.74 $X2=0 $Y2=0
cc_198 N_A_83_264#_M1012_g N_X_c_615_n 0.00796805f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A_83_264#_c_117_n X 0.0193994f $X=2.155 $Y=1.485 $X2=0 $Y2=0
cc_200 N_A_83_264#_c_123_n X 0.00239242f $X=2.16 $Y=1.485 $X2=0 $Y2=0
cc_201 N_A_83_264#_M1011_g X 0.0225935f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_202 N_A_83_264#_c_117_n X 0.0316313f $X=2.155 $Y=1.485 $X2=0 $Y2=0
cc_203 N_A_83_264#_c_118_n X 0.0100698f $X=2.24 $Y=1.32 $X2=0 $Y2=0
cc_204 N_A_83_264#_c_123_n X 0.00593789f $X=2.16 $Y=1.485 $X2=0 $Y2=0
cc_205 N_A_83_264#_M1006_g N_X_c_621_n 0.0134181f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_206 N_A_83_264#_M1008_g N_X_c_621_n 0.0196409f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_207 N_A_83_264#_c_117_n N_X_c_621_n 0.0150496f $X=2.155 $Y=1.485 $X2=0 $Y2=0
cc_208 N_A_83_264#_c_123_n N_X_c_621_n 0.00233344f $X=2.16 $Y=1.485 $X2=0 $Y2=0
cc_209 N_A_83_264#_c_129_n N_A_499_392#_M1019_d 0.00424694f $X=6.465 $Y=2.035
+ $X2=0 $Y2=0
cc_210 N_A_83_264#_M1011_g N_A_499_392#_c_681_n 0.00189577f $X=1.855 $Y=2.4
+ $X2=0 $Y2=0
cc_211 N_A_83_264#_M1011_g N_A_499_392#_c_682_n 0.00316439f $X=1.855 $Y=2.4
+ $X2=0 $Y2=0
cc_212 N_A_83_264#_c_131_n N_A_499_392#_c_683_n 0.00537253f $X=5.625 $Y=2.07
+ $X2=0 $Y2=0
cc_213 N_A_83_264#_c_131_n N_A_499_392#_c_690_n 0.001246f $X=5.625 $Y=2.07 $X2=0
+ $Y2=0
cc_214 N_A_83_264#_M1000_d N_A_499_392#_c_691_n 0.00329665f $X=5.325 $Y=1.96
+ $X2=0 $Y2=0
cc_215 N_A_83_264#_c_129_n N_A_499_392#_c_691_n 0.0257153f $X=6.465 $Y=2.035
+ $X2=0 $Y2=0
cc_216 N_A_83_264#_c_131_n N_A_499_392#_c_691_n 0.0157372f $X=5.625 $Y=2.07
+ $X2=0 $Y2=0
cc_217 N_A_83_264#_c_129_n N_A_499_392#_c_685_n 0.0248692f $X=6.465 $Y=2.035
+ $X2=0 $Y2=0
cc_218 N_A_83_264#_c_129_n N_A_965_392#_M1002_s 0.00193659f $X=6.465 $Y=2.035
+ $X2=0 $Y2=0
cc_219 N_A_83_264#_M1000_d N_A_965_392#_c_779_n 0.0016881f $X=5.325 $Y=1.96
+ $X2=0 $Y2=0
cc_220 N_A_83_264#_c_134_p N_VGND_M1012_d 0.0122153f $X=2.92 $Y=0.875 $X2=0
+ $Y2=0
cc_221 N_A_83_264#_c_141_p N_VGND_M1013_d 0.0370525f $X=4.77 $Y=0.875 $X2=0
+ $Y2=0
cc_222 N_A_83_264#_c_121_n N_VGND_M1009_d 0.00286681f $X=6.465 $Y=1.11 $X2=0
+ $Y2=0
cc_223 N_A_83_264#_M1001_g N_VGND_c_793_n 0.0184904f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_224 N_A_83_264#_c_123_n N_VGND_c_793_n 2.14484e-19 $X=2.16 $Y=1.485 $X2=0
+ $Y2=0
cc_225 N_A_83_264#_M1007_g N_VGND_c_794_n 0.00417204f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_226 N_A_83_264#_M1010_g N_VGND_c_794_n 0.0125758f $X=1.495 $Y=0.74 $X2=0
+ $Y2=0
cc_227 N_A_83_264#_M1012_g N_VGND_c_795_n 0.00516167f $X=2.25 $Y=0.74 $X2=0
+ $Y2=0
cc_228 N_A_83_264#_c_134_p N_VGND_c_795_n 0.0282828f $X=2.92 $Y=0.875 $X2=0
+ $Y2=0
cc_229 N_A_83_264#_c_119_n N_VGND_c_795_n 0.0104464f $X=3.085 $Y=0.515 $X2=0
+ $Y2=0
cc_230 N_A_83_264#_M1001_g N_VGND_c_796_n 0.00434272f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_231 N_A_83_264#_M1007_g N_VGND_c_796_n 0.00434272f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_232 N_A_83_264#_M1010_g N_VGND_c_797_n 0.00383152f $X=1.495 $Y=0.74 $X2=0
+ $Y2=0
cc_233 N_A_83_264#_M1012_g N_VGND_c_797_n 0.00461464f $X=2.25 $Y=0.74 $X2=0
+ $Y2=0
cc_234 N_A_83_264#_M1001_g N_VGND_c_799_n 0.00823934f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_235 N_A_83_264#_M1007_g N_VGND_c_799_n 0.00820718f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_236 N_A_83_264#_M1010_g N_VGND_c_799_n 0.00759969f $X=1.495 $Y=0.74 $X2=0
+ $Y2=0
cc_237 N_A_83_264#_M1012_g N_VGND_c_799_n 0.0045489f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A_83_264#_c_134_p N_VGND_c_799_n 0.00886098f $X=2.92 $Y=0.875 $X2=0
+ $Y2=0
cc_239 N_A_83_264#_c_262_p N_VGND_c_799_n 0.00583874f $X=2.325 $Y=0.875 $X2=0
+ $Y2=0
cc_240 N_A_83_264#_c_119_n N_VGND_c_799_n 0.0118382f $X=3.085 $Y=0.515 $X2=0
+ $Y2=0
cc_241 N_A_83_264#_c_141_p N_VGND_c_799_n 0.0151942f $X=4.77 $Y=0.875 $X2=0
+ $Y2=0
cc_242 N_A_83_264#_c_120_n N_VGND_c_799_n 0.0119984f $X=4.935 $Y=0.515 $X2=0
+ $Y2=0
cc_243 N_A_83_264#_c_119_n N_VGND_c_802_n 0.014379f $X=3.085 $Y=0.515 $X2=0
+ $Y2=0
cc_244 N_A_83_264#_c_119_n N_VGND_c_803_n 0.010535f $X=3.085 $Y=0.515 $X2=0
+ $Y2=0
cc_245 N_A_83_264#_c_141_p N_VGND_c_803_n 0.091374f $X=4.77 $Y=0.875 $X2=0 $Y2=0
cc_246 N_A_83_264#_c_120_n N_VGND_c_803_n 0.010535f $X=4.935 $Y=0.515 $X2=0
+ $Y2=0
cc_247 N_A_83_264#_c_120_n N_VGND_c_804_n 0.0145639f $X=4.935 $Y=0.515 $X2=0
+ $Y2=0
cc_248 N_A_83_264#_c_120_n N_VGND_c_805_n 0.0146527f $X=4.935 $Y=0.515 $X2=0
+ $Y2=0
cc_249 N_A_83_264#_c_121_n N_VGND_c_805_n 0.0390715f $X=6.465 $Y=1.11 $X2=0
+ $Y2=0
cc_250 N_B_c_275_n N_A_M1013_g 0.013775f $X=2.87 $Y=1.22 $X2=0 $Y2=0
cc_251 N_B_c_277_n N_A_M1013_g 0.0118516f $X=4.065 $Y=1.215 $X2=0 $Y2=0
cc_252 N_B_c_278_n N_A_M1013_g 0.0120208f $X=3.235 $Y=1.215 $X2=0 $Y2=0
cc_253 N_B_c_279_n N_A_M1013_g 9.8879e-19 $X=4.23 $Y=1.215 $X2=0 $Y2=0
cc_254 N_B_c_280_n N_A_M1013_g 0.0040104f $X=4.23 $Y=1.385 $X2=0 $Y2=0
cc_255 N_B_M1014_g N_A_M1016_g 0.0215622f $X=2.865 $Y=2.46 $X2=0 $Y2=0
cc_256 N_B_c_273_n A 0.00117519f $X=2.865 $Y=1.64 $X2=0 $Y2=0
cc_257 N_B_M1018_g A 0.00124635f $X=4.235 $Y=2.46 $X2=0 $Y2=0
cc_258 N_B_c_277_n A 0.0247729f $X=4.065 $Y=1.215 $X2=0 $Y2=0
cc_259 N_B_c_278_n A 0.00633894f $X=3.235 $Y=1.215 $X2=0 $Y2=0
cc_260 N_B_c_279_n A 0.00352889f $X=4.23 $Y=1.215 $X2=0 $Y2=0
cc_261 N_B_c_280_n A 2.32886e-19 $X=4.23 $Y=1.385 $X2=0 $Y2=0
cc_262 N_B_c_273_n N_A_c_358_n 0.0353371f $X=2.865 $Y=1.64 $X2=0 $Y2=0
cc_263 N_B_M1018_g N_A_c_358_n 0.0380832f $X=4.235 $Y=2.46 $X2=0 $Y2=0
cc_264 N_B_c_277_n N_A_c_358_n 0.00704512f $X=4.065 $Y=1.215 $X2=0 $Y2=0
cc_265 N_B_c_278_n N_A_c_358_n 0.00241908f $X=3.235 $Y=1.215 $X2=0 $Y2=0
cc_266 N_B_c_279_n N_A_c_358_n 3.40206e-19 $X=4.23 $Y=1.215 $X2=0 $Y2=0
cc_267 N_B_c_280_n N_A_c_358_n 0.00523467f $X=4.23 $Y=1.385 $X2=0 $Y2=0
cc_268 N_B_c_279_n N_C_M1015_g 0.00316947f $X=4.23 $Y=1.215 $X2=0 $Y2=0
cc_269 N_B_c_280_n N_C_M1015_g 0.0114999f $X=4.23 $Y=1.385 $X2=0 $Y2=0
cc_270 N_B_M1018_g N_C_M1003_g 0.0142312f $X=4.235 $Y=2.46 $X2=0 $Y2=0
cc_271 N_B_M1018_g N_C_c_404_n 0.00926972f $X=4.235 $Y=2.46 $X2=0 $Y2=0
cc_272 N_B_c_280_n N_C_c_404_n 0.00691933f $X=4.23 $Y=1.385 $X2=0 $Y2=0
cc_273 N_B_M1018_g N_C_c_407_n 0.00138903f $X=4.235 $Y=2.46 $X2=0 $Y2=0
cc_274 N_B_c_279_n N_C_c_407_n 0.012807f $X=4.23 $Y=1.215 $X2=0 $Y2=0
cc_275 N_B_c_280_n N_C_c_407_n 8.90064e-19 $X=4.23 $Y=1.385 $X2=0 $Y2=0
cc_276 N_B_M1014_g N_VPWR_c_530_n 0.00395619f $X=2.865 $Y=2.46 $X2=0 $Y2=0
cc_277 N_B_M1014_g N_VPWR_c_531_n 6.13527e-19 $X=2.865 $Y=2.46 $X2=0 $Y2=0
cc_278 N_B_M1018_g N_VPWR_c_531_n 6.12882e-19 $X=4.235 $Y=2.46 $X2=0 $Y2=0
cc_279 N_B_M1014_g N_VPWR_c_534_n 0.005209f $X=2.865 $Y=2.46 $X2=0 $Y2=0
cc_280 N_B_M1018_g N_VPWR_c_535_n 0.005209f $X=4.235 $Y=2.46 $X2=0 $Y2=0
cc_281 N_B_M1014_g N_VPWR_c_526_n 0.00988607f $X=2.865 $Y=2.46 $X2=0 $Y2=0
cc_282 N_B_M1018_g N_VPWR_c_526_n 0.00984228f $X=4.235 $Y=2.46 $X2=0 $Y2=0
cc_283 N_B_M1014_g X 0.00396899f $X=2.865 $Y=2.46 $X2=0 $Y2=0
cc_284 N_B_c_273_n N_A_499_392#_c_681_n 0.00111452f $X=2.865 $Y=1.64 $X2=0 $Y2=0
cc_285 N_B_M1014_g N_A_499_392#_c_681_n 0.00438165f $X=2.865 $Y=2.46 $X2=0 $Y2=0
cc_286 N_B_c_278_n N_A_499_392#_c_681_n 0.012069f $X=3.235 $Y=1.215 $X2=0 $Y2=0
cc_287 N_B_M1014_g N_A_499_392#_c_682_n 4.78926e-19 $X=2.865 $Y=2.46 $X2=0 $Y2=0
cc_288 N_B_M1014_g N_A_499_392#_c_699_n 0.0133421f $X=2.865 $Y=2.46 $X2=0 $Y2=0
cc_289 N_B_M1018_g N_A_499_392#_c_699_n 0.0158765f $X=4.235 $Y=2.46 $X2=0 $Y2=0
cc_290 N_B_c_277_n N_A_499_392#_c_699_n 0.0118008f $X=4.065 $Y=1.215 $X2=0 $Y2=0
cc_291 N_B_c_278_n N_A_499_392#_c_699_n 0.0147824f $X=3.235 $Y=1.215 $X2=0 $Y2=0
cc_292 N_B_c_279_n N_A_499_392#_c_699_n 0.00858702f $X=4.23 $Y=1.215 $X2=0 $Y2=0
cc_293 N_B_c_280_n N_A_499_392#_c_699_n 2.76808e-19 $X=4.23 $Y=1.385 $X2=0 $Y2=0
cc_294 N_B_M1018_g N_A_499_392#_c_683_n 5.59553e-19 $X=4.235 $Y=2.46 $X2=0 $Y2=0
cc_295 N_B_c_279_n N_A_499_392#_c_683_n 0.0022688f $X=4.23 $Y=1.215 $X2=0 $Y2=0
cc_296 N_B_c_280_n N_A_499_392#_c_683_n 3.46941e-19 $X=4.23 $Y=1.385 $X2=0 $Y2=0
cc_297 N_B_M1014_g N_A_591_392#_c_753_n 0.00282106f $X=2.865 $Y=2.46 $X2=0 $Y2=0
cc_298 N_B_M1014_g N_A_591_392#_c_751_n 0.0053845f $X=2.865 $Y=2.46 $X2=0 $Y2=0
cc_299 N_B_M1018_g N_A_591_392#_c_755_n 0.00323047f $X=4.235 $Y=2.46 $X2=0 $Y2=0
cc_300 N_B_M1018_g N_A_591_392#_c_752_n 0.00548193f $X=4.235 $Y=2.46 $X2=0 $Y2=0
cc_301 N_B_c_275_n N_VGND_c_795_n 0.00508528f $X=2.87 $Y=1.22 $X2=0 $Y2=0
cc_302 N_B_c_275_n N_VGND_c_799_n 0.00436349f $X=2.87 $Y=1.22 $X2=0 $Y2=0
cc_303 N_B_c_275_n N_VGND_c_802_n 0.00434272f $X=2.87 $Y=1.22 $X2=0 $Y2=0
cc_304 N_A_M1016_g N_VPWR_c_531_n 0.00741692f $X=3.315 $Y=2.46 $X2=0 $Y2=0
cc_305 N_A_M1017_g N_VPWR_c_531_n 0.00757291f $X=3.765 $Y=2.46 $X2=0 $Y2=0
cc_306 N_A_M1016_g N_VPWR_c_534_n 0.00460063f $X=3.315 $Y=2.46 $X2=0 $Y2=0
cc_307 N_A_M1017_g N_VPWR_c_535_n 0.00460063f $X=3.765 $Y=2.46 $X2=0 $Y2=0
cc_308 N_A_M1016_g N_VPWR_c_526_n 0.00443357f $X=3.315 $Y=2.46 $X2=0 $Y2=0
cc_309 N_A_M1017_g N_VPWR_c_526_n 0.00443494f $X=3.765 $Y=2.46 $X2=0 $Y2=0
cc_310 N_A_M1016_g N_A_499_392#_c_681_n 3.81471e-19 $X=3.315 $Y=2.46 $X2=0 $Y2=0
cc_311 N_A_M1016_g N_A_499_392#_c_699_n 0.0145647f $X=3.315 $Y=2.46 $X2=0 $Y2=0
cc_312 N_A_M1017_g N_A_499_392#_c_699_n 0.0135178f $X=3.765 $Y=2.46 $X2=0 $Y2=0
cc_313 A N_A_499_392#_c_699_n 0.0200765f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_314 N_A_c_358_n N_A_499_392#_c_699_n 6.34453e-19 $X=3.765 $Y=1.635 $X2=0
+ $Y2=0
cc_315 N_A_M1016_g N_A_591_392#_c_757_n 0.0121339f $X=3.315 $Y=2.46 $X2=0 $Y2=0
cc_316 N_A_M1017_g N_A_591_392#_c_757_n 0.0104445f $X=3.765 $Y=2.46 $X2=0 $Y2=0
cc_317 N_A_M1016_g N_A_591_392#_c_755_n 2.38225e-19 $X=3.315 $Y=2.46 $X2=0 $Y2=0
cc_318 N_A_M1017_g N_A_591_392#_c_755_n 0.00256315f $X=3.765 $Y=2.46 $X2=0 $Y2=0
cc_319 N_A_M1017_g N_A_591_392#_c_752_n 3.01048e-19 $X=3.765 $Y=2.46 $X2=0 $Y2=0
cc_320 N_A_M1013_g N_VGND_c_799_n 0.00439727f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_321 N_A_M1013_g N_VGND_c_802_n 0.00434272f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_322 N_A_M1013_g N_VGND_c_803_n 0.0103115f $X=3.3 $Y=0.74 $X2=0 $Y2=0
cc_323 N_C_M1015_g N_D_c_470_n 0.0280437f $X=4.72 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_324 N_C_M1003_g N_D_M1000_g 0.039082f $X=4.735 $Y=2.46 $X2=0 $Y2=0
cc_325 N_C_c_407_n N_D_M1000_g 0.0156495f $X=5.34 $Y=1.572 $X2=0 $Y2=0
cc_326 N_C_M1019_g N_D_M1002_g 0.0476229f $X=6.135 $Y=2.46 $X2=0 $Y2=0
cc_327 N_C_c_406_n N_D_M1002_g 0.0135482f $X=6.15 $Y=1.53 $X2=0 $Y2=0
cc_328 N_C_c_405_n N_D_c_474_n 0.00672114f $X=6.15 $Y=1.53 $X2=0 $Y2=0
cc_329 N_C_c_404_n N_D_c_476_n 0.0213325f $X=4.77 $Y=1.605 $X2=0 $Y2=0
cc_330 N_C_c_405_n N_D_c_476_n 0.0268774f $X=6.15 $Y=1.53 $X2=0 $Y2=0
cc_331 N_C_c_406_n N_D_c_476_n 0.0139321f $X=6.15 $Y=1.53 $X2=0 $Y2=0
cc_332 N_C_c_407_n N_D_c_476_n 0.00645108f $X=5.34 $Y=1.572 $X2=0 $Y2=0
cc_333 N_C_M1003_g N_VPWR_c_535_n 0.005209f $X=4.735 $Y=2.46 $X2=0 $Y2=0
cc_334 N_C_M1019_g N_VPWR_c_535_n 0.00519794f $X=6.135 $Y=2.46 $X2=0 $Y2=0
cc_335 N_C_M1003_g N_VPWR_c_526_n 0.00525164f $X=4.735 $Y=2.46 $X2=0 $Y2=0
cc_336 N_C_M1019_g N_VPWR_c_526_n 0.00529098f $X=6.135 $Y=2.46 $X2=0 $Y2=0
cc_337 N_C_M1003_g N_A_499_392#_c_683_n 0.00469374f $X=4.735 $Y=2.46 $X2=0 $Y2=0
cc_338 N_C_c_404_n N_A_499_392#_c_683_n 3.16589e-19 $X=4.77 $Y=1.605 $X2=0 $Y2=0
cc_339 N_C_c_407_n N_A_499_392#_c_683_n 0.00588104f $X=5.34 $Y=1.572 $X2=0 $Y2=0
cc_340 N_C_M1003_g N_A_499_392#_c_690_n 0.00433969f $X=4.735 $Y=2.46 $X2=0 $Y2=0
cc_341 N_C_M1003_g N_A_499_392#_c_684_n 0.00700212f $X=4.735 $Y=2.46 $X2=0 $Y2=0
cc_342 N_C_M1003_g N_A_499_392#_c_691_n 0.0118812f $X=4.735 $Y=2.46 $X2=0 $Y2=0
cc_343 N_C_M1019_g N_A_499_392#_c_691_n 0.0113948f $X=6.135 $Y=2.46 $X2=0 $Y2=0
cc_344 N_C_c_404_n N_A_499_392#_c_691_n 3.81825e-19 $X=4.77 $Y=1.605 $X2=0 $Y2=0
cc_345 N_C_c_407_n N_A_499_392#_c_691_n 0.0162987f $X=5.34 $Y=1.572 $X2=0 $Y2=0
cc_346 N_C_M1003_g N_A_499_392#_c_722_n 4.64231e-19 $X=4.735 $Y=2.46 $X2=0 $Y2=0
cc_347 N_C_M1019_g N_A_499_392#_c_685_n 5.01354e-19 $X=6.135 $Y=2.46 $X2=0 $Y2=0
cc_348 N_C_M1019_g N_A_965_392#_c_779_n 0.00418558f $X=6.135 $Y=2.46 $X2=0 $Y2=0
cc_349 N_C_M1015_g N_VGND_c_799_n 0.00440341f $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_350 N_C_M1015_g N_VGND_c_803_n 0.00868136f $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_351 N_C_M1015_g N_VGND_c_804_n 0.00434272f $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_352 N_C_M1015_g N_VGND_c_805_n 4.32194e-19 $X=4.72 $Y=0.74 $X2=0 $Y2=0
cc_353 N_D_M1000_g N_VPWR_c_535_n 0.00349978f $X=5.235 $Y=2.46 $X2=0 $Y2=0
cc_354 N_D_M1002_g N_VPWR_c_535_n 0.00349978f $X=5.685 $Y=2.46 $X2=0 $Y2=0
cc_355 N_D_M1000_g N_VPWR_c_526_n 0.00430085f $X=5.235 $Y=2.46 $X2=0 $Y2=0
cc_356 N_D_M1002_g N_VPWR_c_526_n 0.00429629f $X=5.685 $Y=2.46 $X2=0 $Y2=0
cc_357 N_D_M1000_g N_A_499_392#_c_683_n 6.22289e-19 $X=5.235 $Y=2.46 $X2=0 $Y2=0
cc_358 N_D_M1000_g N_A_499_392#_c_690_n 9.44887e-19 $X=5.235 $Y=2.46 $X2=0 $Y2=0
cc_359 N_D_M1000_g N_A_499_392#_c_684_n 6.53319e-19 $X=5.235 $Y=2.46 $X2=0 $Y2=0
cc_360 N_D_M1000_g N_A_499_392#_c_691_n 0.0138666f $X=5.235 $Y=2.46 $X2=0 $Y2=0
cc_361 N_D_M1002_g N_A_499_392#_c_691_n 0.0120289f $X=5.685 $Y=2.46 $X2=0 $Y2=0
cc_362 N_D_M1000_g N_A_965_392#_c_779_n 0.0123947f $X=5.235 $Y=2.46 $X2=0 $Y2=0
cc_363 N_D_M1002_g N_A_965_392#_c_779_n 0.0123953f $X=5.685 $Y=2.46 $X2=0 $Y2=0
cc_364 N_D_c_474_n N_VGND_c_798_n 0.0025954f $X=6.285 $Y=0.85 $X2=0 $Y2=0
cc_365 N_D_c_477_n N_VGND_c_798_n 0.00213166f $X=6.45 $Y=0.42 $X2=0 $Y2=0
cc_366 N_D_c_478_n N_VGND_c_798_n 0.0221582f $X=6.45 $Y=0.42 $X2=0 $Y2=0
cc_367 N_D_c_470_n N_VGND_c_799_n 0.00753637f $X=5.22 $Y=1.185 $X2=0 $Y2=0
cc_368 N_D_c_474_n N_VGND_c_799_n 0.00358943f $X=6.285 $Y=0.85 $X2=0 $Y2=0
cc_369 N_D_c_478_n N_VGND_c_799_n 0.0125166f $X=6.45 $Y=0.42 $X2=0 $Y2=0
cc_370 N_D_c_470_n N_VGND_c_804_n 0.00230732f $X=5.22 $Y=1.185 $X2=0 $Y2=0
cc_371 N_D_c_470_n N_VGND_c_805_n 0.00971517f $X=5.22 $Y=1.185 $X2=0 $Y2=0
cc_372 N_D_c_475_n N_VGND_c_805_n 0.013425f $X=5.775 $Y=0.85 $X2=0 $Y2=0
cc_373 N_D_c_476_n N_VGND_c_805_n 8.10942e-19 $X=5.7 $Y=1.335 $X2=0 $Y2=0
cc_374 N_D_c_477_n N_VGND_c_805_n 0.00987736f $X=6.45 $Y=0.42 $X2=0 $Y2=0
cc_375 N_D_c_478_n N_VGND_c_805_n 0.0357573f $X=6.45 $Y=0.42 $X2=0 $Y2=0
cc_376 N_VPWR_M1005_s N_X_c_613_n 0.00418363f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_377 N_VPWR_c_528_n N_X_c_613_n 0.0234556f $X=0.28 $Y=2.405 $X2=0 $Y2=0
cc_378 N_VPWR_c_528_n N_X_c_617_n 0.0255132f $X=0.28 $Y=2.405 $X2=0 $Y2=0
cc_379 N_VPWR_c_529_n N_X_c_617_n 0.0255132f $X=1.18 $Y=2.405 $X2=0 $Y2=0
cc_380 N_VPWR_c_532_n N_X_c_617_n 0.0101736f $X=1.015 $Y=3.33 $X2=0 $Y2=0
cc_381 N_VPWR_c_526_n N_X_c_617_n 0.0084208f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_382 N_VPWR_c_529_n N_X_c_618_n 0.0255132f $X=1.18 $Y=2.405 $X2=0 $Y2=0
cc_383 N_VPWR_c_530_n N_X_c_618_n 0.0255132f $X=2.08 $Y=2.405 $X2=0 $Y2=0
cc_384 N_VPWR_c_533_n N_X_c_618_n 0.0101736f $X=1.915 $Y=3.33 $X2=0 $Y2=0
cc_385 N_VPWR_c_526_n N_X_c_618_n 0.0084208f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_386 N_VPWR_M1011_s X 0.00412975f $X=1.945 $Y=1.84 $X2=0 $Y2=0
cc_387 N_VPWR_c_530_n X 0.0229451f $X=2.08 $Y=2.405 $X2=0 $Y2=0
cc_388 N_VPWR_M1006_s N_X_c_621_n 0.00169251f $X=1.045 $Y=1.84 $X2=0 $Y2=0
cc_389 N_VPWR_c_529_n N_X_c_621_n 0.0178311f $X=1.18 $Y=2.405 $X2=0 $Y2=0
cc_390 N_VPWR_c_530_n N_A_499_392#_c_682_n 0.0439497f $X=2.08 $Y=2.405 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_534_n N_A_499_392#_c_682_n 0.0124046f $X=3.375 $Y=3.33 $X2=0
+ $Y2=0
cc_392 N_VPWR_c_526_n N_A_499_392#_c_682_n 0.0102675f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_393 N_VPWR_M1016_d N_A_499_392#_c_699_n 0.00331313f $X=3.405 $Y=1.96 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_535_n N_A_499_392#_c_684_n 0.014549f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_395 N_VPWR_c_526_n N_A_499_392#_c_684_n 0.0119743f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_526_n N_A_499_392#_c_691_n 0.0116647f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_535_n N_A_499_392#_c_685_n 0.0146513f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_526_n N_A_499_392#_c_685_n 0.0121202f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_531_n N_A_591_392#_c_751_n 0.0101517f $X=3.54 $Y=2.815 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_534_n N_A_591_392#_c_751_n 0.0122358f $X=3.375 $Y=3.33 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_526_n N_A_591_392#_c_751_n 0.0100955f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_402 N_VPWR_M1016_d N_A_591_392#_c_757_n 0.00339373f $X=3.405 $Y=1.96 $X2=0
+ $Y2=0
cc_403 N_VPWR_c_531_n N_A_591_392#_c_757_n 0.016727f $X=3.54 $Y=2.815 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_526_n N_A_591_392#_c_757_n 0.00999888f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_526_n N_A_591_392#_c_755_n 0.00241362f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_531_n N_A_591_392#_c_752_n 0.00929382f $X=3.54 $Y=2.815 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_535_n N_A_591_392#_c_752_n 0.0123047f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_408 N_VPWR_c_526_n N_A_591_392#_c_752_n 0.0101224f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_409 N_VPWR_c_535_n N_A_965_392#_c_779_n 0.0502919f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_526_n N_A_965_392#_c_779_n 0.0422533f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_411 X N_A_499_392#_c_681_n 0.0172799f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_412 N_X_c_614_n N_VGND_M1007_d 0.00250873f $X=1.615 $Y=1.065 $X2=0 $Y2=0
cc_413 N_X_c_612_n N_VGND_c_793_n 0.0243921f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_414 N_X_c_613_n N_VGND_c_793_n 0.0370015f $X=0.73 $Y=2.15 $X2=0 $Y2=0
cc_415 N_X_c_612_n N_VGND_c_794_n 0.0180508f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_416 N_X_c_614_n N_VGND_c_794_n 0.0210288f $X=1.615 $Y=1.065 $X2=0 $Y2=0
cc_417 N_X_c_615_n N_VGND_c_794_n 0.0180508f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_418 N_X_c_615_n N_VGND_c_795_n 0.00585761f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_419 N_X_c_612_n N_VGND_c_796_n 0.0144922f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_420 N_X_c_615_n N_VGND_c_797_n 0.0146357f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_421 N_X_c_612_n N_VGND_c_799_n 0.0118826f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_422 N_X_c_615_n N_VGND_c_799_n 0.0121141f $X=1.78 $Y=0.515 $X2=0 $Y2=0
cc_423 N_A_499_392#_c_699_n N_A_591_392#_M1014_d 0.00442093f $X=4.345 $Y=2.055
+ $X2=-0.19 $Y2=1.66
cc_424 N_A_499_392#_c_699_n N_A_591_392#_M1017_s 0.00539923f $X=4.345 $Y=2.055
+ $X2=0 $Y2=0
cc_425 N_A_499_392#_c_699_n N_A_591_392#_c_753_n 0.01221f $X=4.345 $Y=2.055
+ $X2=0 $Y2=0
cc_426 N_A_499_392#_c_682_n N_A_591_392#_c_751_n 0.0161022f $X=2.64 $Y=2.445
+ $X2=0 $Y2=0
cc_427 N_A_499_392#_c_699_n N_A_591_392#_c_757_n 0.0278551f $X=4.345 $Y=2.055
+ $X2=0 $Y2=0
cc_428 N_A_499_392#_c_699_n N_A_591_392#_c_755_n 0.0186128f $X=4.345 $Y=2.055
+ $X2=0 $Y2=0
cc_429 N_A_499_392#_c_684_n N_A_591_392#_c_752_n 0.0161216f $X=4.51 $Y=2.815
+ $X2=0 $Y2=0
cc_430 N_A_499_392#_c_691_n N_A_965_392#_M1003_s 0.00604471f $X=6.245 $Y=2.445
+ $X2=-0.19 $Y2=1.66
cc_431 N_A_499_392#_c_691_n N_A_965_392#_M1002_s 0.00353365f $X=6.245 $Y=2.445
+ $X2=0 $Y2=0
cc_432 N_A_499_392#_c_684_n N_A_965_392#_c_779_n 0.0113199f $X=4.51 $Y=2.815
+ $X2=0 $Y2=0
cc_433 N_A_499_392#_c_691_n N_A_965_392#_c_779_n 0.0646086f $X=6.245 $Y=2.445
+ $X2=0 $Y2=0
cc_434 N_A_499_392#_c_685_n N_A_965_392#_c_779_n 0.0124625f $X=6.41 $Y=2.455
+ $X2=0 $Y2=0

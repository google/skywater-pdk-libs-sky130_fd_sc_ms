* File: sky130_fd_sc_ms__dfrtp_1.spice
* Created: Fri Aug 28 17:22:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dfrtp_1.pex.spice"
.subckt sky130_fd_sc_ms__dfrtp_1  VNB VPB D CLK RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* CLK	CLK
* D	D
* VPB	VPB
* VNB	VNB
MM1026 A_117_78# N_D_M1026_g N_A_30_78#_M1026_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_RESET_B_M1009_g A_117_78# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_CLK_M1023_g N_A_299_387#_M1023_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.13745 AS=0.245475 PD=1.115 PS=2.15 NRD=7.296 NRS=7.296 M=1
+ R=4.93333 SA=75000.3 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1001 N_A_493_387#_M1001_d N_A_299_387#_M1001_g N_VGND_M1023_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2262 AS=0.13745 PD=2.14 PS=1.115 NRD=4.044 NRS=7.296 M=1
+ R=4.93333 SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_A_701_463#_M1007_d N_A_299_387#_M1007_g N_A_30_78#_M1007_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.07035 AS=0.1344 PD=0.755 PS=1.48 NRD=8.568 NRS=11.424 M=1
+ R=2.8 SA=75000.2 SB=75003.6 A=0.063 P=1.14 MULT=1
MM1002 A_821_138# N_A_493_387#_M1002_g N_A_701_463#_M1007_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.04515 AS=0.07035 PD=0.635 PS=0.755 NRD=14.988 NRS=7.14 M=1 R=2.8
+ SA=75000.7 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1012 A_894_138# N_A_833_400#_M1012_g A_821_138# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.04515 PD=0.66 PS=0.635 NRD=18.564 NRS=14.988 M=1 R=2.8
+ SA=75001.1 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_RESET_B_M1006_g A_894_138# VNB NLOWVT L=0.15 W=0.42
+ AD=0.152965 AS=0.0504 PD=1.05 PS=0.66 NRD=88.332 NRS=18.564 M=1 R=2.8
+ SA=75001.5 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1031 N_A_833_400#_M1031_d N_A_701_463#_M1031_g N_VGND_M1006_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.24605 AS=0.26951 PD=1.405 PS=1.85 NRD=22.296 NRS=50.136 M=1
+ R=4.93333 SA=75001.4 SB=75002.3 A=0.111 P=1.78 MULT=1
MM1027 N_A_1266_74#_M1027_d N_A_493_387#_M1027_g N_A_833_400#_M1031_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.292172 AS=0.24605 PD=2.09241 PS=1.405 NRD=2.424 NRS=8.916
+ M=1 R=4.93333 SA=75002.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1016 A_1476_81# N_A_299_387#_M1016_g N_A_1266_74#_M1027_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.165828 PD=0.66 PS=1.18759 NRD=18.564 NRS=49.992 M=1
+ R=2.8 SA=75002.8 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_1518_203#_M1013_g A_1476_81# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0756 AS=0.0504 PD=0.78 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75003.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 A_1656_81# N_RESET_B_M1000_g N_VGND_M1013_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0756 PD=0.63 PS=0.78 NRD=14.28 NRS=22.848 M=1 R=2.8 SA=75003.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1017 N_A_1518_203#_M1017_d N_A_1266_74#_M1017_g A_1656_81# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75004.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1028 N_A_1867_409#_M1028_d N_A_1266_74#_M1028_g N_VGND_M1028_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.15675 AS=0.15675 PD=1.67 PS=1.67 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1003 N_VGND_M1003_d N_A_1867_409#_M1003_g N_Q_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1018 N_A_30_78#_M1018_d N_D_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.18 W=0.42
+ AD=0.0567 AS=0.1134 PD=0.69 PS=1.38 NRD=0 NRS=0 M=1 R=2.33333 SA=90000.2
+ SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1019 N_VPWR_M1019_d N_RESET_B_M1019_g N_A_30_78#_M1018_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1176 AS=0.0567 PD=1.4 PS=0.69 NRD=0 NRS=0 M=1 R=2.33333 SA=90000.6
+ SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1021 N_VPWR_M1021_d N_CLK_M1021_g N_A_299_387#_M1021_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.31375 PD=1.39 PS=2.92 NRD=0 NRS=13.1793 M=1 R=6.22222
+ SA=90000.2 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1025 N_A_493_387#_M1025_d N_A_299_387#_M1025_g N_VPWR_M1021_d VPB PSHORT
+ L=0.18 W=1.12 AD=0.3024 AS=0.1512 PD=2.78 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1014 N_A_701_463#_M1014_d N_A_493_387#_M1014_g N_A_30_78#_M1014_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0567 AS=0.1176 PD=0.69 PS=1.4 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90001.6 A=0.0756 P=1.2 MULT=1
MM1022 A_791_463# N_A_299_387#_M1022_g N_A_701_463#_M1014_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0441 AS=0.0567 PD=0.63 PS=0.69 NRD=23.443 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1008 N_VPWR_M1008_d N_A_833_400#_M1008_g A_791_463# VPB PSHORT L=0.18 W=0.42
+ AD=0.123625 AS=0.0441 PD=1.095 PS=0.63 NRD=112.251 NRS=23.443 M=1 R=2.33333
+ SA=90001 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1030 N_A_701_463#_M1030_d N_RESET_B_M1030_g N_VPWR_M1008_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1176 AS=0.123625 PD=1.4 PS=1.095 NRD=0 NRS=112.251 M=1 R=2.33333
+ SA=90001.6 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1029 N_A_833_400#_M1029_d N_A_701_463#_M1029_g N_VPWR_M1029_s VPB PSHORT
+ L=0.18 W=1 AD=0.175625 AS=0.29 PD=1.475 PS=2.58 NRD=6.8753 NRS=0.9653 M=1
+ R=5.55556 SA=90000.2 SB=90001.4 A=0.18 P=2.36 MULT=1
MM1004 N_A_1266_74#_M1004_d N_A_299_387#_M1004_g N_A_833_400#_M1029_d VPB PSHORT
+ L=0.18 W=1 AD=0.309155 AS=0.175625 PD=2.39437 PS=1.475 NRD=5.8903 NRS=1.9503
+ M=1 R=5.55556 SA=90000.6 SB=90001.4 A=0.18 P=2.36 MULT=1
MM1010 A_1471_493# N_A_493_387#_M1010_g N_A_1266_74#_M1004_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.129845 PD=0.66 PS=1.00563 NRD=30.4759 NRS=0 M=1
+ R=2.33333 SA=90001.4 SB=90002.2 A=0.0756 P=1.2 MULT=1
MM1015 N_VPWR_M1015_d N_A_1518_203#_M1015_g A_1471_493# VPB PSHORT L=0.18 W=0.42
+ AD=0.08295 AS=0.0504 PD=0.815 PS=0.66 NRD=25.7873 NRS=30.4759 M=1 R=2.33333
+ SA=90001.8 SB=90001.8 A=0.0756 P=1.2 MULT=1
MM1020 N_A_1518_203#_M1020_d N_RESET_B_M1020_g N_VPWR_M1015_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0567 AS=0.08295 PD=0.69 PS=0.815 NRD=0 NRS=28.1316 M=1 R=2.33333
+ SA=90002.4 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1024 N_VPWR_M1024_d N_A_1266_74#_M1024_g N_A_1518_203#_M1020_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.0889 AS=0.0567 PD=0.796667 PS=0.69 NRD=37.5088 NRS=0 M=1
+ R=2.33333 SA=90002.8 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1011 N_A_1867_409#_M1011_d N_A_1266_74#_M1011_g N_VPWR_M1024_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2352 AS=0.1778 PD=2.24 PS=1.59333 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90001.8 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1005 N_VPWR_M1005_d N_A_1867_409#_M1005_g N_Q_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3192 AS=0.364 PD=2.81 PS=2.89 NRD=0 NRS=7.0329 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX32_noxref VNB VPB NWDIODE A=20.9584 P=26.96
c_231 VPB 0 1.4888e-19 $X=0 $Y=3.085
c_1682 A_1471_493# 0 1.00866e-19 $X=7.355 $Y=2.465
*
.include "sky130_fd_sc_ms__dfrtp_1.pxi.spice"
*
.ends
*
*

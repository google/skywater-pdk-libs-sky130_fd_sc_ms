* File: sky130_fd_sc_ms__o2bb2a_4.pex.spice
* Created: Wed Sep  2 12:24:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O2BB2A_4%B1 3 7 11 15 17 18 28 29
c56 11 0 1.0107e-19 $X=1.025 $Y=2.46
c57 3 0 1.72779e-19 $X=0.495 $Y=0.69
r58 29 30 5.93231 $w=3.25e-07 $l=4e-08 $layer=POLY_cond $X=1.025 $Y=1.425
+ $X2=1.065 $Y2=1.425
r59 27 29 11.1231 $w=3.25e-07 $l=7.5e-08 $layer=POLY_cond $X=0.95 $Y=1.425
+ $X2=1.025 $Y2=1.425
r60 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.95
+ $Y=1.425 $X2=0.95 $Y2=1.425
r61 25 27 55.6154 $w=3.25e-07 $l=3.75e-07 $layer=POLY_cond $X=0.575 $Y=1.425
+ $X2=0.95 $Y2=1.425
r62 24 25 11.8646 $w=3.25e-07 $l=8e-08 $layer=POLY_cond $X=0.495 $Y=1.425
+ $X2=0.575 $Y2=1.425
r63 22 24 33.3692 $w=3.25e-07 $l=2.25e-07 $layer=POLY_cond $X=0.27 $Y=1.425
+ $X2=0.495 $Y2=1.425
r64 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.425 $X2=0.27 $Y2=1.425
r65 18 28 5.39408 $w=5.08e-07 $l=2.3e-07 $layer=LI1_cond $X=0.72 $Y=1.515
+ $X2=0.95 $Y2=1.515
r66 18 23 10.5536 $w=5.08e-07 $l=4.5e-07 $layer=LI1_cond $X=0.72 $Y=1.515
+ $X2=0.27 $Y2=1.515
r67 17 23 0.703576 $w=5.08e-07 $l=3e-08 $layer=LI1_cond $X=0.24 $Y=1.515
+ $X2=0.27 $Y2=1.515
r68 13 30 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=1.26
+ $X2=1.065 $Y2=1.425
r69 13 15 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.065 $Y=1.26
+ $X2=1.065 $Y2=0.69
r70 9 29 16.5763 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.025 $Y=1.59
+ $X2=1.025 $Y2=1.425
r71 9 11 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=1.025 $Y=1.59
+ $X2=1.025 $Y2=2.46
r72 5 25 16.5763 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.575 $Y=1.59
+ $X2=0.575 $Y2=1.425
r73 5 7 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=0.575 $Y=1.59
+ $X2=0.575 $Y2=2.46
r74 1 24 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.26
+ $X2=0.495 $Y2=1.425
r75 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=0.495 $Y=1.26
+ $X2=0.495 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2A_4%B2 3 7 11 15 17 18 28
c56 28 0 1.82144e-19 $X=1.995 $Y=1.615
c57 18 0 5.33865e-20 $X=2.16 $Y=1.665
c58 11 0 5.55308e-20 $X=1.925 $Y=2.46
c59 3 0 8.35716e-20 $X=1.475 $Y=2.46
r60 26 28 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.975 $Y=1.615
+ $X2=1.995 $Y2=1.615
r61 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.975
+ $Y=1.615 $X2=1.975 $Y2=1.615
r62 24 26 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=1.925 $Y=1.615
+ $X2=1.975 $Y2=1.615
r63 23 24 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.495 $Y=1.615
+ $X2=1.925 $Y2=1.615
r64 21 23 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.475 $Y=1.615
+ $X2=1.495 $Y2=1.615
r65 18 27 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.16 $Y=1.615
+ $X2=1.975 $Y2=1.615
r66 17 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.68 $Y=1.615
+ $X2=1.975 $Y2=1.615
r67 13 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.995 $Y=1.45
+ $X2=1.995 $Y2=1.615
r68 13 15 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.995 $Y=1.45
+ $X2=1.995 $Y2=0.69
r69 9 24 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.78
+ $X2=1.925 $Y2=1.615
r70 9 11 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=1.925 $Y=1.78
+ $X2=1.925 $Y2=2.46
r71 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.495 $Y=1.45
+ $X2=1.495 $Y2=1.615
r72 5 7 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.495 $Y=1.45
+ $X2=1.495 $Y2=0.69
r73 1 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.475 $Y=1.78
+ $X2=1.475 $Y2=1.615
r74 1 3 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=1.475 $Y=1.78
+ $X2=1.475 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2A_4%A_476_48# 1 2 9 13 17 19 21 22 23 31 32 34
+ 35 37 42 43
c85 34 0 1.74227e-19 $X=3.59 $Y=1.95
c86 23 0 1.82144e-19 $X=3.505 $Y=1.465
c87 9 0 7.85372e-20 $X=2.455 $Y=0.69
r88 47 48 2.41806 $w=2.99e-07 $l=1.5e-08 $layer=POLY_cond $X=2.92 $Y=1.465
+ $X2=2.935 $Y2=1.465
r89 43 48 13.6699 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.025 $Y=1.465
+ $X2=2.935 $Y2=1.465
r90 35 37 21.8266 $w=3.28e-07 $l=6.25e-07 $layer=LI1_cond $X=3.675 $Y=2.115
+ $X2=4.3 $Y2=2.115
r91 34 35 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.59 $Y=1.95
+ $X2=3.675 $Y2=2.115
r92 33 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.59 $Y=1.63
+ $X2=3.59 $Y2=1.465
r93 33 34 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.59 $Y=1.63 $X2=3.59
+ $Y2=1.95
r94 32 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.59 $Y=1.3 $X2=3.59
+ $Y2=1.465
r95 31 41 9.62299 $w=3.74e-07 $l=4.00231e-07 $layer=LI1_cond $X=3.59 $Y=1.13
+ $X2=3.885 $Y2=0.882
r96 31 32 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.59 $Y=1.13
+ $X2=3.59 $Y2=1.3
r97 30 43 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=3.35 $Y=1.465
+ $X2=3.025 $Y2=1.465
r98 29 30 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.35
+ $Y=1.465 $X2=3.35 $Y2=1.465
r99 26 47 42.7191 $w=2.99e-07 $l=2.65e-07 $layer=POLY_cond $X=2.655 $Y=1.465
+ $X2=2.92 $Y2=1.465
r100 25 29 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.655 $Y=1.465
+ $X2=3.35 $Y2=1.465
r101 25 26 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.655
+ $Y=1.465 $X2=2.655 $Y2=1.465
r102 23 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.505 $Y=1.465
+ $X2=3.59 $Y2=1.465
r103 23 29 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.505 $Y=1.465
+ $X2=3.35 $Y2=1.465
r104 22 30 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.365 $Y=1.465
+ $X2=3.35 $Y2=1.465
r105 19 22 14.8326 $w=5.17e-07 $l=2.96606e-07 $layer=POLY_cond $X=3.455 $Y=1.72
+ $X2=3.365 $Y2=1.465
r106 19 21 144.6 $w=1.8e-07 $l=5.4e-07 $layer=POLY_cond $X=3.455 $Y=1.72
+ $X2=3.455 $Y2=2.26
r107 15 48 14.6425 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.935 $Y=1.63
+ $X2=2.935 $Y2=1.465
r108 15 17 244.887 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=2.935 $Y=1.63
+ $X2=2.935 $Y2=2.26
r109 11 47 18.89 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.92 $Y=1.3 $X2=2.92
+ $Y2=1.465
r110 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.92 $Y=1.3
+ $X2=2.92 $Y2=0.69
r111 7 26 32.2408 $w=2.99e-07 $l=2.70185e-07 $layer=POLY_cond $X=2.455 $Y=1.3
+ $X2=2.655 $Y2=1.465
r112 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.455 $Y=1.3
+ $X2=2.455 $Y2=0.69
r113 2 37 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=4.165
+ $Y=1.84 $X2=4.3 $Y2=2.115
r114 1 41 182 $w=1.7e-07 $l=4.04166e-07 $layer=licon1_NDIFF $count=1 $X=3.72
+ $Y=0.47 $X2=3.885 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2A_4%A2_N 3 7 9 12 13
c40 7 0 1.762e-19 $X=4.1 $Y=0.79
r41 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.01 $Y=1.515
+ $X2=4.01 $Y2=1.68
r42 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.01 $Y=1.515
+ $X2=4.01 $Y2=1.35
r43 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.01
+ $Y=1.515 $X2=4.01 $Y2=1.515
r44 9 13 4.93904 $w=3.48e-07 $l=1.5e-07 $layer=LI1_cond $X=4.02 $Y=1.665
+ $X2=4.02 $Y2=1.515
r45 7 14 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.1 $Y=0.79 $X2=4.1
+ $Y2=1.35
r46 3 15 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=4.075 $Y=2.26
+ $X2=4.075 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2A_4%A1_N 3 7 9 12 13
r39 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.58 $Y=1.515
+ $X2=4.58 $Y2=1.68
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.58 $Y=1.515
+ $X2=4.58 $Y2=1.35
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.58
+ $Y=1.515 $X2=4.58 $Y2=1.515
r42 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.58 $Y=1.665
+ $X2=4.58 $Y2=1.515
r43 7 15 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=4.525 $Y=2.26
+ $X2=4.525 $Y2=1.68
r44 3 14 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.49 $Y=0.79 $X2=4.49
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2A_4%A_313_392# 1 2 3 10 12 15 17 21 23 25 28 30
+ 32 33 35 37 40 42 47 50 51 52 54 55 56 58 62 64 68 69 76 77 79 88
c177 68 0 8.35716e-20 $X=1.7 $Y=2.115
c178 56 0 2.65681e-20 $X=4.37 $Y=1.035
c179 47 0 7.85372e-20 $X=4.2 $Y=0.34
r180 87 88 31.3483 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=6.205 $Y=1.385
+ $X2=6.285 $Y2=1.385
r181 86 87 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=6.195 $Y=1.385
+ $X2=6.205 $Y2=1.385
r182 83 84 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=5.695 $Y=1.385
+ $X2=5.705 $Y2=1.385
r183 75 77 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=1.985
+ $X2=3.25 $Y2=1.985
r184 75 76 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.165 $Y=1.985
+ $X2=2.995 $Y2=1.985
r185 69 72 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=2.67 $Y=0.34
+ $X2=2.67 $Y2=0.52
r186 65 86 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=5.9 $Y=1.385
+ $X2=6.195 $Y2=1.385
r187 65 84 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=5.9 $Y=1.385
+ $X2=5.705 $Y2=1.385
r188 64 65 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.9
+ $Y=1.385 $X2=5.9 $Y2=1.385
r189 61 64 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.22 $Y=1.385
+ $X2=5.9 $Y2=1.385
r190 61 62 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.22
+ $Y=1.385 $X2=5.22 $Y2=1.385
r191 59 79 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5 $Y=1.385 $X2=5
+ $Y2=1.035
r192 59 61 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=5.085 $Y=1.385
+ $X2=5.22 $Y2=1.385
r193 57 59 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5 $Y=1.55 $X2=5
+ $Y2=1.385
r194 57 58 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=5 $Y=1.55 $X2=5
+ $Y2=2.45
r195 55 79 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=1.035
+ $X2=5 $Y2=1.035
r196 55 56 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=4.915 $Y=1.035
+ $X2=4.37 $Y2=1.035
r197 54 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.285 $Y=0.95
+ $X2=4.37 $Y2=1.035
r198 53 54 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=4.285 $Y=0.425
+ $X2=4.285 $Y2=0.95
r199 51 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.915 $Y=2.535
+ $X2=5 $Y2=2.45
r200 51 52 103.08 $w=1.68e-07 $l=1.58e-06 $layer=LI1_cond $X=4.915 $Y=2.535
+ $X2=3.335 $Y2=2.535
r201 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.25 $Y=2.45
+ $X2=3.335 $Y2=2.535
r202 49 77 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.25 $Y=2.15
+ $X2=3.25 $Y2=1.985
r203 49 50 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.25 $Y=2.15 $X2=3.25
+ $Y2=2.45
r204 48 69 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=0.34
+ $X2=2.67 $Y2=0.34
r205 47 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.2 $Y=0.34
+ $X2=4.285 $Y2=0.425
r206 47 48 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=4.2 $Y=0.34
+ $X2=2.835 $Y2=0.34
r207 46 68 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=2.035
+ $X2=1.7 $Y2=2.035
r208 46 76 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=1.785 $Y=2.035
+ $X2=2.995 $Y2=2.035
r209 38 42 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=6.65 $Y=1.37
+ $X2=6.65 $Y2=1.295
r210 38 40 400.371 $w=1.8e-07 $l=1.03e-06 $layer=POLY_cond $X=6.65 $Y=1.37
+ $X2=6.65 $Y2=2.4
r211 35 42 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=6.635 $Y=1.22
+ $X2=6.65 $Y2=1.295
r212 35 37 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.635 $Y=1.22
+ $X2=6.635 $Y2=0.74
r213 33 42 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.56 $Y=1.295
+ $X2=6.65 $Y2=1.295
r214 33 88 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=6.56 $Y=1.295
+ $X2=6.285 $Y2=1.295
r215 30 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.205 $Y=1.22
+ $X2=6.205 $Y2=1.385
r216 30 32 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.205 $Y=1.22
+ $X2=6.205 $Y2=0.74
r217 26 86 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.195 $Y=1.55
+ $X2=6.195 $Y2=1.385
r218 26 28 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=6.195 $Y=1.55
+ $X2=6.195 $Y2=2.4
r219 23 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.705 $Y=1.22
+ $X2=5.705 $Y2=1.385
r220 23 25 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.705 $Y=1.22
+ $X2=5.705 $Y2=0.74
r221 19 83 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.695 $Y=1.55
+ $X2=5.695 $Y2=1.385
r222 19 21 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=5.695 $Y=1.55
+ $X2=5.695 $Y2=2.4
r223 18 62 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.235 $Y=1.385
+ $X2=5.145 $Y2=1.385
r224 17 83 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.605 $Y=1.385
+ $X2=5.695 $Y2=1.385
r225 17 18 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=5.605 $Y=1.385
+ $X2=5.235 $Y2=1.385
r226 13 62 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=5.145 $Y=1.55
+ $X2=5.145 $Y2=1.385
r227 13 15 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=5.145 $Y=1.55
+ $X2=5.145 $Y2=2.4
r228 10 62 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=5.13 $Y=1.22
+ $X2=5.145 $Y2=1.385
r229 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.13 $Y=1.22
+ $X2=5.13 $Y2=0.74
r230 3 75 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.025
+ $Y=1.84 $X2=3.165 $Y2=1.985
r231 2 68 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=1.565
+ $Y=1.96 $X2=1.7 $Y2=2.115
r232 1 72 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=2.53
+ $Y=0.37 $X2=2.67 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2A_4%A_41_392# 1 2 3 10 12 14 16 19 20 21 24
c48 16 0 5.55308e-20 $X=1.25 $Y=2.12
c49 10 0 4.76839e-20 $X=0.35 $Y=2.12
r50 22 24 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.15 $Y=2.905
+ $X2=2.15 $Y2=2.455
r51 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.985 $Y=2.99
+ $X2=2.15 $Y2=2.905
r52 20 21 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.985 $Y=2.99
+ $X2=1.415 $Y2=2.99
r53 17 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.25 $Y=2.905
+ $X2=1.415 $Y2=2.99
r54 17 19 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.25 $Y=2.905 $X2=1.25
+ $Y2=2.815
r55 16 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=2.12 $X2=1.25
+ $Y2=2.035
r56 16 19 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.25 $Y=2.12
+ $X2=1.25 $Y2=2.815
r57 15 27 5.07788 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=0.515 $Y=2.035
+ $X2=0.35 $Y2=2.03
r58 14 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.085 $Y=2.035
+ $X2=1.25 $Y2=2.035
r59 14 15 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.085 $Y=2.035
+ $X2=0.515 $Y2=2.035
r60 10 27 2.68829 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=0.35 $Y=2.12 $X2=0.35
+ $Y2=2.03
r61 10 12 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.35 $Y=2.12
+ $X2=0.35 $Y2=2.815
r62 3 24 300 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=2 $X=2.015
+ $Y=1.96 $X2=2.15 $Y2=2.455
r63 2 29 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=1.115
+ $Y=1.96 $X2=1.25 $Y2=2.115
r64 2 19 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.115
+ $Y=1.96 $X2=1.25 $Y2=2.815
r65 1 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.96 $X2=0.35 $Y2=2.105
r66 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.96 $X2=0.35 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2A_4%VPWR 1 2 3 4 5 6 23 27 29 33 37 41 45 47 52
+ 53 54 56 68 72 78 81 84 87 91
r97 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r98 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r99 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r100 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r101 76 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r102 76 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r103 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r104 73 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.085 $Y=3.33
+ $X2=5.92 $Y2=3.33
r105 73 75 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.085 $Y=3.33
+ $X2=6.48 $Y2=3.33
r106 72 90 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.755 $Y=3.33
+ $X2=6.977 $Y2=3.33
r107 72 75 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=3.33
+ $X2=6.48 $Y2=3.33
r108 71 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r109 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r110 68 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.755 $Y=3.33
+ $X2=5.92 $Y2=3.33
r111 68 70 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.755 $Y=3.33
+ $X2=5.52 $Y2=3.33
r112 67 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r113 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r114 64 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.93 $Y=3.33
+ $X2=3.765 $Y2=3.33
r115 64 66 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.93 $Y=3.33
+ $X2=4.56 $Y2=3.33
r116 63 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r117 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r118 60 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r119 60 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r120 59 62 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r121 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r122 57 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=0.8 $Y2=3.33
r123 57 59 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=3.33
+ $X2=1.2 $Y2=3.33
r124 56 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=3.33
+ $X2=2.71 $Y2=3.33
r125 56 62 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.545 $Y=3.33
+ $X2=2.16 $Y2=3.33
r126 54 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r127 54 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r128 54 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r129 52 66 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=4.67 $Y=3.33
+ $X2=4.56 $Y2=3.33
r130 52 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.67 $Y=3.33
+ $X2=4.835 $Y2=3.33
r131 51 70 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5 $Y=3.33 $X2=5.52
+ $Y2=3.33
r132 51 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5 $Y=3.33 $X2=4.835
+ $Y2=3.33
r133 47 50 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=6.92 $Y=1.985
+ $X2=6.92 $Y2=2.815
r134 45 90 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.92 $Y=3.245
+ $X2=6.977 $Y2=3.33
r135 45 50 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.92 $Y=3.245
+ $X2=6.92 $Y2=2.815
r136 41 44 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.92 $Y=2.145
+ $X2=5.92 $Y2=2.825
r137 39 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=3.245
+ $X2=5.92 $Y2=3.33
r138 39 44 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=5.92 $Y=3.245
+ $X2=5.92 $Y2=2.825
r139 35 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.835 $Y=3.245
+ $X2=4.835 $Y2=3.33
r140 35 37 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=4.835 $Y=3.245
+ $X2=4.835 $Y2=2.955
r141 31 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.765 $Y=3.245
+ $X2=3.765 $Y2=3.33
r142 31 33 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=3.765 $Y=3.245
+ $X2=3.765 $Y2=2.955
r143 30 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=3.33
+ $X2=2.71 $Y2=3.33
r144 29 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=3.765 $Y2=3.33
r145 29 30 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=2.875 $Y2=3.33
r146 25 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=3.245
+ $X2=2.71 $Y2=3.33
r147 25 27 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=2.71 $Y=3.245
+ $X2=2.71 $Y2=2.51
r148 21 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=3.245 $X2=0.8
+ $Y2=3.33
r149 21 23 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.8 $Y=3.245
+ $X2=0.8 $Y2=2.455
r150 6 50 400 $w=1.7e-07 $l=1.06119e-06 $layer=licon1_PDIFF $count=1 $X=6.74
+ $Y=1.84 $X2=6.92 $Y2=2.815
r151 6 47 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=6.74
+ $Y=1.84 $X2=6.92 $Y2=1.985
r152 5 44 400 $w=1.7e-07 $l=1.05033e-06 $layer=licon1_PDIFF $count=1 $X=5.785
+ $Y=1.84 $X2=5.92 $Y2=2.825
r153 5 41 400 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_PDIFF $count=1 $X=5.785
+ $Y=1.84 $X2=5.92 $Y2=2.145
r154 4 37 600 $w=1.7e-07 $l=1.22005e-06 $layer=licon1_PDIFF $count=1 $X=4.615
+ $Y=1.84 $X2=4.835 $Y2=2.955
r155 3 33 600 $w=1.7e-07 $l=1.22005e-06 $layer=licon1_PDIFF $count=1 $X=3.545
+ $Y=1.84 $X2=3.765 $Y2=2.955
r156 2 27 600 $w=1.7e-07 $l=7.38952e-07 $layer=licon1_PDIFF $count=1 $X=2.565
+ $Y=1.84 $X2=2.71 $Y2=2.51
r157 1 23 300 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=2 $X=0.665
+ $Y=1.96 $X2=0.8 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2A_4%X 1 2 3 4 13 15 19 23 24 27 30 33 37 38 39
+ 40 41
r67 40 45 4.07572 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=5.42 $Y=0.93
+ $X2=5.585 $Y2=0.93
r68 40 41 19.4475 $w=2.38e-07 $l=4.05e-07 $layer=LI1_cond $X=5.595 $Y=0.93 $X2=6
+ $Y2=0.93
r69 40 45 0.480185 $w=2.38e-07 $l=1e-08 $layer=LI1_cond $X=5.595 $Y=0.93
+ $X2=5.585 $Y2=0.93
r70 37 41 12.2447 $w=2.38e-07 $l=2.55e-07 $layer=LI1_cond $X=6.255 $Y=0.93 $X2=6
+ $Y2=0.93
r71 37 38 2.51069 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=6.255 $Y=0.93
+ $X2=6.42 $Y2=0.93
r72 33 35 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=6.42 $Y=1.985
+ $X2=6.42 $Y2=2.815
r73 31 39 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=1.89 $X2=6.42
+ $Y2=1.805
r74 31 33 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=6.42 $Y=1.89
+ $X2=6.42 $Y2=1.985
r75 30 39 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=1.72 $X2=6.42
+ $Y2=1.805
r76 29 38 3.93362 $w=3.3e-07 $l=1.2e-07 $layer=LI1_cond $X=6.42 $Y=1.05 $X2=6.42
+ $Y2=0.93
r77 29 30 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=6.42 $Y=1.05
+ $X2=6.42 $Y2=1.72
r78 25 38 3.93362 $w=3.3e-07 $l=1.2e-07 $layer=LI1_cond $X=6.42 $Y=0.81 $X2=6.42
+ $Y2=0.93
r79 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.42 $Y=0.81
+ $X2=6.42 $Y2=0.515
r80 23 39 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.255 $Y=1.805
+ $X2=6.42 $Y2=1.805
r81 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.255 $Y=1.805
+ $X2=5.585 $Y2=1.805
r82 19 21 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=5.42 $Y=1.985
+ $X2=5.42 $Y2=2.815
r83 17 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.42 $Y=1.89
+ $X2=5.585 $Y2=1.805
r84 17 19 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=5.42 $Y=1.89
+ $X2=5.42 $Y2=1.985
r85 13 40 2.96416 $w=3.3e-07 $l=1.2e-07 $layer=LI1_cond $X=5.42 $Y=0.81 $X2=5.42
+ $Y2=0.93
r86 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.42 $Y=0.81
+ $X2=5.42 $Y2=0.515
r87 4 35 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.285
+ $Y=1.84 $X2=6.42 $Y2=2.815
r88 4 33 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.285
+ $Y=1.84 $X2=6.42 $Y2=1.985
r89 3 21 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=5.235
+ $Y=1.84 $X2=5.42 $Y2=2.815
r90 3 19 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=5.235
+ $Y=1.84 $X2=5.42 $Y2=1.985
r91 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.28
+ $Y=0.37 $X2=6.42 $Y2=0.515
r92 1 15 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=5.205
+ $Y=0.37 $X2=5.42 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2A_4%A_27_74# 1 2 3 4 15 17 18 21 23 27 29
c53 21 0 1.72779e-19 $X=1.28 $Y=0.515
r54 29 31 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.17 $Y=0.81
+ $X2=3.17 $Y2=0.935
r55 24 27 6.67463 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=0.935
+ $X2=1.28 $Y2=0.935
r56 24 26 28.997 $w=3.08e-07 $l=7.8e-07 $layer=LI1_cond $X=1.445 $Y=0.935
+ $X2=2.225 $Y2=0.935
r57 23 31 1.09485 $w=3.1e-07 $l=1.65e-07 $layer=LI1_cond $X=3.005 $Y=0.935
+ $X2=3.17 $Y2=0.935
r58 23 26 28.997 $w=3.08e-07 $l=7.8e-07 $layer=LI1_cond $X=3.005 $Y=0.935
+ $X2=2.225 $Y2=0.935
r59 19 27 0.225187 $w=3.3e-07 $l=1.55e-07 $layer=LI1_cond $X=1.28 $Y=0.78
+ $X2=1.28 $Y2=0.935
r60 19 21 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=1.28 $Y=0.78
+ $X2=1.28 $Y2=0.515
r61 17 27 6.67463 $w=2.4e-07 $l=1.96914e-07 $layer=LI1_cond $X=1.115 $Y=1.005
+ $X2=1.28 $Y2=0.935
r62 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=1.005
+ $X2=0.445 $Y2=1.005
r63 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.92
+ $X2=0.445 $Y2=1.005
r64 13 15 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=0.28 $Y=0.92
+ $X2=0.28 $Y2=0.515
r65 4 29 182 $w=1.7e-07 $l=5.20192e-07 $layer=licon1_NDIFF $count=1 $X=2.995
+ $Y=0.37 $X2=3.17 $Y2=0.81
r66 3 26 182 $w=1.7e-07 $l=5.6723e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.37 $X2=2.225 $Y2=0.865
r67 2 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.14
+ $Y=0.37 $X2=1.28 $Y2=0.515
r68 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2A_4%VGND 1 2 3 4 5 18 20 24 28 32 34 36 38 40
+ 45 50 55 61 64 67 70 74
c86 28 0 1.762e-19 $X=4.81 $Y=0.64
r87 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r88 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r89 67 68 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r90 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r91 62 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r92 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r93 59 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r94 59 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r95 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r96 56 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.085 $Y=0 $X2=5.92
+ $Y2=0
r97 56 58 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.085 $Y=0 $X2=6.48
+ $Y2=0
r98 55 73 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.977
+ $Y2=0
r99 55 58 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=0 $X2=6.48
+ $Y2=0
r100 54 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r101 54 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r102 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r103 51 67 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=4.81
+ $Y2=0
r104 51 53 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=5.52
+ $Y2=0
r105 50 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.755 $Y=0 $X2=5.92
+ $Y2=0
r106 50 53 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.755 $Y=0
+ $X2=5.52 $Y2=0
r107 49 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r108 48 49 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r109 46 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=1.78
+ $Y2=0
r110 46 48 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.945 $Y=0
+ $X2=2.16 $Y2=0
r111 45 67 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=4.54 $Y=0 $X2=4.81
+ $Y2=0
r112 45 48 155.273 $w=1.68e-07 $l=2.38e-06 $layer=LI1_cond $X=4.54 $Y=0 $X2=2.16
+ $Y2=0
r113 43 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r114 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r115 40 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r116 40 42 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r117 38 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r118 38 49 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.16
+ $Y2=0
r119 34 73 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.977 $Y2=0
r120 34 36 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.92 $Y=0.085
+ $X2=6.92 $Y2=0.515
r121 30 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0
r122 30 32 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=5.92 $Y=0.085
+ $X2=5.92 $Y2=0.535
r123 26 67 2.26835 $w=5.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.81 $Y=0.085
+ $X2=4.81 $Y2=0
r124 26 28 12.293 $w=5.38e-07 $l=5.55e-07 $layer=LI1_cond $X=4.81 $Y=0.085
+ $X2=4.81 $Y2=0.64
r125 22 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0
r126 22 24 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0.52
r127 21 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r128 20 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.615 $Y=0 $X2=1.78
+ $Y2=0
r129 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=0
+ $X2=0.945 $Y2=0
r130 16 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r131 16 18 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.55
r132 5 36 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=6.71
+ $Y=0.37 $X2=6.92 $Y2=0.515
r133 4 32 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=5.78
+ $Y=0.37 $X2=5.92 $Y2=0.535
r134 3 28 182 $w=1.7e-07 $l=3.18865e-07 $layer=licon1_NDIFF $count=1 $X=4.565
+ $Y=0.47 $X2=4.81 $Y2=0.64
r135 2 24 182 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.37 $X2=1.78 $Y2=0.52
r136 1 18 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.55
.ends


* File: sky130_fd_sc_ms__nand4bb_4.pex.spice
* Created: Wed Sep  2 12:15:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NAND4BB_4%A_N 1 3 6 9 10 12 18 21
c47 21 0 1.99278e-19 $X=0.605 $Y=1.615
r48 21 23 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.595 $Y=1.615
+ $X2=0.595 $Y2=1.45
r49 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.605
+ $Y=1.615 $X2=0.605 $Y2=1.615
r50 18 22 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.72 $Y=1.615
+ $X2=0.605 $Y2=1.615
r51 10 12 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=0.955 $Y=2.045
+ $X2=0.955 $Y2=2.54
r52 9 10 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=0.595 $Y=1.97
+ $X2=0.955 $Y2=1.97
r53 8 21 1.64869 $w=3.5e-07 $l=1e-08 $layer=POLY_cond $X=0.595 $Y=1.625
+ $X2=0.595 $Y2=1.615
r54 8 9 44.5147 $w=3.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.595 $Y=1.625
+ $X2=0.595 $Y2=1.895
r55 6 23 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.495 $Y=0.94
+ $X2=0.495 $Y2=1.45
r56 1 9 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.97 $X2=0.595
+ $Y2=1.97
r57 1 3 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=0.505 $Y=2.045
+ $X2=0.505 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4BB_4%B_N 3 5 6 9 11 13 14 18
c58 14 0 9.63788e-20 $X=1.68 $Y=1.665
r59 14 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=1.715 $X2=1.63 $Y2=1.715
r60 11 18 26.8441 $w=4.04e-07 $l=3.7081e-07 $layer=POLY_cond $X=1.855 $Y=2.055
+ $X2=1.63 $Y2=1.78
r61 11 13 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=1.855 $Y=2.055
+ $X2=1.855 $Y2=2.54
r62 7 18 26.8441 $w=4.04e-07 $l=2.25e-07 $layer=POLY_cond $X=1.405 $Y=1.78
+ $X2=1.63 $Y2=1.78
r63 7 9 223.508 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.405 $Y=1.965
+ $X2=1.405 $Y2=2.54
r64 5 7 30.7166 $w=4.04e-07 $l=2.40832e-07 $layer=POLY_cond $X=1.315 $Y=1.58
+ $X2=1.405 $Y2=1.78
r65 5 6 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.315 $Y=1.58
+ $X2=1.16 $Y2=1.58
r66 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.085 $Y=1.505
+ $X2=1.16 $Y2=1.58
r67 1 3 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=1.085 $Y=1.505
+ $X2=1.085 $Y2=0.94
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4BB_4%A_27_114# 1 2 7 9 10 12 13 15 16 18 19 21
+ 22 24 27 29 30 31 33 34 35 37 38 39 40 44 47 49 50 55 60 61
c158 27 0 1.79504e-19 $X=3.635 $Y=0.74
c159 19 0 7.06753e-20 $X=3.205 $Y=1.22
c160 13 0 7.06753e-20 $X=2.765 $Y=1.22
c161 10 0 9.63788e-20 $X=2.575 $Y=1.725
r162 68 69 32.4716 $w=4.75e-07 $l=3.2e-07 $layer=POLY_cond $X=3.205 $Y=1.472
+ $X2=3.525 $Y2=1.472
r163 67 68 13.1916 $w=4.75e-07 $l=1.3e-07 $layer=POLY_cond $X=3.075 $Y=1.472
+ $X2=3.205 $Y2=1.472
r164 62 63 35.0084 $w=4.75e-07 $l=3.45e-07 $layer=POLY_cond $X=2.23 $Y=1.472
+ $X2=2.575 $Y2=1.472
r165 56 67 7.61053 $w=4.75e-07 $l=7.5e-08 $layer=POLY_cond $X=3 $Y=1.472
+ $X2=3.075 $Y2=1.472
r166 56 65 23.8463 $w=4.75e-07 $l=2.35e-07 $layer=POLY_cond $X=3 $Y=1.472
+ $X2=2.765 $Y2=1.472
r167 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3
+ $Y=1.385 $X2=3 $Y2=1.385
r168 53 65 10.6547 $w=4.75e-07 $l=1.05e-07 $layer=POLY_cond $X=2.66 $Y=1.472
+ $X2=2.765 $Y2=1.472
r169 53 63 8.62526 $w=4.75e-07 $l=8.5e-08 $layer=POLY_cond $X=2.66 $Y=1.472
+ $X2=2.575 $Y2=1.472
r170 52 55 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=2.66 $Y=1.38 $X2=3
+ $Y2=1.38
r171 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.66
+ $Y=1.385 $X2=2.66 $Y2=1.385
r172 50 61 14.4036 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=2.495 $Y=1.38
+ $X2=2.155 $Y2=1.38
r173 50 52 5.59274 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.495 $Y=1.38
+ $X2=2.66 $Y2=1.38
r174 49 61 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.76 $Y=1.295
+ $X2=2.155 $Y2=1.295
r175 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.675 $Y=1.21
+ $X2=1.76 $Y2=1.295
r176 46 47 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.675 $Y=0.83
+ $X2=1.675 $Y2=1.21
r177 42 44 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.73 $Y=2.12
+ $X2=0.73 $Y2=2.265
r178 41 59 4.8908 $w=1.7e-07 $l=1.98605e-07 $layer=LI1_cond $X=0.445 $Y=0.745
+ $X2=0.272 $Y2=0.69
r179 40 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.59 $Y=0.745
+ $X2=1.675 $Y2=0.83
r180 40 41 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=1.59 $Y=0.745
+ $X2=0.445 $Y2=0.745
r181 38 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.645 $Y=2.035
+ $X2=0.73 $Y2=2.12
r182 38 39 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.645 $Y=2.035
+ $X2=0.27 $Y2=2.035
r183 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.185 $Y=1.95
+ $X2=0.27 $Y2=2.035
r184 37 60 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.185 $Y=1.95
+ $X2=0.185 $Y2=1.28
r185 35 60 8.71323 $w=3.43e-07 $l=1.72e-07 $layer=LI1_cond $X=0.272 $Y=1.108
+ $X2=0.272 $Y2=1.28
r186 34 59 3.00312 $w=3.45e-07 $l=1.4e-07 $layer=LI1_cond $X=0.272 $Y=0.83
+ $X2=0.272 $Y2=0.69
r187 34 35 9.28635 $w=3.43e-07 $l=2.78e-07 $layer=LI1_cond $X=0.272 $Y=0.83
+ $X2=0.272 $Y2=1.108
r188 31 33 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.975 $Y=1.725
+ $X2=3.975 $Y2=2.4
r189 29 31 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.885 $Y=1.65
+ $X2=3.975 $Y2=1.725
r190 29 30 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=3.885 $Y=1.65
+ $X2=3.71 $Y2=1.65
r191 25 30 32.1576 $w=4.75e-07 $l=2.12212e-07 $layer=POLY_cond $X=3.635 $Y=1.472
+ $X2=3.71 $Y2=1.65
r192 25 69 11.1621 $w=4.75e-07 $l=1.1e-07 $layer=POLY_cond $X=3.635 $Y=1.472
+ $X2=3.525 $Y2=1.472
r193 25 27 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=3.635 $Y=1.325
+ $X2=3.635 $Y2=0.74
r194 22 69 25.6061 $w=1.8e-07 $l=2.53e-07 $layer=POLY_cond $X=3.525 $Y=1.725
+ $X2=3.525 $Y2=1.472
r195 22 24 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.525 $Y=1.725
+ $X2=3.525 $Y2=2.4
r196 19 68 30.117 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=3.205 $Y=1.22
+ $X2=3.205 $Y2=1.472
r197 19 21 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.205 $Y=1.22
+ $X2=3.205 $Y2=0.74
r198 16 67 25.6061 $w=1.8e-07 $l=2.53e-07 $layer=POLY_cond $X=3.075 $Y=1.725
+ $X2=3.075 $Y2=1.472
r199 16 18 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.075 $Y=1.725
+ $X2=3.075 $Y2=2.4
r200 13 65 30.117 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=2.765 $Y=1.22
+ $X2=2.765 $Y2=1.472
r201 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.765 $Y=1.22
+ $X2=2.765 $Y2=0.74
r202 10 63 25.6061 $w=1.8e-07 $l=2.53e-07 $layer=POLY_cond $X=2.575 $Y=1.725
+ $X2=2.575 $Y2=1.472
r203 10 12 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=2.575 $Y=1.725
+ $X2=2.575 $Y2=2.4
r204 7 62 30.117 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=2.23 $Y=1.22
+ $X2=2.23 $Y2=1.472
r205 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.23 $Y=1.22 $X2=2.23
+ $Y2=0.74
r206 2 44 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=2.12 $X2=0.73 $Y2=2.265
r207 1 59 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.57 $X2=0.28 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4BB_4%A_232_114# 1 2 7 9 10 11 14 16 18 21 23 25
+ 28 30 32 35 38 39 40 43 46 47 48 49 54 60 63 76
c175 38 0 1.99278e-19 $X=1.21 $Y=2.05
c176 21 0 6.32537e-21 $X=4.875 $Y=2.4
r177 75 76 15.9151 $w=4.24e-07 $l=1.4e-07 $layer=POLY_cond $X=5.375 $Y=1.432
+ $X2=5.515 $Y2=1.432
r178 72 73 5.68396 $w=4.24e-07 $l=5e-08 $layer=POLY_cond $X=4.875 $Y=1.432
+ $X2=4.925 $Y2=1.432
r179 69 70 7.95755 $w=4.24e-07 $l=7e-08 $layer=POLY_cond $X=4.425 $Y=1.432
+ $X2=4.495 $Y2=1.432
r180 57 60 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=1.21 $Y=1.165
+ $X2=1.315 $Y2=1.165
r181 55 75 22.1675 $w=4.24e-07 $l=1.95e-07 $layer=POLY_cond $X=5.18 $Y=1.432
+ $X2=5.375 $Y2=1.432
r182 55 73 28.9882 $w=4.24e-07 $l=2.55e-07 $layer=POLY_cond $X=5.18 $Y=1.432
+ $X2=4.925 $Y2=1.432
r183 54 55 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.18
+ $Y=1.515 $X2=5.18 $Y2=1.515
r184 52 72 42.6297 $w=4.24e-07 $l=3.75e-07 $layer=POLY_cond $X=4.5 $Y=1.432
+ $X2=4.875 $Y2=1.432
r185 52 70 0.568396 $w=4.24e-07 $l=5e-09 $layer=POLY_cond $X=4.5 $Y=1.432
+ $X2=4.495 $Y2=1.432
r186 51 54 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=4.5 $Y=1.555
+ $X2=5.18 $Y2=1.555
r187 51 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.5
+ $Y=1.515 $X2=4.5 $Y2=1.515
r188 49 67 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.23 $Y=1.555
+ $X2=4.23 $Y2=1.805
r189 49 51 8.52808 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=4.315 $Y=1.555
+ $X2=4.5 $Y2=1.555
r190 47 67 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.145 $Y=1.805
+ $X2=4.23 $Y2=1.805
r191 47 48 131.134 $w=1.68e-07 $l=2.01e-06 $layer=LI1_cond $X=4.145 $Y=1.805
+ $X2=2.135 $Y2=1.805
r192 46 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=2.05
+ $X2=2.05 $Y2=2.135
r193 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.05 $Y=1.89
+ $X2=2.135 $Y2=1.805
r194 45 46 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.05 $Y=1.89
+ $X2=2.05 $Y2=2.05
r195 41 63 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.655 $Y=2.135
+ $X2=2.05 $Y2=2.135
r196 41 43 1.85214 $w=2.78e-07 $l=4.5e-08 $layer=LI1_cond $X=1.655 $Y=2.22
+ $X2=1.655 $Y2=2.265
r197 39 41 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.515 $Y=2.135
+ $X2=1.655 $Y2=2.135
r198 39 40 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.515 $Y=2.135
+ $X2=1.295 $Y2=2.135
r199 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.21 $Y=2.05
+ $X2=1.295 $Y2=2.135
r200 37 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.21 $Y=1.33
+ $X2=1.21 $Y2=1.165
r201 37 38 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.21 $Y=1.33
+ $X2=1.21 $Y2=2.05
r202 33 76 35.2406 $w=4.24e-07 $l=4.15909e-07 $layer=POLY_cond $X=5.825 $Y=1.68
+ $X2=5.515 $Y2=1.432
r203 33 35 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.825 $Y=1.68
+ $X2=5.825 $Y2=2.4
r204 30 76 27.2926 $w=1.5e-07 $l=2.47e-07 $layer=POLY_cond $X=5.515 $Y=1.185
+ $X2=5.515 $Y2=1.432
r205 30 32 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.515 $Y=1.185
+ $X2=5.515 $Y2=0.74
r206 26 75 22.8561 $w=1.8e-07 $l=2.48e-07 $layer=POLY_cond $X=5.375 $Y=1.68
+ $X2=5.375 $Y2=1.432
r207 26 28 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.375 $Y=1.68
+ $X2=5.375 $Y2=2.4
r208 23 73 27.2926 $w=1.5e-07 $l=2.47e-07 $layer=POLY_cond $X=4.925 $Y=1.185
+ $X2=4.925 $Y2=1.432
r209 23 25 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.925 $Y=1.185
+ $X2=4.925 $Y2=0.74
r210 19 72 22.8561 $w=1.8e-07 $l=2.48e-07 $layer=POLY_cond $X=4.875 $Y=1.68
+ $X2=4.875 $Y2=1.432
r211 19 21 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.875 $Y=1.68
+ $X2=4.875 $Y2=2.4
r212 16 70 27.2926 $w=1.5e-07 $l=2.47e-07 $layer=POLY_cond $X=4.495 $Y=1.185
+ $X2=4.495 $Y2=1.432
r213 16 18 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.495 $Y=1.185
+ $X2=4.495 $Y2=0.74
r214 12 69 22.8561 $w=1.8e-07 $l=2.48e-07 $layer=POLY_cond $X=4.425 $Y=1.68
+ $X2=4.425 $Y2=1.432
r215 12 14 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.425 $Y=1.68
+ $X2=4.425 $Y2=2.4
r216 10 69 31.5592 $w=4.24e-07 $l=2.12283e-07 $layer=POLY_cond $X=4.335 $Y=1.26
+ $X2=4.425 $Y2=1.432
r217 10 11 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=4.335 $Y=1.26
+ $X2=4.14 $Y2=1.26
r218 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.065 $Y=1.185
+ $X2=4.14 $Y2=1.26
r219 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.065 $Y=1.185
+ $X2=4.065 $Y2=0.74
r220 2 43 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=2.12 $X2=1.63 $Y2=2.265
r221 1 60 182 $w=1.7e-07 $l=6.68019e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.57 $X2=1.315 $Y2=1.165
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4BB_4%C 3 7 11 15 19 23 27 31 40 43 53 56 58
c98 58 0 1.90128e-19 $X=7.075 $Y=1.55
c99 11 0 1.16661e-20 $X=6.725 $Y=2.4
r100 53 54 10.4136 $w=3.24e-07 $l=7e-08 $layer=POLY_cond $X=7.725 $Y=1.485
+ $X2=7.795 $Y2=1.485
r101 50 51 13.3889 $w=3.24e-07 $l=9e-08 $layer=POLY_cond $X=7.275 $Y=1.485
+ $X2=7.365 $Y2=1.485
r102 49 50 50.5802 $w=3.24e-07 $l=3.4e-07 $layer=POLY_cond $X=6.935 $Y=1.485
+ $X2=7.275 $Y2=1.485
r103 48 49 31.2407 $w=3.24e-07 $l=2.1e-07 $layer=POLY_cond $X=6.725 $Y=1.485
+ $X2=6.935 $Y2=1.485
r104 47 48 32.7284 $w=3.24e-07 $l=2.2e-07 $layer=POLY_cond $X=6.505 $Y=1.485
+ $X2=6.725 $Y2=1.485
r105 43 58 3.96409 $w=4.58e-07 $l=1.15e-07 $layer=LI1_cond $X=6.96 $Y=1.55
+ $X2=7.075 $Y2=1.55
r106 43 56 3.96409 $w=4.58e-07 $l=1.15e-07 $layer=LI1_cond $X=6.96 $Y=1.55
+ $X2=6.845 $Y2=1.55
r107 41 53 41.6543 $w=3.24e-07 $l=2.8e-07 $layer=POLY_cond $X=7.445 $Y=1.485
+ $X2=7.725 $Y2=1.485
r108 41 51 11.9012 $w=3.24e-07 $l=8e-08 $layer=POLY_cond $X=7.445 $Y=1.485
+ $X2=7.365 $Y2=1.485
r109 40 58 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=7.445 $Y=1.485
+ $X2=7.075 $Y2=1.485
r110 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.445
+ $Y=1.485 $X2=7.445 $Y2=1.485
r111 36 47 11.9012 $w=3.24e-07 $l=8e-08 $layer=POLY_cond $X=6.425 $Y=1.485
+ $X2=6.505 $Y2=1.485
r112 36 45 22.3148 $w=3.24e-07 $l=1.5e-07 $layer=POLY_cond $X=6.425 $Y=1.485
+ $X2=6.275 $Y2=1.485
r113 35 56 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=6.425 $Y=1.485
+ $X2=6.845 $Y2=1.485
r114 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.425
+ $Y=1.485 $X2=6.425 $Y2=1.485
r115 29 54 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.795 $Y=1.32
+ $X2=7.795 $Y2=1.485
r116 29 31 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.795 $Y=1.32
+ $X2=7.795 $Y2=0.74
r117 25 53 16.5046 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.725 $Y=1.65
+ $X2=7.725 $Y2=1.485
r118 25 27 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=7.725 $Y=1.65
+ $X2=7.725 $Y2=2.4
r119 21 51 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.365 $Y=1.32
+ $X2=7.365 $Y2=1.485
r120 21 23 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.365 $Y=1.32
+ $X2=7.365 $Y2=0.74
r121 17 50 16.5046 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.275 $Y=1.65
+ $X2=7.275 $Y2=1.485
r122 17 19 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=7.275 $Y=1.65
+ $X2=7.275 $Y2=2.4
r123 13 49 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.935 $Y=1.32
+ $X2=6.935 $Y2=1.485
r124 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.935 $Y=1.32
+ $X2=6.935 $Y2=0.74
r125 9 48 16.5046 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.725 $Y=1.65
+ $X2=6.725 $Y2=1.485
r126 9 11 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=6.725 $Y=1.65
+ $X2=6.725 $Y2=2.4
r127 5 47 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.505 $Y=1.32
+ $X2=6.505 $Y2=1.485
r128 5 7 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.505 $Y=1.32
+ $X2=6.505 $Y2=0.74
r129 1 45 16.5046 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.275 $Y=1.65
+ $X2=6.275 $Y2=1.485
r130 1 3 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=6.275 $Y=1.65
+ $X2=6.275 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4BB_4%D 3 7 11 15 19 23 27 31 33 34 35 36 50
r89 52 53 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=9.765
+ $Y=1.465 $X2=9.765 $Y2=1.465
r90 50 52 26.4512 $w=3.28e-07 $l=1.8e-07 $layer=POLY_cond $X=9.585 $Y=1.465
+ $X2=9.765 $Y2=1.465
r91 49 50 1.46951 $w=3.28e-07 $l=1e-08 $layer=POLY_cond $X=9.575 $Y=1.465
+ $X2=9.585 $Y2=1.465
r92 48 49 66.1281 $w=3.28e-07 $l=4.5e-07 $layer=POLY_cond $X=9.125 $Y=1.465
+ $X2=9.575 $Y2=1.465
r93 47 48 5.87805 $w=3.28e-07 $l=4e-08 $layer=POLY_cond $X=9.085 $Y=1.465
+ $X2=9.125 $Y2=1.465
r94 46 47 60.25 $w=3.28e-07 $l=4.1e-07 $layer=POLY_cond $X=8.675 $Y=1.465
+ $X2=9.085 $Y2=1.465
r95 45 46 2.93902 $w=3.28e-07 $l=2e-08 $layer=POLY_cond $X=8.655 $Y=1.465
+ $X2=8.675 $Y2=1.465
r96 43 45 36.7378 $w=3.28e-07 $l=2.5e-07 $layer=POLY_cond $X=8.405 $Y=1.465
+ $X2=8.655 $Y2=1.465
r97 43 44 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=8.405
+ $Y=1.465 $X2=8.405 $Y2=1.465
r98 41 43 26.4512 $w=3.28e-07 $l=1.8e-07 $layer=POLY_cond $X=8.225 $Y=1.465
+ $X2=8.405 $Y2=1.465
r99 36 53 1.86887 $w=4.78e-07 $l=7.5e-08 $layer=LI1_cond $X=9.84 $Y=1.54
+ $X2=9.765 $Y2=1.54
r100 35 53 10.0919 $w=4.78e-07 $l=4.05e-07 $layer=LI1_cond $X=9.36 $Y=1.54
+ $X2=9.765 $Y2=1.54
r101 34 35 11.9608 $w=4.78e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.54
+ $X2=9.36 $Y2=1.54
r102 34 44 11.8362 $w=4.78e-07 $l=4.75e-07 $layer=LI1_cond $X=8.88 $Y=1.54
+ $X2=8.405 $Y2=1.54
r103 33 44 0.124591 $w=4.78e-07 $l=5e-09 $layer=LI1_cond $X=8.4 $Y=1.54
+ $X2=8.405 $Y2=1.54
r104 29 50 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.585 $Y=1.3
+ $X2=9.585 $Y2=1.465
r105 29 31 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=9.585 $Y=1.3
+ $X2=9.585 $Y2=0.74
r106 25 49 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.575 $Y=1.63
+ $X2=9.575 $Y2=1.465
r107 25 27 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=9.575 $Y=1.63
+ $X2=9.575 $Y2=2.4
r108 21 48 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.125 $Y=1.63
+ $X2=9.125 $Y2=1.465
r109 21 23 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=9.125 $Y=1.63
+ $X2=9.125 $Y2=2.4
r110 17 47 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.085 $Y=1.3
+ $X2=9.085 $Y2=1.465
r111 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=9.085 $Y=1.3
+ $X2=9.085 $Y2=0.74
r112 13 46 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.675 $Y=1.63
+ $X2=8.675 $Y2=1.465
r113 13 15 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=8.675 $Y=1.63
+ $X2=8.675 $Y2=2.4
r114 9 45 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.655 $Y=1.3
+ $X2=8.655 $Y2=1.465
r115 9 11 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.655 $Y=1.3
+ $X2=8.655 $Y2=0.74
r116 5 41 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.225 $Y=1.3
+ $X2=8.225 $Y2=1.465
r117 5 7 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.225 $Y=1.3
+ $X2=8.225 $Y2=0.74
r118 1 41 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.225 $Y=1.63
+ $X2=8.225 $Y2=1.465
r119 1 3 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=8.225 $Y=1.63
+ $X2=8.225 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4BB_4%VPWR 1 2 3 4 5 6 7 8 9 10 11 34 36 40 44
+ 48 50 54 56 60 64 68 70 74 76 80 82 84 88 89 90 92 97 106 111 116 125 128 131
+ 134 137 140 143 146 150
r173 149 150 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r174 146 147 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r175 144 147 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r176 143 144 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r177 141 144 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r178 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r179 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r180 131 132 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r181 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r182 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r183 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r184 120 150 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r185 120 147 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r186 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r187 117 146 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.985 $Y=3.33
+ $X2=8.9 $Y2=3.33
r188 117 119 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.985 $Y=3.33
+ $X2=9.36 $Y2=3.33
r189 116 149 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=9.715 $Y=3.33
+ $X2=9.897 $Y2=3.33
r190 116 119 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=9.715 $Y=3.33
+ $X2=9.36 $Y2=3.33
r191 115 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r192 115 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r193 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r194 112 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.135 $Y=3.33
+ $X2=6.01 $Y2=3.33
r195 112 114 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.135 $Y=3.33
+ $X2=6.48 $Y2=3.33
r196 111 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.835 $Y=3.33
+ $X2=7 $Y2=3.33
r197 111 114 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.835 $Y=3.33
+ $X2=6.48 $Y2=3.33
r198 110 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r199 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r200 107 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.15 $Y2=3.33
r201 107 109 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.52 $Y2=3.33
r202 106 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.885 $Y=3.33
+ $X2=6.01 $Y2=3.33
r203 106 109 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.885 $Y=3.33
+ $X2=5.52 $Y2=3.33
r204 105 132 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r205 105 129 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r206 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r207 102 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=2.17 $Y2=3.33
r208 102 104 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=3.12 $Y2=3.33
r209 101 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r210 101 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r211 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r212 98 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.18 $Y2=3.33
r213 98 100 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r214 97 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=3.33
+ $X2=2.17 $Y2=3.33
r215 97 100 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.005 $Y=3.33
+ $X2=1.68 $Y2=3.33
r216 96 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r217 96 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r218 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r219 93 122 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r220 93 95 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r221 92 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.18 $Y2=3.33
r222 92 95 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r223 90 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r224 90 132 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.08 $Y2=3.33
r225 90 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r226 88 104 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.135 $Y=3.33
+ $X2=3.12 $Y2=3.33
r227 88 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=3.33
+ $X2=3.3 $Y2=3.33
r228 84 87 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=9.84 $Y=2.115
+ $X2=9.84 $Y2=2.815
r229 82 149 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.84 $Y=3.245
+ $X2=9.897 $Y2=3.33
r230 82 87 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.84 $Y=3.245
+ $X2=9.84 $Y2=2.815
r231 78 146 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.9 $Y=3.245
+ $X2=8.9 $Y2=3.33
r232 78 80 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=8.9 $Y=3.245
+ $X2=8.9 $Y2=2.455
r233 77 143 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.115 $Y=3.33
+ $X2=7.99 $Y2=3.33
r234 76 146 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.815 $Y=3.33
+ $X2=8.9 $Y2=3.33
r235 76 77 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=8.815 $Y=3.33
+ $X2=8.115 $Y2=3.33
r236 72 143 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.99 $Y=3.245
+ $X2=7.99 $Y2=3.33
r237 72 74 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=7.99 $Y=3.245
+ $X2=7.99 $Y2=2.455
r238 71 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.165 $Y=3.33
+ $X2=7 $Y2=3.33
r239 70 143 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.865 $Y=3.33
+ $X2=7.99 $Y2=3.33
r240 70 71 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=7.865 $Y=3.33
+ $X2=7.165 $Y2=3.33
r241 66 140 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7 $Y=3.245 $X2=7
+ $Y2=3.33
r242 66 68 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=7 $Y=3.245 $X2=7
+ $Y2=2.455
r243 62 137 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.01 $Y=3.245
+ $X2=6.01 $Y2=3.33
r244 62 64 42.4099 $w=2.48e-07 $l=9.2e-07 $layer=LI1_cond $X=6.01 $Y=3.245
+ $X2=6.01 $Y2=2.325
r245 58 134 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.15 $Y=3.245
+ $X2=5.15 $Y2=3.33
r246 58 60 31.081 $w=3.28e-07 $l=8.9e-07 $layer=LI1_cond $X=5.15 $Y=3.245
+ $X2=5.15 $Y2=2.355
r247 57 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.365 $Y=3.33
+ $X2=4.2 $Y2=3.33
r248 56 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.985 $Y=3.33
+ $X2=5.15 $Y2=3.33
r249 56 57 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.985 $Y=3.33
+ $X2=4.365 $Y2=3.33
r250 52 131 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.2 $Y=3.245
+ $X2=4.2 $Y2=3.33
r251 52 54 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=4.2 $Y=3.245
+ $X2=4.2 $Y2=2.495
r252 51 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=3.33
+ $X2=3.3 $Y2=3.33
r253 50 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.035 $Y=3.33
+ $X2=4.2 $Y2=3.33
r254 50 51 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.035 $Y=3.33
+ $X2=3.465 $Y2=3.33
r255 46 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=3.245 $X2=3.3
+ $Y2=3.33
r256 46 48 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=3.3 $Y=3.245
+ $X2=3.3 $Y2=2.495
r257 42 128 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=3.33
r258 42 44 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=2.495
r259 38 125 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r260 38 40 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.495
r261 34 122 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r262 34 36 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.455
r263 11 87 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.665
+ $Y=1.84 $X2=9.8 $Y2=2.815
r264 11 84 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=9.665
+ $Y=1.84 $X2=9.8 $Y2=2.115
r265 10 80 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=8.765
+ $Y=1.84 $X2=8.9 $Y2=2.455
r266 9 74 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=7.815
+ $Y=1.84 $X2=7.95 $Y2=2.455
r267 8 68 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=6.815
+ $Y=1.84 $X2=7 $Y2=2.455
r268 7 64 300 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=2 $X=5.915
+ $Y=1.84 $X2=6.05 $Y2=2.325
r269 6 60 300 $w=1.7e-07 $l=6.00417e-07 $layer=licon1_PDIFF $count=2 $X=4.965
+ $Y=1.84 $X2=5.15 $Y2=2.355
r270 5 54 300 $w=1.7e-07 $l=7.1934e-07 $layer=licon1_PDIFF $count=2 $X=4.065
+ $Y=1.84 $X2=4.2 $Y2=2.495
r271 4 48 300 $w=1.7e-07 $l=7.1934e-07 $layer=licon1_PDIFF $count=2 $X=3.165
+ $Y=1.84 $X2=3.3 $Y2=2.495
r272 3 44 300 $w=1.7e-07 $l=4.74342e-07 $layer=licon1_PDIFF $count=2 $X=1.945
+ $Y=2.12 $X2=2.17 $Y2=2.495
r273 2 40 300 $w=1.7e-07 $l=4.37321e-07 $layer=licon1_PDIFF $count=2 $X=1.045
+ $Y=2.12 $X2=1.18 $Y2=2.495
r274 1 36 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4BB_4%Y 1 2 3 4 5 6 7 8 9 10 31 33 35 38 42 44
+ 48 50 53 56 58 62 64 68 70 74 76 78 80 83 87 90 94 95 102 103 109 111 114 115
c199 58 0 1.16661e-20 $X=6.335 $Y=1.905
c200 44 0 6.32537e-21 $X=4.485 $Y=2.145
c201 38 0 2.42988e-20 $X=5.515 $Y=1.175
r202 115 121 7.59565 $w=4.38e-07 $l=2.9e-07 $layer=LI1_cond $X=2.745 $Y=2.775
+ $X2=2.745 $Y2=2.485
r203 114 121 2.09535 $w=4.38e-07 $l=8e-08 $layer=LI1_cond $X=2.745 $Y=2.405
+ $X2=2.745 $Y2=2.485
r204 106 107 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=6.5 $Y=1.985
+ $X2=6.5 $Y2=2.035
r205 103 106 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=6.5 $Y=1.905 $X2=6.5
+ $Y2=1.985
r206 99 100 3.26614 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.65 $Y=2.145
+ $X2=4.65 $Y2=2.23
r207 98 99 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=4.65 $Y=2.015
+ $X2=4.65 $Y2=2.145
r208 95 98 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.65 $Y=1.935 $X2=4.65
+ $Y2=2.015
r209 90 91 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.42 $Y=0.955
+ $X2=3.42 $Y2=1.175
r210 87 114 4.58358 $w=4.38e-07 $l=1.75e-07 $layer=LI1_cond $X=2.745 $Y=2.23
+ $X2=2.745 $Y2=2.405
r211 87 89 2.42973 $w=4.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.745 $Y=2.23
+ $X2=2.745 $Y2=2.145
r212 83 85 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=2.485 $Y=0.815
+ $X2=2.485 $Y2=0.955
r213 78 113 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.35 $Y=2.12
+ $X2=9.35 $Y2=2.035
r214 78 80 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=9.35 $Y=2.12
+ $X2=9.35 $Y2=2.815
r215 77 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.615 $Y=2.035
+ $X2=8.45 $Y2=2.035
r216 76 113 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.185 $Y=2.035
+ $X2=9.35 $Y2=2.035
r217 76 77 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=9.185 $Y=2.035
+ $X2=8.615 $Y2=2.035
r218 72 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.45 $Y=2.12
+ $X2=8.45 $Y2=2.035
r219 72 74 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=8.45 $Y=2.12
+ $X2=8.45 $Y2=2.815
r220 71 109 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=7.665 $Y=2.035
+ $X2=7.5 $Y2=1.97
r221 70 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.285 $Y=2.035
+ $X2=8.45 $Y2=2.035
r222 70 71 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=8.285 $Y=2.035
+ $X2=7.665 $Y2=2.035
r223 66 109 0.89609 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=7.5 $Y=2.12 $X2=7.5
+ $Y2=1.97
r224 66 68 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=7.5 $Y=2.12
+ $X2=7.5 $Y2=2.815
r225 65 107 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.665 $Y=2.035
+ $X2=6.5 $Y2=2.035
r226 64 109 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=7.335 $Y=2.035
+ $X2=7.5 $Y2=1.97
r227 64 65 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.335 $Y=2.035
+ $X2=6.665 $Y2=2.035
r228 60 107 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=6.5 $Y=2.12
+ $X2=6.5 $Y2=2.035
r229 60 62 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=6.5 $Y=2.12
+ $X2=6.5 $Y2=2.815
r230 59 102 3.05 $w=1.7e-07 $l=9.21954e-08 $layer=LI1_cond $X=5.685 $Y=1.905
+ $X2=5.6 $Y2=1.92
r231 58 103 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.335 $Y=1.905
+ $X2=6.5 $Y2=1.905
r232 58 59 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.335 $Y=1.905
+ $X2=5.685 $Y2=1.905
r233 54 102 3.05 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=5.6 $Y=2.02 $X2=5.6
+ $Y2=1.92
r234 54 56 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=5.6 $Y=2.02
+ $X2=5.6 $Y2=2.815
r235 53 102 3.05 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=5.6 $Y=1.82 $X2=5.6
+ $Y2=1.92
r236 52 53 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.6 $Y=1.26 $X2=5.6
+ $Y2=1.82
r237 51 95 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.815 $Y=1.935
+ $X2=4.65 $Y2=1.935
r238 50 102 3.05 $w=1.7e-07 $l=9.21954e-08 $layer=LI1_cond $X=5.515 $Y=1.935
+ $X2=5.6 $Y2=1.92
r239 50 51 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.515 $Y=1.935
+ $X2=4.815 $Y2=1.935
r240 48 100 7.61436 $w=2.78e-07 $l=1.85e-07 $layer=LI1_cond $X=4.675 $Y=2.415
+ $X2=4.675 $Y2=2.23
r241 45 94 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.865 $Y=2.145
+ $X2=3.75 $Y2=2.145
r242 44 99 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.485 $Y=2.145
+ $X2=4.65 $Y2=2.145
r243 44 45 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.485 $Y=2.145
+ $X2=3.865 $Y2=2.145
r244 40 94 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.75 $Y=2.23
+ $X2=3.75 $Y2=2.145
r245 40 42 12.7771 $w=2.28e-07 $l=2.55e-07 $layer=LI1_cond $X=3.75 $Y=2.23
+ $X2=3.75 $Y2=2.485
r246 39 91 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.505 $Y=1.175
+ $X2=3.42 $Y2=1.175
r247 38 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.515 $Y=1.175
+ $X2=5.6 $Y2=1.26
r248 38 39 131.134 $w=1.68e-07 $l=2.01e-06 $layer=LI1_cond $X=5.515 $Y=1.175
+ $X2=3.505 $Y2=1.175
r249 35 90 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=0.87
+ $X2=3.42 $Y2=0.955
r250 35 37 0.717647 $w=1.7e-07 $l=1e-08 $layer=LI1_cond $X=3.42 $Y=0.87 $X2=3.42
+ $Y2=0.86
r251 34 89 6.28872 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=2.965 $Y=2.145
+ $X2=2.745 $Y2=2.145
r252 33 94 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.635 $Y=2.145
+ $X2=3.75 $Y2=2.145
r253 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.635 $Y=2.145
+ $X2=2.965 $Y2=2.145
r254 32 85 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.65 $Y=0.955
+ $X2=2.485 $Y2=0.955
r255 31 90 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=0.955
+ $X2=3.42 $Y2=0.955
r256 31 32 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.335 $Y=0.955
+ $X2=2.65 $Y2=0.955
r257 10 113 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=9.215
+ $Y=1.84 $X2=9.35 $Y2=2.115
r258 10 80 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.215
+ $Y=1.84 $X2=9.35 $Y2=2.815
r259 9 111 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=8.315
+ $Y=1.84 $X2=8.45 $Y2=2.115
r260 9 74 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.315
+ $Y=1.84 $X2=8.45 $Y2=2.815
r261 8 109 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.365
+ $Y=1.84 $X2=7.5 $Y2=1.985
r262 8 68 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.365
+ $Y=1.84 $X2=7.5 $Y2=2.815
r263 7 106 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.365
+ $Y=1.84 $X2=6.5 $Y2=1.985
r264 7 62 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.365
+ $Y=1.84 $X2=6.5 $Y2=2.815
r265 6 102 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.465
+ $Y=1.84 $X2=5.6 $Y2=1.985
r266 6 56 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.465
+ $Y=1.84 $X2=5.6 $Y2=2.815
r267 5 98 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.515
+ $Y=1.84 $X2=4.65 $Y2=2.015
r268 5 48 300 $w=1.7e-07 $l=6.38944e-07 $layer=licon1_PDIFF $count=2 $X=4.515
+ $Y=1.84 $X2=4.65 $Y2=2.415
r269 4 94 600 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_PDIFF $count=1 $X=3.615
+ $Y=1.84 $X2=3.75 $Y2=2.145
r270 4 42 300 $w=1.7e-07 $l=7.09295e-07 $layer=licon1_PDIFF $count=2 $X=3.615
+ $Y=1.84 $X2=3.75 $Y2=2.485
r271 3 121 300 $w=1.7e-07 $l=7.09295e-07 $layer=licon1_PDIFF $count=2 $X=2.665
+ $Y=1.84 $X2=2.8 $Y2=2.485
r272 3 89 600 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_PDIFF $count=1 $X=2.665
+ $Y=1.84 $X2=2.8 $Y2=2.145
r273 2 37 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=3.28
+ $Y=0.37 $X2=3.42 $Y2=0.86
r274 1 83 182 $w=1.7e-07 $l=5.27376e-07 $layer=licon1_NDIFF $count=1 $X=2.305
+ $Y=0.37 $X2=2.485 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4BB_4%VGND 1 2 3 12 16 20 22 24 29 37 44 45 48
+ 51 54
r94 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r95 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r96 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r97 45 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r98 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r99 42 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.465 $Y=0 $X2=9.3
+ $Y2=0
r100 42 44 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=9.465 $Y=0
+ $X2=9.84 $Y2=0
r101 41 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r102 41 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r103 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r104 38 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.605 $Y=0 $X2=8.44
+ $Y2=0
r105 38 40 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.605 $Y=0
+ $X2=8.88 $Y2=0
r106 37 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.135 $Y=0 $X2=9.3
+ $Y2=0
r107 37 40 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=9.135 $Y=0
+ $X2=8.88 $Y2=0
r108 36 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r109 35 36 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r110 33 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r111 32 35 438.417 $w=1.68e-07 $l=6.72e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=7.92
+ $Y2=0
r112 32 33 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r113 30 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r114 30 32 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r115 29 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.275 $Y=0 $X2=8.44
+ $Y2=0
r116 29 35 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.275 $Y=0
+ $X2=7.92 $Y2=0
r117 27 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r118 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r119 24 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r120 24 26 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r121 22 36 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=7.92 $Y2=0
r122 22 33 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=1.2
+ $Y2=0
r123 18 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.3 $Y=0.085 $X2=9.3
+ $Y2=0
r124 18 20 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=9.3 $Y=0.085
+ $X2=9.3 $Y2=0.57
r125 14 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.44 $Y=0.085
+ $X2=8.44 $Y2=0
r126 14 16 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=8.44 $Y=0.085
+ $X2=8.44 $Y2=0.57
r127 10 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0
r128 10 12 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0.325
r129 3 20 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=9.16
+ $Y=0.37 $X2=9.3 $Y2=0.57
r130 2 16 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=8.3
+ $Y=0.37 $X2=8.44 $Y2=0.57
r131 1 12 182 $w=1.7e-07 $l=3.37528e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.57 $X2=0.79 $Y2=0.325
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4BB_4%A_374_74# 1 2 3 4 5 18 20 21 22 27 28 29
+ 32 38
c63 22 0 7.06753e-20 $X=3.685 $Y=0.34
c64 20 0 7.06753e-20 $X=2.82 $Y=0.34
r65 38 40 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=5.73 $Y=0.715
+ $X2=5.73 $Y2=0.835
r66 32 35 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.985 $Y=0.34
+ $X2=2.985 $Y2=0.525
r67 29 31 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=3.935 $Y=0.835
+ $X2=4.71 $Y2=0.835
r68 28 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.565 $Y=0.835
+ $X2=5.73 $Y2=0.835
r69 28 31 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=5.565 $Y=0.835
+ $X2=4.71 $Y2=0.835
r70 25 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.81 $Y=0.75
+ $X2=3.935 $Y2=0.835
r71 25 27 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=3.81 $Y=0.75
+ $X2=3.81 $Y2=0.635
r72 24 27 9.68052 $w=2.48e-07 $l=2.1e-07 $layer=LI1_cond $X=3.81 $Y=0.425
+ $X2=3.81 $Y2=0.635
r73 23 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.15 $Y=0.34
+ $X2=2.985 $Y2=0.34
r74 22 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.685 $Y=0.34
+ $X2=3.81 $Y2=0.425
r75 22 23 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.685 $Y=0.34
+ $X2=3.15 $Y2=0.34
r76 20 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.82 $Y=0.34
+ $X2=2.985 $Y2=0.34
r77 20 21 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=2.82 $Y=0.34 $X2=2.1
+ $Y2=0.34
r78 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.015 $Y=0.425
+ $X2=2.1 $Y2=0.34
r79 16 18 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.015 $Y=0.425
+ $X2=2.015 $Y2=0.515
r80 5 38 182 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_NDIFF $count=1 $X=5.59
+ $Y=0.37 $X2=5.73 $Y2=0.715
r81 4 31 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=4.57
+ $Y=0.37 $X2=4.71 $Y2=0.835
r82 3 27 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=3.71
+ $Y=0.37 $X2=3.85 $Y2=0.635
r83 2 35 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=2.84
+ $Y=0.37 $X2=2.985 $Y2=0.525
r84 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.87
+ $Y=0.37 $X2=2.015 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4BB_4%A_828_74# 1 2 3 4 13 19 23 25 29 31 32
c51 19 0 2.42988e-20 $X=6.555 $Y=0.34
c52 13 0 1.79504e-19 $X=5.223 $Y=0.417
r53 27 29 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=7.58 $Y=0.425
+ $X2=7.58 $Y2=0.58
r54 26 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.885 $Y=0.34
+ $X2=6.72 $Y2=0.34
r55 25 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.415 $Y=0.34
+ $X2=7.58 $Y2=0.425
r56 25 26 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.415 $Y=0.34
+ $X2=6.885 $Y2=0.34
r57 21 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.72 $Y=0.425
+ $X2=6.72 $Y2=0.34
r58 21 23 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=6.72 $Y=0.425
+ $X2=6.72 $Y2=0.58
r59 19 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.555 $Y=0.34
+ $X2=6.72 $Y2=0.34
r60 19 31 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=6.555 $Y=0.34
+ $X2=5.385 $Y2=0.34
r61 15 18 33.3322 $w=3.23e-07 $l=9.4e-07 $layer=LI1_cond $X=4.28 $Y=0.417
+ $X2=5.22 $Y2=0.417
r62 13 31 8.35379 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=5.223 $Y=0.417
+ $X2=5.385 $Y2=0.417
r63 13 18 0.106379 $w=3.23e-07 $l=3e-09 $layer=LI1_cond $X=5.223 $Y=0.417
+ $X2=5.22 $Y2=0.417
r64 4 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.44
+ $Y=0.37 $X2=7.58 $Y2=0.58
r65 3 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.58
+ $Y=0.37 $X2=6.72 $Y2=0.58
r66 2 18 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=5 $Y=0.37
+ $X2=5.22 $Y2=0.495
r67 1 15 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.14
+ $Y=0.37 $X2=4.28 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4BB_4%A_1229_74# 1 2 3 4 5 18 20 21 24 26 30 32
+ 36 38 42 44 45 46
r73 40 42 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=9.8 $Y=0.96 $X2=9.8
+ $Y2=0.515
r74 39 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.955 $Y=1.045
+ $X2=8.87 $Y2=1.045
r75 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.635 $Y=1.045
+ $X2=9.8 $Y2=0.96
r76 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.635 $Y=1.045
+ $X2=8.955 $Y2=1.045
r77 34 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.87 $Y=0.96 $X2=8.87
+ $Y2=1.045
r78 34 36 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=8.87 $Y=0.96
+ $X2=8.87 $Y2=0.515
r79 33 45 5.16603 $w=1.7e-07 $l=8.9861e-08 $layer=LI1_cond $X=8.095 $Y=1.045
+ $X2=8.01 $Y2=1.055
r80 32 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.785 $Y=1.045
+ $X2=8.87 $Y2=1.045
r81 32 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.785 $Y=1.045
+ $X2=8.095 $Y2=1.045
r82 28 45 1.34256 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.01 $Y=0.96 $X2=8.01
+ $Y2=1.055
r83 28 30 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=8.01 $Y=0.96
+ $X2=8.01 $Y2=0.515
r84 27 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.235 $Y=1.065
+ $X2=7.15 $Y2=1.065
r85 26 45 5.16603 $w=1.7e-07 $l=8.9861e-08 $layer=LI1_cond $X=7.925 $Y=1.065
+ $X2=8.01 $Y2=1.055
r86 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.925 $Y=1.065
+ $X2=7.235 $Y2=1.065
r87 22 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.15 $Y=0.98 $X2=7.15
+ $Y2=1.065
r88 22 24 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=7.15 $Y=0.98
+ $X2=7.15 $Y2=0.86
r89 20 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.065 $Y=1.065
+ $X2=7.15 $Y2=1.065
r90 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.065 $Y=1.065
+ $X2=6.375 $Y2=1.065
r91 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.25 $Y=0.98
+ $X2=6.375 $Y2=1.065
r92 16 18 5.53173 $w=2.48e-07 $l=1.2e-07 $layer=LI1_cond $X=6.25 $Y=0.98
+ $X2=6.25 $Y2=0.86
r93 5 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.66
+ $Y=0.37 $X2=9.8 $Y2=0.515
r94 4 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.73
+ $Y=0.37 $X2=8.87 $Y2=0.515
r95 3 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.87
+ $Y=0.37 $X2=8.01 $Y2=0.515
r96 2 24 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=7.01
+ $Y=0.37 $X2=7.15 $Y2=0.86
r97 1 18 182 $w=1.7e-07 $l=5.57808e-07 $layer=licon1_NDIFF $count=1 $X=6.145
+ $Y=0.37 $X2=6.29 $Y2=0.86
.ends


* File: sky130_fd_sc_ms__a221oi_1.spice
* Created: Wed Sep  2 11:52:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a221oi_1.pex.spice"
.subckt sky130_fd_sc_ms__a221oi_1  VNB VPB C1 B2 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* C1	C1
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_C1_M1003_g N_Y_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.4477 PD=1.13 PS=2.69 NRD=14.592 NRS=0 M=1 R=4.93333 SA=75000.5
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1008 A_351_74# N_B2_M1008_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74 AD=0.0777
+ AS=0.1443 PD=0.95 PS=1.13 NRD=8.1 NRS=3.24 M=1 R=4.93333 SA=75001.1 SB=75001.6
+ A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_B1_M1000_g A_351_74# VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.0777 PD=1.31 PS=0.95 NRD=19.452 NRS=8.1 M=1 R=4.93333 SA=75001.4
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1006 A_567_74# N_A1_M1006_g N_Y_M1000_d VNB NLOWVT L=0.15 W=0.74 AD=0.0777
+ AS=0.2109 PD=0.95 PS=1.31 NRD=8.1 NRS=27.564 M=1 R=4.93333 SA=75002.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g A_567_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1961
+ AS=0.0777 PD=2.01 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333 SA=75002.5 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1009 N_A_121_368#_M1009_d N_C1_M1009_g N_Y_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2912 AS=0.2912 PD=2.76 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1001 N_A_121_368#_M1001_d N_B2_M1001_g N_A_263_368#_M1001_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1004 N_A_263_368#_M1004_d N_B1_M1004_g N_A_121_368#_M1001_d VPB PSHORT L=0.18
+ W=1.12 AD=0.168 AS=0.1512 PD=1.42 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_263_368#_M1004_d VPB PSHORT L=0.18 W=1.12
+ AD=0.2016 AS=0.168 PD=1.48 PS=1.42 NRD=4.3931 NRS=4.3931 M=1 R=6.22222
+ SA=90001.1 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1005 N_A_263_368#_M1005_d N_A2_M1005_g N_VPWR_M1002_d VPB PSHORT L=0.18 W=1.12
+ AD=0.2912 AS=0.2016 PD=2.76 PS=1.48 NRD=0 NRS=9.6727 M=1 R=6.22222 SA=90001.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ms__a221oi_1.pxi.spice"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 VPWR a_113_98# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 a_27_392# A4 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X2 VGND a_113_98# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VPWR A3 a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X4 a_1205_74# A4 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_27_392# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X6 a_113_98# B1 a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X7 a_113_98# A1 a_751_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_27_392# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X9 X a_113_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_751_74# A1 a_113_98# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 VPWR A1 a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X12 VPWR A4 a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X13 VGND a_113_98# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 X a_113_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 a_751_74# A2 a_1010_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 X a_113_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X17 VPWR A2 a_27_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X18 a_113_98# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 X a_113_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 VGND B1 a_113_98# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 a_27_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X22 a_1010_74# A2 a_751_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 a_1010_74# A3 a_1205_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 a_27_392# B1 a_113_98# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X25 VPWR a_113_98# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X26 a_1205_74# A3 a_1010_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 VGND A4 a_1205_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

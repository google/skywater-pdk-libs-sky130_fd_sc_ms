* NGSPICE file created from sky130_fd_sc_ms__dlxbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__dlxbp_1 D GATE VGND VNB VPB VPWR Q Q_N
M1000 VPWR a_231_74# a_373_82# VPB pshort w=840000u l=180000u
+  ad=1.95315e+12p pd=1.524e+07u as=2.352e+11p ps=2.24e+06u
M1001 a_589_392# a_27_413# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.1e+11p pd=2.42e+06u as=0p ps=0u
M1002 a_231_74# GATE VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.4685e+12p ps=1.184e+07u
M1003 a_815_124# a_231_74# a_667_80# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.028e+11p ps=2.46e+06u
M1004 a_863_98# a_667_80# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1005 VGND D a_27_413# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1006 VPWR a_863_98# a_773_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.995e+11p ps=1.79e+06u
M1007 a_863_98# a_667_80# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1008 Q_N a_1350_116# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1009 Q_N a_1350_116# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.08e+11p pd=2.79e+06u as=0p ps=0u
M1010 VPWR D a_27_413# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.31e+11p ps=2.23e+06u
M1011 a_667_80# a_373_82# a_589_80# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1012 a_589_80# a_27_413# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_231_74# GATE VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1014 a_1350_116# a_863_98# VPWR VPB pshort w=840000u l=180000u
+  ad=2.31e+11p pd=2.23e+06u as=0p ps=0u
M1015 VGND a_863_98# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1016 a_667_80# a_231_74# a_589_392# VPB pshort w=1e+06u l=180000u
+  ad=3.065e+11p pd=2.7e+06u as=0p ps=0u
M1017 VPWR a_863_98# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1018 a_1350_116# a_863_98# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1019 VGND a_231_74# a_373_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1020 VGND a_863_98# a_815_124# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_773_508# a_373_82# a_667_80# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fah_2 A B CI VGND VNB VPB VPWR COUT SUM
X0 a_1692_424# a_852_424# a_1898_424# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X1 a_852_424# a_481_379# a_416_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 VPWR a_1454_424# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 a_1898_424# a_852_424# a_2055_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X4 a_2055_424# a_1692_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X5 VPWR a_1898_424# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X6 VPWR A a_416_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X7 VPWR CI a_1692_424# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X8 VGND CI a_1692_424# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 a_517_424# B a_117_368# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X10 a_852_424# B a_416_392# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X11 VPWR B a_481_379# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X12 a_117_368# B a_852_424# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 a_481_379# a_517_424# a_1454_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X14 VGND A a_416_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 VGND B a_481_379# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 SUM a_1898_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 a_81_260# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X18 VGND a_1898_424# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_1898_424# a_517_424# a_2055_424# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X20 a_481_379# a_852_424# a_1454_424# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X21 a_416_392# B a_517_424# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X22 COUT a_1454_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X23 COUT a_1454_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 a_1692_424# a_517_424# a_1898_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X25 VGND a_81_260# a_117_368# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 a_416_392# a_481_379# a_517_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X27 VGND a_1454_424# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X28 a_1454_424# a_517_424# a_1692_424# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X29 a_2055_424# a_1692_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X30 a_81_260# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X31 a_1454_424# a_852_424# a_1692_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X32 a_517_424# a_481_379# a_117_368# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X33 a_117_368# a_481_379# a_852_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X34 SUM a_1898_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X35 VPWR a_81_260# a_117_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
.ends

* File: sky130_fd_sc_ms__xor2_4.pxi.spice
* Created: Fri Aug 28 18:19:09 2020
* 
x_PM_SKY130_FD_SC_MS__XOR2_4%A N_A_M1004_g N_A_M1001_g N_A_M1009_g N_A_M1022_g
+ N_A_M1003_g N_A_M1015_g N_A_M1006_g N_A_M1016_g N_A_M1021_g N_A_M1025_g
+ N_A_c_148_n N_A_M1026_g N_A_M1027_g N_A_c_151_n N_A_c_152_n N_A_c_153_n
+ N_A_c_318_p N_A_c_154_n N_A_c_183_p N_A_c_175_p N_A_c_178_p N_A_c_200_p
+ N_A_c_208_p N_A_c_155_n N_A_c_204_p N_A_c_176_p A A A A N_A_c_157_n
+ N_A_c_158_n N_A_c_159_n N_A_c_160_n PM_SKY130_FD_SC_MS__XOR2_4%A
x_PM_SKY130_FD_SC_MS__XOR2_4%B N_B_c_384_n N_B_M1007_g N_B_M1023_g N_B_c_385_n
+ N_B_M1011_g N_B_M1028_g N_B_c_371_n N_B_M1000_g N_B_M1010_g N_B_c_374_n
+ N_B_c_375_n N_B_M1012_g N_B_M1002_g N_B_M1005_g N_B_M1020_g N_B_M1008_g
+ N_B_c_378_n N_B_M1024_g N_B_c_380_n N_B_c_381_n N_B_c_392_n N_B_c_393_n
+ N_B_c_407_n N_B_c_382_n N_B_c_394_n N_B_c_422_n B B B B B N_B_c_383_n B
+ PM_SKY130_FD_SC_MS__XOR2_4%B
x_PM_SKY130_FD_SC_MS__XOR2_4%A_160_98# N_A_160_98#_M1001_d N_A_160_98#_M1023_d
+ N_A_160_98#_M1007_d N_A_160_98#_c_568_n N_A_160_98#_M1014_g
+ N_A_160_98#_M1013_g N_A_160_98#_M1017_g N_A_160_98#_c_569_n
+ N_A_160_98#_M1029_g N_A_160_98#_M1018_g N_A_160_98#_c_570_n
+ N_A_160_98#_c_571_n N_A_160_98#_M1019_g N_A_160_98#_c_600_n
+ N_A_160_98#_c_572_n N_A_160_98#_c_608_n N_A_160_98#_c_573_n
+ N_A_160_98#_c_574_n N_A_160_98#_c_611_n N_A_160_98#_c_575_n
+ N_A_160_98#_c_620_n PM_SKY130_FD_SC_MS__XOR2_4%A_160_98#
x_PM_SKY130_FD_SC_MS__XOR2_4%A_36_392# N_A_36_392#_M1004_d N_A_36_392#_M1009_d
+ N_A_36_392#_M1011_s N_A_36_392#_c_698_n N_A_36_392#_c_699_n
+ N_A_36_392#_c_700_n N_A_36_392#_c_713_n N_A_36_392#_c_701_n
+ N_A_36_392#_c_702_n N_A_36_392#_c_703_n PM_SKY130_FD_SC_MS__XOR2_4%A_36_392#
x_PM_SKY130_FD_SC_MS__XOR2_4%VPWR N_VPWR_M1004_s N_VPWR_M1003_s N_VPWR_M1021_s
+ N_VPWR_M1000_d N_VPWR_M1005_d N_VPWR_c_742_n N_VPWR_c_743_n N_VPWR_c_744_n
+ VPWR N_VPWR_c_745_n N_VPWR_c_746_n N_VPWR_c_747_n N_VPWR_c_748_n
+ N_VPWR_c_749_n N_VPWR_c_741_n N_VPWR_c_751_n N_VPWR_c_752_n N_VPWR_c_753_n
+ N_VPWR_c_754_n N_VPWR_c_755_n PM_SKY130_FD_SC_MS__XOR2_4%VPWR
x_PM_SKY130_FD_SC_MS__XOR2_4%A_514_368# N_A_514_368#_M1013_s
+ N_A_514_368#_M1017_s N_A_514_368#_M1019_s N_A_514_368#_M1006_d
+ N_A_514_368#_M1026_d N_A_514_368#_M1002_s N_A_514_368#_M1008_s
+ N_A_514_368#_c_858_n N_A_514_368#_c_859_n N_A_514_368#_c_860_n
+ N_A_514_368#_c_965_p N_A_514_368#_c_861_n N_A_514_368#_c_868_n
+ N_A_514_368#_c_956_p N_A_514_368#_c_862_n N_A_514_368#_c_887_n
+ N_A_514_368#_c_889_n N_A_514_368#_c_863_n N_A_514_368#_c_864_n
+ N_A_514_368#_c_873_n N_A_514_368#_c_865_n N_A_514_368#_c_866_n
+ N_A_514_368#_c_867_n PM_SKY130_FD_SC_MS__XOR2_4%A_514_368#
x_PM_SKY130_FD_SC_MS__XOR2_4%X N_X_M1014_s N_X_M1010_d N_X_M1020_d N_X_M1013_d
+ N_X_M1018_d N_X_c_968_n N_X_c_969_n N_X_c_987_n N_X_c_970_n N_X_c_971_n
+ N_X_c_1004_n N_X_c_978_n N_X_c_1007_n N_X_c_1009_n N_X_c_972_n N_X_c_1126_p
+ N_X_c_973_n N_X_c_974_n N_X_c_1044_n N_X_c_975_n N_X_c_976_n N_X_c_977_n X
+ N_X_c_1051_n N_X_c_1013_n PM_SKY130_FD_SC_MS__XOR2_4%X
x_PM_SKY130_FD_SC_MS__XOR2_4%VGND N_VGND_M1001_s N_VGND_M1022_s N_VGND_M1028_s
+ N_VGND_M1029_d N_VGND_M1015_d N_VGND_M1025_d N_VGND_c_1132_n N_VGND_c_1133_n
+ N_VGND_c_1134_n N_VGND_c_1135_n N_VGND_c_1136_n N_VGND_c_1137_n
+ N_VGND_c_1138_n N_VGND_c_1139_n N_VGND_c_1140_n N_VGND_c_1141_n VGND
+ N_VGND_c_1142_n N_VGND_c_1143_n N_VGND_c_1144_n N_VGND_c_1145_n
+ N_VGND_c_1146_n N_VGND_c_1147_n N_VGND_c_1148_n N_VGND_c_1149_n
+ PM_SKY130_FD_SC_MS__XOR2_4%VGND
x_PM_SKY130_FD_SC_MS__XOR2_4%A_877_74# N_A_877_74#_M1015_s N_A_877_74#_M1016_s
+ N_A_877_74#_M1027_s N_A_877_74#_M1012_s N_A_877_74#_M1024_s
+ N_A_877_74#_c_1261_n N_A_877_74#_c_1263_n N_A_877_74#_c_1254_n
+ N_A_877_74#_c_1255_n N_A_877_74#_c_1278_n N_A_877_74#_c_1256_n
+ N_A_877_74#_c_1257_n N_A_877_74#_c_1258_n N_A_877_74#_c_1268_n
+ N_A_877_74#_c_1259_n N_A_877_74#_c_1260_n PM_SKY130_FD_SC_MS__XOR2_4%A_877_74#
cc_1 VNB N_A_M1001_g 0.0234074f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.86
cc_2 VNB N_A_M1022_g 0.0225154f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=0.86
cc_3 VNB N_A_M1015_g 0.0328409f $X=-0.19 $Y=-0.245 $X2=4.745 $Y2=0.74
cc_4 VNB N_A_M1016_g 0.025165f $X=-0.19 $Y=-0.245 $X2=5.335 $Y2=0.74
cc_5 VNB N_A_M1025_g 0.025165f $X=-0.19 $Y=-0.245 $X2=5.765 $Y2=0.74
cc_6 VNB N_A_c_148_n 0.0241073f $X=-0.19 $Y=-0.245 $X2=6.255 $Y2=1.485
cc_7 VNB N_A_M1026_g 0.00193523f $X=-0.19 $Y=-0.245 $X2=6.345 $Y2=2.4
cc_8 VNB N_A_M1027_g 0.025058f $X=-0.19 $Y=-0.245 $X2=6.355 $Y2=0.74
cc_9 VNB N_A_c_151_n 0.0153274f $X=-0.19 $Y=-0.245 $X2=4.712 $Y2=1.515
cc_10 VNB N_A_c_152_n 0.00875513f $X=-0.19 $Y=-0.245 $X2=6.345 $Y2=1.485
cc_11 VNB N_A_c_153_n 0.00598948f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.42
cc_12 VNB N_A_c_154_n 0.0125135f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.585
cc_13 VNB N_A_c_155_n 0.00557768f $X=-0.19 $Y=-0.245 $X2=3.85 $Y2=1.35
cc_14 VNB A 0.00199724f $X=-0.19 $Y=-0.245 $X2=5.435 $Y2=1.58
cc_15 VNB N_A_c_157_n 0.0196122f $X=-0.19 $Y=-0.245 $X2=5.225 $Y2=1.515
cc_16 VNB N_A_c_158_n 0.0422363f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=1.585
cc_17 VNB N_A_c_159_n 0.023877f $X=-0.19 $Y=-0.245 $X2=5.855 $Y2=1.515
cc_18 VNB N_A_c_160_n 0.00798232f $X=-0.19 $Y=-0.245 $X2=4.39 $Y2=1.562
cc_19 VNB N_B_M1023_g 0.0256964f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.86
cc_20 VNB N_B_M1028_g 0.0260782f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.42
cc_21 VNB N_B_c_371_n 0.00565832f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=0.86
cc_22 VNB N_B_M1000_g 0.0179606f $X=-0.19 $Y=-0.245 $X2=4.725 $Y2=1.68
cc_23 VNB N_B_M1010_g 0.00619066f $X=-0.19 $Y=-0.245 $X2=4.745 $Y2=0.74
cc_24 VNB N_B_c_374_n 0.0283688f $X=-0.19 $Y=-0.245 $X2=4.745 $Y2=0.74
cc_25 VNB N_B_c_375_n 0.0115262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B_M1012_g 0.00656268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B_M1020_g 0.0230909f $X=-0.19 $Y=-0.245 $X2=5.765 $Y2=0.74
cc_28 VNB N_B_c_378_n 0.0683506f $X=-0.19 $Y=-0.245 $X2=6.345 $Y2=2.4
cc_29 VNB N_B_M1024_g 0.0260971f $X=-0.19 $Y=-0.245 $X2=6.355 $Y2=1.35
cc_30 VNB N_B_c_380_n 0.00100736f $X=-0.19 $Y=-0.245 $X2=4.712 $Y2=1.515
cc_31 VNB N_B_c_381_n 0.0378961f $X=-0.19 $Y=-0.245 $X2=6.345 $Y2=1.485
cc_32 VNB N_B_c_382_n 4.22572e-19 $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.585
cc_33 VNB N_B_c_383_n 0.00498375f $X=-0.19 $Y=-0.245 $X2=5.315 $Y2=1.515
cc_34 VNB N_A_160_98#_c_568_n 0.020942f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=2.46
cc_35 VNB N_A_160_98#_c_569_n 0.020159f $X=-0.19 $Y=-0.245 $X2=4.745 $Y2=1.35
cc_36 VNB N_A_160_98#_c_570_n 0.0202979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_160_98#_c_571_n 0.069959f $X=-0.19 $Y=-0.245 $X2=5.335 $Y2=1.35
cc_38 VNB N_A_160_98#_c_572_n 0.00258679f $X=-0.19 $Y=-0.245 $X2=5.765 $Y2=0.74
cc_39 VNB N_A_160_98#_c_573_n 0.00234522f $X=-0.19 $Y=-0.245 $X2=6.345 $Y2=2.4
cc_40 VNB N_A_160_98#_c_574_n 0.00241736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_160_98#_c_575_n 0.00188856f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.665
cc_42 VNB N_VPWR_c_741_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.585
cc_43 VNB N_X_c_968_n 0.00435724f $X=-0.19 $Y=-0.245 $X2=4.725 $Y2=2.4
cc_44 VNB N_X_c_969_n 0.00276895f $X=-0.19 $Y=-0.245 $X2=4.745 $Y2=1.35
cc_45 VNB N_X_c_970_n 0.0209692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_X_c_971_n 0.00207986f $X=-0.19 $Y=-0.245 $X2=5.315 $Y2=1.68
cc_47 VNB N_X_c_972_n 0.0025951f $X=-0.19 $Y=-0.245 $X2=5.765 $Y2=2.4
cc_48 VNB N_X_c_973_n 0.0112366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_X_c_974_n 0.0222851f $X=-0.19 $Y=-0.245 $X2=6.345 $Y2=1.62
cc_50 VNB N_X_c_975_n 0.00345724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_X_c_976_n 0.00253527f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.75
cc_52 VNB N_X_c_977_n 0.00124931f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.42
cc_53 VNB N_VGND_c_1132_n 0.01004f $X=-0.19 $Y=-0.245 $X2=4.725 $Y2=2.4
cc_54 VNB N_VGND_c_1133_n 0.0567336f $X=-0.19 $Y=-0.245 $X2=4.745 $Y2=1.35
cc_55 VNB N_VGND_c_1134_n 0.015878f $X=-0.19 $Y=-0.245 $X2=5.315 $Y2=1.68
cc_56 VNB N_VGND_c_1135_n 0.015091f $X=-0.19 $Y=-0.245 $X2=5.335 $Y2=1.35
cc_57 VNB N_VGND_c_1136_n 0.00790705f $X=-0.19 $Y=-0.245 $X2=5.765 $Y2=1.68
cc_58 VNB N_VGND_c_1137_n 0.0075298f $X=-0.19 $Y=-0.245 $X2=5.765 $Y2=1.35
cc_59 VNB N_VGND_c_1138_n 0.0218315f $X=-0.19 $Y=-0.245 $X2=5.765 $Y2=0.74
cc_60 VNB N_VGND_c_1139_n 0.0260634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1140_n 0.026797f $X=-0.19 $Y=-0.245 $X2=6.355 $Y2=1.35
cc_62 VNB N_VGND_c_1141_n 0.00795087f $X=-0.19 $Y=-0.245 $X2=6.355 $Y2=0.74
cc_63 VNB N_VGND_c_1142_n 0.0216203f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.42
cc_64 VNB N_VGND_c_1143_n 0.0202269f $X=-0.19 $Y=-0.245 $X2=2.87 $Y2=0.685
cc_65 VNB N_VGND_c_1144_n 0.0178371f $X=-0.19 $Y=-0.245 $X2=3.765 $Y2=1.105
cc_66 VNB N_VGND_c_1145_n 0.0576436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1146_n 0.471044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1147_n 0.00631222f $X=-0.19 $Y=-0.245 $X2=5.11 $Y2=1.515
cc_69 VNB N_VGND_c_1148_n 0.00631651f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.585
cc_70 VNB N_VGND_c_1149_n 0.00631651f $X=-0.19 $Y=-0.245 $X2=5.315 $Y2=1.515
cc_71 VNB N_A_877_74#_c_1254_n 6.9777e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_877_74#_c_1255_n 0.00163372f $X=-0.19 $Y=-0.245 $X2=5.315 $Y2=1.68
cc_73 VNB N_A_877_74#_c_1256_n 0.011697f $X=-0.19 $Y=-0.245 $X2=5.335 $Y2=0.74
cc_74 VNB N_A_877_74#_c_1257_n 0.0164799f $X=-0.19 $Y=-0.245 $X2=5.765 $Y2=2.4
cc_75 VNB N_A_877_74#_c_1258_n 0.00217595f $X=-0.19 $Y=-0.245 $X2=5.765 $Y2=1.35
cc_76 VNB N_A_877_74#_c_1259_n 0.00239138f $X=-0.19 $Y=-0.245 $X2=6.255
+ $Y2=1.485
cc_77 VNB N_A_877_74#_c_1260_n 0.00220733f $X=-0.19 $Y=-0.245 $X2=6.345 $Y2=2.4
cc_78 VPB N_A_M1004_g 0.0337676f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=2.46
cc_79 VPB N_A_M1009_g 0.0242742f $X=-0.19 $Y=1.66 $X2=1.05 $Y2=2.46
cc_80 VPB N_A_M1003_g 0.0217564f $X=-0.19 $Y=1.66 $X2=4.725 $Y2=2.4
cc_81 VPB N_A_M1006_g 0.0219548f $X=-0.19 $Y=1.66 $X2=5.315 $Y2=2.4
cc_82 VPB N_A_M1021_g 0.0218933f $X=-0.19 $Y=1.66 $X2=5.765 $Y2=2.4
cc_83 VPB N_A_M1026_g 0.0233105f $X=-0.19 $Y=1.66 $X2=6.345 $Y2=2.4
cc_84 VPB N_A_c_151_n 0.00154547f $X=-0.19 $Y=1.66 $X2=4.712 $Y2=1.515
cc_85 VPB N_A_c_154_n 0.00380335f $X=-0.19 $Y=1.66 $X2=0.685 $Y2=1.585
cc_86 VPB A 0.00880428f $X=-0.19 $Y=1.66 $X2=5.435 $Y2=1.58
cc_87 VPB N_A_c_157_n 0.00743058f $X=-0.19 $Y=1.66 $X2=5.225 $Y2=1.515
cc_88 VPB N_A_c_158_n 0.0153572f $X=-0.19 $Y=1.66 $X2=1.05 $Y2=1.585
cc_89 VPB N_A_c_159_n 0.0042616f $X=-0.19 $Y=1.66 $X2=5.855 $Y2=1.515
cc_90 VPB N_A_c_160_n 0.00330362f $X=-0.19 $Y=1.66 $X2=4.39 $Y2=1.562
cc_91 VPB N_B_c_384_n 0.0150006f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=1.75
cc_92 VPB N_B_c_385_n 0.0214133f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_B_M1000_g 0.0211867f $X=-0.19 $Y=1.66 $X2=4.725 $Y2=1.68
cc_94 VPB N_B_M1002_g 0.020498f $X=-0.19 $Y=1.66 $X2=5.335 $Y2=0.74
cc_95 VPB N_B_M1005_g 0.0204965f $X=-0.19 $Y=1.66 $X2=5.765 $Y2=2.4
cc_96 VPB N_B_M1008_g 0.025344f $X=-0.19 $Y=1.66 $X2=6.345 $Y2=1.62
cc_97 VPB N_B_c_378_n 0.00820157f $X=-0.19 $Y=1.66 $X2=6.345 $Y2=2.4
cc_98 VPB N_B_c_381_n 0.0423235f $X=-0.19 $Y=1.66 $X2=6.345 $Y2=1.485
cc_99 VPB N_B_c_392_n 0.00968953f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.42
cc_100 VPB N_B_c_393_n 0.00115796f $X=-0.19 $Y=1.66 $X2=1.275 $Y2=0.665
cc_101 VPB N_B_c_394_n 6.1801e-19 $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.585
cc_102 VPB N_B_c_383_n 0.013618f $X=-0.19 $Y=1.66 $X2=5.315 $Y2=1.515
cc_103 VPB N_A_160_98#_M1013_g 0.0240583f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=0.86
cc_104 VPB N_A_160_98#_M1017_g 0.0204563f $X=-0.19 $Y=1.66 $X2=4.725 $Y2=2.4
cc_105 VPB N_A_160_98#_M1018_g 0.0204319f $X=-0.19 $Y=1.66 $X2=5.315 $Y2=2.4
cc_106 VPB N_A_160_98#_c_570_n 0.0037599f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_160_98#_c_571_n 0.0141901f $X=-0.19 $Y=1.66 $X2=5.335 $Y2=1.35
cc_108 VPB N_A_160_98#_M1019_g 0.0197764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_160_98#_c_572_n 0.00106568f $X=-0.19 $Y=1.66 $X2=5.765 $Y2=0.74
cc_110 VPB N_A_160_98#_c_574_n 0.00170979f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_36_392#_c_698_n 0.0363954f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_36_392#_c_699_n 0.00927999f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_36_392#_c_700_n 0.014412f $X=-0.19 $Y=1.66 $X2=4.725 $Y2=1.68
cc_114 VPB N_A_36_392#_c_701_n 0.00632687f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_36_392#_c_702_n 0.00160153f $X=-0.19 $Y=1.66 $X2=5.315 $Y2=1.68
cc_116 VPB N_A_36_392#_c_703_n 0.00668387f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_742_n 0.00845772f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_743_n 0.00495786f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_744_n 0.00797179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_745_n 0.0908753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_746_n 0.018101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_747_n 0.0175244f $X=-0.19 $Y=1.66 $X2=6.345 $Y2=2.4
cc_123 VPB N_VPWR_c_748_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_749_n 0.0197879f $X=-0.19 $Y=1.66 $X2=0.685 $Y2=0.665
cc_125 VPB N_VPWR_c_741_n 0.0960064f $X=-0.19 $Y=1.66 $X2=0.685 $Y2=1.585
cc_126 VPB N_VPWR_c_751_n 0.0263173f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.585
cc_127 VPB N_VPWR_c_752_n 0.0141186f $X=-0.19 $Y=1.66 $X2=1.445 $Y2=0.685
cc_128 VPB N_VPWR_c_753_n 0.0138857f $X=-0.19 $Y=1.66 $X2=1.275 $Y2=0.675
cc_129 VPB N_VPWR_c_754_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_755_n 0.00324402f $X=-0.19 $Y=1.66 $X2=5.225 $Y2=1.515
cc_131 VPB N_A_514_368#_c_858_n 0.00658249f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_514_368#_c_859_n 0.0026202f $X=-0.19 $Y=1.66 $X2=5.315 $Y2=2.4
cc_133 VPB N_A_514_368#_c_860_n 0.00369664f $X=-0.19 $Y=1.66 $X2=5.315 $Y2=2.4
cc_134 VPB N_A_514_368#_c_861_n 0.00284344f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_514_368#_c_862_n 0.00173277f $X=-0.19 $Y=1.66 $X2=5.765 $Y2=0.74
cc_136 VPB N_A_514_368#_c_863_n 0.00121438f $X=-0.19 $Y=1.66 $X2=6.355 $Y2=0.74
cc_137 VPB N_A_514_368#_c_864_n 0.0017942f $X=-0.19 $Y=1.66 $X2=6.355 $Y2=0.74
cc_138 VPB N_A_514_368#_c_865_n 0.0022923f $X=-0.19 $Y=1.66 $X2=0.685 $Y2=1.585
cc_139 VPB N_A_514_368#_c_866_n 0.00231675f $X=-0.19 $Y=1.66 $X2=1.445 $Y2=0.685
cc_140 VPB N_A_514_368#_c_867_n 0.0308267f $X=-0.19 $Y=1.66 $X2=2.955 $Y2=1.02
cc_141 VPB N_X_c_978_n 0.00692367f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_X_c_974_n 0.00832134f $X=-0.19 $Y=1.66 $X2=6.345 $Y2=1.62
cc_143 N_A_M1022_g N_B_M1023_g 0.0289814f $X=1.155 $Y=0.86 $X2=0 $Y2=0
cc_144 N_A_c_175_p N_B_M1023_g 0.0124999f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_145 N_A_c_176_p N_B_M1023_g 5.1812e-19 $X=1.445 $Y=0.675 $X2=0 $Y2=0
cc_146 N_A_c_175_p N_B_M1028_g 0.0125312f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_147 N_A_c_178_p N_B_M1028_g 9.06409e-19 $X=2.955 $Y=1.02 $X2=0 $Y2=0
cc_148 N_A_M1027_g N_B_c_371_n 0.00858677f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A_c_152_n N_B_M1000_g 0.0501047f $X=6.345 $Y=1.485 $X2=0 $Y2=0
cc_150 N_A_M1027_g N_B_c_375_n 0.024894f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A_M1009_g N_B_c_381_n 0.013241f $X=1.05 $Y=2.46 $X2=0 $Y2=0
cc_152 N_A_c_183_p N_B_c_381_n 0.00117645f $X=0.945 $Y=1.585 $X2=0 $Y2=0
cc_153 N_A_c_158_n N_B_c_381_n 0.0182552f $X=1.05 $Y=1.585 $X2=0 $Y2=0
cc_154 N_A_M1003_g N_B_c_407_n 0.0123498f $X=4.725 $Y=2.4 $X2=0 $Y2=0
cc_155 N_A_M1006_g N_B_c_407_n 0.0123635f $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A_M1021_g N_B_c_407_n 0.0145288f $X=5.765 $Y=2.4 $X2=0 $Y2=0
cc_157 N_A_M1026_g N_B_c_407_n 6.7865e-19 $X=6.345 $Y=2.4 $X2=0 $Y2=0
cc_158 A N_B_c_407_n 0.0865621f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_159 N_A_c_157_n N_B_c_407_n 0.00126836f $X=5.225 $Y=1.515 $X2=0 $Y2=0
cc_160 N_A_c_159_n N_B_c_407_n 4.96096e-19 $X=5.855 $Y=1.515 $X2=0 $Y2=0
cc_161 N_A_c_160_n N_B_c_407_n 0.0365387f $X=4.39 $Y=1.562 $X2=0 $Y2=0
cc_162 N_A_M1021_g N_B_c_382_n 0.00286779f $X=5.765 $Y=2.4 $X2=0 $Y2=0
cc_163 N_A_c_148_n N_B_c_382_n 0.00798799f $X=6.255 $Y=1.485 $X2=0 $Y2=0
cc_164 A N_B_c_382_n 0.031682f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_165 N_A_c_159_n N_B_c_382_n 0.00453713f $X=5.855 $Y=1.515 $X2=0 $Y2=0
cc_166 N_A_M1006_g N_B_c_394_n 8.17229e-19 $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_167 N_A_M1021_g N_B_c_394_n 0.00465905f $X=5.765 $Y=2.4 $X2=0 $Y2=0
cc_168 N_A_M1026_g N_B_c_394_n 0.0031513f $X=6.345 $Y=2.4 $X2=0 $Y2=0
cc_169 N_A_c_200_p N_B_c_422_n 0.00146645f $X=3.765 $Y=1.105 $X2=0 $Y2=0
cc_170 N_A_c_148_n N_B_c_383_n 0.0122919f $X=6.255 $Y=1.485 $X2=0 $Y2=0
cc_171 N_A_M1026_g N_B_c_383_n 0.00951454f $X=6.345 $Y=2.4 $X2=0 $Y2=0
cc_172 N_A_c_152_n N_B_c_383_n 0.0101955f $X=6.345 $Y=1.485 $X2=0 $Y2=0
cc_173 N_A_c_204_p N_A_160_98#_M1001_d 0.00439657f $X=1.275 $Y=0.675 $X2=-0.19
+ $Y2=-0.245
cc_174 N_A_c_175_p N_A_160_98#_M1023_d 0.00782857f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_175 N_A_c_175_p N_A_160_98#_c_568_n 0.0115801f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_176 N_A_c_178_p N_A_160_98#_c_568_n 0.00775701f $X=2.955 $Y=1.02 $X2=0 $Y2=0
cc_177 N_A_c_208_p N_A_160_98#_c_568_n 0.00681965f $X=3.04 $Y=1.105 $X2=0 $Y2=0
cc_178 N_A_c_178_p N_A_160_98#_c_569_n 0.00271318f $X=2.955 $Y=1.02 $X2=0 $Y2=0
cc_179 N_A_c_200_p N_A_160_98#_c_569_n 0.0140661f $X=3.765 $Y=1.105 $X2=0 $Y2=0
cc_180 N_A_c_155_n N_A_160_98#_c_569_n 0.00585519f $X=3.85 $Y=1.35 $X2=0 $Y2=0
cc_181 N_A_c_160_n N_A_160_98#_M1018_g 0.00302426f $X=4.39 $Y=1.562 $X2=0 $Y2=0
cc_182 N_A_c_151_n N_A_160_98#_c_570_n 0.00831704f $X=4.712 $Y=1.515 $X2=0 $Y2=0
cc_183 N_A_c_160_n N_A_160_98#_c_570_n 0.0191404f $X=4.39 $Y=1.562 $X2=0 $Y2=0
cc_184 N_A_c_175_p N_A_160_98#_c_571_n 0.00181746f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_185 N_A_c_200_p N_A_160_98#_c_571_n 0.0125306f $X=3.765 $Y=1.105 $X2=0 $Y2=0
cc_186 N_A_c_160_n N_A_160_98#_c_571_n 0.0129583f $X=4.39 $Y=1.562 $X2=0 $Y2=0
cc_187 N_A_M1003_g N_A_160_98#_M1019_g 0.0523968f $X=4.725 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A_c_160_n N_A_160_98#_M1019_g 0.0060375f $X=4.39 $Y=1.562 $X2=0 $Y2=0
cc_189 N_A_M1022_g N_A_160_98#_c_600_n 0.0139847f $X=1.155 $Y=0.86 $X2=0 $Y2=0
cc_190 N_A_c_183_p N_A_160_98#_c_600_n 2.60315e-19 $X=0.945 $Y=1.585 $X2=0 $Y2=0
cc_191 N_A_c_204_p N_A_160_98#_c_600_n 0.00795398f $X=1.275 $Y=0.675 $X2=0 $Y2=0
cc_192 N_A_c_176_p N_A_160_98#_c_600_n 0.0204402f $X=1.445 $Y=0.675 $X2=0 $Y2=0
cc_193 N_A_M1009_g N_A_160_98#_c_572_n 2.76068e-19 $X=1.05 $Y=2.46 $X2=0 $Y2=0
cc_194 N_A_M1022_g N_A_160_98#_c_572_n 0.00431001f $X=1.155 $Y=0.86 $X2=0 $Y2=0
cc_195 N_A_c_183_p N_A_160_98#_c_572_n 0.0118099f $X=0.945 $Y=1.585 $X2=0 $Y2=0
cc_196 N_A_c_158_n N_A_160_98#_c_572_n 0.00186962f $X=1.05 $Y=1.585 $X2=0 $Y2=0
cc_197 N_A_c_175_p N_A_160_98#_c_608_n 0.053955f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_198 N_A_c_178_p N_A_160_98#_c_608_n 0.00628036f $X=2.955 $Y=1.02 $X2=0 $Y2=0
cc_199 N_A_c_208_p N_A_160_98#_c_608_n 0.0148586f $X=3.04 $Y=1.105 $X2=0 $Y2=0
cc_200 N_A_c_175_p N_A_160_98#_c_611_n 0.00371196f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_201 N_A_c_200_p N_A_160_98#_c_611_n 0.0385816f $X=3.765 $Y=1.105 $X2=0 $Y2=0
cc_202 N_A_c_208_p N_A_160_98#_c_611_n 0.0111271f $X=3.04 $Y=1.105 $X2=0 $Y2=0
cc_203 N_A_c_160_n N_A_160_98#_c_611_n 0.0213902f $X=4.39 $Y=1.562 $X2=0 $Y2=0
cc_204 N_A_M1022_g N_A_160_98#_c_575_n 0.00279462f $X=1.155 $Y=0.86 $X2=0 $Y2=0
cc_205 N_A_c_153_n N_A_160_98#_c_575_n 0.0118907f $X=0.6 $Y=1.42 $X2=0 $Y2=0
cc_206 N_A_c_183_p N_A_160_98#_c_575_n 0.0196847f $X=0.945 $Y=1.585 $X2=0 $Y2=0
cc_207 N_A_c_204_p N_A_160_98#_c_575_n 0.0144338f $X=1.275 $Y=0.675 $X2=0 $Y2=0
cc_208 N_A_c_158_n N_A_160_98#_c_575_n 0.00267222f $X=1.05 $Y=1.585 $X2=0 $Y2=0
cc_209 N_A_c_175_p N_A_160_98#_c_620_n 0.0149765f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_210 N_A_M1004_g N_A_36_392#_c_698_n 0.0127027f $X=0.55 $Y=2.46 $X2=0 $Y2=0
cc_211 N_A_M1009_g N_A_36_392#_c_698_n 6.46187e-19 $X=1.05 $Y=2.46 $X2=0 $Y2=0
cc_212 N_A_M1004_g N_A_36_392#_c_699_n 0.013221f $X=0.55 $Y=2.46 $X2=0 $Y2=0
cc_213 N_A_M1009_g N_A_36_392#_c_699_n 0.0155386f $X=1.05 $Y=2.46 $X2=0 $Y2=0
cc_214 N_A_c_154_n N_A_36_392#_c_699_n 0.0148795f $X=0.685 $Y=1.585 $X2=0 $Y2=0
cc_215 N_A_c_183_p N_A_36_392#_c_699_n 0.0313107f $X=0.945 $Y=1.585 $X2=0 $Y2=0
cc_216 N_A_c_158_n N_A_36_392#_c_699_n 0.00728628f $X=1.05 $Y=1.585 $X2=0 $Y2=0
cc_217 N_A_M1004_g N_A_36_392#_c_700_n 0.00168649f $X=0.55 $Y=2.46 $X2=0 $Y2=0
cc_218 N_A_c_154_n N_A_36_392#_c_700_n 0.00410213f $X=0.685 $Y=1.585 $X2=0 $Y2=0
cc_219 N_A_M1004_g N_A_36_392#_c_713_n 6.01834e-19 $X=0.55 $Y=2.46 $X2=0 $Y2=0
cc_220 N_A_M1009_g N_A_36_392#_c_713_n 0.0106703f $X=1.05 $Y=2.46 $X2=0 $Y2=0
cc_221 N_A_M1009_g N_A_36_392#_c_702_n 0.00337536f $X=1.05 $Y=2.46 $X2=0 $Y2=0
cc_222 N_A_M1004_g N_VPWR_c_742_n 0.00306788f $X=0.55 $Y=2.46 $X2=0 $Y2=0
cc_223 N_A_M1009_g N_VPWR_c_742_n 0.00137311f $X=1.05 $Y=2.46 $X2=0 $Y2=0
cc_224 N_A_M1026_g N_VPWR_c_743_n 3.90993e-19 $X=6.345 $Y=2.4 $X2=0 $Y2=0
cc_225 N_A_M1009_g N_VPWR_c_745_n 0.00517089f $X=1.05 $Y=2.46 $X2=0 $Y2=0
cc_226 N_A_M1003_g N_VPWR_c_745_n 0.00371808f $X=4.725 $Y=2.4 $X2=0 $Y2=0
cc_227 N_A_M1006_g N_VPWR_c_746_n 0.0037329f $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_228 N_A_M1021_g N_VPWR_c_746_n 0.00422125f $X=5.765 $Y=2.4 $X2=0 $Y2=0
cc_229 N_A_M1026_g N_VPWR_c_747_n 0.00377953f $X=6.345 $Y=2.4 $X2=0 $Y2=0
cc_230 N_A_M1004_g N_VPWR_c_741_n 0.00986643f $X=0.55 $Y=2.46 $X2=0 $Y2=0
cc_231 N_A_M1009_g N_VPWR_c_741_n 0.00977404f $X=1.05 $Y=2.46 $X2=0 $Y2=0
cc_232 N_A_M1003_g N_VPWR_c_741_n 0.00459002f $X=4.725 $Y=2.4 $X2=0 $Y2=0
cc_233 N_A_M1006_g N_VPWR_c_741_n 0.00460941f $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_234 N_A_M1021_g N_VPWR_c_741_n 0.00633653f $X=5.765 $Y=2.4 $X2=0 $Y2=0
cc_235 N_A_M1026_g N_VPWR_c_741_n 0.00467157f $X=6.345 $Y=2.4 $X2=0 $Y2=0
cc_236 N_A_M1004_g N_VPWR_c_751_n 0.005209f $X=0.55 $Y=2.46 $X2=0 $Y2=0
cc_237 N_A_M1003_g N_VPWR_c_752_n 0.00151179f $X=4.725 $Y=2.4 $X2=0 $Y2=0
cc_238 N_A_M1006_g N_VPWR_c_752_n 0.00339137f $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_239 N_A_M1021_g N_VPWR_c_753_n 0.00339727f $X=5.765 $Y=2.4 $X2=0 $Y2=0
cc_240 N_A_M1026_g N_VPWR_c_753_n 0.00196535f $X=6.345 $Y=2.4 $X2=0 $Y2=0
cc_241 N_A_M1021_g N_A_514_368#_c_868_n 0.00887184f $X=5.765 $Y=2.4 $X2=0 $Y2=0
cc_242 N_A_M1026_g N_A_514_368#_c_868_n 0.0124647f $X=6.345 $Y=2.4 $X2=0 $Y2=0
cc_243 N_A_M1026_g N_A_514_368#_c_862_n 2.2826e-19 $X=6.345 $Y=2.4 $X2=0 $Y2=0
cc_244 N_A_M1003_g N_A_514_368#_c_864_n 0.00733114f $X=4.725 $Y=2.4 $X2=0 $Y2=0
cc_245 N_A_M1006_g N_A_514_368#_c_864_n 8.68995e-19 $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_246 N_A_M1003_g N_A_514_368#_c_873_n 0.0102985f $X=4.725 $Y=2.4 $X2=0 $Y2=0
cc_247 N_A_M1006_g N_A_514_368#_c_873_n 0.00975355f $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_248 N_A_M1003_g N_A_514_368#_c_865_n 7.69308e-19 $X=4.725 $Y=2.4 $X2=0 $Y2=0
cc_249 N_A_M1006_g N_A_514_368#_c_865_n 0.00511754f $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_250 N_A_M1021_g N_A_514_368#_c_865_n 0.00508969f $X=5.765 $Y=2.4 $X2=0 $Y2=0
cc_251 N_A_M1026_g N_A_514_368#_c_865_n 7.72861e-19 $X=6.345 $Y=2.4 $X2=0 $Y2=0
cc_252 N_A_c_175_p N_X_M1014_s 0.00223669f $X=2.87 $Y=0.685 $X2=-0.19 $Y2=-0.245
cc_253 N_A_c_178_p N_X_M1014_s 0.00327917f $X=2.955 $Y=1.02 $X2=-0.19 $Y2=-0.245
cc_254 N_A_c_200_p N_X_M1014_s 0.0144824f $X=3.765 $Y=1.105 $X2=-0.19 $Y2=-0.245
cc_255 N_A_c_208_p N_X_M1014_s 3.64502e-19 $X=3.04 $Y=1.105 $X2=-0.19 $Y2=-0.245
cc_256 N_A_c_200_p N_X_c_968_n 0.0250503f $X=3.765 $Y=1.105 $X2=0 $Y2=0
cc_257 N_A_c_160_n N_X_c_968_n 0.00617915f $X=4.39 $Y=1.562 $X2=0 $Y2=0
cc_258 N_A_M1015_g N_X_c_969_n 0.00402271f $X=4.745 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A_M1003_g N_X_c_987_n 0.0123486f $X=4.725 $Y=2.4 $X2=0 $Y2=0
cc_260 N_A_M1006_g N_X_c_987_n 0.0124022f $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_261 N_A_M1021_g N_X_c_987_n 0.0122933f $X=5.765 $Y=2.4 $X2=0 $Y2=0
cc_262 N_A_c_148_n N_X_c_987_n 8.01427e-19 $X=6.255 $Y=1.485 $X2=0 $Y2=0
cc_263 N_A_M1026_g N_X_c_987_n 0.00584183f $X=6.345 $Y=2.4 $X2=0 $Y2=0
cc_264 N_A_M1015_g N_X_c_970_n 0.0131565f $X=4.745 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A_M1016_g N_X_c_970_n 0.0112941f $X=5.335 $Y=0.74 $X2=0 $Y2=0
cc_266 N_A_M1025_g N_X_c_970_n 0.0150594f $X=5.765 $Y=0.74 $X2=0 $Y2=0
cc_267 N_A_c_148_n N_X_c_970_n 0.00506351f $X=6.255 $Y=1.485 $X2=0 $Y2=0
cc_268 N_A_M1027_g N_X_c_970_n 0.0112465f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A_c_151_n N_X_c_970_n 0.00159523f $X=4.712 $Y=1.515 $X2=0 $Y2=0
cc_270 A N_X_c_970_n 0.0950924f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_271 N_A_c_157_n N_X_c_970_n 0.00596724f $X=5.225 $Y=1.515 $X2=0 $Y2=0
cc_272 N_A_c_159_n N_X_c_970_n 0.00230115f $X=5.855 $Y=1.515 $X2=0 $Y2=0
cc_273 N_A_c_160_n N_X_c_970_n 0.00930879f $X=4.39 $Y=1.562 $X2=0 $Y2=0
cc_274 N_A_c_200_p N_X_c_971_n 0.0144259f $X=3.765 $Y=1.105 $X2=0 $Y2=0
cc_275 N_A_c_160_n N_X_c_971_n 0.0150081f $X=4.39 $Y=1.562 $X2=0 $Y2=0
cc_276 N_A_M1021_g N_X_c_1004_n 0.00311332f $X=5.765 $Y=2.4 $X2=0 $Y2=0
cc_277 N_A_M1026_g N_X_c_1004_n 0.00473876f $X=6.345 $Y=2.4 $X2=0 $Y2=0
cc_278 N_A_M1026_g N_X_c_978_n 0.00837972f $X=6.345 $Y=2.4 $X2=0 $Y2=0
cc_279 N_A_M1021_g N_X_c_1007_n 6.65006e-19 $X=5.765 $Y=2.4 $X2=0 $Y2=0
cc_280 N_A_M1026_g N_X_c_1007_n 0.00332621f $X=6.345 $Y=2.4 $X2=0 $Y2=0
cc_281 N_A_M1027_g N_X_c_1009_n 7.61432e-19 $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_282 N_A_c_175_p N_X_c_975_n 0.0144777f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_283 N_A_c_178_p N_X_c_975_n 0.00607737f $X=2.955 $Y=1.02 $X2=0 $Y2=0
cc_284 N_A_c_200_p N_X_c_975_n 0.0208829f $X=3.765 $Y=1.105 $X2=0 $Y2=0
cc_285 N_A_M1003_g N_X_c_1013_n 7.68112e-19 $X=4.725 $Y=2.4 $X2=0 $Y2=0
cc_286 N_A_c_153_n N_VGND_M1001_s 0.00510428f $X=0.6 $Y=1.42 $X2=-0.19
+ $Y2=-0.245
cc_287 N_A_c_318_p N_VGND_M1001_s 0.00321586f $X=0.685 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_288 N_A_c_175_p N_VGND_M1022_s 0.00394843f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_289 N_A_c_176_p N_VGND_M1022_s 0.00392577f $X=1.445 $Y=0.675 $X2=0 $Y2=0
cc_290 N_A_c_175_p N_VGND_M1028_s 0.00765915f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_291 N_A_c_200_p N_VGND_M1029_d 0.00594424f $X=3.765 $Y=1.105 $X2=0 $Y2=0
cc_292 N_A_c_155_n N_VGND_M1029_d 0.0021153f $X=3.85 $Y=1.35 $X2=0 $Y2=0
cc_293 N_A_M1001_g N_VGND_c_1133_n 0.0103672f $X=0.725 $Y=0.86 $X2=0 $Y2=0
cc_294 N_A_c_153_n N_VGND_c_1133_n 0.0374154f $X=0.6 $Y=1.42 $X2=0 $Y2=0
cc_295 N_A_c_318_p N_VGND_c_1133_n 0.0141996f $X=0.685 $Y=0.665 $X2=0 $Y2=0
cc_296 N_A_c_175_p N_VGND_c_1134_n 0.0247182f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_297 N_A_M1015_g N_VGND_c_1135_n 0.00348294f $X=4.745 $Y=0.74 $X2=0 $Y2=0
cc_298 N_A_M1015_g N_VGND_c_1136_n 0.00416335f $X=4.745 $Y=0.74 $X2=0 $Y2=0
cc_299 N_A_M1016_g N_VGND_c_1136_n 0.00418252f $X=5.335 $Y=0.74 $X2=0 $Y2=0
cc_300 N_A_M1025_g N_VGND_c_1137_n 0.00418252f $X=5.765 $Y=0.74 $X2=0 $Y2=0
cc_301 N_A_M1027_g N_VGND_c_1137_n 0.00231005f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_302 N_A_M1022_g N_VGND_c_1138_n 0.0014541f $X=1.155 $Y=0.86 $X2=0 $Y2=0
cc_303 N_A_c_175_p N_VGND_c_1138_n 0.0114916f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_304 N_A_c_176_p N_VGND_c_1138_n 0.0119842f $X=1.445 $Y=0.675 $X2=0 $Y2=0
cc_305 N_A_M1001_g N_VGND_c_1139_n 0.00374701f $X=0.725 $Y=0.86 $X2=0 $Y2=0
cc_306 N_A_M1022_g N_VGND_c_1139_n 0.00374721f $X=1.155 $Y=0.86 $X2=0 $Y2=0
cc_307 N_A_c_318_p N_VGND_c_1139_n 0.00306302f $X=0.685 $Y=0.665 $X2=0 $Y2=0
cc_308 N_A_c_204_p N_VGND_c_1139_n 0.0101323f $X=1.275 $Y=0.675 $X2=0 $Y2=0
cc_309 N_A_c_175_p N_VGND_c_1140_n 0.00464991f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_310 N_A_c_175_p N_VGND_c_1142_n 0.0129334f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_311 N_A_M1015_g N_VGND_c_1143_n 0.00324657f $X=4.745 $Y=0.74 $X2=0 $Y2=0
cc_312 N_A_M1016_g N_VGND_c_1144_n 0.00323547f $X=5.335 $Y=0.74 $X2=0 $Y2=0
cc_313 N_A_M1025_g N_VGND_c_1144_n 0.00323547f $X=5.765 $Y=0.74 $X2=0 $Y2=0
cc_314 N_A_M1027_g N_VGND_c_1145_n 0.00321293f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_315 N_A_M1001_g N_VGND_c_1146_n 0.00508379f $X=0.725 $Y=0.86 $X2=0 $Y2=0
cc_316 N_A_M1022_g N_VGND_c_1146_n 0.00508379f $X=1.155 $Y=0.86 $X2=0 $Y2=0
cc_317 N_A_M1015_g N_VGND_c_1146_n 0.00416139f $X=4.745 $Y=0.74 $X2=0 $Y2=0
cc_318 N_A_M1016_g N_VGND_c_1146_n 0.00412104f $X=5.335 $Y=0.74 $X2=0 $Y2=0
cc_319 N_A_M1025_g N_VGND_c_1146_n 0.00412104f $X=5.765 $Y=0.74 $X2=0 $Y2=0
cc_320 N_A_M1027_g N_VGND_c_1146_n 0.0041125f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_321 N_A_c_318_p N_VGND_c_1146_n 0.00533032f $X=0.685 $Y=0.665 $X2=0 $Y2=0
cc_322 N_A_c_175_p N_VGND_c_1146_n 0.0344715f $X=2.87 $Y=0.685 $X2=0 $Y2=0
cc_323 N_A_c_204_p N_VGND_c_1146_n 0.0176507f $X=1.275 $Y=0.675 $X2=0 $Y2=0
cc_324 N_A_c_176_p N_VGND_c_1146_n 7.98341e-19 $X=1.445 $Y=0.675 $X2=0 $Y2=0
cc_325 N_A_M1025_g N_A_877_74#_c_1261_n 0.00927675f $X=5.765 $Y=0.74 $X2=0 $Y2=0
cc_326 N_A_M1027_g N_A_877_74#_c_1261_n 0.00927675f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_327 N_A_M1025_g N_A_877_74#_c_1263_n 7.8287e-19 $X=5.765 $Y=0.74 $X2=0 $Y2=0
cc_328 N_A_M1027_g N_A_877_74#_c_1263_n 0.00539834f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_329 N_A_M1027_g N_A_877_74#_c_1255_n 0.0039285f $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_330 N_A_M1015_g N_A_877_74#_c_1258_n 0.00838898f $X=4.745 $Y=0.74 $X2=0 $Y2=0
cc_331 N_A_M1016_g N_A_877_74#_c_1258_n 7.98198e-19 $X=5.335 $Y=0.74 $X2=0 $Y2=0
cc_332 N_A_M1015_g N_A_877_74#_c_1268_n 0.00927675f $X=4.745 $Y=0.74 $X2=0 $Y2=0
cc_333 N_A_M1016_g N_A_877_74#_c_1268_n 0.00927675f $X=5.335 $Y=0.74 $X2=0 $Y2=0
cc_334 N_A_M1015_g N_A_877_74#_c_1259_n 7.98516e-19 $X=4.745 $Y=0.74 $X2=0 $Y2=0
cc_335 N_A_M1016_g N_A_877_74#_c_1259_n 0.00763599f $X=5.335 $Y=0.74 $X2=0 $Y2=0
cc_336 N_A_M1025_g N_A_877_74#_c_1259_n 0.00763599f $X=5.765 $Y=0.74 $X2=0 $Y2=0
cc_337 N_A_M1027_g N_A_877_74#_c_1259_n 7.98516e-19 $X=6.355 $Y=0.74 $X2=0 $Y2=0
cc_338 N_B_M1028_g N_A_160_98#_c_568_n 0.0239678f $X=2.285 $Y=0.86 $X2=0 $Y2=0
cc_339 N_B_c_380_n N_A_160_98#_M1013_g 0.00103996f $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_340 N_B_c_381_n N_A_160_98#_M1013_g 0.00491551f $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_341 N_B_c_392_n N_A_160_98#_M1013_g 0.0183584f $X=3.485 $Y=1.935 $X2=0 $Y2=0
cc_342 N_B_c_392_n N_A_160_98#_M1017_g 0.0108123f $X=3.485 $Y=1.935 $X2=0 $Y2=0
cc_343 N_B_c_407_n N_A_160_98#_M1018_g 0.0123863f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_344 N_B_c_422_n N_A_160_98#_M1018_g 0.00248464f $X=3.57 $Y=1.935 $X2=0 $Y2=0
cc_345 N_B_c_407_n N_A_160_98#_c_570_n 5.02183e-19 $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_346 N_B_M1028_g N_A_160_98#_c_571_n 0.0193036f $X=2.285 $Y=0.86 $X2=0 $Y2=0
cc_347 N_B_c_380_n N_A_160_98#_c_571_n 2.34086e-19 $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_348 N_B_c_392_n N_A_160_98#_c_571_n 0.00586816f $X=3.485 $Y=1.935 $X2=0 $Y2=0
cc_349 N_B_c_422_n N_A_160_98#_c_571_n 0.00266507f $X=3.57 $Y=1.935 $X2=0 $Y2=0
cc_350 N_B_c_407_n N_A_160_98#_M1019_g 0.0115787f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_351 N_B_c_381_n N_A_160_98#_c_600_n 0.00539411f $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_352 N_B_c_384_n N_A_160_98#_c_572_n 0.0115982f $X=1.5 $Y=1.9 $X2=0 $Y2=0
cc_353 N_B_M1023_g N_A_160_98#_c_572_n 0.0104353f $X=1.745 $Y=0.86 $X2=0 $Y2=0
cc_354 N_B_M1028_g N_A_160_98#_c_572_n 0.00149841f $X=2.285 $Y=0.86 $X2=0 $Y2=0
cc_355 N_B_c_380_n N_A_160_98#_c_572_n 0.0229023f $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_356 N_B_c_381_n N_A_160_98#_c_572_n 0.0265559f $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_357 N_B_c_393_n N_A_160_98#_c_572_n 0.00946087f $X=2.36 $Y=1.935 $X2=0 $Y2=0
cc_358 N_B_M1023_g N_A_160_98#_c_608_n 6.6817e-19 $X=1.745 $Y=0.86 $X2=0 $Y2=0
cc_359 N_B_M1028_g N_A_160_98#_c_608_n 0.0117669f $X=2.285 $Y=0.86 $X2=0 $Y2=0
cc_360 N_B_c_380_n N_A_160_98#_c_608_n 0.0158037f $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_361 N_B_c_381_n N_A_160_98#_c_608_n 0.00522409f $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_362 N_B_c_392_n N_A_160_98#_c_608_n 0.00402169f $X=3.485 $Y=1.935 $X2=0 $Y2=0
cc_363 N_B_M1028_g N_A_160_98#_c_573_n 0.0037313f $X=2.285 $Y=0.86 $X2=0 $Y2=0
cc_364 N_B_M1028_g N_A_160_98#_c_574_n 0.0044251f $X=2.285 $Y=0.86 $X2=0 $Y2=0
cc_365 N_B_c_380_n N_A_160_98#_c_574_n 0.01771f $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_366 N_B_c_392_n N_A_160_98#_c_574_n 0.0136221f $X=3.485 $Y=1.935 $X2=0 $Y2=0
cc_367 N_B_c_392_n N_A_160_98#_c_611_n 0.0499776f $X=3.485 $Y=1.935 $X2=0 $Y2=0
cc_368 N_B_c_422_n N_A_160_98#_c_611_n 0.00693899f $X=3.57 $Y=1.935 $X2=0 $Y2=0
cc_369 N_B_M1023_g N_A_160_98#_c_620_n 0.0093952f $X=1.745 $Y=0.86 $X2=0 $Y2=0
cc_370 N_B_c_393_n N_A_36_392#_M1011_s 0.00223196f $X=2.36 $Y=1.935 $X2=0 $Y2=0
cc_371 N_B_c_384_n N_A_36_392#_c_699_n 3.48606e-19 $X=1.5 $Y=1.9 $X2=0 $Y2=0
cc_372 N_B_c_384_n N_A_36_392#_c_701_n 0.0139961f $X=1.5 $Y=1.9 $X2=0 $Y2=0
cc_373 N_B_c_385_n N_A_36_392#_c_701_n 0.014552f $X=1.95 $Y=1.845 $X2=0 $Y2=0
cc_374 N_B_c_384_n N_A_36_392#_c_703_n 6.51491e-19 $X=1.5 $Y=1.9 $X2=0 $Y2=0
cc_375 N_B_c_385_n N_A_36_392#_c_703_n 0.0124236f $X=1.95 $Y=1.845 $X2=0 $Y2=0
cc_376 N_B_c_381_n N_A_36_392#_c_703_n 0.00143058f $X=2.195 $Y=1.635 $X2=0 $Y2=0
cc_377 N_B_c_393_n N_A_36_392#_c_703_n 0.0223657f $X=2.36 $Y=1.935 $X2=0 $Y2=0
cc_378 N_B_c_407_n N_VPWR_M1003_s 0.00631727f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_379 N_B_c_407_n N_VPWR_M1021_s 0.00225758f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_380 N_B_c_394_n N_VPWR_M1021_s 0.00131423f $X=5.89 $Y=1.945 $X2=0 $Y2=0
cc_381 N_B_M1000_g N_VPWR_c_743_n 0.00847535f $X=6.795 $Y=2.4 $X2=0 $Y2=0
cc_382 N_B_M1002_g N_VPWR_c_743_n 0.002979f $X=7.245 $Y=2.4 $X2=0 $Y2=0
cc_383 N_B_M1005_g N_VPWR_c_744_n 0.0027763f $X=7.695 $Y=2.4 $X2=0 $Y2=0
cc_384 N_B_M1008_g N_VPWR_c_744_n 0.0027763f $X=8.145 $Y=2.4 $X2=0 $Y2=0
cc_385 N_B_c_384_n N_VPWR_c_745_n 0.00333926f $X=1.5 $Y=1.9 $X2=0 $Y2=0
cc_386 N_B_c_385_n N_VPWR_c_745_n 0.00333896f $X=1.95 $Y=1.845 $X2=0 $Y2=0
cc_387 N_B_M1000_g N_VPWR_c_747_n 0.00460063f $X=6.795 $Y=2.4 $X2=0 $Y2=0
cc_388 N_B_M1002_g N_VPWR_c_748_n 0.005209f $X=7.245 $Y=2.4 $X2=0 $Y2=0
cc_389 N_B_M1005_g N_VPWR_c_748_n 0.005209f $X=7.695 $Y=2.4 $X2=0 $Y2=0
cc_390 N_B_M1008_g N_VPWR_c_749_n 0.005209f $X=8.145 $Y=2.4 $X2=0 $Y2=0
cc_391 N_B_c_384_n N_VPWR_c_741_n 0.00422798f $X=1.5 $Y=1.9 $X2=0 $Y2=0
cc_392 N_B_c_385_n N_VPWR_c_741_n 0.00427818f $X=1.95 $Y=1.845 $X2=0 $Y2=0
cc_393 N_B_M1000_g N_VPWR_c_741_n 0.00908665f $X=6.795 $Y=2.4 $X2=0 $Y2=0
cc_394 N_B_M1002_g N_VPWR_c_741_n 0.00982266f $X=7.245 $Y=2.4 $X2=0 $Y2=0
cc_395 N_B_M1005_g N_VPWR_c_741_n 0.00982266f $X=7.695 $Y=2.4 $X2=0 $Y2=0
cc_396 N_B_M1008_g N_VPWR_c_741_n 0.00985972f $X=8.145 $Y=2.4 $X2=0 $Y2=0
cc_397 N_B_c_392_n N_A_514_368#_M1013_s 0.00473172f $X=3.485 $Y=1.935 $X2=-0.19
+ $Y2=-0.245
cc_398 N_B_c_407_n N_A_514_368#_M1017_s 0.00153118f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_399 N_B_c_422_n N_A_514_368#_M1017_s 0.0045141f $X=3.57 $Y=1.935 $X2=0 $Y2=0
cc_400 N_B_c_407_n N_A_514_368#_M1019_s 0.00332471f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_401 N_B_c_407_n N_A_514_368#_M1006_d 0.00314624f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_402 N_B_c_385_n N_A_514_368#_c_858_n 0.00123081f $X=1.95 $Y=1.845 $X2=0 $Y2=0
cc_403 N_B_c_392_n N_A_514_368#_c_858_n 0.0197942f $X=3.485 $Y=1.935 $X2=0 $Y2=0
cc_404 N_B_c_385_n N_A_514_368#_c_860_n 5.90446e-19 $X=1.95 $Y=1.845 $X2=0 $Y2=0
cc_405 N_B_M1000_g N_A_514_368#_c_887_n 0.0140196f $X=6.795 $Y=2.4 $X2=0 $Y2=0
cc_406 N_B_M1002_g N_A_514_368#_c_887_n 0.0126573f $X=7.245 $Y=2.4 $X2=0 $Y2=0
cc_407 N_B_M1005_g N_A_514_368#_c_889_n 0.012696f $X=7.695 $Y=2.4 $X2=0 $Y2=0
cc_408 N_B_M1008_g N_A_514_368#_c_889_n 0.012696f $X=8.145 $Y=2.4 $X2=0 $Y2=0
cc_409 N_B_M1000_g N_A_514_368#_c_866_n 5.87938e-19 $X=6.795 $Y=2.4 $X2=0 $Y2=0
cc_410 N_B_M1002_g N_A_514_368#_c_866_n 0.00896953f $X=7.245 $Y=2.4 $X2=0 $Y2=0
cc_411 N_B_M1005_g N_A_514_368#_c_866_n 0.00877121f $X=7.695 $Y=2.4 $X2=0 $Y2=0
cc_412 N_B_M1008_g N_A_514_368#_c_866_n 5.64228e-19 $X=8.145 $Y=2.4 $X2=0 $Y2=0
cc_413 N_B_M1005_g N_A_514_368#_c_867_n 5.64228e-19 $X=7.695 $Y=2.4 $X2=0 $Y2=0
cc_414 N_B_M1008_g N_A_514_368#_c_867_n 0.00893344f $X=8.145 $Y=2.4 $X2=0 $Y2=0
cc_415 N_B_c_392_n N_X_M1013_d 0.00311483f $X=3.485 $Y=1.935 $X2=0 $Y2=0
cc_416 N_B_c_407_n N_X_M1018_d 0.00314279f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_417 N_B_c_407_n N_X_c_987_n 0.00883092f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_418 N_B_c_383_n N_X_c_987_n 0.00618698f $X=8 $Y=1.515 $X2=0 $Y2=0
cc_419 N_B_M1010_g N_X_c_970_n 0.00895879f $X=6.785 $Y=0.74 $X2=0 $Y2=0
cc_420 N_B_c_382_n N_X_c_970_n 0.010549f $X=5.89 $Y=1.78 $X2=0 $Y2=0
cc_421 N_B_c_383_n N_X_c_970_n 0.065983f $X=8 $Y=1.515 $X2=0 $Y2=0
cc_422 N_B_M1000_g N_X_c_1004_n 7.76868e-19 $X=6.795 $Y=2.4 $X2=0 $Y2=0
cc_423 N_B_M1000_g N_X_c_978_n 0.0116248f $X=6.795 $Y=2.4 $X2=0 $Y2=0
cc_424 N_B_M1002_g N_X_c_978_n 0.0116623f $X=7.245 $Y=2.4 $X2=0 $Y2=0
cc_425 N_B_M1005_g N_X_c_978_n 0.0116623f $X=7.695 $Y=2.4 $X2=0 $Y2=0
cc_426 N_B_M1008_g N_X_c_978_n 0.0151299f $X=8.145 $Y=2.4 $X2=0 $Y2=0
cc_427 N_B_c_378_n N_X_c_978_n 9.81182e-19 $X=8.145 $Y=1.35 $X2=0 $Y2=0
cc_428 N_B_c_383_n N_X_c_978_n 0.125611f $X=8 $Y=1.515 $X2=0 $Y2=0
cc_429 N_B_c_407_n N_X_c_1007_n 0.0148765f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_430 N_B_c_383_n N_X_c_1007_n 0.0118338f $X=8 $Y=1.515 $X2=0 $Y2=0
cc_431 N_B_M1010_g N_X_c_1009_n 0.00659181f $X=6.785 $Y=0.74 $X2=0 $Y2=0
cc_432 N_B_c_374_n N_X_c_1009_n 5.72926e-19 $X=7.14 $Y=0.22 $X2=0 $Y2=0
cc_433 N_B_M1012_g N_X_c_1009_n 0.00674159f $X=7.215 $Y=0.74 $X2=0 $Y2=0
cc_434 N_B_M1020_g N_X_c_1009_n 7.30686e-19 $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_435 N_B_M1012_g N_X_c_972_n 0.0093986f $X=7.215 $Y=0.74 $X2=0 $Y2=0
cc_436 N_B_M1020_g N_X_c_972_n 0.0124803f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_437 N_B_c_378_n N_X_c_972_n 0.00895685f $X=8.145 $Y=1.35 $X2=0 $Y2=0
cc_438 N_B_c_383_n N_X_c_972_n 0.0510605f $X=8 $Y=1.515 $X2=0 $Y2=0
cc_439 N_B_c_378_n N_X_c_973_n 6.22593e-19 $X=8.145 $Y=1.35 $X2=0 $Y2=0
cc_440 N_B_M1024_g N_X_c_973_n 0.0151483f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_441 N_B_c_383_n N_X_c_973_n 0.0111136f $X=8 $Y=1.515 $X2=0 $Y2=0
cc_442 N_B_c_378_n N_X_c_974_n 0.0179941f $X=8.145 $Y=1.35 $X2=0 $Y2=0
cc_443 N_B_M1024_g N_X_c_974_n 0.00614193f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_444 N_B_c_383_n N_X_c_974_n 0.034159f $X=8 $Y=1.515 $X2=0 $Y2=0
cc_445 N_B_c_392_n N_X_c_1044_n 0.0167216f $X=3.485 $Y=1.935 $X2=0 $Y2=0
cc_446 N_B_c_371_n N_X_c_976_n 8.27088e-19 $X=6.795 $Y=1.275 $X2=0 $Y2=0
cc_447 N_B_M1010_g N_X_c_976_n 0.00277633f $X=6.785 $Y=0.74 $X2=0 $Y2=0
cc_448 N_B_M1012_g N_X_c_976_n 0.00269795f $X=7.215 $Y=0.74 $X2=0 $Y2=0
cc_449 N_B_c_383_n N_X_c_976_n 0.0289344f $X=8 $Y=1.515 $X2=0 $Y2=0
cc_450 N_B_c_378_n N_X_c_977_n 0.00237463f $X=8.145 $Y=1.35 $X2=0 $Y2=0
cc_451 N_B_c_383_n N_X_c_977_n 0.0144276f $X=8 $Y=1.515 $X2=0 $Y2=0
cc_452 N_B_c_392_n N_X_c_1051_n 0.00713119f $X=3.485 $Y=1.935 $X2=0 $Y2=0
cc_453 N_B_c_407_n N_X_c_1051_n 0.115888f $X=5.805 $Y=2.03 $X2=0 $Y2=0
cc_454 N_B_c_422_n N_X_c_1051_n 0.00996656f $X=3.57 $Y=1.935 $X2=0 $Y2=0
cc_455 N_B_M1028_g N_VGND_c_1134_n 0.00203574f $X=2.285 $Y=0.86 $X2=0 $Y2=0
cc_456 N_B_c_375_n N_VGND_c_1137_n 0.00170967f $X=6.86 $Y=0.22 $X2=0 $Y2=0
cc_457 N_B_M1023_g N_VGND_c_1138_n 0.0014541f $X=1.745 $Y=0.86 $X2=0 $Y2=0
cc_458 N_B_M1023_g N_VGND_c_1142_n 0.00376411f $X=1.745 $Y=0.86 $X2=0 $Y2=0
cc_459 N_B_M1028_g N_VGND_c_1142_n 0.00376411f $X=2.285 $Y=0.86 $X2=0 $Y2=0
cc_460 N_B_c_375_n N_VGND_c_1145_n 0.0124522f $X=6.86 $Y=0.22 $X2=0 $Y2=0
cc_461 N_B_M1020_g N_VGND_c_1145_n 0.00278247f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_462 N_B_M1024_g N_VGND_c_1145_n 0.00278247f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_463 N_B_M1023_g N_VGND_c_1146_n 0.00508379f $X=1.745 $Y=0.86 $X2=0 $Y2=0
cc_464 N_B_M1028_g N_VGND_c_1146_n 0.00508379f $X=2.285 $Y=0.86 $X2=0 $Y2=0
cc_465 N_B_c_374_n N_VGND_c_1146_n 0.0121953f $X=7.14 $Y=0.22 $X2=0 $Y2=0
cc_466 N_B_c_375_n N_VGND_c_1146_n 0.00536641f $X=6.86 $Y=0.22 $X2=0 $Y2=0
cc_467 N_B_M1020_g N_VGND_c_1146_n 0.00354085f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_468 N_B_M1024_g N_VGND_c_1146_n 0.00357084f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_469 N_B_M1010_g N_A_877_74#_c_1254_n 0.00852441f $X=6.785 $Y=0.74 $X2=0 $Y2=0
cc_470 N_B_c_374_n N_A_877_74#_c_1254_n 0.00709642f $X=7.14 $Y=0.22 $X2=0 $Y2=0
cc_471 N_B_c_375_n N_A_877_74#_c_1254_n 0.00216415f $X=6.86 $Y=0.22 $X2=0 $Y2=0
cc_472 N_B_M1012_g N_A_877_74#_c_1254_n 0.0088595f $X=7.215 $Y=0.74 $X2=0 $Y2=0
cc_473 N_B_M1020_g N_A_877_74#_c_1278_n 0.00646522f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_474 N_B_M1024_g N_A_877_74#_c_1278_n 5.7278e-19 $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_475 N_B_M1020_g N_A_877_74#_c_1256_n 0.00792642f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_476 N_B_M1024_g N_A_877_74#_c_1256_n 0.0118796f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_477 N_B_M1020_g N_A_877_74#_c_1257_n 5.7278e-19 $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_478 N_B_M1024_g N_A_877_74#_c_1257_n 0.00690717f $X=8.145 $Y=0.74 $X2=0 $Y2=0
cc_479 N_B_M1020_g N_A_877_74#_c_1260_n 0.00294698f $X=7.715 $Y=0.74 $X2=0 $Y2=0
cc_480 N_A_160_98#_c_572_n N_A_36_392#_c_699_n 0.00700951f $X=1.725 $Y=2.105
+ $X2=0 $Y2=0
cc_481 N_A_160_98#_M1007_d N_A_36_392#_c_701_n 0.00165831f $X=1.59 $Y=1.96 $X2=0
+ $Y2=0
cc_482 N_A_160_98#_M1013_g N_A_36_392#_c_701_n 5.84324e-19 $X=2.925 $Y=2.4 $X2=0
+ $Y2=0
cc_483 N_A_160_98#_c_572_n N_A_36_392#_c_701_n 0.0139027f $X=1.725 $Y=2.105
+ $X2=0 $Y2=0
cc_484 N_A_160_98#_M1013_g N_VPWR_c_745_n 0.00333926f $X=2.925 $Y=2.4 $X2=0
+ $Y2=0
cc_485 N_A_160_98#_M1017_g N_VPWR_c_745_n 0.00333926f $X=3.375 $Y=2.4 $X2=0
+ $Y2=0
cc_486 N_A_160_98#_M1018_g N_VPWR_c_745_n 0.00333926f $X=3.825 $Y=2.4 $X2=0
+ $Y2=0
cc_487 N_A_160_98#_M1019_g N_VPWR_c_745_n 0.00333926f $X=4.275 $Y=2.4 $X2=0
+ $Y2=0
cc_488 N_A_160_98#_M1013_g N_VPWR_c_741_n 0.0042782f $X=2.925 $Y=2.4 $X2=0 $Y2=0
cc_489 N_A_160_98#_M1017_g N_VPWR_c_741_n 0.00422687f $X=3.375 $Y=2.4 $X2=0
+ $Y2=0
cc_490 N_A_160_98#_M1018_g N_VPWR_c_741_n 0.00422687f $X=3.825 $Y=2.4 $X2=0
+ $Y2=0
cc_491 N_A_160_98#_M1019_g N_VPWR_c_741_n 0.00422798f $X=4.275 $Y=2.4 $X2=0
+ $Y2=0
cc_492 N_A_160_98#_M1013_g N_A_514_368#_c_859_n 0.0149887f $X=2.925 $Y=2.4 $X2=0
+ $Y2=0
cc_493 N_A_160_98#_M1017_g N_A_514_368#_c_859_n 0.0108701f $X=3.375 $Y=2.4 $X2=0
+ $Y2=0
cc_494 N_A_160_98#_M1018_g N_A_514_368#_c_861_n 0.0108462f $X=3.825 $Y=2.4 $X2=0
+ $Y2=0
cc_495 N_A_160_98#_M1019_g N_A_514_368#_c_861_n 0.01005f $X=4.275 $Y=2.4 $X2=0
+ $Y2=0
cc_496 N_A_160_98#_M1019_g N_A_514_368#_c_864_n 2.29065e-19 $X=4.275 $Y=2.4
+ $X2=0 $Y2=0
cc_497 N_A_160_98#_c_569_n N_X_c_968_n 0.0108146f $X=3.59 $Y=1.35 $X2=0 $Y2=0
cc_498 N_A_160_98#_c_570_n N_X_c_968_n 5.69335e-19 $X=4.185 $Y=1.605 $X2=0 $Y2=0
cc_499 N_A_160_98#_c_569_n N_X_c_969_n 0.00409433f $X=3.59 $Y=1.35 $X2=0 $Y2=0
cc_500 N_A_160_98#_M1019_g N_X_c_987_n 0.00978447f $X=4.275 $Y=2.4 $X2=0 $Y2=0
cc_501 N_A_160_98#_c_570_n N_X_c_970_n 4.05724e-19 $X=4.185 $Y=1.605 $X2=0 $Y2=0
cc_502 N_A_160_98#_c_569_n N_X_c_971_n 0.00102704f $X=3.59 $Y=1.35 $X2=0 $Y2=0
cc_503 N_A_160_98#_c_570_n N_X_c_971_n 8.40444e-19 $X=4.185 $Y=1.605 $X2=0 $Y2=0
cc_504 N_A_160_98#_M1013_g N_X_c_1044_n 0.00762274f $X=2.925 $Y=2.4 $X2=0 $Y2=0
cc_505 N_A_160_98#_M1017_g N_X_c_1044_n 0.00813468f $X=3.375 $Y=2.4 $X2=0 $Y2=0
cc_506 N_A_160_98#_M1018_g N_X_c_1044_n 0.00102153f $X=3.825 $Y=2.4 $X2=0 $Y2=0
cc_507 N_A_160_98#_c_568_n N_X_c_975_n 0.00391079f $X=2.875 $Y=1.35 $X2=0 $Y2=0
cc_508 N_A_160_98#_c_569_n N_X_c_975_n 0.00967015f $X=3.59 $Y=1.35 $X2=0 $Y2=0
cc_509 N_A_160_98#_M1017_g N_X_c_1051_n 0.0114028f $X=3.375 $Y=2.4 $X2=0 $Y2=0
cc_510 N_A_160_98#_M1018_g N_X_c_1051_n 0.00982318f $X=3.825 $Y=2.4 $X2=0 $Y2=0
cc_511 N_A_160_98#_M1017_g N_X_c_1013_n 4.89439e-19 $X=3.375 $Y=2.4 $X2=0 $Y2=0
cc_512 N_A_160_98#_M1018_g N_X_c_1013_n 0.00655324f $X=3.825 $Y=2.4 $X2=0 $Y2=0
cc_513 N_A_160_98#_M1019_g N_X_c_1013_n 0.00653767f $X=4.275 $Y=2.4 $X2=0 $Y2=0
cc_514 N_A_160_98#_c_600_n N_VGND_M1022_s 0.0110596f $X=1.56 $Y=1.065 $X2=0
+ $Y2=0
cc_515 N_A_160_98#_c_572_n N_VGND_M1022_s 4.81637e-19 $X=1.725 $Y=2.105 $X2=0
+ $Y2=0
cc_516 N_A_160_98#_c_620_n N_VGND_M1022_s 5.87954e-19 $X=1.685 $Y=1.065 $X2=0
+ $Y2=0
cc_517 N_A_160_98#_c_608_n N_VGND_M1028_s 0.00947801f $X=2.53 $Y=1.065 $X2=0
+ $Y2=0
cc_518 N_A_160_98#_c_573_n N_VGND_M1028_s 8.87448e-19 $X=2.615 $Y=1.36 $X2=0
+ $Y2=0
cc_519 N_A_160_98#_c_568_n N_VGND_c_1134_n 0.00203574f $X=2.875 $Y=1.35 $X2=0
+ $Y2=0
cc_520 N_A_160_98#_c_569_n N_VGND_c_1135_n 0.00559625f $X=3.59 $Y=1.35 $X2=0
+ $Y2=0
cc_521 N_A_160_98#_c_568_n N_VGND_c_1140_n 0.00376367f $X=2.875 $Y=1.35 $X2=0
+ $Y2=0
cc_522 N_A_160_98#_c_569_n N_VGND_c_1140_n 0.00380789f $X=3.59 $Y=1.35 $X2=0
+ $Y2=0
cc_523 N_A_160_98#_c_568_n N_VGND_c_1146_n 0.00508379f $X=2.875 $Y=1.35 $X2=0
+ $Y2=0
cc_524 N_A_160_98#_c_569_n N_VGND_c_1146_n 0.00508379f $X=3.59 $Y=1.35 $X2=0
+ $Y2=0
cc_525 N_A_36_392#_c_699_n N_VPWR_M1004_s 0.00218982f $X=1.11 $Y=2.005 $X2=-0.19
+ $Y2=1.66
cc_526 N_A_36_392#_c_698_n N_VPWR_c_742_n 0.0243967f $X=0.325 $Y=2.105 $X2=0
+ $Y2=0
cc_527 N_A_36_392#_c_699_n N_VPWR_c_742_n 0.0167599f $X=1.11 $Y=2.005 $X2=0
+ $Y2=0
cc_528 N_A_36_392#_c_702_n N_VPWR_c_742_n 0.0117278f $X=1.36 $Y=2.99 $X2=0 $Y2=0
cc_529 N_A_36_392#_c_701_n N_VPWR_c_745_n 0.0644071f $X=2.01 $Y=2.99 $X2=0 $Y2=0
cc_530 N_A_36_392#_c_702_n N_VPWR_c_745_n 0.0178163f $X=1.36 $Y=2.99 $X2=0 $Y2=0
cc_531 N_A_36_392#_c_698_n N_VPWR_c_741_n 0.0119743f $X=0.325 $Y=2.105 $X2=0
+ $Y2=0
cc_532 N_A_36_392#_c_701_n N_VPWR_c_741_n 0.0356218f $X=2.01 $Y=2.99 $X2=0 $Y2=0
cc_533 N_A_36_392#_c_702_n N_VPWR_c_741_n 0.00958215f $X=1.36 $Y=2.99 $X2=0
+ $Y2=0
cc_534 N_A_36_392#_c_698_n N_VPWR_c_751_n 0.014549f $X=0.325 $Y=2.105 $X2=0
+ $Y2=0
cc_535 N_A_36_392#_c_703_n N_A_514_368#_c_858_n 0.0528782f $X=2.175 $Y=2.355
+ $X2=0 $Y2=0
cc_536 N_A_36_392#_c_701_n N_A_514_368#_c_860_n 0.0144477f $X=2.01 $Y=2.99 $X2=0
+ $Y2=0
cc_537 N_A_36_392#_c_700_n N_VGND_c_1133_n 0.00657381f $X=0.49 $Y=2.005 $X2=0
+ $Y2=0
cc_538 N_VPWR_c_745_n N_A_514_368#_c_859_n 0.0459191f $X=4.855 $Y=3.33 $X2=0
+ $Y2=0
cc_539 N_VPWR_c_741_n N_A_514_368#_c_859_n 0.0258001f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_540 N_VPWR_c_745_n N_A_514_368#_c_860_n 0.0179217f $X=4.855 $Y=3.33 $X2=0
+ $Y2=0
cc_541 N_VPWR_c_741_n N_A_514_368#_c_860_n 0.00971942f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_542 N_VPWR_c_745_n N_A_514_368#_c_861_n 0.0459483f $X=4.855 $Y=3.33 $X2=0
+ $Y2=0
cc_543 N_VPWR_c_741_n N_A_514_368#_c_861_n 0.0258042f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_544 N_VPWR_M1021_s N_A_514_368#_c_868_n 0.00626389f $X=5.855 $Y=1.84 $X2=0
+ $Y2=0
cc_545 N_VPWR_c_746_n N_A_514_368#_c_868_n 0.00253855f $X=5.89 $Y=3.33 $X2=0
+ $Y2=0
cc_546 N_VPWR_c_747_n N_A_514_368#_c_868_n 0.00420254f $X=6.855 $Y=3.33 $X2=0
+ $Y2=0
cc_547 N_VPWR_c_741_n N_A_514_368#_c_868_n 0.0112876f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_548 N_VPWR_c_753_n N_A_514_368#_c_868_n 0.0229497f $X=6.055 $Y=3.05 $X2=0
+ $Y2=0
cc_549 N_VPWR_c_743_n N_A_514_368#_c_862_n 0.0117359f $X=7.02 $Y=2.805 $X2=0
+ $Y2=0
cc_550 N_VPWR_c_747_n N_A_514_368#_c_862_n 0.00759366f $X=6.855 $Y=3.33 $X2=0
+ $Y2=0
cc_551 N_VPWR_c_741_n N_A_514_368#_c_862_n 0.00628181f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_552 N_VPWR_c_753_n N_A_514_368#_c_862_n 8.74611e-19 $X=6.055 $Y=3.05 $X2=0
+ $Y2=0
cc_553 N_VPWR_M1000_d N_A_514_368#_c_887_n 0.00332066f $X=6.885 $Y=1.84 $X2=0
+ $Y2=0
cc_554 N_VPWR_c_743_n N_A_514_368#_c_887_n 0.0148589f $X=7.02 $Y=2.805 $X2=0
+ $Y2=0
cc_555 N_VPWR_M1005_d N_A_514_368#_c_889_n 0.00324075f $X=7.785 $Y=1.84 $X2=0
+ $Y2=0
cc_556 N_VPWR_c_744_n N_A_514_368#_c_889_n 0.0126919f $X=7.92 $Y=2.805 $X2=0
+ $Y2=0
cc_557 N_VPWR_c_745_n N_A_514_368#_c_863_n 0.0118207f $X=4.855 $Y=3.33 $X2=0
+ $Y2=0
cc_558 N_VPWR_c_741_n N_A_514_368#_c_863_n 0.00654074f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_559 N_VPWR_c_745_n N_A_514_368#_c_864_n 0.0171415f $X=4.855 $Y=3.33 $X2=0
+ $Y2=0
cc_560 N_VPWR_c_741_n N_A_514_368#_c_864_n 0.00940804f $X=8.4 $Y=3.33 $X2=0
+ $Y2=0
cc_561 N_VPWR_c_752_n N_A_514_368#_c_864_n 0.00784965f $X=5.02 $Y=3.05 $X2=0
+ $Y2=0
cc_562 N_VPWR_M1003_s N_A_514_368#_c_873_n 0.00657535f $X=4.815 $Y=1.84 $X2=0
+ $Y2=0
cc_563 N_VPWR_c_745_n N_A_514_368#_c_873_n 0.00364766f $X=4.855 $Y=3.33 $X2=0
+ $Y2=0
cc_564 N_VPWR_c_746_n N_A_514_368#_c_873_n 0.00363957f $X=5.89 $Y=3.33 $X2=0
+ $Y2=0
cc_565 N_VPWR_c_741_n N_A_514_368#_c_873_n 0.012114f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_566 N_VPWR_c_752_n N_A_514_368#_c_873_n 0.0232472f $X=5.02 $Y=3.05 $X2=0
+ $Y2=0
cc_567 N_VPWR_c_746_n N_A_514_368#_c_865_n 0.0138332f $X=5.89 $Y=3.33 $X2=0
+ $Y2=0
cc_568 N_VPWR_c_741_n N_A_514_368#_c_865_n 0.0116354f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_569 N_VPWR_c_752_n N_A_514_368#_c_865_n 0.00102354f $X=5.02 $Y=3.05 $X2=0
+ $Y2=0
cc_570 N_VPWR_c_753_n N_A_514_368#_c_865_n 0.0010443f $X=6.055 $Y=3.05 $X2=0
+ $Y2=0
cc_571 N_VPWR_c_743_n N_A_514_368#_c_866_n 0.0122069f $X=7.02 $Y=2.805 $X2=0
+ $Y2=0
cc_572 N_VPWR_c_744_n N_A_514_368#_c_866_n 0.0121684f $X=7.92 $Y=2.805 $X2=0
+ $Y2=0
cc_573 N_VPWR_c_748_n N_A_514_368#_c_866_n 0.0144776f $X=7.835 $Y=3.33 $X2=0
+ $Y2=0
cc_574 N_VPWR_c_741_n N_A_514_368#_c_866_n 0.0118404f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_575 N_VPWR_c_744_n N_A_514_368#_c_867_n 0.0121684f $X=7.92 $Y=2.805 $X2=0
+ $Y2=0
cc_576 N_VPWR_c_749_n N_A_514_368#_c_867_n 0.0145644f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_577 N_VPWR_c_741_n N_A_514_368#_c_867_n 0.0119803f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_578 N_VPWR_M1003_s N_X_c_987_n 0.00656633f $X=4.815 $Y=1.84 $X2=0 $Y2=0
cc_579 N_VPWR_M1021_s N_X_c_987_n 0.0068f $X=5.855 $Y=1.84 $X2=0 $Y2=0
cc_580 N_VPWR_M1021_s N_X_c_1004_n 0.00207781f $X=5.855 $Y=1.84 $X2=0 $Y2=0
cc_581 N_VPWR_M1000_d N_X_c_978_n 0.00332471f $X=6.885 $Y=1.84 $X2=0 $Y2=0
cc_582 N_VPWR_M1005_d N_X_c_978_n 0.0031478f $X=7.785 $Y=1.84 $X2=0 $Y2=0
cc_583 N_VPWR_M1021_s N_X_c_1007_n 0.0021229f $X=5.855 $Y=1.84 $X2=0 $Y2=0
cc_584 N_A_514_368#_c_859_n N_X_M1013_d 0.00165831f $X=3.515 $Y=2.99 $X2=0 $Y2=0
cc_585 N_A_514_368#_c_861_n N_X_M1018_d 0.00166235f $X=4.415 $Y=2.99 $X2=0 $Y2=0
cc_586 N_A_514_368#_M1019_s N_X_c_987_n 0.00332066f $X=4.365 $Y=1.84 $X2=0 $Y2=0
cc_587 N_A_514_368#_M1006_d N_X_c_987_n 0.0032437f $X=5.405 $Y=1.84 $X2=0 $Y2=0
cc_588 N_A_514_368#_c_861_n N_X_c_987_n 0.00458951f $X=4.415 $Y=2.99 $X2=0 $Y2=0
cc_589 N_A_514_368#_c_868_n N_X_c_987_n 0.00866795f $X=6.485 $Y=2.71 $X2=0 $Y2=0
cc_590 N_A_514_368#_c_864_n N_X_c_987_n 0.0143712f $X=4.54 $Y=2.71 $X2=0 $Y2=0
cc_591 N_A_514_368#_c_873_n N_X_c_987_n 0.0854383f $X=5.375 $Y=2.802 $X2=0 $Y2=0
cc_592 N_A_514_368#_M1026_d N_X_c_978_n 0.00332066f $X=6.435 $Y=1.84 $X2=0 $Y2=0
cc_593 N_A_514_368#_M1002_s N_X_c_978_n 0.00314376f $X=7.335 $Y=1.84 $X2=0 $Y2=0
cc_594 N_A_514_368#_M1008_s N_X_c_978_n 0.0124238f $X=8.235 $Y=1.84 $X2=0 $Y2=0
cc_595 N_A_514_368#_c_868_n N_X_c_978_n 0.00331783f $X=6.485 $Y=2.71 $X2=0 $Y2=0
cc_596 N_A_514_368#_c_956_p N_X_c_978_n 0.0127071f $X=6.57 $Y=2.46 $X2=0 $Y2=0
cc_597 N_A_514_368#_c_887_n N_X_c_978_n 0.0336305f $X=7.305 $Y=2.375 $X2=0 $Y2=0
cc_598 N_A_514_368#_c_889_n N_X_c_978_n 0.0315971f $X=8.205 $Y=2.375 $X2=0 $Y2=0
cc_599 N_A_514_368#_c_866_n N_X_c_978_n 0.0171986f $X=7.47 $Y=2.455 $X2=0 $Y2=0
cc_600 N_A_514_368#_c_867_n N_X_c_978_n 0.0209207f $X=8.37 $Y=2.455 $X2=0 $Y2=0
cc_601 N_A_514_368#_M1008_s N_X_c_974_n 0.00591199f $X=8.235 $Y=1.84 $X2=0 $Y2=0
cc_602 N_A_514_368#_c_859_n N_X_c_1044_n 0.0156632f $X=3.515 $Y=2.99 $X2=0 $Y2=0
cc_603 N_A_514_368#_M1017_s N_X_c_1051_n 0.00322588f $X=3.465 $Y=1.84 $X2=0
+ $Y2=0
cc_604 N_A_514_368#_c_859_n N_X_c_1051_n 0.00460492f $X=3.515 $Y=2.99 $X2=0
+ $Y2=0
cc_605 N_A_514_368#_c_965_p N_X_c_1051_n 0.0122761f $X=3.6 $Y=2.8 $X2=0 $Y2=0
cc_606 N_A_514_368#_c_861_n N_X_c_1051_n 0.00458951f $X=4.415 $Y=2.99 $X2=0
+ $Y2=0
cc_607 N_A_514_368#_c_861_n N_X_c_1013_n 0.0155605f $X=4.415 $Y=2.99 $X2=0 $Y2=0
cc_608 N_X_c_968_n N_VGND_M1029_d 0.011365f $X=4.105 $Y=0.765 $X2=0 $Y2=0
cc_609 N_X_c_969_n N_VGND_M1029_d 0.00238572f $X=4.19 $Y=1.01 $X2=0 $Y2=0
cc_610 N_X_c_971_n N_VGND_M1029_d 0.00189155f $X=4.275 $Y=1.095 $X2=0 $Y2=0
cc_611 N_X_c_970_n N_VGND_M1015_d 0.00391227f $X=6.835 $Y=1.095 $X2=0 $Y2=0
cc_612 N_X_c_970_n N_VGND_M1025_d 0.00391227f $X=6.835 $Y=1.095 $X2=0 $Y2=0
cc_613 N_X_c_968_n N_VGND_c_1135_n 0.0320467f $X=4.105 $Y=0.765 $X2=0 $Y2=0
cc_614 N_X_c_975_n N_VGND_c_1135_n 0.00221964f $X=3.375 $Y=0.66 $X2=0 $Y2=0
cc_615 N_X_c_968_n N_VGND_c_1140_n 0.0023127f $X=4.105 $Y=0.765 $X2=0 $Y2=0
cc_616 N_X_c_975_n N_VGND_c_1140_n 0.00937878f $X=3.375 $Y=0.66 $X2=0 $Y2=0
cc_617 N_X_c_968_n N_VGND_c_1143_n 0.00251932f $X=4.105 $Y=0.765 $X2=0 $Y2=0
cc_618 N_X_c_968_n N_VGND_c_1146_n 0.0106811f $X=4.105 $Y=0.765 $X2=0 $Y2=0
cc_619 N_X_c_975_n N_VGND_c_1146_n 0.0109286f $X=3.375 $Y=0.66 $X2=0 $Y2=0
cc_620 N_X_c_970_n N_A_877_74#_M1015_s 0.00463994f $X=6.835 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_621 N_X_c_970_n N_A_877_74#_M1016_s 0.00176891f $X=6.835 $Y=1.095 $X2=0 $Y2=0
cc_622 N_X_c_970_n N_A_877_74#_M1027_s 0.00176461f $X=6.835 $Y=1.095 $X2=0 $Y2=0
cc_623 N_X_c_972_n N_A_877_74#_M1012_s 0.00250873f $X=7.845 $Y=1.095 $X2=0 $Y2=0
cc_624 N_X_c_973_n N_A_877_74#_M1024_s 0.00757941f $X=8.335 $Y=1.095 $X2=0 $Y2=0
cc_625 N_X_c_970_n N_A_877_74#_c_1263_n 0.0151804f $X=6.835 $Y=1.095 $X2=0 $Y2=0
cc_626 N_X_M1010_d N_A_877_74#_c_1254_n 0.00176461f $X=6.86 $Y=0.37 $X2=0 $Y2=0
cc_627 N_X_c_970_n N_A_877_74#_c_1254_n 0.00304353f $X=6.835 $Y=1.095 $X2=0
+ $Y2=0
cc_628 N_X_c_1009_n N_A_877_74#_c_1254_n 0.0157964f $X=7 $Y=0.76 $X2=0 $Y2=0
cc_629 N_X_c_972_n N_A_877_74#_c_1254_n 0.00304353f $X=7.845 $Y=1.095 $X2=0
+ $Y2=0
cc_630 N_X_c_972_n N_A_877_74#_c_1278_n 0.020731f $X=7.845 $Y=1.095 $X2=0 $Y2=0
cc_631 N_X_M1020_d N_A_877_74#_c_1256_n 0.00176461f $X=7.79 $Y=0.37 $X2=0 $Y2=0
cc_632 N_X_c_972_n N_A_877_74#_c_1256_n 0.00304353f $X=7.845 $Y=1.095 $X2=0
+ $Y2=0
cc_633 N_X_c_1126_p N_A_877_74#_c_1256_n 0.0124895f $X=7.93 $Y=0.805 $X2=0 $Y2=0
cc_634 N_X_c_973_n N_A_877_74#_c_1256_n 0.00304353f $X=8.335 $Y=1.095 $X2=0
+ $Y2=0
cc_635 N_X_c_973_n N_A_877_74#_c_1257_n 0.0215474f $X=8.335 $Y=1.095 $X2=0 $Y2=0
cc_636 N_X_c_968_n N_A_877_74#_c_1258_n 0.0147083f $X=4.105 $Y=0.765 $X2=0 $Y2=0
cc_637 N_X_c_970_n N_A_877_74#_c_1258_n 0.0150829f $X=6.835 $Y=1.095 $X2=0 $Y2=0
cc_638 N_X_c_970_n N_A_877_74#_c_1268_n 0.0978095f $X=6.835 $Y=1.095 $X2=0 $Y2=0
cc_639 N_VGND_M1025_d N_A_877_74#_c_1261_n 0.00726893f $X=5.84 $Y=0.37 $X2=0
+ $Y2=0
cc_640 N_VGND_c_1137_n N_A_877_74#_c_1261_n 0.0251188f $X=6.06 $Y=0.335 $X2=0
+ $Y2=0
cc_641 N_VGND_c_1144_n N_A_877_74#_c_1261_n 0.00236055f $X=5.895 $Y=0 $X2=0
+ $Y2=0
cc_642 N_VGND_c_1145_n N_A_877_74#_c_1261_n 0.00236055f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_643 N_VGND_c_1146_n N_A_877_74#_c_1261_n 0.0102106f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_644 N_VGND_c_1145_n N_A_877_74#_c_1254_n 0.0420053f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_645 N_VGND_c_1146_n N_A_877_74#_c_1254_n 0.022853f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_646 N_VGND_c_1137_n N_A_877_74#_c_1255_n 0.0114117f $X=6.06 $Y=0.335 $X2=0
+ $Y2=0
cc_647 N_VGND_c_1145_n N_A_877_74#_c_1255_n 0.0176331f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_648 N_VGND_c_1146_n N_A_877_74#_c_1255_n 0.00956698f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_649 N_VGND_c_1145_n N_A_877_74#_c_1256_n 0.0566663f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_650 N_VGND_c_1146_n N_A_877_74#_c_1256_n 0.0314476f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_651 N_VGND_c_1135_n N_A_877_74#_c_1258_n 0.00853811f $X=3.925 $Y=0.345 $X2=0
+ $Y2=0
cc_652 N_VGND_c_1136_n N_A_877_74#_c_1258_n 0.00591149f $X=5.04 $Y=0.335 $X2=0
+ $Y2=0
cc_653 N_VGND_c_1143_n N_A_877_74#_c_1258_n 0.0107387f $X=4.875 $Y=0 $X2=0 $Y2=0
cc_654 N_VGND_c_1146_n N_A_877_74#_c_1258_n 0.00894442f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_655 N_VGND_M1015_d N_A_877_74#_c_1268_n 0.00726893f $X=4.82 $Y=0.37 $X2=0
+ $Y2=0
cc_656 N_VGND_c_1136_n N_A_877_74#_c_1268_n 0.0251188f $X=5.04 $Y=0.335 $X2=0
+ $Y2=0
cc_657 N_VGND_c_1143_n N_A_877_74#_c_1268_n 0.00236055f $X=4.875 $Y=0 $X2=0
+ $Y2=0
cc_658 N_VGND_c_1144_n N_A_877_74#_c_1268_n 0.00236055f $X=5.895 $Y=0 $X2=0
+ $Y2=0
cc_659 N_VGND_c_1146_n N_A_877_74#_c_1268_n 0.0102106f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_660 N_VGND_c_1136_n N_A_877_74#_c_1259_n 0.0060913f $X=5.04 $Y=0.335 $X2=0
+ $Y2=0
cc_661 N_VGND_c_1137_n N_A_877_74#_c_1259_n 0.0060913f $X=6.06 $Y=0.335 $X2=0
+ $Y2=0
cc_662 N_VGND_c_1144_n N_A_877_74#_c_1259_n 0.0141766f $X=5.895 $Y=0 $X2=0 $Y2=0
cc_663 N_VGND_c_1146_n N_A_877_74#_c_1259_n 0.0118057f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_664 N_VGND_c_1145_n N_A_877_74#_c_1260_n 0.0233048f $X=8.4 $Y=0 $X2=0 $Y2=0
cc_665 N_VGND_c_1146_n N_A_877_74#_c_1260_n 0.0126653f $X=8.4 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__and3_1.spice
* Created: Fri Aug 28 17:11:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__and3_1.pex.spice"
.subckt sky130_fd_sc_ms__and3_1  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1001 A_121_136# N_A_M1001_g N_A_27_398#_M1001_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1312 AS=0.1824 PD=1.05 PS=1.85 NRD=28.116 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1002 A_233_136# N_B_M1002_g A_121_136# VNB NLOWVT L=0.15 W=0.64 AD=0.111
+ AS=0.1312 PD=1.045 PS=1.05 NRD=22.2 NRS=28.116 M=1 R=4.26667 SA=75000.8
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1004 N_VGND_M1004_d N_C_M1004_g A_233_136# VNB NLOWVT L=0.15 W=0.64
+ AD=0.144093 AS=0.111 PD=1.08522 PS=1.045 NRD=15.468 NRS=22.2 M=1 R=4.26667
+ SA=75001.1 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1007 N_X_M1007_d N_A_27_398#_M1007_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.166607 PD=2.05 PS=1.25478 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_A_27_398#_M1006_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1554 AS=0.2352 PD=1.21 PS=2.24 NRD=10.5395 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90002.1 A=0.1512 P=2.04 MULT=1
MM1003 N_A_27_398#_M1003_d N_B_M1003_g N_VPWR_M1006_d VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.1554 PD=1.11 PS=1.21 NRD=0 NRS=10.5395 M=1 R=4.66667 SA=90000.7
+ SB=90001.5 A=0.1512 P=2.04 MULT=1
MM1005 N_VPWR_M1005_d N_C_M1005_g N_A_27_398#_M1003_d VPB PSHORT L=0.18 W=0.84
+ AD=0.298736 AS=0.1134 PD=1.55143 PS=1.11 NRD=6.4419 NRS=0 M=1 R=4.66667
+ SA=90001.2 SB=90001.1 A=0.1512 P=2.04 MULT=1
MM1000 N_X_M1000_d N_A_27_398#_M1000_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.398314 PD=2.8 PS=2.06857 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ms__and3_1.pxi.spice"
*
.ends
*
*

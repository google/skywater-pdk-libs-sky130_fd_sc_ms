* File: sky130_fd_sc_ms__o31a_1.pex.spice
* Created: Wed Sep  2 12:25:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O31A_1%A_84_48# 1 2 9 13 16 17 18 21 25 29 32 35 37
+ 40 41
r85 35 44 40.6969 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.587 $Y=1.485
+ $X2=0.587 $Y2=1.65
r86 35 43 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.587 $Y=1.485
+ $X2=0.587 $Y2=1.32
r87 34 37 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.59 $Y=1.485
+ $X2=0.71 $Y2=1.485
r88 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.485 $X2=0.59 $Y2=1.485
r89 32 41 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=3.17 $Y=1.95
+ $X2=3.17 $Y2=1.13
r90 27 41 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=3.085 $Y=0.96
+ $X2=3.085 $Y2=1.13
r91 27 29 11.6939 $w=3.38e-07 $l=3.45e-07 $layer=LI1_cond $X=3.085 $Y=0.96
+ $X2=3.085 $Y2=0.615
r92 26 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=2.035
+ $X2=2.36 $Y2=2.035
r93 25 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.085 $Y=2.035
+ $X2=3.17 $Y2=1.95
r94 25 26 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.085 $Y=2.035
+ $X2=2.525 $Y2=2.035
r95 21 23 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.36 $Y=2.375
+ $X2=2.36 $Y2=2.715
r96 19 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.36 $Y=2.12 $X2=2.36
+ $Y2=2.035
r97 19 21 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.36 $Y=2.12
+ $X2=2.36 $Y2=2.375
r98 17 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=2.035
+ $X2=2.36 $Y2=2.035
r99 17 18 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=2.195 $Y=2.035
+ $X2=0.795 $Y2=2.035
r100 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.71 $Y=1.95
+ $X2=0.795 $Y2=2.035
r101 15 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.71 $Y=1.65
+ $X2=0.71 $Y2=1.485
r102 15 16 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.71 $Y=1.65 $X2=0.71
+ $Y2=1.95
r103 13 44 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=0.515 $Y=2.4
+ $X2=0.515 $Y2=1.65
r104 9 43 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.495 $Y=0.74
+ $X2=0.495 $Y2=1.32
r105 2 40 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.84 $X2=2.36 $Y2=2.035
r106 2 23 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.84 $X2=2.36 $Y2=2.715
r107 2 21 600 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=1.84 $X2=2.36 $Y2=2.375
r108 1 29 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=2.87
+ $Y=0.47 $X2=3.08 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_1%A1 3 7 9 12 13
c40 7 0 1.19054e-19 $X=1.205 $Y=2.34
r41 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.515
+ $X2=1.13 $Y2=1.68
r42 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.515
+ $X2=1.13 $Y2=1.35
r43 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.515 $X2=1.13 $Y2=1.515
r44 9 13 4.93904 $w=3.48e-07 $l=1.5e-07 $layer=LI1_cond $X=1.14 $Y=1.665
+ $X2=1.14 $Y2=1.515
r45 7 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.205 $Y=2.34
+ $X2=1.205 $Y2=1.68
r46 3 14 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.075 $Y=0.79
+ $X2=1.075 $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_1%A2 3 7 9 12 13
c35 7 0 1.59866e-19 $X=1.625 $Y=2.34
r36 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.67 $Y=1.465
+ $X2=1.67 $Y2=1.63
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.67 $Y=1.465
+ $X2=1.67 $Y2=1.3
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.67
+ $Y=1.465 $X2=1.67 $Y2=1.465
r39 9 13 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=1.67 $Y=1.665 $X2=1.67
+ $Y2=1.465
r40 7 15 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=1.625 $Y=2.34
+ $X2=1.625 $Y2=1.63
r41 3 14 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.58 $Y=0.79 $X2=1.58
+ $Y2=1.3
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_1%A3 3 7 9 12 13
c38 13 0 1.59866e-19 $X=2.21 $Y=1.515
r39 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.515
+ $X2=2.21 $Y2=1.68
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.515
+ $X2=2.21 $Y2=1.35
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.21
+ $Y=1.515 $X2=2.21 $Y2=1.515
r42 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.21 $Y=1.665
+ $X2=2.21 $Y2=1.515
r43 7 14 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.3 $Y=0.79 $X2=2.3
+ $Y2=1.35
r44 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.135 $Y=2.34
+ $X2=2.135 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_1%B1 3 7 9 12 13
r32 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.75 $Y=1.515
+ $X2=2.75 $Y2=1.68
r33 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.75 $Y=1.515
+ $X2=2.75 $Y2=1.35
r34 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.75
+ $Y=1.515 $X2=2.75 $Y2=1.515
r35 9 13 4.67207 $w=3.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.73 $Y=1.665
+ $X2=2.73 $Y2=1.515
r36 7 14 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.795 $Y=0.79
+ $X2=2.795 $Y2=1.35
r37 3 15 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=2.675 $Y=2.26
+ $X2=2.675 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_1%X 1 2 9 13 14 15 16 23 32
c25 14 0 1.19054e-19 $X=0.155 $Y=1.95
r26 21 23 0.934413 $w=3.68e-07 $l=3e-08 $layer=LI1_cond $X=0.27 $Y=2.005
+ $X2=0.27 $Y2=2.035
r27 15 16 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.27 $Y=2.405
+ $X2=0.27 $Y2=2.775
r28 14 21 0.872119 $w=3.68e-07 $l=2.8e-08 $layer=LI1_cond $X=0.27 $Y=1.977
+ $X2=0.27 $Y2=2.005
r29 14 32 8.28963 $w=3.68e-07 $l=1.57e-07 $layer=LI1_cond $X=0.27 $Y=1.977
+ $X2=0.27 $Y2=1.82
r30 14 15 10.6835 $w=3.68e-07 $l=3.43e-07 $layer=LI1_cond $X=0.27 $Y=2.062
+ $X2=0.27 $Y2=2.405
r31 14 23 0.840972 $w=3.68e-07 $l=2.7e-08 $layer=LI1_cond $X=0.27 $Y=2.062
+ $X2=0.27 $Y2=2.035
r32 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.17 $Y=1.13 $X2=0.17
+ $Y2=1.82
r33 7 13 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.265 $Y=0.95
+ $X2=0.265 $Y2=1.13
r34 7 9 13.9254 $w=3.58e-07 $l=4.35e-07 $layer=LI1_cond $X=0.265 $Y=0.95
+ $X2=0.265 $Y2=0.515
r35 2 14 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.29 $Y2=1.985
r36 2 16 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.29 $Y2=2.815
r37 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_1%VPWR 1 2 9 13 16 17 18 20 33 34 37
r38 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 31 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 27 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r45 25 37 10.8012 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=1.09 $Y=3.33
+ $X2=0.857 $Y2=3.33
r46 25 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.09 $Y=3.33 $X2=1.2
+ $Y2=3.33
r47 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 20 37 10.8012 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.857 $Y2=3.33
r50 20 22 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 18 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 18 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 16 30 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.735 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 16 17 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=2.735 $Y=3.33
+ $X2=2.892 $Y2=3.33
r55 15 33 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.05 $Y=3.33 $X2=3.12
+ $Y2=3.33
r56 15 17 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=3.05 $Y=3.33
+ $X2=2.892 $Y2=3.33
r57 11 17 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.892 $Y=3.245
+ $X2=2.892 $Y2=3.33
r58 11 13 28.9025 $w=3.13e-07 $l=7.9e-07 $layer=LI1_cond $X=2.892 $Y=3.245
+ $X2=2.892 $Y2=2.455
r59 7 37 1.88438 $w=4.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.857 $Y=3.245
+ $X2=0.857 $Y2=3.33
r60 7 9 21.478 $w=4.63e-07 $l=8.35e-07 $layer=LI1_cond $X=0.857 $Y=3.245
+ $X2=0.857 $Y2=2.41
r61 2 13 600 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=1 $X=2.765
+ $Y=1.84 $X2=2.9 $Y2=2.455
r62 1 9 300 $w=1.7e-07 $l=7.1225e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.84 $X2=0.925 $Y2=2.41
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_1%VGND 1 2 9 15 18 19 20 22 35 36 39
r39 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r41 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r42 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r43 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r44 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r45 27 29 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.68
+ $Y2=0
r46 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r47 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r49 22 24 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r50 20 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r51 20 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r52 20 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r53 18 29 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=0 $X2=1.68
+ $Y2=0
r54 18 19 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=1.765 $Y=0 $X2=1.947
+ $Y2=0
r55 17 32 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.13 $Y=0 $X2=2.16
+ $Y2=0
r56 17 19 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=2.13 $Y=0 $X2=1.947
+ $Y2=0
r57 13 19 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.947 $Y=0.085
+ $X2=1.947 $Y2=0
r58 13 15 16.7341 $w=3.63e-07 $l=5.3e-07 $layer=LI1_cond $X=1.947 $Y=0.085
+ $X2=1.947 $Y2=0.615
r59 9 11 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.78 $Y=0.515
+ $X2=0.78 $Y2=0.965
r60 7 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0
r61 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0.515
r62 2 15 182 $w=1.7e-07 $l=3.55176e-07 $layer=licon1_NDIFF $count=1 $X=1.655
+ $Y=0.47 $X2=1.945 $Y2=0.615
r63 1 11 182 $w=1.7e-07 $l=6.9208e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.965
r64 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_1%A_230_94# 1 2 9 11 12 15
r32 13 15 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.58 $Y=0.96
+ $X2=2.58 $Y2=0.615
r33 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.415 $Y=1.045
+ $X2=2.58 $Y2=0.96
r34 11 12 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=2.415 $Y=1.045
+ $X2=1.46 $Y2=1.045
r35 7 12 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=1.292 $Y=0.96
+ $X2=1.46 $Y2=1.045
r36 7 9 11.8684 $w=3.33e-07 $l=3.45e-07 $layer=LI1_cond $X=1.292 $Y=0.96
+ $X2=1.292 $Y2=0.615
r37 2 15 91 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=2 $X=2.375
+ $Y=0.47 $X2=2.58 $Y2=0.615
r38 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.15
+ $Y=0.47 $X2=1.29 $Y2=0.615
.ends


* File: sky130_fd_sc_ms__a311o_2.spice
* Created: Wed Sep  2 11:54:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a311o_2.pex.spice"
.subckt sky130_fd_sc_ms__a311o_2  VNB VPB A3 A2 A1 B1 C1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_21_270#_M1002_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_21_270#_M1007_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=17.016 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1005 A_351_74# N_A3_M1005_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.74 AD=0.0777
+ AS=0.1554 PD=0.95 PS=1.16 NRD=8.1 NRS=5.664 M=1 R=4.93333 SA=75001.2
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1001 A_423_74# N_A2_M1001_g A_351_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1443
+ AS=0.0777 PD=1.13 PS=0.95 NRD=22.692 NRS=8.1 M=1 R=4.93333 SA=75001.6
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1011 N_A_21_270#_M1011_d N_A1_M1011_g A_423_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.1443 PD=1.13 PS=1.13 NRD=3.24 NRS=22.692 M=1 R=4.93333
+ SA=75002.1 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_B1_M1004_g N_A_21_270#_M1011_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.1443 PD=1.13 PS=1.13 NRD=3.24 NRS=14.592 M=1 R=4.93333
+ SA=75002.6 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1006 N_A_21_270#_M1006_d N_C1_M1006_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1443 PD=2.01 PS=1.13 NRD=0 NRS=14.592 M=1 R=4.93333 SA=75003.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_A_21_270#_M1000_g N_X_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2912 AS=0.1512 PD=2.76 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90002.9 A=0.2016 P=2.6 MULT=1
MM1012 N_VPWR_M1012_d N_A_21_270#_M1012_g N_X_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.196106 AS=0.1512 PD=1.54264 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90002.5 A=0.2016 P=2.6 MULT=1
MM1010 N_A_333_392#_M1010_d N_A3_M1010_g N_VPWR_M1012_d VPB PSHORT L=0.18 W=1
+ AD=0.15 AS=0.175094 PD=1.3 PS=1.37736 NRD=0 NRS=12.7853 M=1 R=5.55556
+ SA=90001.1 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_A2_M1008_g N_A_333_392#_M1010_d VPB PSHORT L=0.18 W=1
+ AD=0.255 AS=0.15 PD=1.51 PS=1.3 NRD=22.6353 NRS=4.9053 M=1 R=5.55556
+ SA=90001.6 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1009 N_A_333_392#_M1009_d N_A1_M1009_g N_VPWR_M1008_d VPB PSHORT L=0.18 W=1
+ AD=0.15 AS=0.255 PD=1.3 PS=1.51 NRD=4.9053 NRS=22.6353 M=1 R=5.55556
+ SA=90002.3 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1003 A_663_392# N_B1_M1003_g N_A_333_392#_M1009_d VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.15 PD=1.24 PS=1.3 NRD=12.7853 NRS=0 M=1 R=5.55556 SA=90002.8
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1013 N_A_21_270#_M1013_d N_C1_M1013_g A_663_392# VPB PSHORT L=0.18 W=1 AD=0.26
+ AS=0.12 PD=2.52 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556 SA=90003.2 SB=90000.2
+ A=0.18 P=2.36 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__a311o_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__o31ai_1.spice
* Created: Wed Sep  2 12:25:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o31ai_1.pex.spice"
.subckt sky130_fd_sc_ms__o31ai_1  VNB VPB A1 A2 A3 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1005 N_A_114_74#_M1005_d N_A1_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g N_A_114_74#_M1005_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.3492 AS=0.1036 PD=1.7 PS=1.02 NRD=13.776 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1001 N_A_114_74#_M1001_d N_A3_M1001_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.111 AS=0.3492 PD=1.04 PS=1.7 NRD=0 NRS=13.776 M=1 R=4.93333 SA=75001.6
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_B1_M1002_g N_A_114_74#_M1001_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2479 AS=0.111 PD=2.15 PS=1.04 NRD=8.1 NRS=3.24 M=1 R=4.93333 SA=75002.1
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1003 A_122_368# N_A1_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12 AD=0.1344
+ AS=0.3136 PD=1.36 PS=2.8 NRD=11.426 NRS=0 M=1 R=6.22222 SA=90000.2 SB=90002
+ A=0.2016 P=2.6 MULT=1
MM1000 A_206_368# N_A2_M1000_g A_122_368# VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.1344 PD=1.51 PS=1.36 NRD=24.6053 NRS=11.426 M=1 R=6.22222 SA=90000.6
+ SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1007 N_Y_M1007_d N_A3_M1007_g A_206_368# VPB PSHORT L=0.18 W=1.12 AD=0.3696
+ AS=0.2184 PD=1.78 PS=1.51 NRD=0 NRS=24.6053 M=1 R=6.22222 SA=90001.2 SB=90001
+ A=0.2016 P=2.6 MULT=1
MM1004 N_VPWR_M1004_d N_B1_M1004_g N_Y_M1007_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.3696 PD=2.8 PS=1.78 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ms__o31ai_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__o2bb2ai_2.pxi.spice
* Created: Wed Sep  2 12:24:35 2020
* 
x_PM_SKY130_FD_SC_MS__O2BB2AI_2%A1_N N_A1_N_M1001_g N_A1_N_M1007_g
+ N_A1_N_c_104_n N_A1_N_M1012_g N_A1_N_c_105_n N_A1_N_M1014_g N_A1_N_c_106_n
+ N_A1_N_c_107_n N_A1_N_c_115_n N_A1_N_c_122_p N_A1_N_c_116_n N_A1_N_c_165_p
+ N_A1_N_c_123_p N_A1_N_c_108_n A1_N N_A1_N_c_109_n A1_N
+ PM_SKY130_FD_SC_MS__O2BB2AI_2%A1_N
x_PM_SKY130_FD_SC_MS__O2BB2AI_2%A2_N N_A2_N_M1008_g N_A2_N_M1003_g
+ N_A2_N_M1019_g N_A2_N_M1018_g A2_N N_A2_N_c_202_n
+ PM_SKY130_FD_SC_MS__O2BB2AI_2%A2_N
x_PM_SKY130_FD_SC_MS__O2BB2AI_2%A_136_387# N_A_136_387#_M1008_d
+ N_A_136_387#_M1001_d N_A_136_387#_M1018_s N_A_136_387#_M1011_g
+ N_A_136_387#_M1000_g N_A_136_387#_c_264_n N_A_136_387#_M1016_g
+ N_A_136_387#_M1006_g N_A_136_387#_c_282_n N_A_136_387#_c_267_n
+ N_A_136_387#_c_268_n N_A_136_387#_c_356_p N_A_136_387#_c_269_n
+ N_A_136_387#_c_270_n N_A_136_387#_c_293_n N_A_136_387#_c_298_n
+ N_A_136_387#_c_271_n PM_SKY130_FD_SC_MS__O2BB2AI_2%A_136_387#
x_PM_SKY130_FD_SC_MS__O2BB2AI_2%B1 N_B1_M1010_g N_B1_M1004_g N_B1_M1013_g
+ N_B1_M1017_g N_B1_c_366_n N_B1_c_367_n N_B1_c_374_n N_B1_c_375_n B1
+ N_B1_c_369_n PM_SKY130_FD_SC_MS__O2BB2AI_2%B1
x_PM_SKY130_FD_SC_MS__O2BB2AI_2%B2 N_B2_c_451_n N_B2_M1002_g N_B2_M1005_g
+ N_B2_M1009_g N_B2_c_454_n N_B2_M1015_g B2 N_B2_c_456_n
+ PM_SKY130_FD_SC_MS__O2BB2AI_2%B2
x_PM_SKY130_FD_SC_MS__O2BB2AI_2%VPWR N_VPWR_M1001_s N_VPWR_M1003_d
+ N_VPWR_M1014_s N_VPWR_M1016_s N_VPWR_M1013_s N_VPWR_c_508_n N_VPWR_c_509_n
+ N_VPWR_c_510_n N_VPWR_c_511_n N_VPWR_c_512_n N_VPWR_c_513_n N_VPWR_c_514_n
+ N_VPWR_c_515_n VPWR N_VPWR_c_516_n N_VPWR_c_517_n N_VPWR_c_518_n
+ N_VPWR_c_519_n N_VPWR_c_520_n N_VPWR_c_521_n N_VPWR_c_507_n
+ PM_SKY130_FD_SC_MS__O2BB2AI_2%VPWR
x_PM_SKY130_FD_SC_MS__O2BB2AI_2%Y N_Y_M1000_d N_Y_M1011_d N_Y_M1005_d
+ N_Y_c_587_n N_Y_c_593_n N_Y_c_608_n Y Y Y Y Y Y
+ PM_SKY130_FD_SC_MS__O2BB2AI_2%Y
x_PM_SKY130_FD_SC_MS__O2BB2AI_2%A_799_368# N_A_799_368#_M1004_d
+ N_A_799_368#_M1009_s N_A_799_368#_c_634_n N_A_799_368#_c_630_n
+ N_A_799_368#_c_631_n N_A_799_368#_c_637_n
+ PM_SKY130_FD_SC_MS__O2BB2AI_2%A_799_368#
x_PM_SKY130_FD_SC_MS__O2BB2AI_2%VGND N_VGND_M1007_s N_VGND_M1012_s
+ N_VGND_M1010_s N_VGND_M1015_d N_VGND_c_658_n N_VGND_c_659_n N_VGND_c_660_n
+ N_VGND_c_661_n N_VGND_c_662_n VGND N_VGND_c_663_n N_VGND_c_664_n
+ N_VGND_c_665_n N_VGND_c_666_n N_VGND_c_667_n N_VGND_c_668_n N_VGND_c_669_n
+ N_VGND_c_670_n PM_SKY130_FD_SC_MS__O2BB2AI_2%VGND
x_PM_SKY130_FD_SC_MS__O2BB2AI_2%A_134_74# N_A_134_74#_M1007_d
+ N_A_134_74#_M1019_s N_A_134_74#_c_732_n N_A_134_74#_c_730_n
+ N_A_134_74#_c_731_n N_A_134_74#_c_735_n
+ PM_SKY130_FD_SC_MS__O2BB2AI_2%A_134_74#
x_PM_SKY130_FD_SC_MS__O2BB2AI_2%A_518_74# N_A_518_74#_M1000_s
+ N_A_518_74#_M1006_s N_A_518_74#_M1002_s N_A_518_74#_M1017_d
+ N_A_518_74#_c_754_n N_A_518_74#_c_755_n N_A_518_74#_c_756_n
+ N_A_518_74#_c_767_n N_A_518_74#_c_768_n N_A_518_74#_c_757_n
+ N_A_518_74#_c_758_n N_A_518_74#_c_774_n N_A_518_74#_c_759_n
+ N_A_518_74#_c_760_n N_A_518_74#_c_788_n
+ PM_SKY130_FD_SC_MS__O2BB2AI_2%A_518_74#
cc_1 VNB N_A1_N_M1007_g 0.033863f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.69
cc_2 VNB N_A1_N_c_104_n 0.0160204f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.085
cc_3 VNB N_A1_N_c_105_n 0.0468589f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=1.68
cc_4 VNB N_A1_N_c_106_n 0.0444554f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.465
cc_5 VNB N_A1_N_c_107_n 0.0133717f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.3
cc_6 VNB N_A1_N_c_108_n 0.00491898f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=1.515
cc_7 VNB N_A1_N_c_109_n 0.0131935f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.465
cc_8 VNB A1_N 0.00134219f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.665
cc_9 VNB N_A2_N_M1008_g 0.0323868f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.355
cc_10 VNB N_A2_N_M1019_g 0.0339291f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=0.69
cc_11 VNB A2_N 0.00179472f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.3
cc_12 VNB N_A2_N_c_202_n 0.0316384f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=2.517
cc_13 VNB N_A_136_387#_M1011_g 0.00183388f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=1.68
cc_14 VNB N_A_136_387#_M1000_g 0.0224193f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.465
cc_15 VNB N_A_136_387#_c_264_n 0.0680725f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.5
cc_16 VNB N_A_136_387#_M1016_g 0.00270766f $X=-0.19 $Y=-0.245 $X2=2.165
+ $Y2=2.535
cc_17 VNB N_A_136_387#_M1006_g 0.0209341f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=2.415
cc_18 VNB N_A_136_387#_c_267_n 0.00267999f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=1.515
cc_19 VNB N_A_136_387#_c_268_n 0.00262414f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=1.515
cc_20 VNB N_A_136_387#_c_269_n 0.0264071f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.465
cc_21 VNB N_A_136_387#_c_270_n 0.00454919f $X=-0.19 $Y=-0.245 $X2=2.09 $Y2=1.515
cc_22 VNB N_A_136_387#_c_271_n 0.0140213f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.465
cc_23 VNB N_B1_M1010_g 0.0255172f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.355
cc_24 VNB N_B1_M1017_g 0.0337117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B1_c_366_n 0.00205059f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=2.5
cc_26 VNB N_B1_c_367_n 0.0270624f $X=-0.19 $Y=-0.245 $X2=2.165 $Y2=2.535
cc_27 VNB B1 0.0201105f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=2.415
cc_28 VNB N_B1_c_369_n 0.0288675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B2_c_451_n 0.0176191f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.72
cc_30 VNB N_B2_M1005_g 0.00584866f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.69
cc_31 VNB N_B2_M1009_g 0.00596185f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=0.69
cc_32 VNB N_B2_c_454_n 0.0172889f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=1.68
cc_33 VNB B2 0.00363541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_B2_c_456_n 0.0420234f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=2.415
cc_35 VNB N_VPWR_c_507_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB Y 0.00205679f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=2.535
cc_37 VNB N_VGND_c_658_n 0.01317f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=2.26
cc_38 VNB N_VGND_c_659_n 0.0407813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_660_n 0.0126674f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=2.5
cc_40 VNB N_VGND_c_661_n 0.00533463f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=2.45
cc_41 VNB N_VGND_c_662_n 0.00330537f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=1.515
cc_42 VNB N_VGND_c_663_n 0.0385965f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=1.515
cc_43 VNB N_VGND_c_664_n 0.0396346f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=1.465
cc_44 VNB N_VGND_c_665_n 0.0163741f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.69
cc_45 VNB N_VGND_c_666_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_667_n 0.322373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_668_n 0.00499734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_669_n 0.00615422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_670_n 0.00629135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_134_74#_c_730_n 0.0045598f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=0.69
cc_51 VNB N_A_134_74#_c_731_n 0.00203831f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=1.68
cc_52 VNB N_A_518_74#_c_754_n 0.00365422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_518_74#_c_755_n 0.00459841f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.3
cc_54 VNB N_A_518_74#_c_756_n 0.0037722f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.5
cc_55 VNB N_A_518_74#_c_757_n 0.01028f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=2.415
cc_56 VNB N_A_518_74#_c_758_n 0.00225496f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=1.515
cc_57 VNB N_A_518_74#_c_759_n 0.0217561f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=1.515
cc_58 VNB N_A_518_74#_c_760_n 0.0177969f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_59 VPB N_A1_N_M1001_g 0.0246879f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=2.355
cc_60 VPB N_A1_N_c_105_n 0.0086743f $X=-0.19 $Y=1.66 $X2=2.205 $Y2=1.68
cc_61 VPB N_A1_N_M1014_g 0.0242927f $X=-0.19 $Y=1.66 $X2=2.205 $Y2=2.26
cc_62 VPB N_A1_N_c_107_n 0.00326705f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.3
cc_63 VPB N_A1_N_c_115_n 0.00702792f $X=-0.19 $Y=1.66 $X2=0.355 $Y2=2.5
cc_64 VPB N_A1_N_c_116_n 0.00191281f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=2.45
cc_65 VPB N_A1_N_c_108_n 4.59347e-19 $X=-0.19 $Y=1.66 $X2=2.25 $Y2=1.515
cc_66 VPB A1_N 0.0300805f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.665
cc_67 VPB N_A2_N_M1003_g 0.02199f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=0.69
cc_68 VPB N_A2_N_M1018_g 0.026223f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB A2_N 0.00320605f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.3
cc_70 VPB N_A2_N_c_202_n 0.0197771f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=2.517
cc_71 VPB N_A_136_387#_M1011_g 0.0256048f $X=-0.19 $Y=1.66 $X2=2.205 $Y2=1.68
cc_72 VPB N_A_136_387#_M1016_g 0.0232625f $X=-0.19 $Y=1.66 $X2=2.165 $Y2=2.535
cc_73 VPB N_B1_M1004_g 0.0207306f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=0.69
cc_74 VPB N_B1_M1013_g 0.0243541f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=0.69
cc_75 VPB N_B1_c_366_n 7.62107e-19 $X=-0.19 $Y=1.66 $X2=0.355 $Y2=2.5
cc_76 VPB N_B1_c_367_n 0.00564782f $X=-0.19 $Y=1.66 $X2=2.165 $Y2=2.535
cc_77 VPB N_B1_c_374_n 0.0124295f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=1.68
cc_78 VPB N_B1_c_375_n 0.00104096f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=2.45
cc_79 VPB B1 0.00978549f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=2.415
cc_80 VPB N_B1_c_369_n 0.00581884f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_B2_M1005_g 0.0206071f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=0.69
cc_82 VPB N_B2_M1009_g 0.0206233f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=0.69
cc_83 VPB N_VPWR_c_508_n 0.0121899f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.465
cc_84 VPB N_VPWR_c_509_n 0.0282721f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=2.5
cc_85 VPB N_VPWR_c_510_n 0.0207138f $X=-0.19 $Y=1.66 $X2=2.165 $Y2=2.535
cc_86 VPB N_VPWR_c_511_n 0.0231606f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=2.415
cc_87 VPB N_VPWR_c_512_n 0.0187296f $X=-0.19 $Y=1.66 $X2=2.13 $Y2=1.515
cc_88 VPB N_VPWR_c_513_n 0.00855808f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_514_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.315 $Y2=1.465
cc_90 VPB N_VPWR_c_515_n 0.0498488f $X=-0.19 $Y=1.66 $X2=0.315 $Y2=1.465
cc_91 VPB N_VPWR_c_516_n 0.0283053f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.69
cc_92 VPB N_VPWR_c_517_n 0.0174051f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_518_n 0.0389302f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_519_n 0.00631873f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_520_n 0.00613202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_521_n 0.00631973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_507_n 0.0834902f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_Y_c_587_n 0.00247671f $X=-0.19 $Y=1.66 $X2=2.205 $Y2=1.68
cc_99 VPB Y 0.00179517f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=2.535
cc_100 VPB N_A_799_368#_c_630_n 0.00388794f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=0.69
cc_101 VPB N_A_799_368#_c_631_n 0.00196526f $X=-0.19 $Y=1.66 $X2=2.205 $Y2=1.68
cc_102 N_A1_N_M1007_g N_A2_N_M1008_g 0.0169811f $X=0.595 $Y=0.69 $X2=0 $Y2=0
cc_103 N_A1_N_c_109_n N_A2_N_M1008_g 2.01039e-19 $X=0.315 $Y=1.465 $X2=0 $Y2=0
cc_104 N_A1_N_M1001_g N_A2_N_M1003_g 0.0226382f $X=0.59 $Y=2.355 $X2=0 $Y2=0
cc_105 N_A1_N_c_122_p N_A2_N_M1003_g 0.0141495f $X=2.165 $Y=2.535 $X2=0 $Y2=0
cc_106 N_A1_N_c_123_p N_A2_N_M1003_g 9.76371e-19 $X=0.82 $Y=2.517 $X2=0 $Y2=0
cc_107 N_A1_N_c_104_n N_A2_N_M1019_g 0.0276245f $X=1.96 $Y=1.085 $X2=0 $Y2=0
cc_108 N_A1_N_c_105_n N_A2_N_M1019_g 0.00733936f $X=2.205 $Y=1.68 $X2=0 $Y2=0
cc_109 N_A1_N_c_108_n N_A2_N_M1019_g 5.52541e-19 $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_110 N_A1_N_c_122_p N_A2_N_M1018_g 0.0146368f $X=2.165 $Y=2.535 $X2=0 $Y2=0
cc_111 N_A1_N_c_116_n N_A2_N_M1018_g 0.00175829f $X=2.25 $Y=2.45 $X2=0 $Y2=0
cc_112 N_A1_N_c_105_n A2_N 8.01605e-19 $X=2.205 $Y=1.68 $X2=0 $Y2=0
cc_113 N_A1_N_M1014_g A2_N 7.32208e-19 $X=2.205 $Y=2.26 $X2=0 $Y2=0
cc_114 N_A1_N_c_116_n A2_N 0.00428262f $X=2.25 $Y=2.45 $X2=0 $Y2=0
cc_115 N_A1_N_c_108_n A2_N 0.0191382f $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_116 N_A1_N_c_105_n N_A2_N_c_202_n 0.0148825f $X=2.205 $Y=1.68 $X2=0 $Y2=0
cc_117 N_A1_N_M1014_g N_A2_N_c_202_n 0.0314509f $X=2.205 $Y=2.26 $X2=0 $Y2=0
cc_118 N_A1_N_c_107_n N_A2_N_c_202_n 0.0396193f $X=0.5 $Y=1.3 $X2=0 $Y2=0
cc_119 N_A1_N_c_108_n N_A2_N_c_202_n 2.63377e-19 $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_120 N_A1_N_c_122_p N_A_136_387#_M1001_d 0.0021896f $X=2.165 $Y=2.535 $X2=0
+ $Y2=0
cc_121 N_A1_N_c_123_p N_A_136_387#_M1001_d 0.00292161f $X=0.82 $Y=2.517 $X2=0
+ $Y2=0
cc_122 N_A1_N_c_122_p N_A_136_387#_M1018_s 0.00919441f $X=2.165 $Y=2.535 $X2=0
+ $Y2=0
cc_123 N_A1_N_c_105_n N_A_136_387#_M1011_g 0.0128346f $X=2.205 $Y=1.68 $X2=0
+ $Y2=0
cc_124 N_A1_N_c_116_n N_A_136_387#_M1011_g 0.00112177f $X=2.25 $Y=2.45 $X2=0
+ $Y2=0
cc_125 N_A1_N_c_108_n N_A_136_387#_M1011_g 4.11777e-19 $X=2.25 $Y=1.515 $X2=0
+ $Y2=0
cc_126 N_A1_N_c_105_n N_A_136_387#_c_264_n 0.0196063f $X=2.205 $Y=1.68 $X2=0
+ $Y2=0
cc_127 N_A1_N_c_108_n N_A_136_387#_c_264_n 9.3018e-19 $X=2.25 $Y=1.515 $X2=0
+ $Y2=0
cc_128 N_A1_N_M1001_g N_A_136_387#_c_282_n 0.0106935f $X=0.59 $Y=2.355 $X2=0
+ $Y2=0
cc_129 N_A1_N_M1007_g N_A_136_387#_c_282_n 0.00125799f $X=0.595 $Y=0.69 $X2=0
+ $Y2=0
cc_130 N_A1_N_c_107_n N_A_136_387#_c_282_n 0.0117293f $X=0.5 $Y=1.3 $X2=0 $Y2=0
cc_131 N_A1_N_c_122_p N_A_136_387#_c_282_n 0.00702775f $X=2.165 $Y=2.535 $X2=0
+ $Y2=0
cc_132 N_A1_N_c_123_p N_A_136_387#_c_282_n 0.00903475f $X=0.82 $Y=2.517 $X2=0
+ $Y2=0
cc_133 N_A1_N_c_109_n N_A_136_387#_c_282_n 0.0248813f $X=0.315 $Y=1.465 $X2=0
+ $Y2=0
cc_134 A1_N N_A_136_387#_c_282_n 0.0317177f $X=0.24 $Y=1.665 $X2=0 $Y2=0
cc_135 N_A1_N_M1007_g N_A_136_387#_c_268_n 0.0102229f $X=0.595 $Y=0.69 $X2=0
+ $Y2=0
cc_136 N_A1_N_c_104_n N_A_136_387#_c_269_n 0.00951367f $X=1.96 $Y=1.085 $X2=0
+ $Y2=0
cc_137 N_A1_N_c_105_n N_A_136_387#_c_269_n 0.0163257f $X=2.205 $Y=1.68 $X2=0
+ $Y2=0
cc_138 N_A1_N_c_108_n N_A_136_387#_c_269_n 0.0274115f $X=2.25 $Y=1.515 $X2=0
+ $Y2=0
cc_139 N_A1_N_c_105_n N_A_136_387#_c_293_n 7.47741e-19 $X=2.205 $Y=1.68 $X2=0
+ $Y2=0
cc_140 N_A1_N_M1014_g N_A_136_387#_c_293_n 0.00267534f $X=2.205 $Y=2.26 $X2=0
+ $Y2=0
cc_141 N_A1_N_c_122_p N_A_136_387#_c_293_n 0.0164722f $X=2.165 $Y=2.535 $X2=0
+ $Y2=0
cc_142 N_A1_N_c_116_n N_A_136_387#_c_293_n 0.0256974f $X=2.25 $Y=2.45 $X2=0
+ $Y2=0
cc_143 N_A1_N_c_108_n N_A_136_387#_c_293_n 0.00163364f $X=2.25 $Y=1.515 $X2=0
+ $Y2=0
cc_144 N_A1_N_c_122_p N_A_136_387#_c_298_n 0.0397144f $X=2.165 $Y=2.535 $X2=0
+ $Y2=0
cc_145 N_A1_N_c_105_n N_A_136_387#_c_271_n 0.00394852f $X=2.205 $Y=1.68 $X2=0
+ $Y2=0
cc_146 N_A1_N_c_108_n N_A_136_387#_c_271_n 0.0225013f $X=2.25 $Y=1.515 $X2=0
+ $Y2=0
cc_147 N_A1_N_c_115_n N_VPWR_M1001_s 0.00410969f $X=0.355 $Y=2.5 $X2=-0.19
+ $Y2=-0.245
cc_148 N_A1_N_c_165_p N_VPWR_M1001_s 0.00422357f $X=0.65 $Y=2.517 $X2=-0.19
+ $Y2=-0.245
cc_149 A1_N N_VPWR_M1001_s 0.0107166f $X=0.24 $Y=1.665 $X2=-0.19 $Y2=-0.245
cc_150 N_A1_N_c_122_p N_VPWR_M1003_d 0.00766107f $X=2.165 $Y=2.535 $X2=0 $Y2=0
cc_151 N_A1_N_M1001_g N_VPWR_c_509_n 0.00594909f $X=0.59 $Y=2.355 $X2=0 $Y2=0
cc_152 N_A1_N_c_115_n N_VPWR_c_509_n 0.0199258f $X=0.355 $Y=2.5 $X2=0 $Y2=0
cc_153 N_A1_N_c_165_p N_VPWR_c_509_n 0.00688446f $X=0.65 $Y=2.517 $X2=0 $Y2=0
cc_154 N_A1_N_M1001_g N_VPWR_c_510_n 0.00428077f $X=0.59 $Y=2.355 $X2=0 $Y2=0
cc_155 N_A1_N_c_165_p N_VPWR_c_510_n 0.00231342f $X=0.65 $Y=2.517 $X2=0 $Y2=0
cc_156 N_A1_N_c_123_p N_VPWR_c_510_n 0.00658386f $X=0.82 $Y=2.517 $X2=0 $Y2=0
cc_157 N_A1_N_c_122_p N_VPWR_c_511_n 0.0255558f $X=2.165 $Y=2.535 $X2=0 $Y2=0
cc_158 N_A1_N_M1014_g N_VPWR_c_512_n 0.00772614f $X=2.205 $Y=2.26 $X2=0 $Y2=0
cc_159 N_A1_N_c_116_n N_VPWR_c_512_n 0.0260112f $X=2.25 $Y=2.45 $X2=0 $Y2=0
cc_160 N_A1_N_M1014_g N_VPWR_c_516_n 0.00378744f $X=2.205 $Y=2.26 $X2=0 $Y2=0
cc_161 N_A1_N_c_122_p N_VPWR_c_516_n 0.010552f $X=2.165 $Y=2.535 $X2=0 $Y2=0
cc_162 N_A1_N_M1001_g N_VPWR_c_507_n 0.00587053f $X=0.59 $Y=2.355 $X2=0 $Y2=0
cc_163 N_A1_N_M1014_g N_VPWR_c_507_n 0.00555093f $X=2.205 $Y=2.26 $X2=0 $Y2=0
cc_164 N_A1_N_c_115_n N_VPWR_c_507_n 9.6483e-19 $X=0.355 $Y=2.5 $X2=0 $Y2=0
cc_165 N_A1_N_c_122_p N_VPWR_c_507_n 0.023291f $X=2.165 $Y=2.535 $X2=0 $Y2=0
cc_166 N_A1_N_c_165_p N_VPWR_c_507_n 0.00557097f $X=0.65 $Y=2.517 $X2=0 $Y2=0
cc_167 N_A1_N_c_123_p N_VPWR_c_507_n 0.0142518f $X=0.82 $Y=2.517 $X2=0 $Y2=0
cc_168 N_A1_N_c_116_n Y 0.00415404f $X=2.25 $Y=2.45 $X2=0 $Y2=0
cc_169 N_A1_N_c_108_n Y 0.0015446f $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_170 N_A1_N_M1007_g N_VGND_c_659_n 0.0164257f $X=0.595 $Y=0.69 $X2=0 $Y2=0
cc_171 N_A1_N_c_106_n N_VGND_c_659_n 0.00713769f $X=0.5 $Y=1.465 $X2=0 $Y2=0
cc_172 N_A1_N_c_109_n N_VGND_c_659_n 0.0196148f $X=0.315 $Y=1.465 $X2=0 $Y2=0
cc_173 N_A1_N_c_104_n N_VGND_c_660_n 0.00500836f $X=1.96 $Y=1.085 $X2=0 $Y2=0
cc_174 N_A1_N_M1007_g N_VGND_c_663_n 0.00430908f $X=0.595 $Y=0.69 $X2=0 $Y2=0
cc_175 N_A1_N_c_104_n N_VGND_c_663_n 0.00430908f $X=1.96 $Y=1.085 $X2=0 $Y2=0
cc_176 N_A1_N_M1007_g N_VGND_c_667_n 0.0081951f $X=0.595 $Y=0.69 $X2=0 $Y2=0
cc_177 N_A1_N_c_104_n N_VGND_c_667_n 0.00820555f $X=1.96 $Y=1.085 $X2=0 $Y2=0
cc_178 N_A1_N_M1007_g N_A_134_74#_c_732_n 0.00569679f $X=0.595 $Y=0.69 $X2=0
+ $Y2=0
cc_179 N_A1_N_c_104_n N_A_134_74#_c_730_n 0.00393598f $X=1.96 $Y=1.085 $X2=0
+ $Y2=0
cc_180 N_A1_N_M1007_g N_A_134_74#_c_731_n 0.00327745f $X=0.595 $Y=0.69 $X2=0
+ $Y2=0
cc_181 N_A1_N_c_104_n N_A_134_74#_c_735_n 0.00505485f $X=1.96 $Y=1.085 $X2=0
+ $Y2=0
cc_182 N_A2_N_M1008_g N_A_136_387#_c_282_n 0.00529294f $X=1.025 $Y=0.69 $X2=0
+ $Y2=0
cc_183 N_A2_N_M1003_g N_A_136_387#_c_282_n 0.00674994f $X=1.04 $Y=2.355 $X2=0
+ $Y2=0
cc_184 N_A2_N_M1019_g N_A_136_387#_c_282_n 8.01327e-19 $X=1.53 $Y=0.69 $X2=0
+ $Y2=0
cc_185 N_A2_N_M1018_g N_A_136_387#_c_282_n 7.56691e-19 $X=1.66 $Y=2.355 $X2=0
+ $Y2=0
cc_186 A2_N N_A_136_387#_c_282_n 0.0129425f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_187 N_A2_N_c_202_n N_A_136_387#_c_282_n 0.0121389f $X=1.66 $Y=1.61 $X2=0
+ $Y2=0
cc_188 N_A2_N_M1008_g N_A_136_387#_c_267_n 0.0127505f $X=1.025 $Y=0.69 $X2=0
+ $Y2=0
cc_189 N_A2_N_M1008_g N_A_136_387#_c_268_n 0.00312194f $X=1.025 $Y=0.69 $X2=0
+ $Y2=0
cc_190 N_A2_N_M1019_g N_A_136_387#_c_269_n 0.0128475f $X=1.53 $Y=0.69 $X2=0
+ $Y2=0
cc_191 A2_N N_A_136_387#_c_269_n 0.0206507f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_192 N_A2_N_c_202_n N_A_136_387#_c_269_n 0.00356193f $X=1.66 $Y=1.61 $X2=0
+ $Y2=0
cc_193 N_A2_N_M1008_g N_A_136_387#_c_270_n 0.00307017f $X=1.025 $Y=0.69 $X2=0
+ $Y2=0
cc_194 N_A2_N_M1019_g N_A_136_387#_c_270_n 0.00311703f $X=1.53 $Y=0.69 $X2=0
+ $Y2=0
cc_195 A2_N N_A_136_387#_c_270_n 0.00253019f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_196 N_A2_N_c_202_n N_A_136_387#_c_270_n 0.00538053f $X=1.66 $Y=1.61 $X2=0
+ $Y2=0
cc_197 N_A2_N_M1018_g N_A_136_387#_c_293_n 0.00234576f $X=1.66 $Y=2.355 $X2=0
+ $Y2=0
cc_198 N_A2_N_M1003_g N_A_136_387#_c_298_n 0.0155662f $X=1.04 $Y=2.355 $X2=0
+ $Y2=0
cc_199 N_A2_N_M1018_g N_A_136_387#_c_298_n 0.0134019f $X=1.66 $Y=2.355 $X2=0
+ $Y2=0
cc_200 A2_N N_A_136_387#_c_298_n 0.028811f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_201 N_A2_N_c_202_n N_A_136_387#_c_298_n 0.00515598f $X=1.66 $Y=1.61 $X2=0
+ $Y2=0
cc_202 N_A2_N_M1003_g N_VPWR_c_510_n 0.00425758f $X=1.04 $Y=2.355 $X2=0 $Y2=0
cc_203 N_A2_N_M1003_g N_VPWR_c_511_n 0.00337464f $X=1.04 $Y=2.355 $X2=0 $Y2=0
cc_204 N_A2_N_M1018_g N_VPWR_c_511_n 0.00337464f $X=1.66 $Y=2.355 $X2=0 $Y2=0
cc_205 N_A2_N_M1018_g N_VPWR_c_516_n 0.00425758f $X=1.66 $Y=2.355 $X2=0 $Y2=0
cc_206 N_A2_N_M1003_g N_VPWR_c_507_n 0.00587053f $X=1.04 $Y=2.355 $X2=0 $Y2=0
cc_207 N_A2_N_M1018_g N_VPWR_c_507_n 0.00587053f $X=1.66 $Y=2.355 $X2=0 $Y2=0
cc_208 N_A2_N_M1008_g N_VGND_c_663_n 0.00278247f $X=1.025 $Y=0.69 $X2=0 $Y2=0
cc_209 N_A2_N_M1019_g N_VGND_c_663_n 0.00278247f $X=1.53 $Y=0.69 $X2=0 $Y2=0
cc_210 N_A2_N_M1008_g N_VGND_c_667_n 0.00354226f $X=1.025 $Y=0.69 $X2=0 $Y2=0
cc_211 N_A2_N_M1019_g N_VGND_c_667_n 0.00354226f $X=1.53 $Y=0.69 $X2=0 $Y2=0
cc_212 N_A2_N_M1008_g N_A_134_74#_c_732_n 0.00719216f $X=1.025 $Y=0.69 $X2=0
+ $Y2=0
cc_213 N_A2_N_M1019_g N_A_134_74#_c_732_n 6.34304e-19 $X=1.53 $Y=0.69 $X2=0
+ $Y2=0
cc_214 N_A2_N_M1008_g N_A_134_74#_c_730_n 0.0104897f $X=1.025 $Y=0.69 $X2=0
+ $Y2=0
cc_215 N_A2_N_M1019_g N_A_134_74#_c_730_n 0.010847f $X=1.53 $Y=0.69 $X2=0 $Y2=0
cc_216 N_A2_N_M1008_g N_A_134_74#_c_731_n 0.00184341f $X=1.025 $Y=0.69 $X2=0
+ $Y2=0
cc_217 N_A2_N_M1008_g N_A_134_74#_c_735_n 5.5881e-19 $X=1.025 $Y=0.69 $X2=0
+ $Y2=0
cc_218 N_A2_N_M1019_g N_A_134_74#_c_735_n 0.00648761f $X=1.53 $Y=0.69 $X2=0
+ $Y2=0
cc_219 N_A_136_387#_M1006_g N_B1_M1010_g 0.017351f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A_136_387#_M1016_g N_B1_M1004_g 0.0233811f $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_221 N_A_136_387#_c_264_n N_B1_c_366_n 0.00145822f $X=3.365 $Y=1.605 $X2=0
+ $Y2=0
cc_222 N_A_136_387#_M1016_g N_B1_c_366_n 3.41312e-19 $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_223 N_A_136_387#_c_264_n N_B1_c_367_n 0.0183309f $X=3.365 $Y=1.605 $X2=0
+ $Y2=0
cc_224 N_A_136_387#_M1016_g N_B1_c_375_n 0.00163413f $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_225 N_A_136_387#_c_298_n N_VPWR_M1003_d 0.00921087f $X=1.72 $Y=2.115 $X2=0
+ $Y2=0
cc_226 N_A_136_387#_M1011_g N_VPWR_c_512_n 0.0192271f $X=2.9 $Y=2.4 $X2=0 $Y2=0
cc_227 N_A_136_387#_c_264_n N_VPWR_c_512_n 0.00237199f $X=3.365 $Y=1.605 $X2=0
+ $Y2=0
cc_228 N_A_136_387#_M1016_g N_VPWR_c_512_n 6.65254e-19 $X=3.365 $Y=2.4 $X2=0
+ $Y2=0
cc_229 N_A_136_387#_c_271_n N_VPWR_c_512_n 0.0260338f $X=2.67 $Y=1.095 $X2=0
+ $Y2=0
cc_230 N_A_136_387#_M1016_g N_VPWR_c_513_n 0.00202402f $X=3.365 $Y=2.4 $X2=0
+ $Y2=0
cc_231 N_A_136_387#_M1011_g N_VPWR_c_517_n 0.00475445f $X=2.9 $Y=2.4 $X2=0 $Y2=0
cc_232 N_A_136_387#_M1016_g N_VPWR_c_517_n 0.00537895f $X=3.365 $Y=2.4 $X2=0
+ $Y2=0
cc_233 N_A_136_387#_M1011_g N_VPWR_c_507_n 0.00938812f $X=2.9 $Y=2.4 $X2=0 $Y2=0
cc_234 N_A_136_387#_M1016_g N_VPWR_c_507_n 0.0103734f $X=3.365 $Y=2.4 $X2=0
+ $Y2=0
cc_235 N_A_136_387#_M1011_g N_Y_c_587_n 2.8281e-19 $X=2.9 $Y=2.4 $X2=0 $Y2=0
cc_236 N_A_136_387#_M1016_g N_Y_c_587_n 0.0097592f $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_237 N_A_136_387#_M1016_g N_Y_c_593_n 0.0194965f $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_238 N_A_136_387#_M1000_g Y 0.0139043f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_239 N_A_136_387#_M1006_g Y 0.00541215f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A_136_387#_c_271_n Y 0.00600767f $X=2.67 $Y=1.095 $X2=0 $Y2=0
cc_241 N_A_136_387#_M1000_g Y 0.0040844f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A_136_387#_c_264_n Y 0.0251256f $X=3.365 $Y=1.605 $X2=0 $Y2=0
cc_243 N_A_136_387#_M1016_g Y 0.00995211f $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_244 N_A_136_387#_c_271_n Y 0.0326778f $X=2.67 $Y=1.095 $X2=0 $Y2=0
cc_245 N_A_136_387#_M1016_g Y 4.77e-19 $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_246 N_A_136_387#_M1000_g N_VGND_c_660_n 0.00164546f $X=2.95 $Y=0.74 $X2=0
+ $Y2=0
cc_247 N_A_136_387#_c_269_n N_VGND_c_660_n 0.0196286f $X=2.505 $Y=1.095 $X2=0
+ $Y2=0
cc_248 N_A_136_387#_M1000_g N_VGND_c_664_n 0.00278271f $X=2.95 $Y=0.74 $X2=0
+ $Y2=0
cc_249 N_A_136_387#_M1006_g N_VGND_c_664_n 0.00278271f $X=3.38 $Y=0.74 $X2=0
+ $Y2=0
cc_250 N_A_136_387#_M1000_g N_VGND_c_667_n 0.00358427f $X=2.95 $Y=0.74 $X2=0
+ $Y2=0
cc_251 N_A_136_387#_M1006_g N_VGND_c_667_n 0.00353799f $X=3.38 $Y=0.74 $X2=0
+ $Y2=0
cc_252 N_A_136_387#_c_268_n N_A_134_74#_c_732_n 0.0242411f $X=0.98 $Y=1.19 $X2=0
+ $Y2=0
cc_253 N_A_136_387#_M1008_d N_A_134_74#_c_730_n 0.00262408f $X=1.1 $Y=0.37 $X2=0
+ $Y2=0
cc_254 N_A_136_387#_c_356_p N_A_134_74#_c_730_n 0.0174435f $X=1.24 $Y=0.78 $X2=0
+ $Y2=0
cc_255 N_A_136_387#_c_269_n N_A_134_74#_c_730_n 0.00382546f $X=2.505 $Y=1.095
+ $X2=0 $Y2=0
cc_256 N_A_136_387#_c_269_n N_A_134_74#_c_735_n 0.020073f $X=2.505 $Y=1.095
+ $X2=0 $Y2=0
cc_257 N_A_136_387#_c_271_n N_A_518_74#_M1000_s 0.00259532f $X=2.67 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_258 N_A_136_387#_c_264_n N_A_518_74#_c_754_n 0.00137075f $X=3.365 $Y=1.605
+ $X2=0 $Y2=0
cc_259 N_A_136_387#_c_271_n N_A_518_74#_c_754_n 0.0139685f $X=2.67 $Y=1.095
+ $X2=0 $Y2=0
cc_260 N_A_136_387#_M1000_g N_A_518_74#_c_755_n 0.0144222f $X=2.95 $Y=0.74 $X2=0
+ $Y2=0
cc_261 N_A_136_387#_M1006_g N_A_518_74#_c_755_n 0.0131461f $X=3.38 $Y=0.74 $X2=0
+ $Y2=0
cc_262 N_B1_M1010_g N_B2_c_451_n 0.0307135f $X=3.84 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_263 N_B1_M1004_g N_B2_M1005_g 0.0361308f $X=3.905 $Y=2.4 $X2=0 $Y2=0
cc_264 N_B1_c_366_n N_B2_M1005_g 8.48493e-19 $X=3.86 $Y=1.515 $X2=0 $Y2=0
cc_265 N_B1_c_374_n N_B2_M1005_g 0.0140695f $X=4.925 $Y=1.805 $X2=0 $Y2=0
cc_266 N_B1_M1013_g N_B2_M1009_g 0.0167293f $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_267 N_B1_c_374_n N_B2_M1009_g 0.021404f $X=4.925 $Y=1.805 $X2=0 $Y2=0
cc_268 N_B1_M1017_g N_B2_c_454_n 0.0337897f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_269 N_B1_M1010_g B2 8.65119e-19 $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_270 N_B1_M1017_g B2 5.30633e-19 $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_271 N_B1_c_366_n B2 0.0090454f $X=3.86 $Y=1.515 $X2=0 $Y2=0
cc_272 N_B1_c_367_n B2 6.51756e-19 $X=3.86 $Y=1.515 $X2=0 $Y2=0
cc_273 N_B1_c_374_n B2 0.0246222f $X=4.925 $Y=1.805 $X2=0 $Y2=0
cc_274 B1 B2 0.0124556f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_275 N_B1_c_366_n N_B2_c_456_n 0.00172432f $X=3.86 $Y=1.515 $X2=0 $Y2=0
cc_276 N_B1_c_367_n N_B2_c_456_n 0.0183886f $X=3.86 $Y=1.515 $X2=0 $Y2=0
cc_277 N_B1_c_374_n N_B2_c_456_n 6.34453e-19 $X=4.925 $Y=1.805 $X2=0 $Y2=0
cc_278 B1 N_B2_c_456_n 0.0075901f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_279 N_B1_c_369_n N_B2_c_456_n 0.0167293f $X=5.33 $Y=1.515 $X2=0 $Y2=0
cc_280 N_B1_c_375_n N_VPWR_M1016_s 0.00132909f $X=4.025 $Y=1.805 $X2=0 $Y2=0
cc_281 N_B1_M1004_g N_VPWR_c_513_n 0.0014841f $X=3.905 $Y=2.4 $X2=0 $Y2=0
cc_282 N_B1_M1013_g N_VPWR_c_515_n 0.00330306f $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_283 B1 N_VPWR_c_515_n 0.00852165f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_284 N_B1_c_369_n N_VPWR_c_515_n 5.93922e-19 $X=5.33 $Y=1.515 $X2=0 $Y2=0
cc_285 N_B1_M1004_g N_VPWR_c_518_n 0.00517089f $X=3.905 $Y=2.4 $X2=0 $Y2=0
cc_286 N_B1_M1013_g N_VPWR_c_518_n 0.00517089f $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_287 N_B1_M1004_g N_VPWR_c_507_n 0.0097793f $X=3.905 $Y=2.4 $X2=0 $Y2=0
cc_288 N_B1_M1013_g N_VPWR_c_507_n 0.0098133f $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_289 N_B1_c_374_n N_Y_M1005_d 0.00165831f $X=4.925 $Y=1.805 $X2=0 $Y2=0
cc_290 N_B1_M1004_g N_Y_c_587_n 6.29912e-19 $X=3.905 $Y=2.4 $X2=0 $Y2=0
cc_291 N_B1_M1004_g N_Y_c_593_n 0.0166787f $X=3.905 $Y=2.4 $X2=0 $Y2=0
cc_292 N_B1_c_367_n N_Y_c_593_n 4.27666e-19 $X=3.86 $Y=1.515 $X2=0 $Y2=0
cc_293 N_B1_c_374_n N_Y_c_593_n 0.0234974f $X=4.925 $Y=1.805 $X2=0 $Y2=0
cc_294 N_B1_c_375_n N_Y_c_593_n 0.0184822f $X=4.025 $Y=1.805 $X2=0 $Y2=0
cc_295 N_B1_c_374_n N_Y_c_608_n 0.0126843f $X=4.925 $Y=1.805 $X2=0 $Y2=0
cc_296 N_B1_M1010_g Y 2.22458e-19 $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_297 N_B1_M1004_g Y 9.48722e-19 $X=3.905 $Y=2.4 $X2=0 $Y2=0
cc_298 N_B1_c_366_n Y 0.0137607f $X=3.86 $Y=1.515 $X2=0 $Y2=0
cc_299 N_B1_c_367_n Y 9.46247e-19 $X=3.86 $Y=1.515 $X2=0 $Y2=0
cc_300 N_B1_c_375_n Y 0.00734143f $X=4.025 $Y=1.805 $X2=0 $Y2=0
cc_301 N_B1_c_374_n N_A_799_368#_M1004_d 0.00166235f $X=4.925 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_302 B1 N_A_799_368#_M1009_s 0.00222333f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_303 N_B1_M1004_g N_A_799_368#_c_634_n 0.00617601f $X=3.905 $Y=2.4 $X2=0 $Y2=0
cc_304 N_B1_M1013_g N_A_799_368#_c_630_n 0.00358808f $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_305 N_B1_M1004_g N_A_799_368#_c_631_n 0.00340097f $X=3.905 $Y=2.4 $X2=0 $Y2=0
cc_306 N_B1_M1013_g N_A_799_368#_c_637_n 0.0111002f $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_307 N_B1_c_374_n N_A_799_368#_c_637_n 0.00216696f $X=4.925 $Y=1.805 $X2=0
+ $Y2=0
cc_308 B1 N_A_799_368#_c_637_n 0.0167959f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_309 N_B1_M1010_g N_VGND_c_661_n 0.00293683f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_310 N_B1_M1017_g N_VGND_c_662_n 0.00981808f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_311 N_B1_M1010_g N_VGND_c_664_n 0.00430908f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_312 N_B1_M1017_g N_VGND_c_666_n 0.00383152f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_313 N_B1_M1010_g N_VGND_c_667_n 0.00445932f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_314 N_B1_M1017_g N_VGND_c_667_n 0.00372886f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_315 N_B1_M1010_g N_A_518_74#_c_755_n 0.00332495f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_316 N_B1_M1010_g N_A_518_74#_c_767_n 0.00642991f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_317 N_B1_M1010_g N_A_518_74#_c_768_n 0.00963801f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_318 N_B1_c_366_n N_A_518_74#_c_768_n 0.00900162f $X=3.86 $Y=1.515 $X2=0 $Y2=0
cc_319 N_B1_c_367_n N_A_518_74#_c_768_n 4.87923e-19 $X=3.86 $Y=1.515 $X2=0 $Y2=0
cc_320 N_B1_M1010_g N_A_518_74#_c_757_n 0.00333924f $X=3.84 $Y=0.74 $X2=0 $Y2=0
cc_321 N_B1_c_366_n N_A_518_74#_c_757_n 0.00667011f $X=3.86 $Y=1.515 $X2=0 $Y2=0
cc_322 N_B1_c_367_n N_A_518_74#_c_757_n 5.28989e-19 $X=3.86 $Y=1.515 $X2=0 $Y2=0
cc_323 N_B1_M1017_g N_A_518_74#_c_774_n 0.0107539f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_324 B1 N_A_518_74#_c_774_n 0.0167053f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_325 N_B1_M1017_g N_A_518_74#_c_759_n 0.00412046f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_326 B1 N_A_518_74#_c_759_n 0.0124005f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_327 N_B1_c_369_n N_A_518_74#_c_759_n 0.00115984f $X=5.33 $Y=1.515 $X2=0 $Y2=0
cc_328 N_B1_M1017_g N_A_518_74#_c_760_n 0.00130587f $X=5.265 $Y=0.74 $X2=0 $Y2=0
cc_329 N_B2_M1005_g N_VPWR_c_518_n 0.00333896f $X=4.355 $Y=2.4 $X2=0 $Y2=0
cc_330 N_B2_M1009_g N_VPWR_c_518_n 0.00333896f $X=4.805 $Y=2.4 $X2=0 $Y2=0
cc_331 N_B2_M1005_g N_VPWR_c_507_n 0.00422796f $X=4.355 $Y=2.4 $X2=0 $Y2=0
cc_332 N_B2_M1009_g N_VPWR_c_507_n 0.00422796f $X=4.805 $Y=2.4 $X2=0 $Y2=0
cc_333 N_B2_M1005_g N_Y_c_593_n 0.0119021f $X=4.355 $Y=2.4 $X2=0 $Y2=0
cc_334 N_B2_M1005_g N_A_799_368#_c_634_n 0.00738921f $X=4.355 $Y=2.4 $X2=0 $Y2=0
cc_335 N_B2_M1009_g N_A_799_368#_c_634_n 5.23376e-19 $X=4.805 $Y=2.4 $X2=0 $Y2=0
cc_336 N_B2_M1005_g N_A_799_368#_c_630_n 0.00936332f $X=4.355 $Y=2.4 $X2=0 $Y2=0
cc_337 N_B2_M1009_g N_A_799_368#_c_630_n 0.0135505f $X=4.805 $Y=2.4 $X2=0 $Y2=0
cc_338 N_B2_M1005_g N_A_799_368#_c_631_n 0.00191106f $X=4.355 $Y=2.4 $X2=0 $Y2=0
cc_339 N_B2_M1005_g N_A_799_368#_c_637_n 5.69844e-19 $X=4.355 $Y=2.4 $X2=0 $Y2=0
cc_340 N_B2_M1009_g N_A_799_368#_c_637_n 0.0111705f $X=4.805 $Y=2.4 $X2=0 $Y2=0
cc_341 N_B2_c_451_n N_VGND_c_661_n 0.00773369f $X=4.34 $Y=1.22 $X2=0 $Y2=0
cc_342 N_B2_c_454_n N_VGND_c_661_n 4.19327e-19 $X=4.82 $Y=1.22 $X2=0 $Y2=0
cc_343 N_B2_c_451_n N_VGND_c_662_n 4.00885e-19 $X=4.34 $Y=1.22 $X2=0 $Y2=0
cc_344 N_B2_c_454_n N_VGND_c_662_n 0.00702777f $X=4.82 $Y=1.22 $X2=0 $Y2=0
cc_345 N_B2_c_451_n N_VGND_c_665_n 0.00383152f $X=4.34 $Y=1.22 $X2=0 $Y2=0
cc_346 N_B2_c_454_n N_VGND_c_665_n 0.00383152f $X=4.82 $Y=1.22 $X2=0 $Y2=0
cc_347 N_B2_c_451_n N_VGND_c_667_n 0.00384446f $X=4.34 $Y=1.22 $X2=0 $Y2=0
cc_348 N_B2_c_454_n N_VGND_c_667_n 0.00369749f $X=4.82 $Y=1.22 $X2=0 $Y2=0
cc_349 N_B2_c_451_n N_A_518_74#_c_767_n 6.25243e-19 $X=4.34 $Y=1.22 $X2=0 $Y2=0
cc_350 N_B2_c_451_n N_A_518_74#_c_768_n 0.0124209f $X=4.34 $Y=1.22 $X2=0 $Y2=0
cc_351 B2 N_A_518_74#_c_768_n 0.00730648f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_352 N_B2_c_451_n N_A_518_74#_c_757_n 5.68029e-19 $X=4.34 $Y=1.22 $X2=0 $Y2=0
cc_353 N_B2_c_451_n N_A_518_74#_c_758_n 2.53282e-19 $X=4.34 $Y=1.22 $X2=0 $Y2=0
cc_354 N_B2_c_454_n N_A_518_74#_c_758_n 2.53282e-19 $X=4.82 $Y=1.22 $X2=0 $Y2=0
cc_355 N_B2_c_454_n N_A_518_74#_c_774_n 0.0162195f $X=4.82 $Y=1.22 $X2=0 $Y2=0
cc_356 N_B2_c_454_n N_A_518_74#_c_759_n 5.82428e-19 $X=4.82 $Y=1.22 $X2=0 $Y2=0
cc_357 B2 N_A_518_74#_c_788_n 0.0177874f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_358 N_B2_c_456_n N_A_518_74#_c_788_n 0.00105185f $X=4.82 $Y=1.385 $X2=0 $Y2=0
cc_359 N_VPWR_c_512_n N_Y_c_587_n 0.0289149f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_360 N_VPWR_c_513_n N_Y_c_587_n 0.0220702f $X=3.625 $Y=2.485 $X2=0 $Y2=0
cc_361 N_VPWR_c_517_n N_Y_c_587_n 0.0125859f $X=3.46 $Y=3.33 $X2=0 $Y2=0
cc_362 N_VPWR_c_507_n N_Y_c_587_n 0.0103846f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_363 N_VPWR_M1016_s N_Y_c_593_n 0.0101591f $X=3.455 $Y=1.84 $X2=0 $Y2=0
cc_364 N_VPWR_c_513_n N_Y_c_593_n 0.0200142f $X=3.625 $Y=2.485 $X2=0 $Y2=0
cc_365 N_VPWR_c_512_n Y 0.0097785f $X=2.67 $Y=1.985 $X2=0 $Y2=0
cc_366 N_VPWR_c_515_n N_A_799_368#_c_630_n 0.0103534f $X=5.48 $Y=2.115 $X2=0
+ $Y2=0
cc_367 N_VPWR_c_518_n N_A_799_368#_c_630_n 0.0592384f $X=5.395 $Y=3.33 $X2=0
+ $Y2=0
cc_368 N_VPWR_c_507_n N_A_799_368#_c_630_n 0.0326137f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_369 N_VPWR_c_513_n N_A_799_368#_c_631_n 0.011661f $X=3.625 $Y=2.485 $X2=0
+ $Y2=0
cc_370 N_VPWR_c_518_n N_A_799_368#_c_631_n 0.0234328f $X=5.395 $Y=3.33 $X2=0
+ $Y2=0
cc_371 N_VPWR_c_507_n N_A_799_368#_c_631_n 0.0125526f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_372 N_Y_c_593_n N_A_799_368#_M1004_d 0.00332066f $X=4.465 $Y=2.145 $X2=-0.19
+ $Y2=-0.245
cc_373 N_Y_c_593_n N_A_799_368#_c_634_n 0.0170155f $X=4.465 $Y=2.145 $X2=0 $Y2=0
cc_374 N_Y_M1005_d N_A_799_368#_c_630_n 0.00165831f $X=4.445 $Y=1.84 $X2=0 $Y2=0
cc_375 N_Y_c_593_n N_A_799_368#_c_630_n 0.00318644f $X=4.465 $Y=2.145 $X2=0
+ $Y2=0
cc_376 N_Y_c_608_n N_A_799_368#_c_630_n 0.0118669f $X=4.58 $Y=2.225 $X2=0 $Y2=0
cc_377 N_Y_M1000_d N_A_518_74#_c_755_n 0.00176461f $X=3.025 $Y=0.37 $X2=0 $Y2=0
cc_378 Y N_A_518_74#_c_755_n 0.0143448f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_379 Y N_A_518_74#_c_757_n 0.00157293f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_380 N_VGND_c_660_n N_A_134_74#_c_730_n 0.0117551f $X=2.175 $Y=0.66 $X2=0
+ $Y2=0
cc_381 N_VGND_c_663_n N_A_134_74#_c_730_n 0.0613668f $X=2.08 $Y=0 $X2=0 $Y2=0
cc_382 N_VGND_c_667_n N_A_134_74#_c_730_n 0.0341446f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_383 N_VGND_c_659_n N_A_134_74#_c_731_n 0.011924f $X=0.31 $Y=0.515 $X2=0 $Y2=0
cc_384 N_VGND_c_663_n N_A_134_74#_c_731_n 0.0234809f $X=2.08 $Y=0 $X2=0 $Y2=0
cc_385 N_VGND_c_667_n N_A_134_74#_c_731_n 0.0126009f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_386 N_VGND_c_660_n N_A_518_74#_c_754_n 0.025902f $X=2.175 $Y=0.66 $X2=0 $Y2=0
cc_387 N_VGND_c_661_n N_A_518_74#_c_755_n 0.011924f $X=4.125 $Y=0.55 $X2=0 $Y2=0
cc_388 N_VGND_c_664_n N_A_518_74#_c_755_n 0.0638649f $X=3.96 $Y=0 $X2=0 $Y2=0
cc_389 N_VGND_c_667_n N_A_518_74#_c_755_n 0.0354046f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_390 N_VGND_c_660_n N_A_518_74#_c_756_n 0.0119579f $X=2.175 $Y=0.66 $X2=0
+ $Y2=0
cc_391 N_VGND_c_664_n N_A_518_74#_c_756_n 0.0176866f $X=3.96 $Y=0 $X2=0 $Y2=0
cc_392 N_VGND_c_667_n N_A_518_74#_c_756_n 0.00967523f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_393 N_VGND_M1010_s N_A_518_74#_c_768_n 0.0101164f $X=3.915 $Y=0.37 $X2=0
+ $Y2=0
cc_394 N_VGND_c_661_n N_A_518_74#_c_768_n 0.0205261f $X=4.125 $Y=0.55 $X2=0
+ $Y2=0
cc_395 N_VGND_c_667_n N_A_518_74#_c_768_n 0.0113542f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_396 N_VGND_c_661_n N_A_518_74#_c_758_n 0.0121832f $X=4.125 $Y=0.55 $X2=0
+ $Y2=0
cc_397 N_VGND_c_662_n N_A_518_74#_c_758_n 0.0097355f $X=5.04 $Y=0.515 $X2=0
+ $Y2=0
cc_398 N_VGND_c_665_n N_A_518_74#_c_758_n 0.00970617f $X=4.87 $Y=0 $X2=0 $Y2=0
cc_399 N_VGND_c_667_n N_A_518_74#_c_758_n 0.00804326f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_400 N_VGND_M1015_d N_A_518_74#_c_774_n 0.00460082f $X=4.895 $Y=0.37 $X2=0
+ $Y2=0
cc_401 N_VGND_c_662_n N_A_518_74#_c_774_n 0.0181964f $X=5.04 $Y=0.515 $X2=0
+ $Y2=0
cc_402 N_VGND_c_667_n N_A_518_74#_c_774_n 0.0101909f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_403 N_VGND_c_667_n N_A_518_74#_c_759_n 0.00293094f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_404 N_VGND_c_662_n N_A_518_74#_c_760_n 0.00974948f $X=5.04 $Y=0.515 $X2=0
+ $Y2=0
cc_405 N_VGND_c_666_n N_A_518_74#_c_760_n 0.011066f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_406 N_VGND_c_667_n N_A_518_74#_c_760_n 0.00915947f $X=5.52 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__nand3_4.spice
* Created: Wed Sep  2 12:13:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nand3_4.pex.spice"
.subckt sky130_fd_sc_ms__nand3_4  VNB VPB A B C VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1007 N_Y_M1007_d N_A_M1007_g N_A_27_82#_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.19525 PD=1.02 PS=2.03 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1014 N_Y_M1007_d N_A_M1014_g N_A_27_82#_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1015 N_Y_M1015_d N_A_M1015_g N_A_27_82#_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1017 N_Y_M1015_d N_A_M1017_g N_A_27_82#_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1002 N_A_27_82#_M1017_s N_B_M1002_g N_A_456_82#_M1002_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.9 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1003 N_A_27_82#_M1003_d N_B_M1003_g N_A_456_82#_M1002_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.3 SB=75001 A=0.111 P=1.78 MULT=1
MM1012 N_A_27_82#_M1003_d N_B_M1012_g N_A_456_82#_M1012_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.8 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1016 N_A_27_82#_M1016_d N_B_M1016_g N_A_456_82#_M1012_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.19525 AS=0.1036 PD=2.03 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_456_82#_M1000_d N_C_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2035 PD=1.02 PS=2.03 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1001 N_A_456_82#_M1000_d N_C_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1009 N_A_456_82#_M1009_d N_C_M1009_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1013 N_A_456_82#_M1009_d N_C_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2035 PD=1.02 PS=2.03 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12 AD=0.4424
+ AS=0.3136 PD=1.91 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2 SB=90005.1
+ A=0.2016 P=2.6 MULT=1
MM1006 N_Y_M1005_d N_A_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12 AD=0.4424
+ AS=0.1792 PD=1.91 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.2 SB=90004.1
+ A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1004_d N_B_M1004_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.7 SB=90003.6
+ A=0.2016 P=2.6 MULT=1
MM1008 N_Y_M1004_d N_B_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.7252 PD=1.39 PS=2.415 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.1 SB=90003.1
+ A=0.2016 P=2.6 MULT=1
MM1010 N_Y_M1010_d N_C_M1010_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.7252 PD=1.39 PS=2.415 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.6 SB=90001.7
+ A=0.2016 P=2.6 MULT=1
MM1011 N_Y_M1010_d N_C_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=1.4672 PD=1.39 PS=4.86 NRD=0 NRS=0 M=1 R=6.22222 SA=90004 SB=90001.2
+ A=0.2016 P=2.6 MULT=1
DX18_noxref VNB VPB NWDIODE A=12.3132 P=16.96
*
.include "sky130_fd_sc_ms__nand3_4.pxi.spice"
*
.ends
*
*

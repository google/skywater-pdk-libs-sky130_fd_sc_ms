* NGSPICE file created from sky130_fd_sc_ms__a2111oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 VGND C1 Y VNB nlowvt w=740000u l=150000u
+  ad=7.141e+11p pd=6.37e+06u as=6.919e+11p ps=6.31e+06u
M1001 a_722_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=5.994e+11p pd=6.06e+06u as=0p ps=0u
M1002 a_533_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.1872e+12p pd=1.108e+07u as=6.048e+11p ps=5.56e+06u
M1003 Y D1 a_69_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=8.848e+11p ps=8.3e+06u
M1004 a_69_368# D1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_722_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_337_368# C1 a_69_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1007 Y D1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_69_368# C1 a_337_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_337_368# B1 a_533_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_533_368# B1 a_337_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A1 a_533_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A2 a_722_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y A1 a_722_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_533_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A2 a_533_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


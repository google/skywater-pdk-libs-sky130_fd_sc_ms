* File: sky130_fd_sc_ms__inv_4.pex.spice
* Created: Fri Aug 28 17:38:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__INV_4%A 3 7 11 15 19 23 27 31 33 34 35 36 55
r76 54 55 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.89 $Y=1.515
+ $X2=1.905 $Y2=1.515
r77 52 54 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=1.635 $Y=1.515
+ $X2=1.89 $Y2=1.515
r78 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.635
+ $Y=1.515 $X2=1.635 $Y2=1.515
r79 50 52 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=1.475 $Y=1.515
+ $X2=1.635 $Y2=1.515
r80 49 50 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=1.44 $Y=1.515
+ $X2=1.475 $Y2=1.515
r81 48 49 77.8133 $w=3.3e-07 $l=4.45e-07 $layer=POLY_cond $X=0.995 $Y=1.515
+ $X2=1.44 $Y2=1.515
r82 47 48 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=0.99 $Y=1.515
+ $X2=0.995 $Y2=1.515
r83 45 47 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=0.615 $Y=1.515
+ $X2=0.99 $Y2=1.515
r84 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.615
+ $Y=1.515 $X2=0.615 $Y2=1.515
r85 43 45 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.54 $Y=1.515
+ $X2=0.615 $Y2=1.515
r86 41 43 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.525 $Y=1.515
+ $X2=0.54 $Y2=1.515
r87 36 53 1.20605 $w=4.28e-07 $l=4.5e-08 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.635 $Y2=1.565
r88 35 53 11.6584 $w=4.28e-07 $l=4.35e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.635 $Y2=1.565
r89 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r90 34 46 2.81411 $w=4.28e-07 $l=1.05e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.615 $Y2=1.565
r91 33 46 10.0504 $w=4.28e-07 $l=3.75e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.615 $Y2=1.565
r92 29 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.35
+ $X2=1.905 $Y2=1.515
r93 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.905 $Y=1.35
+ $X2=1.905 $Y2=0.74
r94 25 54 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=1.68
+ $X2=1.89 $Y2=1.515
r95 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.89 $Y=1.68
+ $X2=1.89 $Y2=2.4
r96 21 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.475 $Y=1.35
+ $X2=1.475 $Y2=1.515
r97 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.475 $Y=1.35
+ $X2=1.475 $Y2=0.74
r98 17 49 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.44 $Y=1.68
+ $X2=1.44 $Y2=1.515
r99 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.44 $Y=1.68
+ $X2=1.44 $Y2=2.4
r100 13 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=1.515
r101 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=0.74
r102 9 47 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=1.68
+ $X2=0.99 $Y2=1.515
r103 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.99 $Y=1.68
+ $X2=0.99 $Y2=2.4
r104 5 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.68
+ $X2=0.54 $Y2=1.515
r105 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.54 $Y=1.68 $X2=0.54
+ $Y2=2.4
r106 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.35
+ $X2=0.525 $Y2=1.515
r107 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.525 $Y=1.35
+ $X2=0.525 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__INV_4%VPWR 1 2 3 10 12 16 20 22 24 26 28 37 41
r36 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r38 32 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r40 29 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=3.33 $X2=1.215
+ $Y2=3.33
r41 29 31 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.3 $Y=3.33 $X2=1.68
+ $Y2=3.33
r42 28 40 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.03 $Y=3.33
+ $X2=2.215 $Y2=3.33
r43 28 31 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.03 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 26 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r46 26 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r47 22 40 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=2.155 $Y=3.245
+ $X2=2.215 $Y2=3.33
r48 22 24 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=2.155 $Y=3.245
+ $X2=2.155 $Y2=2.455
r49 18 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=3.245
+ $X2=1.215 $Y2=3.33
r50 18 20 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.215 $Y=3.245
+ $X2=1.215 $Y2=2.455
r51 17 34 3.96842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.4 $Y=3.33 $X2=0.2
+ $Y2=3.33
r52 16 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=3.33
+ $X2=1.215 $Y2=3.33
r53 16 17 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.13 $Y=3.33 $X2=0.4
+ $Y2=3.33
r54 12 15 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=0.275 $Y=2.115
+ $X2=0.275 $Y2=2.815
r55 10 34 3.17474 $w=2.5e-07 $l=1.16619e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.2 $Y2=3.33
r56 10 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.275 $Y2=2.815
r57 3 24 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.98
+ $Y=1.84 $X2=2.115 $Y2=2.455
r58 2 20 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.08
+ $Y=1.84 $X2=1.215 $Y2=2.455
r59 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.17
+ $Y=1.84 $X2=0.315 $Y2=2.815
r60 1 12 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.17
+ $Y=1.84 $X2=0.315 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__INV_4%Y 1 2 3 4 13 15 19 21 22 23 27 31 33 35 40 41
+ 44
r73 43 44 32.8196 $w=2.28e-07 $l=6.55e-07 $layer=LI1_cond $X=2.16 $Y=1.95
+ $X2=2.16 $Y2=1.295
r74 42 44 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.16 $Y=1.18
+ $X2=2.16 $Y2=1.295
r75 36 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.83 $Y=2.035
+ $X2=1.665 $Y2=2.035
r76 35 43 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.045 $Y=2.035
+ $X2=2.16 $Y2=1.95
r77 35 36 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.045 $Y=2.035
+ $X2=1.83 $Y2=2.035
r78 34 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.775 $Y=1.095
+ $X2=1.69 $Y2=1.095
r79 33 42 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.045 $Y=1.095
+ $X2=2.16 $Y2=1.18
r80 33 34 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.045 $Y=1.095
+ $X2=1.775 $Y2=1.095
r81 29 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.69 $Y=1.01 $X2=1.69
+ $Y2=1.095
r82 29 31 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.69 $Y=1.01
+ $X2=1.69 $Y2=0.515
r83 25 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=2.12
+ $X2=1.665 $Y2=2.035
r84 25 27 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.665 $Y=2.12
+ $X2=1.665 $Y2=2.815
r85 24 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.93 $Y=2.035
+ $X2=0.765 $Y2=2.035
r86 23 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.5 $Y=2.035
+ $X2=1.665 $Y2=2.035
r87 23 24 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.5 $Y=2.035
+ $X2=0.93 $Y2=2.035
r88 21 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=1.095
+ $X2=1.69 $Y2=1.095
r89 21 22 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.605 $Y=1.095
+ $X2=0.865 $Y2=1.095
r90 17 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.74 $Y=1.01
+ $X2=0.865 $Y2=1.095
r91 17 19 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.74 $Y=1.01
+ $X2=0.74 $Y2=0.515
r92 13 38 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=2.12
+ $X2=0.765 $Y2=2.035
r93 13 15 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.765 $Y=2.12
+ $X2=0.765 $Y2=2.815
r94 4 40 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.84 $X2=1.665 $Y2=2.115
r95 4 27 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.84 $X2=1.665 $Y2=2.815
r96 3 38 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.84 $X2=0.765 $Y2=2.115
r97 3 15 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.84 $X2=0.765 $Y2=2.815
r98 2 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.55
+ $Y=0.37 $X2=1.69 $Y2=0.515
r99 1 19 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=0.6
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__INV_4%VGND 1 2 3 10 12 16 18 20 22 24 29 38 42
r37 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r38 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r39 33 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r40 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r41 30 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.21
+ $Y2=0
r42 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.68
+ $Y2=0
r43 29 41 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=1.955 $Y=0 $X2=2.177
+ $Y2=0
r44 29 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.955 $Y=0 $X2=1.68
+ $Y2=0
r45 28 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r46 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r47 25 35 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r48 25 27 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r49 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.21
+ $Y2=0
r50 24 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=0.72
+ $Y2=0
r51 22 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r52 22 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r53 22 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 18 41 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=2.12 $Y=0.085
+ $X2=2.177 $Y2=0
r55 18 20 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=2.12 $Y=0.085
+ $X2=2.12 $Y2=0.595
r56 14 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0
r57 14 16 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0.595
r58 10 35 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r59 10 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.515
r60 3 20 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=1.98
+ $Y=0.37 $X2=2.12 $Y2=0.595
r61 2 16 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.21 $Y2=0.595
r62 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends


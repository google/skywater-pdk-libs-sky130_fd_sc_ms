* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__maj3_2 A B C VGND VNB VPB VPWR X
X0 a_793_368# C a_87_264# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X1 a_87_264# B a_587_347# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X2 a_587_347# C VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X3 a_87_264# B a_577_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VPWR A a_793_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X5 a_413_74# B a_87_264# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_793_74# C a_87_264# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 X a_87_264# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 VGND a_87_264# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 VGND A a_413_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 VGND A a_793_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 VPWR A a_396_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X12 a_396_368# B a_87_264# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X13 a_577_74# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 X a_87_264# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 VPWR a_87_264# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
.ends

* File: sky130_fd_sc_ms__dlclkp_2.spice
* Created: Fri Aug 28 17:26:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dlclkp_2.pex.spice"
.subckt sky130_fd_sc_ms__dlclkp_2  VNB VPB GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* VPB	VPB
* VNB	VNB
MM1021 N_VGND_M1021_d N_A_83_244#_M1021_g N_A_27_74#_M1021_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.224467 AS=0.2109 PD=1.45319 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1014 A_267_74# N_GATE_M1014_g N_VGND_M1021_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.194133 PD=0.88 PS=1.25681 NRD=12.18 NRS=62.808 M=1 R=4.26667
+ SA=75001 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1013 N_A_83_244#_M1013_d N_A_315_48#_M1013_g A_267_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.184091 AS=0.0768 PD=1.49132 PS=0.88 NRD=22.488 NRS=12.18 M=1
+ R=4.26667 SA=75001.4 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1007 A_494_118# N_A_315_338#_M1007_g N_A_83_244#_M1013_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0774375 AS=0.120809 PD=0.85 PS=0.978679 NRD=36.96 NRS=55.704 M=1
+ R=2.8 SA=75002.1 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_27_74#_M1010_g A_494_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.125529 AS=0.0774375 PD=0.99569 PS=0.85 NRD=0 NRS=36.96 M=1 R=2.8 SA=75002
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1011 N_A_315_338#_M1011_d N_A_315_48#_M1011_g N_VGND_M1010_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.221171 PD=2.05 PS=1.75431 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_CLK_M1015_g N_A_315_48#_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1019 A_1044_119# N_CLK_M1019_g N_VGND_M1015_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.0777 AS=0.1295 PD=0.95 PS=1.09 NRD=8.1 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1017 N_A_1044_387#_M1017_d N_A_27_74#_M1017_g A_1044_119# VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.0777 PD=2.05 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333
+ SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_GCLK_M1003_d N_A_1044_387#_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.21835 PD=1.02 PS=2.21 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1009 N_GCLK_M1003_d N_A_1044_387#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_VPWR_M1004_d N_A_83_244#_M1004_g N_A_27_74#_M1004_s VPB PSHORT L=0.18
+ W=1.12 AD=0.311698 AS=0.3136 PD=1.77509 PS=2.8 NRD=25.4918 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90001.9 A=0.2016 P=2.6 MULT=1
MM1020 A_267_392# N_GATE_M1020_g N_VPWR_M1004_d VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.278302 PD=1.24 PS=1.58491 NRD=12.7853 NRS=26.5753 M=1 R=5.55556
+ SA=90000.9 SB=90001.4 A=0.18 P=2.36 MULT=1
MM1000 N_A_83_244#_M1000_d N_A_315_338#_M1000_g A_267_392# VPB PSHORT L=0.18 W=1
+ AD=0.285493 AS=0.12 PD=2.28169 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556
+ SA=90001.3 SB=90001 A=0.18 P=2.36 MULT=1
MM1002 A_511_508# N_A_315_48#_M1002_g N_A_83_244#_M1000_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.119907 PD=0.66 PS=0.95831 NRD=30.4759 NRS=0 M=1
+ R=2.33333 SA=90002.1 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1006 N_VPWR_M1006_d N_A_27_74#_M1006_g A_511_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.1092 AS=0.0504 PD=0.913333 PS=0.66 NRD=46.886 NRS=30.4759 M=1 R=2.33333
+ SA=90002.6 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1008 N_A_315_338#_M1008_d N_A_315_48#_M1008_g N_VPWR_M1006_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.2184 PD=2.24 PS=1.82667 NRD=0 NRS=35.1645 M=1 R=4.66667
+ SA=90001.7 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1012 N_VPWR_M1012_d N_CLK_M1012_g N_A_315_48#_M1012_s VPB PSHORT L=0.18 W=0.84
+ AD=0.142891 AS=0.252 PD=1.20978 PS=2.28 NRD=5.8509 NRS=3.5066 M=1 R=4.66667
+ SA=90000.2 SB=90002.7 A=0.1512 P=2.04 MULT=1
MM1001 N_A_1044_387#_M1001_d N_CLK_M1001_g N_VPWR_M1012_d VPB PSHORT L=0.18 W=1
+ AD=0.1475 AS=0.170109 PD=1.295 PS=1.44022 NRD=3.9203 NRS=3.9203 M=1 R=5.55556
+ SA=90000.6 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_A_27_74#_M1005_g N_A_1044_387#_M1001_d VPB PSHORT L=0.18
+ W=1 AD=0.458255 AS=0.1475 PD=1.9434 PS=1.295 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90001.1 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1016 N_GCLK_M1016_d N_A_1044_387#_M1016_g N_VPWR_M1005_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.513245 PD=1.39 PS=2.1766 NRD=0 NRS=4.3931 M=1 R=6.22222
+ SA=90002 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1018 N_GCLK_M1016_d N_A_1044_387#_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX22_noxref VNB VPB NWDIODE A=14.4324 P=20.08
*
.include "sky130_fd_sc_ms__dlclkp_2.pxi.spice"
*
.ends
*
*

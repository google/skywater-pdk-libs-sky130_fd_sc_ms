* File: sky130_fd_sc_ms__dlrtn_1.spice
* Created: Wed Sep  2 12:05:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dlrtn_1.pex.spice"
.subckt sky130_fd_sc_ms__dlrtn_1  VNB VPB D GATE_N RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1013 N_VGND_M1013_d N_D_M1013_g N_A_27_136#_M1013_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.171076 AS=0.15675 PD=1.27054 PS=1.67 NRD=55.86 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1000 N_A_232_98#_M1000_d N_GATE_N_M1000_g N_VGND_M1013_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1961 AS=0.230174 PD=2.01 PS=1.70946 NRD=0 NRS=41.52 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1016_d N_A_232_98#_M1016_g N_A_357_392#_M1016_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.426921 AS=0.2109 PD=2.06449 PS=2.05 NRD=84.624 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1010 A_681_74# N_A_27_136#_M1010_g N_VGND_M1016_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.369229 PD=0.88 PS=1.78551 NRD=12.18 NRS=15.936 M=1 R=4.26667
+ SA=75001.3 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1017 N_A_657_392#_M1017_d N_A_232_98#_M1017_g A_681_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.115623 AS=0.0768 PD=1.16528 PS=0.88 NRD=8.436 NRS=12.18 M=1
+ R=4.26667 SA=75001.7 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1003 A_854_74# N_A_357_392#_M1003_g N_A_657_392#_M1017_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.05775 AS=0.0758774 PD=0.695 PS=0.764717 NRD=23.568 NRS=0 M=1 R=2.8
+ SA=75002.1 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_897_406#_M1001_g A_854_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1239 AS=0.05775 PD=1.43 PS=0.695 NRD=1.428 NRS=23.568 M=1 R=2.8
+ SA=75002.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1014 A_1139_74# N_A_657_392#_M1014_g N_A_897_406#_M1014_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_RESET_B_M1008_g A_1139_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.163525 AS=0.0888 PD=1.185 PS=0.98 NRD=12.972 NRS=10.536 M=1 R=4.93333
+ SA=75000.6 SB=75000.9 A=0.111 P=1.78 MULT=1
MM1015 N_Q_M1015_d N_A_897_406#_M1015_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2701 AS=0.163525 PD=2.21 PS=1.185 NRD=12.972 NRS=12.972 M=1 R=4.93333
+ SA=75001.2 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1012 N_VPWR_M1012_d N_D_M1012_g N_A_27_136#_M1012_s VPB PSHORT L=0.18 W=0.84
+ AD=0.185525 AS=0.2352 PD=1.285 PS=2.24 NRD=18.7544 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1005 N_A_232_98#_M1005_d N_GATE_N_M1005_g N_VPWR_M1012_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.185525 PD=2.24 PS=1.285 NRD=0 NRS=18.7544 M=1 R=4.66667
+ SA=90000.8 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1009 N_VPWR_M1009_d N_A_232_98#_M1009_g N_A_357_392#_M1009_s VPB PSHORT L=0.18
+ W=0.84 AD=0.212602 AS=0.2352 PD=1.43348 PS=2.24 NRD=46.4526 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90002.3 A=0.1512 P=2.04 MULT=1
MM1004 A_573_392# N_A_27_136#_M1004_g N_VPWR_M1009_d VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.253098 PD=1.24 PS=1.70652 NRD=12.7853 NRS=16.7253 M=1 R=5.55556
+ SA=90000.7 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1018 N_A_657_392#_M1018_d N_A_357_392#_M1018_g A_573_392# VPB PSHORT L=0.18
+ W=1 AD=0.268732 AS=0.12 PD=2.1338 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556
+ SA=90001.1 SB=90001.4 A=0.18 P=2.36 MULT=1
MM1006 A_796_508# N_A_232_98#_M1006_g N_A_657_392#_M1018_d VPB PSHORT L=0.18
+ W=0.42 AD=0.10605 AS=0.112868 PD=0.925 PS=0.896197 NRD=92.6294 NRS=100.234 M=1
+ R=2.33333 SA=90001.7 SB=90002.4 A=0.0756 P=1.2 MULT=1
MM1007 N_VPWR_M1007_d N_A_897_406#_M1007_g A_796_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.125852 AS=0.10605 PD=1.09732 PS=0.925 NRD=0 NRS=92.6294 M=1 R=2.33333
+ SA=90002.4 SB=90001.7 A=0.0756 P=1.2 MULT=1
MM1019 N_A_897_406#_M1019_d N_A_657_392#_M1019_g N_VPWR_M1007_d VPB PSHORT
+ L=0.18 W=1 AD=0.22 AS=0.299648 PD=1.44 PS=2.61268 NRD=15.7403 NRS=0 M=1
+ R=5.55556 SA=90001.1 SB=90001.4 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1011_d N_RESET_B_M1011_g N_A_897_406#_M1019_d VPB PSHORT L=0.18
+ W=1 AD=0.209717 AS=0.22 PD=1.43868 PS=1.44 NRD=16.0752 NRS=15.7403 M=1
+ R=5.55556 SA=90001.8 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1002 N_Q_M1002_d N_A_897_406#_M1002_g N_VPWR_M1011_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.234883 PD=2.8 PS=1.61132 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90002.1 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX20_noxref VNB VPB NWDIODE A=14.0988 P=18.88
*
.include "sky130_fd_sc_ms__dlrtn_1.pxi.spice"
*
.ends
*
*

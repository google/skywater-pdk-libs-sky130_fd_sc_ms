* File: sky130_fd_sc_ms__or4_1.pex.spice
* Created: Fri Aug 28 18:08:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__OR4_1%D 3 5 7 8 12
c27 12 0 3.48794e-20 $X=0.485 $Y=1.585
r28 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.485
+ $Y=1.585 $X2=0.485 $Y2=1.585
r29 8 12 7.84301 $w=3.58e-07 $l=2.45e-07 $layer=LI1_cond $X=0.24 $Y=1.6
+ $X2=0.485 $Y2=1.6
r30 5 11 48.8089 $w=2.97e-07 $l=2.96606e-07 $layer=POLY_cond $X=0.59 $Y=1.84
+ $X2=0.5 $Y2=1.585
r31 5 7 166.022 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=0.59 $Y=1.84 $X2=0.59
+ $Y2=2.46
r32 1 11 38.5662 $w=2.97e-07 $l=1.94808e-07 $layer=POLY_cond $X=0.565 $Y=1.42
+ $X2=0.5 $Y2=1.585
r33 1 3 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=0.565 $Y=1.42
+ $X2=0.565 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__OR4_1%C 3 7 9 12
c33 7 0 6.19511e-20 $X=1.01 $Y=2.46
r34 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.585
+ $X2=1.085 $Y2=1.75
r35 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.585
+ $X2=1.085 $Y2=1.42
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.085
+ $Y=1.585 $X2=1.085 $Y2=1.585
r37 9 13 3.68142 $w=3.58e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.6 $X2=1.085
+ $Y2=1.6
r38 7 15 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=1.01 $Y=2.46 $X2=1.01
+ $Y2=1.75
r39 3 14 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=0.995 $Y=0.835
+ $X2=0.995 $Y2=1.42
.ends

.subckt PM_SKY130_FD_SC_MS__OR4_1%B 3 7 9 12
c33 9 0 1.43521e-19 $X=1.68 $Y=1.665
c34 3 0 8.7203e-20 $X=1.58 $Y=2.46
r35 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.655 $Y=1.585
+ $X2=1.655 $Y2=1.75
r36 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.655 $Y=1.585
+ $X2=1.655 $Y2=1.42
r37 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.655
+ $Y=1.585 $X2=1.655 $Y2=1.585
r38 7 14 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=1.73 $Y=0.835
+ $X2=1.73 $Y2=1.42
r39 3 15 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=1.58 $Y=2.46 $X2=1.58
+ $Y2=1.75
.ends

.subckt PM_SKY130_FD_SC_MS__OR4_1%A 3 7 9 15 16
c40 15 0 8.7203e-20 $X=2.225 $Y=1.515
c41 3 0 2.35487e-19 $X=2.15 $Y=2.46
r42 14 16 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=2.225 $Y=1.515
+ $X2=2.32 $Y2=1.515
r43 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.225
+ $Y=1.515 $X2=2.225 $Y2=1.515
r44 11 14 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.15 $Y=1.515
+ $X2=2.225 $Y2=1.515
r45 9 15 5.01062 $w=3.43e-07 $l=1.5e-07 $layer=LI1_cond $X=2.217 $Y=1.665
+ $X2=2.217 $Y2=1.515
r46 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.32 $Y=1.35
+ $X2=2.32 $Y2=1.515
r47 5 7 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=2.32 $Y=1.35 $X2=2.32
+ $Y2=0.835
r48 1 11 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.68
+ $X2=2.15 $Y2=1.515
r49 1 3 303.194 $w=1.8e-07 $l=7.8e-07 $layer=POLY_cond $X=2.15 $Y=1.68 $X2=2.15
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__OR4_1%A_44_392# 1 2 3 12 16 18 20 22 26 28 29 32 34
+ 36 37 40 44
c102 44 0 3.9013e-20 $X=2.77 $Y=1.465
r103 44 47 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.465
+ $X2=2.77 $Y2=1.63
r104 44 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.465
+ $X2=2.77 $Y2=1.3
r105 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.465 $X2=2.77 $Y2=1.465
r106 36 43 9.06394 $w=2.79e-07 $l=2.09893e-07 $layer=LI1_cond $X=2.645 $Y=1.63
+ $X2=2.747 $Y2=1.465
r107 36 37 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.645 $Y=1.63
+ $X2=2.645 $Y2=1.95
r108 35 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.19 $Y=1.095
+ $X2=2.025 $Y2=1.095
r109 34 43 16.1792 $w=2.79e-07 $l=4.53971e-07 $layer=LI1_cond $X=2.56 $Y=1.095
+ $X2=2.747 $Y2=1.465
r110 34 35 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.56 $Y=1.095
+ $X2=2.19 $Y2=1.095
r111 30 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=1.01
+ $X2=2.025 $Y2=1.095
r112 30 32 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=2.025 $Y=1.01
+ $X2=2.025 $Y2=0.835
r113 28 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.86 $Y=1.095
+ $X2=2.025 $Y2=1.095
r114 28 29 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=1.86 $Y=1.095
+ $X2=0.945 $Y2=1.095
r115 24 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.78 $Y=1.01
+ $X2=0.945 $Y2=1.095
r116 24 26 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=0.78 $Y=1.01
+ $X2=0.78 $Y2=0.835
r117 23 39 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.53 $Y=2.035
+ $X2=0.365 $Y2=2.035
r118 22 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.56 $Y=2.035
+ $X2=2.645 $Y2=1.95
r119 22 23 132.439 $w=1.68e-07 $l=2.03e-06 $layer=LI1_cond $X=2.56 $Y=2.035
+ $X2=0.53 $Y2=2.035
r120 18 39 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.365 $Y=2.12
+ $X2=0.365 $Y2=2.035
r121 18 20 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.365 $Y=2.12
+ $X2=0.365 $Y2=2.815
r122 16 46 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.83 $Y=0.74
+ $X2=2.83 $Y2=1.3
r123 12 47 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=2.84 $Y=2.4
+ $X2=2.84 $Y2=1.63
r124 3 39 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=0.22
+ $Y=1.96 $X2=0.365 $Y2=2.115
r125 3 20 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.22
+ $Y=1.96 $X2=0.365 $Y2=2.815
r126 2 32 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.56 $X2=2.025 $Y2=0.835
r127 1 26 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.64
+ $Y=0.56 $X2=0.78 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__OR4_1%VPWR 1 6 8 10 17 18 21
r27 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r28 18 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r29 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r30 15 21 10.0494 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=2.565 $Y=3.33
+ $X2=2.357 $Y2=3.33
r31 15 17 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.565 $Y=3.33
+ $X2=3.12 $Y2=3.33
r32 12 13 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 10 21 10.0494 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=2.15 $Y=3.33
+ $X2=2.357 $Y2=3.33
r34 10 12 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=2.15 $Y=3.33
+ $X2=0.24 $Y2=3.33
r35 8 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r36 8 13 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r37 4 21 1.57254 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.357 $Y=3.245
+ $X2=2.357 $Y2=3.33
r38 4 6 21.9381 $w=4.13e-07 $l=7.9e-07 $layer=LI1_cond $X=2.357 $Y=3.245
+ $X2=2.357 $Y2=2.455
r39 1 6 300 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=2 $X=2.24
+ $Y=1.96 $X2=2.375 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__OR4_1%X 1 2 9 13 14 15 16 23 32
c24 14 0 1.58051e-19 $X=3.035 $Y=1.95
r25 21 23 0.860491 $w=3.73e-07 $l=2.8e-08 $layer=LI1_cond $X=3.087 $Y=2.007
+ $X2=3.087 $Y2=2.035
r26 15 16 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=3.087 $Y=2.405
+ $X2=3.087 $Y2=2.775
r27 14 21 0.891223 $w=3.73e-07 $l=2.9e-08 $layer=LI1_cond $X=3.087 $Y=1.978
+ $X2=3.087 $Y2=2.007
r28 14 32 8.33934 $w=3.73e-07 $l=1.58e-07 $layer=LI1_cond $X=3.087 $Y=1.978
+ $X2=3.087 $Y2=1.82
r29 14 15 10.5103 $w=3.73e-07 $l=3.42e-07 $layer=LI1_cond $X=3.087 $Y=2.063
+ $X2=3.087 $Y2=2.405
r30 14 23 0.860491 $w=3.73e-07 $l=2.8e-08 $layer=LI1_cond $X=3.087 $Y=2.063
+ $X2=3.087 $Y2=2.035
r31 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.19 $Y=1.13 $X2=3.19
+ $Y2=1.82
r32 7 13 8.16989 $w=3.13e-07 $l=1.57e-07 $layer=LI1_cond $X=3.117 $Y=0.973
+ $X2=3.117 $Y2=1.13
r33 7 9 16.7562 $w=3.13e-07 $l=4.58e-07 $layer=LI1_cond $X=3.117 $Y=0.973
+ $X2=3.117 $Y2=0.515
r34 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.84 $X2=3.065 $Y2=1.985
r35 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.93
+ $Y=1.84 $X2=3.065 $Y2=2.815
r36 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.905
+ $Y=0.37 $X2=3.045 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR4_1%VGND 1 2 3 10 12 14 18 22 24 26 33 34 40 43
r46 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r47 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r48 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r49 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r50 34 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r51 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r52 31 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.78 $Y=0 $X2=2.615
+ $Y2=0
r53 31 33 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.78 $Y=0 $X2=3.12
+ $Y2=0
r54 30 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r55 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r56 27 40 10.9443 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=1.6 $Y=0 $X2=1.362
+ $Y2=0
r57 27 29 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.6 $Y=0 $X2=2.16
+ $Y2=0
r58 26 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.45 $Y=0 $X2=2.615
+ $Y2=0
r59 26 29 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.45 $Y=0 $X2=2.16
+ $Y2=0
r60 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r61 24 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r62 20 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=0.085
+ $X2=2.615 $Y2=0
r63 20 22 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=2.615 $Y=0.085
+ $X2=2.615 $Y2=0.675
r64 16 40 1.94084 $w=4.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.362 $Y=0.085
+ $X2=1.362 $Y2=0
r65 16 18 14.8566 $w=4.73e-07 $l=5.9e-07 $layer=LI1_cond $X=1.362 $Y=0.085
+ $X2=1.362 $Y2=0.675
r66 15 37 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r67 14 40 10.9443 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=1.125 $Y=0 $X2=1.362
+ $Y2=0
r68 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.125 $Y=0 $X2=0.445
+ $Y2=0
r69 10 37 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r70 10 12 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.835
r71 3 22 182 $w=1.7e-07 $l=2.71477e-07 $layer=licon1_NDIFF $count=1 $X=2.395
+ $Y=0.56 $X2=2.615 $Y2=0.675
r72 2 18 182 $w=1.7e-07 $l=3.4271e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.56 $X2=1.36 $Y2=0.675
r73 1 12 182 $w=1.7e-07 $l=3.67083e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.35 $Y2=0.835
.ends


* File: sky130_fd_sc_ms__a311o_4.pex.spice
* Created: Fri Aug 28 17:05:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A311O_4%C1 3 7 11 15 17 24
r60 24 25 8.33429 $w=3.47e-07 $l=6e-08 $layer=POLY_cond $X=1.145 $Y=1.62
+ $X2=1.205 $Y2=1.62
r61 23 24 51.3948 $w=3.47e-07 $l=3.7e-07 $layer=POLY_cond $X=0.775 $Y=1.62
+ $X2=1.145 $Y2=1.62
r62 22 23 11.1124 $w=3.47e-07 $l=8e-08 $layer=POLY_cond $X=0.695 $Y=1.62
+ $X2=0.775 $Y2=1.62
r63 20 22 4.86167 $w=3.47e-07 $l=3.5e-08 $layer=POLY_cond $X=0.66 $Y=1.62
+ $X2=0.695 $Y2=1.62
r64 17 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.66
+ $Y=1.635 $X2=0.66 $Y2=1.635
r65 13 25 22.4223 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.205 $Y=1.44
+ $X2=1.205 $Y2=1.62
r66 13 15 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.205 $Y=1.44
+ $X2=1.205 $Y2=0.73
r67 9 24 18.1053 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=1.145 $Y=1.8
+ $X2=1.145 $Y2=1.62
r68 9 11 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.145 $Y=1.8
+ $X2=1.145 $Y2=2.46
r69 5 23 22.4223 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.775 $Y=1.44
+ $X2=0.775 $Y2=1.62
r70 5 7 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.775 $Y=1.44
+ $X2=0.775 $Y2=0.73
r71 1 22 18.1053 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=0.695 $Y=1.8
+ $X2=0.695 $Y2=1.62
r72 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=0.695 $Y=1.8 $X2=0.695
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_4%B1 3 7 11 15 17 24
c60 3 0 1.44144e-19 $X=1.595 $Y=2.46
r61 24 25 2.93902 $w=3.28e-07 $l=2e-08 $layer=POLY_cond $X=2.045 $Y=1.635
+ $X2=2.065 $Y2=1.635
r62 22 24 50.6982 $w=3.28e-07 $l=3.45e-07 $layer=POLY_cond $X=1.7 $Y=1.635
+ $X2=2.045 $Y2=1.635
r63 20 22 9.55183 $w=3.28e-07 $l=6.5e-08 $layer=POLY_cond $X=1.635 $Y=1.635
+ $X2=1.7 $Y2=1.635
r64 19 20 5.87805 $w=3.28e-07 $l=4e-08 $layer=POLY_cond $X=1.595 $Y=1.635
+ $X2=1.635 $Y2=1.635
r65 17 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.7
+ $Y=1.635 $X2=1.7 $Y2=1.635
r66 13 25 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.065 $Y=1.47
+ $X2=2.065 $Y2=1.635
r67 13 15 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.065 $Y=1.47
+ $X2=2.065 $Y2=0.73
r68 9 24 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.045 $Y=1.8
+ $X2=2.045 $Y2=1.635
r69 9 11 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.045 $Y=1.8
+ $X2=2.045 $Y2=2.46
r70 5 20 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.635 $Y=1.47
+ $X2=1.635 $Y2=1.635
r71 5 7 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.635 $Y=1.47
+ $X2=1.635 $Y2=0.73
r72 1 19 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.595 $Y=1.8
+ $X2=1.595 $Y2=1.635
r73 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.595 $Y=1.8 $X2=1.595
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_4%A_157_392# 1 2 3 4 15 19 21 23 26 28 30 33
+ 35 37 38 40 42 45 48 49 53 56 60 63 64 65 67 71 73 76 78 82 94
c209 71 0 1.0161e-19 $X=1.08 $Y=2.105
c210 64 0 5.59968e-20 $X=5.545 $Y=2.035
c211 63 0 1.44209e-19 $X=4.56 $Y=1.95
c212 53 0 1.88456e-19 $X=1.85 $Y=0.555
c213 48 0 4.25334e-20 $X=1.08 $Y=2.02
c214 40 0 1.38345e-19 $X=4.365 $Y=1.75
c215 38 0 1.45634e-19 $X=4.275 $Y=1.675
r216 93 94 36.7053 $w=4.3e-07 $l=9e-08 $layer=POLY_cond $X=3.915 $Y=1.535
+ $X2=4.005 $Y2=1.535
r217 92 93 5.17352 $w=4.3e-07 $l=4e-08 $layer=POLY_cond $X=3.875 $Y=1.535
+ $X2=3.915 $Y2=1.535
r218 89 90 2.58676 $w=4.3e-07 $l=2e-08 $layer=POLY_cond $X=3.445 $Y=1.535
+ $X2=3.465 $Y2=1.535
r219 88 89 55.6154 $w=4.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.015 $Y=1.535
+ $X2=3.445 $Y2=1.535
r220 87 88 5.82021 $w=4.3e-07 $l=4.5e-08 $layer=POLY_cond $X=2.97 $Y=1.535
+ $X2=3.015 $Y2=1.535
r221 79 82 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=5.63 $Y=1.1
+ $X2=6.02 $Y2=1.1
r222 77 92 17.4606 $w=4.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.74 $Y=1.535
+ $X2=3.875 $Y2=1.535
r223 77 90 35.568 $w=4.3e-07 $l=2.75e-07 $layer=POLY_cond $X=3.74 $Y=1.535
+ $X2=3.465 $Y2=1.535
r224 76 78 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.74 $Y=1.485
+ $X2=3.905 $Y2=1.485
r225 76 77 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.74
+ $Y=1.485 $X2=3.74 $Y2=1.485
r226 69 71 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=0.92 $Y=2.105
+ $X2=1.08 $Y2=2.105
r227 66 79 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.63 $Y=1.265
+ $X2=5.63 $Y2=1.1
r228 66 67 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=5.63 $Y=1.265
+ $X2=5.63 $Y2=1.95
r229 64 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.545 $Y=2.035
+ $X2=5.63 $Y2=1.95
r230 64 65 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=5.545 $Y=2.035
+ $X2=4.645 $Y2=2.035
r231 63 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.56 $Y=1.95
+ $X2=4.645 $Y2=2.035
r232 62 63 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.56 $Y=1.65 $X2=4.56
+ $Y2=1.95
r233 60 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.475 $Y=1.565
+ $X2=4.56 $Y2=1.65
r234 60 78 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.475 $Y=1.565
+ $X2=3.905 $Y2=1.565
r235 59 87 32.3345 $w=4.3e-07 $l=2.5e-07 $layer=POLY_cond $X=2.72 $Y=1.535
+ $X2=2.97 $Y2=1.535
r236 59 84 23.2809 $w=4.3e-07 $l=1.8e-07 $layer=POLY_cond $X=2.72 $Y=1.535
+ $X2=2.54 $Y2=1.535
r237 58 76 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=2.72 $Y=1.485
+ $X2=3.74 $Y2=1.485
r238 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.72
+ $Y=1.485 $X2=2.72 $Y2=1.485
r239 56 58 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=2.325 $Y=1.485
+ $X2=2.72 $Y2=1.485
r240 51 56 17.4806 $w=3.35e-07 $l=6.33088e-07 $layer=LI1_cond $X=1.845 $Y=1.13
+ $X2=2.325 $Y2=1.485
r241 51 53 35.4293 $w=1.78e-07 $l=5.75e-07 $layer=LI1_cond $X=1.845 $Y=1.13
+ $X2=1.845 $Y2=0.555
r242 50 73 1.44715 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.165 $Y=1.215
+ $X2=1.035 $Y2=1.215
r243 49 51 6.23108 $w=3.35e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.755 $Y=1.215
+ $X2=1.845 $Y2=1.13
r244 49 50 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.755 $Y=1.215
+ $X2=1.165 $Y2=1.215
r245 48 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.08 $Y=2.02
+ $X2=1.08 $Y2=2.105
r246 47 73 5.04255 $w=1.75e-07 $l=1.05119e-07 $layer=LI1_cond $X=1.08 $Y=1.3
+ $X2=1.035 $Y2=1.215
r247 47 48 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.08 $Y=1.3
+ $X2=1.08 $Y2=2.02
r248 43 73 5.04255 $w=1.75e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.995 $Y=1.13
+ $X2=1.035 $Y2=1.215
r249 43 45 35.4293 $w=1.78e-07 $l=5.75e-07 $layer=LI1_cond $X=0.995 $Y=1.13
+ $X2=0.995 $Y2=0.555
r250 40 42 174.056 $w=1.8e-07 $l=6.5e-07 $layer=POLY_cond $X=4.365 $Y=1.75
+ $X2=4.365 $Y2=2.4
r251 38 40 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.275 $Y=1.675
+ $X2=4.365 $Y2=1.75
r252 38 94 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.275 $Y=1.675
+ $X2=4.005 $Y2=1.675
r253 35 93 23.194 $w=1.8e-07 $l=2.15e-07 $layer=POLY_cond $X=3.915 $Y=1.75
+ $X2=3.915 $Y2=1.535
r254 35 37 174.056 $w=1.8e-07 $l=6.5e-07 $layer=POLY_cond $X=3.915 $Y=1.75
+ $X2=3.915 $Y2=2.4
r255 31 92 27.6395 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=3.875 $Y=1.32
+ $X2=3.875 $Y2=1.535
r256 31 33 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=3.875 $Y=1.32
+ $X2=3.875 $Y2=0.795
r257 28 90 23.194 $w=1.8e-07 $l=2.15e-07 $layer=POLY_cond $X=3.465 $Y=1.75
+ $X2=3.465 $Y2=1.535
r258 28 30 174.056 $w=1.8e-07 $l=6.5e-07 $layer=POLY_cond $X=3.465 $Y=1.75
+ $X2=3.465 $Y2=2.4
r259 24 89 27.6395 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=3.445 $Y=1.32
+ $X2=3.445 $Y2=1.535
r260 24 26 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=3.445 $Y=1.32
+ $X2=3.445 $Y2=0.795
r261 21 88 23.194 $w=1.8e-07 $l=2.15e-07 $layer=POLY_cond $X=3.015 $Y=1.75
+ $X2=3.015 $Y2=1.535
r262 21 23 174.056 $w=1.8e-07 $l=6.5e-07 $layer=POLY_cond $X=3.015 $Y=1.75
+ $X2=3.015 $Y2=2.4
r263 17 87 27.6395 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=2.97 $Y=1.32
+ $X2=2.97 $Y2=1.535
r264 17 19 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.97 $Y=1.32
+ $X2=2.97 $Y2=0.78
r265 13 84 27.6395 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=2.54 $Y=1.32
+ $X2=2.54 $Y2=1.535
r266 13 15 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.54 $Y=1.32
+ $X2=2.54 $Y2=0.78
r267 4 69 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.785
+ $Y=1.96 $X2=0.92 $Y2=2.105
r268 3 82 182 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_NDIFF $count=1 $X=5.88
+ $Y=0.585 $X2=6.02 $Y2=1.1
r269 2 53 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.71
+ $Y=0.41 $X2=1.85 $Y2=0.555
r270 1 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.85
+ $Y=0.41 $X2=0.99 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_4%A3 1 3 4 5 6 8 11 15 17 22 23
c62 23 0 9.17238e-20 $X=5.13 $Y=1.585
r63 22 24 27.5429 $w=3.5e-07 $l=2e-07 $layer=POLY_cond $X=5.13 $Y=1.495 $X2=5.33
+ $Y2=1.495
r64 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.13
+ $Y=1.585 $X2=5.13 $Y2=1.585
r65 20 22 34.4286 $w=3.5e-07 $l=2.5e-07 $layer=POLY_cond $X=4.88 $Y=1.495
+ $X2=5.13 $Y2=1.495
r66 19 20 11.7057 $w=3.5e-07 $l=8.5e-08 $layer=POLY_cond $X=4.795 $Y=1.495
+ $X2=4.88 $Y2=1.495
r67 17 23 2.88111 $w=3.58e-07 $l=9e-08 $layer=LI1_cond $X=5.04 $Y=1.6 $X2=5.13
+ $Y2=1.6
r68 13 24 18.307 $w=1.8e-07 $l=2.55e-07 $layer=POLY_cond $X=5.33 $Y=1.75
+ $X2=5.33 $Y2=1.495
r69 13 15 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=5.33 $Y=1.75
+ $X2=5.33 $Y2=2.46
r70 9 20 18.307 $w=1.8e-07 $l=2.55e-07 $layer=POLY_cond $X=4.88 $Y=1.75 $X2=4.88
+ $Y2=1.495
r71 9 11 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=4.88 $Y=1.75 $X2=4.88
+ $Y2=2.46
r72 6 19 22.6286 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=4.795 $Y=1.24
+ $X2=4.795 $Y2=1.495
r73 6 8 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.795 $Y=1.24
+ $X2=4.795 $Y2=0.845
r74 4 19 26.3896 $w=3.5e-07 $l=2.14243e-07 $layer=POLY_cond $X=4.72 $Y=1.315
+ $X2=4.795 $Y2=1.495
r75 4 5 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.72 $Y=1.315 $X2=4.44
+ $Y2=1.315
r76 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.365 $Y=1.24
+ $X2=4.44 $Y2=1.315
r77 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.365 $Y=1.24
+ $X2=4.365 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_4%A1 3 7 11 15 17 18 19 29
c52 11 0 2.03712e-19 $X=6.23 $Y=2.46
c53 7 0 8.35615e-20 $X=5.805 $Y=0.905
c54 3 0 3.22225e-19 $X=5.78 $Y=2.46
r55 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.245
+ $Y=1.615 $X2=6.245 $Y2=1.615
r56 27 29 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=6.235 $Y=1.615
+ $X2=6.245 $Y2=1.615
r57 26 27 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=6.23 $Y=1.615
+ $X2=6.235 $Y2=1.615
r58 25 26 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=5.805 $Y=1.615
+ $X2=6.23 $Y2=1.615
r59 23 25 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=5.78 $Y=1.615
+ $X2=5.805 $Y2=1.615
r60 18 19 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.615
+ $X2=6.96 $Y2=1.615
r61 18 30 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=6.48 $Y=1.615
+ $X2=6.245 $Y2=1.615
r62 17 30 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=6 $Y=1.615
+ $X2=6.245 $Y2=1.615
r63 13 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.235 $Y=1.45
+ $X2=6.235 $Y2=1.615
r64 13 15 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=6.235 $Y=1.45
+ $X2=6.235 $Y2=0.905
r65 9 26 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.23 $Y=1.78
+ $X2=6.23 $Y2=1.615
r66 9 11 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=6.23 $Y=1.78 $X2=6.23
+ $Y2=2.46
r67 5 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.805 $Y=1.45
+ $X2=5.805 $Y2=1.615
r68 5 7 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=5.805 $Y=1.45
+ $X2=5.805 $Y2=0.905
r69 1 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.78 $Y=1.78
+ $X2=5.78 $Y2=1.615
r70 1 3 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=5.78 $Y=1.78 $X2=5.78
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_4%A2 3 7 11 15 17 22
c37 11 0 2.31472e-19 $X=7.16 $Y=2.46
c38 3 0 1.47716e-19 $X=6.71 $Y=2.46
r39 22 24 37.0769 $w=3.25e-07 $l=2.5e-07 $layer=POLY_cond $X=7.16 $Y=1.615
+ $X2=7.41 $Y2=1.615
r40 21 22 0.741538 $w=3.25e-07 $l=5e-09 $layer=POLY_cond $X=7.155 $Y=1.615
+ $X2=7.16 $Y2=1.615
r41 20 21 63.7723 $w=3.25e-07 $l=4.3e-07 $layer=POLY_cond $X=6.725 $Y=1.615
+ $X2=7.155 $Y2=1.615
r42 19 20 2.22462 $w=3.25e-07 $l=1.5e-08 $layer=POLY_cond $X=6.71 $Y=1.615
+ $X2=6.725 $Y2=1.615
r43 17 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.41
+ $Y=1.615 $X2=7.41 $Y2=1.615
r44 13 21 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.155 $Y=1.45
+ $X2=7.155 $Y2=1.615
r45 13 15 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=7.155 $Y=1.45
+ $X2=7.155 $Y2=0.905
r46 9 22 16.5763 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.16 $Y=1.78
+ $X2=7.16 $Y2=1.615
r47 9 11 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=7.16 $Y=1.78 $X2=7.16
+ $Y2=2.46
r48 5 20 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.725 $Y=1.45
+ $X2=6.725 $Y2=1.615
r49 5 7 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=6.725 $Y=1.45
+ $X2=6.725 $Y2=0.905
r50 1 19 16.5763 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.71 $Y=1.78
+ $X2=6.71 $Y2=1.615
r51 1 3 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=6.71 $Y=1.78 $X2=6.71
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_4%A_69_392# 1 2 3 14 18 19 21
r36 21 23 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.27 $Y=2.78
+ $X2=2.27 $Y2=2.99
r37 17 19 8.55446 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.37 $Y=2.887
+ $X2=1.535 $Y2=2.887
r38 17 18 5.8355 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.37 $Y=2.887
+ $X2=1.205 $Y2=2.887
r39 14 23 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.105 $Y=2.99
+ $X2=2.27 $Y2=2.99
r40 14 19 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.105 $Y=2.99
+ $X2=1.535 $Y2=2.99
r41 12 18 30.2516 $w=2.78e-07 $l=7.35e-07 $layer=LI1_cond $X=0.47 $Y=2.84
+ $X2=1.205 $Y2=2.84
r42 3 21 600 $w=1.7e-07 $l=8.84929e-07 $layer=licon1_PDIFF $count=1 $X=2.135
+ $Y=1.96 $X2=2.27 $Y2=2.78
r43 2 17 600 $w=1.7e-07 $l=9.04986e-07 $layer=licon1_PDIFF $count=1 $X=1.235
+ $Y=1.96 $X2=1.37 $Y2=2.8
r44 1 12 600 $w=1.7e-07 $l=9.00333e-07 $layer=licon1_PDIFF $count=1 $X=0.345
+ $Y=1.96 $X2=0.47 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_4%A_337_392# 1 2 3 4 13 17 19 23 25 27 29 31
+ 37
c69 37 0 2.28359e-19 $X=5.105 $Y=2.455
c70 29 0 2.95431e-19 $X=6.935 $Y=2.815
c71 27 0 8.37567e-20 $X=6.935 $Y=2.12
c72 23 0 2.95431e-19 $X=6.005 $Y=2.465
c73 19 0 8.44955e-20 $X=6.005 $Y=2.12
r74 31 34 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.82 $Y=2.405
+ $X2=1.82 $Y2=2.52
r75 27 42 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.935 $Y=2.12
+ $X2=6.935 $Y2=2.035
r76 27 29 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.935 $Y=2.12
+ $X2=6.935 $Y2=2.815
r77 26 39 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.09 $Y=2.035
+ $X2=6.005 $Y2=2.035
r78 25 42 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.85 $Y=2.035
+ $X2=6.935 $Y2=2.035
r79 25 26 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=6.85 $Y=2.035
+ $X2=6.09 $Y2=2.035
r80 21 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=2.46
+ $X2=6.005 $Y2=2.375
r81 21 23 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.005 $Y=2.46
+ $X2=6.005 $Y2=2.465
r82 20 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=2.29
+ $X2=6.005 $Y2=2.375
r83 19 39 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.005 $Y=2.12
+ $X2=6.005 $Y2=2.035
r84 19 20 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.005 $Y=2.12
+ $X2=6.005 $Y2=2.29
r85 18 37 8.61065 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=5.27 $Y=2.375
+ $X2=5.105 $Y2=2.39
r86 17 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=2.375
+ $X2=6.005 $Y2=2.375
r87 17 18 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.92 $Y=2.375
+ $X2=5.27 $Y2=2.375
r88 14 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.905 $Y=2.405
+ $X2=1.82 $Y2=2.405
r89 13 37 8.61065 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=4.94 $Y=2.405
+ $X2=5.105 $Y2=2.39
r90 13 14 198.005 $w=1.68e-07 $l=3.035e-06 $layer=LI1_cond $X=4.94 $Y=2.405
+ $X2=1.905 $Y2=2.405
r91 4 42 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=6.8
+ $Y=1.96 $X2=6.935 $Y2=2.115
r92 4 29 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.8
+ $Y=1.96 $X2=6.935 $Y2=2.815
r93 3 39 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=5.87
+ $Y=1.96 $X2=6.005 $Y2=2.115
r94 3 23 300 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_PDIFF $count=2 $X=5.87
+ $Y=1.96 $X2=6.005 $Y2=2.465
r95 2 37 300 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=2 $X=4.97
+ $Y=1.96 $X2=5.105 $Y2=2.455
r96 1 34 600 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=1 $X=1.685
+ $Y=1.96 $X2=1.82 $Y2=2.52
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_4%VPWR 1 2 3 4 5 6 21 23 27 31 33 37 41 43 45
+ 49 51 56 61 66 72 75 78 81 84 88
r109 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r110 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r111 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r112 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r113 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r114 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r115 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r116 72 73 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r117 70 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r118 70 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r119 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r120 67 84 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=6.65 $Y=3.33
+ $X2=6.47 $Y2=3.33
r121 67 69 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.65 $Y=3.33
+ $X2=6.96 $Y2=3.33
r122 66 87 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=7.22 $Y=3.33
+ $X2=7.45 $Y2=3.33
r123 66 69 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.22 $Y=3.33
+ $X2=6.96 $Y2=3.33
r124 65 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r125 65 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r126 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r127 62 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.72 $Y=3.33
+ $X2=5.595 $Y2=3.33
r128 62 64 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.72 $Y=3.33 $X2=6
+ $Y2=3.33
r129 61 84 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=6.29 $Y=3.33
+ $X2=6.47 $Y2=3.33
r130 61 64 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.29 $Y=3.33 $X2=6
+ $Y2=3.33
r131 60 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r132 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r133 57 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=3.69 $Y2=3.33
r134 57 59 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=4.08 $Y2=3.33
r135 56 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.59 $Y2=3.33
r136 56 59 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.08 $Y2=3.33
r137 54 73 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=2.64 $Y2=3.33
r138 53 54 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r139 51 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.625 $Y=3.33
+ $X2=2.79 $Y2=3.33
r140 51 53 155.599 $w=1.68e-07 $l=2.385e-06 $layer=LI1_cond $X=2.625 $Y=3.33
+ $X2=0.24 $Y2=3.33
r141 49 60 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.08 $Y2=3.33
r142 49 76 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r143 45 48 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=7.385 $Y=2.115
+ $X2=7.385 $Y2=2.815
r144 43 87 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=7.385 $Y=3.245
+ $X2=7.45 $Y2=3.33
r145 43 48 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.385 $Y=3.245
+ $X2=7.385 $Y2=2.815
r146 39 84 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.47 $Y=3.245
+ $X2=6.47 $Y2=3.33
r147 39 41 25.2897 $w=3.58e-07 $l=7.9e-07 $layer=LI1_cond $X=6.47 $Y=3.245
+ $X2=6.47 $Y2=2.455
r148 35 81 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.595 $Y=3.245
+ $X2=5.595 $Y2=3.33
r149 35 37 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=5.595 $Y=3.245
+ $X2=5.595 $Y2=2.805
r150 34 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.755 $Y=3.33
+ $X2=4.59 $Y2=3.33
r151 33 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.47 $Y=3.33
+ $X2=5.595 $Y2=3.33
r152 33 34 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=5.47 $Y=3.33
+ $X2=4.755 $Y2=3.33
r153 29 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.59 $Y=3.245
+ $X2=4.59 $Y2=3.33
r154 29 31 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.59 $Y=3.245
+ $X2=4.59 $Y2=2.78
r155 25 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=3.245
+ $X2=3.69 $Y2=3.33
r156 25 27 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.69 $Y=3.245
+ $X2=3.69 $Y2=2.78
r157 24 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.955 $Y=3.33
+ $X2=2.79 $Y2=3.33
r158 23 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.525 $Y=3.33
+ $X2=3.69 $Y2=3.33
r159 23 24 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.525 $Y=3.33
+ $X2=2.955 $Y2=3.33
r160 19 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.79 $Y=3.245
+ $X2=2.79 $Y2=3.33
r161 19 21 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.79 $Y=3.245
+ $X2=2.79 $Y2=2.78
r162 6 48 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.25
+ $Y=1.96 $X2=7.385 $Y2=2.815
r163 6 45 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=7.25
+ $Y=1.96 $X2=7.385 $Y2=2.115
r164 5 41 300 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=2 $X=6.32
+ $Y=1.96 $X2=6.47 $Y2=2.455
r165 4 37 600 $w=1.7e-07 $l=9.1e-07 $layer=licon1_PDIFF $count=1 $X=5.42 $Y=1.96
+ $X2=5.555 $Y2=2.805
r166 3 31 600 $w=1.7e-07 $l=1.00524e-06 $layer=licon1_PDIFF $count=1 $X=4.455
+ $Y=1.84 $X2=4.59 $Y2=2.78
r167 2 27 600 $w=1.7e-07 $l=1.00524e-06 $layer=licon1_PDIFF $count=1 $X=3.555
+ $Y=1.84 $X2=3.69 $Y2=2.78
r168 1 21 600 $w=1.7e-07 $l=1.00055e-06 $layer=licon1_PDIFF $count=1 $X=2.665
+ $Y=1.84 $X2=2.79 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_4%X 1 2 3 4 14 15 16 18 20 21 25 27 28 31 33
+ 35 36 38 41 44 48
c133 44 0 1.88456e-19 $X=2.755 $Y=0.555
r134 48 51 6.56993 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.24 $Y=0.925
+ $X2=0.24 $Y2=1.04
r135 41 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0.925
+ $X2=0.24 $Y2=0.925
r136 39 44 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=2.727 $Y=0.925
+ $X2=2.727 $Y2=0.555
r137 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0.925
+ $X2=2.64 $Y2=0.925
r138 36 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.385 $Y=0.925
+ $X2=0.24 $Y2=0.925
r139 35 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.495 $Y=0.925
+ $X2=2.64 $Y2=0.925
r140 35 36 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=2.495 $Y=0.925
+ $X2=0.385 $Y2=0.925
r141 34 39 1.64635 $w=3.83e-07 $l=5.5e-08 $layer=LI1_cond $X=2.727 $Y=0.98
+ $X2=2.727 $Y2=0.925
r142 29 31 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=3.62 $Y=0.98
+ $X2=3.62 $Y2=0.57
r143 28 34 8.24022 $w=1.7e-07 $l=2.31633e-07 $layer=LI1_cond $X=2.92 $Y=1.065
+ $X2=2.727 $Y2=0.98
r144 27 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.495 $Y=1.065
+ $X2=3.62 $Y2=0.98
r145 27 28 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=3.495 $Y=1.065
+ $X2=2.92 $Y2=1.065
r146 23 25 31.4303 $w=3.28e-07 $l=9e-07 $layer=LI1_cond $X=3.24 $Y=1.985
+ $X2=4.14 $Y2=1.985
r147 21 33 8.16218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=1.985
+ $X2=2.525 $Y2=1.985
r148 21 23 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=2.69 $Y=1.985
+ $X2=3.24 $Y2=1.985
r149 20 33 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=1.505 $Y=2.055
+ $X2=2.525 $Y2=2.055
r150 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.42 $Y=2.14
+ $X2=1.505 $Y2=2.055
r151 17 18 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.42 $Y=2.14
+ $X2=1.42 $Y2=2.36
r152 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.335 $Y=2.445
+ $X2=1.42 $Y2=2.36
r153 15 16 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=1.335 $Y=2.445
+ $X2=0.295 $Y2=2.445
r154 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.21 $Y=2.36
+ $X2=0.295 $Y2=2.445
r155 14 51 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=0.21 $Y=2.36
+ $X2=0.21 $Y2=1.04
r156 4 25 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.84 $X2=4.14 $Y2=1.985
r157 3 23 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.105
+ $Y=1.84 $X2=3.24 $Y2=1.985
r158 2 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.52
+ $Y=0.425 $X2=3.66 $Y2=0.57
r159 1 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.615
+ $Y=0.41 $X2=2.755 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_4%VGND 1 2 3 4 5 6 21 25 27 31 33 37 42 43 45
+ 48 49 50 51 53 62 72 73 76 79 82
c107 45 0 5.39098e-20 $X=5.01 $Y=1.02
r108 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r109 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r110 77 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r111 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r112 72 73 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r113 70 73 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=7.44 $Y2=0
r114 70 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r115 69 72 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=7.44
+ $Y2=0
r116 69 70 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r117 67 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.175 $Y=0 $X2=4.05
+ $Y2=0
r118 67 69 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.175 $Y=0
+ $X2=4.56 $Y2=0
r119 66 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r120 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r121 63 79 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=3.315 $Y=0
+ $X2=3.207 $Y2=0
r122 63 65 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.315 $Y=0 $X2=3.6
+ $Y2=0
r123 62 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.925 $Y=0 $X2=4.05
+ $Y2=0
r124 62 65 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.925 $Y=0 $X2=3.6
+ $Y2=0
r125 61 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r126 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r127 57 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r128 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r129 53 83 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=4.08 $Y2=0
r130 53 66 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r131 50 60 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.2
+ $Y2=0
r132 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.42
+ $Y2=0
r133 48 56 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.395 $Y=0
+ $X2=0.24 $Y2=0
r134 48 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.56
+ $Y2=0
r135 47 60 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=0.725 $Y=0 $X2=1.2
+ $Y2=0
r136 47 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=0 $X2=0.56
+ $Y2=0
r137 43 52 18.3822 $w=2.5e-07 $l=3.75e-07 $layer=LI1_cond $X=4.425 $Y=1.06
+ $X2=4.05 $Y2=1.06
r138 43 45 26.9672 $w=2.48e-07 $l=5.85e-07 $layer=LI1_cond $X=4.425 $Y=1.06
+ $X2=5.01 $Y2=1.06
r139 40 52 0.255588 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=4.05 $Y=0.935
+ $X2=4.05 $Y2=1.06
r140 40 42 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=4.05 $Y=0.935
+ $X2=4.05 $Y2=0.57
r141 39 82 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.05 $Y=0.085
+ $X2=4.05 $Y2=0
r142 39 42 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=4.05 $Y=0.085
+ $X2=4.05 $Y2=0.57
r143 35 79 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.207 $Y=0.085
+ $X2=3.207 $Y2=0
r144 35 37 27.873 $w=2.13e-07 $l=5.2e-07 $layer=LI1_cond $X=3.207 $Y=0.085
+ $X2=3.207 $Y2=0.605
r145 34 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.365 $Y=0 $X2=2.24
+ $Y2=0
r146 33 79 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=3.1 $Y=0 $X2=3.207
+ $Y2=0
r147 33 34 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=3.1 $Y=0 $X2=2.365
+ $Y2=0
r148 29 76 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=0.085
+ $X2=2.24 $Y2=0
r149 29 31 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=2.24 $Y=0.085
+ $X2=2.24 $Y2=0.795
r150 28 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.585 $Y=0 $X2=1.42
+ $Y2=0
r151 27 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=2.24
+ $Y2=0
r152 27 28 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.115 $Y=0
+ $X2=1.585 $Y2=0
r153 23 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.42 $Y=0.085
+ $X2=1.42 $Y2=0
r154 23 25 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.42 $Y=0.085
+ $X2=1.42 $Y2=0.535
r155 19 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.56 $Y=0.085
+ $X2=0.56 $Y2=0
r156 19 21 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.56 $Y=0.085
+ $X2=0.56 $Y2=0.555
r157 6 45 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=4.87
+ $Y=0.525 $X2=5.01 $Y2=1.02
r158 5 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.95
+ $Y=0.425 $X2=4.09 $Y2=0.57
r159 4 37 182 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_NDIFF $count=1 $X=3.045
+ $Y=0.41 $X2=3.205 $Y2=0.605
r160 3 31 182 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_NDIFF $count=1 $X=2.14
+ $Y=0.41 $X2=2.28 $Y2=0.795
r161 2 25 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.28
+ $Y=0.41 $X2=1.42 $Y2=0.535
r162 1 21 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.435
+ $Y=0.41 $X2=0.56 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_4%A_888_105# 1 2 12 14 15
r30 14 15 9.26861 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=6.94 $Y=0.705
+ $X2=6.775 $Y2=0.705
r31 12 15 132.439 $w=1.68e-07 $l=2.03e-06 $layer=LI1_cond $X=4.745 $Y=0.68
+ $X2=6.775 $Y2=0.68
r32 10 12 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.58 $Y=0.635
+ $X2=4.745 $Y2=0.635
r33 2 14 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.8
+ $Y=0.585 $X2=6.94 $Y2=0.73
r34 1 10 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=4.44
+ $Y=0.525 $X2=4.58 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_4%A_1081_39# 1 2 3 10 14 19 21
c30 14 0 8.35615e-20 $X=7.285 $Y=1.115
r31 19 23 3.47681 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=7.41 $Y=0.985
+ $X2=7.41 $Y2=1.115
r32 19 21 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=7.41 $Y=0.985
+ $X2=7.41 $Y2=0.73
r33 18 21 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=7.41 $Y=0.425
+ $X2=7.41 $Y2=0.73
r34 14 23 3.34309 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=7.285 $Y=1.115
+ $X2=7.41 $Y2=1.115
r35 14 16 37.0112 $w=2.58e-07 $l=8.35e-07 $layer=LI1_cond $X=7.285 $Y=1.115
+ $X2=6.45 $Y2=1.115
r36 10 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.285 $Y=0.34
+ $X2=7.41 $Y2=0.425
r37 10 12 114.497 $w=1.68e-07 $l=1.755e-06 $layer=LI1_cond $X=7.285 $Y=0.34
+ $X2=5.53 $Y2=0.34
r38 3 23 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=7.23
+ $Y=0.585 $X2=7.37 $Y2=1.08
r39 3 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.23
+ $Y=0.585 $X2=7.37 $Y2=0.73
r40 2 16 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=6.31
+ $Y=0.585 $X2=6.45 $Y2=1.075
r41 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=5.405
+ $Y=0.195 $X2=5.53 $Y2=0.34
.ends


* File: sky130_fd_sc_ms__dfxbp_2.pex.spice
* Created: Fri Aug 28 17:24:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DFXBP_2%CLK 3 7 8 11 12 13
c31 12 0 8.40497e-20 $X=0.42 $Y=1.385
r32 11 14 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.425 $Y=1.385
+ $X2=0.425 $Y2=1.55
r33 11 13 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.425 $Y=1.385
+ $X2=0.425 $Y2=1.22
r34 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.42
+ $Y=1.385 $X2=0.42 $Y2=1.385
r35 8 12 5.60648 $w=3.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.24 $Y=1.365
+ $X2=0.42 $Y2=1.365
r36 7 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=0.74
+ $X2=0.495 $Y2=1.22
r37 3 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.505 $Y=2.4
+ $X2=0.505 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_2%A_27_74# 1 2 9 11 13 14 16 18 21 25 27 28 30
+ 31 36 39 41 44 48 52 53 54 55 57 59 60 63 64 65 67 69 70 73 74 75 77 80 83 85
+ 94 95 99 107 112 114
c266 107 0 1.39464e-19 $X=1.14 $Y=1.385
c267 85 0 4.88492e-20 $X=0.97 $Y=1.385
c268 80 0 6.69395e-20 $X=6.075 $Y=0.365
c269 59 0 1.39925e-19 $X=0.84 $Y=1.72
c270 54 0 7.68583e-20 $X=0.755 $Y=1.805
c271 39 0 2.47898e-20 $X=3.12 $Y=1.165
c272 31 0 2.58209e-19 $X=6.09 $Y=1.245
c273 21 0 1.22749e-19 $X=3.435 $Y=2.435
c274 11 0 1.50442e-19 $X=1.14 $Y=1.22
r275 100 117 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.68 $Y=1.335
+ $X2=5.68 $Y2=1.5
r276 100 114 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.68 $Y=1.335
+ $X2=5.68 $Y2=1.245
r277 99 100 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.68
+ $Y=1.335 $X2=5.68 $Y2=1.335
r278 96 99 6.1738 $w=2.78e-07 $l=1.5e-07 $layer=LI1_cond $X=5.53 $Y=1.31
+ $X2=5.68 $Y2=1.31
r279 90 112 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=3.39 $Y=1.9
+ $X2=3.435 $Y2=1.9
r280 90 109 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=3.39 $Y=1.9
+ $X2=3.12 $Y2=1.9
r281 89 90 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.39
+ $Y=1.9 $X2=3.39 $Y2=1.9
r282 86 107 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=0.97 $Y=1.385
+ $X2=1.14 $Y2=1.385
r283 86 104 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.97 $Y=1.385
+ $X2=0.955 $Y2=1.385
r284 85 87 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=0.927 $Y=1.385
+ $X2=0.927 $Y2=1.55
r285 85 86 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=1.385 $X2=0.97 $Y2=1.385
r286 80 81 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.075
+ $Y=0.365 $X2=6.075 $Y2=0.365
r287 78 95 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=5.615 $Y=0.392
+ $X2=5.53 $Y2=0.392
r288 78 80 19.2772 $w=2.73e-07 $l=4.6e-07 $layer=LI1_cond $X=5.615 $Y=0.392
+ $X2=6.075 $Y2=0.392
r289 77 96 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.53 $Y=1.17
+ $X2=5.53 $Y2=1.31
r290 76 95 3.11956 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=5.53 $Y=0.53
+ $X2=5.53 $Y2=0.392
r291 76 77 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.53 $Y=0.53
+ $X2=5.53 $Y2=1.17
r292 74 95 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=5.445 $Y=0.392
+ $X2=5.53 $Y2=0.392
r293 74 75 26.4014 $w=2.73e-07 $l=6.3e-07 $layer=LI1_cond $X=5.445 $Y=0.392
+ $X2=4.815 $Y2=0.392
r294 72 75 7.32204 $w=2.75e-07 $l=1.75425e-07 $layer=LI1_cond $X=4.73 $Y=0.53
+ $X2=4.815 $Y2=0.392
r295 72 73 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.73 $Y=0.53
+ $X2=4.73 $Y2=0.78
r296 71 94 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=0.865
+ $X2=3.555 $Y2=0.865
r297 70 73 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.645 $Y=0.865
+ $X2=4.73 $Y2=0.78
r298 70 71 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=4.645 $Y=0.865
+ $X2=3.64 $Y2=0.865
r299 69 89 6.03661 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=1.907
+ $X2=3.39 $Y2=1.907
r300 68 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.555 $Y=0.95
+ $X2=3.555 $Y2=0.865
r301 68 69 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=3.555 $Y=0.95
+ $X2=3.555 $Y2=1.75
r302 67 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.555 $Y=0.78
+ $X2=3.555 $Y2=0.865
r303 66 67 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.555 $Y=0.425
+ $X2=3.555 $Y2=0.78
r304 64 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.47 $Y=0.34
+ $X2=3.555 $Y2=0.425
r305 64 65 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.47 $Y=0.34
+ $X2=2.53 $Y2=0.34
r306 62 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.445 $Y=0.425
+ $X2=2.53 $Y2=0.34
r307 62 63 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.445 $Y=0.425
+ $X2=2.445 $Y2=0.73
r308 61 83 7.25401 $w=2.25e-07 $l=1.98605e-07 $layer=LI1_cond $X=1.1 $Y=0.815
+ $X2=0.927 $Y2=0.87
r309 60 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.36 $Y=0.815
+ $X2=2.445 $Y2=0.73
r310 60 61 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=2.36 $Y=0.815
+ $X2=1.1 $Y2=0.815
r311 59 87 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.84 $Y=1.72
+ $X2=0.84 $Y2=1.55
r312 57 85 0.233829 $w=3.43e-07 $l=7e-09 $layer=LI1_cond $X=0.927 $Y=1.378
+ $X2=0.927 $Y2=1.385
r313 56 83 0.140858 $w=3.45e-07 $l=1.4e-07 $layer=LI1_cond $X=0.927 $Y=1.01
+ $X2=0.927 $Y2=0.87
r314 56 57 12.2927 $w=3.43e-07 $l=3.68e-07 $layer=LI1_cond $X=0.927 $Y=1.01
+ $X2=0.927 $Y2=1.378
r315 54 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.755 $Y=1.805
+ $X2=0.84 $Y2=1.72
r316 54 55 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.755 $Y=1.805
+ $X2=0.445 $Y2=1.805
r317 52 83 7.25401 $w=2.25e-07 $l=1.72e-07 $layer=LI1_cond $X=0.755 $Y=0.87
+ $X2=0.927 $Y2=0.87
r318 52 53 12.7592 $w=2.78e-07 $l=3.1e-07 $layer=LI1_cond $X=0.755 $Y=0.87
+ $X2=0.445 $Y2=0.87
r319 48 50 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r320 46 55 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.89
+ $X2=0.445 $Y2=1.805
r321 46 48 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.28 $Y=1.89
+ $X2=0.28 $Y2=1.985
r322 42 53 6.87623 $w=2.8e-07 $l=2.24332e-07 $layer=LI1_cond $X=0.28 $Y=0.73
+ $X2=0.445 $Y2=0.87
r323 42 44 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=0.28 $Y=0.73
+ $X2=0.28 $Y2=0.515
r324 41 81 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.09 $Y=0.365
+ $X2=6.075 $Y2=0.365
r325 37 39 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=3 $Y=1.165 $X2=3.12
+ $Y2=1.165
r326 34 36 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.165 $Y=1.17
+ $X2=6.165 $Y2=0.85
r327 33 41 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=6.165 $Y=0.53
+ $X2=6.09 $Y2=0.365
r328 33 36 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.165 $Y=0.53
+ $X2=6.165 $Y2=0.85
r329 32 114 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.845 $Y=1.245
+ $X2=5.68 $Y2=1.245
r330 31 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.09 $Y=1.245
+ $X2=6.165 $Y2=1.17
r331 31 32 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=6.09 $Y=1.245
+ $X2=5.845 $Y2=1.245
r332 30 117 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.59 $Y=1.69
+ $X2=5.59 $Y2=1.5
r333 27 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.515 $Y=1.765
+ $X2=5.59 $Y2=1.69
r334 27 28 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=5.515 $Y=1.765
+ $X2=5.015 $Y2=1.765
r335 23 28 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.925 $Y=1.84
+ $X2=5.015 $Y2=1.765
r336 23 25 272.097 $w=1.8e-07 $l=7e-07 $layer=POLY_cond $X=4.925 $Y=1.84
+ $X2=4.925 $Y2=2.54
r337 19 112 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.435 $Y=2.065
+ $X2=3.435 $Y2=1.9
r338 19 21 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=3.435 $Y=2.065
+ $X2=3.435 $Y2=2.435
r339 18 109 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.12 $Y=1.735
+ $X2=3.12 $Y2=1.9
r340 17 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.12 $Y=1.24
+ $X2=3.12 $Y2=1.165
r341 17 18 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.12 $Y=1.24
+ $X2=3.12 $Y2=1.735
r342 14 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3 $Y=1.09 $X2=3
+ $Y2=1.165
r343 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3 $Y=1.09 $X2=3
+ $Y2=0.805
r344 11 107 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.22
+ $X2=1.14 $Y2=1.385
r345 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.14 $Y=1.22
+ $X2=1.14 $Y2=0.74
r346 7 104 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.55
+ $X2=0.955 $Y2=1.385
r347 7 9 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.955 $Y=1.55
+ $X2=0.955 $Y2=2.4
r348 2 50 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r349 2 48 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r350 1 44 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_2%D 3 5 7 11 13 15 16 22 25 34
c55 34 0 6.95252e-20 $X=2.16 $Y=1.665
c56 25 0 3.91626e-20 $X=2.21 $Y=1.29
c57 15 0 4.82751e-20 $X=2.16 $Y=1.295
r58 28 34 2.36399 $w=3.88e-07 $l=8e-08 $layer=LI1_cond $X=2.18 $Y=1.585 $X2=2.18
+ $Y2=1.665
r59 16 36 7.07103 $w=3.88e-07 $l=1.13e-07 $layer=LI1_cond $X=2.18 $Y=1.667
+ $X2=2.18 $Y2=1.78
r60 16 34 0.0590996 $w=3.88e-07 $l=2e-09 $layer=LI1_cond $X=2.18 $Y=1.667
+ $X2=2.18 $Y2=1.665
r61 16 28 0.0886495 $w=3.88e-07 $l=3e-09 $layer=LI1_cond $X=2.18 $Y=1.582
+ $X2=2.18 $Y2=1.585
r62 15 16 8.62855 $w=3.88e-07 $l=2.92e-07 $layer=LI1_cond $X=2.18 $Y=1.29
+ $X2=2.18 $Y2=1.582
r63 15 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.21
+ $Y=1.29 $X2=2.21 $Y2=1.29
r64 13 36 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.07 $Y=2.025
+ $X2=2.07 $Y2=1.78
r65 12 22 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=1.99 $Y=2.19
+ $X2=2.18 $Y2=2.19
r66 11 13 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.99 $Y=2.19
+ $X2=1.99 $Y2=2.025
r67 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.99
+ $Y=2.19 $X2=1.99 $Y2=2.19
r68 5 25 69.6867 $w=2.49e-07 $l=4.34741e-07 $layer=POLY_cond $X=2.57 $Y=1.125
+ $X2=2.21 $Y2=1.29
r69 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.57 $Y=1.125 $X2=2.57
+ $Y2=0.805
r70 1 22 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.18 $Y=2.355
+ $X2=2.18 $Y2=2.19
r71 1 3 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=2.18 $Y=2.355 $X2=2.18
+ $Y2=2.725
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_2%A_209_368# 1 2 9 10 11 15 19 23 27 30 33 35
+ 38 39 43 44 49 52 56 57 60 64
c184 52 0 2.65632e-19 $X=1.65 $Y=1.65
c185 43 0 1.39777e-19 $X=6.04 $Y=2.07
r186 60 61 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.12 $Y=2.71
+ $X2=5.12 $Y2=2.88
r187 57 67 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.14 $Y=1.285
+ $X2=5.015 $Y2=1.285
r188 56 59 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=5.13 $Y=1.285
+ $X2=5.13 $Y2=1.45
r189 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.14
+ $Y=1.285 $X2=5.14 $Y2=1.285
r190 52 65 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.65 $Y=1.65 $X2=1.65
+ $Y2=1.74
r191 52 64 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.65 $Y=1.65
+ $X2=1.65 $Y2=1.485
r192 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.65 $X2=1.65 $Y2=1.65
r193 49 51 7.9006 $w=3.32e-07 $l=2.15e-07 $layer=LI1_cond $X=1.435 $Y=1.736
+ $X2=1.65 $Y2=1.736
r194 44 73 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.04 $Y=2.07
+ $X2=6.04 $Y2=2.235
r195 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.04
+ $Y=2.07 $X2=6.04 $Y2=2.07
r196 41 43 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=6.04 $Y=2.795
+ $X2=6.04 $Y2=2.07
r197 40 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.205 $Y=2.88
+ $X2=5.12 $Y2=2.88
r198 39 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.875 $Y=2.88
+ $X2=6.04 $Y2=2.795
r199 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.875 $Y=2.88
+ $X2=5.205 $Y2=2.88
r200 38 60 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.12 $Y=2.625
+ $X2=5.12 $Y2=2.71
r201 38 59 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=5.12 $Y=2.625
+ $X2=5.12 $Y2=1.45
r202 36 54 4.73278 $w=1.7e-07 $l=2.14114e-07 $layer=LI1_cond $X=1.44 $Y=2.71
+ $X2=1.267 $Y2=2.802
r203 35 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.035 $Y=2.71
+ $X2=5.12 $Y2=2.71
r204 35 36 234.54 $w=1.68e-07 $l=3.595e-06 $layer=LI1_cond $X=5.035 $Y=2.71
+ $X2=1.44 $Y2=2.71
r205 31 49 0.753319 $w=3.3e-07 $l=2.51e-07 $layer=LI1_cond $X=1.435 $Y=1.485
+ $X2=1.435 $Y2=1.736
r206 31 33 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.435 $Y=1.485
+ $X2=1.435 $Y2=1.155
r207 30 54 3.16114 $w=3.45e-07 $l=1.77e-07 $layer=LI1_cond $X=1.267 $Y=2.625
+ $X2=1.267 $Y2=2.802
r208 29 49 6.17349 $w=3.32e-07 $l=3.24298e-07 $layer=LI1_cond $X=1.267 $Y=1.987
+ $X2=1.435 $Y2=1.736
r209 29 47 3.19699 $w=3.32e-07 $l=8.79943e-08 $layer=LI1_cond $X=1.267 $Y=1.987
+ $X2=1.18 $Y2=1.985
r210 29 30 21.3118 $w=3.43e-07 $l=6.38e-07 $layer=LI1_cond $X=1.267 $Y=1.987
+ $X2=1.267 $Y2=2.625
r211 27 73 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=5.965 $Y=2.605
+ $X2=5.965 $Y2=2.235
r212 21 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.015 $Y=1.12
+ $X2=5.015 $Y2=1.285
r213 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.015 $Y=1.12
+ $X2=5.015 $Y2=0.655
r214 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.51 $Y=0.255
+ $X2=3.51 $Y2=0.72
r215 13 15 241 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=2.715 $Y=1.815
+ $X2=2.715 $Y2=2.435
r216 12 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.74
+ $X2=1.65 $Y2=1.74
r217 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.625 $Y=1.74
+ $X2=2.715 $Y2=1.815
r218 11 12 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.625 $Y=1.74
+ $X2=1.815 $Y2=1.74
r219 9 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.435 $Y=0.18
+ $X2=3.51 $Y2=0.255
r220 9 10 835.809 $w=1.5e-07 $l=1.63e-06 $layer=POLY_cond $X=3.435 $Y=0.18
+ $X2=1.805 $Y2=0.18
r221 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.73 $Y=0.255
+ $X2=1.805 $Y2=0.18
r222 7 64 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=1.73 $Y=0.255
+ $X2=1.73 $Y2=1.485
r223 2 54 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.815
r224 2 47 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=1.985
r225 1 33 182 $w=1.7e-07 $l=8.88214e-07 $layer=licon1_NDIFF $count=1 $X=1.215
+ $Y=0.37 $X2=1.435 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_2%A_753_284# 1 2 7 9 13 15 20 21
c55 13 0 3.89984e-20 $X=3.9 $Y=0.72
r56 21 23 1.25721 $w=2.73e-07 $l=3e-08 $layer=LI1_cond $X=4.73 $Y=2.317 $X2=4.7
+ $Y2=2.317
r57 20 28 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.73 $Y=1.45
+ $X2=4.73 $Y2=1.285
r58 20 21 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.73 $Y=1.45
+ $X2=4.73 $Y2=2.18
r59 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.975
+ $Y=1.255 $X2=3.975 $Y2=1.255
r60 15 28 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.645 $Y=1.285
+ $X2=4.73 $Y2=1.285
r61 15 17 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=4.645 $Y=1.285
+ $X2=3.975 $Y2=1.285
r62 11 18 38.532 $w=3.09e-07 $l=1.89222e-07 $layer=POLY_cond $X=3.9 $Y=1.09
+ $X2=3.952 $Y2=1.255
r63 11 13 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.9 $Y=1.09 $X2=3.9
+ $Y2=0.72
r64 7 18 48.107 $w=3.09e-07 $l=2.996e-07 $layer=POLY_cond $X=3.855 $Y=1.51
+ $X2=3.952 $Y2=1.255
r65 7 9 359.556 $w=1.8e-07 $l=9.25e-07 $layer=POLY_cond $X=3.855 $Y=1.51
+ $X2=3.855 $Y2=2.435
r66 2 23 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=4.565
+ $Y=2.12 $X2=4.7 $Y2=2.275
r67 1 28 182 $w=1.7e-07 $l=1.00902e-06 $layer=licon1_NDIFF $count=1 $X=4.5
+ $Y=0.38 $X2=4.72 $Y2=1.285
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_2%A_561_445# 1 2 9 13 16 17 19 21 22 26 32 33
c79 19 0 1.01646e-19 $X=3.215 $Y=0.815
r80 33 38 40.172 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=4.36 $Y=1.795
+ $X2=4.36 $Y2=1.96
r81 33 37 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=4.36 $Y=1.795
+ $X2=4.36 $Y2=1.63
r82 32 35 8.46025 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=4.315 $Y=1.795
+ $X2=4.315 $Y2=1.96
r83 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.32
+ $Y=1.795 $X2=4.32 $Y2=1.795
r84 26 35 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.24 $Y=2.285
+ $X2=4.24 $Y2=1.96
r85 22 24 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=3.055 $Y=2.37
+ $X2=3.085 $Y2=2.37
r86 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.155 $Y=2.37
+ $X2=4.24 $Y2=2.285
r87 21 24 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=4.155 $Y=2.37
+ $X2=3.085 $Y2=2.37
r88 17 27 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.175 $Y=1.495
+ $X2=2.97 $Y2=1.495
r89 17 19 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=3.175 $Y=1.41
+ $X2=3.175 $Y2=0.815
r90 16 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.97 $Y=2.285
+ $X2=3.055 $Y2=2.37
r91 15 27 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=1.58
+ $X2=2.97 $Y2=1.495
r92 15 16 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.97 $Y=1.58
+ $X2=2.97 $Y2=2.285
r93 13 38 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=4.475 $Y=2.54
+ $X2=4.475 $Y2=1.96
r94 9 37 499.947 $w=1.5e-07 $l=9.75e-07 $layer=POLY_cond $X=4.425 $Y=0.655
+ $X2=4.425 $Y2=1.63
r95 2 24 600 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_PDIFF $count=1 $X=2.805
+ $Y=2.225 $X2=3.085 $Y2=2.37
r96 1 19 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=3.075
+ $Y=0.595 $X2=3.215 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_2%A_1290_102# 1 2 7 9 12 14 18 22 24 28 32 36
+ 40 43 44 45 47 48 49 50 53 59 61 64 65 69 73 76 77
c158 7 0 6.69395e-20 $X=6.525 $Y=1.17
r159 75 76 5.26419 $w=2.78e-07 $l=8.5e-08 $layer=LI1_cond $X=7.84 $Y=2.27
+ $X2=7.925 $Y2=2.27
r160 73 75 21.1967 $w=2.78e-07 $l=5.15e-07 $layer=LI1_cond $X=7.325 $Y=2.27
+ $X2=7.84 $Y2=2.27
r161 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.85
+ $Y=1.485 $X2=8.85 $Y2=1.485
r162 67 69 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=8.85 $Y=2.24
+ $X2=8.85 $Y2=1.485
r163 65 67 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.685 $Y=2.325
+ $X2=8.85 $Y2=2.24
r164 65 76 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=8.685 $Y=2.325
+ $X2=7.925 $Y2=2.325
r165 64 75 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=7.84 $Y=2.13
+ $X2=7.84 $Y2=2.27
r166 63 64 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=7.84 $Y=1.5
+ $X2=7.84 $Y2=2.13
r167 62 77 5.16603 $w=2.5e-07 $l=1.60078e-07 $layer=LI1_cond $X=7.465 $Y=1.415
+ $X2=7.34 $Y2=1.335
r168 61 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.755 $Y=1.415
+ $X2=7.84 $Y2=1.5
r169 61 62 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=7.755 $Y=1.415
+ $X2=7.465 $Y2=1.415
r170 57 77 1.34256 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=7.34 $Y=1.17
+ $X2=7.34 $Y2=1.335
r171 57 59 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=7.34 $Y=1.17
+ $X2=7.34 $Y2=0.535
r172 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.88
+ $Y=1.335 $X2=6.88 $Y2=1.335
r173 50 77 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=7.215 $Y=1.335
+ $X2=7.34 $Y2=1.335
r174 50 52 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.215 $Y=1.335
+ $X2=6.88 $Y2=1.335
r175 48 70 105.791 $w=3.3e-07 $l=6.05e-07 $layer=POLY_cond $X=9.455 $Y=1.485
+ $X2=8.85 $Y2=1.485
r176 48 49 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.455 $Y=1.485
+ $X2=9.545 $Y2=1.485
r177 46 70 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=8.625 $Y=1.485
+ $X2=8.85 $Y2=1.485
r178 46 47 7.86782 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=8.625 $Y=1.485
+ $X2=8.525 $Y2=1.485
r179 42 53 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=6.6 $Y=1.335
+ $X2=6.88 $Y2=1.335
r180 42 43 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.6 $Y=1.335
+ $X2=6.525 $Y2=1.335
r181 38 49 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=9.56 $Y=1.32
+ $X2=9.545 $Y2=1.485
r182 38 40 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=9.56 $Y=1.32
+ $X2=9.56 $Y2=0.835
r183 34 49 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=9.545 $Y=1.65
+ $X2=9.545 $Y2=1.485
r184 34 36 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=9.545 $Y=1.65
+ $X2=9.545 $Y2=2.34
r185 30 47 16.8416 $w=1.8e-07 $l=1.69926e-07 $layer=POLY_cond $X=8.535 $Y=1.65
+ $X2=8.525 $Y2=1.485
r186 30 32 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=8.535 $Y=1.65
+ $X2=8.535 $Y2=2.4
r187 26 47 16.8416 $w=1.5e-07 $l=1.77059e-07 $layer=POLY_cond $X=8.5 $Y=1.32
+ $X2=8.525 $Y2=1.485
r188 26 28 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.5 $Y=1.32 $X2=8.5
+ $Y2=0.76
r189 25 45 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.175 $Y=1.395
+ $X2=8.085 $Y2=1.395
r190 24 47 7.86782 $w=1.5e-07 $l=1.3784e-07 $layer=POLY_cond $X=8.425 $Y=1.395
+ $X2=8.525 $Y2=1.485
r191 24 25 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.425 $Y=1.395
+ $X2=8.175 $Y2=1.395
r192 20 45 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=8.085 $Y=1.47
+ $X2=8.085 $Y2=1.395
r193 20 22 361.5 $w=1.8e-07 $l=9.3e-07 $layer=POLY_cond $X=8.085 $Y=1.47
+ $X2=8.085 $Y2=2.4
r194 16 45 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=8.07 $Y=1.32
+ $X2=8.085 $Y2=1.395
r195 16 18 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.07 $Y=1.32
+ $X2=8.07 $Y2=0.76
r196 12 44 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.54 $Y=1.83 $X2=6.54
+ $Y2=1.74
r197 12 14 301.25 $w=1.8e-07 $l=7.75e-07 $layer=POLY_cond $X=6.54 $Y=1.83
+ $X2=6.54 $Y2=2.605
r198 10 43 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.525 $Y=1.5
+ $X2=6.525 $Y2=1.335
r199 10 44 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=6.525 $Y=1.5
+ $X2=6.525 $Y2=1.74
r200 7 43 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.525 $Y=1.17
+ $X2=6.525 $Y2=1.335
r201 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.525 $Y=1.17
+ $X2=6.525 $Y2=0.85
r202 2 73 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=7.19
+ $Y=2.12 $X2=7.325 $Y2=2.295
r203 1 59 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=7.235
+ $Y=0.39 $X2=7.38 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_2%A_1003_424# 1 2 9 13 17 21 23 24 26 31 37 39
+ 40 41 44
c107 37 0 1.18432e-19 $X=6.1 $Y=0.825
r108 44 45 8.24715 $w=2.63e-07 $l=4.5e-08 $layer=POLY_cond $X=7.55 $Y=1.795
+ $X2=7.595 $Y2=1.795
r109 40 41 8.71257 $w=2.88e-07 $l=1.7e-07 $layer=LI1_cond $X=6.375 $Y=1.79
+ $X2=6.545 $Y2=1.79
r110 35 37 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=5.95 $Y=0.825
+ $X2=6.1 $Y2=0.825
r111 32 44 23.8251 $w=2.63e-07 $l=1.3e-07 $layer=POLY_cond $X=7.42 $Y=1.795
+ $X2=7.55 $Y2=1.795
r112 31 41 34.772 $w=2.88e-07 $l=8.75e-07 $layer=LI1_cond $X=7.42 $Y=1.815
+ $X2=6.545 $Y2=1.815
r113 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.42
+ $Y=1.795 $X2=7.42 $Y2=1.795
r114 28 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.185 $Y=1.705
+ $X2=6.1 $Y2=1.705
r115 28 40 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=6.185 $Y=1.705
+ $X2=6.375 $Y2=1.705
r116 26 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.1 $Y=1.62 $X2=6.1
+ $Y2=1.705
r117 25 37 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.1 $Y=0.95 $X2=6.1
+ $Y2=0.825
r118 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.1 $Y=0.95 $X2=6.1
+ $Y2=1.62
r119 23 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.015 $Y=1.705
+ $X2=6.1 $Y2=1.705
r120 23 24 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.015 $Y=1.705
+ $X2=5.705 $Y2=1.705
r121 19 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.54 $Y=1.79
+ $X2=5.705 $Y2=1.705
r122 19 21 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=5.54 $Y=1.79
+ $X2=5.54 $Y2=2.54
r123 15 45 15.8942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.595 $Y=1.63
+ $X2=7.595 $Y2=1.795
r124 15 17 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=7.595 $Y=1.63
+ $X2=7.595 $Y2=0.76
r125 11 44 11.6845 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.55 $Y=1.96
+ $X2=7.55 $Y2=1.795
r126 11 13 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=7.55 $Y=1.96
+ $X2=7.55 $Y2=2.54
r127 7 32 58.6464 $w=2.63e-07 $l=3.93954e-07 $layer=POLY_cond $X=7.1 $Y=1.96
+ $X2=7.42 $Y2=1.795
r128 7 9 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=7.1 $Y=1.96 $X2=7.1
+ $Y2=2.54
r129 2 21 600 $w=1.7e-07 $l=7.04361e-07 $layer=licon1_PDIFF $count=1 $X=5.015
+ $Y=2.12 $X2=5.54 $Y2=2.54
r130 1 35 182 $w=1.7e-07 $l=1.04302e-06 $layer=licon1_NDIFF $count=1 $X=5.09
+ $Y=0.38 $X2=5.95 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_2%A_1835_368# 1 2 9 13 17 21 25 29 35 38 44
c70 29 0 8.25183e-20 $X=9.32 $Y=1.985
r71 43 44 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=10.53 $Y=1.465
+ $X2=10.545 $Y2=1.465
r72 42 43 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=10.115 $Y=1.465
+ $X2=10.53 $Y2=1.465
r73 41 42 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=10.08 $Y=1.465
+ $X2=10.115 $Y2=1.465
r74 36 41 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=10.01 $Y=1.465
+ $X2=10.08 $Y2=1.465
r75 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.01
+ $Y=1.465 $X2=10.01 $Y2=1.465
r76 33 38 0.533013 $w=3.3e-07 $l=1.38e-07 $layer=LI1_cond $X=9.51 $Y=1.465
+ $X2=9.372 $Y2=1.465
r77 33 35 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=9.51 $Y=1.465
+ $X2=10.01 $Y2=1.465
r78 29 31 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=9.36 $Y=1.985
+ $X2=9.36 $Y2=2.695
r79 27 38 6.22203 $w=2.62e-07 $l=1.70895e-07 $layer=LI1_cond $X=9.36 $Y=1.63
+ $X2=9.372 $Y2=1.465
r80 27 29 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=9.36 $Y=1.63
+ $X2=9.36 $Y2=1.985
r81 23 38 6.22203 $w=2.62e-07 $l=1.65e-07 $layer=LI1_cond $X=9.372 $Y=1.3
+ $X2=9.372 $Y2=1.465
r82 23 25 19.4868 $w=2.73e-07 $l=4.65e-07 $layer=LI1_cond $X=9.372 $Y=1.3
+ $X2=9.372 $Y2=0.835
r83 19 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.545 $Y=1.3
+ $X2=10.545 $Y2=1.465
r84 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=10.545 $Y=1.3
+ $X2=10.545 $Y2=0.74
r85 15 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.53 $Y=1.63
+ $X2=10.53 $Y2=1.465
r86 15 17 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=10.53 $Y=1.63
+ $X2=10.53 $Y2=2.4
r87 11 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.115 $Y=1.3
+ $X2=10.115 $Y2=1.465
r88 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=10.115 $Y=1.3
+ $X2=10.115 $Y2=0.74
r89 7 41 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.08 $Y=1.63
+ $X2=10.08 $Y2=1.465
r90 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=10.08 $Y=1.63
+ $X2=10.08 $Y2=2.4
r91 2 31 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=9.175
+ $Y=1.84 $X2=9.32 $Y2=2.695
r92 2 29 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=9.175
+ $Y=1.84 $X2=9.32 $Y2=1.985
r93 1 25 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=9.2
+ $Y=0.56 $X2=9.345 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_2%VPWR 1 2 3 4 5 6 7 8 29 33 37 41 45 49 51 56
+ 57 59 60 61 68 80 88 92 98 103 106 108 115 118 122
c118 29 0 1.39464e-19 $X=0.73 $Y=2.225
r119 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r120 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r121 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r122 111 112 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r123 108 111 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=4.165 $Y=3.05
+ $X2=4.165 $Y2=3.33
r124 105 106 10.9518 $w=4.48e-07 $l=2.3e-07 $layer=LI1_cond $X=1.805 $Y=3.19
+ $X2=2.035 $Y2=3.19
r125 101 105 3.32244 $w=4.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.68 $Y=3.19
+ $X2=1.805 $Y2=3.19
r126 101 103 7.62935 $w=4.48e-07 $l=1.05e-07 $layer=LI1_cond $X=1.68 $Y=3.19
+ $X2=1.575 $Y2=3.19
r127 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r128 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r129 96 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r130 96 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r131 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r132 93 118 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.94 $Y=3.33
+ $X2=9.815 $Y2=3.33
r133 93 95 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.94 $Y=3.33
+ $X2=10.32 $Y2=3.33
r134 92 121 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=10.675 $Y=3.33
+ $X2=10.857 $Y2=3.33
r135 92 95 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=10.675 $Y=3.33
+ $X2=10.32 $Y2=3.33
r136 91 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r137 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r138 88 118 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.69 $Y=3.33
+ $X2=9.815 $Y2=3.33
r139 88 90 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.69 $Y=3.33
+ $X2=9.36 $Y2=3.33
r140 87 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r141 87 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r142 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r143 84 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=7.86 $Y2=3.33
r144 84 86 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=8.4 $Y2=3.33
r145 83 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r146 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r147 80 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.695 $Y=3.33
+ $X2=7.86 $Y2=3.33
r148 80 82 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.695 $Y=3.33
+ $X2=7.44 $Y2=3.33
r149 79 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r150 78 79 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r151 76 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r152 75 78 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r153 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r154 73 111 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=3.33
+ $X2=4.165 $Y2=3.33
r155 73 75 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.33 $Y=3.33
+ $X2=4.56 $Y2=3.33
r156 72 112 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r157 72 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r158 71 106 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=2.035 $Y2=3.33
r159 71 72 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r160 68 111 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4 $Y=3.33
+ $X2=4.165 $Y2=3.33
r161 68 71 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4 $Y=3.33 $X2=2.16
+ $Y2=3.33
r162 67 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r163 67 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r164 66 103 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=1.575 $Y2=3.33
r165 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r166 64 98 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.77 $Y2=3.33
r167 64 66 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r168 61 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r169 61 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r170 59 86 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=8.595 $Y=3.33
+ $X2=8.4 $Y2=3.33
r171 59 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.595 $Y=3.33
+ $X2=8.76 $Y2=3.33
r172 58 90 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=8.925 $Y=3.33
+ $X2=9.36 $Y2=3.33
r173 58 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.925 $Y=3.33
+ $X2=8.76 $Y2=3.33
r174 56 78 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=6.6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r175 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.6 $Y=3.33
+ $X2=6.765 $Y2=3.33
r176 55 82 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.93 $Y=3.33
+ $X2=7.44 $Y2=3.33
r177 55 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.93 $Y=3.33
+ $X2=6.765 $Y2=3.33
r178 51 54 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=10.8 $Y=1.985
+ $X2=10.8 $Y2=2.815
r179 49 121 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.8 $Y=3.245
+ $X2=10.857 $Y2=3.33
r180 49 54 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.8 $Y=3.245
+ $X2=10.8 $Y2=2.815
r181 45 48 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=9.815 $Y=1.985
+ $X2=9.815 $Y2=2.815
r182 43 118 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.815 $Y=3.245
+ $X2=9.815 $Y2=3.33
r183 43 48 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.815 $Y=3.245
+ $X2=9.815 $Y2=2.815
r184 39 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.76 $Y=3.245
+ $X2=8.76 $Y2=3.33
r185 39 41 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=8.76 $Y=3.245
+ $X2=8.76 $Y2=2.78
r186 35 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.86 $Y=3.245
+ $X2=7.86 $Y2=3.33
r187 35 37 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=7.86 $Y=3.245
+ $X2=7.86 $Y2=2.78
r188 31 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.765 $Y=3.245
+ $X2=6.765 $Y2=3.33
r189 31 33 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=6.765 $Y=3.245
+ $X2=6.765 $Y2=2.605
r190 27 98 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=3.245
+ $X2=0.77 $Y2=3.33
r191 27 29 47.0197 $w=2.48e-07 $l=1.02e-06 $layer=LI1_cond $X=0.77 $Y=3.245
+ $X2=0.77 $Y2=2.225
r192 8 54 400 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=1 $X=10.62
+ $Y=1.84 $X2=10.76 $Y2=2.815
r193 8 51 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.62
+ $Y=1.84 $X2=10.76 $Y2=1.985
r194 7 48 600 $w=1.7e-07 $l=1.07941e-06 $layer=licon1_PDIFF $count=1 $X=9.635
+ $Y=1.84 $X2=9.855 $Y2=2.815
r195 7 45 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=9.635
+ $Y=1.84 $X2=9.855 $Y2=1.985
r196 6 41 600 $w=1.7e-07 $l=1.00524e-06 $layer=licon1_PDIFF $count=1 $X=8.625
+ $Y=1.84 $X2=8.76 $Y2=2.78
r197 5 37 600 $w=1.7e-07 $l=7.62102e-07 $layer=licon1_PDIFF $count=1 $X=7.64
+ $Y=2.12 $X2=7.86 $Y2=2.78
r198 4 33 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=6.63
+ $Y=2.395 $X2=6.765 $Y2=2.605
r199 3 108 600 $w=1.7e-07 $l=9.28507e-07 $layer=licon1_PDIFF $count=1 $X=3.945
+ $Y=2.225 $X2=4.165 $Y2=3.05
r200 2 105 600 $w=1.7e-07 $l=6.31328e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=2.515 $X2=1.805 $Y2=3.05
r201 1 29 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_2%A_454_503# 1 2 8 11 16 20
c35 16 0 1.22749e-19 $X=2.63 $Y=2.33
r36 18 20 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.63 $Y=1.155
+ $X2=2.785 $Y2=1.155
r37 14 16 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=2.49 $Y=2.33
+ $X2=2.63 $Y2=2.33
r38 9 20 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.785 $Y=1.07
+ $X2=2.785 $Y2=1.155
r39 9 11 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.785 $Y=1.07
+ $X2=2.785 $Y2=0.815
r40 8 16 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.63 $Y=2.205
+ $X2=2.63 $Y2=2.33
r41 7 18 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=1.24 $X2=2.63
+ $Y2=1.155
r42 7 8 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=2.63 $Y=1.24 $X2=2.63
+ $Y2=2.205
r43 2 14 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=2.515 $X2=2.49 $Y2=2.37
r44 1 11 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.595 $X2=2.785 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_2%Q 1 2 9 11
r21 11 17 9.96707 $w=3.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.33 $Y=1.665
+ $X2=8.33 $Y2=1.985
r22 11 14 3.97169 $w=3.68e-07 $l=1.15e-07 $layer=LI1_cond $X=8.33 $Y=1.665
+ $X2=8.33 $Y2=1.55
r23 9 14 38.3518 $w=3.03e-07 $l=1.015e-06 $layer=LI1_cond $X=8.297 $Y=0.535
+ $X2=8.297 $Y2=1.55
r24 2 17 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.175
+ $Y=1.84 $X2=8.31 $Y2=1.985
r25 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.145
+ $Y=0.39 $X2=8.285 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_2%Q_N 1 2 9 13 14 15 16 23 32
r31 21 23 1.04193 $w=3.63e-07 $l=3.3e-08 $layer=LI1_cond $X=10.322 $Y=2.002
+ $X2=10.322 $Y2=2.035
r32 15 16 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=10.322 $Y=2.405
+ $X2=10.322 $Y2=2.775
r33 14 21 0.820918 $w=3.63e-07 $l=2.6e-08 $layer=LI1_cond $X=10.322 $Y=1.976
+ $X2=10.322 $Y2=2.002
r34 14 32 8.24014 $w=3.63e-07 $l=1.56e-07 $layer=LI1_cond $X=10.322 $Y=1.976
+ $X2=10.322 $Y2=1.82
r35 14 15 10.8614 $w=3.63e-07 $l=3.44e-07 $layer=LI1_cond $X=10.322 $Y=2.061
+ $X2=10.322 $Y2=2.405
r36 14 23 0.820918 $w=3.63e-07 $l=2.6e-08 $layer=LI1_cond $X=10.322 $Y=2.061
+ $X2=10.322 $Y2=2.035
r37 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=10.42 $Y=1.13
+ $X2=10.42 $Y2=1.82
r38 7 13 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=10.335 $Y=0.96
+ $X2=10.335 $Y2=1.13
r39 7 9 15.0834 $w=3.38e-07 $l=4.45e-07 $layer=LI1_cond $X=10.335 $Y=0.96
+ $X2=10.335 $Y2=0.515
r40 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.17
+ $Y=1.84 $X2=10.305 $Y2=1.985
r41 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.17
+ $Y=1.84 $X2=10.305 $Y2=2.815
r42 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.19
+ $Y=0.37 $X2=10.33 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFXBP_2%VGND 1 2 3 4 5 6 7 8 27 31 33 37 41 45 49 53
+ 57 59 62 63 65 66 68 69 70 72 77 95 99 105 108 111 114 118
c141 31 0 6.63922e-20 $X=2.025 $Y=0.475
r142 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r143 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r144 111 112 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r145 109 112 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=4.08 $Y2=0
r146 108 109 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r147 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r148 103 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r149 103 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r150 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r151 100 114 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.985 $Y=0
+ $X2=9.86 $Y2=0
r152 100 102 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.985 $Y=0
+ $X2=10.32 $Y2=0
r153 99 117 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=10.675 $Y=0
+ $X2=10.857 $Y2=0
r154 99 102 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=10.675 $Y=0
+ $X2=10.32 $Y2=0
r155 98 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r156 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r157 95 114 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.735 $Y=0
+ $X2=9.86 $Y2=0
r158 95 97 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=9.735 $Y=0
+ $X2=9.36 $Y2=0
r159 94 98 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r160 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r161 91 94 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=8.4
+ $Y2=0
r162 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r163 88 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r164 87 88 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r165 85 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=4.08 $Y2=0
r166 84 87 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6.48
+ $Y2=0
r167 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r168 82 111 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.37 $Y=0 $X2=4.2
+ $Y2=0
r169 82 84 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.37 $Y=0 $X2=4.56
+ $Y2=0
r170 81 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r171 81 106 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=0.72 $Y2=0
r172 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r173 78 105 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.01 $Y=0
+ $X2=0.817 $Y2=0
r174 78 80 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=1.68
+ $Y2=0
r175 77 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.86 $Y=0
+ $X2=2.025 $Y2=0
r176 77 80 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=1.68
+ $Y2=0
r177 75 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r178 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r179 72 105 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.817 $Y2=0
r180 72 74 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r181 70 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r182 70 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r183 68 93 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.62 $Y=0 $X2=8.4
+ $Y2=0
r184 68 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.62 $Y=0 $X2=8.785
+ $Y2=0
r185 67 97 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=8.95 $Y=0 $X2=9.36
+ $Y2=0
r186 67 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.95 $Y=0 $X2=8.785
+ $Y2=0
r187 65 90 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.645 $Y=0
+ $X2=7.44 $Y2=0
r188 65 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.645 $Y=0 $X2=7.81
+ $Y2=0
r189 64 93 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=7.975 $Y=0 $X2=8.4
+ $Y2=0
r190 64 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.975 $Y=0 $X2=7.81
+ $Y2=0
r191 62 87 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.655 $Y=0
+ $X2=6.48 $Y2=0
r192 62 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.655 $Y=0 $X2=6.82
+ $Y2=0
r193 61 90 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=6.985 $Y=0
+ $X2=7.44 $Y2=0
r194 61 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.985 $Y=0 $X2=6.82
+ $Y2=0
r195 57 117 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.8 $Y=0.085
+ $X2=10.857 $Y2=0
r196 57 59 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.8 $Y=0.085
+ $X2=10.8 $Y2=0.515
r197 53 55 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=9.86 $Y=0.515
+ $X2=9.86 $Y2=0.965
r198 51 114 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.86 $Y=0.085
+ $X2=9.86 $Y2=0
r199 51 53 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.86 $Y=0.085
+ $X2=9.86 $Y2=0.515
r200 47 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.785 $Y=0.085
+ $X2=8.785 $Y2=0
r201 47 49 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=8.785 $Y=0.085
+ $X2=8.785 $Y2=0.535
r202 43 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.81 $Y=0.085
+ $X2=7.81 $Y2=0
r203 43 45 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=7.81 $Y=0.085
+ $X2=7.81 $Y2=0.535
r204 39 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.82 $Y=0.085
+ $X2=6.82 $Y2=0
r205 39 41 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=6.82 $Y=0.085
+ $X2=6.82 $Y2=0.81
r206 35 111 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.2 $Y=0.085
+ $X2=4.2 $Y2=0
r207 35 37 14.914 $w=3.38e-07 $l=4.4e-07 $layer=LI1_cond $X=4.2 $Y=0.085 $X2=4.2
+ $Y2=0.525
r208 34 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.19 $Y=0
+ $X2=2.025 $Y2=0
r209 33 111 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.03 $Y=0 $X2=4.2
+ $Y2=0
r210 33 34 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.03 $Y=0 $X2=2.19
+ $Y2=0
r211 29 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0
r212 29 31 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0.475
r213 25 105 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.817 $Y=0.085
+ $X2=0.817 $Y2=0
r214 25 27 9.27941 $w=3.83e-07 $l=3.1e-07 $layer=LI1_cond $X=0.817 $Y=0.085
+ $X2=0.817 $Y2=0.395
r215 8 59 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.62
+ $Y=0.37 $X2=10.76 $Y2=0.515
r216 7 55 182 $w=1.7e-07 $l=5.20913e-07 $layer=licon1_NDIFF $count=1 $X=9.635
+ $Y=0.56 $X2=9.9 $Y2=0.965
r217 7 53 182 $w=1.7e-07 $l=2.86618e-07 $layer=licon1_NDIFF $count=1 $X=9.635
+ $Y=0.56 $X2=9.9 $Y2=0.515
r218 6 49 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=8.575
+ $Y=0.39 $X2=8.785 $Y2=0.535
r219 5 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.67
+ $Y=0.39 $X2=7.81 $Y2=0.535
r220 4 41 182 $w=1.7e-07 $l=2.92916e-07 $layer=licon1_NDIFF $count=1 $X=6.6
+ $Y=0.64 $X2=6.82 $Y2=0.81
r221 3 37 182 $w=1.7e-07 $l=2.32379e-07 $layer=licon1_NDIFF $count=1 $X=3.975
+ $Y=0.51 $X2=4.2 $Y2=0.525
r222 2 31 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=1.88
+ $Y=0.33 $X2=2.025 $Y2=0.475
r223 1 27 182 $w=1.7e-07 $l=2.57196e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.815 $Y2=0.395
.ends


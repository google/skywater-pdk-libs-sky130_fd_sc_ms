* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 a_511_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 VGND A2 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 VGND A2 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VPWR A1 a_1291_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X4 Y C1 a_27_84# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_27_84# B1 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_1291_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 a_483_74# B1 a_27_84# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_483_74# B2 a_27_84# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X11 Y B2 a_511_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X12 a_483_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_483_74# B1 a_27_84# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 VPWR A1 a_1291_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 a_1291_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X16 a_511_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X17 a_27_84# B2 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 a_1291_368# A2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X19 VPWR B1 a_511_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X20 a_511_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X21 a_511_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X22 a_1291_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X23 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X24 a_27_84# C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X26 a_483_74# B2 a_27_84# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 a_483_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X28 a_483_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X29 a_27_84# C1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X30 VPWR B1 a_511_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X31 Y A2 a_1291_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X32 Y C1 a_27_84# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X33 VGND A1 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X34 VGND A1 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X35 Y B2 a_511_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X36 a_27_84# B2 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X37 a_27_84# B1 a_483_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X38 a_483_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X39 Y A2 a_1291_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
.ends

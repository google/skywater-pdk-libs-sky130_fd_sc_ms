* File: sky130_fd_sc_ms__sdfxtp_1.spice
* Created: Fri Aug 28 18:14:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdfxtp_1.pex.spice"
.subckt sky130_fd_sc_ms__sdfxtp_1  VNB VPB SCE D SCD CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_SCE_M1006_g N_A_35_74#_M1006_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.07455 AS=0.1197 PD=0.775 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1020 A_223_74# N_A_35_74#_M1020_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.07455 PD=0.66 PS=0.775 NRD=18.564 NRS=21.42 M=1 R=2.8
+ SA=75000.7 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1021 N_A_301_74#_M1021_d N_D_M1021_g A_223_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.12495 AS=0.0504 PD=1.015 PS=0.66 NRD=48.564 NRS=18.564 M=1 R=2.8
+ SA=75001.1 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1029 A_450_74# N_SCE_M1029_g N_A_301_74#_M1021_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.12495 PD=0.66 PS=1.015 NRD=18.564 NRS=41.424 M=1 R=2.8
+ SA=75001.8 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1028 N_VGND_M1028_d N_SCD_M1028_g A_450_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0877655 AS=0.0504 PD=0.796552 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8
+ SA=75002.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1003 N_A_630_74#_M1003_d N_CLK_M1003_g N_VGND_M1028_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.154634 PD=2.05 PS=1.40345 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1018 N_A_828_74#_M1018_d N_A_630_74#_M1018_g N_VGND_M1018_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1961 AS=0.2109 PD=2.01 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_A_1018_100#_M1007_d N_A_630_74#_M1007_g N_A_301_74#_M1007_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1113 PD=0.95 PS=1.37 NRD=71.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.8 A=0.063 P=1.14 MULT=1
MM1030 A_1154_100# N_A_828_74#_M1030_g N_A_1018_100#_M1007_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.08925 AS=0.1113 PD=0.845 PS=0.95 NRD=45 NRS=0 M=1 R=2.8 SA=75000.9
+ SB=75004.1 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_A_1239_74#_M1024_g A_1154_100# VNB NLOWVT L=0.15 W=0.42
+ AD=0.174387 AS=0.08925 PD=1.19505 PS=0.845 NRD=102.912 NRS=45 M=1 R=2.8
+ SA=75001.4 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1011 N_A_1239_74#_M1011_d N_A_1018_100#_M1011_g N_VGND_M1024_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.078375 AS=0.228363 PD=0.835 PS=1.56495 NRD=1.08 NRS=72 M=1
+ R=3.66667 SA=75001.9 SB=75002.2 A=0.0825 P=1.4 MULT=1
MM1000 N_A_1520_74#_M1000_d N_A_828_74#_M1000_g N_A_1239_74#_M1011_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.182747 AS=0.078375 PD=1.40619 PS=0.835 NRD=89.448 NRS=0 M=1
+ R=3.66667 SA=75002.3 SB=75001.8 A=0.0825 P=1.4 MULT=1
MM1023 A_1688_100# N_A_630_74#_M1023_g N_A_1520_74#_M1000_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.139553 PD=0.66 PS=1.07381 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75003.5 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_1736_74#_M1005_g A_1688_100# VNB NLOWVT L=0.15 W=0.42
+ AD=0.140462 AS=0.0504 PD=1.07814 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75003.9
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1009 N_A_1736_74#_M1009_d N_A_1520_74#_M1009_g N_VGND_M1005_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.14575 AS=0.183938 PD=1.63 PS=1.41186 NRD=0 NRS=15.264 M=1
+ R=3.66667 SA=75003.7 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1017 N_Q_M1017_d N_A_1736_74#_M1017_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2035 AS=0.1998 PD=2.03 PS=2.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1014 N_VPWR_M1014_d N_SCE_M1014_g N_A_35_74#_M1014_s VPB PSHORT L=0.18 W=0.64
+ AD=0.1024 AS=0.1792 PD=0.96 PS=1.84 NRD=13.8491 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90002.8 A=0.1152 P=1.64 MULT=1
MM1012 A_241_464# N_SCE_M1012_g N_VPWR_M1014_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.1024 PD=0.88 PS=0.96 NRD=19.9955 NRS=0 M=1 R=3.55556 SA=90000.7
+ SB=90002.3 A=0.1152 P=1.64 MULT=1
MM1025 N_A_301_74#_M1025_d N_D_M1025_g A_241_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.0864 AS=0.0768 PD=0.91 PS=0.88 NRD=0 NRS=19.9955 M=1 R=3.55556 SA=90001.1
+ SB=90001.9 A=0.1152 P=1.64 MULT=1
MM1027 A_415_464# N_A_35_74#_M1027_g N_A_301_74#_M1025_d VPB PSHORT L=0.18
+ W=0.64 AD=0.1152 AS=0.0864 PD=1 PS=0.91 NRD=38.4741 NRS=0 M=1 R=3.55556
+ SA=90001.6 SB=90001.4 A=0.1152 P=1.64 MULT=1
MM1002 N_VPWR_M1002_d N_SCD_M1002_g A_415_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.166982 AS=0.1152 PD=1.2 PS=1 NRD=50.7866 NRS=38.4741 M=1 R=3.55556
+ SA=90002.1 SB=90000.9 A=0.1152 P=1.64 MULT=1
MM1004 N_A_630_74#_M1004_d N_CLK_M1004_g N_VPWR_M1002_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.292218 PD=2.8 PS=2.1 NRD=0 NRS=14.9326 M=1 R=6.22222 SA=90001.7
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1008 N_A_828_74#_M1008_d N_A_630_74#_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.5152 PD=2.8 PS=3.16 NRD=0 NRS=14.9326 M=1 R=6.22222
+ SA=90000.4 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1015 N_A_1018_100#_M1015_d N_A_828_74#_M1015_g N_A_301_74#_M1015_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0672 AS=0.1176 PD=0.74 PS=1.4 NRD=21.0987 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90004.3 A=0.0756 P=1.2 MULT=1
MM1013 A_1205_508# N_A_630_74#_M1013_g N_A_1018_100#_M1015_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0462 AS=0.0672 PD=0.64 PS=0.74 NRD=25.7873 NRS=0 M=1 R=2.33333
+ SA=90000.7 SB=90003.8 A=0.0756 P=1.2 MULT=1
MM1019 N_VPWR_M1019_d N_A_1239_74#_M1019_g A_1205_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.1169 AS=0.0462 PD=0.993333 PS=0.64 NRD=39.8531 NRS=25.7873 M=1 R=2.33333
+ SA=90001.1 SB=90003.4 A=0.0756 P=1.2 MULT=1
MM1016 N_A_1239_74#_M1016_d N_A_1018_100#_M1016_g N_VPWR_M1019_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2205 AS=0.2338 PD=1.365 PS=1.98667 NRD=0 NRS=52.3626 M=1
+ R=4.66667 SA=90000.9 SB=90001.9 A=0.1512 P=2.04 MULT=1
MM1026 N_A_1520_74#_M1026_d N_A_630_74#_M1026_g N_A_1239_74#_M1016_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2492 AS=0.2205 PD=1.82 PS=1.365 NRD=18.7544 NRS=55.1009 M=1
+ R=4.66667 SA=90001.6 SB=90001.2 A=0.1512 P=2.04 MULT=1
MM1010 A_1691_508# N_A_828_74#_M1010_g N_A_1520_74#_M1026_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.1246 PD=0.66 PS=0.91 NRD=30.4759 NRS=77.3816 M=1
+ R=2.33333 SA=90003.1 SB=90001.4 A=0.0756 P=1.2 MULT=1
MM1022 N_VPWR_M1022_d N_A_1736_74#_M1022_g A_1691_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.1141 AS=0.0504 PD=0.936667 PS=0.66 NRD=53.9386 NRS=30.4759 M=1 R=2.33333
+ SA=90003.5 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1031 N_A_1736_74#_M1031_d N_A_1520_74#_M1031_g N_VPWR_M1022_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2352 AS=0.2282 PD=2.24 PS=1.87333 NRD=0 NRS=39.8531 M=1
+ R=4.66667 SA=90002.2 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1001 N_Q_M1001_d N_A_1736_74#_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.308 AS=0.3136 PD=2.79 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX32_noxref VNB VPB NWDIODE A=21.2412 P=26.56
c_125 VNB 0 2.44411e-19 $X=0 $Y=0
c_225 VPB 0 3.09632e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__sdfxtp_1.pxi.spice"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
X0 Y a_62_94# a_241_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 VGND a_62_94# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 VPWR A1 a_241_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 VPWR B1_N a_62_94# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X4 a_436_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_62_94# B1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 VPWR A2 a_241_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 Y A1 a_436_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_241_368# a_62_94# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X9 VGND A2 a_436_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_241_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X11 a_241_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X12 Y a_62_94# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_436_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

* File: sky130_fd_sc_ms__sdfrtp_2.pex.spice
* Created: Wed Sep  2 12:30:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SDFRTP_2%A_27_74# 1 2 7 9 11 14 18 21 24 28 31 33 34
+ 36 37 41
c83 31 0 3.64595e-20 $X=2.375 $Y=2.09
c84 9 0 3.56444e-20 $X=1.485 $Y=0.935
r85 37 47 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.5 $Y=1.995
+ $X2=2.5 $Y2=2.16
r86 36 39 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.54 $Y=1.995
+ $X2=2.54 $Y2=2.09
r87 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.5
+ $Y=1.995 $X2=2.5 $Y2=1.995
r88 32 34 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.09
+ $X2=0.28 $Y2=2.09
r89 31 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=2.09
+ $X2=2.54 $Y2=2.09
r90 31 32 125.914 $w=1.68e-07 $l=1.93e-06 $layer=LI1_cond $X=2.375 $Y=2.09
+ $X2=0.445 $Y2=2.09
r91 29 41 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.975 $Y=1.1 $X2=0.975
+ $Y2=1.01
r92 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.1 $X2=0.975 $Y2=1.1
r93 26 33 0.221902 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=1.1
+ $X2=0.24 $Y2=1.1
r94 26 28 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=0.365 $Y=1.1
+ $X2=0.975 $Y2=1.1
r95 22 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.175
+ $X2=0.28 $Y2=2.09
r96 22 24 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=0.28 $Y=2.175
+ $X2=0.28 $Y2=2.465
r97 21 34 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.2 $Y=2.005
+ $X2=0.28 $Y2=2.09
r98 20 33 7.38875 $w=2.1e-07 $l=1.83916e-07 $layer=LI1_cond $X=0.2 $Y=1.265
+ $X2=0.24 $Y2=1.1
r99 20 21 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.2 $Y=1.265 $X2=0.2
+ $Y2=2.005
r100 16 33 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=0.935
+ $X2=0.24 $Y2=1.1
r101 16 18 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=0.24 $Y=0.935
+ $X2=0.24 $Y2=0.58
r102 14 47 223.508 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.495 $Y=2.735
+ $X2=2.495 $Y2=2.16
r103 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.485 $Y=0.935
+ $X2=1.485 $Y2=0.615
r104 8 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.01
+ $X2=0.975 $Y2=1.01
r105 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.41 $Y=1.01
+ $X2=1.485 $Y2=0.935
r106 7 8 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.41 $Y=1.01 $X2=1.14
+ $Y2=1.01
r107 2 24 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.465
r108 1 18 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_2%SCE 3 7 11 17 19 20 21 22 23 26 27 31 32 33
+ 45 47 56 58
c85 27 0 3.38289e-19 $X=2.5 $Y=1.425
r86 47 56 1.90404 $w=3.43e-07 $l=5.7e-08 $layer=LI1_cond $X=1.623 $Y=1.662
+ $X2=1.68 $Y2=1.662
r87 42 43 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.45
+ $Y=1.67 $X2=1.45 $Y2=1.67
r88 39 42 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=0.77 $Y=1.67
+ $X2=1.45 $Y2=1.67
r89 33 58 6.34154 $w=3.43e-07 $l=1.01e-07 $layer=LI1_cond $X=1.694 $Y=1.662
+ $X2=1.795 $Y2=1.662
r90 33 56 0.467658 $w=3.43e-07 $l=1.4e-08 $layer=LI1_cond $X=1.694 $Y=1.662
+ $X2=1.68 $Y2=1.662
r91 33 47 0.467658 $w=3.43e-07 $l=1.4e-08 $layer=LI1_cond $X=1.609 $Y=1.662
+ $X2=1.623 $Y2=1.662
r92 33 43 5.31126 $w=3.43e-07 $l=1.59e-07 $layer=LI1_cond $X=1.609 $Y=1.662
+ $X2=1.45 $Y2=1.662
r93 32 43 8.35104 $w=3.43e-07 $l=2.5e-07 $layer=LI1_cond $X=1.2 $Y=1.662
+ $X2=1.45 $Y2=1.662
r94 31 32 16.034 $w=3.43e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.662 $X2=1.2
+ $Y2=1.662
r95 31 39 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.77
+ $Y=1.67 $X2=0.77 $Y2=1.67
r96 27 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.5 $Y=1.425
+ $X2=2.5 $Y2=1.26
r97 26 29 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.54 $Y=1.425
+ $X2=2.54 $Y2=1.575
r98 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.5
+ $Y=1.425 $X2=2.5 $Y2=1.425
r99 23 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=1.575
+ $X2=2.54 $Y2=1.575
r100 23 58 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=2.375 $Y=1.575
+ $X2=1.795 $Y2=1.575
r101 22 45 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.59 $Y=1.05
+ $X2=2.59 $Y2=1.26
r102 21 22 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.625 $Y=0.9
+ $X2=2.625 $Y2=1.05
r103 20 42 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=1.535 $Y=1.67
+ $X2=1.45 $Y2=1.67
r104 18 39 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=0.595 $Y=1.67
+ $X2=0.77 $Y2=1.67
r105 18 19 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.595 $Y=1.67
+ $X2=0.505 $Y2=1.67
r106 17 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.66 $Y=0.615
+ $X2=2.66 $Y2=0.9
r107 9 20 30.0773 $w=3.3e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.625 $Y=1.835
+ $X2=1.535 $Y2=1.67
r108 9 11 349.839 $w=1.8e-07 $l=9e-07 $layer=POLY_cond $X=1.625 $Y=1.835
+ $X2=1.625 $Y2=2.735
r109 5 19 34.7346 $w=1.65e-07 $l=1.69926e-07 $layer=POLY_cond $X=0.495 $Y=1.505
+ $X2=0.505 $Y2=1.67
r110 5 7 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.495 $Y=1.505
+ $X2=0.495 $Y2=0.58
r111 1 19 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.835
+ $X2=0.505 $Y2=1.67
r112 1 3 312.911 $w=1.8e-07 $l=8.05e-07 $layer=POLY_cond $X=0.505 $Y=1.835
+ $X2=0.505 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_2%D 3 6 8 11 12 13
r44 11 14 40.8147 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.947 $Y=1.1
+ $X2=1.947 $Y2=1.265
r45 11 13 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.947 $Y=1.1
+ $X2=1.947 $Y2=0.935
r46 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.1 $X2=1.935 $Y2=1.1
r47 8 12 6.7033 $w=4.53e-07 $l=2.55e-07 $layer=LI1_cond $X=1.68 $Y=1.037
+ $X2=1.935 $Y2=1.037
r48 6 14 571.403 $w=1.8e-07 $l=1.47e-06 $layer=POLY_cond $X=2.035 $Y=2.735
+ $X2=2.035 $Y2=1.265
r49 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.875 $Y=0.615
+ $X2=1.875 $Y2=0.935
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_2%SCD 3 7 11 12 13 14 18
c48 13 0 1.16038e-19 $X=3.12 $Y=1.665
c49 3 0 8.88027e-20 $X=3.035 $Y=2.735
r50 13 14 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=3.11 $Y=1.645
+ $X2=3.11 $Y2=2.035
r51 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.04
+ $Y=1.645 $X2=3.04 $Y2=1.645
r52 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.04 $Y=1.985
+ $X2=3.04 $Y2=1.645
r53 11 12 34.9753 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.04 $Y=1.985
+ $X2=3.04 $Y2=2.15
r54 10 18 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.04 $Y=1.48
+ $X2=3.04 $Y2=1.645
r55 7 10 443.543 $w=1.5e-07 $l=8.65e-07 $layer=POLY_cond $X=3.05 $Y=0.615
+ $X2=3.05 $Y2=1.48
r56 3 12 227.395 $w=1.8e-07 $l=5.85e-07 $layer=POLY_cond $X=3.035 $Y=2.735
+ $X2=3.035 $Y2=2.15
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_2%CLK 1 5 8 10 13 18 19
c60 19 0 1.40651e-19 $X=4.565 $Y=1.41
c61 18 0 3.36092e-20 $X=4.565 $Y=1.51
c62 13 0 1.8717e-19 $X=3.94 $Y=1.445
c63 10 0 2.36685e-20 $X=4.08 $Y=1.295
r64 21 23 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=4.565 $Y=1.61
+ $X2=4.565 $Y2=1.775
r65 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.56
+ $Y=1.61 $X2=4.56 $Y2=1.61
r66 18 21 16.9718 $w=3.4e-07 $l=1e-07 $layer=POLY_cond $X=4.565 $Y=1.51
+ $X2=4.565 $Y2=1.61
r67 18 19 35.2748 $w=3.4e-07 $l=1e-07 $layer=POLY_cond $X=4.565 $Y=1.51
+ $X2=4.565 $Y2=1.41
r68 13 16 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=3.94 $Y=1.445
+ $X2=3.94 $Y2=1.51
r69 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.94
+ $Y=1.445 $X2=3.94 $Y2=1.445
r70 10 22 10.6473 $w=5.5e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=1.395
+ $X2=4.56 $Y2=1.395
r71 10 14 3.10545 $w=5.5e-07 $l=1.4e-07 $layer=LI1_cond $X=4.08 $Y=1.395
+ $X2=3.94 $Y2=1.395
r72 8 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.645 $Y=2.495
+ $X2=4.645 $Y2=1.775
r73 5 19 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.54 $Y=0.965
+ $X2=4.54 $Y2=1.41
r74 2 16 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.105 $Y=1.51 $X2=3.94
+ $Y2=1.51
r75 1 18 15.178 $w=2e-07 $l=1.7e-07 $layer=POLY_cond $X=4.395 $Y=1.51 $X2=4.565
+ $Y2=1.51
r76 1 2 96.1574 $w=2e-07 $l=2.9e-07 $layer=POLY_cond $X=4.395 $Y=1.51 $X2=4.105
+ $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_2%A_1037_119# 1 2 9 11 13 15 17 19 20 21 24
+ 30 32 33 34 37 40 43 44 45 47 48 49 52 55 60 62 65 69 79
c214 60 0 1.82923e-19 $X=5.32 $Y=1.11
c215 52 0 8.16714e-20 $X=9.645 $Y=1.17
c216 49 0 6.41644e-20 $X=9.26 $Y=1.17
c217 48 0 1.18082e-19 $X=9.785 $Y=1.17
c218 34 0 9.49943e-20 $X=5.42 $Y=0.365
c219 33 0 1.34587e-19 $X=7.015 $Y=0.365
c220 32 0 3.36092e-20 $X=5.502 $Y=1.635
c221 24 0 7.04642e-20 $X=10.11 $Y=2.75
c222 20 0 6.19065e-20 $X=9.48 $Y=1.26
r223 65 67 14.4055 $w=2.38e-07 $l=3e-07 $layer=LI1_cond $X=7.135 $Y=0.365
+ $X2=7.135 $Y2=0.665
r224 62 64 11.426 $w=3.31e-07 $l=3.1e-07 $layer=LI1_cond $X=5.387 $Y=1.8
+ $X2=5.387 $Y2=2.11
r225 60 61 8.16324 $w=2.72e-07 $l=1.82e-07 $layer=LI1_cond $X=5.32 $Y=1.07
+ $X2=5.502 $Y2=1.07
r226 58 60 1.12132 $w=2.72e-07 $l=2.5e-08 $layer=LI1_cond $X=5.295 $Y=1.07
+ $X2=5.32 $Y2=1.07
r227 56 79 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=9.95 $Y=2.165
+ $X2=10.11 $Y2=2.165
r228 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.95
+ $Y=2.165 $X2=9.95 $Y2=2.165
r229 53 55 36.0954 $w=2.63e-07 $l=8.3e-07 $layer=LI1_cond $X=9.917 $Y=1.335
+ $X2=9.917 $Y2=2.165
r230 52 75 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.645 $Y=1.17
+ $X2=9.645 $Y2=1.26
r231 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.645
+ $Y=1.17 $X2=9.645 $Y2=1.17
r232 49 51 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=9.26 $Y=1.17
+ $X2=9.645 $Y2=1.17
r233 48 53 6.92284 $w=3.3e-07 $l=2.21371e-07 $layer=LI1_cond $X=9.785 $Y=1.17
+ $X2=9.917 $Y2=1.335
r234 48 51 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=9.785 $Y=1.17
+ $X2=9.645 $Y2=1.17
r235 47 49 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.175 $Y=1.005
+ $X2=9.26 $Y2=1.17
r236 46 47 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=9.175 $Y=0.425
+ $X2=9.175 $Y2=1.005
r237 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.09 $Y=0.34
+ $X2=9.175 $Y2=0.425
r238 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.09 $Y=0.34
+ $X2=8.42 $Y2=0.34
r239 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.335 $Y=0.425
+ $X2=8.42 $Y2=0.34
r240 42 43 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=8.335 $Y=0.425
+ $X2=8.335 $Y2=0.58
r241 41 67 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.255 $Y=0.665
+ $X2=7.135 $Y2=0.665
r242 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.25 $Y=0.665
+ $X2=8.335 $Y2=0.58
r243 40 41 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=8.25 $Y=0.665
+ $X2=7.255 $Y2=0.665
r244 38 72 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.065 $Y=1.8
+ $X2=6.065 $Y2=1.965
r245 38 69 20.6336 $w=3.3e-07 $l=1.18e-07 $layer=POLY_cond $X=6.065 $Y=1.8
+ $X2=6.065 $Y2=1.682
r246 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.065
+ $Y=1.8 $X2=6.065 $Y2=1.8
r247 35 62 0.734941 $w=3.3e-07 $l=2.33e-07 $layer=LI1_cond $X=5.62 $Y=1.8
+ $X2=5.387 $Y2=1.8
r248 35 37 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=5.62 $Y=1.8
+ $X2=6.065 $Y2=1.8
r249 33 65 1.80669 $w=2e-07 $l=1.2e-07 $layer=LI1_cond $X=7.015 $Y=0.365
+ $X2=7.135 $Y2=0.365
r250 33 34 88.45 $w=1.98e-07 $l=1.595e-06 $layer=LI1_cond $X=7.015 $Y=0.365
+ $X2=5.42 $Y2=0.365
r251 32 62 7.12462 $w=3.31e-07 $l=2.14942e-07 $layer=LI1_cond $X=5.502 $Y=1.635
+ $X2=5.387 $Y2=1.8
r252 31 61 1.61602 $w=2.35e-07 $l=1.5e-07 $layer=LI1_cond $X=5.502 $Y=1.22
+ $X2=5.502 $Y2=1.07
r253 31 32 20.3517 $w=2.33e-07 $l=4.15e-07 $layer=LI1_cond $X=5.502 $Y=1.22
+ $X2=5.502 $Y2=1.635
r254 28 58 1.22563 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=5.295 $Y=0.92
+ $X2=5.295 $Y2=1.07
r255 28 30 8.29759 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=5.295 $Y=0.92
+ $X2=5.295 $Y2=0.74
r256 27 34 6.92652 $w=2e-07 $l=1.67705e-07 $layer=LI1_cond $X=5.295 $Y=0.465
+ $X2=5.42 $Y2=0.365
r257 27 30 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=5.295 $Y=0.465
+ $X2=5.295 $Y2=0.74
r258 22 79 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.11 $Y=2.33
+ $X2=10.11 $Y2=2.165
r259 22 24 163.258 $w=1.8e-07 $l=4.2e-07 $layer=POLY_cond $X=10.11 $Y=2.33
+ $X2=10.11 $Y2=2.75
r260 20 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.48 $Y=1.26
+ $X2=9.645 $Y2=1.26
r261 20 21 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=9.48 $Y=1.26
+ $X2=9.12 $Y2=1.26
r262 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.045 $Y=1.185
+ $X2=9.12 $Y2=1.26
r263 17 19 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=9.045 $Y=1.185
+ $X2=9.045 $Y2=0.74
r264 13 26 74.7716 $w=2.28e-07 $l=3.62566e-07 $layer=POLY_cond $X=6.695 $Y=1.355
+ $X2=6.62 $Y2=1.682
r265 13 15 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.695 $Y=1.355
+ $X2=6.695 $Y2=0.805
r266 12 69 13.99 $w=2.05e-07 $l=1.65e-07 $layer=POLY_cond $X=6.23 $Y=1.682
+ $X2=6.065 $Y2=1.682
r267 11 26 5.46652 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=6.47 $Y=1.682
+ $X2=6.62 $Y2=1.682
r268 11 12 77.6376 $w=2.05e-07 $l=2.4e-07 $layer=POLY_cond $X=6.47 $Y=1.682
+ $X2=6.23 $Y2=1.682
r269 9 72 206.016 $w=1.8e-07 $l=5.3e-07 $layer=POLY_cond $X=6.135 $Y=2.495
+ $X2=6.135 $Y2=1.965
r270 2 64 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=5.185
+ $Y=1.935 $X2=5.32 $Y2=2.11
r271 1 60 182 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_NDIFF $count=1 $X=5.185
+ $Y=0.595 $X2=5.32 $Y2=1.11
r272 1 30 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.185
+ $Y=0.595 $X2=5.32 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_2%A_1383_349# 1 2 9 13 17 18 20 21 26 29 34
+ 35
c92 21 0 1.25732e-19 $X=7.315 $Y=1.005
c93 13 0 1.40848e-19 $X=7.085 $Y=0.805
r94 36 38 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=7.005 $Y=1.91
+ $X2=7.085 $Y2=1.91
r95 34 35 8.52431 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=8.932 $Y=1.88
+ $X2=8.932 $Y2=1.715
r96 32 35 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=8.835 $Y=1.13
+ $X2=8.835 $Y2=1.715
r97 31 32 7.06528 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=8.755 $Y=1.005
+ $X2=8.755 $Y2=1.13
r98 29 31 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=8.755 $Y=0.86
+ $X2=8.755 $Y2=1.005
r99 24 34 0.536754 $w=3.63e-07 $l=1.7e-08 $layer=LI1_cond $X=8.932 $Y=1.897
+ $X2=8.932 $Y2=1.88
r100 24 26 10.6719 $w=3.63e-07 $l=3.38e-07 $layer=LI1_cond $X=8.932 $Y=1.897
+ $X2=8.932 $Y2=2.235
r101 20 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.59 $Y=1.005
+ $X2=8.755 $Y2=1.005
r102 20 21 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=8.59 $Y=1.005
+ $X2=7.315 $Y2=1.005
r103 18 38 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=7.165 $Y=1.91
+ $X2=7.085 $Y2=1.91
r104 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.165
+ $Y=1.91 $X2=7.165 $Y2=1.91
r105 15 21 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=7.177 $Y=1.09
+ $X2=7.315 $Y2=1.005
r106 15 17 34.3638 $w=2.73e-07 $l=8.2e-07 $layer=LI1_cond $X=7.177 $Y=1.09
+ $X2=7.177 $Y2=1.91
r107 11 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.085 $Y=1.745
+ $X2=7.085 $Y2=1.91
r108 11 13 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=7.085 $Y=1.745
+ $X2=7.085 $Y2=0.805
r109 7 36 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.005 $Y=2.075
+ $X2=7.005 $Y2=1.91
r110 7 9 163.258 $w=1.8e-07 $l=4.2e-07 $layer=POLY_cond $X=7.005 $Y=2.075
+ $X2=7.005 $Y2=2.495
r111 2 34 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=8.73
+ $Y=1.735 $X2=8.95 $Y2=1.88
r112 2 26 300 $w=1.7e-07 $l=6e-07 $layer=licon1_PDIFF $count=2 $X=8.73 $Y=1.735
+ $X2=8.95 $Y2=2.235
r113 1 29 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=8.615
+ $Y=0.37 $X2=8.755 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_2%RESET_B 2 5 10 11 12 16 19 22 25 29 32 34
+ 37 39 40 41 42 49 50 53 54 60 65 76
c220 41 0 1.13179e-19 $X=11.135 $Y=2.035
c221 11 0 1.68004e-19 $X=7.4 $Y=0.18
r222 65 67 11.8137 $w=3.06e-07 $l=7.5e-08 $layer=POLY_cond $X=11.275 $Y=2.07
+ $X2=11.35 $Y2=2.07
r223 65 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.275
+ $Y=2.07 $X2=11.275 $Y2=2.07
r224 63 65 22.0523 $w=3.06e-07 $l=1.4e-07 $layer=POLY_cond $X=11.135 $Y=2.07
+ $X2=11.275 $Y2=2.07
r225 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.975
+ $Y=1.96 $X2=7.975 $Y2=1.96
r226 58 60 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=7.645 $Y=1.96
+ $X2=7.975 $Y2=1.96
r227 56 58 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.63 $Y=1.96
+ $X2=7.645 $Y2=1.96
r228 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.995 $X2=3.95 $Y2=1.995
r229 50 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=2.035
+ $X2=11.28 $Y2=2.035
r230 49 61 13.7969 $w=3.53e-07 $l=4.25e-07 $layer=LI1_cond $X=8.4 $Y=1.972
+ $X2=7.975 $Y2=1.972
r231 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=2.035
+ $X2=8.4 $Y2=2.035
r232 44 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=2.035
+ $X2=4.08 $Y2=2.035
r233 42 48 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.545 $Y=2.035
+ $X2=8.4 $Y2=2.035
r234 41 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.135 $Y=2.035
+ $X2=11.28 $Y2=2.035
r235 41 42 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=11.135 $Y=2.035
+ $X2=8.545 $Y2=2.035
r236 40 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=2.035
+ $X2=4.08 $Y2=2.035
r237 39 48 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=2.035
+ $X2=8.4 $Y2=2.035
r238 39 40 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=8.255 $Y=2.035
+ $X2=4.225 $Y2=2.035
r239 35 37 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=7.475 $Y=1.26
+ $X2=7.645 $Y2=1.26
r240 33 53 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=3.595 $Y=1.995
+ $X2=3.95 $Y2=1.995
r241 33 34 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.595 $Y=1.995
+ $X2=3.505 $Y2=1.995
r242 31 32 69.9677 $w=1.75e-07 $l=1.75e-07 $layer=POLY_cond $X=3.502 $Y=0.9
+ $X2=3.502 $Y2=1.075
r243 27 67 15.178 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=11.35 $Y=2.235
+ $X2=11.35 $Y2=2.07
r244 27 29 200.185 $w=1.8e-07 $l=5.15e-07 $layer=POLY_cond $X=11.35 $Y=2.235
+ $X2=11.35 $Y2=2.75
r245 23 63 19.4347 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.135 $Y=1.905
+ $X2=11.135 $Y2=2.07
r246 23 25 679.415 $w=1.5e-07 $l=1.325e-06 $layer=POLY_cond $X=11.135 $Y=1.905
+ $X2=11.135 $Y2=0.58
r247 22 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.645 $Y=1.795
+ $X2=7.645 $Y2=1.96
r248 21 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.645 $Y=1.335
+ $X2=7.645 $Y2=1.26
r249 21 22 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=7.645 $Y=1.335
+ $X2=7.645 $Y2=1.795
r250 17 56 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.63 $Y=2.125
+ $X2=7.63 $Y2=1.96
r251 17 19 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=7.63 $Y=2.125
+ $X2=7.63 $Y2=2.495
r252 14 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.475 $Y=1.185
+ $X2=7.475 $Y2=1.26
r253 14 16 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=7.475 $Y=1.185
+ $X2=7.475 $Y2=0.805
r254 13 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7.475 $Y=0.255
+ $X2=7.475 $Y2=0.805
r255 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.4 $Y=0.18
+ $X2=7.475 $Y2=0.255
r256 11 12 1953.64 $w=1.5e-07 $l=3.81e-06 $layer=POLY_cond $X=7.4 $Y=0.18
+ $X2=3.59 $Y2=0.18
r257 10 31 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.515 $Y=0.615
+ $X2=3.515 $Y2=0.9
r258 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.515 $Y=0.255
+ $X2=3.59 $Y2=0.18
r259 7 10 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.515 $Y=0.255
+ $X2=3.515 $Y2=0.615
r260 3 34 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=3.505 $Y=2.16
+ $X2=3.505 $Y2=1.995
r261 3 5 223.508 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.505 $Y=2.16
+ $X2=3.505 $Y2=2.735
r262 2 34 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=3.49 $Y=1.83
+ $X2=3.505 $Y2=1.995
r263 2 32 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=3.49 $Y=1.83
+ $X2=3.49 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_2%A_1235_119# 1 2 3 12 16 18 19 20 25 26 29
+ 30 32 36 38
c119 20 0 1.28673e-19 $X=6.7 $Y=2.6
c120 19 0 1.13179e-19 $X=8.465 $Y=1.245
c121 12 0 6.41644e-20 $X=8.54 $Y=0.74
r122 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.255
+ $Y=1.41 $X2=8.255 $Y2=1.41
r123 30 32 21.9513 $w=3.13e-07 $l=6e-07 $layer=LI1_cond $X=7.655 $Y=1.417
+ $X2=8.255 $Y2=1.417
r124 29 41 11.0732 $w=3.14e-07 $l=3.72552e-07 $layer=LI1_cond $X=7.57 $Y=2.32
+ $X2=7.855 $Y2=2.522
r125 28 30 7.64049 $w=3.15e-07 $l=1.95944e-07 $layer=LI1_cond $X=7.57 $Y=1.575
+ $X2=7.655 $Y2=1.417
r126 28 29 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=7.57 $Y=1.575
+ $X2=7.57 $Y2=2.32
r127 27 38 4.3182 $w=2.1e-07 $l=1.53734e-07 $layer=LI1_cond $X=6.87 $Y=2.405
+ $X2=6.785 $Y2=2.522
r128 26 29 5.85116 $w=3.14e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.485 $Y=2.405
+ $X2=7.57 $Y2=2.32
r129 26 27 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=7.485 $Y=2.405
+ $X2=6.87 $Y2=2.405
r130 25 38 2.11342 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=6.785 $Y=2.32
+ $X2=6.785 $Y2=2.522
r131 24 36 10.5113 $w=3.54e-07 $l=4.07707e-07 $layer=LI1_cond $X=6.785 $Y=1.125
+ $X2=6.48 $Y2=0.885
r132 24 25 77.9626 $w=1.68e-07 $l=1.195e-06 $layer=LI1_cond $X=6.785 $Y=1.125
+ $X2=6.785 $Y2=2.32
r133 20 38 4.3182 $w=2.1e-07 $l=1.17707e-07 $layer=LI1_cond $X=6.7 $Y=2.6
+ $X2=6.785 $Y2=2.522
r134 20 22 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=6.7 $Y=2.6 $X2=6.36
+ $Y2=2.6
r135 18 33 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=8.465 $Y=1.41
+ $X2=8.255 $Y2=1.41
r136 18 19 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.465 $Y=1.41
+ $X2=8.465 $Y2=1.245
r137 14 19 34.7346 $w=1.65e-07 $l=4.08228e-07 $layer=POLY_cond $X=8.64 $Y=1.575
+ $X2=8.465 $Y2=1.245
r138 14 16 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=8.64 $Y=1.575
+ $X2=8.64 $Y2=2.235
r139 10 19 34.7346 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=8.54 $Y=1.245
+ $X2=8.465 $Y2=1.245
r140 10 12 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=8.54 $Y=1.245
+ $X2=8.54 $Y2=0.74
r141 3 41 600 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_PDIFF $count=1 $X=7.72
+ $Y=2.285 $X2=7.855 $Y2=2.52
r142 2 22 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=6.225
+ $Y=2.285 $X2=6.36 $Y2=2.56
r143 1 36 182 $w=1.7e-07 $l=3.98246e-07 $layer=licon1_NDIFF $count=1 $X=6.175
+ $Y=0.595 $X2=6.48 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_2%A_837_119# 1 2 9 12 13 16 19 20 21 22 23 24
+ 25 27 30 32 37 38 39 41 44 46 47 48 51 53 55 58 60 62 64 72 75 76 78
c203 76 0 9.49943e-20 $X=5.13 $Y=1.41
c204 75 0 4.95374e-20 $X=5.13 $Y=1.485
c205 60 0 1.21651e-19 $X=4.9 $Y=1.945
c206 20 0 1.28673e-19 $X=5.61 $Y=3.075
r207 75 76 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.13 $Y=1.485
+ $X2=5.13 $Y2=1.41
r208 73 78 55.5535 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=5.13 $Y=1.61
+ $X2=5.13 $Y2=1.86
r209 73 75 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.13 $Y=1.61
+ $X2=5.13 $Y2=1.485
r210 72 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.13
+ $Y=1.61 $X2=5.13 $Y2=1.61
r211 69 72 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=4.9 $Y=1.61
+ $X2=5.13 $Y2=1.61
r212 64 67 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.46 $Y=2.03 $X2=4.46
+ $Y2=2.11
r213 59 69 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.9 $Y=1.775
+ $X2=4.9 $Y2=1.61
r214 59 60 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.9 $Y=1.775
+ $X2=4.9 $Y2=1.945
r215 58 69 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.9 $Y=1.445
+ $X2=4.9 $Y2=1.61
r216 57 58 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.9 $Y=1.09
+ $X2=4.9 $Y2=1.445
r217 56 64 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.585 $Y=2.03
+ $X2=4.46 $Y2=2.03
r218 55 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.815 $Y=2.03
+ $X2=4.9 $Y2=1.945
r219 55 56 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.815 $Y=2.03
+ $X2=4.585 $Y2=2.03
r220 54 62 9.86469 $w=3.03e-07 $l=3.34978e-07 $layer=LI1_cond $X=4.57 $Y=1.005
+ $X2=4.357 $Y2=0.76
r221 53 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.815 $Y=1.005
+ $X2=4.9 $Y2=1.09
r222 53 54 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.815 $Y=1.005
+ $X2=4.57 $Y2=1.005
r223 49 51 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=10.125 $Y=1.055
+ $X2=10.315 $Y2=1.055
r224 42 51 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.315 $Y=0.98
+ $X2=10.315 $Y2=1.055
r225 42 44 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=10.315 $Y=0.98
+ $X2=10.315 $Y2=0.58
r226 40 49 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.125 $Y=1.13
+ $X2=10.125 $Y2=1.055
r227 40 41 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=10.125 $Y=1.13
+ $X2=10.125 $Y2=1.575
r228 38 41 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.05 $Y=1.65
+ $X2=10.125 $Y2=1.575
r229 38 39 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=10.05 $Y=1.65
+ $X2=9.35 $Y2=1.65
r230 35 37 289.589 $w=1.8e-07 $l=7.45e-07 $layer=POLY_cond $X=9.26 $Y=3.075
+ $X2=9.26 $Y2=2.33
r231 34 39 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=9.26 $Y=1.725
+ $X2=9.35 $Y2=1.65
r232 34 37 235.169 $w=1.8e-07 $l=6.05e-07 $layer=POLY_cond $X=9.26 $Y=1.725
+ $X2=9.26 $Y2=2.33
r233 33 48 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.695 $Y=3.15
+ $X2=6.605 $Y2=3.15
r234 32 35 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=9.17 $Y=3.15
+ $X2=9.26 $Y2=3.075
r235 32 33 1269.1 $w=1.5e-07 $l=2.475e-06 $layer=POLY_cond $X=9.17 $Y=3.15
+ $X2=6.695 $Y2=3.15
r236 28 48 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=6.605 $Y=3.075
+ $X2=6.605 $Y2=3.15
r237 28 30 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=6.605 $Y=3.075
+ $X2=6.605 $Y2=2.495
r238 25 27 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.1 $Y=1.09 $X2=6.1
+ $Y2=0.805
r239 23 48 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.515 $Y=3.15
+ $X2=6.605 $Y2=3.15
r240 23 24 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=6.515 $Y=3.15
+ $X2=5.69 $Y2=3.15
r241 21 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.025 $Y=1.165
+ $X2=6.1 $Y2=1.09
r242 21 22 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=6.025 $Y=1.165
+ $X2=5.68 $Y2=1.165
r243 20 24 26.9672 $w=1.5e-07 $l=1.11355e-07 $layer=POLY_cond $X=5.61 $Y=3.075
+ $X2=5.69 $Y2=3.15
r244 19 47 37.4638 $w=1.6e-07 $l=8e-08 $layer=POLY_cond $X=5.61 $Y=2.275
+ $X2=5.61 $Y2=2.195
r245 19 20 370.769 $w=1.6e-07 $l=8e-07 $layer=POLY_cond $X=5.61 $Y=2.275
+ $X2=5.61 $Y2=3.075
r246 17 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.605 $Y=1.56
+ $X2=5.605 $Y2=1.485
r247 17 47 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=5.605 $Y=1.56
+ $X2=5.605 $Y2=2.195
r248 16 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.605 $Y=1.41
+ $X2=5.605 $Y2=1.485
r249 15 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.605 $Y=1.24
+ $X2=5.68 $Y2=1.165
r250 15 16 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=5.605 $Y=1.24
+ $X2=5.605 $Y2=1.41
r251 14 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.295 $Y=1.485
+ $X2=5.13 $Y2=1.485
r252 13 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.53 $Y=1.485
+ $X2=5.605 $Y2=1.485
r253 13 14 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=5.53 $Y=1.485
+ $X2=5.295 $Y2=1.485
r254 12 76 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.11 $Y=0.965
+ $X2=5.11 $Y2=1.41
r255 9 78 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=5.095 $Y=2.495
+ $X2=5.095 $Y2=1.86
r256 2 67 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.275
+ $Y=1.935 $X2=4.42 $Y2=2.11
r257 1 62 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=4.185
+ $Y=0.595 $X2=4.31 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_2%A_2082_446# 1 2 9 13 17 21 22 23 25 26 29
+ 33 35 36 38 40 41
c119 26 0 7.04642e-20 $X=10.85 $Y=2.475
c120 21 0 1.13484e-19 $X=10.685 $Y=2.215
c121 13 0 1.18082e-19 $X=10.705 $Y=0.58
r122 41 44 5.42589 $w=4.1e-07 $l=4e-08 $layer=POLY_cond $X=10.645 $Y=1.535
+ $X2=10.645 $Y2=1.575
r123 41 47 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=10.645 $Y=1.535
+ $X2=10.645 $Y2=1.37
r124 40 43 5.16612 $w=2.88e-07 $l=1.3e-07 $layer=LI1_cond $X=10.705 $Y=1.535
+ $X2=10.705 $Y2=1.665
r125 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=10.685
+ $Y=1.535 $X2=10.685 $Y2=1.535
r126 37 38 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=12.145 $Y=0.94
+ $X2=12.145 $Y2=1.58
r127 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.06 $Y=0.855
+ $X2=12.145 $Y2=0.94
r128 35 36 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=12.06 $Y=0.855
+ $X2=11.875 $Y2=0.855
r129 31 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.71 $Y=0.77
+ $X2=11.875 $Y2=0.855
r130 31 33 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=11.71 $Y=0.77
+ $X2=11.71 $Y2=0.58
r131 27 29 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=11.575 $Y=2.56
+ $X2=11.575 $Y2=2.75
r132 25 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.41 $Y=2.475
+ $X2=11.575 $Y2=2.56
r133 25 26 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=11.41 $Y=2.475
+ $X2=10.85 $Y2=2.475
r134 24 43 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=10.85 $Y=1.665
+ $X2=10.705 $Y2=1.665
r135 23 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.06 $Y=1.665
+ $X2=12.145 $Y2=1.58
r136 23 24 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=12.06 $Y=1.665
+ $X2=10.85 $Y2=1.665
r137 22 44 86.8143 $w=4.1e-07 $l=6.4e-07 $layer=POLY_cond $X=10.645 $Y=2.215
+ $X2=10.645 $Y2=1.575
r138 21 22 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=10.685
+ $Y=2.215 $X2=10.685 $Y2=2.215
r139 19 26 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=10.705 $Y=2.39
+ $X2=10.85 $Y2=2.475
r140 19 21 6.9544 $w=2.88e-07 $l=1.75e-07 $layer=LI1_cond $X=10.705 $Y=2.39
+ $X2=10.705 $Y2=2.215
r141 18 43 3.37785 $w=2.88e-07 $l=8.5e-08 $layer=LI1_cond $X=10.705 $Y=1.75
+ $X2=10.705 $Y2=1.665
r142 18 21 18.4788 $w=2.88e-07 $l=4.65e-07 $layer=LI1_cond $X=10.705 $Y=1.75
+ $X2=10.705 $Y2=2.215
r143 16 22 2.03471 $w=4.1e-07 $l=1.5e-08 $layer=POLY_cond $X=10.645 $Y=2.23
+ $X2=10.645 $Y2=2.215
r144 16 17 38.1373 $w=4.1e-07 $l=1.5e-07 $layer=POLY_cond $X=10.63 $Y=2.23
+ $X2=10.63 $Y2=2.38
r145 13 47 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=10.705 $Y=0.58
+ $X2=10.705 $Y2=1.37
r146 9 17 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=10.5 $Y=2.75
+ $X2=10.5 $Y2=2.38
r147 2 29 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=11.44
+ $Y=2.54 $X2=11.575 $Y2=2.75
r148 1 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.57
+ $Y=0.37 $X2=11.71 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_2%A_1824_74# 1 2 9 11 13 17 18 21 23 25 26 27
+ 30 32 36 37 41 43 48 51 52 53
c137 51 0 6.53658e-20 $X=10.305 $Y=1.115
c138 41 0 1.63056e-20 $X=10.305 $Y=1.03
c139 30 0 6.19065e-20 $X=9.485 $Y=2.005
c140 26 0 6.36774e-20 $X=11.8 $Y=1.665
r141 52 53 8.67671 $w=2.98e-07 $l=1.7e-07 $layer=LI1_cond $X=11.02 $Y=1.22
+ $X2=11.19 $Y2=1.22
r142 49 56 15.7174 $w=2.76e-07 $l=9e-08 $layer=POLY_cond $X=11.725 $Y=1.26
+ $X2=11.815 $Y2=1.26
r143 48 53 20.5519 $w=2.98e-07 $l=5.35e-07 $layer=LI1_cond $X=11.725 $Y=1.26
+ $X2=11.19 $Y2=1.26
r144 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.725
+ $Y=1.26 $X2=11.725 $Y2=1.26
r145 45 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.39 $Y=1.115
+ $X2=10.305 $Y2=1.115
r146 45 52 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=10.39 $Y=1.115
+ $X2=11.02 $Y2=1.115
r147 42 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.305 $Y=1.2
+ $X2=10.305 $Y2=1.115
r148 42 43 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=10.305 $Y=1.2
+ $X2=10.305 $Y2=2.52
r149 41 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.305 $Y=1.03
+ $X2=10.305 $Y2=1.115
r150 40 41 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=10.305 $Y=0.81
+ $X2=10.305 $Y2=1.03
r151 37 39 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=9.6 $Y=2.685
+ $X2=9.885 $Y2=2.685
r152 36 43 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.22 $Y=2.685
+ $X2=10.305 $Y2=2.52
r153 36 39 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=10.22 $Y=2.685
+ $X2=9.885 $Y2=2.685
r154 32 40 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.22 $Y=0.645
+ $X2=10.305 $Y2=0.81
r155 32 34 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=10.22 $Y=0.645
+ $X2=10.1 $Y2=0.645
r156 28 37 6.87623 $w=3.3e-07 $l=2.24332e-07 $layer=LI1_cond $X=9.46 $Y=2.52
+ $X2=9.6 $Y2=2.685
r157 28 30 21.1967 $w=2.78e-07 $l=5.15e-07 $layer=LI1_cond $X=9.46 $Y=2.52
+ $X2=9.46 $Y2=2.005
r158 23 27 34.7346 $w=1.65e-07 $l=1.9e-07 $layer=POLY_cond $X=12.485 $Y=1.095
+ $X2=12.295 $Y2=1.095
r159 23 25 130.14 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=12.485 $Y=1.095
+ $X2=12.485 $Y2=0.69
r160 19 27 34.7346 $w=1.65e-07 $l=3.7229e-07 $layer=POLY_cond $X=12.385 $Y=1.425
+ $X2=12.295 $Y2=1.095
r161 19 21 402.315 $w=1.8e-07 $l=1.035e-06 $layer=POLY_cond $X=12.385 $Y=1.425
+ $X2=12.385 $Y2=2.46
r162 18 56 12.3868 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=11.89 $Y=1.26
+ $X2=11.815 $Y2=1.26
r163 17 27 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.295 $Y=1.26
+ $X2=12.295 $Y2=1.095
r164 17 18 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=12.295 $Y=1.26
+ $X2=11.89 $Y2=1.26
r165 15 56 17.0164 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.815 $Y=1.425
+ $X2=11.815 $Y2=1.26
r166 15 26 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=11.815 $Y=1.425
+ $X2=11.815 $Y2=1.665
r167 11 26 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.8 $Y=1.755
+ $X2=11.8 $Y2=1.665
r168 11 13 386.766 $w=1.8e-07 $l=9.95e-07 $layer=POLY_cond $X=11.8 $Y=1.755
+ $X2=11.8 $Y2=2.75
r169 7 49 40.1667 $w=2.76e-07 $l=3.01413e-07 $layer=POLY_cond $X=11.495 $Y=1.095
+ $X2=11.725 $Y2=1.26
r170 7 9 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=11.495 $Y=1.095
+ $X2=11.495 $Y2=0.58
r171 2 39 300 $w=1.7e-07 $l=1.09016e-06 $layer=licon1_PDIFF $count=2 $X=9.35
+ $Y=1.83 $X2=9.885 $Y2=2.685
r172 2 30 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=9.35
+ $Y=1.83 $X2=9.485 $Y2=2.005
r173 1 34 91 $w=1.7e-07 $l=1.10901e-06 $layer=licon1_NDIFF $count=2 $X=9.12
+ $Y=0.37 $X2=10.1 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_2%A_2495_392# 1 2 9 13 17 21 25 27 31 37 40
+ 41 45
r62 45 46 9.00935 $w=3.21e-07 $l=6e-08 $layer=POLY_cond $X=13.845 $Y=1.465
+ $X2=13.905 $Y2=1.465
r63 44 45 55.5576 $w=3.21e-07 $l=3.7e-07 $layer=POLY_cond $X=13.475 $Y=1.465
+ $X2=13.845 $Y2=1.465
r64 43 44 12.0125 $w=3.21e-07 $l=8e-08 $layer=POLY_cond $X=13.395 $Y=1.465
+ $X2=13.475 $Y2=1.465
r65 38 43 30.7819 $w=3.21e-07 $l=2.05e-07 $layer=POLY_cond $X=13.19 $Y=1.465
+ $X2=13.395 $Y2=1.465
r66 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.19
+ $Y=1.465 $X2=13.19 $Y2=1.465
r67 35 41 0.144206 $w=3.3e-07 $l=1.3e-07 $layer=LI1_cond $X=12.865 $Y=1.465
+ $X2=12.735 $Y2=1.465
r68 35 37 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=12.865 $Y=1.465
+ $X2=13.19 $Y2=1.465
r69 33 41 7.25953 $w=2.15e-07 $l=1.86145e-07 $layer=LI1_cond $X=12.69 $Y=1.63
+ $X2=12.735 $Y2=1.465
r70 33 40 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=12.69 $Y=1.63
+ $X2=12.69 $Y2=1.94
r71 29 41 7.25953 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=12.735 $Y=1.3
+ $X2=12.735 $Y2=1.465
r72 29 31 34.7949 $w=2.58e-07 $l=7.85e-07 $layer=LI1_cond $X=12.735 $Y=1.3
+ $X2=12.735 $Y2=0.515
r73 25 40 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.61 $Y=2.105
+ $X2=12.61 $Y2=1.94
r74 25 27 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=12.61 $Y=2.105
+ $X2=12.61 $Y2=2.815
r75 19 46 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.905 $Y=1.3
+ $X2=13.905 $Y2=1.465
r76 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.905 $Y=1.3
+ $X2=13.905 $Y2=0.74
r77 15 45 16.2883 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=13.845 $Y=1.63
+ $X2=13.845 $Y2=1.465
r78 15 17 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=13.845 $Y=1.63
+ $X2=13.845 $Y2=2.4
r79 11 44 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.475 $Y=1.3
+ $X2=13.475 $Y2=1.465
r80 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.475 $Y=1.3
+ $X2=13.475 $Y2=0.74
r81 7 43 16.2883 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=13.395 $Y=1.63
+ $X2=13.395 $Y2=1.465
r82 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=13.395 $Y=1.63
+ $X2=13.395 $Y2=2.4
r83 2 27 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=12.475
+ $Y=1.96 $X2=12.61 $Y2=2.815
r84 2 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=12.475
+ $Y=1.96 $X2=12.61 $Y2=2.105
r85 1 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.56
+ $Y=0.37 $X2=12.7 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_2%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 52 56
+ 58 63 64 66 67 69 70 71 73 78 96 100 112 116 122 131 134 137 144 148
c170 3 0 1.21651e-19 $X=4.735 $Y=1.935
r171 147 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r172 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r173 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r174 137 140 9.05853 $w=6.78e-07 $l=5.15e-07 $layer=LI1_cond $X=10.9 $Y=2.815
+ $X2=10.9 $Y2=3.33
r175 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r176 131 132 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r177 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r178 125 127 5.39368 $w=9.48e-07 $l=4.2e-07 $layer=LI1_cond $X=1.09 $Y=2.91
+ $X2=1.09 $Y2=3.33
r179 122 125 5.71474 $w=9.48e-07 $l=4.45e-07 $layer=LI1_cond $X=1.09 $Y=2.465
+ $X2=1.09 $Y2=2.91
r180 120 148 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.16 $Y2=3.33
r181 120 145 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=13.2 $Y2=3.33
r182 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r183 117 144 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.335 $Y=3.33
+ $X2=13.17 $Y2=3.33
r184 117 119 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=13.335 $Y=3.33
+ $X2=13.68 $Y2=3.33
r185 116 147 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=13.955 $Y=3.33
+ $X2=14.177 $Y2=3.33
r186 116 119 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=13.955 $Y=3.33
+ $X2=13.68 $Y2=3.33
r187 115 145 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r188 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r189 112 144 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.005 $Y=3.33
+ $X2=13.17 $Y2=3.33
r190 112 114 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=13.005 $Y=3.33
+ $X2=12.72 $Y2=3.33
r191 111 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.72 $Y2=3.33
r192 111 141 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=10.8 $Y2=3.33
r193 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r194 108 140 9.13095 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=11.24 $Y=3.33
+ $X2=10.9 $Y2=3.33
r195 108 110 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=11.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r196 107 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r197 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r198 104 107 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r199 104 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r200 103 106 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r201 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r202 101 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.58 $Y=3.33
+ $X2=8.415 $Y2=3.33
r203 101 103 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=8.58 $Y=3.33
+ $X2=8.88 $Y2=3.33
r204 100 140 9.13095 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=10.56 $Y=3.33
+ $X2=10.9 $Y2=3.33
r205 100 106 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=10.56 $Y=3.33
+ $X2=10.32 $Y2=3.33
r206 99 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r207 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r208 96 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.25 $Y=3.33
+ $X2=8.415 $Y2=3.33
r209 96 98 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.25 $Y=3.33
+ $X2=7.92 $Y2=3.33
r210 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r211 92 95 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r212 91 94 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r213 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r214 89 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r215 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r216 86 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r217 86 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r218 85 88 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r219 85 86 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r220 83 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.26 $Y2=3.33
r221 83 85 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.6 $Y2=3.33
r222 82 132 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r223 82 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r224 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r225 79 127 11.3727 $w=1.7e-07 $l=4.75e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.09 $Y2=3.33
r226 79 81 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.68 $Y2=3.33
r227 78 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=3.26 $Y2=3.33
r228 78 81 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=1.68 $Y2=3.33
r229 76 128 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r230 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r231 73 127 11.3727 $w=1.7e-07 $l=4.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=1.09 $Y2=3.33
r232 73 75 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r233 71 99 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=7.92 $Y2=3.33
r234 71 95 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=6.96 $Y2=3.33
r235 69 110 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=11.945 $Y=3.33
+ $X2=11.76 $Y2=3.33
r236 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.945 $Y=3.33
+ $X2=12.11 $Y2=3.33
r237 68 114 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=12.275 $Y=3.33
+ $X2=12.72 $Y2=3.33
r238 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.275 $Y=3.33
+ $X2=12.11 $Y2=3.33
r239 66 94 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=7.15 $Y=3.33
+ $X2=6.96 $Y2=3.33
r240 66 67 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=7.15 $Y=3.33
+ $X2=7.317 $Y2=3.33
r241 65 98 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.485 $Y=3.33
+ $X2=7.92 $Y2=3.33
r242 65 67 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=7.485 $Y=3.33
+ $X2=7.317 $Y2=3.33
r243 63 88 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.56 $Y2=3.33
r244 63 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.87 $Y2=3.33
r245 62 91 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=5.04 $Y2=3.33
r246 62 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=4.87 $Y2=3.33
r247 58 61 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=14.12 $Y=1.985
+ $X2=14.12 $Y2=2.815
r248 56 147 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=14.12 $Y=3.245
+ $X2=14.177 $Y2=3.33
r249 56 61 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=14.12 $Y=3.245
+ $X2=14.12 $Y2=2.815
r250 52 55 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=13.17 $Y=1.985
+ $X2=13.17 $Y2=2.815
r251 50 144 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.17 $Y=3.245
+ $X2=13.17 $Y2=3.33
r252 50 55 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.17 $Y=3.245
+ $X2=13.17 $Y2=2.815
r253 46 49 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=12.11 $Y=2.105
+ $X2=12.11 $Y2=2.815
r254 44 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.11 $Y=3.245
+ $X2=12.11 $Y2=3.33
r255 44 49 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=12.11 $Y=3.245
+ $X2=12.11 $Y2=2.815
r256 40 134 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.415 $Y=3.245
+ $X2=8.415 $Y2=3.33
r257 40 42 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=8.415 $Y=3.245
+ $X2=8.415 $Y2=2.535
r258 36 67 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=7.317 $Y=3.245
+ $X2=7.317 $Y2=3.33
r259 36 38 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=7.317 $Y=3.245
+ $X2=7.317 $Y2=2.825
r260 32 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=3.33
r261 32 34 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=2.88
r262 28 131 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=3.33
r263 28 30 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=2.79
r264 9 61 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=13.935
+ $Y=1.84 $X2=14.12 $Y2=2.815
r265 9 58 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=13.935
+ $Y=1.84 $X2=14.12 $Y2=1.985
r266 8 55 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=13.025
+ $Y=1.84 $X2=13.17 $Y2=2.815
r267 8 52 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=13.025
+ $Y=1.84 $X2=13.17 $Y2=1.985
r268 7 49 600 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_PDIFF $count=1 $X=11.89
+ $Y=2.54 $X2=12.11 $Y2=2.815
r269 7 46 300 $w=1.7e-07 $l=5.33784e-07 $layer=licon1_PDIFF $count=2 $X=11.89
+ $Y=2.54 $X2=12.11 $Y2=2.105
r270 6 137 300 $w=1.7e-07 $l=6.07124e-07 $layer=licon1_PDIFF $count=2 $X=10.59
+ $Y=2.54 $X2=11.075 $Y2=2.815
r271 5 42 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=8.27
+ $Y=2.34 $X2=8.415 $Y2=2.535
r272 4 38 600 $w=1.7e-07 $l=6.40625e-07 $layer=licon1_PDIFF $count=1 $X=7.095
+ $Y=2.285 $X2=7.315 $Y2=2.825
r273 3 34 600 $w=1.7e-07 $l=1.01025e-06 $layer=licon1_PDIFF $count=1 $X=4.735
+ $Y=1.935 $X2=4.87 $Y2=2.88
r274 2 30 600 $w=1.7e-07 $l=4.37321e-07 $layer=licon1_PDIFF $count=1 $X=3.125
+ $Y=2.415 $X2=3.26 $Y2=2.79
r275 1 125 300 $w=1.7e-07 $l=1.05971e-06 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=2.32 $X2=1.4 $Y2=2.91
r276 1 122 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=2.32 $X2=0.78 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_2%A_390_81# 1 2 3 4 5 18 20 24 25 27 28 29 31
+ 34 37 40 42 43 44 45 47 51
c167 51 0 8.88027e-20 $X=3.83 $Y=2.56
c168 34 0 2.36685e-20 $X=5.745 $Y=2.535
c169 29 0 1.85791e-19 $X=3.045 $Y=1.225
c170 28 0 1.8717e-19 $X=3.445 $Y=1.225
r171 49 51 0.627572 $w=4.86e-07 $l=2.5e-08 $layer=LI1_cond $X=3.72 $Y=2.535
+ $X2=3.72 $Y2=2.56
r172 48 49 2.6358 $w=4.86e-07 $l=1.05e-07 $layer=LI1_cond $X=3.72 $Y=2.43
+ $X2=3.72 $Y2=2.535
r173 46 47 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.445 $Y=1.465
+ $X2=6.445 $Y2=2.135
r174 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.36 $Y=1.38
+ $X2=6.445 $Y2=1.465
r175 44 45 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.36 $Y=1.38
+ $X2=6.115 $Y2=1.38
r176 42 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.36 $Y=2.22
+ $X2=6.445 $Y2=2.135
r177 42 43 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.36 $Y=2.22
+ $X2=5.995 $Y2=2.22
r178 38 45 7.72402 $w=1.7e-07 $l=2.01057e-07 $layer=LI1_cond $X=5.952 $Y=1.295
+ $X2=6.115 $Y2=1.38
r179 38 40 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=5.952 $Y=1.295
+ $X2=5.952 $Y2=0.815
r180 37 53 3.13516 $w=2.5e-07 $l=1.4e-07 $layer=LI1_cond $X=5.87 $Y=2.445
+ $X2=5.87 $Y2=2.585
r181 36 43 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.87 $Y=2.305
+ $X2=5.995 $Y2=2.22
r182 36 37 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=5.87 $Y=2.305
+ $X2=5.87 $Y2=2.445
r183 35 49 6.62291 $w=1.8e-07 $l=2.75e-07 $layer=LI1_cond $X=3.995 $Y=2.535
+ $X2=3.72 $Y2=2.535
r184 34 53 3.91895 $w=1.8e-07 $l=1.47902e-07 $layer=LI1_cond $X=5.745 $Y=2.535
+ $X2=5.87 $Y2=2.585
r185 34 35 107.828 $w=1.78e-07 $l=1.75e-06 $layer=LI1_cond $X=5.745 $Y=2.535
+ $X2=3.995 $Y2=2.535
r186 31 48 7.98911 $w=4.86e-07 $l=2.34734e-07 $layer=LI1_cond $X=3.53 $Y=2.33
+ $X2=3.72 $Y2=2.43
r187 30 31 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=3.53 $Y=1.31
+ $X2=3.53 $Y2=2.33
r188 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.445 $Y=1.225
+ $X2=3.53 $Y2=1.31
r189 28 29 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.445 $Y=1.225
+ $X2=3.045 $Y2=1.225
r190 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.96 $Y=1.14
+ $X2=3.045 $Y2=1.225
r191 26 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.96 $Y=0.845
+ $X2=2.96 $Y2=1.14
r192 24 48 6.97875 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=3.445 $Y=2.43
+ $X2=3.72 $Y2=2.43
r193 24 25 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.445 $Y=2.43
+ $X2=2.435 $Y2=2.43
r194 20 26 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.875 $Y=0.72
+ $X2=2.96 $Y2=0.845
r195 20 22 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=2.875 $Y=0.72
+ $X2=2.44 $Y2=0.72
r196 16 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.27 $Y=2.515
+ $X2=2.435 $Y2=2.43
r197 16 18 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=2.27 $Y=2.515
+ $X2=2.27 $Y2=2.56
r198 5 53 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=5.765
+ $Y=2.285 $X2=5.91 $Y2=2.495
r199 4 51 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=3.595
+ $Y=2.415 $X2=3.83 $Y2=2.56
r200 3 18 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=2.125
+ $Y=2.415 $X2=2.27 $Y2=2.56
r201 2 40 182 $w=1.7e-07 $l=2.89137e-07 $layer=licon1_NDIFF $count=1 $X=5.725
+ $Y=0.595 $X2=5.885 $Y2=0.815
r202 1 22 182 $w=1.7e-07 $l=6.1225e-07 $layer=licon1_NDIFF $count=1 $X=1.95
+ $Y=0.405 $X2=2.44 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_2%Q 1 2 9 13 14 15 29
r21 20 29 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=13.69 $Y=1.245
+ $X2=13.69 $Y2=1.295
r22 15 31 3.97298 $w=3.28e-07 $l=9.8e-08 $layer=LI1_cond $X=13.69 $Y=1.312
+ $X2=13.69 $Y2=1.41
r23 15 29 0.593683 $w=3.28e-07 $l=1.7e-08 $layer=LI1_cond $X=13.69 $Y=1.312
+ $X2=13.69 $Y2=1.295
r24 15 20 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=13.69 $Y=1.227
+ $X2=13.69 $Y2=1.245
r25 14 15 10.5466 $w=3.28e-07 $l=3.02e-07 $layer=LI1_cond $X=13.69 $Y=0.925
+ $X2=13.69 $Y2=1.227
r26 13 14 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=13.69 $Y=0.515
+ $X2=13.69 $Y2=0.925
r27 9 11 36.7895 $w=2.58e-07 $l=8.3e-07 $layer=LI1_cond $X=13.655 $Y=1.985
+ $X2=13.655 $Y2=2.815
r28 9 31 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=13.655 $Y=1.985
+ $X2=13.655 $Y2=1.41
r29 2 11 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=13.485
+ $Y=1.84 $X2=13.62 $Y2=2.815
r30 2 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=13.485
+ $Y=1.84 $X2=13.62 $Y2=1.985
r31 1 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.55
+ $Y=0.37 $X2=13.69 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_2%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 49
+ 51 54 55 57 58 59 61 76 83 88 93 98 104 114 117 120 124
c136 124 0 4.1906e-20 $X=14.16 $Y=0
c137 35 0 4.95374e-20 $X=4.825 $Y=0.585
r138 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r139 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r140 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r141 114 115 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r142 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r143 102 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=14.16 $Y2=0
r144 102 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r145 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r146 99 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.345 $Y=0
+ $X2=13.22 $Y2=0
r147 99 101 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=13.345 $Y=0
+ $X2=13.68 $Y2=0
r148 98 123 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=14.035 $Y=0
+ $X2=14.217 $Y2=0
r149 98 101 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=14.035 $Y=0
+ $X2=13.68 $Y2=0
r150 97 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r151 97 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r152 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r153 94 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.435 $Y=0
+ $X2=12.27 $Y2=0
r154 94 96 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=12.435 $Y=0
+ $X2=12.72 $Y2=0
r155 93 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.095 $Y=0
+ $X2=13.22 $Y2=0
r156 93 96 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.095 $Y=0
+ $X2=12.72 $Y2=0
r157 92 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r158 92 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=10.8 $Y2=0
r159 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r160 89 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.085 $Y=0
+ $X2=10.92 $Y2=0
r161 89 91 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=11.085 $Y=0
+ $X2=11.76 $Y2=0
r162 88 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.105 $Y=0
+ $X2=12.27 $Y2=0
r163 88 91 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=12.105 $Y=0
+ $X2=11.76 $Y2=0
r164 87 115 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.4 $Y=0 $X2=10.8
+ $Y2=0
r165 87 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r166 86 87 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r167 84 86 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.08 $Y=0 $X2=8.4
+ $Y2=0
r168 83 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.755 $Y=0
+ $X2=10.92 $Y2=0
r169 83 86 153.642 $w=1.68e-07 $l=2.355e-06 $layer=LI1_cond $X=10.755 $Y=0
+ $X2=8.4 $Y2=0
r170 82 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r171 81 82 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r172 78 81 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=7.44
+ $Y2=0
r173 78 79 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r174 76 111 8.18369 $w=4.73e-07 $l=3.25e-07 $layer=LI1_cond $X=7.842 $Y=0
+ $X2=7.842 $Y2=0.325
r175 76 84 6.83586 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=7.842 $Y=0 $X2=8.08
+ $Y2=0
r176 76 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r177 76 81 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.605 $Y=0
+ $X2=7.44 $Y2=0
r178 75 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r179 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r180 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r181 71 72 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r182 69 72 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r183 69 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r184 68 71 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r185 68 69 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r186 66 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0
+ $X2=0.71 $Y2=0
r187 66 68 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r188 64 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r189 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r190 61 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.71 $Y2=0
r191 61 63 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r192 59 82 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=0 $X2=7.44
+ $Y2=0
r193 59 79 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=7.2 $Y=0 $X2=5.04
+ $Y2=0
r194 57 74 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=4.56
+ $Y2=0
r195 57 58 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=4.87
+ $Y2=0
r196 56 78 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=5 $Y=0 $X2=5.04 $Y2=0
r197 56 58 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5 $Y=0 $X2=4.87
+ $Y2=0
r198 54 71 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.665 $Y=0 $X2=3.6
+ $Y2=0
r199 54 55 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.665 $Y=0 $X2=3.815
+ $Y2=0
r200 53 74 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.965 $Y=0
+ $X2=4.56 $Y2=0
r201 53 55 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.965 $Y=0 $X2=3.815
+ $Y2=0
r202 49 123 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=14.16 $Y=0.085
+ $X2=14.217 $Y2=0
r203 49 51 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=14.16 $Y=0.085
+ $X2=14.16 $Y2=0.515
r204 45 120 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.22 $Y=0.085
+ $X2=13.22 $Y2=0
r205 45 47 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=13.22 $Y=0.085
+ $X2=13.22 $Y2=0.515
r206 41 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.27 $Y=0.085
+ $X2=12.27 $Y2=0
r207 41 43 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=12.27 $Y=0.085
+ $X2=12.27 $Y2=0.515
r208 37 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.92 $Y=0.085
+ $X2=10.92 $Y2=0
r209 37 39 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.92 $Y=0.085
+ $X2=10.92 $Y2=0.58
r210 33 58 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=0.085
+ $X2=4.87 $Y2=0
r211 33 35 22.1624 $w=2.58e-07 $l=5e-07 $layer=LI1_cond $X=4.87 $Y=0.085
+ $X2=4.87 $Y2=0.585
r212 29 55 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.815 $Y=0.085
+ $X2=3.815 $Y2=0
r213 29 31 20.3598 $w=2.98e-07 $l=5.3e-07 $layer=LI1_cond $X=3.815 $Y=0.085
+ $X2=3.815 $Y2=0.615
r214 25 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r215 25 27 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.555
r216 8 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.98
+ $Y=0.37 $X2=14.12 $Y2=0.515
r217 7 47 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=13.115
+ $Y=0.37 $X2=13.26 $Y2=0.515
r218 6 43 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=12.125
+ $Y=0.37 $X2=12.27 $Y2=0.515
r219 5 39 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.78
+ $Y=0.37 $X2=10.92 $Y2=0.58
r220 4 111 182 $w=1.7e-07 $l=4.02989e-07 $layer=licon1_NDIFF $count=1 $X=7.55
+ $Y=0.595 $X2=7.84 $Y2=0.325
r221 3 35 182 $w=1.7e-07 $l=2.14942e-07 $layer=licon1_NDIFF $count=1 $X=4.615
+ $Y=0.595 $X2=4.825 $Y2=0.585
r222 2 31 182 $w=1.7e-07 $l=2.93428e-07 $layer=licon1_NDIFF $count=1 $X=3.59
+ $Y=0.405 $X2=3.79 $Y2=0.615
r223 1 27 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_2%noxref_24 1 2 7 11 13
r26 13 16 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.27 $Y=0.34
+ $X2=1.27 $Y2=0.55
r27 9 11 10.5364 $w=1.98e-07 $l=1.9e-07 $layer=LI1_cond $X=3.315 $Y=0.425
+ $X2=3.315 $Y2=0.615
r28 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.435 $Y=0.34
+ $X2=1.27 $Y2=0.34
r29 7 9 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.215 $Y=0.34
+ $X2=3.315 $Y2=0.425
r30 7 8 116.128 $w=1.68e-07 $l=1.78e-06 $layer=LI1_cond $X=3.215 $Y=0.34
+ $X2=1.435 $Y2=0.34
r31 2 11 182 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_NDIFF $count=1 $X=3.125
+ $Y=0.405 $X2=3.3 $Y2=0.615
r32 1 16 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.405 $X2=1.27 $Y2=0.55
.ends


* File: sky130_fd_sc_ms__maj3_1.pex.spice
* Created: Wed Sep  2 12:11:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__MAJ3_1%A_84_74# 1 2 3 4 15 18 20 21 24 28 31 32 33
+ 34 36 38 43 48 50 57
c115 36 0 9.62704e-20 $X=3.56 $Y=2.12
r116 50 52 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.535 $Y=1.05
+ $X2=3.535 $Y2=1.175
r117 43 58 40.6969 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.587 $Y=1.515
+ $X2=0.587 $Y2=1.68
r118 43 57 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.587 $Y=1.515
+ $X2=0.587 $Y2=1.35
r119 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.515 $X2=0.59 $Y2=1.515
r120 36 55 2.73254 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.56 $Y=2.12
+ $X2=3.56 $Y2=2.025
r121 36 38 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=3.56 $Y=2.12
+ $X2=3.56 $Y2=2.775
r122 35 48 2.76166 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=2.065 $Y=2.035
+ $X2=1.815 $Y2=2.035
r123 34 55 5.03363 $w=1.7e-07 $l=1.69926e-07 $layer=LI1_cond $X=3.395 $Y=2.035
+ $X2=3.56 $Y2=2.025
r124 34 35 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=3.395 $Y=2.035
+ $X2=2.065 $Y2=2.035
r125 33 46 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=1.175
+ $X2=1.98 $Y2=1.175
r126 32 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.37 $Y=1.175
+ $X2=3.535 $Y2=1.175
r127 32 33 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=3.37 $Y=1.175
+ $X2=2.065 $Y2=1.175
r128 31 48 3.70735 $w=2.5e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.98 $Y=1.95
+ $X2=1.815 $Y2=2.035
r129 30 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=1.26
+ $X2=1.98 $Y2=1.175
r130 30 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.98 $Y=1.26
+ $X2=1.98 $Y2=1.95
r131 26 48 3.70735 $w=2.5e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.73 $Y=2.12
+ $X2=1.815 $Y2=2.035
r132 26 28 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=1.73 $Y=2.12
+ $X2=1.73 $Y2=2.775
r133 22 46 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.645 $Y=1.175
+ $X2=1.98 $Y2=1.175
r134 22 24 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.645 $Y=1.09
+ $X2=1.645 $Y2=0.745
r135 21 42 15.029 $w=2.76e-07 $l=4.20476e-07 $layer=LI1_cond $X=0.785 $Y=1.175
+ $X2=0.605 $Y2=1.515
r136 20 22 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.48 $Y=1.175
+ $X2=1.645 $Y2=1.175
r137 20 21 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.48 $Y=1.175
+ $X2=0.785 $Y2=1.175
r138 18 58 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.55 $Y=2.4
+ $X2=0.55 $Y2=1.68
r139 15 57 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=0.87
+ $X2=0.495 $Y2=1.35
r140 4 55 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=1.92 $X2=3.56 $Y2=2.095
r141 4 38 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=1.92 $X2=3.56 $Y2=2.775
r142 3 48 400 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_PDIFF $count=1 $X=1.565
+ $Y=1.92 $X2=1.73 $Y2=2.095
r143 3 28 400 $w=1.7e-07 $l=9.33863e-07 $layer=licon1_PDIFF $count=1 $X=1.565
+ $Y=1.92 $X2=1.73 $Y2=2.775
r144 2 50 182 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_NDIFF $count=1 $X=3.395
+ $Y=0.68 $X2=3.535 $Y2=1.05
r145 1 22 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.6 $X2=1.645 $Y2=1.095
r146 1 24 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.6 $X2=1.645 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_1%B 3 7 9 11 14 16 23 25
c51 14 0 2.22981e-20 $X=1.955 $Y=2.42
r52 24 25 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.94 $Y=1.595
+ $X2=1.955 $Y2=1.595
r53 22 24 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=1.52 $Y=1.595
+ $X2=1.94 $Y2=1.595
r54 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.52
+ $Y=1.595 $X2=1.52 $Y2=1.595
r55 20 22 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=1.475 $Y=1.595
+ $X2=1.52 $Y2=1.595
r56 18 20 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=1.43 $Y=1.595
+ $X2=1.475 $Y2=1.595
r57 16 23 10.5366 $w=3.48e-07 $l=3.2e-07 $layer=LI1_cond $X=1.2 $Y=1.605
+ $X2=1.52 $Y2=1.605
r58 12 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.955 $Y=1.76
+ $X2=1.955 $Y2=1.595
r59 12 14 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.955 $Y=1.76
+ $X2=1.955 $Y2=2.42
r60 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.94 $Y=1.43
+ $X2=1.94 $Y2=1.595
r61 9 11 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.94 $Y=1.43 $X2=1.94
+ $Y2=1
r62 5 20 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.475 $Y=1.76
+ $X2=1.475 $Y2=1.595
r63 5 7 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.475 $Y=1.76
+ $X2=1.475 $Y2=2.42
r64 1 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.43 $Y=1.43
+ $X2=1.43 $Y2=1.595
r65 1 3 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.43 $Y=1.43 $X2=1.43
+ $Y2=0.92
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_1%C 3 6 10 13 17 18 20 23 25 28 34
c60 34 0 2.22981e-20 $X=2.755 $Y=1.605
c61 25 0 2.11268e-20 $X=2.435 $Y=1.4
r62 23 26 40.8642 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.435 $Y=1.595
+ $X2=2.435 $Y2=1.76
r63 23 25 51.3914 $w=3.6e-07 $l=1.95e-07 $layer=POLY_cond $X=2.435 $Y=1.595
+ $X2=2.435 $Y2=1.4
r64 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.45
+ $Y=1.595 $X2=2.45 $Y2=1.595
r65 20 34 3.83775 $w=3.48e-07 $l=1.15e-07 $layer=LI1_cond $X=2.64 $Y=1.605
+ $X2=2.755 $Y2=1.605
r66 20 24 6.25612 $w=3.48e-07 $l=1.9e-07 $layer=LI1_cond $X=2.64 $Y=1.605
+ $X2=2.45 $Y2=1.605
r67 18 29 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=1.595
+ $X2=3.41 $Y2=1.76
r68 18 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.41 $Y=1.595
+ $X2=3.41 $Y2=1.43
r69 17 34 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=3.41 $Y=1.595
+ $X2=2.755 $Y2=1.595
r70 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.41
+ $Y=1.595 $X2=3.41 $Y2=1.595
r71 13 29 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.335 $Y=2.42
+ $X2=3.335 $Y2=1.76
r72 10 28 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.32 $Y=1 $X2=3.32
+ $Y2=1.43
r73 6 26 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.375 $Y=2.42
+ $X2=2.375 $Y2=1.76
r74 3 25 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.33 $Y=1 $X2=2.33
+ $Y2=1.4
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_1%A 4 5 7 9 10 14 15 17 26 28 33
c73 33 0 2.11268e-20 $X=3.485 $Y=0.462
c74 17 0 9.62704e-20 $X=2.915 $Y=2.42
c75 4 0 5.99351e-20 $X=1.04 $Y=0.92
r76 26 33 3.89033 $w=4.13e-07 $l=1.15e-07 $layer=LI1_cond $X=3.6 $Y=0.462
+ $X2=3.485 $Y2=0.462
r77 24 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.81 $Y=0.405
+ $X2=2.81 $Y2=0.57
r78 24 28 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=2.81 $Y=0.405
+ $X2=2.81 $Y2=0.185
r79 23 33 24.6952 $w=3.13e-07 $l=6.75e-07 $layer=LI1_cond $X=2.81 $Y=0.412
+ $X2=3.485 $Y2=0.412
r80 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.81
+ $Y=0.405 $X2=2.81 $Y2=0.405
r81 15 20 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.915 $Y=1.485
+ $X2=2.915 $Y2=1.395
r82 15 17 363.444 $w=1.8e-07 $l=9.35e-07 $layer=POLY_cond $X=2.915 $Y=1.485
+ $X2=2.915 $Y2=2.42
r83 14 20 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.9 $Y=1 $X2=2.9
+ $Y2=1.395
r84 14 31 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.9 $Y=1 $X2=2.9
+ $Y2=0.57
r85 9 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=0.185
+ $X2=2.81 $Y2=0.185
r86 9 10 784.532 $w=1.5e-07 $l=1.53e-06 $layer=POLY_cond $X=2.645 $Y=0.185
+ $X2=1.115 $Y2=0.185
r87 5 19 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.055 $Y=1.405
+ $X2=1.055 $Y2=1.315
r88 5 7 394.54 $w=1.8e-07 $l=1.015e-06 $layer=POLY_cond $X=1.055 $Y=1.405
+ $X2=1.055 $Y2=2.42
r89 4 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.04 $Y=0.92
+ $X2=1.04 $Y2=1.315
r90 1 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.04 $Y=0.26
+ $X2=1.115 $Y2=0.185
r91 1 4 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.04 $Y=0.26 $X2=1.04
+ $Y2=0.92
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_1%X 1 2 9 13 14 15 16 30
c21 13 0 5.99351e-20 $X=0.265 $Y=1.18
r22 15 16 10.5285 $w=4.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.287 $Y=2.405
+ $X2=0.287 $Y2=2.775
r23 14 21 1.45122 $w=4.03e-07 $l=5.1e-08 $layer=LI1_cond $X=0.287 $Y=2.001
+ $X2=0.287 $Y2=2.052
r24 14 30 8.27043 $w=4.03e-07 $l=1.51e-07 $layer=LI1_cond $X=0.287 $Y=2.001
+ $X2=0.287 $Y2=1.85
r25 14 15 9.07727 $w=4.03e-07 $l=3.19e-07 $layer=LI1_cond $X=0.287 $Y=2.086
+ $X2=0.287 $Y2=2.405
r26 14 21 0.967483 $w=4.03e-07 $l=3.4e-08 $layer=LI1_cond $X=0.287 $Y=2.086
+ $X2=0.287 $Y2=2.052
r27 13 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.17 $Y=1.18
+ $X2=0.17 $Y2=1.85
r28 7 13 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.265 $Y=1 $X2=0.265
+ $Y2=1.18
r29 7 9 11.3644 $w=3.58e-07 $l=3.55e-07 $layer=LI1_cond $X=0.265 $Y=1 $X2=0.265
+ $Y2=0.645
r30 2 14 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.18
+ $Y=1.84 $X2=0.325 $Y2=2.015
r31 2 16 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.18
+ $Y=1.84 $X2=0.325 $Y2=2.815
r32 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.5 $X2=0.28 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_1%VPWR 1 2 11 17 19 21 31 32 35 38
r44 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 32 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r48 29 38 9.89127 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=2.84 $Y=3.33
+ $X2=2.637 $Y2=3.33
r49 29 31 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.84 $Y=3.33 $X2=3.6
+ $Y2=3.33
r50 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 25 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 24 27 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r54 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r55 22 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=3.33
+ $X2=0.825 $Y2=3.33
r56 22 24 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.99 $Y=3.33 $X2=1.2
+ $Y2=3.33
r57 21 38 9.89127 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=2.435 $Y=3.33
+ $X2=2.637 $Y2=3.33
r58 21 27 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.435 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 19 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r60 19 25 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r61 15 38 1.50354 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.637 $Y=3.245
+ $X2=2.637 $Y2=3.33
r62 15 17 24.7562 $w=4.03e-07 $l=8.7e-07 $layer=LI1_cond $X=2.637 $Y=3.245
+ $X2=2.637 $Y2=2.375
r63 11 14 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.825 $Y=2.095
+ $X2=0.825 $Y2=2.775
r64 9 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=3.245
+ $X2=0.825 $Y2=3.33
r65 9 14 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.825 $Y=3.245
+ $X2=0.825 $Y2=2.775
r66 2 17 300 $w=1.7e-07 $l=5.35397e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=1.92 $X2=2.64 $Y2=2.375
r67 1 14 400 $w=1.7e-07 $l=1.02333e-06 $layer=licon1_PDIFF $count=1 $X=0.64
+ $Y=1.84 $X2=0.825 $Y2=2.775
r68 1 11 400 $w=1.7e-07 $l=3.34963e-07 $layer=licon1_PDIFF $count=1 $X=0.64
+ $Y=1.84 $X2=0.825 $Y2=2.095
.ends

.subckt PM_SKY130_FD_SC_MS__MAJ3_1%VGND 1 2 9 12 13 15 18 19 20 22 38 39 42
r54 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r55 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r56 36 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r57 35 38 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r58 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r59 33 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r60 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r61 30 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r62 29 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r63 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r64 27 42 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.802
+ $Y2=0
r65 27 29 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.2
+ $Y2=0
r66 25 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r67 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r68 22 42 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.802
+ $Y2=0
r69 22 24 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r70 20 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r71 20 30 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r72 18 32 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.16
+ $Y2=0
r73 18 19 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.39
+ $Y2=0
r74 17 35 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.64
+ $Y2=0
r75 17 19 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.39
+ $Y2=0
r76 13 15 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.475 $Y=0.825
+ $X2=2.615 $Y2=0.825
r77 12 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.39 $Y=0.74
+ $X2=2.475 $Y2=0.825
r78 11 19 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.39 $Y=0.085
+ $X2=2.39 $Y2=0
r79 11 12 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.39 $Y=0.085
+ $X2=2.39 $Y2=0.74
r80 7 42 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.802 $Y=0.085
+ $X2=0.802 $Y2=0
r81 7 9 21.0513 $w=3.73e-07 $l=6.85e-07 $layer=LI1_cond $X=0.802 $Y=0.085
+ $X2=0.802 $Y2=0.77
r82 2 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.405
+ $Y=0.68 $X2=2.615 $Y2=0.825
r83 1 9 182 $w=1.7e-07 $l=3.67423e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.5 $X2=0.8 $Y2=0.77
.ends


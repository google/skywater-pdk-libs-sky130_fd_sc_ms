* File: sky130_fd_sc_ms__nand4b_1.pxi.spice
* Created: Fri Aug 28 17:45:07 2020
* 
x_PM_SKY130_FD_SC_MS__NAND4B_1%A_N N_A_N_M1004_g N_A_N_M1006_g A_N N_A_N_c_59_n
+ N_A_N_c_60_n PM_SKY130_FD_SC_MS__NAND4B_1%A_N
x_PM_SKY130_FD_SC_MS__NAND4B_1%D N_D_M1005_g N_D_M1008_g D N_D_c_88_n N_D_c_89_n
+ PM_SKY130_FD_SC_MS__NAND4B_1%D
x_PM_SKY130_FD_SC_MS__NAND4B_1%C N_C_M1009_g N_C_M1007_g C N_C_c_121_n
+ N_C_c_122_n PM_SKY130_FD_SC_MS__NAND4B_1%C
x_PM_SKY130_FD_SC_MS__NAND4B_1%B N_B_M1002_g N_B_M1000_g B N_B_c_154_n
+ N_B_c_155_n PM_SKY130_FD_SC_MS__NAND4B_1%B
x_PM_SKY130_FD_SC_MS__NAND4B_1%A_27_112# N_A_27_112#_M1006_s N_A_27_112#_M1004_s
+ N_A_27_112#_M1003_g N_A_27_112#_M1001_g N_A_27_112#_c_188_n
+ N_A_27_112#_c_197_n N_A_27_112#_c_189_n N_A_27_112#_c_195_n
+ N_A_27_112#_c_190_n N_A_27_112#_c_205_n N_A_27_112#_c_207_n
+ N_A_27_112#_c_191_n N_A_27_112#_c_192_n N_A_27_112#_c_193_n
+ PM_SKY130_FD_SC_MS__NAND4B_1%A_27_112#
x_PM_SKY130_FD_SC_MS__NAND4B_1%VPWR N_VPWR_M1004_d N_VPWR_M1007_d N_VPWR_M1001_d
+ N_VPWR_c_261_n N_VPWR_c_262_n N_VPWR_c_263_n N_VPWR_c_264_n N_VPWR_c_265_n
+ N_VPWR_c_266_n N_VPWR_c_267_n N_VPWR_c_268_n VPWR N_VPWR_c_269_n
+ N_VPWR_c_260_n PM_SKY130_FD_SC_MS__NAND4B_1%VPWR
x_PM_SKY130_FD_SC_MS__NAND4B_1%Y N_Y_M1003_d N_Y_M1005_d N_Y_M1000_d N_Y_c_309_n
+ N_Y_c_310_n N_Y_c_311_n N_Y_c_312_n N_Y_c_306_n N_Y_c_307_n N_Y_c_314_n
+ N_Y_c_315_n N_Y_c_308_n Y PM_SKY130_FD_SC_MS__NAND4B_1%Y
x_PM_SKY130_FD_SC_MS__NAND4B_1%VGND N_VGND_M1006_d N_VGND_c_365_n N_VGND_c_366_n
+ N_VGND_c_367_n VGND N_VGND_c_368_n N_VGND_c_369_n
+ PM_SKY130_FD_SC_MS__NAND4B_1%VGND
cc_1 VNB N_A_N_M1004_g 0.0073206f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.26
cc_2 VNB A_N 0.00846479f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_A_N_c_59_n 0.0346483f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_4 VNB N_A_N_c_60_n 0.0224562f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.22
cc_5 VNB N_D_M1005_g 0.00672475f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=2.26
cc_6 VNB D 0.00411297f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_7 VNB N_D_c_88_n 0.0318649f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_8 VNB N_D_c_89_n 0.0189071f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.22
cc_9 VNB N_C_M1007_g 0.00667073f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.835
cc_10 VNB C 0.00365302f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_11 VNB N_C_c_121_n 0.0318254f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_12 VNB N_C_c_122_n 0.0178699f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.22
cc_13 VNB N_B_M1000_g 0.00667073f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.835
cc_14 VNB B 0.00602028f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_15 VNB N_B_c_154_n 0.0297189f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_16 VNB N_B_c_155_n 0.0191804f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.22
cc_17 VNB N_A_27_112#_M1001_g 0.00688438f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_18 VNB N_A_27_112#_c_188_n 0.0140131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_112#_c_189_n 0.0011463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_112#_c_190_n 0.0298066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_112#_c_191_n 0.0055235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_112#_c_192_n 0.036431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_112#_c_193_n 0.0220447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_260_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_306_n 0.0241427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_307_n 0.028403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_308_n 0.00739565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_365_n 0.013703f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.835
cc_29 VNB N_VGND_c_366_n 0.0271358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_367_n 0.00616254f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_31 VNB N_VGND_c_368_n 0.0683234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_369_n 0.219095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VPB N_A_N_M1004_g 0.0291097f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=2.26
cc_34 VPB N_D_M1005_g 0.0246993f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=2.26
cc_35 VPB N_C_M1007_g 0.023934f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=0.835
cc_36 VPB N_B_M1000_g 0.0233443f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=0.835
cc_37 VPB N_A_27_112#_M1001_g 0.0247391f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_38 VPB N_A_27_112#_c_195_n 0.0532882f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_A_27_112#_c_190_n 0.0080854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_261_n 0.0282836f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_41 VPB N_VPWR_c_262_n 0.00900218f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_263_n 0.0156997f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_264_n 0.0476283f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_265_n 0.0249968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_266_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_267_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_268_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_269_n 0.019175f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_260_n 0.0678844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_Y_c_309_n 0.00943334f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_51 VPB N_Y_c_310_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_52 VPB N_Y_c_311_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_Y_c_312_n 0.0178895f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_Y_c_307_n 0.00301454f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_Y_c_314_n 0.00837886f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_Y_c_315_n 0.00769224f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 N_A_N_M1004_g N_D_M1005_g 0.0210097f $X=0.64 $Y=2.26 $X2=0 $Y2=0
cc_58 A_N D 0.0296943f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_59 N_A_N_c_59_n D 3.7859e-19 $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_60 A_N N_D_c_88_n 0.00187636f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_61 N_A_N_c_59_n N_D_c_88_n 0.0206382f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_62 N_A_N_c_60_n N_D_c_89_n 0.019495f $X=0.61 $Y=1.22 $X2=0 $Y2=0
cc_63 N_A_N_c_60_n N_A_27_112#_c_197_n 0.0089549f $X=0.61 $Y=1.22 $X2=0 $Y2=0
cc_64 N_A_N_M1004_g N_A_27_112#_c_195_n 0.0161412f $X=0.64 $Y=2.26 $X2=0 $Y2=0
cc_65 A_N N_A_27_112#_c_195_n 0.00793195f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_66 N_A_N_c_59_n N_A_27_112#_c_195_n 0.00231314f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_67 N_A_N_M1004_g N_A_27_112#_c_190_n 0.00840278f $X=0.64 $Y=2.26 $X2=0 $Y2=0
cc_68 A_N N_A_27_112#_c_190_n 0.0282012f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_69 N_A_N_c_59_n N_A_27_112#_c_190_n 0.00231928f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_70 N_A_N_c_60_n N_A_27_112#_c_190_n 0.00457953f $X=0.61 $Y=1.22 $X2=0 $Y2=0
cc_71 A_N N_A_27_112#_c_205_n 0.0250429f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_72 N_A_N_c_59_n N_A_27_112#_c_205_n 0.00105368f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_73 N_A_N_c_60_n N_A_27_112#_c_207_n 0.00455786f $X=0.61 $Y=1.22 $X2=0 $Y2=0
cc_74 N_A_N_M1004_g N_VPWR_c_261_n 0.00862531f $X=0.64 $Y=2.26 $X2=0 $Y2=0
cc_75 A_N N_VPWR_c_261_n 0.00187223f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_76 N_A_N_M1004_g N_VPWR_c_265_n 0.00465228f $X=0.64 $Y=2.26 $X2=0 $Y2=0
cc_77 N_A_N_M1004_g N_VPWR_c_260_n 0.00555093f $X=0.64 $Y=2.26 $X2=0 $Y2=0
cc_78 N_A_N_c_60_n N_VGND_c_365_n 0.00662399f $X=0.61 $Y=1.22 $X2=0 $Y2=0
cc_79 N_A_N_c_60_n N_VGND_c_366_n 0.00434489f $X=0.61 $Y=1.22 $X2=0 $Y2=0
cc_80 N_A_N_c_60_n N_VGND_c_369_n 0.00487769f $X=0.61 $Y=1.22 $X2=0 $Y2=0
cc_81 N_D_M1005_g N_C_M1007_g 0.023112f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_82 D C 0.0235844f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_83 N_D_c_88_n C 0.00114936f $X=1.15 $Y=1.385 $X2=0 $Y2=0
cc_84 N_D_c_89_n C 2.19577e-19 $X=1.15 $Y=1.22 $X2=0 $Y2=0
cc_85 D N_C_c_121_n 0.00114936f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_86 N_D_c_88_n N_C_c_121_n 0.0201104f $X=1.15 $Y=1.385 $X2=0 $Y2=0
cc_87 N_D_c_89_n N_C_c_122_n 0.0541207f $X=1.15 $Y=1.22 $X2=0 $Y2=0
cc_88 D N_A_27_112#_c_197_n 0.0228656f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_89 N_D_c_88_n N_A_27_112#_c_197_n 0.001011f $X=1.15 $Y=1.385 $X2=0 $Y2=0
cc_90 N_D_c_89_n N_A_27_112#_c_197_n 0.0119277f $X=1.15 $Y=1.22 $X2=0 $Y2=0
cc_91 N_D_c_89_n N_A_27_112#_c_207_n 5.7889e-19 $X=1.15 $Y=1.22 $X2=0 $Y2=0
cc_92 N_D_M1005_g N_VPWR_c_261_n 0.00446697f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_93 D N_VPWR_c_261_n 0.00773068f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_94 N_D_c_88_n N_VPWR_c_261_n 9.57671e-19 $X=1.15 $Y=1.385 $X2=0 $Y2=0
cc_95 N_D_M1005_g N_VPWR_c_267_n 0.005209f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_96 N_D_M1005_g N_VPWR_c_260_n 0.00986837f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_97 N_D_M1005_g N_Y_c_309_n 0.00512816f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_98 D N_Y_c_309_n 0.00161552f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_99 N_D_M1005_g N_Y_c_310_n 0.0105788f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_100 N_D_c_89_n N_VGND_c_365_n 0.0107451f $X=1.15 $Y=1.22 $X2=0 $Y2=0
cc_101 N_D_c_89_n N_VGND_c_368_n 0.00398535f $X=1.15 $Y=1.22 $X2=0 $Y2=0
cc_102 N_D_c_89_n N_VGND_c_369_n 0.00398847f $X=1.15 $Y=1.22 $X2=0 $Y2=0
cc_103 N_C_M1007_g N_B_M1000_g 0.0323105f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_104 C B 0.0272327f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_105 N_C_c_121_n B 0.00188716f $X=1.69 $Y=1.385 $X2=0 $Y2=0
cc_106 C N_B_c_154_n 3.99347e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_107 N_C_c_121_n N_B_c_154_n 0.0206935f $X=1.69 $Y=1.385 $X2=0 $Y2=0
cc_108 N_C_c_122_n N_B_c_155_n 0.037909f $X=1.69 $Y=1.22 $X2=0 $Y2=0
cc_109 C N_A_27_112#_c_197_n 0.0218012f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_110 N_C_c_121_n N_A_27_112#_c_197_n 8.19391e-19 $X=1.69 $Y=1.385 $X2=0 $Y2=0
cc_111 N_C_c_122_n N_A_27_112#_c_197_n 0.0119829f $X=1.69 $Y=1.22 $X2=0 $Y2=0
cc_112 N_C_M1007_g N_VPWR_c_262_n 0.00220017f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_113 N_C_M1007_g N_VPWR_c_267_n 0.005209f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_114 N_C_M1007_g N_VPWR_c_260_n 0.00982843f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_115 N_C_M1007_g N_Y_c_309_n 0.0252947f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_116 C N_Y_c_309_n 0.022292f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_117 N_C_c_121_n N_Y_c_309_n 9.3191e-19 $X=1.69 $Y=1.385 $X2=0 $Y2=0
cc_118 N_C_M1007_g N_Y_c_310_n 0.0121838f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_119 N_C_M1007_g N_Y_c_311_n 4.09773e-19 $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_120 C N_Y_c_314_n 0.00192199f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_121 N_C_c_122_n N_VGND_c_365_n 0.00212642f $X=1.69 $Y=1.22 $X2=0 $Y2=0
cc_122 N_C_c_122_n N_VGND_c_368_n 0.00461464f $X=1.69 $Y=1.22 $X2=0 $Y2=0
cc_123 N_C_c_122_n N_VGND_c_369_n 0.00465092f $X=1.69 $Y=1.22 $X2=0 $Y2=0
cc_124 N_B_M1000_g N_A_27_112#_M1001_g 0.0230827f $X=2.245 $Y=2.4 $X2=0 $Y2=0
cc_125 B N_A_27_112#_c_197_n 0.0237469f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_126 N_B_c_154_n N_A_27_112#_c_197_n 0.00100354f $X=2.23 $Y=1.385 $X2=0 $Y2=0
cc_127 N_B_c_155_n N_A_27_112#_c_197_n 0.0127995f $X=2.23 $Y=1.22 $X2=0 $Y2=0
cc_128 B N_A_27_112#_c_189_n 0.00318562f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_129 N_B_c_155_n N_A_27_112#_c_189_n 0.00162255f $X=2.23 $Y=1.22 $X2=0 $Y2=0
cc_130 B N_A_27_112#_c_191_n 0.0264357f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_131 N_B_c_154_n N_A_27_112#_c_191_n 0.00187066f $X=2.23 $Y=1.385 $X2=0 $Y2=0
cc_132 B N_A_27_112#_c_192_n 3.77186e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_133 N_B_c_154_n N_A_27_112#_c_192_n 0.02065f $X=2.23 $Y=1.385 $X2=0 $Y2=0
cc_134 N_B_c_155_n N_A_27_112#_c_193_n 0.0312011f $X=2.23 $Y=1.22 $X2=0 $Y2=0
cc_135 N_B_M1000_g N_VPWR_c_262_n 0.00722785f $X=2.245 $Y=2.4 $X2=0 $Y2=0
cc_136 N_B_M1000_g N_VPWR_c_269_n 0.0049824f $X=2.245 $Y=2.4 $X2=0 $Y2=0
cc_137 N_B_M1000_g N_VPWR_c_260_n 0.00909917f $X=2.245 $Y=2.4 $X2=0 $Y2=0
cc_138 N_B_M1000_g N_Y_c_310_n 6.58927e-19 $X=2.245 $Y=2.4 $X2=0 $Y2=0
cc_139 N_B_M1000_g N_Y_c_311_n 0.013526f $X=2.245 $Y=2.4 $X2=0 $Y2=0
cc_140 N_B_M1000_g N_Y_c_314_n 0.0198387f $X=2.245 $Y=2.4 $X2=0 $Y2=0
cc_141 B N_Y_c_314_n 0.0190624f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_142 N_B_c_154_n N_Y_c_314_n 6.72676e-19 $X=2.23 $Y=1.385 $X2=0 $Y2=0
cc_143 N_B_M1000_g N_Y_c_315_n 0.00406763f $X=2.245 $Y=2.4 $X2=0 $Y2=0
cc_144 B N_Y_c_315_n 0.00908459f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_145 N_B_c_154_n N_Y_c_315_n 4.66969e-19 $X=2.23 $Y=1.385 $X2=0 $Y2=0
cc_146 N_B_c_155_n N_VGND_c_368_n 0.00461464f $X=2.23 $Y=1.22 $X2=0 $Y2=0
cc_147 N_B_c_155_n N_VGND_c_369_n 0.00466411f $X=2.23 $Y=1.22 $X2=0 $Y2=0
cc_148 N_A_27_112#_c_195_n N_VPWR_c_261_n 0.0314063f $X=0.415 $Y=1.985 $X2=0
+ $Y2=0
cc_149 N_A_27_112#_M1001_g N_VPWR_c_264_n 0.00534567f $X=2.695 $Y=2.4 $X2=0
+ $Y2=0
cc_150 N_A_27_112#_c_195_n N_VPWR_c_265_n 0.00961163f $X=0.415 $Y=1.985 $X2=0
+ $Y2=0
cc_151 N_A_27_112#_M1001_g N_VPWR_c_269_n 0.005209f $X=2.695 $Y=2.4 $X2=0 $Y2=0
cc_152 N_A_27_112#_M1001_g N_VPWR_c_260_n 0.00985888f $X=2.695 $Y=2.4 $X2=0
+ $Y2=0
cc_153 N_A_27_112#_c_195_n N_VPWR_c_260_n 0.0143718f $X=0.415 $Y=1.985 $X2=0
+ $Y2=0
cc_154 N_A_27_112#_M1001_g N_Y_c_311_n 0.0108099f $X=2.695 $Y=2.4 $X2=0 $Y2=0
cc_155 N_A_27_112#_M1001_g N_Y_c_312_n 0.0147554f $X=2.695 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A_27_112#_c_191_n N_Y_c_312_n 0.0219515f $X=2.77 $Y=1.385 $X2=0 $Y2=0
cc_157 N_A_27_112#_c_192_n N_Y_c_312_n 0.00336308f $X=2.77 $Y=1.385 $X2=0 $Y2=0
cc_158 N_A_27_112#_c_197_n N_Y_c_306_n 0.0140856f $X=2.565 $Y=0.925 $X2=0 $Y2=0
cc_159 N_A_27_112#_c_193_n N_Y_c_306_n 0.0230379f $X=2.77 $Y=1.22 $X2=0 $Y2=0
cc_160 N_A_27_112#_M1001_g N_Y_c_307_n 0.00503397f $X=2.695 $Y=2.4 $X2=0 $Y2=0
cc_161 N_A_27_112#_c_189_n N_Y_c_307_n 0.00669252f $X=2.65 $Y=1.22 $X2=0 $Y2=0
cc_162 N_A_27_112#_c_191_n N_Y_c_307_n 0.0249903f $X=2.77 $Y=1.385 $X2=0 $Y2=0
cc_163 N_A_27_112#_c_192_n N_Y_c_307_n 0.00231223f $X=2.77 $Y=1.385 $X2=0 $Y2=0
cc_164 N_A_27_112#_c_193_n N_Y_c_307_n 0.00289106f $X=2.77 $Y=1.22 $X2=0 $Y2=0
cc_165 N_A_27_112#_M1001_g N_Y_c_315_n 0.0114614f $X=2.695 $Y=2.4 $X2=0 $Y2=0
cc_166 N_A_27_112#_c_191_n N_Y_c_315_n 0.0059332f $X=2.77 $Y=1.385 $X2=0 $Y2=0
cc_167 N_A_27_112#_c_189_n N_Y_c_308_n 0.00295346f $X=2.65 $Y=1.22 $X2=0 $Y2=0
cc_168 N_A_27_112#_c_191_n N_Y_c_308_n 0.00240045f $X=2.77 $Y=1.385 $X2=0 $Y2=0
cc_169 N_A_27_112#_c_192_n N_Y_c_308_n 6.75008e-19 $X=2.77 $Y=1.385 $X2=0 $Y2=0
cc_170 N_A_27_112#_c_197_n N_VGND_M1006_d 0.0103133f $X=2.565 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_171 N_A_27_112#_c_197_n N_VGND_c_365_n 0.0214267f $X=2.565 $Y=0.925 $X2=0
+ $Y2=0
cc_172 N_A_27_112#_c_188_n N_VGND_c_366_n 0.00300961f $X=0.275 $Y=0.845 $X2=0
+ $Y2=0
cc_173 N_A_27_112#_c_205_n N_VGND_c_366_n 0.00572092f $X=0.485 $Y=0.845 $X2=0
+ $Y2=0
cc_174 N_A_27_112#_c_193_n N_VGND_c_368_n 0.00461464f $X=2.77 $Y=1.22 $X2=0
+ $Y2=0
cc_175 N_A_27_112#_c_188_n N_VGND_c_369_n 0.00499017f $X=0.275 $Y=0.845 $X2=0
+ $Y2=0
cc_176 N_A_27_112#_c_197_n N_VGND_c_369_n 0.0577132f $X=2.565 $Y=0.925 $X2=0
+ $Y2=0
cc_177 N_A_27_112#_c_205_n N_VGND_c_369_n 0.0105838f $X=0.485 $Y=0.845 $X2=0
+ $Y2=0
cc_178 N_A_27_112#_c_193_n N_VGND_c_369_n 0.00528843f $X=2.77 $Y=1.22 $X2=0
+ $Y2=0
cc_179 N_A_27_112#_c_197_n A_263_74# 0.00734082f $X=2.565 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_180 N_A_27_112#_c_197_n A_341_74# 0.0116011f $X=2.565 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_181 N_A_27_112#_c_197_n A_443_74# 0.0127373f $X=2.565 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_182 N_VPWR_c_261_n N_Y_c_309_n 0.0146948f $X=0.95 $Y=1.985 $X2=0 $Y2=0
cc_183 N_VPWR_c_262_n N_Y_c_309_n 6.97594e-19 $X=1.95 $Y=2.405 $X2=0 $Y2=0
cc_184 N_VPWR_c_261_n N_Y_c_310_n 0.0318965f $X=0.95 $Y=1.985 $X2=0 $Y2=0
cc_185 N_VPWR_c_262_n N_Y_c_310_n 0.0255552f $X=1.95 $Y=2.405 $X2=0 $Y2=0
cc_186 N_VPWR_c_267_n N_Y_c_310_n 0.0144623f $X=1.785 $Y=3.33 $X2=0 $Y2=0
cc_187 N_VPWR_c_260_n N_Y_c_310_n 0.0118344f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_188 N_VPWR_c_262_n N_Y_c_311_n 0.0257793f $X=1.95 $Y=2.405 $X2=0 $Y2=0
cc_189 N_VPWR_c_264_n N_Y_c_311_n 0.032178f $X=2.97 $Y=2.145 $X2=0 $Y2=0
cc_190 N_VPWR_c_269_n N_Y_c_311_n 0.0152949f $X=2.805 $Y=3.33 $X2=0 $Y2=0
cc_191 N_VPWR_c_260_n N_Y_c_311_n 0.0124766f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_192 N_VPWR_M1001_d N_Y_c_312_n 0.00330044f $X=2.785 $Y=1.84 $X2=0 $Y2=0
cc_193 N_VPWR_c_264_n N_Y_c_312_n 0.0240427f $X=2.97 $Y=2.145 $X2=0 $Y2=0
cc_194 N_VPWR_M1007_d N_Y_c_314_n 0.00343351f $X=1.765 $Y=1.84 $X2=0 $Y2=0
cc_195 N_VPWR_c_262_n N_Y_c_314_n 0.0232166f $X=1.95 $Y=2.405 $X2=0 $Y2=0
cc_196 N_Y_c_306_n N_VGND_c_368_n 0.0164394f $X=2.99 $Y=0.515 $X2=0 $Y2=0
cc_197 N_Y_c_306_n N_VGND_c_369_n 0.0135988f $X=2.99 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__o221ai_1.pxi.spice
* Created: Wed Sep  2 12:23:09 2020
* 
x_PM_SKY130_FD_SC_MS__O221AI_1%C1 N_C1_M1009_g N_C1_M1002_g C1 N_C1_c_62_n
+ N_C1_c_63_n PM_SKY130_FD_SC_MS__O221AI_1%C1
x_PM_SKY130_FD_SC_MS__O221AI_1%B1 N_B1_M1004_g N_B1_M1003_g B1 N_B1_c_89_n
+ N_B1_c_90_n PM_SKY130_FD_SC_MS__O221AI_1%B1
x_PM_SKY130_FD_SC_MS__O221AI_1%B2 N_B2_M1007_g N_B2_M1001_g B2 N_B2_c_124_n
+ N_B2_c_125_n PM_SKY130_FD_SC_MS__O221AI_1%B2
x_PM_SKY130_FD_SC_MS__O221AI_1%A2 N_A2_M1005_g N_A2_M1000_g A2 A2 A2 A2
+ N_A2_c_163_n N_A2_c_164_n A2 PM_SKY130_FD_SC_MS__O221AI_1%A2
x_PM_SKY130_FD_SC_MS__O221AI_1%A1 N_A1_M1008_g N_A1_M1006_g A1 A1 N_A1_c_210_n
+ PM_SKY130_FD_SC_MS__O221AI_1%A1
x_PM_SKY130_FD_SC_MS__O221AI_1%Y N_Y_M1009_s N_Y_M1002_s N_Y_M1007_d N_Y_c_238_n
+ N_Y_c_235_n N_Y_c_256_n N_Y_c_246_n N_Y_c_262_n N_Y_c_240_n Y Y Y N_Y_c_237_n
+ PM_SKY130_FD_SC_MS__O221AI_1%Y
x_PM_SKY130_FD_SC_MS__O221AI_1%VPWR N_VPWR_M1002_d N_VPWR_M1008_d N_VPWR_c_287_n
+ N_VPWR_c_288_n N_VPWR_c_289_n N_VPWR_c_290_n VPWR N_VPWR_c_291_n
+ N_VPWR_c_292_n N_VPWR_c_286_n N_VPWR_c_294_n PM_SKY130_FD_SC_MS__O221AI_1%VPWR
x_PM_SKY130_FD_SC_MS__O221AI_1%A_114_74# N_A_114_74#_M1009_d N_A_114_74#_M1003_d
+ N_A_114_74#_c_325_n N_A_114_74#_c_326_n N_A_114_74#_c_327_n
+ PM_SKY130_FD_SC_MS__O221AI_1%A_114_74#
x_PM_SKY130_FD_SC_MS__O221AI_1%A_239_74# N_A_239_74#_M1003_s N_A_239_74#_M1001_d
+ N_A_239_74#_M1006_d N_A_239_74#_c_348_n N_A_239_74#_c_349_n
+ N_A_239_74#_c_350_n N_A_239_74#_c_351_n N_A_239_74#_c_352_n
+ N_A_239_74#_c_353_n PM_SKY130_FD_SC_MS__O221AI_1%A_239_74#
x_PM_SKY130_FD_SC_MS__O221AI_1%VGND N_VGND_M1000_d N_VGND_c_394_n VGND
+ N_VGND_c_395_n N_VGND_c_396_n N_VGND_c_397_n N_VGND_c_398_n
+ PM_SKY130_FD_SC_MS__O221AI_1%VGND
cc_1 VNB N_C1_M1009_g 0.0339542f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_C1_M1002_g 0.0015305f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.4
cc_3 VNB N_C1_c_62_n 0.00448523f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_4 VNB N_C1_c_63_n 0.0683711f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_5 VNB N_B1_M1003_g 0.0340087f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_6 VNB N_B1_c_89_n 0.0486822f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_7 VNB N_B1_c_90_n 0.0109062f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.63
cc_8 VNB N_B2_M1001_g 0.0259532f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.4
cc_9 VNB N_B2_c_124_n 0.0250975f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_10 VNB N_B2_c_125_n 0.00419897f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_11 VNB N_A2_M1000_g 0.0287203f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.4
cc_12 VNB N_A2_c_163_n 0.0269912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_c_164_n 0.00179855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A1_M1008_g 0.00172115f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_15 VNB N_A1_M1006_g 0.0335202f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.4
cc_16 VNB A1 0.0179013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_c_210_n 0.0638583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_235_n 0.0116419f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.63
cc_19 VNB Y 0.0258829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_237_n 0.00992326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_286_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_114_74#_c_325_n 0.0150295f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.4
cc_23 VNB N_A_114_74#_c_326_n 0.00814237f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_24 VNB N_A_114_74#_c_327_n 0.00262119f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_25 VNB N_A_239_74#_c_348_n 0.00920118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_239_74#_c_349_n 0.00279871f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_27 VNB N_A_239_74#_c_350_n 0.0200423f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_28 VNB N_A_239_74#_c_351_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_239_74#_c_352_n 0.00726397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_239_74#_c_353_n 0.00804404f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_394_n 0.0121692f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.4
cc_32 VNB N_VGND_c_395_n 0.0713008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_396_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_397_n 0.233314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_398_n 0.0105791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_C1_M1002_g 0.0309523f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=2.4
cc_37 VPB N_C1_c_62_n 0.0147418f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_38 VPB N_B1_M1004_g 0.0245611f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.63
cc_39 VPB N_B1_c_89_n 0.016099f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.465
cc_40 VPB N_B1_c_90_n 0.00521524f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.63
cc_41 VPB N_B2_M1007_g 0.0226492f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_42 VPB N_B2_c_124_n 0.00557395f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_43 VPB N_B2_c_125_n 0.00284954f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_44 VPB N_A2_M1005_g 0.0239605f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_45 VPB A2 0.00132234f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_46 VPB N_A2_c_163_n 0.00567265f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A1_M1008_g 0.0281988f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_48 VPB A1 0.0175673f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_Y_c_238_n 0.00262792f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_50 VPB N_Y_c_235_n 0.00180816f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.63
cc_51 VPB N_Y_c_240_n 0.00284634f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_287_n 0.0107847f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_53 VPB N_VPWR_c_288_n 0.0484149f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_54 VPB N_VPWR_c_289_n 0.0465089f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.665
cc_55 VPB N_VPWR_c_290_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_291_n 0.0239133f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_292_n 0.0131219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_286_n 0.0925773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_294_n 0.0153869f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 N_C1_c_63_n N_B1_c_89_n 0.0145415f $X=0.495 $Y=1.465 $X2=0 $Y2=0
cc_61 N_C1_M1002_g N_B1_c_90_n 6.90552e-19 $X=0.635 $Y=2.4 $X2=0 $Y2=0
cc_62 N_C1_c_63_n N_B1_c_90_n 2.28044e-19 $X=0.495 $Y=1.465 $X2=0 $Y2=0
cc_63 N_C1_M1002_g N_Y_c_238_n 0.0161124f $X=0.635 $Y=2.4 $X2=0 $Y2=0
cc_64 N_C1_M1009_g N_Y_c_235_n 0.00950615f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_65 N_C1_M1002_g N_Y_c_235_n 0.0155071f $X=0.635 $Y=2.4 $X2=0 $Y2=0
cc_66 N_C1_c_62_n N_Y_c_235_n 0.0355293f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_67 N_C1_c_63_n N_Y_c_235_n 0.00675118f $X=0.495 $Y=1.465 $X2=0 $Y2=0
cc_68 N_C1_M1002_g N_Y_c_246_n 0.0165981f $X=0.635 $Y=2.4 $X2=0 $Y2=0
cc_69 N_C1_c_62_n N_Y_c_246_n 0.00880161f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_70 N_C1_c_63_n N_Y_c_246_n 0.00361455f $X=0.495 $Y=1.465 $X2=0 $Y2=0
cc_71 N_C1_M1009_g Y 0.0146416f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_72 N_C1_M1009_g N_Y_c_237_n 0.0174061f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_73 N_C1_c_62_n N_Y_c_237_n 0.0247471f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_74 N_C1_c_63_n N_Y_c_237_n 0.00373946f $X=0.495 $Y=1.465 $X2=0 $Y2=0
cc_75 N_C1_M1002_g N_VPWR_c_287_n 0.00585939f $X=0.635 $Y=2.4 $X2=0 $Y2=0
cc_76 N_C1_M1002_g N_VPWR_c_291_n 0.005209f $X=0.635 $Y=2.4 $X2=0 $Y2=0
cc_77 N_C1_M1002_g N_VPWR_c_286_n 0.00990843f $X=0.635 $Y=2.4 $X2=0 $Y2=0
cc_78 N_C1_M1009_g N_A_114_74#_c_326_n 0.00122485f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_79 N_C1_M1009_g N_A_239_74#_c_352_n 0.00471147f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_80 N_C1_M1009_g N_VGND_c_395_n 0.00434272f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_81 N_C1_M1009_g N_VGND_c_397_n 0.00829926f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_82 N_B1_M1004_g N_B2_M1007_g 0.0459087f $X=1.545 $Y=2.4 $X2=0 $Y2=0
cc_83 N_B1_M1003_g N_B2_M1001_g 0.0313505f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_84 N_B1_c_89_n N_B2_c_124_n 0.0459087f $X=1.47 $Y=1.515 $X2=0 $Y2=0
cc_85 N_B1_c_90_n N_B2_c_124_n 0.00153564f $X=1.47 $Y=1.515 $X2=0 $Y2=0
cc_86 N_B1_c_89_n N_B2_c_125_n 0.00171497f $X=1.47 $Y=1.515 $X2=0 $Y2=0
cc_87 N_B1_c_90_n N_B2_c_125_n 0.0262024f $X=1.47 $Y=1.515 $X2=0 $Y2=0
cc_88 N_B1_M1004_g N_Y_c_235_n 0.00264604f $X=1.545 $Y=2.4 $X2=0 $Y2=0
cc_89 N_B1_c_89_n N_Y_c_235_n 0.00235174f $X=1.47 $Y=1.515 $X2=0 $Y2=0
cc_90 N_B1_c_90_n N_Y_c_235_n 0.0318707f $X=1.47 $Y=1.515 $X2=0 $Y2=0
cc_91 N_B1_M1004_g N_Y_c_256_n 0.0158091f $X=1.545 $Y=2.4 $X2=0 $Y2=0
cc_92 N_B1_c_89_n N_Y_c_256_n 0.00255564f $X=1.47 $Y=1.515 $X2=0 $Y2=0
cc_93 N_B1_c_90_n N_Y_c_256_n 0.0501791f $X=1.47 $Y=1.515 $X2=0 $Y2=0
cc_94 N_B1_M1004_g N_Y_c_240_n 0.00270272f $X=1.545 $Y=2.4 $X2=0 $Y2=0
cc_95 N_B1_M1004_g N_VPWR_c_287_n 0.0261357f $X=1.545 $Y=2.4 $X2=0 $Y2=0
cc_96 N_B1_M1004_g N_VPWR_c_289_n 0.00229331f $X=1.545 $Y=2.4 $X2=0 $Y2=0
cc_97 N_B1_M1004_g N_VPWR_c_286_n 0.00457309f $X=1.545 $Y=2.4 $X2=0 $Y2=0
cc_98 N_B1_M1003_g N_A_114_74#_c_325_n 0.0121776f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_99 N_B1_M1003_g N_A_114_74#_c_326_n 0.00672761f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_100 N_B1_M1003_g N_A_114_74#_c_327_n 4.44647e-19 $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_101 N_B1_M1003_g N_A_239_74#_c_348_n 0.00961368f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_102 N_B1_c_90_n N_A_239_74#_c_348_n 0.00947557f $X=1.47 $Y=1.515 $X2=0 $Y2=0
cc_103 N_B1_M1003_g N_A_239_74#_c_352_n 0.00723558f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_104 N_B1_c_89_n N_A_239_74#_c_352_n 0.00227386f $X=1.47 $Y=1.515 $X2=0 $Y2=0
cc_105 N_B1_c_90_n N_A_239_74#_c_352_n 0.0268812f $X=1.47 $Y=1.515 $X2=0 $Y2=0
cc_106 N_B1_M1003_g N_VGND_c_395_n 0.00291649f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_107 N_B1_M1003_g N_VGND_c_397_n 0.00364831f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_108 N_B2_M1007_g N_A2_M1005_g 0.0236726f $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_109 N_B2_M1001_g N_A2_M1000_g 0.0247498f $X=2.055 $Y=0.74 $X2=0 $Y2=0
cc_110 N_B2_M1007_g A2 8.76463e-19 $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_111 N_B2_c_125_n A2 0.00588878f $X=2.04 $Y=1.515 $X2=0 $Y2=0
cc_112 N_B2_c_124_n N_A2_c_163_n 0.0173872f $X=2.04 $Y=1.515 $X2=0 $Y2=0
cc_113 N_B2_c_125_n N_A2_c_163_n 0.0028697f $X=2.04 $Y=1.515 $X2=0 $Y2=0
cc_114 N_B2_c_124_n N_A2_c_164_n 3.65288e-19 $X=2.04 $Y=1.515 $X2=0 $Y2=0
cc_115 N_B2_c_125_n N_A2_c_164_n 0.0265213f $X=2.04 $Y=1.515 $X2=0 $Y2=0
cc_116 N_B2_M1007_g N_Y_c_256_n 0.0126379f $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_117 N_B2_c_125_n N_Y_c_256_n 0.0108932f $X=2.04 $Y=1.515 $X2=0 $Y2=0
cc_118 N_B2_M1007_g N_Y_c_262_n 8.8334e-19 $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_119 N_B2_c_124_n N_Y_c_262_n 7.75071e-19 $X=2.04 $Y=1.515 $X2=0 $Y2=0
cc_120 N_B2_c_125_n N_Y_c_262_n 0.0192914f $X=2.04 $Y=1.515 $X2=0 $Y2=0
cc_121 N_B2_M1007_g N_Y_c_240_n 0.0155906f $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_122 N_B2_M1007_g N_VPWR_c_287_n 0.00282357f $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_123 N_B2_M1007_g N_VPWR_c_289_n 0.005209f $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_124 N_B2_M1007_g N_VPWR_c_286_n 0.00984319f $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_125 N_B2_M1001_g N_A_114_74#_c_327_n 0.00617064f $X=2.055 $Y=0.74 $X2=0 $Y2=0
cc_126 N_B2_M1001_g N_A_239_74#_c_348_n 0.015042f $X=2.055 $Y=0.74 $X2=0 $Y2=0
cc_127 N_B2_c_124_n N_A_239_74#_c_348_n 0.0010384f $X=2.04 $Y=1.515 $X2=0 $Y2=0
cc_128 N_B2_c_125_n N_A_239_74#_c_348_n 0.0224475f $X=2.04 $Y=1.515 $X2=0 $Y2=0
cc_129 N_B2_M1001_g N_A_239_74#_c_349_n 0.00324276f $X=2.055 $Y=0.74 $X2=0 $Y2=0
cc_130 N_B2_M1001_g N_A_239_74#_c_352_n 6.83744e-19 $X=2.055 $Y=0.74 $X2=0 $Y2=0
cc_131 N_B2_c_124_n N_A_239_74#_c_353_n 2.37442e-19 $X=2.04 $Y=1.515 $X2=0 $Y2=0
cc_132 N_B2_c_125_n N_A_239_74#_c_353_n 0.00883898f $X=2.04 $Y=1.515 $X2=0 $Y2=0
cc_133 N_B2_M1001_g N_VGND_c_395_n 0.00434272f $X=2.055 $Y=0.74 $X2=0 $Y2=0
cc_134 N_B2_M1001_g N_VGND_c_397_n 0.00822693f $X=2.055 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A2_M1005_g N_A1_M1008_g 0.038349f $X=2.535 $Y=2.4 $X2=0 $Y2=0
cc_136 A2 N_A1_M1008_g 0.0120458f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_137 N_A2_M1000_g N_A1_M1006_g 0.0111967f $X=2.555 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A2_M1005_g A1 3.31532e-19 $X=2.535 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A2_M1000_g A1 0.00109635f $X=2.555 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A2_c_163_n A1 0.00220148f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_141 N_A2_c_164_n A1 0.0292169f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_142 N_A2_M1000_g N_A1_c_210_n 0.00138545f $X=2.555 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A2_c_163_n N_A1_c_210_n 0.0175988f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_144 N_A2_c_164_n N_A1_c_210_n 4.10694e-19 $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_145 N_A2_M1005_g N_Y_c_262_n 0.00153613f $X=2.535 $Y=2.4 $X2=0 $Y2=0
cc_146 A2 N_Y_c_262_n 0.0137715f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_147 N_A2_M1005_g N_Y_c_240_n 0.00897338f $X=2.535 $Y=2.4 $X2=0 $Y2=0
cc_148 A2 N_Y_c_240_n 0.0585275f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_149 N_A2_M1005_g N_VPWR_c_288_n 0.00173246f $X=2.535 $Y=2.4 $X2=0 $Y2=0
cc_150 A2 N_VPWR_c_288_n 0.0376957f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_151 N_A2_M1005_g N_VPWR_c_289_n 0.00449364f $X=2.535 $Y=2.4 $X2=0 $Y2=0
cc_152 A2 N_VPWR_c_289_n 0.00684978f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_153 N_A2_M1005_g N_VPWR_c_286_n 0.00737192f $X=2.535 $Y=2.4 $X2=0 $Y2=0
cc_154 A2 N_VPWR_c_286_n 0.00815361f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_155 A2 A_525_368# 0.0142598f $X=2.555 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_156 N_A2_M1000_g N_A_239_74#_c_349_n 0.013204f $X=2.555 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A2_M1000_g N_A_239_74#_c_350_n 0.0127283f $X=2.555 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A2_c_163_n N_A_239_74#_c_350_n 9.61123e-19 $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_159 N_A2_c_164_n N_A_239_74#_c_350_n 0.0171097f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_160 N_A2_M1000_g N_A_239_74#_c_353_n 0.00406658f $X=2.555 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A2_c_163_n N_A_239_74#_c_353_n 2.65889e-19 $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_162 N_A2_c_164_n N_A_239_74#_c_353_n 0.00488735f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_163 N_A2_M1000_g N_VGND_c_394_n 0.00450194f $X=2.555 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A2_M1000_g N_VGND_c_395_n 0.00434272f $X=2.555 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A2_M1000_g N_VGND_c_397_n 0.00823337f $X=2.555 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A1_M1008_g N_VPWR_c_288_n 0.0232011f $X=3.105 $Y=2.4 $X2=0 $Y2=0
cc_167 A1 N_VPWR_c_288_n 0.0264613f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_168 N_A1_c_210_n N_VPWR_c_288_n 0.00151458f $X=3.52 $Y=1.465 $X2=0 $Y2=0
cc_169 N_A1_M1008_g N_VPWR_c_289_n 0.00460063f $X=3.105 $Y=2.4 $X2=0 $Y2=0
cc_170 N_A1_M1008_g N_VPWR_c_286_n 0.00909693f $X=3.105 $Y=2.4 $X2=0 $Y2=0
cc_171 N_A1_M1006_g N_A_239_74#_c_350_n 0.0136182f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_172 A1 N_A_239_74#_c_350_n 0.0574315f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_173 N_A1_c_210_n N_A_239_74#_c_350_n 0.0125998f $X=3.52 $Y=1.465 $X2=0 $Y2=0
cc_174 N_A1_M1006_g N_A_239_74#_c_351_n 0.0138506f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A1_M1006_g N_VGND_c_394_n 0.00450194f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A1_M1006_g N_VGND_c_396_n 0.00434272f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A1_M1006_g N_VGND_c_397_n 0.00826283f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_178 N_Y_c_256_n N_VPWR_M1002_d 0.0207554f $X=2.025 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_179 N_Y_c_238_n N_VPWR_c_287_n 0.0256941f $X=0.41 $Y=2.815 $X2=0 $Y2=0
cc_180 N_Y_c_256_n N_VPWR_c_287_n 0.057997f $X=2.025 $Y=2.035 $X2=0 $Y2=0
cc_181 N_Y_c_240_n N_VPWR_c_287_n 0.0242146f $X=2.19 $Y=2.815 $X2=0 $Y2=0
cc_182 N_Y_c_240_n N_VPWR_c_289_n 0.014549f $X=2.19 $Y=2.815 $X2=0 $Y2=0
cc_183 N_Y_c_238_n N_VPWR_c_291_n 0.0109793f $X=0.41 $Y=2.815 $X2=0 $Y2=0
cc_184 N_Y_c_238_n N_VPWR_c_286_n 0.00901959f $X=0.41 $Y=2.815 $X2=0 $Y2=0
cc_185 N_Y_c_240_n N_VPWR_c_286_n 0.0119743f $X=2.19 $Y=2.815 $X2=0 $Y2=0
cc_186 N_Y_c_256_n A_327_368# 0.0096152f $X=2.025 $Y=2.035 $X2=-0.19 $Y2=-0.245
cc_187 N_Y_c_237_n N_A_114_74#_M1009_d 0.00435283f $X=0.69 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_188 Y N_A_114_74#_c_326_n 0.0165499f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_189 N_Y_c_237_n N_A_114_74#_c_326_n 0.01066f $X=0.69 $Y=1.045 $X2=0 $Y2=0
cc_190 N_Y_c_235_n N_A_239_74#_c_352_n 0.00219497f $X=0.69 $Y=1.95 $X2=0 $Y2=0
cc_191 N_Y_c_237_n N_A_239_74#_c_352_n 0.00790447f $X=0.69 $Y=1.045 $X2=0 $Y2=0
cc_192 Y N_VGND_c_395_n 0.0144497f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_193 Y N_VGND_c_397_n 0.0119539f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_194 N_A_114_74#_c_325_n N_A_239_74#_M1003_s 0.00390908f $X=1.675 $Y=0.435
+ $X2=-0.19 $Y2=-0.245
cc_195 N_A_114_74#_M1003_d N_A_239_74#_c_348_n 0.00277863f $X=1.63 $Y=0.37 $X2=0
+ $Y2=0
cc_196 N_A_114_74#_c_325_n N_A_239_74#_c_348_n 0.00357806f $X=1.675 $Y=0.435
+ $X2=0 $Y2=0
cc_197 N_A_114_74#_c_327_n N_A_239_74#_c_348_n 0.0170103f $X=1.84 $Y=0.435 $X2=0
+ $Y2=0
cc_198 N_A_114_74#_c_327_n N_A_239_74#_c_349_n 0.017488f $X=1.84 $Y=0.435 $X2=0
+ $Y2=0
cc_199 N_A_114_74#_c_325_n N_A_239_74#_c_352_n 0.013123f $X=1.675 $Y=0.435 $X2=0
+ $Y2=0
cc_200 N_A_114_74#_c_325_n N_VGND_c_395_n 0.0290838f $X=1.675 $Y=0.435 $X2=0
+ $Y2=0
cc_201 N_A_114_74#_c_326_n N_VGND_c_395_n 0.0141382f $X=0.78 $Y=0.435 $X2=0
+ $Y2=0
cc_202 N_A_114_74#_c_327_n N_VGND_c_395_n 0.0141284f $X=1.84 $Y=0.435 $X2=0
+ $Y2=0
cc_203 N_A_114_74#_c_325_n N_VGND_c_397_n 0.0250986f $X=1.675 $Y=0.435 $X2=0
+ $Y2=0
cc_204 N_A_114_74#_c_326_n N_VGND_c_397_n 0.0119234f $X=0.78 $Y=0.435 $X2=0
+ $Y2=0
cc_205 N_A_114_74#_c_327_n N_VGND_c_397_n 0.0118299f $X=1.84 $Y=0.435 $X2=0
+ $Y2=0
cc_206 N_A_239_74#_c_350_n N_VGND_M1000_d 0.0079007f $X=3.395 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_207 N_A_239_74#_c_349_n N_VGND_c_394_n 0.0173638f $X=2.34 $Y=0.515 $X2=0
+ $Y2=0
cc_208 N_A_239_74#_c_350_n N_VGND_c_394_n 0.0427946f $X=3.395 $Y=1.045 $X2=0
+ $Y2=0
cc_209 N_A_239_74#_c_351_n N_VGND_c_394_n 0.0173638f $X=3.56 $Y=0.515 $X2=0
+ $Y2=0
cc_210 N_A_239_74#_c_349_n N_VGND_c_395_n 0.0145639f $X=2.34 $Y=0.515 $X2=0
+ $Y2=0
cc_211 N_A_239_74#_c_351_n N_VGND_c_396_n 0.0145639f $X=3.56 $Y=0.515 $X2=0
+ $Y2=0
cc_212 N_A_239_74#_c_349_n N_VGND_c_397_n 0.0119984f $X=2.34 $Y=0.515 $X2=0
+ $Y2=0
cc_213 N_A_239_74#_c_351_n N_VGND_c_397_n 0.0119984f $X=3.56 $Y=0.515 $X2=0
+ $Y2=0

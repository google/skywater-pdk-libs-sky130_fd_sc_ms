* File: sky130_fd_sc_ms__dfrtp_1.pex.spice
* Created: Wed Sep  2 12:03:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DFRTP_1%D 2 5 9 11 12 13 18 19 22
r32 22 24 40.9207 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.845
+ $X2=0.402 $Y2=2.01
r33 22 23 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.845 $X2=0.385 $Y2=1.845
r34 18 20 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.165
+ $X2=0.402 $Y2=1
r35 18 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.165 $X2=0.385 $Y2=1.165
r36 13 23 5.61447 $w=3.88e-07 $l=1.9e-07 $layer=LI1_cond $X=0.32 $Y=2.035
+ $X2=0.32 $Y2=1.845
r37 12 23 5.31897 $w=3.88e-07 $l=1.8e-07 $layer=LI1_cond $X=0.32 $Y=1.665
+ $X2=0.32 $Y2=1.845
r38 11 12 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.32 $Y=1.295
+ $X2=0.32 $Y2=1.665
r39 11 19 3.84148 $w=3.88e-07 $l=1.3e-07 $layer=LI1_cond $X=0.32 $Y=1.295
+ $X2=0.32 $Y2=1.165
r40 9 20 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.51 $Y=0.6 $X2=0.51
+ $Y2=1
r41 5 24 316.798 $w=1.8e-07 $l=8.15e-07 $layer=POLY_cond $X=0.495 $Y=2.825
+ $X2=0.495 $Y2=2.01
r42 2 22 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=0.402 $Y=1.828
+ $X2=0.402 $Y2=1.845
r43 1 18 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=0.402 $Y=1.182
+ $X2=0.402 $Y2=1.165
r44 1 2 102.129 $w=3.65e-07 $l=6.46e-07 $layer=POLY_cond $X=0.402 $Y=1.182
+ $X2=0.402 $Y2=1.828
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_1%CLK 3 7 8 11 13
c45 8 0 1.4256e-19 $X=2.16 $Y=1.665
c46 3 0 1.46527e-19 $X=1.925 $Y=2.495
r47 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.91 $Y=1.61
+ $X2=1.91 $Y2=1.775
r48 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.91 $Y=1.61
+ $X2=1.91 $Y2=1.445
r49 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.91
+ $Y=1.61 $X2=1.91 $Y2=1.61
r50 8 12 6.53105 $w=4.67e-07 $l=2.5e-07 $layer=LI1_cond $X=2.16 $Y=1.545
+ $X2=1.91 $Y2=1.545
r51 7 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.955 $Y=0.965
+ $X2=1.955 $Y2=1.445
r52 3 14 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.925 $Y=2.495
+ $X2=1.925 $Y2=1.775
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_1%A_493_387# 1 2 9 11 13 15 17 19 20 21 24 28
+ 29 32 33 34 36 37 38 41 45 48 52 59 62 64 74
c193 64 0 1.8423e-19 $X=3.337 $Y=1.76
c194 48 0 1.4256e-19 $X=2.945 $Y=1.925
c195 38 0 1.54738e-19 $X=5.65 $Y=0.34
c196 21 0 1.90132e-19 $X=6.33 $Y=1.27
c197 13 0 2.46211e-20 $X=4.03 $Y=1.435
c198 9 0 8.14778e-21 $X=3.415 $Y=2.525
r199 61 62 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=7.13 $Y=1.18
+ $X2=7.335 $Y2=1.18
r200 59 70 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.855 $Y=1.18
+ $X2=6.855 $Y2=1.27
r201 58 61 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.855 $Y=1.18
+ $X2=7.13 $Y2=1.18
r202 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.855
+ $Y=1.18 $X2=6.855 $Y2=1.18
r203 55 56 7.05682 $w=4.83e-07 $l=8.5e-08 $layer=LI1_cond $X=2.792 $Y=0.72
+ $X2=2.792 $Y2=0.805
r204 52 55 9.37134 $w=4.83e-07 $l=3.8e-07 $layer=LI1_cond $X=2.792 $Y=0.34
+ $X2=2.792 $Y2=0.72
r205 51 67 40.6969 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=3.337 $Y=1.85
+ $X2=3.337 $Y2=2.015
r206 51 64 15.5026 $w=3.35e-07 $l=9e-08 $layer=POLY_cond $X=3.337 $Y=1.85
+ $X2=3.337 $Y2=1.76
r207 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.335
+ $Y=1.85 $X2=3.335 $Y2=1.85
r208 48 50 10.9885 $w=4.33e-07 $l=3.9e-07 $layer=LI1_cond $X=2.945 $Y=1.925
+ $X2=3.335 $Y2=1.925
r209 47 48 9.72055 $w=4.33e-07 $l=4.2761e-07 $layer=LI1_cond $X=2.6 $Y=2.11
+ $X2=2.945 $Y2=1.925
r210 45 62 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.335 $Y=1.015
+ $X2=7.335 $Y2=1.18
r211 44 45 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.335 $Y=0.425
+ $X2=7.335 $Y2=1.015
r212 42 74 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=7.13 $Y=2.14
+ $X2=7.265 $Y2=2.14
r213 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.13
+ $Y=2.14 $X2=7.13 $Y2=2.14
r214 39 61 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.13 $Y=1.345
+ $X2=7.13 $Y2=1.18
r215 39 41 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=7.13 $Y=1.345
+ $X2=7.13 $Y2=2.14
r216 37 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.25 $Y=0.34
+ $X2=7.335 $Y2=0.425
r217 37 38 104.385 $w=1.68e-07 $l=1.6e-06 $layer=LI1_cond $X=7.25 $Y=0.34
+ $X2=5.65 $Y2=0.34
r218 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.565 $Y=0.425
+ $X2=5.65 $Y2=0.34
r219 35 36 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.565 $Y=0.425
+ $X2=5.565 $Y2=0.565
r220 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.48 $Y=0.65
+ $X2=5.565 $Y2=0.565
r221 33 34 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=5.48 $Y=0.65 $X2=4.48
+ $Y2=0.65
r222 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.395 $Y=0.565
+ $X2=4.48 $Y2=0.65
r223 31 32 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=4.395 $Y=0.425
+ $X2=4.395 $Y2=0.565
r224 30 52 6.96588 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=3.035 $Y=0.34
+ $X2=2.792 $Y2=0.34
r225 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.31 $Y=0.34
+ $X2=4.395 $Y2=0.425
r226 29 30 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=4.31 $Y=0.34
+ $X2=3.035 $Y2=0.34
r227 28 48 5.91304 $w=1.8e-07 $l=3.5e-07 $layer=LI1_cond $X=2.945 $Y=1.575
+ $X2=2.945 $Y2=1.925
r228 28 56 47.4444 $w=1.78e-07 $l=7.7e-07 $layer=LI1_cond $X=2.945 $Y=1.575
+ $X2=2.945 $Y2=0.805
r229 22 74 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.265 $Y=2.305
+ $X2=7.265 $Y2=2.14
r230 22 24 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=7.265 $Y=2.305
+ $X2=7.265 $Y2=2.675
r231 20 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.69 $Y=1.27
+ $X2=6.855 $Y2=1.27
r232 20 21 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=6.69 $Y=1.27
+ $X2=6.33 $Y2=1.27
r233 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.255 $Y=1.195
+ $X2=6.33 $Y2=1.27
r234 17 19 146.207 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=6.255 $Y=1.195
+ $X2=6.255 $Y2=0.74
r235 13 26 82.6988 $w=1.96e-07 $l=3.55106e-07 $layer=POLY_cond $X=4.03 $Y=1.435
+ $X2=3.967 $Y2=1.76
r236 13 15 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=4.03 $Y=1.435
+ $X2=4.03 $Y2=0.9
r237 12 64 21.5811 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=3.505 $Y=1.76
+ $X2=3.337 $Y2=1.76
r238 11 26 9.11062 $w=1.5e-07 $l=1.37e-07 $layer=POLY_cond $X=3.83 $Y=1.76
+ $X2=3.967 $Y2=1.76
r239 11 12 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=3.83 $Y=1.76
+ $X2=3.505 $Y2=1.76
r240 9 67 198.242 $w=1.8e-07 $l=5.1e-07 $layer=POLY_cond $X=3.415 $Y=2.525
+ $X2=3.415 $Y2=2.015
r241 2 47 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.935 $X2=2.6 $Y2=2.11
r242 1 55 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=2.55
+ $Y=0.595 $X2=2.715 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_1%A_833_400# 1 2 7 9 13 17 20 21 26 29 33
c88 21 0 5.33388e-20 $X=4.445 $Y=0.99
c89 20 0 1.06493e-20 $X=5.82 $Y=0.99
c90 9 0 1.36594e-19 $X=4.255 $Y=2.525
r91 32 33 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=6.065 $Y=1.13
+ $X2=6.065 $Y2=1.865
r92 31 32 7.58911 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=5.985 $Y=0.99
+ $X2=5.985 $Y2=1.13
r93 29 31 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=5.985 $Y=0.855
+ $X2=5.985 $Y2=0.99
r94 26 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.145 $Y=2.03
+ $X2=6.145 $Y2=1.865
r95 20 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.82 $Y=0.99
+ $X2=5.985 $Y2=0.99
r96 20 21 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=5.82 $Y=0.99
+ $X2=4.445 $Y2=0.99
r97 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.36
+ $Y=1.96 $X2=4.36 $Y2=1.96
r98 15 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.36 $Y=1.075
+ $X2=4.445 $Y2=0.99
r99 15 17 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=4.36 $Y=1.075
+ $X2=4.36 $Y2=1.96
r100 11 18 38.6889 $w=3.41e-07 $l=1.88348e-07 $layer=POLY_cond $X=4.395 $Y=1.795
+ $X2=4.345 $Y2=1.96
r101 11 13 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=4.395 $Y=1.795
+ $X2=4.395 $Y2=0.9
r102 7 18 34.0112 $w=3.41e-07 $l=2.05122e-07 $layer=POLY_cond $X=4.255 $Y=2.125
+ $X2=4.345 $Y2=1.96
r103 7 9 155.484 $w=1.8e-07 $l=4e-07 $layer=POLY_cond $X=4.255 $Y=2.125
+ $X2=4.255 $Y2=2.525
r104 2 26 300 $w=1.7e-07 $l=3.72357e-07 $layer=licon1_PDIFF $count=2 $X=5.97
+ $Y=1.735 $X2=6.145 $Y2=2.03
r105 1 29 182 $w=1.7e-07 $l=6.8057e-07 $layer=licon1_NDIFF $count=1 $X=5.515
+ $Y=0.37 $X2=5.985 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_1%RESET_B 4 6 9 11 12 16 17 19 21 24 28 32 34
+ 35 36 37 40 42 45 48 49 52 59 60
c214 49 0 1.33156e-19 $X=1.155 $Y=1.295
c215 48 0 1.17243e-19 $X=1.155 $Y=1.295
c216 36 0 4.55276e-20 $X=7.775 $Y=2.035
c217 35 0 1.33709e-20 $X=1.345 $Y=2.035
c218 34 0 2.46211e-20 $X=4.895 $Y=2.035
c219 16 0 1.54738e-19 $X=4.785 $Y=0.9
c220 11 0 6.39881e-20 $X=4.71 $Y=0.18
r221 59 62 40.6969 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=8.182 $Y=2.09
+ $X2=8.182 $Y2=2.255
r222 59 61 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=8.182 $Y=2.09
+ $X2=8.182 $Y2=1.925
r223 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.18
+ $Y=2.09 $X2=8.18 $Y2=2.09
r224 52 54 40.6549 $w=4.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.072 $Y=1.975
+ $X2=1.072 $Y2=2.14
r225 52 53 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.975 $X2=1.155 $Y2=1.975
r226 49 53 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.155 $Y=1.295
+ $X2=1.155 $Y2=1.975
r227 48 50 46.3954 $w=4.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.072 $Y=1.295
+ $X2=1.072 $Y2=1.13
r228 48 49 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.295 $X2=1.155 $Y2=1.295
r229 45 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.035
+ $X2=1.2 $Y2=2.035
r230 43 60 8.94433 $w=3.33e-07 $l=2.6e-07 $layer=LI1_cond $X=7.92 $Y=2.087
+ $X2=8.18 $Y2=2.087
r231 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r232 40 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.12
+ $Y=1.96 $X2=5.12 $Y2=1.96
r233 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=2.035
+ $X2=5.04 $Y2=2.035
r234 37 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=2.035
+ $X2=5.04 $Y2=2.035
r235 36 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r236 36 37 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=5.185 $Y2=2.035
r237 35 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=2.035
+ $X2=1.2 $Y2=2.035
r238 34 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=5.04 $Y2=2.035
r239 34 35 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=1.345 $Y2=2.035
r240 30 32 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.785 $Y=1.26
+ $X2=4.875 $Y2=1.26
r241 28 62 163.258 $w=1.8e-07 $l=4.2e-07 $layer=POLY_cond $X=8.26 $Y=2.675
+ $X2=8.26 $Y2=2.255
r242 24 61 671.723 $w=1.5e-07 $l=1.31e-06 $layer=POLY_cond $X=8.205 $Y=0.615
+ $X2=8.205 $Y2=1.925
r243 21 56 39.7049 $w=4.06e-07 $l=2.28703e-07 $layer=POLY_cond $X=4.875 $Y=1.795
+ $X2=5.027 $Y2=1.96
r244 20 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.875 $Y=1.335
+ $X2=4.875 $Y2=1.26
r245 20 21 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=4.875 $Y=1.335
+ $X2=4.875 $Y2=1.795
r246 17 56 52.5546 $w=4.06e-07 $l=3.89654e-07 $layer=POLY_cond $X=4.86 $Y=2.275
+ $X2=5.027 $Y2=1.96
r247 17 19 66.9444 $w=1.8e-07 $l=2.5e-07 $layer=POLY_cond $X=4.86 $Y=2.275
+ $X2=4.86 $Y2=2.525
r248 14 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.785 $Y=1.185
+ $X2=4.785 $Y2=1.26
r249 14 16 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.785 $Y=1.185
+ $X2=4.785 $Y2=0.9
r250 13 16 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=4.785 $Y=0.255
+ $X2=4.785 $Y2=0.9
r251 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.71 $Y=0.18
+ $X2=4.785 $Y2=0.255
r252 11 12 1915.18 $w=1.5e-07 $l=3.735e-06 $layer=POLY_cond $X=4.71 $Y=0.18
+ $X2=0.975 $Y2=0.18
r253 9 54 266.266 $w=1.8e-07 $l=6.85e-07 $layer=POLY_cond $X=0.945 $Y=2.825
+ $X2=0.945 $Y2=2.14
r254 6 52 8.86311 $w=4.95e-07 $l=8.2e-08 $layer=POLY_cond $X=1.072 $Y=1.893
+ $X2=1.072 $Y2=1.975
r255 5 48 8.86311 $w=4.95e-07 $l=8.2e-08 $layer=POLY_cond $X=1.072 $Y=1.377
+ $X2=1.072 $Y2=1.295
r256 5 6 55.7728 $w=4.95e-07 $l=5.16e-07 $layer=POLY_cond $X=1.072 $Y=1.377
+ $X2=1.072 $Y2=1.893
r257 4 50 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.9 $Y=0.6 $X2=0.9
+ $Y2=1.13
r258 1 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.9 $Y=0.255
+ $X2=0.975 $Y2=0.18
r259 1 4 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=0.9 $Y=0.255 $X2=0.9
+ $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_1%A_701_463# 1 2 3 12 16 18 24 27 29 30 32 33
+ 38 40 41 44 47
c130 41 0 1.83166e-19 $X=4.075 $Y=2.36
c131 40 0 8.14778e-21 $X=4.075 $Y=2.46
c132 24 0 1.06777e-19 $X=4.615 $Y=2.46
c133 18 0 2.25353e-19 $X=3.935 $Y=2.64
r134 44 46 15.8682 $w=2.96e-07 $l=3.85e-07 $layer=LI1_cond $X=4.7 $Y=2.5
+ $X2=5.085 $Y2=2.5
r135 40 42 7.40856 $w=2.78e-07 $l=1.8e-07 $layer=LI1_cond $X=4.075 $Y=2.46
+ $X2=4.075 $Y2=2.64
r136 40 41 5.88157 $w=2.78e-07 $l=1e-07 $layer=LI1_cond $X=4.075 $Y=2.46
+ $X2=4.075 $Y2=2.36
r137 36 38 6.09338 $w=4.33e-07 $l=2.3e-07 $layer=LI1_cond $X=3.79 $Y=0.812
+ $X2=4.02 $Y2=0.812
r138 33 48 9 $w=2.41e-07 $l=4.5e-08 $layer=POLY_cond $X=5.485 $Y=1.41 $X2=5.44
+ $Y2=1.41
r139 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.485
+ $Y=1.41 $X2=5.485 $Y2=1.41
r140 30 47 7.71909 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=5.335 $Y=1.43
+ $X2=5.19 $Y2=1.43
r141 30 32 5.96091 $w=2.88e-07 $l=1.5e-07 $layer=LI1_cond $X=5.335 $Y=1.43
+ $X2=5.485 $Y2=1.43
r142 29 47 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.785 $Y=1.49
+ $X2=5.19 $Y2=1.49
r143 27 44 3.98214 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=4.7 $Y=2.32 $X2=4.7
+ $Y2=2.5
r144 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.7 $Y=1.575
+ $X2=4.785 $Y2=1.49
r145 26 27 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=4.7 $Y=1.575
+ $X2=4.7 $Y2=2.32
r146 25 40 2.70854 $w=2e-07 $l=1.4e-07 $layer=LI1_cond $X=4.215 $Y=2.46
+ $X2=4.075 $Y2=2.46
r147 24 44 4.79272 $w=2.96e-07 $l=1.03078e-07 $layer=LI1_cond $X=4.615 $Y=2.46
+ $X2=4.7 $Y2=2.5
r148 24 25 22.1818 $w=1.98e-07 $l=4e-07 $layer=LI1_cond $X=4.615 $Y=2.46
+ $X2=4.215 $Y2=2.46
r149 22 38 6.29128 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=4.02 $Y=1.03
+ $X2=4.02 $Y2=0.812
r150 22 41 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=4.02 $Y=1.03
+ $X2=4.02 $Y2=2.36
r151 18 42 1.89134 $w=2.3e-07 $l=1.4e-07 $layer=LI1_cond $X=3.935 $Y=2.64
+ $X2=4.075 $Y2=2.64
r152 18 20 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.935 $Y=2.64
+ $X2=3.64 $Y2=2.64
r153 14 33 79 $w=2.41e-07 $l=4.70319e-07 $layer=POLY_cond $X=5.88 $Y=1.575
+ $X2=5.485 $Y2=1.41
r154 14 16 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=5.88 $Y=1.575
+ $X2=5.88 $Y2=2.235
r155 10 48 13.8727 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.44 $Y=1.245
+ $X2=5.44 $Y2=1.41
r156 10 12 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.44 $Y=1.245
+ $X2=5.44 $Y2=0.74
r157 3 46 600 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=4.95
+ $Y=2.315 $X2=5.085 $Y2=2.485
r158 2 20 600 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_PDIFF $count=1 $X=3.505
+ $Y=2.315 $X2=3.64 $Y2=2.61
r159 1 36 182 $w=1.7e-07 $l=2.40416e-07 $layer=licon1_NDIFF $count=1 $X=3.62
+ $Y=0.69 $X2=3.79 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_1%A_299_387# 1 2 9 11 13 15 16 17 18 19 22 26
+ 28 33 34 35 38 40 43 46 47 50 52 56
c177 52 0 1.17243e-19 $X=1.695 $Y=1.055
c178 50 0 4.54223e-20 $X=2.565 $Y=1.43
c179 26 0 1.06777e-19 $X=3.865 $Y=2.525
c180 18 0 1.83166e-19 $X=3.47 $Y=1.4
c181 15 0 8.87588e-20 $X=2.885 $Y=3.075
r182 60 64 38.1583 $w=3.6e-07 $l=2.85e-07 $layer=POLY_cond $X=2.6 $Y=1.55
+ $X2=2.885 $Y2=1.55
r183 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.6
+ $Y=1.61 $X2=2.6 $Y2=1.61
r184 53 56 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=1.54 $Y=2.11 $X2=1.62
+ $Y2=2.11
r185 50 59 9.63385 $w=2.4e-07 $l=1.8e-07 $layer=LI1_cond $X=2.565 $Y=1.43
+ $X2=2.565 $Y2=1.61
r186 49 50 13.9254 $w=2.38e-07 $l=2.9e-07 $layer=LI1_cond $X=2.565 $Y=1.14
+ $X2=2.565 $Y2=1.43
r187 48 52 3.35233 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=1.87 $Y=1.055
+ $X2=1.662 $Y2=1.055
r188 47 49 10.2245 $w=1.41e-07 $l=1.56844e-07 $layer=LI1_cond $X=2.445 $Y=1.055
+ $X2=2.565 $Y2=1.14
r189 47 48 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.445 $Y=1.055
+ $X2=1.87 $Y2=1.055
r190 46 53 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=1.945
+ $X2=1.54 $Y2=2.11
r191 45 52 3.22182 $w=2.92e-07 $l=1.58915e-07 $layer=LI1_cond $X=1.54 $Y=1.14
+ $X2=1.662 $Y2=1.055
r192 45 46 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.54 $Y=1.14
+ $X2=1.54 $Y2=1.945
r193 41 52 3.22182 $w=2.92e-07 $l=8.5e-08 $layer=LI1_cond $X=1.662 $Y=0.97
+ $X2=1.662 $Y2=1.055
r194 41 43 7.08128 $w=4.13e-07 $l=2.55e-07 $layer=LI1_cond $X=1.662 $Y=0.97
+ $X2=1.662 $Y2=0.715
r195 36 38 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=7.305 $Y=1.585
+ $X2=7.305 $Y2=0.615
r196 34 36 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.23 $Y=1.66
+ $X2=7.305 $Y2=1.585
r197 34 35 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=7.23 $Y=1.66
+ $X2=6.475 $Y2=1.66
r198 31 33 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=6.385 $Y=3.075
+ $X2=6.385 $Y2=2.385
r199 30 35 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.385 $Y=1.735
+ $X2=6.475 $Y2=1.66
r200 30 33 252.661 $w=1.8e-07 $l=6.5e-07 $layer=POLY_cond $X=6.385 $Y=1.735
+ $X2=6.385 $Y2=2.385
r201 29 40 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.955 $Y=3.15
+ $X2=3.865 $Y2=3.15
r202 28 31 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.295 $Y=3.15
+ $X2=6.385 $Y2=3.075
r203 28 29 1199.87 $w=1.5e-07 $l=2.34e-06 $layer=POLY_cond $X=6.295 $Y=3.15
+ $X2=3.955 $Y2=3.15
r204 24 40 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.865 $Y=3.075
+ $X2=3.865 $Y2=3.15
r205 24 26 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=3.865 $Y=3.075
+ $X2=3.865 $Y2=2.525
r206 20 22 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=3.545 $Y=1.325
+ $X2=3.545 $Y2=0.9
r207 19 64 37.5714 $w=3.6e-07 $l=2.17428e-07 $layer=POLY_cond $X=3.04 $Y=1.4
+ $X2=2.885 $Y2=1.55
r208 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.47 $Y=1.4
+ $X2=3.545 $Y2=1.325
r209 18 19 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.47 $Y=1.4
+ $X2=3.04 $Y2=1.4
r210 16 40 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.775 $Y=3.15
+ $X2=3.865 $Y2=3.15
r211 16 17 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=3.775 $Y=3.15
+ $X2=2.96 $Y2=3.15
r212 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.885 $Y=3.075
+ $X2=2.96 $Y2=3.15
r213 14 64 23.3057 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.885 $Y=1.775
+ $X2=2.885 $Y2=1.55
r214 14 15 666.596 $w=1.5e-07 $l=1.3e-06 $layer=POLY_cond $X=2.885 $Y=1.775
+ $X2=2.885 $Y2=3.075
r215 11 60 16.7361 $w=3.6e-07 $l=1.25e-07 $layer=POLY_cond $X=2.475 $Y=1.55
+ $X2=2.6 $Y2=1.55
r216 11 61 13.3889 $w=3.6e-07 $l=1e-07 $layer=POLY_cond $X=2.475 $Y=1.55
+ $X2=2.375 $Y2=1.55
r217 11 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.475 $Y=1.41
+ $X2=2.475 $Y2=0.965
r218 7 61 18.9685 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=2.375 $Y=1.775
+ $X2=2.375 $Y2=1.55
r219 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.375 $Y=1.775
+ $X2=2.375 $Y2=2.495
r220 2 56 600 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.935 $X2=1.62 $Y2=2.1
r221 1 52 182 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_NDIFF $count=1 $X=1.55
+ $Y=0.59 $X2=1.695 $Y2=1.055
r222 1 43 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.55
+ $Y=0.59 $X2=1.695 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_1%A_1518_203# 1 2 9 11 15 17 18 24 26 27 29 30
+ 34 37 38 41
r114 37 38 10.5766 $w=3.63e-07 $l=2.3e-07 $layer=LI1_cond $X=8.502 $Y=2.675
+ $X2=8.502 $Y2=2.445
r115 34 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.755 $Y=1.18
+ $X2=7.755 $Y2=1.345
r116 34 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.755 $Y=1.18
+ $X2=7.755 $Y2=1.015
r117 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.755
+ $Y=1.18 $X2=7.755 $Y2=1.18
r118 30 33 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.755 $Y=1.1 $X2=7.755
+ $Y2=1.18
r119 28 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.105 $Y=1.185
+ $X2=9.105 $Y2=1.1
r120 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.105 $Y=1.185
+ $X2=9.105 $Y2=1.855
r121 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.02 $Y=1.94
+ $X2=9.105 $Y2=1.855
r122 26 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.02 $Y=1.94
+ $X2=8.685 $Y2=1.94
r123 22 41 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.78 $Y=1.1
+ $X2=9.105 $Y2=1.1
r124 22 24 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=8.78 $Y=1.015 $X2=8.78
+ $Y2=0.615
r125 20 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.6 $Y=2.025
+ $X2=8.685 $Y2=1.94
r126 20 38 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=8.6 $Y=2.025
+ $X2=8.6 $Y2=2.445
r127 19 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.92 $Y=1.1
+ $X2=7.755 $Y2=1.1
r128 18 22 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=8.615 $Y=1.1
+ $X2=8.78 $Y2=1.1
r129 18 19 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=8.615 $Y=1.1
+ $X2=7.92 $Y2=1.1
r130 17 45 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=7.67 $Y=1.745
+ $X2=7.67 $Y2=1.345
r131 15 44 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=7.695 $Y=0.615
+ $X2=7.695 $Y2=1.015
r132 9 17 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.685 $Y=1.835
+ $X2=7.685 $Y2=1.745
r133 9 11 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=7.685 $Y=1.835
+ $X2=7.685 $Y2=2.675
r134 2 37 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=8.35
+ $Y=2.465 $X2=8.485 $Y2=2.675
r135 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.64
+ $Y=0.405 $X2=8.78 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_1%A_1266_74# 1 2 9 13 15 16 18 21 23 24 25 27
+ 28 29 30 32 35 37 38 42 43 44 49 52
c155 49 0 1.44605e-19 $X=6.565 $Y=1.6
c156 44 0 1.4888e-19 $X=7.635 $Y=1.6
c157 43 0 3.23044e-20 $X=8.52 $Y=1.6
c158 42 0 1.00866e-19 $X=7.55 $Y=2.475
r159 53 59 3.86218 $w=3.12e-07 $l=2.5e-08 $layer=POLY_cond $X=8.685 $Y=1.52
+ $X2=8.71 $Y2=1.52
r160 53 57 18.5385 $w=3.12e-07 $l=1.2e-07 $layer=POLY_cond $X=8.685 $Y=1.52
+ $X2=8.565 $Y2=1.52
r161 52 55 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=8.685 $Y=1.52
+ $X2=8.685 $Y2=1.6
r162 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.685
+ $Y=1.52 $X2=8.685 $Y2=1.52
r163 47 49 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=6.405 $Y=1.6
+ $X2=6.565 $Y2=1.6
r164 43 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.52 $Y=1.6
+ $X2=8.685 $Y2=1.6
r165 43 44 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=8.52 $Y=1.6
+ $X2=7.635 $Y2=1.6
r166 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.55 $Y=1.685
+ $X2=7.635 $Y2=1.6
r167 41 42 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=7.55 $Y=1.685
+ $X2=7.55 $Y2=2.475
r168 38 40 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=6.65 $Y=2.64
+ $X2=7.04 $Y2=2.64
r169 37 42 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.465 $Y=2.64
+ $X2=7.55 $Y2=2.475
r170 37 40 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=7.465 $Y=2.64
+ $X2=7.04 $Y2=2.64
r171 33 46 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.49 $Y=0.72
+ $X2=6.405 $Y2=0.72
r172 33 35 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=6.49 $Y=0.72
+ $X2=6.915 $Y2=0.72
r173 32 38 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.565 $Y=2.475
+ $X2=6.65 $Y2=2.64
r174 31 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.565 $Y=1.685
+ $X2=6.565 $Y2=1.6
r175 31 32 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=6.565 $Y=1.685
+ $X2=6.565 $Y2=2.475
r176 30 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.405 $Y=1.515
+ $X2=6.405 $Y2=1.6
r177 29 46 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.405 $Y=0.845
+ $X2=6.405 $Y2=0.72
r178 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.405 $Y=0.845
+ $X2=6.405 $Y2=1.515
r179 25 27 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=9.555 $Y=0.995
+ $X2=9.555 $Y2=0.645
r180 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.48 $Y=1.07
+ $X2=9.555 $Y2=0.995
r181 23 24 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=9.48 $Y=1.07
+ $X2=9.305 $Y2=1.07
r182 19 28 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=9.245 $Y=1.685
+ $X2=9.245 $Y2=1.52
r183 19 21 303.194 $w=1.8e-07 $l=7.8e-07 $layer=POLY_cond $X=9.245 $Y=1.685
+ $X2=9.245 $Y2=2.465
r184 18 28 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=9.23 $Y=1.355
+ $X2=9.245 $Y2=1.52
r185 17 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.23 $Y=1.145
+ $X2=9.305 $Y2=1.07
r186 17 18 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=9.23 $Y=1.145
+ $X2=9.23 $Y2=1.355
r187 16 59 13.3422 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.8 $Y=1.52 $X2=8.71
+ $Y2=1.52
r188 15 28 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.155 $Y=1.52
+ $X2=9.245 $Y2=1.52
r189 15 16 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=9.155 $Y=1.52
+ $X2=8.8 $Y2=1.52
r190 11 59 15.628 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.71 $Y=1.685
+ $X2=8.71 $Y2=1.52
r191 11 13 384.823 $w=1.8e-07 $l=9.9e-07 $layer=POLY_cond $X=8.71 $Y=1.685
+ $X2=8.71 $Y2=2.675
r192 7 57 19.893 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.565 $Y=1.355
+ $X2=8.565 $Y2=1.52
r193 7 9 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=8.565 $Y=1.355
+ $X2=8.565 $Y2=0.615
r194 2 40 300 $w=1.7e-07 $l=9.98299e-07 $layer=licon1_PDIFF $count=2 $X=6.475
+ $Y=1.885 $X2=7.04 $Y2=2.64
r195 1 46 182 $w=1.7e-07 $l=3.79671e-07 $layer=licon1_NDIFF $count=1 $X=6.33
+ $Y=0.37 $X2=6.485 $Y2=0.68
r196 1 35 182 $w=1.7e-07 $l=7.23585e-07 $layer=licon1_NDIFF $count=1 $X=6.33
+ $Y=0.37 $X2=6.915 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_1%A_1867_409# 1 2 7 9 12 14 15 18 22 27
r51 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.77
+ $Y=1.55 $X2=9.77 $Y2=1.55
r52 24 27 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=9.47 $Y=1.55 $X2=9.77
+ $Y2=1.55
r53 20 27 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.77 $Y=1.385
+ $X2=9.77 $Y2=1.55
r54 20 22 25.8427 $w=3.28e-07 $l=7.4e-07 $layer=LI1_cond $X=9.77 $Y=1.385
+ $X2=9.77 $Y2=0.645
r55 16 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.47 $Y=1.715
+ $X2=9.47 $Y2=1.55
r56 16 18 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=9.47 $Y=1.715
+ $X2=9.47 $Y2=2.19
r57 14 28 117.157 $w=3.3e-07 $l=6.7e-07 $layer=POLY_cond $X=10.44 $Y=1.55
+ $X2=9.77 $Y2=1.55
r58 14 15 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=10.44 $Y=1.55
+ $X2=10.53 $Y2=1.55
r59 10 15 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=10.545 $Y=1.385
+ $X2=10.53 $Y2=1.55
r60 10 12 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=10.545 $Y=1.385
+ $X2=10.545 $Y2=0.74
r61 7 15 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=10.53 $Y=1.715
+ $X2=10.53 $Y2=1.55
r62 7 9 183.428 $w=1.8e-07 $l=6.85e-07 $layer=POLY_cond $X=10.53 $Y=1.715
+ $X2=10.53 $Y2=2.4
r63 2 18 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=9.335
+ $Y=2.045 $X2=9.47 $Y2=2.19
r64 1 22 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=9.63
+ $Y=0.37 $X2=9.77 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_1%VPWR 1 2 3 4 5 6 7 8 25 27 31 35 39 41 45 51
+ 53 57 59 61 65 67 72 77 85 93 105 108 111 114 117 120 124
r137 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r138 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r139 118 121 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r140 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r141 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r142 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r143 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r144 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r145 100 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r146 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r147 97 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r148 97 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r149 96 99 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r150 96 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r151 94 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.185 $Y=3.33
+ $X2=9.02 $Y2=3.33
r152 94 96 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=9.185 $Y=3.33
+ $X2=9.36 $Y2=3.33
r153 93 123 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=10.595 $Y=3.33
+ $X2=10.817 $Y2=3.33
r154 93 99 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.595 $Y=3.33
+ $X2=10.32 $Y2=3.33
r155 92 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r156 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r157 89 92 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=7.44 $Y2=3.33
r158 88 91 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=7.44
+ $Y2=3.33
r159 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r160 86 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.81 $Y=3.33
+ $X2=5.645 $Y2=3.33
r161 86 88 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.81 $Y=3.33 $X2=6
+ $Y2=3.33
r162 85 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.805 $Y=3.33
+ $X2=7.97 $Y2=3.33
r163 85 91 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.805 $Y=3.33
+ $X2=7.44 $Y2=3.33
r164 84 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r165 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r166 81 84 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r167 81 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r168 80 83 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r169 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r170 78 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=2.15 $Y2=3.33
r171 78 80 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=2.64 $Y2=3.33
r172 77 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.39 $Y=3.33
+ $X2=4.555 $Y2=3.33
r173 77 83 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.39 $Y=3.33
+ $X2=4.08 $Y2=3.33
r174 76 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r175 76 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r176 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r177 73 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.17 $Y2=3.33
r178 73 75 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.68 $Y2=3.33
r179 72 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=2.15 $Y2=3.33
r180 72 75 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=1.68 $Y2=3.33
r181 71 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r182 71 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r183 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r184 68 102 4.02368 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.177 $Y2=3.33
r185 68 70 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.72 $Y2=3.33
r186 67 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.17 $Y2=3.33
r187 67 70 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.72 $Y2=3.33
r188 65 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r189 65 112 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r190 65 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r191 61 64 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=10.76 $Y=1.985
+ $X2=10.76 $Y2=2.815
r192 59 123 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.76 $Y=3.245
+ $X2=10.817 $Y2=3.33
r193 59 64 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.76 $Y=3.245
+ $X2=10.76 $Y2=2.815
r194 55 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.02 $Y=3.245
+ $X2=9.02 $Y2=3.33
r195 55 57 30.9064 $w=3.28e-07 $l=8.85e-07 $layer=LI1_cond $X=9.02 $Y=3.245
+ $X2=9.02 $Y2=2.36
r196 54 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.135 $Y=3.33
+ $X2=7.97 $Y2=3.33
r197 53 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.855 $Y=3.33
+ $X2=9.02 $Y2=3.33
r198 53 54 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=8.855 $Y=3.33
+ $X2=8.135 $Y2=3.33
r199 49 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.97 $Y=3.245
+ $X2=7.97 $Y2=3.33
r200 49 51 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=7.97 $Y=3.245
+ $X2=7.97 $Y2=2.675
r201 45 48 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.645 $Y=1.91
+ $X2=5.645 $Y2=2.59
r202 43 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.645 $Y=3.245
+ $X2=5.645 $Y2=3.33
r203 43 48 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=5.645 $Y=3.245
+ $X2=5.645 $Y2=2.59
r204 42 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.72 $Y=3.33
+ $X2=4.555 $Y2=3.33
r205 41 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.48 $Y=3.33
+ $X2=5.645 $Y2=3.33
r206 41 42 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=5.48 $Y=3.33
+ $X2=4.72 $Y2=3.33
r207 37 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.555 $Y=3.245
+ $X2=4.555 $Y2=3.33
r208 37 39 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=4.555 $Y=3.245
+ $X2=4.555 $Y2=2.825
r209 33 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=3.245
+ $X2=2.15 $Y2=3.33
r210 33 35 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=2.15 $Y=3.245
+ $X2=2.15 $Y2=2.87
r211 29 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=3.33
r212 29 31 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=2.89
r213 25 102 3.11948 $w=2.5e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.23 $Y=3.245
+ $X2=0.177 $Y2=3.33
r214 25 27 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=0.23 $Y=3.245
+ $X2=0.23 $Y2=2.82
r215 8 64 400 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=1 $X=10.62
+ $Y=1.84 $X2=10.76 $Y2=2.815
r216 8 61 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.62
+ $Y=1.84 $X2=10.76 $Y2=1.985
r217 7 57 300 $w=1.7e-07 $l=2.67395e-07 $layer=licon1_PDIFF $count=2 $X=8.8
+ $Y=2.465 $X2=9.02 $Y2=2.36
r218 6 51 600 $w=1.7e-07 $l=2.91633e-07 $layer=licon1_PDIFF $count=1 $X=7.775
+ $Y=2.465 $X2=7.97 $Y2=2.675
r219 5 48 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.5
+ $Y=1.735 $X2=5.645 $Y2=2.59
r220 5 45 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.5
+ $Y=1.735 $X2=5.645 $Y2=1.91
r221 4 39 600 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=2.315 $X2=4.555 $Y2=2.825
r222 3 35 600 $w=1.7e-07 $l=1.00022e-06 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.935 $X2=2.15 $Y2=2.87
r223 2 31 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=2.615 $X2=1.17 $Y2=2.89
r224 1 27 600 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.615 $X2=0.27 $Y2=2.82
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_1%A_30_78# 1 2 3 4 13 17 20 21 25 27 30 32 36
+ 38 43
c112 27 0 1.38808e-19 $X=3.595 $Y=2.27
r113 38 40 0.257384 $w=2.37e-07 $l=5e-09 $layer=LI1_cond $X=3.165 $Y=2.53
+ $X2=3.165 $Y2=2.535
r114 37 38 13.384 $w=2.37e-07 $l=2.6e-07 $layer=LI1_cond $X=3.165 $Y=2.27
+ $X2=3.165 $Y2=2.53
r115 32 34 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.295 $Y=0.6
+ $X2=0.295 $Y2=0.745
r116 29 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.68 $Y=1.37
+ $X2=3.68 $Y2=1.285
r117 29 30 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=3.68 $Y=1.37
+ $X2=3.68 $Y2=2.185
r118 28 37 2.684 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.305 $Y=2.27
+ $X2=3.165 $Y2=2.27
r119 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.595 $Y=2.27
+ $X2=3.68 $Y2=2.185
r120 27 28 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.595 $Y=2.27
+ $X2=3.305 $Y2=2.27
r121 23 43 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.35 $Y=1.285
+ $X2=3.68 $Y2=1.285
r122 23 25 11.9218 $w=2.88e-07 $l=3e-07 $layer=LI1_cond $X=3.35 $Y=1.2 $X2=3.35
+ $Y2=0.9
r123 22 36 2.60907 $w=1.7e-07 $l=3.64966e-07 $layer=LI1_cond $X=0.885 $Y=2.53
+ $X2=0.525 $Y2=2.52
r124 21 38 2.684 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.025 $Y=2.53
+ $X2=3.165 $Y2=2.53
r125 21 22 139.615 $w=1.68e-07 $l=2.14e-06 $layer=LI1_cond $X=3.025 $Y=2.53
+ $X2=0.885 $Y2=2.53
r126 20 36 3.84343 $w=2.4e-07 $l=2.8e-07 $layer=LI1_cond $X=0.77 $Y=2.445
+ $X2=0.525 $Y2=2.52
r127 19 20 105.364 $w=1.68e-07 $l=1.615e-06 $layer=LI1_cond $X=0.77 $Y=0.83
+ $X2=0.77 $Y2=2.445
r128 15 36 3.84343 $w=2.4e-07 $l=2.10178e-07 $layer=LI1_cond $X=0.68 $Y=2.65
+ $X2=0.525 $Y2=2.52
r129 15 17 6.31985 $w=3.08e-07 $l=1.7e-07 $layer=LI1_cond $X=0.68 $Y=2.65
+ $X2=0.68 $Y2=2.82
r130 14 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.46 $Y=0.745
+ $X2=0.295 $Y2=0.745
r131 13 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.685 $Y=0.745
+ $X2=0.77 $Y2=0.83
r132 13 14 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.685 $Y=0.745
+ $X2=0.46 $Y2=0.745
r133 4 40 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=3.045
+ $Y=2.315 $X2=3.19 $Y2=2.535
r134 3 17 600 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.615 $X2=0.72 $Y2=2.82
r135 2 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.15
+ $Y=0.69 $X2=3.29 $Y2=0.9
r136 1 32 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.39 $X2=0.295 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_1%Q 1 2 9 13 14 15 16 29
r28 20 32 3.16106 $w=6.98e-07 $l=1.85e-07 $layer=LI1_cond $X=10.075 $Y=2.235
+ $X2=10.075 $Y2=2.05
r29 16 26 0.683473 $w=6.98e-07 $l=4e-08 $layer=LI1_cond $X=10.075 $Y=2.775
+ $X2=10.075 $Y2=2.815
r30 15 16 6.32213 $w=6.98e-07 $l=3.7e-07 $layer=LI1_cond $X=10.075 $Y=2.405
+ $X2=10.075 $Y2=2.775
r31 15 20 2.90476 $w=6.98e-07 $l=1.7e-07 $layer=LI1_cond $X=10.075 $Y=2.405
+ $X2=10.075 $Y2=2.235
r32 14 32 0.256303 $w=6.98e-07 $l=1.5e-08 $layer=LI1_cond $X=10.075 $Y=2.035
+ $X2=10.075 $Y2=2.05
r33 14 29 7.51816 $w=6.98e-07 $l=1.5e-07 $layer=LI1_cond $X=10.075 $Y=2.035
+ $X2=10.075 $Y2=1.885
r34 13 29 33.4652 $w=2.58e-07 $l=7.55e-07 $layer=LI1_cond $X=10.295 $Y=1.13
+ $X2=10.295 $Y2=1.885
r35 7 13 6.31279 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=10.33 $Y=0.965
+ $X2=10.33 $Y2=1.13
r36 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=10.33 $Y=0.965
+ $X2=10.33 $Y2=0.515
r37 2 32 400 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=10.115
+ $Y=1.84 $X2=10.26 $Y2=2.05
r38 2 26 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=10.115
+ $Y=1.84 $X2=10.26 $Y2=2.815
r39 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=10.185
+ $Y=0.37 $X2=10.33 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_1%VGND 1 2 3 4 5 6 21 25 29 33 35 37 40 41 42
+ 48 52 60 68 73 79 89 92 96
c103 29 0 3.23044e-20 $X=7.91 $Y=0.615
r104 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r105 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r106 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r107 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r108 77 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r109 77 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.36 $Y2=0
r110 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r111 74 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.425 $Y=0 $X2=9.3
+ $Y2=0
r112 74 76 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=9.425 $Y=0
+ $X2=10.32 $Y2=0
r113 73 95 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=10.675 $Y=0
+ $X2=10.857 $Y2=0
r114 73 76 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=10.675 $Y=0
+ $X2=10.32 $Y2=0
r115 72 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r116 72 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=7.92
+ $Y2=0
r117 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r118 69 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.075 $Y=0 $X2=7.91
+ $Y2=0
r119 69 71 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=8.075 $Y=0
+ $X2=8.88 $Y2=0
r120 68 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.175 $Y=0 $X2=9.3
+ $Y2=0
r121 68 71 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.175 $Y=0 $X2=8.88
+ $Y2=0
r122 67 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r123 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r124 63 66 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=7.44
+ $Y2=0
r125 61 63 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.31 $Y=0 $X2=5.52
+ $Y2=0
r126 60 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.745 $Y=0 $X2=7.91
+ $Y2=0
r127 60 66 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.44 $Y2=0
r128 59 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r129 58 59 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r130 56 59 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.56 $Y2=0
r131 56 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r132 55 58 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r133 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r134 53 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.38 $Y=0 $X2=2.215
+ $Y2=0
r135 53 55 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.38 $Y=0 $X2=2.64
+ $Y2=0
r136 52 86 9.04449 $w=3.93e-07 $l=3.1e-07 $layer=LI1_cond $X=5.112 $Y=0
+ $X2=5.112 $Y2=0.31
r137 52 61 5.70203 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=5.112 $Y=0 $X2=5.31
+ $Y2=0
r138 52 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r139 52 58 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.915 $Y=0
+ $X2=4.56 $Y2=0
r140 51 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r141 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r142 48 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.05 $Y=0 $X2=2.215
+ $Y2=0
r143 48 50 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.05 $Y=0 $X2=1.68
+ $Y2=0
r144 46 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r145 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r146 42 67 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=7.44 $Y2=0
r147 42 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r148 42 63 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r149 40 45 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=0.72
+ $Y2=0
r150 40 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=1.155
+ $Y2=0
r151 39 50 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.68
+ $Y2=0
r152 39 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.155
+ $Y2=0
r153 35 95 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.8 $Y=0.085
+ $X2=10.857 $Y2=0
r154 35 37 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.8 $Y=0.085
+ $X2=10.8 $Y2=0.515
r155 31 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.3 $Y=0.085
+ $X2=9.3 $Y2=0
r156 31 33 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=9.3 $Y=0.085
+ $X2=9.3 $Y2=0.595
r157 27 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0
r158 27 29 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0.615
r159 23 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.215 $Y=0.085
+ $X2=2.215 $Y2=0
r160 23 25 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=2.215 $Y=0.085
+ $X2=2.215 $Y2=0.715
r161 19 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0
r162 19 21 23.7403 $w=2.48e-07 $l=5.15e-07 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0.6
r163 6 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.62
+ $Y=0.37 $X2=10.76 $Y2=0.515
r164 5 33 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=9.195
+ $Y=0.37 $X2=9.34 $Y2=0.595
r165 4 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.77
+ $Y=0.405 $X2=7.91 $Y2=0.615
r166 3 86 182 $w=1.7e-07 $l=4.89285e-07 $layer=licon1_NDIFF $count=1 $X=4.86
+ $Y=0.69 $X2=5.11 $Y2=0.31
r167 2 25 182 $w=1.7e-07 $l=2.37539e-07 $layer=licon1_NDIFF $count=1 $X=2.03
+ $Y=0.595 $X2=2.215 $Y2=0.715
r168 1 21 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.975
+ $Y=0.39 $X2=1.115 $Y2=0.6
.ends


* File: sky130_fd_sc_ms__dfstp_4.pex.spice
* Created: Wed Sep  2 12:03:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DFSTP_4%D 2 5 9 11 12 16 17 20
c34 17 0 1.42976e-19 $X=0.64 $Y=1.145
r35 20 22 39.7991 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.825
+ $X2=0.61 $Y2=1.99
r36 20 21 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.825 $X2=0.64 $Y2=1.825
r37 16 18 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.145
+ $X2=0.61 $Y2=0.98
r38 16 17 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.145 $X2=0.64 $Y2=1.145
r39 12 21 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=0.64 $Y=1.665
+ $X2=0.64 $Y2=1.825
r40 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.665
r41 11 17 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.145
r42 9 18 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.495 $Y=0.58 $X2=0.495
+ $Y2=0.98
r43 5 22 287.645 $w=1.8e-07 $l=7.4e-07 $layer=POLY_cond $X=0.505 $Y=2.73
+ $X2=0.505 $Y2=1.99
r44 2 20 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=0.61 $Y=1.795 $X2=0.61
+ $Y2=1.825
r45 1 16 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=0.61 $Y=1.175 $X2=0.61
+ $Y2=1.145
r46 1 2 88.4142 $w=3.9e-07 $l=6.2e-07 $layer=POLY_cond $X=0.61 $Y=1.175 $X2=0.61
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_4%CLK 3 6 8 11 13
c38 11 0 2.57177e-19 $X=1.465 $Y=1.385
c39 6 0 1.42976e-19 $X=1.515 $Y=2.4
r40 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.385
+ $X2=1.465 $Y2=1.55
r41 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.385
+ $X2=1.465 $Y2=1.22
r42 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.465
+ $Y=1.385 $X2=1.465 $Y2=1.385
r43 8 12 6.69663 $w=3.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=1.465 $Y2=1.365
r44 6 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.515 $Y=2.4
+ $X2=1.515 $Y2=1.55
r45 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.485 $Y=0.74
+ $X2=1.485 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_4%A_398_74# 1 2 9 11 15 19 22 26 30 32 33 34
+ 35 38 39 45 46 49 50 53 54 55 57 58 59 63 64 65 68 69 71 72 73 76 78 88 92
c261 72 0 8.24247e-20 $X=6.53 $Y=1.285
c262 71 0 2.80241e-20 $X=6.53 $Y=1.285
c263 59 0 1.64109e-19 $X=5.51 $Y=2.18
c264 22 0 1.74759e-19 $X=7.325 $Y=2.75
r265 82 83 97.5202 $w=3.3e-07 $l=4.9e-07 $layer=POLY_cond $X=2.95 $Y=1.635
+ $X2=2.95 $Y2=2.125
r266 77 92 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=7.21 $Y=2.185
+ $X2=7.325 $Y2=2.185
r267 76 78 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.21 $Y=2.185
+ $X2=7.21 $Y2=2.02
r268 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.21
+ $Y=2.185 $X2=7.21 $Y2=2.185
r269 72 88 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.53 $Y=1.285
+ $X2=6.53 $Y2=1.12
r270 71 74 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=6.5 $Y=1.285
+ $X2=6.5 $Y2=1.45
r271 71 73 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=6.5 $Y=1.285
+ $X2=6.5 $Y2=1.12
r272 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.53
+ $Y=1.285 $X2=6.53 $Y2=1.285
r273 66 78 104.059 $w=1.68e-07 $l=1.595e-06 $layer=LI1_cond $X=7.29 $Y=0.425
+ $X2=7.29 $Y2=2.02
r274 64 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.205 $Y=0.34
+ $X2=7.29 $Y2=0.425
r275 64 65 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.205 $Y=0.34
+ $X2=6.475 $Y2=0.34
r276 63 74 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=6.39 $Y=2.095
+ $X2=6.39 $Y2=1.45
r277 60 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.39 $Y=0.425
+ $X2=6.475 $Y2=0.34
r278 60 73 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.39 $Y=0.425
+ $X2=6.39 $Y2=1.12
r279 58 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.305 $Y=2.18
+ $X2=6.39 $Y2=2.095
r280 58 59 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=6.305 $Y=2.18
+ $X2=5.51 $Y2=2.18
r281 56 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.425 $Y=2.265
+ $X2=5.51 $Y2=2.18
r282 56 57 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.425 $Y=2.265
+ $X2=5.425 $Y2=2.905
r283 54 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.34 $Y=2.99
+ $X2=5.425 $Y2=2.905
r284 54 55 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.34 $Y=2.99
+ $X2=4.685 $Y2=2.99
r285 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.6 $Y=2.905
+ $X2=4.685 $Y2=2.99
r286 52 53 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.6 $Y=2.335
+ $X2=4.6 $Y2=2.905
r287 51 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.795 $Y=2.25
+ $X2=3.71 $Y2=2.25
r288 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.515 $Y=2.25
+ $X2=4.6 $Y2=2.335
r289 50 51 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=4.515 $Y=2.25
+ $X2=3.795 $Y2=2.25
r290 48 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.71 $Y=2.335
+ $X2=3.71 $Y2=2.25
r291 48 49 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.71 $Y=2.335
+ $X2=3.71 $Y2=2.905
r292 46 84 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=3.71 $Y=1.635
+ $X2=3.585 $Y2=1.635
r293 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.71
+ $Y=1.635 $X2=3.71 $Y2=1.635
r294 43 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.71 $Y=2.165
+ $X2=3.71 $Y2=2.25
r295 43 45 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.71 $Y=2.165
+ $X2=3.71 $Y2=1.635
r296 41 68 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=3.03 $Y=0.425
+ $X2=3.03 $Y2=1.455
r297 39 82 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.95 $Y=1.62
+ $X2=2.95 $Y2=1.635
r298 38 68 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.95 $Y=1.62
+ $X2=2.95 $Y2=1.455
r299 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.95
+ $Y=1.62 $X2=2.95 $Y2=1.62
r300 34 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.625 $Y=2.99
+ $X2=3.71 $Y2=2.905
r301 34 35 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=3.625 $Y=2.99
+ $X2=2.275 $Y2=2.99
r302 32 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.945 $Y=0.34
+ $X2=3.03 $Y2=0.425
r303 32 33 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.945 $Y=0.34
+ $X2=2.215 $Y2=0.34
r304 28 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.19 $Y=2.905
+ $X2=2.275 $Y2=2.99
r305 28 30 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.19 $Y=2.905
+ $X2=2.19 $Y2=2.575
r306 24 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.13 $Y=0.425
+ $X2=2.215 $Y2=0.34
r307 24 26 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.13 $Y=0.425
+ $X2=2.13 $Y2=0.515
r308 20 92 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.325 $Y=2.35
+ $X2=7.325 $Y2=2.185
r309 20 22 155.484 $w=1.8e-07 $l=4e-07 $layer=POLY_cond $X=7.325 $Y=2.35
+ $X2=7.325 $Y2=2.75
r310 19 88 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.595 $Y=0.69
+ $X2=6.595 $Y2=1.12
r311 13 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.585 $Y=1.47
+ $X2=3.585 $Y2=1.635
r312 13 15 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=3.585 $Y=1.47
+ $X2=3.585 $Y2=0.58
r313 12 82 2.83073 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.115 $Y=1.635
+ $X2=2.95 $Y2=1.635
r314 11 84 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.51 $Y=1.635
+ $X2=3.585 $Y2=1.635
r315 11 12 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=3.51 $Y=1.635
+ $X2=3.115 $Y2=1.635
r316 9 83 155.484 $w=1.8e-07 $l=4e-07 $layer=POLY_cond $X=3.005 $Y=2.525
+ $X2=3.005 $Y2=2.125
r317 2 30 600 $w=1.7e-07 $l=7.99656e-07 $layer=licon1_PDIFF $count=1 $X=2.055
+ $Y=1.84 $X2=2.19 $Y2=2.575
r318 1 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.99
+ $Y=0.37 $X2=2.13 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_4%A_767_402# 1 2 9 11 13 14 15 17 18 21 24 26
+ 33 38
c85 38 0 1.30099e-19 $X=4.395 $Y=0.975
c86 18 0 1.30611e-19 $X=4.855 $Y=1.867
c87 9 0 1.2346e-19 $X=3.925 $Y=2.525
r88 30 33 3.79782 $w=4.38e-07 $l=1.45e-07 $layer=LI1_cond $X=4.94 $Y=2.515
+ $X2=5.085 $Y2=2.515
r89 27 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.395 $Y=1.065
+ $X2=4.395 $Y2=1.23
r90 27 38 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.395 $Y=1.065
+ $X2=4.395 $Y2=0.975
r91 26 29 14.8027 $w=3.75e-07 $l=4.55e-07 $layer=LI1_cond $X=4.395 $Y=0.925
+ $X2=4.85 $Y2=0.925
r92 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.395
+ $Y=1.065 $X2=4.395 $Y2=1.065
r93 24 30 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=4.94 $Y=2.295
+ $X2=4.94 $Y2=2.515
r94 23 24 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.94 $Y=1.995 $X2=4.94
+ $Y2=2.295
r95 21 37 3.80126 $w=3.17e-07 $l=2.5e-08 $layer=POLY_cond $X=4.28 $Y=1.93
+ $X2=4.305 $Y2=1.93
r96 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.28
+ $Y=1.865 $X2=4.28 $Y2=1.865
r97 18 23 7.17723 $w=2.55e-07 $l=1.65118e-07 $layer=LI1_cond $X=4.855 $Y=1.867
+ $X2=4.94 $Y2=1.995
r98 18 20 25.9865 $w=2.53e-07 $l=5.75e-07 $layer=LI1_cond $X=4.855 $Y=1.867
+ $X2=4.28 $Y2=1.867
r99 17 37 20.269 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=4.305 $Y=1.7
+ $X2=4.305 $Y2=1.93
r100 17 41 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=4.305 $Y=1.7 $X2=4.305
+ $Y2=1.23
r101 14 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.23 $Y=0.975
+ $X2=4.395 $Y2=0.975
r102 14 15 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=4.23 $Y=0.975
+ $X2=4.05 $Y2=0.975
r103 11 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.975 $Y=0.9
+ $X2=4.05 $Y2=0.975
r104 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.975 $Y=0.9
+ $X2=3.975 $Y2=0.58
r105 7 21 53.9779 $w=3.17e-07 $l=4.55714e-07 $layer=POLY_cond $X=3.925 $Y=2.16
+ $X2=4.28 $Y2=1.93
r106 7 9 141.879 $w=1.8e-07 $l=3.65e-07 $layer=POLY_cond $X=3.925 $Y=2.16
+ $X2=3.925 $Y2=2.525
r107 2 33 600 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_PDIFF $count=1 $X=4.95
+ $Y=2.315 $X2=5.085 $Y2=2.515
r108 1 29 182 $w=1.7e-07 $l=2.70416e-07 $layer=licon1_NDIFF $count=1 $X=4.67
+ $Y=0.59 $X2=4.85 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_4%A_612_74# 1 2 9 11 13 16 20 24 28 30 32 35
+ 36 38 39 44 49 53 58
c136 44 0 2.27104e-19 $X=4.935 $Y=1.285
c137 35 0 1.2346e-19 $X=3.28 $Y=2.515
c138 9 0 1.64109e-19 $X=4.86 $Y=2.525
r139 53 62 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.97 $Y=1.365
+ $X2=5.97 $Y2=1.53
r140 53 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.97 $Y=1.365
+ $X2=5.97 $Y2=1.2
r141 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.97
+ $Y=1.365 $X2=5.97 $Y2=1.365
r142 49 52 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5.97 $Y=1.285 $X2=5.97
+ $Y2=1.365
r143 45 58 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.935 $Y=1.285
+ $X2=5.1 $Y2=1.285
r144 45 55 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.935 $Y=1.285
+ $X2=4.86 $Y2=1.285
r145 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.935
+ $Y=1.285 $X2=4.935 $Y2=1.285
r146 39 41 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.05 $Y=1.215
+ $X2=4.05 $Y2=1.485
r147 35 36 10.3362 $w=3.38e-07 $l=2.2e-07 $layer=LI1_cond $X=3.285 $Y=2.515
+ $X2=3.285 $Y2=2.295
r148 33 44 3.11056 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=5.025 $Y=1.285
+ $X2=4.897 $Y2=1.285
r149 32 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.805 $Y=1.285
+ $X2=5.97 $Y2=1.285
r150 32 33 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=5.805 $Y=1.285
+ $X2=5.025 $Y2=1.285
r151 31 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.135 $Y=1.485
+ $X2=4.05 $Y2=1.485
r152 30 44 9.03877 $w=2.53e-07 $l=2e-07 $layer=LI1_cond $X=4.897 $Y=1.485
+ $X2=4.897 $Y2=1.285
r153 30 31 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.77 $Y=1.485
+ $X2=4.135 $Y2=1.485
r154 29 38 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.535 $Y=1.215
+ $X2=3.41 $Y2=1.215
r155 28 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.965 $Y=1.215
+ $X2=4.05 $Y2=1.215
r156 28 29 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.965 $Y=1.215
+ $X2=3.535 $Y2=1.215
r157 26 38 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=3.37 $Y=1.3
+ $X2=3.41 $Y2=1.215
r158 26 36 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=3.37 $Y=1.3
+ $X2=3.37 $Y2=2.295
r159 22 38 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.41 $Y=1.13 $X2=3.41
+ $Y2=1.215
r160 22 24 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=3.41 $Y=1.13
+ $X2=3.41 $Y2=0.58
r161 20 61 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=6.05 $Y=0.69
+ $X2=6.05 $Y2=1.2
r162 16 62 274.04 $w=1.8e-07 $l=7.05e-07 $layer=POLY_cond $X=6.025 $Y=2.235
+ $X2=6.025 $Y2=1.53
r163 11 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.1 $Y=1.12
+ $X2=5.1 $Y2=1.285
r164 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.1 $Y=1.12 $X2=5.1
+ $Y2=0.8
r165 7 55 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.86 $Y=1.45
+ $X2=4.86 $Y2=1.285
r166 7 9 417.863 $w=1.8e-07 $l=1.075e-06 $layer=POLY_cond $X=4.86 $Y=1.45
+ $X2=4.86 $Y2=2.525
r167 2 35 600 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_PDIFF $count=1 $X=3.095
+ $Y=2.315 $X2=3.28 $Y2=2.515
r168 1 24 182 $w=1.7e-07 $l=4.01497e-07 $layer=licon1_NDIFF $count=1 $X=3.06
+ $Y=0.37 $X2=3.37 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_4%SET_B 3 7 9 11 12 13 16 18 19 20 25 31 32 37
c127 37 0 1.13172e-19 $X=8.35 $Y=1.345
c128 20 0 9.70053e-20 $X=5.665 $Y=1.665
c129 19 0 2.34318e-20 $X=8.255 $Y=1.665
c130 3 0 1.30611e-19 $X=5.31 $Y=2.525
r131 37 44 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=8.35 $Y=1.345
+ $X2=8.35 $Y2=1.665
r132 30 32 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=5.36 $Y=1.825
+ $X2=5.49 $Y2=1.825
r133 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.36
+ $Y=1.825 $X2=5.36 $Y2=1.825
r134 27 30 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=5.31 $Y=1.825
+ $X2=5.36 $Y2=1.825
r135 25 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=1.665
+ $X2=8.4 $Y2=1.665
r136 22 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.665
+ $X2=5.52 $Y2=1.665
r137 20 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=1.665
+ $X2=5.52 $Y2=1.665
r138 19 25 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=8.4 $Y2=1.665
r139 19 20 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=5.665 $Y2=1.665
r140 16 18 349.839 $w=1.8e-07 $l=9e-07 $layer=POLY_cond $X=8.195 $Y=2.75
+ $X2=8.195 $Y2=1.85
r141 13 18 45.5979 $w=4.1e-07 $l=2.05e-07 $layer=POLY_cond $X=8.31 $Y=1.645
+ $X2=8.31 $Y2=1.85
r142 12 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.35
+ $Y=1.345 $X2=8.35 $Y2=1.345
r143 12 13 35.2683 $w=4.1e-07 $l=2.6e-07 $layer=POLY_cond $X=8.31 $Y=1.385
+ $X2=8.31 $Y2=1.645
r144 9 12 86.4346 $w=2.37e-07 $l=6.27495e-07 $layer=POLY_cond $X=7.885 $Y=0.935
+ $X2=8.31 $Y2=1.385
r145 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.885 $Y=0.935
+ $X2=7.885 $Y2=0.65
r146 5 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.49 $Y=1.66
+ $X2=5.49 $Y2=1.825
r147 5 7 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.49 $Y=1.66 $X2=5.49
+ $Y2=0.8
r148 1 27 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.31 $Y=1.99
+ $X2=5.31 $Y2=1.825
r149 1 3 207.96 $w=1.8e-07 $l=5.35e-07 $layer=POLY_cond $X=5.31 $Y=1.99 $X2=5.31
+ $Y2=2.525
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_4%A_225_74# 1 2 9 13 16 17 19 20 23 27 29 34
+ 35 36 39 42 43 46 47 49 50 54 58 65
c173 54 0 1.60368e-19 $X=2.11 $Y=1.515
c174 35 0 2.80241e-20 $X=7.03 $Y=1.735
c175 27 0 1.25277e-19 $X=3.505 $Y=2.525
c176 16 0 1.99891e-19 $X=2.485 $Y=3.075
r177 64 65 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.29 $Y=1.895
+ $X2=1.455 $Y2=1.895
r178 61 64 7.5732 $w=3.48e-07 $l=2.3e-07 $layer=LI1_cond $X=1.06 $Y=1.895
+ $X2=1.29 $Y2=1.895
r179 58 60 17.8607 $w=4.58e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=0.515
+ $X2=1.205 $Y2=1.01
r180 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.11
+ $Y=1.515 $X2=2.11 $Y2=1.515
r181 52 54 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=2.11 $Y=1.72
+ $X2=2.11 $Y2=1.515
r182 50 52 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.945 $Y=1.805
+ $X2=2.11 $Y2=1.72
r183 50 65 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.945 $Y=1.805
+ $X2=1.455 $Y2=1.805
r184 49 61 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.06 $Y=1.72 $X2=1.06
+ $Y2=1.895
r185 49 60 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.06 $Y=1.72
+ $X2=1.06 $Y2=1.01
r186 46 55 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=2.41 $Y=1.515
+ $X2=2.11 $Y2=1.515
r187 43 46 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=2.485 $Y=1.14
+ $X2=2.485 $Y2=1.515
r188 41 55 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=2.055 $Y=1.515
+ $X2=2.11 $Y2=1.515
r189 41 42 3.90195 $w=3.3e-07 $l=1.08e-07 $layer=POLY_cond $X=2.055 $Y=1.515
+ $X2=1.947 $Y2=1.515
r190 37 39 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=7.105 $Y=1.66
+ $X2=7.105 $Y2=0.65
r191 35 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.03 $Y=1.735
+ $X2=7.105 $Y2=1.66
r192 35 36 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=7.03 $Y=1.735
+ $X2=6.62 $Y2=1.735
r193 32 34 239.056 $w=1.8e-07 $l=6.15e-07 $layer=POLY_cond $X=6.53 $Y=3.075
+ $X2=6.53 $Y2=2.46
r194 31 36 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.53 $Y=1.81
+ $X2=6.62 $Y2=1.735
r195 31 34 252.661 $w=1.8e-07 $l=6.5e-07 $layer=POLY_cond $X=6.53 $Y=1.81
+ $X2=6.53 $Y2=2.46
r196 30 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.595 $Y=3.15
+ $X2=3.505 $Y2=3.15
r197 29 32 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.44 $Y=3.15
+ $X2=6.53 $Y2=3.075
r198 29 30 1458.82 $w=1.5e-07 $l=2.845e-06 $layer=POLY_cond $X=6.44 $Y=3.15
+ $X2=3.595 $Y2=3.15
r199 25 47 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.505 $Y=3.075
+ $X2=3.505 $Y2=3.15
r200 25 27 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=3.505 $Y=3.075
+ $X2=3.505 $Y2=2.525
r201 21 23 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=2.985 $Y=1.065
+ $X2=2.985 $Y2=0.58
r202 19 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.415 $Y=3.15
+ $X2=3.505 $Y2=3.15
r203 19 20 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=3.415 $Y=3.15
+ $X2=2.56 $Y2=3.15
r204 18 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.56 $Y=1.14
+ $X2=2.485 $Y2=1.14
r205 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.91 $Y=1.14
+ $X2=2.985 $Y2=1.065
r206 17 18 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.91 $Y=1.14
+ $X2=2.56 $Y2=1.14
r207 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.485 $Y=3.075
+ $X2=2.56 $Y2=3.15
r208 15 46 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.485 $Y=1.68
+ $X2=2.485 $Y2=1.515
r209 15 16 715.309 $w=1.5e-07 $l=1.395e-06 $layer=POLY_cond $X=2.485 $Y=1.68
+ $X2=2.485 $Y2=3.075
r210 11 42 34.7346 $w=1.65e-07 $l=1.73767e-07 $layer=POLY_cond $X=1.965 $Y=1.68
+ $X2=1.947 $Y2=1.515
r211 11 13 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.965 $Y=1.68
+ $X2=1.965 $Y2=2.4
r212 7 42 34.7346 $w=1.65e-07 $l=1.80291e-07 $layer=POLY_cond $X=1.915 $Y=1.35
+ $X2=1.947 $Y2=1.515
r213 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.915 $Y=1.35
+ $X2=1.915 $Y2=0.74
r214 2 64 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.84 $X2=1.29 $Y2=1.985
r215 1 58 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.125
+ $Y=0.37 $X2=1.27 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_4%A_1484_62# 1 2 9 13 17 20 21 24 28 30 31 36
c82 36 0 1.90022e-19 $X=7.745 $Y=1.49
c83 13 0 2.73146e-19 $X=7.745 $Y=2.75
c84 9 0 1.13172e-19 $X=7.495 $Y=0.65
r85 30 31 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.395 $Y=2.815
+ $X2=9.395 $Y2=2.65
r86 26 28 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=9.365 $Y=1.01
+ $X2=9.285 $Y2=0.925
r87 26 31 106.995 $w=1.68e-07 $l=1.64e-06 $layer=LI1_cond $X=9.365 $Y=1.01
+ $X2=9.365 $Y2=2.65
r88 22 28 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.285 $Y=0.84
+ $X2=9.285 $Y2=0.925
r89 22 24 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=9.285 $Y=0.84
+ $X2=9.285 $Y2=0.65
r90 20 28 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.12 $Y=0.925
+ $X2=9.285 $Y2=0.925
r91 20 21 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=9.12 $Y=0.925
+ $X2=7.875 $Y2=0.925
r92 18 36 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=7.71 $Y=1.49
+ $X2=7.745 $Y2=1.49
r93 18 33 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=7.71 $Y=1.49
+ $X2=7.495 $Y2=1.49
r94 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.71
+ $Y=1.49 $X2=7.71 $Y2=1.49
r95 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.71 $Y=1.01
+ $X2=7.875 $Y2=0.925
r96 15 17 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.71 $Y=1.01
+ $X2=7.71 $Y2=1.49
r97 11 36 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.745 $Y=1.655
+ $X2=7.745 $Y2=1.49
r98 11 13 425.637 $w=1.8e-07 $l=1.095e-06 $layer=POLY_cond $X=7.745 $Y=1.655
+ $X2=7.745 $Y2=2.75
r99 7 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.495 $Y=1.325
+ $X2=7.495 $Y2=1.49
r100 7 9 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=7.495 $Y=1.325
+ $X2=7.495 $Y2=0.65
r101 2 30 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=9.26
+ $Y=2.54 $X2=9.395 $Y2=2.815
r102 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.145
+ $Y=0.44 $X2=9.285 $Y2=0.65
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_4%A_1324_392# 1 2 3 11 14 18 20 24 26 28 29 31
+ 33 34 38 40 41 42 43 47 49 53 54 58 65 69 71 75
c162 71 0 1.74759e-19 $X=7.63 $Y=2.395
c163 69 0 5.89928e-20 $X=6.95 $Y=1.705
c164 43 0 1.90022e-19 $X=8.255 $Y=2.395
c165 41 0 1.96733e-19 $X=7.545 $Y=2.565
c166 29 0 2.80689e-21 $X=10.505 $Y=1.69
c167 24 0 2.91921e-19 $X=10.13 $Y=0.74
r168 71 73 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.63 $Y=2.395
+ $X2=7.63 $Y2=2.565
r169 67 69 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.755 $Y=1.705
+ $X2=6.95 $Y2=1.705
r170 63 65 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=6.81 $Y=0.76
+ $X2=6.95 $Y2=0.76
r171 59 61 8.78706 $w=4.79e-07 $l=3.45e-07 $layer=LI1_cond $X=6.755 $Y=2.73
+ $X2=7.1 $Y2=2.73
r172 58 78 40.2621 $w=4.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.02 $Y=2.215
+ $X2=9.02 $Y2=2.38
r173 57 58 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.945
+ $Y=2.215 $X2=8.945 $Y2=2.215
r174 53 57 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=8.945 $Y=1.535
+ $X2=8.945 $Y2=2.215
r175 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.945
+ $Y=1.535 $X2=8.945 $Y2=1.535
r176 51 57 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=8.945 $Y=2.31
+ $X2=8.945 $Y2=2.215
r177 50 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.585 $Y=2.395
+ $X2=8.42 $Y2=2.395
r178 49 51 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.78 $Y=2.395
+ $X2=8.945 $Y2=2.31
r179 49 50 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=8.78 $Y=2.395
+ $X2=8.585 $Y2=2.395
r180 45 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.42 $Y=2.48
+ $X2=8.42 $Y2=2.395
r181 45 47 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=8.42 $Y=2.48
+ $X2=8.42 $Y2=2.75
r182 44 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.715 $Y=2.395
+ $X2=7.63 $Y2=2.395
r183 43 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.255 $Y=2.395
+ $X2=8.42 $Y2=2.395
r184 43 44 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=8.255 $Y=2.395
+ $X2=7.715 $Y2=2.395
r185 42 61 9.57821 $w=4.79e-07 $l=2.33345e-07 $layer=LI1_cond $X=7.265 $Y=2.565
+ $X2=7.1 $Y2=2.73
r186 41 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.545 $Y=2.565
+ $X2=7.63 $Y2=2.565
r187 41 42 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.545 $Y=2.565
+ $X2=7.265 $Y2=2.565
r188 40 69 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.95 $Y=1.62
+ $X2=6.95 $Y2=1.705
r189 39 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.95 $Y=0.925
+ $X2=6.95 $Y2=0.76
r190 39 40 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.95 $Y=0.925
+ $X2=6.95 $Y2=1.62
r191 36 59 6.88815 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=6.755 $Y=2.48
+ $X2=6.755 $Y2=2.73
r192 36 38 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.755 $Y=2.48
+ $X2=6.755 $Y2=2.135
r193 35 67 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.755 $Y=1.79
+ $X2=6.755 $Y2=1.705
r194 35 38 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.755 $Y=1.79
+ $X2=6.755 $Y2=2.135
r195 31 33 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=10.595 $Y=1.765
+ $X2=10.595 $Y2=2.26
r196 30 34 9.95731 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=10.235 $Y=1.69
+ $X2=10.055 $Y2=1.37
r197 29 31 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=10.505 $Y=1.69
+ $X2=10.595 $Y2=1.765
r198 29 30 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=10.505 $Y=1.69
+ $X2=10.235 $Y2=1.69
r199 26 34 14.284 $w=1.8e-07 $l=4.37693e-07 $layer=POLY_cond $X=10.145 $Y=1.765
+ $X2=10.055 $Y2=1.37
r200 26 28 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=10.145 $Y=1.765
+ $X2=10.145 $Y2=2.26
r201 22 34 14.284 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.13 $Y=1.37
+ $X2=10.055 $Y2=1.37
r202 22 24 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=10.13 $Y=1.37
+ $X2=10.13 $Y2=0.74
r203 21 54 8.93404 $w=2.45e-07 $l=2.4e-07 $layer=POLY_cond $X=9.26 $Y=1.492
+ $X2=9.02 $Y2=1.492
r204 20 34 9.95731 $w=2.45e-07 $l=1.22e-07 $layer=POLY_cond $X=10.055 $Y=1.492
+ $X2=10.055 $Y2=1.37
r205 20 21 201.552 $w=2.45e-07 $l=7.95e-07 $layer=POLY_cond $X=10.055 $Y=1.492
+ $X2=9.26 $Y2=1.492
r206 18 78 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=9.17 $Y=2.75
+ $X2=9.17 $Y2=2.38
r207 12 54 16.4793 $w=3.15e-07 $l=1.44859e-07 $layer=POLY_cond $X=9.07 $Y=1.37
+ $X2=9.02 $Y2=1.492
r208 12 14 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=9.07 $Y=1.37
+ $X2=9.07 $Y2=0.65
r209 11 58 8.35984 $w=4.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.02 $Y=2.14
+ $X2=9.02 $Y2=2.215
r210 10 54 16.4793 $w=3.15e-07 $l=1.23e-07 $layer=POLY_cond $X=9.02 $Y=1.615
+ $X2=9.02 $Y2=1.492
r211 10 11 58.5188 $w=4.8e-07 $l=5.25e-07 $layer=POLY_cond $X=9.02 $Y=1.615
+ $X2=9.02 $Y2=2.14
r212 3 47 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=8.285
+ $Y=2.54 $X2=8.42 $Y2=2.75
r213 2 61 300 $w=1.7e-07 $l=1.06837e-06 $layer=licon1_PDIFF $count=2 $X=6.62
+ $Y=1.96 $X2=7.1 $Y2=2.815
r214 2 38 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=6.62
+ $Y=1.96 $X2=6.755 $Y2=2.135
r215 1 63 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=6.67
+ $Y=0.37 $X2=6.81 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_4%A_1940_74# 1 2 7 9 10 11 12 14 17 21 23 25
+ 28 30 32 36 40 42 43 46 53 56
r117 62 63 12.0184 $w=3.81e-07 $l=9.5e-08 $layer=POLY_cond $X=11.92 $Y=1.437
+ $X2=12.015 $Y2=1.437
r118 57 58 6.95801 $w=3.81e-07 $l=5.5e-08 $layer=POLY_cond $X=11.06 $Y=1.437
+ $X2=11.115 $Y2=1.437
r119 54 62 11.3858 $w=3.81e-07 $l=9e-08 $layer=POLY_cond $X=11.83 $Y=1.437
+ $X2=11.92 $Y2=1.437
r120 54 60 33.5249 $w=3.81e-07 $l=2.65e-07 $layer=POLY_cond $X=11.83 $Y=1.437
+ $X2=11.565 $Y2=1.437
r121 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.83
+ $Y=1.485 $X2=11.83 $Y2=1.485
r122 51 60 52.5013 $w=3.81e-07 $l=4.15e-07 $layer=POLY_cond $X=11.15 $Y=1.437
+ $X2=11.565 $Y2=1.437
r123 51 58 4.42782 $w=3.81e-07 $l=3.5e-08 $layer=POLY_cond $X=11.15 $Y=1.437
+ $X2=11.115 $Y2=1.437
r124 50 53 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=11.15 $Y=1.485
+ $X2=11.83 $Y2=1.485
r125 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.15
+ $Y=1.485 $X2=11.15 $Y2=1.485
r126 48 56 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=10.535 $Y=1.485
+ $X2=10.37 $Y2=1.485
r127 48 50 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=10.535 $Y=1.485
+ $X2=11.15 $Y2=1.485
r128 44 56 0.364692 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=10.37 $Y=1.65
+ $X2=10.37 $Y2=1.485
r129 44 46 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=10.37 $Y=1.65
+ $X2=10.37 $Y2=1.985
r130 42 56 6.46576 $w=2.5e-07 $l=2.0106e-07 $layer=LI1_cond $X=10.205 $Y=1.405
+ $X2=10.37 $Y2=1.485
r131 42 43 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=10.205 $Y=1.405
+ $X2=10.01 $Y2=1.405
r132 38 43 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.845 $Y=1.32
+ $X2=10.01 $Y2=1.405
r133 38 40 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=9.845 $Y=1.32
+ $X2=9.845 $Y2=0.515
r134 34 65 20.3063 $w=1.8e-07 $l=2.13e-07 $layer=POLY_cond $X=12.465 $Y=1.65
+ $X2=12.465 $Y2=1.437
r135 34 36 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=12.465 $Y=1.65
+ $X2=12.465 $Y2=2.4
r136 30 65 8.85564 $w=3.81e-07 $l=7e-08 $layer=POLY_cond $X=12.395 $Y=1.437
+ $X2=12.465 $Y2=1.437
r137 30 63 48.0735 $w=3.81e-07 $l=3.8e-07 $layer=POLY_cond $X=12.395 $Y=1.437
+ $X2=12.015 $Y2=1.437
r138 30 32 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=12.395 $Y=1.32
+ $X2=12.395 $Y2=0.74
r139 26 63 20.3063 $w=1.8e-07 $l=2.13e-07 $layer=POLY_cond $X=12.015 $Y=1.65
+ $X2=12.015 $Y2=1.437
r140 26 28 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=12.015 $Y=1.65
+ $X2=12.015 $Y2=2.4
r141 23 62 24.6764 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=11.92 $Y=1.225
+ $X2=11.92 $Y2=1.437
r142 23 25 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=11.92 $Y=1.225
+ $X2=11.92 $Y2=0.74
r143 19 60 20.3063 $w=1.8e-07 $l=2.13e-07 $layer=POLY_cond $X=11.565 $Y=1.65
+ $X2=11.565 $Y2=1.437
r144 19 21 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=11.565 $Y=1.65
+ $X2=11.565 $Y2=2.4
r145 15 58 20.3063 $w=1.8e-07 $l=2.13e-07 $layer=POLY_cond $X=11.115 $Y=1.65
+ $X2=11.115 $Y2=1.437
r146 15 17 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=11.115 $Y=1.65
+ $X2=11.115 $Y2=2.4
r147 12 57 24.6764 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=11.06 $Y=1.225
+ $X2=11.06 $Y2=1.437
r148 12 14 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=11.06 $Y=1.225
+ $X2=11.06 $Y2=0.74
r149 10 57 27.8494 $w=3.81e-07 $l=1.70423e-07 $layer=POLY_cond $X=10.985 $Y=1.3
+ $X2=11.06 $Y2=1.437
r150 10 11 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=10.985 $Y=1.3
+ $X2=10.705 $Y2=1.3
r151 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.63 $Y=1.225
+ $X2=10.705 $Y2=1.3
r152 7 9 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=10.63 $Y=1.225
+ $X2=10.63 $Y2=0.74
r153 2 46 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=10.235
+ $Y=1.84 $X2=10.37 $Y2=1.985
r154 1 40 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=9.7
+ $Y=0.37 $X2=9.845 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_4%A_27_74# 1 2 3 4 15 18 21 23 25 28 29 30 31
+ 38
c69 25 0 1.25277e-19 $X=2.445 $Y=2.155
r70 35 38 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.53 $Y=0.76 $X2=2.69
+ $Y2=0.76
r71 31 33 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.71 $Y=2.155
+ $X2=1.71 $Y2=2.325
r72 27 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.53 $Y=0.925
+ $X2=2.53 $Y2=0.76
r73 27 28 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=2.53 $Y=0.925
+ $X2=2.53 $Y2=2.07
r74 26 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=2.155
+ $X2=1.71 $Y2=2.155
r75 25 42 11.3196 $w=3.88e-07 $l=4.68615e-07 $layer=LI1_cond $X=2.445 $Y=2.155
+ $X2=2.695 $Y2=2.515
r76 25 28 6.58872 $w=3.88e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.445 $Y=2.155
+ $X2=2.53 $Y2=2.07
r77 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.445 $Y=2.155
+ $X2=1.795 $Y2=2.155
r78 24 30 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=2.325
+ $X2=0.24 $Y2=2.325
r79 23 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=2.325
+ $X2=1.71 $Y2=2.325
r80 23 24 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=1.625 $Y=2.325
+ $X2=0.365 $Y2=2.325
r81 19 30 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.41 $X2=0.24
+ $Y2=2.325
r82 19 21 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=0.24 $Y=2.41
+ $X2=0.24 $Y2=2.73
r83 18 30 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.2 $Y=2.24
+ $X2=0.24 $Y2=2.325
r84 18 29 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=0.2 $Y=2.24 $X2=0.2
+ $Y2=0.81
r85 13 29 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=0.685
+ $X2=0.24 $Y2=0.81
r86 13 15 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=0.24 $Y=0.685
+ $X2=0.24 $Y2=0.58
r87 4 42 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=2.635
+ $Y=2.315 $X2=2.78 $Y2=2.515
r88 3 21 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.52 $X2=0.28 $Y2=2.73
r89 2 38 182 $w=1.7e-07 $l=4.56782e-07 $layer=licon1_NDIFF $count=1 $X=2.545
+ $Y=0.37 $X2=2.69 $Y2=0.76
r90 1 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_4%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 40 43 47 51
+ 55 57 61 67 69 71 76 79 80 81 83 88 93 105 109 114 119 124 130 133 136 139 142
+ 145 148 151 155
c174 37 0 1.99891e-19 $X=1.74 $Y=2.74
r175 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r176 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r177 148 149 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r178 146 149 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.8 $Y2=3.33
r179 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r180 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r181 139 140 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r182 136 137 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r183 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r184 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r185 128 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r186 128 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r187 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r188 125 151 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.955 $Y=3.33
+ $X2=11.79 $Y2=3.33
r189 125 127 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=11.955 $Y=3.33
+ $X2=12.24 $Y2=3.33
r190 124 154 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=12.525 $Y=3.33
+ $X2=12.742 $Y2=3.33
r191 124 127 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=12.525 $Y=3.33
+ $X2=12.24 $Y2=3.33
r192 123 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r193 123 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r194 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r195 120 148 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=11.005 $Y=3.33
+ $X2=10.865 $Y2=3.33
r196 120 122 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.005 $Y=3.33
+ $X2=11.28 $Y2=3.33
r197 119 151 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.625 $Y=3.33
+ $X2=11.79 $Y2=3.33
r198 119 122 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=11.625 $Y=3.33
+ $X2=11.28 $Y2=3.33
r199 118 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r200 118 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r201 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r202 115 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.03 $Y=3.33
+ $X2=8.905 $Y2=3.33
r203 115 117 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.03 $Y=3.33
+ $X2=9.36 $Y2=3.33
r204 114 145 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.755 $Y=3.33
+ $X2=9.88 $Y2=3.33
r205 114 117 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=9.755 $Y=3.33
+ $X2=9.36 $Y2=3.33
r206 113 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r207 113 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r208 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r209 110 139 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.055 $Y=3.33
+ $X2=7.97 $Y2=3.33
r210 110 112 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.055 $Y=3.33
+ $X2=8.4 $Y2=3.33
r211 109 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.78 $Y=3.33
+ $X2=8.905 $Y2=3.33
r212 109 112 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=8.78 $Y=3.33
+ $X2=8.4 $Y2=3.33
r213 107 108 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r214 105 139 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.885 $Y=3.33
+ $X2=7.97 $Y2=3.33
r215 105 107 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=7.885 $Y=3.33
+ $X2=6 $Y2=3.33
r216 104 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r217 104 137 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.08 $Y2=3.33
r218 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r219 101 136 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.155 $Y=3.33
+ $X2=4.07 $Y2=3.33
r220 101 103 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=4.155 $Y=3.33
+ $X2=5.52 $Y2=3.33
r221 100 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r222 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r223 97 100 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r224 97 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r225 96 99 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r226 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r227 94 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=1.74 $Y2=3.33
r228 94 96 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=2.16 $Y2=3.33
r229 93 136 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.985 $Y=3.33
+ $X2=4.07 $Y2=3.33
r230 93 99 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.985 $Y=3.33
+ $X2=3.6 $Y2=3.33
r231 92 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r232 92 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r233 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r234 89 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r235 89 91 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r236 88 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.74 $Y2=3.33
r237 88 91 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.2 $Y2=3.33
r238 86 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r239 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r240 83 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r241 83 85 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r242 81 140 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.92 $Y2=3.33
r243 81 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r244 79 103 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.68 $Y=3.33
+ $X2=5.52 $Y2=3.33
r245 79 80 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.68 $Y=3.33
+ $X2=5.81 $Y2=3.33
r246 78 107 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=5.94 $Y=3.33 $X2=6
+ $Y2=3.33
r247 78 80 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.94 $Y=3.33
+ $X2=5.81 $Y2=3.33
r248 73 76 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=4.07 $Y=2.63
+ $X2=4.165 $Y2=2.63
r249 69 154 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=12.69 $Y=3.245
+ $X2=12.742 $Y2=3.33
r250 69 71 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=12.69 $Y=3.245
+ $X2=12.69 $Y2=2.405
r251 65 151 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.79 $Y=3.245
+ $X2=11.79 $Y2=3.33
r252 65 67 31.7795 $w=3.28e-07 $l=9.1e-07 $layer=LI1_cond $X=11.79 $Y=3.245
+ $X2=11.79 $Y2=2.335
r253 61 64 34.1617 $w=2.78e-07 $l=8.3e-07 $layer=LI1_cond $X=10.865 $Y=1.985
+ $X2=10.865 $Y2=2.815
r254 59 148 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=10.865 $Y=3.245
+ $X2=10.865 $Y2=3.33
r255 59 64 17.6982 $w=2.78e-07 $l=4.3e-07 $layer=LI1_cond $X=10.865 $Y=3.245
+ $X2=10.865 $Y2=2.815
r256 58 145 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.005 $Y=3.33
+ $X2=9.88 $Y2=3.33
r257 57 148 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=10.725 $Y=3.33
+ $X2=10.865 $Y2=3.33
r258 57 58 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=10.725 $Y=3.33
+ $X2=10.005 $Y2=3.33
r259 53 145 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.88 $Y=3.245
+ $X2=9.88 $Y2=3.33
r260 53 55 58.0831 $w=2.48e-07 $l=1.26e-06 $layer=LI1_cond $X=9.88 $Y=3.245
+ $X2=9.88 $Y2=1.985
r261 49 142 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.905 $Y=3.245
+ $X2=8.905 $Y2=3.33
r262 49 51 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.905 $Y=3.245
+ $X2=8.905 $Y2=2.815
r263 45 139 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.97 $Y=3.245
+ $X2=7.97 $Y2=3.33
r264 45 47 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=7.97 $Y=3.245
+ $X2=7.97 $Y2=2.815
r265 41 80 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.81 $Y=3.245
+ $X2=5.81 $Y2=3.33
r266 41 43 28.5895 $w=2.58e-07 $l=6.45e-07 $layer=LI1_cond $X=5.81 $Y=3.245
+ $X2=5.81 $Y2=2.6
r267 40 136 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.07 $Y=3.245
+ $X2=4.07 $Y2=3.33
r268 39 73 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.07 $Y=2.755
+ $X2=4.07 $Y2=2.63
r269 39 40 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=4.07 $Y=2.755
+ $X2=4.07 $Y2=3.245
r270 35 133 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=3.245
+ $X2=1.74 $Y2=3.33
r271 35 37 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=1.74 $Y=3.245
+ $X2=1.74 $Y2=2.74
r272 31 130 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r273 31 33 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.73
r274 10 71 300 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=2 $X=12.555
+ $Y=1.84 $X2=12.69 $Y2=2.405
r275 9 67 300 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=2 $X=11.655
+ $Y=1.84 $X2=11.79 $Y2=2.335
r276 8 64 600 $w=1.7e-07 $l=1.07261e-06 $layer=licon1_PDIFF $count=1 $X=10.685
+ $Y=1.84 $X2=10.89 $Y2=2.815
r277 8 61 300 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=2 $X=10.685
+ $Y=1.84 $X2=10.89 $Y2=1.985
r278 7 55 300 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=2 $X=9.79
+ $Y=1.84 $X2=9.92 $Y2=1.985
r279 6 51 600 $w=1.7e-07 $l=3.33729e-07 $layer=licon1_PDIFF $count=1 $X=8.815
+ $Y=2.54 $X2=8.945 $Y2=2.815
r280 5 47 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=7.835
+ $Y=2.54 $X2=7.97 $Y2=2.815
r281 4 43 600 $w=1.7e-07 $l=4.92291e-07 $layer=licon1_PDIFF $count=1 $X=5.4
+ $Y=2.315 $X2=5.77 $Y2=2.6
r282 3 76 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=4.015
+ $Y=2.315 $X2=4.165 $Y2=2.59
r283 2 37 600 $w=1.7e-07 $l=9.65142e-07 $layer=licon1_PDIFF $count=1 $X=1.605
+ $Y=1.84 $X2=1.74 $Y2=2.74
r284 1 33 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=2.52 $X2=0.73 $Y2=2.73
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_4%Q 1 2 3 4 15 17 18 19 21 27 31 33 37 39 40
+ 41 52
c72 18 0 1.09277e-19 $X=11.01 $Y=1.065
c73 15 0 1.85451e-19 $X=10.845 $Y=0.515
r74 51 52 4.56667 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=12.24 $Y=1.985
+ $X2=12.125 $Y2=1.985
r75 41 51 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=12.72 $Y=1.985
+ $X2=12.24 $Y2=1.985
r76 41 45 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=12.72 $Y=1.985
+ $X2=12.72 $Y2=1.82
r77 40 45 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=12.72 $Y=1.665
+ $X2=12.72 $Y2=1.82
r78 39 40 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.72 $Y=1.295
+ $X2=12.72 $Y2=1.665
r79 38 39 7.2654 $w=2.28e-07 $l=1.45e-07 $layer=LI1_cond $X=12.72 $Y=1.15
+ $X2=12.72 $Y2=1.295
r80 34 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.345 $Y=1.065
+ $X2=12.18 $Y2=1.065
r81 33 38 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=12.605 $Y=1.065
+ $X2=12.72 $Y2=1.15
r82 33 34 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=12.605 $Y=1.065
+ $X2=12.345 $Y2=1.065
r83 29 51 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=12.24 $Y=2.15
+ $X2=12.24 $Y2=1.985
r84 29 31 11.775 $w=2.28e-07 $l=2.35e-07 $layer=LI1_cond $X=12.24 $Y=2.15
+ $X2=12.24 $Y2=2.385
r85 25 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.18 $Y=0.98
+ $X2=12.18 $Y2=1.065
r86 25 27 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=12.18 $Y=0.98
+ $X2=12.18 $Y2=0.515
r87 24 36 3.54079 $w=2.6e-07 $l=1.4e-07 $layer=LI1_cond $X=11.455 $Y=1.95
+ $X2=11.315 $Y2=1.95
r88 24 52 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=11.455 $Y=1.95
+ $X2=12.125 $Y2=1.95
r89 19 36 3.28787 $w=2.8e-07 $l=1.3e-07 $layer=LI1_cond $X=11.315 $Y=2.08
+ $X2=11.315 $Y2=1.95
r90 19 21 12.5534 $w=2.78e-07 $l=3.05e-07 $layer=LI1_cond $X=11.315 $Y=2.08
+ $X2=11.315 $Y2=2.385
r91 17 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.015 $Y=1.065
+ $X2=12.18 $Y2=1.065
r92 17 18 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=12.015 $Y=1.065
+ $X2=11.01 $Y2=1.065
r93 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.845 $Y=0.98
+ $X2=11.01 $Y2=1.065
r94 13 15 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=10.845 $Y=0.98
+ $X2=10.845 $Y2=0.515
r95 4 51 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=12.105
+ $Y=1.84 $X2=12.24 $Y2=1.985
r96 4 31 300 $w=1.7e-07 $l=6.08769e-07 $layer=licon1_PDIFF $count=2 $X=12.105
+ $Y=1.84 $X2=12.24 $Y2=2.385
r97 3 36 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=11.205
+ $Y=1.84 $X2=11.34 $Y2=1.985
r98 3 21 300 $w=1.7e-07 $l=6.08769e-07 $layer=licon1_PDIFF $count=2 $X=11.205
+ $Y=1.84 $X2=11.34 $Y2=2.385
r99 2 27 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=11.995
+ $Y=0.37 $X2=12.18 $Y2=0.515
r100 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.705
+ $Y=0.37 $X2=10.845 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_4%VGND 1 2 3 4 5 6 7 8 27 29 33 37 41 45 49 51
+ 53 56 57 58 60 65 84 89 94 100 103 106 110 119 121 124 130
c144 33 0 9.68091e-20 $X=1.7 $Y=0.495
r145 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r146 125 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r147 124 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r148 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r149 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r150 117 119 9.64943 $w=7.53e-07 $l=7e-08 $layer=LI1_cond $X=8.88 $Y=0.292
+ $X2=8.95 $Y2=0.292
r151 117 118 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r152 115 117 1.505 $w=7.53e-07 $l=9.5e-08 $layer=LI1_cond $X=8.785 $Y=0.292
+ $X2=8.88 $Y2=0.292
r153 113 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=8.88 $Y2=0
r154 112 115 6.09921 $w=7.53e-07 $l=3.85e-07 $layer=LI1_cond $X=8.4 $Y=0.292
+ $X2=8.785 $Y2=0.292
r155 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r156 109 112 4.75263 $w=7.53e-07 $l=3e-07 $layer=LI1_cond $X=8.1 $Y=0.292
+ $X2=8.4 $Y2=0.292
r157 109 110 11.1544 $w=7.53e-07 $l=1.65e-07 $layer=LI1_cond $X=8.1 $Y=0.292
+ $X2=7.935 $Y2=0.292
r158 106 107 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r159 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r160 101 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=1.68 $Y2=0
r161 100 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r162 98 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r163 98 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r164 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r165 95 124 13.2917 $w=1.7e-07 $l=3.33e-07 $layer=LI1_cond $X=11.845 $Y=0
+ $X2=11.512 $Y2=0
r166 95 97 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=11.845 $Y=0
+ $X2=12.24 $Y2=0
r167 94 129 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=12.515 $Y=0
+ $X2=12.737 $Y2=0
r168 94 97 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=12.515 $Y=0
+ $X2=12.24 $Y2=0
r169 93 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r170 93 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r171 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r172 90 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.51 $Y=0
+ $X2=10.345 $Y2=0
r173 90 92 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=10.51 $Y=0 $X2=10.8
+ $Y2=0
r174 89 124 13.2917 $w=1.7e-07 $l=3.32e-07 $layer=LI1_cond $X=11.18 $Y=0
+ $X2=11.512 $Y2=0
r175 89 92 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=11.18 $Y=0 $X2=10.8
+ $Y2=0
r176 88 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r177 88 118 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=8.88 $Y2=0
r178 87 119 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=9.84 $Y=0 $X2=8.95
+ $Y2=0
r179 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r180 84 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.18 $Y=0
+ $X2=10.345 $Y2=0
r181 84 87 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=10.18 $Y=0 $X2=9.84
+ $Y2=0
r182 83 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r183 82 110 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=7.92 $Y=0
+ $X2=7.935 $Y2=0
r184 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r185 79 82 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6 $Y=0 $X2=7.92
+ $Y2=0
r186 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r187 76 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r188 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r189 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r190 73 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=4.08 $Y2=0
r191 72 75 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r192 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r193 70 106 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=4.42 $Y=0
+ $X2=4.222 $Y2=0
r194 70 72 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=4.42 $Y=0 $X2=4.56
+ $Y2=0
r195 69 107 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=4.08 $Y2=0
r196 69 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r197 68 69 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r198 66 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.865 $Y=0
+ $X2=1.74 $Y2=0
r199 66 68 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.16
+ $Y2=0
r200 65 106 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=4.025 $Y=0
+ $X2=4.222 $Y2=0
r201 65 68 121.674 $w=1.68e-07 $l=1.865e-06 $layer=LI1_cond $X=4.025 $Y=0
+ $X2=2.16 $Y2=0
r202 63 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r203 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r204 60 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.67 $Y2=0
r205 60 62 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r206 58 83 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=7.92 $Y2=0
r207 58 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r208 57 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.835 $Y=0 $X2=6
+ $Y2=0
r209 56 75 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=5.67 $Y=0 $X2=5.52
+ $Y2=0
r210 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.67 $Y=0 $X2=5.835
+ $Y2=0
r211 51 129 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=12.68 $Y=0.085
+ $X2=12.737 $Y2=0
r212 51 53 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=12.68 $Y=0.085
+ $X2=12.68 $Y2=0.645
r213 47 124 2.7522 $w=6.65e-07 $l=8.5e-08 $layer=LI1_cond $X=11.512 $Y=0.085
+ $X2=11.512 $Y2=0
r214 47 49 9.89238 $w=6.63e-07 $l=5.5e-07 $layer=LI1_cond $X=11.512 $Y=0.085
+ $X2=11.512 $Y2=0.635
r215 43 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.345 $Y=0.085
+ $X2=10.345 $Y2=0
r216 43 45 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.345 $Y=0.085
+ $X2=10.345 $Y2=0.515
r217 39 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.835 $Y=0.085
+ $X2=5.835 $Y2=0
r218 39 41 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.835 $Y=0.085
+ $X2=5.835 $Y2=0.515
r219 35 106 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=4.222 $Y=0.085
+ $X2=4.222 $Y2=0
r220 35 37 12.5456 $w=3.93e-07 $l=4.3e-07 $layer=LI1_cond $X=4.222 $Y=0.085
+ $X2=4.222 $Y2=0.515
r221 31 103 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=0.085
+ $X2=1.74 $Y2=0
r222 31 33 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=1.74 $Y=0.085
+ $X2=1.74 $Y2=0.495
r223 30 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=0
+ $X2=0.67 $Y2=0
r224 29 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.615 $Y=0
+ $X2=1.74 $Y2=0
r225 29 30 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=1.615 $Y=0
+ $X2=0.795 $Y2=0
r226 25 100 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0
r227 25 27 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0.58
r228 8 53 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=12.47
+ $Y=0.37 $X2=12.68 $Y2=0.645
r229 7 49 91 $w=1.7e-07 $l=6.89891e-07 $layer=licon1_NDIFF $count=2 $X=11.135
+ $Y=0.37 $X2=11.705 $Y2=0.635
r230 6 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.205
+ $Y=0.37 $X2=10.345 $Y2=0.515
r231 5 115 121.333 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_NDIFF $count=1
+ $X=7.96 $Y=0.44 $X2=8.785 $Y2=0.585
r232 5 109 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1
+ $X=7.96 $Y=0.44 $X2=8.1 $Y2=0.585
r233 4 41 91 $w=1.7e-07 $l=3.05205e-07 $layer=licon1_NDIFF $count=2 $X=5.565
+ $Y=0.59 $X2=5.835 $Y2=0.515
r234 3 37 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=4.05
+ $Y=0.37 $X2=4.22 $Y2=0.515
r235 2 33 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.56
+ $Y=0.37 $X2=1.7 $Y2=0.495
r236 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.58
.ends


* File: sky130_fd_sc_ms__a22o_1.pxi.spice
* Created: Fri Aug 28 17:02:29 2020
* 
x_PM_SKY130_FD_SC_MS__A22O_1%A2 N_A2_c_60_n N_A2_M1005_g N_A2_M1001_g A2
+ N_A2_c_64_n PM_SKY130_FD_SC_MS__A22O_1%A2
x_PM_SKY130_FD_SC_MS__A22O_1%B2 N_B2_M1006_g N_B2_M1003_g B2 B2 N_B2_c_90_n
+ N_B2_c_91_n PM_SKY130_FD_SC_MS__A22O_1%B2
x_PM_SKY130_FD_SC_MS__A22O_1%B1 N_B1_M1000_g N_B1_M1004_g N_B1_c_126_n
+ N_B1_c_127_n B1 N_B1_c_129_n N_B1_c_130_n PM_SKY130_FD_SC_MS__A22O_1%B1
x_PM_SKY130_FD_SC_MS__A22O_1%A1 N_A1_c_167_n N_A1_M1007_g N_A1_c_168_n
+ N_A1_M1009_g A1 N_A1_c_169_n PM_SKY130_FD_SC_MS__A22O_1%A1
x_PM_SKY130_FD_SC_MS__A22O_1%A_225_392# N_A_225_392#_M1000_d
+ N_A_225_392#_M1006_d N_A_225_392#_M1002_g N_A_225_392#_M1008_g
+ N_A_225_392#_c_221_n N_A_225_392#_c_211_n N_A_225_392#_c_212_n
+ N_A_225_392#_c_217_n N_A_225_392#_c_213_n N_A_225_392#_c_214_n
+ PM_SKY130_FD_SC_MS__A22O_1%A_225_392#
x_PM_SKY130_FD_SC_MS__A22O_1%VPWR N_VPWR_M1005_s N_VPWR_M1009_d N_VPWR_c_275_n
+ N_VPWR_c_276_n N_VPWR_c_277_n VPWR N_VPWR_c_278_n N_VPWR_c_279_n
+ N_VPWR_c_274_n N_VPWR_c_281_n PM_SKY130_FD_SC_MS__A22O_1%VPWR
x_PM_SKY130_FD_SC_MS__A22O_1%A_135_392# N_A_135_392#_M1005_d
+ N_A_135_392#_M1004_d N_A_135_392#_c_311_n N_A_135_392#_c_309_n
+ N_A_135_392#_c_310_n N_A_135_392#_c_315_n
+ PM_SKY130_FD_SC_MS__A22O_1%A_135_392#
x_PM_SKY130_FD_SC_MS__A22O_1%X N_X_M1008_d N_X_M1002_d X X X X X X X
+ PM_SKY130_FD_SC_MS__A22O_1%X
x_PM_SKY130_FD_SC_MS__A22O_1%A_52_123# N_A_52_123#_M1001_s N_A_52_123#_M1007_d
+ N_A_52_123#_c_343_n N_A_52_123#_c_344_n N_A_52_123#_c_345_n
+ N_A_52_123#_c_346_n N_A_52_123#_c_347_n PM_SKY130_FD_SC_MS__A22O_1%A_52_123#
x_PM_SKY130_FD_SC_MS__A22O_1%VGND N_VGND_M1001_d N_VGND_M1008_s N_VGND_c_386_n
+ N_VGND_c_387_n N_VGND_c_388_n N_VGND_c_389_n VGND N_VGND_c_390_n
+ N_VGND_c_391_n N_VGND_c_392_n N_VGND_c_393_n PM_SKY130_FD_SC_MS__A22O_1%VGND
cc_1 VNB N_A2_c_60_n 0.0086683f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.42
cc_2 VNB N_A2_M1005_g 0.015328f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.46
cc_3 VNB N_A2_M1001_g 0.0113873f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.935
cc_4 VNB A2 0.0232559f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_5 VNB N_A2_c_64_n 0.0570677f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.34
cc_6 VNB N_B2_M1003_g 0.0316329f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.935
cc_7 VNB N_B2_c_90_n 0.0149356f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=0.34
cc_8 VNB N_B2_c_91_n 0.0183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B1_c_126_n 0.0137133f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_10 VNB N_B1_c_127_n 0.0133794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB B1 0.00283269f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=0.34
cc_12 VNB N_B1_c_129_n 0.0152763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B1_c_130_n 0.0120262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A1_c_167_n 0.0163683f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.42
cc_15 VNB N_A1_c_168_n 0.0588574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A1_c_169_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=0.34
cc_17 VNB N_A_225_392#_M1002_g 0.00169179f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.33
cc_18 VNB N_A_225_392#_M1008_g 0.0295424f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=0.34
cc_19 VNB N_A_225_392#_c_211_n 0.0190281f $X=-0.19 $Y=-0.245 $X2=0.342 $Y2=0.555
cc_20 VNB N_A_225_392#_c_212_n 0.00233602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_225_392#_c_213_n 0.00179529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_225_392#_c_214_n 0.0470336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_274_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB X 0.0565573f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.935
cc_25 VNB N_A_52_123#_c_343_n 0.00794929f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.935
cc_26 VNB N_A_52_123#_c_344_n 5.74149e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_27 VNB N_A_52_123#_c_345_n 0.00120814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_52_123#_c_346_n 0.00843668f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=0.34
cc_29 VNB N_A_52_123#_c_347_n 0.0209393f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.34
cc_30 VNB N_VGND_c_386_n 0.0106411f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.33
cc_31 VNB N_VGND_c_387_n 0.0161981f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=0.34
cc_32 VNB N_VGND_c_388_n 0.021055f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.34
cc_33 VNB N_VGND_c_389_n 0.00413177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_390_n 0.0408693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_391_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_392_n 0.221318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_393_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_A2_M1005_g 0.0350814f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=2.46
cc_39 VPB N_B2_M1006_g 0.021441f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=2.46
cc_40 VPB N_B2_c_90_n 0.0127759f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=0.34
cc_41 VPB N_B2_c_91_n 0.0163607f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_B1_M1004_g 0.0223968f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=0.935
cc_43 VPB B1 0.00222003f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=0.34
cc_44 VPB N_B1_c_129_n 0.0113568f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A1_c_168_n 0.0057612f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A1_M1009_g 0.0320693f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.33
cc_47 VPB N_A1_c_169_n 0.00217856f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=0.34
cc_48 VPB N_A_225_392#_M1002_g 0.0278634f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.33
cc_49 VPB N_A_225_392#_c_212_n 0.00156669f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_275_n 0.013204f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=0.935
cc_51 VPB N_VPWR_c_276_n 0.0494329f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.33
cc_52 VPB N_VPWR_c_277_n 0.0083905f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_278_n 0.0414344f $X=-0.19 $Y=1.66 $X2=0.342 $Y2=0.555
cc_54 VPB N_VPWR_c_279_n 0.0196299f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_274_n 0.0623191f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_281_n 0.0105477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_135_392#_c_309_n 0.0051056f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=0.34
cc_58 VPB N_A_135_392#_c_310_n 0.00160153f $X=-0.19 $Y=1.66 $X2=0.395 $Y2=0.34
cc_59 VPB X 0.0604727f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=0.935
cc_60 N_A2_M1005_g N_B2_M1006_g 0.0147971f $X=0.585 $Y=2.46 $X2=0 $Y2=0
cc_61 N_A2_c_64_n N_B2_M1003_g 0.0292353f $X=0.6 $Y=0.34 $X2=0 $Y2=0
cc_62 N_A2_M1005_g N_B2_c_90_n 0.0213587f $X=0.585 $Y=2.46 $X2=0 $Y2=0
cc_63 N_A2_M1005_g N_B2_c_91_n 0.0254147f $X=0.585 $Y=2.46 $X2=0 $Y2=0
cc_64 N_A2_M1005_g N_VPWR_c_276_n 0.00330306f $X=0.585 $Y=2.46 $X2=0 $Y2=0
cc_65 N_A2_M1005_g N_VPWR_c_278_n 0.00517089f $X=0.585 $Y=2.46 $X2=0 $Y2=0
cc_66 N_A2_M1005_g N_VPWR_c_274_n 0.00981577f $X=0.585 $Y=2.46 $X2=0 $Y2=0
cc_67 N_A2_M1005_g N_A_135_392#_c_311_n 0.012102f $X=0.585 $Y=2.46 $X2=0 $Y2=0
cc_68 N_A2_M1005_g N_A_135_392#_c_310_n 0.00358808f $X=0.585 $Y=2.46 $X2=0 $Y2=0
cc_69 A2 N_A_52_123#_M1001_s 0.00167987f $X=0.155 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_70 N_A2_M1001_g N_A_52_123#_c_343_n 0.011742f $X=0.6 $Y=0.935 $X2=0 $Y2=0
cc_71 A2 N_A_52_123#_c_343_n 2.3751e-19 $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_72 N_A2_M1001_g N_A_52_123#_c_344_n 5.89712e-19 $X=0.6 $Y=0.935 $X2=0 $Y2=0
cc_73 N_A2_c_60_n N_A_52_123#_c_347_n 9.56069e-19 $X=0.585 $Y=1.42 $X2=0 $Y2=0
cc_74 N_A2_M1001_g N_A_52_123#_c_347_n 0.00748439f $X=0.6 $Y=0.935 $X2=0 $Y2=0
cc_75 A2 N_A_52_123#_c_347_n 0.0179561f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_76 N_A2_c_64_n N_A_52_123#_c_347_n 0.00159699f $X=0.6 $Y=0.34 $X2=0 $Y2=0
cc_77 A2 N_VGND_c_386_n 0.0257619f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_78 N_A2_c_64_n N_VGND_c_386_n 0.00658794f $X=0.6 $Y=0.34 $X2=0 $Y2=0
cc_79 A2 N_VGND_c_388_n 0.0285096f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_80 N_A2_c_64_n N_VGND_c_388_n 0.010364f $X=0.6 $Y=0.34 $X2=0 $Y2=0
cc_81 A2 N_VGND_c_392_n 0.0151033f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_82 N_A2_c_64_n N_VGND_c_392_n 0.0170069f $X=0.6 $Y=0.34 $X2=0 $Y2=0
cc_83 N_B2_M1006_g N_B1_M1004_g 0.0227754f $X=1.035 $Y=2.46 $X2=0 $Y2=0
cc_84 N_B2_M1003_g N_B1_c_126_n 0.0600955f $X=1.075 $Y=0.715 $X2=0 $Y2=0
cc_85 N_B2_c_90_n B1 4.14342e-19 $X=1.05 $Y=1.635 $X2=0 $Y2=0
cc_86 N_B2_c_91_n B1 0.0223685f $X=1.05 $Y=1.635 $X2=0 $Y2=0
cc_87 N_B2_c_90_n N_B1_c_129_n 0.0214313f $X=1.05 $Y=1.635 $X2=0 $Y2=0
cc_88 N_B2_c_91_n N_B1_c_129_n 4.10923e-19 $X=1.05 $Y=1.635 $X2=0 $Y2=0
cc_89 N_B2_M1003_g N_B1_c_130_n 0.0103623f $X=1.075 $Y=0.715 $X2=0 $Y2=0
cc_90 N_B2_M1006_g N_A_225_392#_c_217_n 0.0103926f $X=1.035 $Y=2.46 $X2=0 $Y2=0
cc_91 N_B2_c_90_n N_A_225_392#_c_217_n 0.00202153f $X=1.05 $Y=1.635 $X2=0 $Y2=0
cc_92 N_B2_c_91_n N_A_225_392#_c_217_n 0.00722671f $X=1.05 $Y=1.635 $X2=0 $Y2=0
cc_93 N_B2_M1003_g N_A_225_392#_c_213_n 3.18622e-19 $X=1.075 $Y=0.715 $X2=0
+ $Y2=0
cc_94 N_B2_c_91_n N_VPWR_c_276_n 0.0212991f $X=1.05 $Y=1.635 $X2=0 $Y2=0
cc_95 N_B2_M1006_g N_VPWR_c_278_n 0.00333926f $X=1.035 $Y=2.46 $X2=0 $Y2=0
cc_96 N_B2_M1006_g N_VPWR_c_274_n 0.00423187f $X=1.035 $Y=2.46 $X2=0 $Y2=0
cc_97 N_B2_c_91_n N_A_135_392#_c_311_n 0.0183935f $X=1.05 $Y=1.635 $X2=0 $Y2=0
cc_98 N_B2_M1006_g N_A_135_392#_c_309_n 0.0141334f $X=1.035 $Y=2.46 $X2=0 $Y2=0
cc_99 N_B2_M1006_g N_A_135_392#_c_315_n 8.23621e-19 $X=1.035 $Y=2.46 $X2=0 $Y2=0
cc_100 N_B2_M1003_g N_A_52_123#_c_343_n 0.0126441f $X=1.075 $Y=0.715 $X2=0 $Y2=0
cc_101 N_B2_c_90_n N_A_52_123#_c_343_n 0.00430928f $X=1.05 $Y=1.635 $X2=0 $Y2=0
cc_102 N_B2_c_91_n N_A_52_123#_c_343_n 0.0506736f $X=1.05 $Y=1.635 $X2=0 $Y2=0
cc_103 N_B2_M1003_g N_A_52_123#_c_344_n 0.00951806f $X=1.075 $Y=0.715 $X2=0
+ $Y2=0
cc_104 N_B2_M1003_g N_A_52_123#_c_345_n 0.00535541f $X=1.075 $Y=0.715 $X2=0
+ $Y2=0
cc_105 N_B2_M1003_g N_A_52_123#_c_347_n 6.05736e-19 $X=1.075 $Y=0.715 $X2=0
+ $Y2=0
cc_106 N_B2_c_91_n N_A_52_123#_c_347_n 0.0278161f $X=1.05 $Y=1.635 $X2=0 $Y2=0
cc_107 N_B2_M1003_g N_VGND_c_386_n 0.00384771f $X=1.075 $Y=0.715 $X2=0 $Y2=0
cc_108 N_B2_M1003_g N_VGND_c_390_n 0.00522295f $X=1.075 $Y=0.715 $X2=0 $Y2=0
cc_109 N_B2_M1003_g N_VGND_c_392_n 0.00537853f $X=1.075 $Y=0.715 $X2=0 $Y2=0
cc_110 N_B1_c_126_n N_A1_c_167_n 0.0232104f $X=1.467 $Y=1.11 $X2=-0.19
+ $Y2=-0.245
cc_111 N_B1_c_127_n N_A1_c_168_n 0.00974511f $X=1.467 $Y=1.26 $X2=0 $Y2=0
cc_112 B1 N_A1_c_168_n 0.00230058f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_113 N_B1_c_129_n N_A1_c_168_n 0.020306f $X=1.59 $Y=1.635 $X2=0 $Y2=0
cc_114 N_B1_c_130_n N_A1_c_168_n 0.00726285f $X=1.59 $Y=1.47 $X2=0 $Y2=0
cc_115 N_B1_M1004_g N_A1_M1009_g 0.0219744f $X=1.515 $Y=2.46 $X2=0 $Y2=0
cc_116 B1 N_A1_c_169_n 0.0247613f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_117 N_B1_c_129_n N_A1_c_169_n 3.55055e-19 $X=1.59 $Y=1.635 $X2=0 $Y2=0
cc_118 N_B1_c_130_n N_A1_c_169_n 6.90997e-19 $X=1.59 $Y=1.47 $X2=0 $Y2=0
cc_119 N_B1_M1004_g N_A_225_392#_c_221_n 0.0153186f $X=1.515 $Y=2.46 $X2=0 $Y2=0
cc_120 B1 N_A_225_392#_c_221_n 0.0249441f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_121 N_B1_c_129_n N_A_225_392#_c_221_n 0.00323803f $X=1.59 $Y=1.635 $X2=0
+ $Y2=0
cc_122 N_B1_c_126_n N_A_225_392#_c_213_n 0.00452641f $X=1.467 $Y=1.11 $X2=0
+ $Y2=0
cc_123 N_B1_c_127_n N_A_225_392#_c_213_n 0.00482129f $X=1.467 $Y=1.26 $X2=0
+ $Y2=0
cc_124 B1 N_A_225_392#_c_213_n 0.0164626f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_125 N_B1_c_129_n N_A_225_392#_c_213_n 0.00392531f $X=1.59 $Y=1.635 $X2=0
+ $Y2=0
cc_126 N_B1_M1004_g N_VPWR_c_278_n 0.00333916f $X=1.515 $Y=2.46 $X2=0 $Y2=0
cc_127 N_B1_M1004_g N_VPWR_c_274_n 0.00423978f $X=1.515 $Y=2.46 $X2=0 $Y2=0
cc_128 N_B1_M1004_g N_A_135_392#_c_309_n 0.0149019f $X=1.515 $Y=2.46 $X2=0 $Y2=0
cc_129 N_B1_M1004_g N_A_135_392#_c_315_n 0.00741027f $X=1.515 $Y=2.46 $X2=0
+ $Y2=0
cc_130 N_B1_c_127_n N_A_52_123#_c_343_n 0.00280224f $X=1.467 $Y=1.26 $X2=0 $Y2=0
cc_131 N_B1_c_130_n N_A_52_123#_c_343_n 0.00113592f $X=1.59 $Y=1.47 $X2=0 $Y2=0
cc_132 N_B1_c_126_n N_A_52_123#_c_344_n 0.00585891f $X=1.467 $Y=1.11 $X2=0 $Y2=0
cc_133 N_B1_c_126_n N_A_52_123#_c_346_n 0.016242f $X=1.467 $Y=1.11 $X2=0 $Y2=0
cc_134 N_B1_c_126_n N_VGND_c_390_n 0.00399513f $X=1.467 $Y=1.11 $X2=0 $Y2=0
cc_135 N_B1_c_126_n N_VGND_c_392_n 0.00537853f $X=1.467 $Y=1.11 $X2=0 $Y2=0
cc_136 N_A1_c_168_n N_A_225_392#_M1002_g 0.00129392f $X=2.055 $Y=1.68 $X2=0
+ $Y2=0
cc_137 N_A1_M1009_g N_A_225_392#_M1002_g 0.0172894f $X=2.055 $Y=2.46 $X2=0 $Y2=0
cc_138 N_A1_c_169_n N_A_225_392#_M1002_g 3.32709e-19 $X=2.13 $Y=1.515 $X2=0
+ $Y2=0
cc_139 N_A1_c_168_n N_A_225_392#_M1008_g 0.00183582f $X=2.055 $Y=1.68 $X2=0
+ $Y2=0
cc_140 N_A1_c_168_n N_A_225_392#_c_221_n 6.94101e-19 $X=2.055 $Y=1.68 $X2=0
+ $Y2=0
cc_141 N_A1_M1009_g N_A_225_392#_c_221_n 0.0180088f $X=2.055 $Y=2.46 $X2=0 $Y2=0
cc_142 N_A1_c_169_n N_A_225_392#_c_221_n 0.0210878f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_143 N_A1_c_167_n N_A_225_392#_c_211_n 0.00648271f $X=1.865 $Y=1.11 $X2=0
+ $Y2=0
cc_144 N_A1_c_168_n N_A_225_392#_c_211_n 0.0153039f $X=2.055 $Y=1.68 $X2=0 $Y2=0
cc_145 N_A1_c_169_n N_A_225_392#_c_211_n 0.0247243f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_146 N_A1_c_168_n N_A_225_392#_c_212_n 0.00408954f $X=2.055 $Y=1.68 $X2=0
+ $Y2=0
cc_147 N_A1_M1009_g N_A_225_392#_c_212_n 0.00405738f $X=2.055 $Y=2.46 $X2=0
+ $Y2=0
cc_148 N_A1_c_169_n N_A_225_392#_c_212_n 0.0277121f $X=2.13 $Y=1.515 $X2=0 $Y2=0
cc_149 N_A1_c_167_n N_A_225_392#_c_213_n 0.0110654f $X=1.865 $Y=1.11 $X2=0 $Y2=0
cc_150 N_A1_c_168_n N_A_225_392#_c_213_n 0.00186216f $X=2.055 $Y=1.68 $X2=0
+ $Y2=0
cc_151 N_A1_c_168_n N_A_225_392#_c_214_n 0.0190434f $X=2.055 $Y=1.68 $X2=0 $Y2=0
cc_152 N_A1_c_169_n N_A_225_392#_c_214_n 0.00100886f $X=2.13 $Y=1.515 $X2=0
+ $Y2=0
cc_153 N_A1_M1009_g N_VPWR_c_277_n 0.00403102f $X=2.055 $Y=2.46 $X2=0 $Y2=0
cc_154 N_A1_M1009_g N_VPWR_c_278_n 0.00517089f $X=2.055 $Y=2.46 $X2=0 $Y2=0
cc_155 N_A1_M1009_g N_VPWR_c_274_n 0.00979911f $X=2.055 $Y=2.46 $X2=0 $Y2=0
cc_156 N_A1_M1009_g N_A_135_392#_c_309_n 0.00374867f $X=2.055 $Y=2.46 $X2=0
+ $Y2=0
cc_157 N_A1_M1009_g N_A_135_392#_c_315_n 0.00738125f $X=2.055 $Y=2.46 $X2=0
+ $Y2=0
cc_158 N_A1_c_167_n N_A_52_123#_c_346_n 0.01135f $X=1.865 $Y=1.11 $X2=0 $Y2=0
cc_159 N_A1_c_168_n N_A_52_123#_c_346_n 7.37405e-19 $X=2.055 $Y=1.68 $X2=0 $Y2=0
cc_160 N_A1_c_167_n N_VGND_c_387_n 0.00705117f $X=1.865 $Y=1.11 $X2=0 $Y2=0
cc_161 N_A1_c_167_n N_VGND_c_390_n 0.00399513f $X=1.865 $Y=1.11 $X2=0 $Y2=0
cc_162 N_A1_c_167_n N_VGND_c_392_n 0.00537853f $X=1.865 $Y=1.11 $X2=0 $Y2=0
cc_163 N_A_225_392#_c_221_n N_VPWR_M1009_d 0.0152819f $X=2.505 $Y=2.055 $X2=0
+ $Y2=0
cc_164 N_A_225_392#_c_212_n N_VPWR_M1009_d 0.00189894f $X=2.67 $Y=1.465 $X2=0
+ $Y2=0
cc_165 N_A_225_392#_M1002_g N_VPWR_c_277_n 0.0227873f $X=2.785 $Y=2.4 $X2=0
+ $Y2=0
cc_166 N_A_225_392#_c_221_n N_VPWR_c_277_n 0.0389741f $X=2.505 $Y=2.055 $X2=0
+ $Y2=0
cc_167 N_A_225_392#_c_214_n N_VPWR_c_277_n 4.83456e-19 $X=2.785 $Y=1.465 $X2=0
+ $Y2=0
cc_168 N_A_225_392#_M1002_g N_VPWR_c_279_n 0.00460063f $X=2.785 $Y=2.4 $X2=0
+ $Y2=0
cc_169 N_A_225_392#_M1002_g N_VPWR_c_274_n 0.00912516f $X=2.785 $Y=2.4 $X2=0
+ $Y2=0
cc_170 N_A_225_392#_c_221_n N_A_135_392#_M1004_d 0.00813118f $X=2.505 $Y=2.055
+ $X2=0 $Y2=0
cc_171 N_A_225_392#_M1006_d N_A_135_392#_c_309_n 0.00197722f $X=1.125 $Y=1.96
+ $X2=0 $Y2=0
cc_172 N_A_225_392#_c_217_n N_A_135_392#_c_309_n 0.0161861f $X=1.26 $Y=2.135
+ $X2=0 $Y2=0
cc_173 N_A_225_392#_c_221_n N_A_135_392#_c_315_n 0.0227906f $X=2.505 $Y=2.055
+ $X2=0 $Y2=0
cc_174 N_A_225_392#_c_217_n N_A_135_392#_c_315_n 0.0322329f $X=1.26 $Y=2.135
+ $X2=0 $Y2=0
cc_175 N_A_225_392#_M1008_g X 0.0214406f $X=2.875 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A_225_392#_c_211_n X 0.00962585f $X=2.505 $Y=1.095 $X2=0 $Y2=0
cc_177 N_A_225_392#_c_212_n X 0.0550462f $X=2.67 $Y=1.465 $X2=0 $Y2=0
cc_178 N_A_225_392#_c_214_n X 0.0172494f $X=2.785 $Y=1.465 $X2=0 $Y2=0
cc_179 N_A_225_392#_c_211_n N_A_52_123#_M1007_d 0.00358528f $X=2.505 $Y=1.095
+ $X2=0 $Y2=0
cc_180 N_A_225_392#_c_217_n N_A_52_123#_c_343_n 0.00236654f $X=1.26 $Y=2.135
+ $X2=0 $Y2=0
cc_181 N_A_225_392#_c_213_n N_A_52_123#_c_343_n 0.00373163f $X=1.65 $Y=0.885
+ $X2=0 $Y2=0
cc_182 N_A_225_392#_c_213_n N_A_52_123#_c_344_n 0.0218843f $X=1.65 $Y=0.885
+ $X2=0 $Y2=0
cc_183 N_A_225_392#_M1000_d N_A_52_123#_c_346_n 0.00177578f $X=1.51 $Y=0.395
+ $X2=0 $Y2=0
cc_184 N_A_225_392#_c_211_n N_A_52_123#_c_346_n 0.014733f $X=2.505 $Y=1.095
+ $X2=0 $Y2=0
cc_185 N_A_225_392#_c_213_n N_A_52_123#_c_346_n 0.0162725f $X=1.65 $Y=0.885
+ $X2=0 $Y2=0
cc_186 N_A_225_392#_c_211_n N_VGND_M1008_s 0.00345306f $X=2.505 $Y=1.095 $X2=0
+ $Y2=0
cc_187 N_A_225_392#_M1008_g N_VGND_c_387_n 0.00698798f $X=2.875 $Y=0.74 $X2=0
+ $Y2=0
cc_188 N_A_225_392#_c_211_n N_VGND_c_387_n 0.0222869f $X=2.505 $Y=1.095 $X2=0
+ $Y2=0
cc_189 N_A_225_392#_c_214_n N_VGND_c_387_n 9.99596e-19 $X=2.785 $Y=1.465 $X2=0
+ $Y2=0
cc_190 N_A_225_392#_M1008_g N_VGND_c_391_n 0.00434272f $X=2.875 $Y=0.74 $X2=0
+ $Y2=0
cc_191 N_A_225_392#_M1008_g N_VGND_c_392_n 0.00828906f $X=2.875 $Y=0.74 $X2=0
+ $Y2=0
cc_192 N_VPWR_c_277_n N_A_135_392#_c_309_n 0.01232f $X=2.56 $Y=2.43 $X2=0 $Y2=0
cc_193 N_VPWR_c_278_n N_A_135_392#_c_309_n 0.07252f $X=2.165 $Y=3.33 $X2=0 $Y2=0
cc_194 N_VPWR_c_274_n N_A_135_392#_c_309_n 0.0400816f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_195 N_VPWR_c_276_n N_A_135_392#_c_310_n 0.0103534f $X=0.36 $Y=2.135 $X2=0
+ $Y2=0
cc_196 N_VPWR_c_278_n N_A_135_392#_c_310_n 0.0178163f $X=2.165 $Y=3.33 $X2=0
+ $Y2=0
cc_197 N_VPWR_c_274_n N_A_135_392#_c_310_n 0.00958215f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_198 N_VPWR_c_277_n X 0.0246374f $X=2.56 $Y=2.43 $X2=0 $Y2=0
cc_199 N_VPWR_c_279_n X 0.0146357f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_200 N_VPWR_c_274_n X 0.0121141f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_201 X N_VGND_c_387_n 0.0182902f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_202 X N_VGND_c_391_n 0.0145639f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_203 X N_VGND_c_392_n 0.0119984f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_204 N_A_52_123#_c_343_n N_VGND_M1001_d 0.00205163f $X=1.115 $Y=1.215
+ $X2=-0.19 $Y2=-0.245
cc_205 N_A_52_123#_c_343_n N_VGND_c_386_n 0.0172284f $X=1.115 $Y=1.215 $X2=0
+ $Y2=0
cc_206 N_A_52_123#_c_345_n N_VGND_c_386_n 0.011275f $X=1.285 $Y=0.5 $X2=0 $Y2=0
cc_207 N_A_52_123#_c_346_n N_VGND_c_387_n 0.0164198f $X=2.08 $Y=0.54 $X2=0 $Y2=0
cc_208 N_A_52_123#_c_345_n N_VGND_c_390_n 0.00679203f $X=1.285 $Y=0.5 $X2=0
+ $Y2=0
cc_209 N_A_52_123#_c_346_n N_VGND_c_390_n 0.0353785f $X=2.08 $Y=0.54 $X2=0 $Y2=0
cc_210 N_A_52_123#_c_345_n N_VGND_c_392_n 0.00615299f $X=1.285 $Y=0.5 $X2=0
+ $Y2=0
cc_211 N_A_52_123#_c_346_n N_VGND_c_392_n 0.033495f $X=2.08 $Y=0.54 $X2=0 $Y2=0
cc_212 N_A_52_123#_c_344_n A_230_79# 0.00395173f $X=1.2 $Y=1.13 $X2=-0.19
+ $Y2=-0.245
cc_213 N_A_52_123#_c_346_n A_230_79# 6.79616e-19 $X=2.08 $Y=0.54 $X2=-0.19
+ $Y2=-0.245

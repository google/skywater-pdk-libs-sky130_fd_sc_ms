* File: sky130_fd_sc_ms__dfxtp_2.pex.spice
* Created: Fri Aug 28 17:25:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DFXTP_2%CLK 3 7 9 13 16
r35 15 16 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.465
+ $X2=0.505 $Y2=1.465
r36 12 15 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=0.34 $Y=1.465
+ $X2=0.495 $Y2=1.465
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.34
+ $Y=1.465 $X2=0.34 $Y2=1.465
r38 9 13 6.06549 $w=3.78e-07 $l=2e-07 $layer=LI1_cond $X=0.315 $Y=1.665
+ $X2=0.315 $Y2=1.465
r39 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.465
r40 5 7 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.74
r41 1 16 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=1.465
r42 1 3 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_2%A_27_74# 1 2 9 13 16 20 24 26 27 31 34 36 38
+ 40 41 42 45 48 49 51 52 53 55 56 57 59 61 63 64 67 69 72 73 76 86 90 91 92 95
+ 98
c263 98 0 6.76432e-20 $X=3.145 $Y=1.92
c264 90 0 6.36416e-20 $X=5.725 $Y=0.345
c265 88 0 2.82287e-20 $X=3.67 $Y=0.775
c266 61 0 1.41143e-20 $X=3.67 $Y=0.69
c267 16 0 5.64678e-20 $X=2.99 $Y=0.805
c268 9 0 8.25497e-20 $X=0.955 $Y=2.4
r269 91 102 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.725 $Y=0.345
+ $X2=5.725 $Y2=0.51
r270 90 92 8.74048 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=5.725 $Y=0.382
+ $X2=5.56 $Y2=0.382
r271 90 91 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.725
+ $Y=0.345 $X2=5.725 $Y2=0.345
r272 84 86 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.455 $Y=1.37
+ $X2=3.67 $Y2=1.37
r273 80 98 27.1549 $w=2.84e-07 $l=1.6e-07 $layer=POLY_cond $X=3.305 $Y=1.92
+ $X2=3.145 $Y2=1.92
r274 79 80 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.305
+ $Y=1.92 $X2=3.305 $Y2=1.92
r275 76 96 40.8147 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.982 $Y=1.385
+ $X2=0.982 $Y2=1.55
r276 76 95 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.982 $Y=1.385
+ $X2=0.982 $Y2=1.22
r277 75 77 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=1.385
+ $X2=0.905 $Y2=1.55
r278 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.97
+ $Y=1.385 $X2=0.97 $Y2=1.385
r279 72 75 8.84058 $w=4.58e-07 $l=3.4e-07 $layer=LI1_cond $X=0.905 $Y=1.045
+ $X2=0.905 $Y2=1.385
r280 72 73 7.19996 $w=4.58e-07 $l=8.5e-08 $layer=LI1_cond $X=0.905 $Y=1.045
+ $X2=0.905 $Y2=0.96
r281 69 92 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=4.575 $Y=0.34
+ $X2=5.56 $Y2=0.34
r282 66 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.49 $Y=0.425
+ $X2=4.575 $Y2=0.34
r283 66 67 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.49 $Y=0.425
+ $X2=4.49 $Y2=0.69
r284 65 88 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.755 $Y=0.775
+ $X2=3.67 $Y2=0.775
r285 64 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.405 $Y=0.775
+ $X2=4.49 $Y2=0.69
r286 64 65 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.405 $Y=0.775
+ $X2=3.755 $Y2=0.775
r287 63 86 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=1.285
+ $X2=3.67 $Y2=1.37
r288 62 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=0.86
+ $X2=3.67 $Y2=0.775
r289 62 63 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.67 $Y=0.86
+ $X2=3.67 $Y2=1.285
r290 61 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=0.69
+ $X2=3.67 $Y2=0.775
r291 60 61 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.67 $Y=0.425
+ $X2=3.67 $Y2=0.69
r292 59 79 6.77908 $w=2.53e-07 $l=1.5e-07 $layer=LI1_cond $X=3.455 $Y=1.957
+ $X2=3.305 $Y2=1.957
r293 58 84 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.455 $Y=1.455
+ $X2=3.455 $Y2=1.37
r294 58 59 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.455 $Y=1.455
+ $X2=3.455 $Y2=1.83
r295 56 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.585 $Y=0.34
+ $X2=3.67 $Y2=0.425
r296 56 57 69.4813 $w=1.68e-07 $l=1.065e-06 $layer=LI1_cond $X=3.585 $Y=0.34
+ $X2=2.52 $Y2=0.34
r297 54 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.435 $Y=0.425
+ $X2=2.52 $Y2=0.34
r298 54 55 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.435 $Y=0.425
+ $X2=2.435 $Y2=0.81
r299 52 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.35 $Y=0.895
+ $X2=2.435 $Y2=0.81
r300 52 53 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.35 $Y=0.895
+ $X2=1.815 $Y2=0.895
r301 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.73 $Y=0.81
+ $X2=1.815 $Y2=0.895
r302 50 51 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.73 $Y=0.425
+ $X2=1.73 $Y2=0.81
r303 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.645 $Y=0.34
+ $X2=1.73 $Y2=0.425
r304 48 49 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.645 $Y=0.34
+ $X2=1.135 $Y2=0.34
r305 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.05 $Y=0.425
+ $X2=1.135 $Y2=0.34
r306 46 73 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=1.05 $Y=0.425
+ $X2=1.05 $Y2=0.96
r307 45 77 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=0.76 $Y=1.95 $X2=0.76
+ $Y2=1.55
r308 43 71 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.035
+ $X2=0.28 $Y2=2.035
r309 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.675 $Y=2.035
+ $X2=0.76 $Y2=1.95
r310 42 43 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.675 $Y=2.035
+ $X2=0.445 $Y2=2.035
r311 40 72 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.675 $Y=1.045
+ $X2=0.905 $Y2=1.045
r312 40 41 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.675 $Y=1.045
+ $X2=0.365 $Y2=1.045
r313 36 71 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.12 $X2=0.28
+ $Y2=2.035
r314 36 38 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.28 $Y=2.12
+ $X2=0.28 $Y2=2.815
r315 32 41 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.96
+ $X2=0.365 $Y2=1.045
r316 32 34 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.24 $Y=0.96
+ $X2=0.24 $Y2=0.515
r317 31 102 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.785 $Y=0.83
+ $X2=5.785 $Y2=0.51
r318 29 31 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=5.785 $Y=1.69
+ $X2=5.785 $Y2=0.83
r319 26 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.71 $Y=1.765
+ $X2=5.785 $Y2=1.69
r320 26 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.71 $Y=1.765 $X2=5.11
+ $Y2=1.765
r321 22 27 33.7919 $w=1.32e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.02 $Y=1.84
+ $X2=5.11 $Y2=1.765
r322 22 24 272.097 $w=1.8e-07 $l=7e-07 $layer=POLY_cond $X=5.02 $Y=1.84 $X2=5.02
+ $Y2=2.54
r323 18 98 13.4541 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.145 $Y=2.085
+ $X2=3.145 $Y2=1.92
r324 18 20 250.718 $w=1.8e-07 $l=6.45e-07 $layer=POLY_cond $X=3.145 $Y=2.085
+ $X2=3.145 $Y2=2.73
r325 14 98 26.3063 $w=2.84e-07 $l=2.29783e-07 $layer=POLY_cond $X=2.99 $Y=1.755
+ $X2=3.145 $Y2=1.92
r326 14 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.99 $Y=1.755
+ $X2=2.99 $Y2=0.805
r327 13 95 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.085 $Y=0.74
+ $X2=1.085 $Y2=1.22
r328 9 96 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.955 $Y=2.4
+ $X2=0.955 $Y2=1.55
r329 2 71 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r330 2 38 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r331 1 34 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_2%D 3 5 9 14 16 18 22 24
c62 24 0 1.22251e-19 $X=2.165 $Y=1.225
c63 18 0 5.64678e-20 $X=2.16 $Y=1.295
c64 14 0 2.06364e-19 $X=1.89 $Y=2.215
c65 5 0 1.77322e-19 $X=2.485 $Y=1.225
r66 24 27 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.165 $Y=1.225
+ $X2=2.165 $Y2=1.315
r67 18 30 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.16 $Y=1.315
+ $X2=1.97 $Y2=1.315
r68 18 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.165
+ $Y=1.315 $X2=2.165 $Y2=1.315
r69 15 22 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=1.89 $Y=2.215
+ $X2=2.08 $Y2=2.215
r70 14 16 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.89 $Y=2.215
+ $X2=1.89 $Y2=2.05
r71 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.89
+ $Y=2.215 $X2=1.89 $Y2=2.215
r72 11 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.97 $Y=1.48
+ $X2=1.97 $Y2=1.315
r73 11 16 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.97 $Y=1.48
+ $X2=1.97 $Y2=2.05
r74 7 9 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=2.56 $Y=1.15 $X2=2.56
+ $Y2=0.805
r75 6 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.33 $Y=1.225
+ $X2=2.165 $Y2=1.225
r76 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.485 $Y=1.225
+ $X2=2.56 $Y2=1.15
r77 5 6 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=2.485 $Y=1.225
+ $X2=2.33 $Y2=1.225
r78 1 22 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.08 $Y=2.38
+ $X2=2.08 $Y2=2.215
r79 1 3 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=2.08 $Y=2.38 $X2=2.08
+ $Y2=2.75
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_2%A_209_368# 1 2 9 10 11 15 19 23 27 30 32 35
+ 37 39 41 43 44 45 49 50 53 56 59 63 70 71 75
c223 70 0 4.0193e-19 $X=5.25 $Y=1.315
c224 53 0 1.22251e-19 $X=1.39 $Y=1.65
c225 50 0 1.43814e-19 $X=5.71 $Y=2.215
c226 15 0 1.23815e-19 $X=2.615 $Y=2.355
r227 71 72 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.905 $Y=2.71
+ $X2=4.905 $Y2=2.99
r228 70 78 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=5.25 $Y=1.315
+ $X2=5.125 $Y2=1.315
r229 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.25
+ $Y=1.315 $X2=5.25 $Y2=1.315
r230 63 65 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.455 $Y=2.71
+ $X2=3.455 $Y2=2.84
r231 59 61 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.19 $Y=2.71
+ $X2=2.19 $Y2=2.84
r232 56 76 40.0724 $w=3.6e-07 $l=2.5e-07 $layer=POLY_cond $X=1.58 $Y=1.515
+ $X2=1.58 $Y2=1.765
r233 56 75 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.58 $Y=1.515
+ $X2=1.58 $Y2=1.35
r234 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.565
+ $Y=1.515 $X2=1.565 $Y2=1.515
r235 53 55 5.81744 $w=3.67e-07 $l=1.75e-07 $layer=LI1_cond $X=1.39 $Y=1.65
+ $X2=1.565 $Y2=1.65
r236 50 82 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=5.71 $Y=2.215
+ $X2=5.55 $Y2=2.215
r237 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.71
+ $Y=2.215 $X2=5.71 $Y2=2.215
r238 47 49 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=5.71 $Y=2.905
+ $X2=5.71 $Y2=2.215
r239 46 72 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.99 $Y=2.99
+ $X2=4.905 $Y2=2.99
r240 45 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.545 $Y=2.99
+ $X2=5.71 $Y2=2.905
r241 45 46 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=5.545 $Y=2.99
+ $X2=4.99 $Y2=2.99
r242 44 71 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.905 $Y=2.625
+ $X2=4.905 $Y2=2.71
r243 43 69 14.4144 $w=2.92e-07 $l=4.31625e-07 $layer=LI1_cond $X=4.905 $Y=1.54
+ $X2=5.25 $Y2=1.345
r244 43 44 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=4.905 $Y=1.54
+ $X2=4.905 $Y2=2.625
r245 42 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=2.71
+ $X2=3.455 $Y2=2.71
r246 41 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.82 $Y=2.71
+ $X2=4.905 $Y2=2.71
r247 41 42 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=4.82 $Y=2.71
+ $X2=3.54 $Y2=2.71
r248 40 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=2.84
+ $X2=2.19 $Y2=2.84
r249 39 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.37 $Y=2.84
+ $X2=3.455 $Y2=2.84
r250 39 40 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=3.37 $Y=2.84
+ $X2=2.275 $Y2=2.84
r251 38 58 5.73712 $w=1.7e-07 $l=2.7214e-07 $layer=LI1_cond $X=1.475 $Y=2.71
+ $X2=1.245 $Y2=2.802
r252 37 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=2.71
+ $X2=2.19 $Y2=2.71
r253 37 38 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.105 $Y=2.71
+ $X2=1.475 $Y2=2.71
r254 33 53 5.25812 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=1.39 $Y=1.35 $X2=1.39
+ $Y2=1.65
r255 33 35 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.39 $Y=1.35
+ $X2=1.39 $Y2=0.86
r256 30 58 3.15363 $w=4.6e-07 $l=1.77e-07 $layer=LI1_cond $X=1.245 $Y=2.625
+ $X2=1.245 $Y2=2.802
r257 30 32 16.6411 $w=4.58e-07 $l=6.4e-07 $layer=LI1_cond $X=1.245 $Y=2.625
+ $X2=1.245 $Y2=1.985
r258 29 53 4.82016 $w=3.67e-07 $l=3.65377e-07 $layer=LI1_cond $X=1.245 $Y=1.95
+ $X2=1.39 $Y2=1.65
r259 29 32 0.91006 $w=4.58e-07 $l=3.5e-08 $layer=LI1_cond $X=1.245 $Y=1.95
+ $X2=1.245 $Y2=1.985
r260 25 82 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.55 $Y=2.38
+ $X2=5.55 $Y2=2.215
r261 25 27 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=5.55 $Y=2.38
+ $X2=5.55 $Y2=2.75
r262 21 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.125 $Y=1.15
+ $X2=5.125 $Y2=1.315
r263 21 23 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=5.125 $Y=1.15
+ $X2=5.125 $Y2=0.65
r264 17 19 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=3.465 $Y=0.255
+ $X2=3.465 $Y2=0.715
r265 13 15 200.185 $w=1.8e-07 $l=5.15e-07 $layer=POLY_cond $X=2.615 $Y=1.84
+ $X2=2.615 $Y2=2.355
r266 12 76 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.76 $Y=1.765
+ $X2=1.58 $Y2=1.765
r267 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.525 $Y=1.765
+ $X2=2.615 $Y2=1.84
r268 11 12 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=2.525 $Y=1.765
+ $X2=1.76 $Y2=1.765
r269 9 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.39 $Y=0.18
+ $X2=3.465 $Y2=0.255
r270 9 10 835.809 $w=1.5e-07 $l=1.63e-06 $layer=POLY_cond $X=3.39 $Y=0.18
+ $X2=1.76 $Y2=0.18
r271 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.685 $Y=0.255
+ $X2=1.76 $Y2=0.18
r272 7 75 561.479 $w=1.5e-07 $l=1.095e-06 $layer=POLY_cond $X=1.685 $Y=0.255
+ $X2=1.685 $Y2=1.35
r273 2 58 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.815
r274 2 32 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=1.985
r275 1 35 182 $w=1.7e-07 $l=5.9397e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.37 $X2=1.39 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_2%A_695_459# 1 2 7 9 11 14 18 20 25 26 30 36
c85 26 0 1.31176e-19 $X=4.565 $Y=2.125
c86 14 0 1.80864e-19 $X=3.855 $Y=0.715
c87 11 0 5.9515e-20 $X=3.755 $Y=2.295
r88 28 30 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.475 $Y=2.29
+ $X2=4.565 $Y2=2.29
r89 26 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.565 $Y=2.125
+ $X2=4.565 $Y2=2.29
r90 25 26 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.565 $Y=1.415
+ $X2=4.565 $Y2=2.125
r91 23 36 38.0101 $w=2.98e-07 $l=2.35e-07 $layer=POLY_cond $X=4.09 $Y=1.25
+ $X2=3.855 $Y2=1.25
r92 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.09
+ $Y=1.25 $X2=4.09 $Y2=1.25
r93 20 25 10.1681 $w=2.93e-07 $l=2.31633e-07 $layer=LI1_cond $X=4.48 $Y=1.222
+ $X2=4.565 $Y2=1.415
r94 20 33 18.8205 $w=2.93e-07 $l=5.81849e-07 $layer=LI1_cond $X=4.48 $Y=1.222
+ $X2=4.777 $Y2=0.77
r95 20 22 11.6741 $w=3.83e-07 $l=3.9e-07 $layer=LI1_cond $X=4.48 $Y=1.222
+ $X2=4.09 $Y2=1.222
r96 12 36 18.8112 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.855 $Y=1.085
+ $X2=3.855 $Y2=1.25
r97 12 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.855 $Y=1.085
+ $X2=3.855 $Y2=0.715
r98 11 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.755 $Y=2.295
+ $X2=3.755 $Y2=2.37
r99 10 36 16.1745 $w=2.98e-07 $l=2.09105e-07 $layer=POLY_cond $X=3.755 $Y=1.415
+ $X2=3.855 $Y2=1.25
r100 10 11 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=3.755 $Y=1.415
+ $X2=3.755 $Y2=2.295
r101 7 18 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.565 $Y=2.37
+ $X2=3.755 $Y2=2.37
r102 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.565 $Y=2.445
+ $X2=3.565 $Y2=2.73
r103 2 28 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=4.335
+ $Y=2.12 $X2=4.475 $Y2=2.29
r104 1 33 182 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_NDIFF $count=1 $X=4.77
+ $Y=0.375 $X2=4.91 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_2%A_541_429# 1 2 9 12 13 15 18 22 25 27 28 29
+ 35 40 45 51
c102 40 0 1.80864e-19 $X=3.225 $Y=0.78
c103 25 0 2.36837e-19 $X=3.115 $Y=1.49
r104 50 51 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=4.245 $Y=1.79
+ $X2=4.57 $Y2=1.79
r105 46 50 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=4.205 $Y=1.79
+ $X2=4.245 $Y2=1.79
r106 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.205
+ $Y=1.79 $X2=4.205 $Y2=1.79
r107 42 45 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=4.05 $Y=1.79
+ $X2=4.205 $Y2=1.79
r108 37 40 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.115 $Y=0.78
+ $X2=3.225 $Y2=0.78
r109 33 35 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.87 $Y=1.575
+ $X2=3.115 $Y2=1.575
r110 28 31 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=2.855 $Y=2.34
+ $X2=2.855 $Y2=2.355
r111 28 29 12.2041 $w=1.98e-07 $l=2.15e-07 $layer=LI1_cond $X=2.855 $Y=2.34
+ $X2=2.855 $Y2=2.125
r112 26 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.05 $Y=1.955
+ $X2=4.05 $Y2=1.79
r113 26 27 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.05 $Y=1.955
+ $X2=4.05 $Y2=2.255
r114 25 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=1.49
+ $X2=3.115 $Y2=1.575
r115 24 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.115 $Y=0.945
+ $X2=3.115 $Y2=0.78
r116 24 25 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=3.115 $Y=0.945
+ $X2=3.115 $Y2=1.49
r117 23 28 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.955 $Y=2.34
+ $X2=2.855 $Y2=2.34
r118 22 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.965 $Y=2.34
+ $X2=4.05 $Y2=2.255
r119 22 23 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.965 $Y=2.34
+ $X2=2.955 $Y2=2.34
r120 20 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=1.66
+ $X2=2.87 $Y2=1.575
r121 20 29 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.87 $Y=1.66
+ $X2=2.87 $Y2=2.125
r122 16 18 64.0957 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=4.57 $Y=1.075
+ $X2=4.695 $Y2=1.075
r123 13 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.695 $Y=1
+ $X2=4.695 $Y2=1.075
r124 13 15 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.695 $Y=1
+ $X2=4.695 $Y2=0.65
r125 12 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.57 $Y=1.625
+ $X2=4.57 $Y2=1.79
r126 11 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.57 $Y=1.15
+ $X2=4.57 $Y2=1.075
r127 11 12 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=4.57 $Y=1.15
+ $X2=4.57 $Y2=1.625
r128 7 50 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.245 $Y=1.955
+ $X2=4.245 $Y2=1.79
r129 7 9 227.395 $w=1.8e-07 $l=5.85e-07 $layer=POLY_cond $X=4.245 $Y=1.955
+ $X2=4.245 $Y2=2.54
r130 2 31 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=2.705
+ $Y=2.145 $X2=2.84 $Y2=2.355
r131 1 40 182 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.595 $X2=3.225 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_2%A_1217_314# 1 2 9 13 17 21 23 25 28 32 33 36
+ 40 44 48 50 51 55 56 57 59 61 68
c133 68 0 1.78913e-19 $X=8.135 $Y=1.56
c134 56 0 2.92783e-19 $X=6.25 $Y=1.735
c135 13 0 6.36416e-20 $X=6.175 $Y=0.83
r136 68 69 1.38109 $w=3.49e-07 $l=1e-08 $layer=POLY_cond $X=8.135 $Y=1.56
+ $X2=8.145 $Y2=1.56
r137 67 68 58.0057 $w=3.49e-07 $l=4.2e-07 $layer=POLY_cond $X=7.715 $Y=1.56
+ $X2=8.135 $Y2=1.56
r138 59 62 8.8128 $w=3.38e-07 $l=2.6e-07 $layer=LI1_cond $X=7.595 $Y=1.515
+ $X2=7.595 $Y2=1.775
r139 59 61 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=7.595 $Y=1.515
+ $X2=7.595 $Y2=1.35
r140 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.645
+ $Y=1.515 $X2=7.645 $Y2=1.515
r141 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.25
+ $Y=1.735 $X2=6.25 $Y2=1.735
r142 52 61 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.51 $Y=1.02
+ $X2=7.51 $Y2=1.35
r143 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.425 $Y=0.935
+ $X2=7.51 $Y2=1.02
r144 50 51 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=7.425 $Y=0.935
+ $X2=7.115 $Y2=0.935
r145 49 57 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.04 $Y=1.775
+ $X2=6.915 $Y2=1.775
r146 48 62 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=7.425 $Y=1.775
+ $X2=7.595 $Y2=1.775
r147 48 49 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=7.425 $Y=1.775
+ $X2=7.04 $Y2=1.775
r148 44 46 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=6.915 $Y=1.985
+ $X2=6.915 $Y2=2.695
r149 42 57 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.915 $Y=1.86
+ $X2=6.915 $Y2=1.775
r150 42 44 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.915 $Y=1.86
+ $X2=6.915 $Y2=1.985
r151 38 51 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.95 $Y=0.85
+ $X2=7.115 $Y2=0.935
r152 38 40 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=6.95 $Y=0.85
+ $X2=6.95 $Y2=0.645
r153 37 55 4.72267 $w=1.7e-07 $l=1.92678e-07 $layer=LI1_cond $X=6.415 $Y=1.775
+ $X2=6.25 $Y2=1.715
r154 36 57 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.79 $Y=1.775
+ $X2=6.915 $Y2=1.775
r155 36 37 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.79 $Y=1.775
+ $X2=6.415 $Y2=1.775
r156 32 56 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.25 $Y=2.075
+ $X2=6.25 $Y2=1.735
r157 32 33 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.25 $Y=2.075
+ $X2=6.25 $Y2=2.24
r158 31 56 43.7316 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.25 $Y=1.57
+ $X2=6.25 $Y2=1.735
r159 26 69 22.56 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=8.145 $Y=1.35
+ $X2=8.145 $Y2=1.56
r160 26 28 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.145 $Y=1.35
+ $X2=8.145 $Y2=0.74
r161 23 68 18.24 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=8.135 $Y=1.77
+ $X2=8.135 $Y2=1.56
r162 23 25 168.7 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=8.135 $Y=1.77
+ $X2=8.135 $Y2=2.4
r163 19 67 22.56 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.715 $Y=1.35
+ $X2=7.715 $Y2=1.56
r164 19 21 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.715 $Y=1.35
+ $X2=7.715 $Y2=0.74
r165 15 67 4.14327 $w=3.49e-07 $l=3e-08 $layer=POLY_cond $X=7.685 $Y=1.56
+ $X2=7.715 $Y2=1.56
r166 15 60 5.52436 $w=3.49e-07 $l=4e-08 $layer=POLY_cond $X=7.685 $Y=1.56
+ $X2=7.645 $Y2=1.56
r167 15 17 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.685 $Y=1.68
+ $X2=7.685 $Y2=2.4
r168 13 31 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.175 $Y=0.83
+ $X2=6.175 $Y2=1.57
r169 9 33 198.242 $w=1.8e-07 $l=5.1e-07 $layer=POLY_cond $X=6.175 $Y=2.75
+ $X2=6.175 $Y2=2.24
r170 2 46 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.81
+ $Y=1.84 $X2=6.955 $Y2=2.695
r171 2 44 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=6.81
+ $Y=1.84 $X2=6.955 $Y2=1.985
r172 1 40 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=6.805
+ $Y=0.37 $X2=6.95 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_2%A_1022_424# 1 2 9 13 17 19 23 24 26 28 31 33
+ 34 35
c102 35 0 1.43814e-19 $X=6.91 $Y=1.355
c103 33 0 1.78913e-19 $X=7.075 $Y=1.355
c104 28 0 1.52685e-19 $X=5.67 $Y=1.71
c105 24 0 1.79753e-19 $X=5.33 $Y=1.795
c106 23 0 2.31098e-19 $X=5.585 $Y=1.795
c107 9 0 2.55617e-20 $X=7.165 $Y=0.645
r108 34 39 40.8642 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=7.09 $Y=1.355
+ $X2=7.09 $Y2=1.52
r109 34 38 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=7.09 $Y=1.355
+ $X2=7.09 $Y2=1.19
r110 33 35 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.075 $Y=1.355
+ $X2=6.91 $Y2=1.355
r111 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.075
+ $Y=1.355 $X2=7.075 $Y2=1.355
r112 30 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.755 $Y=1.315
+ $X2=5.67 $Y2=1.315
r113 30 35 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=5.755 $Y=1.315
+ $X2=6.91 $Y2=1.315
r114 27 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.67 $Y=1.4 $X2=5.67
+ $Y2=1.315
r115 27 28 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.67 $Y=1.4
+ $X2=5.67 $Y2=1.71
r116 26 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.67 $Y=1.23
+ $X2=5.67 $Y2=1.315
r117 25 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.67 $Y=0.945
+ $X2=5.67 $Y2=1.23
r118 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.585 $Y=1.795
+ $X2=5.67 $Y2=1.71
r119 23 24 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.585 $Y=1.795
+ $X2=5.33 $Y2=1.795
r120 19 25 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.585 $Y=0.82
+ $X2=5.67 $Y2=0.945
r121 19 21 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=5.585 $Y=0.82
+ $X2=5.49 $Y2=0.82
r122 15 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.245 $Y=1.88
+ $X2=5.33 $Y2=1.795
r123 15 17 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=5.245 $Y=1.88
+ $X2=5.245 $Y2=2.495
r124 13 39 318.742 $w=1.8e-07 $l=8.2e-07 $layer=POLY_cond $X=7.18 $Y=2.34
+ $X2=7.18 $Y2=1.52
r125 9 38 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=7.165 $Y=0.645
+ $X2=7.165 $Y2=1.19
r126 2 17 600 $w=1.7e-07 $l=4.37321e-07 $layer=licon1_PDIFF $count=1 $X=5.11
+ $Y=2.12 $X2=5.245 $Y2=2.495
r127 1 21 182 $w=1.7e-07 $l=5.30542e-07 $layer=licon1_NDIFF $count=1 $X=5.2
+ $Y=0.375 $X2=5.49 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_2%VPWR 1 2 3 4 5 6 23 27 31 33 35 39 41 46 54
+ 59 64 70 73 80 87 90 94
r103 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r104 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r105 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r106 83 84 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r107 80 83 8.27395 $w=3.88e-07 $l=2.8e-07 $layer=LI1_cond $X=3.905 $Y=3.05
+ $X2=3.905 $Y2=3.33
r108 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r109 73 76 8.96345 $w=3.58e-07 $l=2.8e-07 $layer=LI1_cond $X=1.755 $Y=3.05
+ $X2=1.755 $Y2=3.33
r110 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r111 68 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r112 68 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r113 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r114 65 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.57 $Y=3.33
+ $X2=7.405 $Y2=3.33
r115 65 67 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.57 $Y=3.33
+ $X2=7.92 $Y2=3.33
r116 64 93 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=8.275 $Y=3.33
+ $X2=8.457 $Y2=3.33
r117 64 67 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.275 $Y=3.33
+ $X2=7.92 $Y2=3.33
r118 63 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r119 63 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r120 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r121 60 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.565 $Y=3.33
+ $X2=6.4 $Y2=3.33
r122 60 62 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.565 $Y=3.33
+ $X2=6.96 $Y2=3.33
r123 59 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.24 $Y=3.33
+ $X2=7.405 $Y2=3.33
r124 59 62 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.24 $Y=3.33
+ $X2=6.96 $Y2=3.33
r125 58 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r126 57 58 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r127 55 83 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.1 $Y=3.33
+ $X2=3.905 $Y2=3.33
r128 55 57 123.957 $w=1.68e-07 $l=1.9e-06 $layer=LI1_cond $X=4.1 $Y=3.33 $X2=6
+ $Y2=3.33
r129 54 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.235 $Y=3.33
+ $X2=6.4 $Y2=3.33
r130 54 57 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.235 $Y=3.33
+ $X2=6 $Y2=3.33
r131 53 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r132 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r133 50 53 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r134 50 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r135 49 52 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r136 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r137 47 76 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.935 $Y=3.33
+ $X2=1.755 $Y2=3.33
r138 47 49 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.935 $Y=3.33
+ $X2=2.16 $Y2=3.33
r139 46 83 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=3.71 $Y=3.33
+ $X2=3.905 $Y2=3.33
r140 46 52 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.71 $Y=3.33
+ $X2=3.6 $Y2=3.33
r141 45 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r142 45 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r143 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r144 42 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.73 $Y2=3.33
r145 42 44 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=1.2 $Y2=3.33
r146 41 76 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.755 $Y2=3.33
r147 41 44 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.2 $Y2=3.33
r148 39 58 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=6 $Y2=3.33
r149 39 84 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r150 35 38 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=8.4 $Y=1.985
+ $X2=8.4 $Y2=2.815
r151 33 93 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.4 $Y=3.245
+ $X2=8.457 $Y2=3.33
r152 33 38 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.4 $Y=3.245 $X2=8.4
+ $Y2=2.815
r153 29 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.405 $Y=3.245
+ $X2=7.405 $Y2=3.33
r154 29 31 36.6686 $w=3.28e-07 $l=1.05e-06 $layer=LI1_cond $X=7.405 $Y=3.245
+ $X2=7.405 $Y2=2.195
r155 25 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.4 $Y=3.245 $X2=6.4
+ $Y2=3.33
r156 25 27 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=6.4 $Y=3.245
+ $X2=6.4 $Y2=2.75
r157 21 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r158 21 23 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.455
r159 6 38 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.225
+ $Y=1.84 $X2=8.36 $Y2=2.815
r160 6 35 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.225
+ $Y=1.84 $X2=8.36 $Y2=1.985
r161 5 31 300 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_PDIFF $count=2 $X=7.27
+ $Y=1.84 $X2=7.405 $Y2=2.195
r162 4 27 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=6.265
+ $Y=2.54 $X2=6.4 $Y2=2.75
r163 3 80 600 $w=1.7e-07 $l=6.42962e-07 $layer=licon1_PDIFF $count=1 $X=3.655
+ $Y=2.52 $X2=3.905 $Y2=3.05
r164 2 73 600 $w=1.7e-07 $l=5.84551e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=2.54 $X2=1.755 $Y2=3.05
r165 1 23 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_2%A_434_508# 1 2 9 15 17 18 21
c44 9 0 6.76432e-20 $X=2.39 $Y=2.29
r45 19 21 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.53 $Y=1.235
+ $X2=2.775 $Y2=1.235
r46 17 18 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.42 $Y=1.65
+ $X2=2.42 $Y2=1.82
r47 13 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=1.15
+ $X2=2.775 $Y2=1.235
r48 13 15 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.775 $Y=1.15
+ $X2=2.775 $Y2=0.815
r49 11 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=1.32
+ $X2=2.53 $Y2=1.235
r50 11 17 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.53 $Y=1.32
+ $X2=2.53 $Y2=1.65
r51 9 18 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=2.39 $Y=2.29 $X2=2.39
+ $Y2=1.82
r52 2 9 600 $w=1.7e-07 $l=3.42783e-07 $layer=licon1_PDIFF $count=1 $X=2.17
+ $Y=2.54 $X2=2.39 $Y2=2.29
r53 1 15 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=2.635
+ $Y=0.595 $X2=2.775 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_2%Q 1 2 9 15 16 17 18 19
c35 17 0 2.55617e-20 $X=7.935 $Y=1.13
r36 18 19 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=7.925 $Y=2.405
+ $X2=7.925 $Y2=2.775
r37 16 17 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=8.02 $Y=2.03 $X2=8.02
+ $Y2=1.13
r38 15 16 6.59029 $w=3.58e-07 $l=1.05e-07 $layer=LI1_cond $X=7.925 $Y=2.135
+ $X2=7.925 $Y2=2.03
r39 13 18 6.2424 $w=3.58e-07 $l=1.95e-07 $layer=LI1_cond $X=7.925 $Y=2.21
+ $X2=7.925 $Y2=2.405
r40 13 15 2.40092 $w=3.58e-07 $l=7.5e-08 $layer=LI1_cond $X=7.925 $Y=2.21
+ $X2=7.925 $Y2=2.135
r41 7 17 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=7.935 $Y=0.96
+ $X2=7.935 $Y2=1.13
r42 7 9 15.0834 $w=3.38e-07 $l=4.45e-07 $layer=LI1_cond $X=7.935 $Y=0.96
+ $X2=7.935 $Y2=0.515
r43 2 19 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.775
+ $Y=1.84 $X2=7.91 $Y2=2.815
r44 2 15 400 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_PDIFF $count=1 $X=7.775
+ $Y=1.84 $X2=7.91 $Y2=2.135
r45 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.79
+ $Y=0.37 $X2=7.93 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFXTP_2%VGND 1 2 3 4 5 6 21 25 29 33 37 39 41 44 45
+ 46 48 53 58 70 74 80 83 86 89 93
r116 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r117 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r118 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r119 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r120 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r121 78 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r122 78 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r123 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r124 75 89 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=7.595 $Y=0
+ $X2=7.447 $Y2=0
r125 75 77 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.595 $Y=0
+ $X2=7.92 $Y2=0
r126 74 92 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=8.275 $Y=0
+ $X2=8.457 $Y2=0
r127 74 77 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.275 $Y=0
+ $X2=7.92 $Y2=0
r128 73 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r129 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r130 70 89 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=7.3 $Y=0 $X2=7.447
+ $Y2=0
r131 70 72 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.3 $Y=0 $X2=6.96
+ $Y2=0
r132 69 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r133 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r134 66 69 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=6
+ $Y2=0
r135 65 68 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6
+ $Y2=0
r136 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r137 63 86 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.235 $Y=0 $X2=4.11
+ $Y2=0
r138 63 65 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.235 $Y=0
+ $X2=4.56 $Y2=0
r139 62 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r140 62 84 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.16
+ $Y2=0
r141 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r142 59 83 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.082
+ $Y2=0
r143 59 61 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=2.18 $Y=0 $X2=3.6
+ $Y2=0
r144 58 86 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.985 $Y=0 $X2=4.11
+ $Y2=0
r145 58 61 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.985 $Y=0 $X2=3.6
+ $Y2=0
r146 57 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r147 57 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r148 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r149 54 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.67
+ $Y2=0
r150 54 56 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=1.68
+ $Y2=0
r151 53 83 5.78184 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=1.985 $Y=0 $X2=2.082
+ $Y2=0
r152 53 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=0
+ $X2=1.68 $Y2=0
r153 51 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r154 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r155 48 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.67
+ $Y2=0
r156 48 50 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r157 46 66 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.56 $Y2=0
r158 46 87 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.08 $Y2=0
r159 44 68 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.225 $Y=0 $X2=6
+ $Y2=0
r160 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.225 $Y=0 $X2=6.39
+ $Y2=0
r161 43 72 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=6.555 $Y=0
+ $X2=6.96 $Y2=0
r162 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.555 $Y=0 $X2=6.39
+ $Y2=0
r163 39 92 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.4 $Y=0.085
+ $X2=8.457 $Y2=0
r164 39 41 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.4 $Y=0.085 $X2=8.4
+ $Y2=0.515
r165 35 89 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=7.447 $Y=0.085
+ $X2=7.447 $Y2=0
r166 35 37 16.7983 $w=2.93e-07 $l=4.3e-07 $layer=LI1_cond $X=7.447 $Y=0.085
+ $X2=7.447 $Y2=0.515
r167 31 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.39 $Y=0.085
+ $X2=6.39 $Y2=0
r168 31 33 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=6.39 $Y=0.085
+ $X2=6.39 $Y2=0.83
r169 27 86 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=0.085
+ $X2=4.11 $Y2=0
r170 27 29 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=4.11 $Y=0.085
+ $X2=4.11 $Y2=0.355
r171 23 83 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.082 $Y=0.085
+ $X2=2.082 $Y2=0
r172 23 25 22.1818 $w=1.93e-07 $l=3.9e-07 $layer=LI1_cond $X=2.082 $Y=0.085
+ $X2=2.082 $Y2=0.475
r173 19 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0
r174 19 21 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0.57
r175 6 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.22
+ $Y=0.37 $X2=8.36 $Y2=0.515
r176 5 37 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=7.24
+ $Y=0.37 $X2=7.405 $Y2=0.515
r177 4 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.25
+ $Y=0.62 $X2=6.39 $Y2=0.83
r178 3 29 182 $w=1.7e-07 $l=2.85307e-07 $layer=licon1_NDIFF $count=1 $X=3.93
+ $Y=0.505 $X2=4.15 $Y2=0.355
r179 2 25 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=1.925
+ $Y=0.33 $X2=2.08 $Y2=0.475
r180 1 21 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.57
.ends


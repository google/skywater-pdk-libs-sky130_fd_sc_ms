* NGSPICE file created from sky130_fd_sc_ms__nand2_4.ext - technology: sky130A

.subckt sky130_fd_sc_ms__nand2_4 A B VGND VNB VPB VPWR Y
M1000 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=1.0472e+12p pd=8.59e+06u as=2.6824e+12p ps=9.27e+06u
M1001 Y B VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=5.365e+11p pd=4.41e+06u as=1.1581e+12p ps=1.053e+07u
M1003 a_27_74# A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND B a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=0p ps=0u
M1005 Y A a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_74# A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND B a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_74# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__mux2_1.pex.spice
* Created: Fri Aug 28 17:39:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__MUX2_1%S 3 7 11 15 18 19 20 21 25
c56 15 0 1.07726e-19 $X=1.055 $Y=0.74
c57 3 0 3.23367e-20 $X=0.505 $Y=2.26
r58 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.67
+ $Y=1.515 $X2=0.67 $Y2=1.515
r59 21 25 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.67 $Y=1.665
+ $X2=0.67 $Y2=1.515
r60 19 24 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=0.95 $Y=1.515
+ $X2=0.67 $Y2=1.515
r61 19 20 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.95 $Y=1.515 $X2=1.04
+ $Y2=1.515
r62 17 24 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.595 $Y=1.515
+ $X2=0.67 $Y2=1.515
r63 17 18 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.595 $Y=1.515
+ $X2=0.505 $Y2=1.515
r64 13 20 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=1.055 $Y=1.35
+ $X2=1.04 $Y2=1.515
r65 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.055 $Y=1.35
+ $X2=1.055 $Y2=0.74
r66 9 20 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.04 $Y=1.68
+ $X2=1.04 $Y2=1.515
r67 9 11 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.04 $Y=1.68 $X2=1.04
+ $Y2=2.34
r68 5 18 34.7346 $w=1.65e-07 $l=1.69926e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.505 $Y2=1.515
r69 5 7 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.835
r70 1 18 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.68
+ $X2=0.505 $Y2=1.515
r71 1 3 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=0.505 $Y=1.68
+ $X2=0.505 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2_1%A1 3 6 9 10 11 14 16 18 19 24 27 31
c65 24 0 1.32486e-19 $X=1.51 $Y=1.22
c66 11 0 1.07726e-19 $X=1.685 $Y=0.895
r67 27 30 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.62 $Y=1.385
+ $X2=2.62 $Y2=1.55
r68 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.62
+ $Y=1.385 $X2=2.62 $Y2=1.385
r69 19 28 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.62 $Y=1.295 $X2=2.62
+ $Y2=1.385
r70 18 31 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=0.895 $X2=2.62
+ $Y2=0.98
r71 18 19 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=2.62 $Y=0.995 $X2=2.62
+ $Y2=1.295
r72 18 31 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.62 $Y=0.995
+ $X2=2.62 $Y2=0.98
r73 14 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.51 $Y=1.385
+ $X2=1.51 $Y2=1.22
r74 13 16 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.51 $Y=1.385 $X2=1.6
+ $Y2=1.385
r75 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.51
+ $Y=1.385 $X2=1.51 $Y2=1.385
r76 10 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.455 $Y=0.895
+ $X2=2.62 $Y2=0.895
r77 10 11 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.455 $Y=0.895
+ $X2=1.685 $Y2=0.895
r78 9 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.6 $Y=1.22 $X2=1.6
+ $Y2=1.385
r79 8 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.6 $Y=0.98
+ $X2=1.685 $Y2=0.895
r80 8 9 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.6 $Y=0.98 $X2=1.6
+ $Y2=1.22
r81 6 30 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=2.545 $Y=2.34
+ $X2=2.545 $Y2=1.55
r82 3 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.445 $Y=0.74
+ $X2=1.445 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2_1%A0 3 7 8 11 13
c32 8 0 1.1756e-19 $X=2.16 $Y=1.295
r33 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.05 $Y=1.385
+ $X2=2.05 $Y2=1.55
r34 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.05 $Y=1.385
+ $X2=2.05 $Y2=1.22
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.05
+ $Y=1.385 $X2=2.05 $Y2=1.385
r36 8 12 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.16 $Y=1.365
+ $X2=2.05 $Y2=1.365
r37 7 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.14 $Y=0.74 $X2=2.14
+ $Y2=1.22
r38 3 14 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=2.005 $Y=2.34
+ $X2=2.005 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2_1%A_27_112# 1 2 9 13 17 20 23 26 27 28 30 31 33
+ 37 38
c94 37 0 1.1743e-19 $X=3.19 $Y=1.485
c95 9 0 8.6251e-20 $X=3.1 $Y=0.74
r96 38 42 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.19 $Y=1.485
+ $X2=3.19 $Y2=1.65
r97 38 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.19 $Y=1.485
+ $X2=3.19 $Y2=1.32
r98 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.19
+ $Y=1.485 $X2=3.19 $Y2=1.485
r99 34 37 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.04 $Y=1.485
+ $X2=3.19 $Y2=1.485
r100 29 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.04 $Y=1.65
+ $X2=3.04 $Y2=1.485
r101 29 30 81.877 $w=1.68e-07 $l=1.255e-06 $layer=LI1_cond $X=3.04 $Y=1.65
+ $X2=3.04 $Y2=2.905
r102 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.955 $Y=2.99
+ $X2=3.04 $Y2=2.905
r103 27 28 106.668 $w=1.68e-07 $l=1.635e-06 $layer=LI1_cond $X=2.955 $Y=2.99
+ $X2=1.32 $Y2=2.99
r104 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.235 $Y=2.905
+ $X2=1.32 $Y2=2.99
r105 25 26 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.235 $Y=2.23
+ $X2=1.235 $Y2=2.905
r106 24 33 2.76166 $w=1.7e-07 $l=1.90526e-07 $layer=LI1_cond $X=0.445 $Y=2.145
+ $X2=0.28 $Y2=2.09
r107 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.15 $Y=2.145
+ $X2=1.235 $Y2=2.23
r108 23 24 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=1.15 $Y=2.145
+ $X2=0.445 $Y2=2.145
r109 20 33 3.70735 $w=2.5e-07 $l=1.75499e-07 $layer=LI1_cond $X=0.2 $Y=1.95
+ $X2=0.28 $Y2=2.09
r110 20 31 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.2 $Y=1.95 $X2=0.2
+ $Y2=1.13
r111 15 31 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=0.965
+ $X2=0.28 $Y2=1.13
r112 15 17 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.28 $Y=0.965
+ $X2=0.28 $Y2=0.835
r113 13 42 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=3.115 $Y=2.34
+ $X2=3.115 $Y2=1.65
r114 9 41 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.1 $Y=0.74 $X2=3.1
+ $Y2=1.32
r115 2 33 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.06
r116 1 17 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.28 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2_1%A_304_74# 1 2 9 13 16 18 19 20 21 22 27 30 31
+ 32 34 37 42 43
c109 43 0 1.16478e-19 $X=3.73 $Y=1.465
c110 16 0 3.23367e-20 $X=1.09 $Y=1.72
c111 9 0 1.1743e-19 $X=3.735 $Y=2.4
r112 43 47 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=1.465
+ $X2=3.73 $Y2=1.63
r113 43 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=1.465
+ $X2=3.73 $Y2=1.3
r114 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.73
+ $Y=1.465 $X2=3.73 $Y2=1.465
r115 39 42 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=3.61 $Y=1.465
+ $X2=3.73 $Y2=1.465
r116 35 37 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.09 $Y=0.935
+ $X2=1.26 $Y2=0.935
r117 34 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.61 $Y=1.3
+ $X2=3.61 $Y2=1.465
r118 33 34 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.61 $Y=1.15
+ $X2=3.61 $Y2=1.3
r119 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.525 $Y=1.065
+ $X2=3.61 $Y2=1.15
r120 31 32 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.525 $Y=1.065
+ $X2=3.125 $Y2=1.065
r121 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.04 $Y=0.98
+ $X2=3.125 $Y2=1.065
r122 29 30 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.04 $Y=0.64
+ $X2=3.04 $Y2=0.98
r123 25 27 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.23 $Y=1.89
+ $X2=2.23 $Y2=1.985
r124 22 24 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=1.345 $Y=0.515
+ $X2=1.79 $Y2=0.515
r125 21 29 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.955 $Y=0.515
+ $X2=3.04 $Y2=0.64
r126 21 24 53.7038 $w=2.48e-07 $l=1.165e-06 $layer=LI1_cond $X=2.955 $Y=0.515
+ $X2=1.79 $Y2=0.515
r127 19 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.065 $Y=1.805
+ $X2=2.23 $Y2=1.89
r128 19 20 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=2.065 $Y=1.805
+ $X2=1.175 $Y2=1.805
r129 18 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.26 $Y=0.85
+ $X2=1.26 $Y2=0.935
r130 17 22 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.26 $Y=0.64
+ $X2=1.345 $Y2=0.515
r131 17 18 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.26 $Y=0.64
+ $X2=1.26 $Y2=0.85
r132 16 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.09 $Y=1.72
+ $X2=1.175 $Y2=1.805
r133 15 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.09 $Y=1.02
+ $X2=1.09 $Y2=0.935
r134 15 16 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.09 $Y=1.02 $X2=1.09
+ $Y2=1.72
r135 13 46 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.815 $Y=0.74
+ $X2=3.815 $Y2=1.3
r136 9 47 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=3.735 $Y=2.4
+ $X2=3.735 $Y2=1.63
r137 2 27 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.095
+ $Y=1.84 $X2=2.23 $Y2=1.985
r138 1 24 182 $w=1.7e-07 $l=3.505e-07 $layer=licon1_NDIFF $count=1 $X=1.52
+ $Y=0.37 $X2=1.79 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2_1%VPWR 1 2 11 15 20 21 22 32 33 36
r43 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r45 30 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r46 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 27 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 26 29 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 26 27 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 24 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r51 24 26 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33 $X2=1.2
+ $Y2=3.33
r52 22 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r53 22 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r54 20 29 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.295 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=3.33
+ $X2=3.46 $Y2=3.33
r56 19 32 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.625 $Y=3.33
+ $X2=4.08 $Y2=3.33
r57 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.625 $Y=3.33
+ $X2=3.46 $Y2=3.33
r58 15 18 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.46 $Y=1.985
+ $X2=3.46 $Y2=2.815
r59 13 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=3.245
+ $X2=3.46 $Y2=3.33
r60 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.46 $Y=3.245
+ $X2=3.46 $Y2=2.815
r61 9 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r62 9 11 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.51
r63 2 18 600 $w=1.7e-07 $l=1.0951e-06 $layer=licon1_PDIFF $count=1 $X=3.205
+ $Y=1.84 $X2=3.46 $Y2=2.815
r64 2 15 300 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=2 $X=3.205
+ $Y=1.84 $X2=3.46 $Y2=1.985
r65 1 11 600 $w=1.7e-07 $l=7.72205e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.815 $Y2=2.51
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2_1%X 1 2 9 13 14 15 16 31 32 35
c26 13 0 2.02729e-19 $X=4.05 $Y=1.13
r27 31 32 8.83531 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=4.015 $Y=1.985
+ $X2=4.015 $Y2=1.82
r28 21 35 0.130959 $w=4.38e-07 $l=5e-09 $layer=LI1_cond $X=4.015 $Y=2.04
+ $X2=4.015 $Y2=2.035
r29 16 28 1.04768 $w=4.38e-07 $l=4e-08 $layer=LI1_cond $X=4.015 $Y=2.775
+ $X2=4.015 $Y2=2.815
r30 15 16 9.691 $w=4.38e-07 $l=3.7e-07 $layer=LI1_cond $X=4.015 $Y=2.405
+ $X2=4.015 $Y2=2.775
r31 14 35 1.04768 $w=4.38e-07 $l=4e-08 $layer=LI1_cond $X=4.015 $Y=1.995
+ $X2=4.015 $Y2=2.035
r32 14 31 0.261919 $w=4.38e-07 $l=1e-08 $layer=LI1_cond $X=4.015 $Y=1.995
+ $X2=4.015 $Y2=1.985
r33 14 15 8.51236 $w=4.38e-07 $l=3.25e-07 $layer=LI1_cond $X=4.015 $Y=2.08
+ $X2=4.015 $Y2=2.405
r34 14 21 1.04768 $w=4.38e-07 $l=4e-08 $layer=LI1_cond $X=4.015 $Y=2.08
+ $X2=4.015 $Y2=2.04
r35 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.15 $Y=1.13 $X2=4.15
+ $Y2=1.82
r36 7 13 9.16175 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.05 $Y=0.945
+ $X2=4.05 $Y2=1.13
r37 7 9 13.3933 $w=3.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.05 $Y=0.945 $X2=4.05
+ $Y2=0.515
r38 2 31 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.825
+ $Y=1.84 $X2=3.96 $Y2=1.985
r39 2 28 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.825
+ $Y=1.84 $X2=3.96 $Y2=2.815
r40 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.89
+ $Y=0.37 $X2=4.03 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__MUX2_1%VGND 1 2 8 11 15 18 21 22 23 25 38 39 42
c51 18 0 1.49261e-20 $X=0.815 $Y=0.515
r52 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r53 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r54 36 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r55 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r56 33 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r57 32 35 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r58 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r59 30 42 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=0.815
+ $Y2=0
r60 30 32 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=1.2
+ $Y2=0
r61 28 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r62 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r63 25 42 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.815
+ $Y2=0
r64 25 27 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.24
+ $Y2=0
r65 23 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r66 23 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r67 21 35 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.295 $Y=0 $X2=3.12
+ $Y2=0
r68 21 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=0 $X2=3.46
+ $Y2=0
r69 20 38 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.625 $Y=0 $X2=4.08
+ $Y2=0
r70 20 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.625 $Y=0 $X2=3.46
+ $Y2=0
r71 18 19 7.29301 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=0.815 $Y=0.515
+ $X2=0.815 $Y2=0.68
r72 13 22 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=0.085
+ $X2=3.46 $Y2=0
r73 13 15 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=3.46 $Y=0.085
+ $X2=3.46 $Y2=0.645
r74 11 19 15.0519 $w=2.08e-07 $l=2.85e-07 $layer=LI1_cond $X=0.73 $Y=0.965
+ $X2=0.73 $Y2=0.68
r75 8 18 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=0.815 $Y=0.49
+ $X2=0.815 $Y2=0.515
r76 7 42 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0
r77 7 8 12.2826 $w=3.78e-07 $l=4.05e-07 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0.49
r78 2 15 182 $w=1.7e-07 $l=3.995e-07 $layer=licon1_NDIFF $count=1 $X=3.175
+ $Y=0.37 $X2=3.46 $Y2=0.645
r79 1 18 182 $w=1.7e-07 $l=2.66552e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.56 $X2=0.815 $Y2=0.515
r80 1 11 182 $w=1.7e-07 $l=4.76235e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.56 $X2=0.725 $Y2=0.965
.ends


* File: sky130_fd_sc_ms__a22oi_4.spice
* Created: Wed Sep  2 11:53:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a22oi_4.pex.spice"
.subckt sky130_fd_sc_ms__a22oi_4  VNB VPB B2 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_B2_M1005_g N_A_48_74#_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1005_d N_B2_M1010_g N_A_48_74#_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1014_d N_B2_M1014_g N_A_48_74#_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1028 N_VGND_M1014_d N_B2_M1028_g N_A_48_74#_M1028_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1001 N_A_48_74#_M1028_s N_B1_M1001_g N_Y_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1002 N_A_48_74#_M1002_d N_B1_M1002_g N_Y_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1024 N_A_48_74#_M1002_d N_B1_M1024_g N_Y_M1024_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1025 N_A_48_74#_M1025_d N_B1_M1025_g N_Y_M1024_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_A_840_74#_M1009_d N_A1_M1009_g N_Y_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1017 N_A_840_74#_M1017_d N_A1_M1017_g N_Y_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1027 N_A_840_74#_M1017_d N_A1_M1027_g N_Y_M1027_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1030 N_A_840_74#_M1030_d N_A1_M1030_g N_Y_M1027_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_A2_M1012_g N_A_840_74#_M1030_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1012_d N_A2_M1013_g N_A_840_74#_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_A2_M1015_g N_A_840_74#_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1029 N_VGND_M1015_d N_A2_M1029_g N_A_840_74#_M1029_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1003_d N_B2_M1003_g N_A_45_368#_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90007.1 A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1003_d N_B2_M1004_g N_A_45_368#_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90006.7 A=0.2016 P=2.6 MULT=1
MM1006 N_Y_M1006_d N_B2_M1006_g N_A_45_368#_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90006.2 A=0.2016 P=2.6 MULT=1
MM1007 N_Y_M1006_d N_B2_M1007_g N_A_45_368#_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90005.8 A=0.2016 P=2.6 MULT=1
MM1008 N_Y_M1008_d N_B1_M1008_g N_A_45_368#_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90005.3 A=0.2016 P=2.6 MULT=1
MM1011 N_Y_M1008_d N_B1_M1011_g N_A_45_368#_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.4
+ SB=90004.9 A=0.2016 P=2.6 MULT=1
MM1016 N_Y_M1016_d N_B1_M1016_g N_A_45_368#_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.9
+ SB=90004.4 A=0.2016 P=2.6 MULT=1
MM1019 N_Y_M1016_d N_B1_M1019_g N_A_45_368#_M1019_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.3
+ SB=90004 A=0.2016 P=2.6 MULT=1
MM1018 N_A_45_368#_M1019_s N_A1_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.8
+ SB=90003.5 A=0.2016 P=2.6 MULT=1
MM1020 N_A_45_368#_M1020_d N_A1_M1020_g N_VPWR_M1018_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.2
+ SB=90003.1 A=0.2016 P=2.6 MULT=1
MM1022 N_A_45_368#_M1020_d N_A1_M1022_g N_VPWR_M1022_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.28 PD=1.39 PS=1.62 NRD=0 NRS=19.3454 M=1 R=6.22222 SA=90004.7
+ SB=90002.6 A=0.2016 P=2.6 MULT=1
MM1031 N_A_45_368#_M1031_d N_A1_M1031_g N_VPWR_M1022_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.28 PD=1.39 PS=1.62 NRD=0 NRS=19.3454 M=1 R=6.22222 SA=90005.3
+ SB=90002 A=0.2016 P=2.6 MULT=1
MM1000 N_A_45_368#_M1031_d N_A2_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90005.8
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1021 N_A_45_368#_M1021_d N_A2_M1021_g N_VPWR_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90006.2
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1023 N_A_45_368#_M1021_d N_A2_M1023_g N_VPWR_M1023_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90006.7
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1026 N_A_45_368#_M1026_d N_A2_M1026_g N_VPWR_M1023_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2912 AS=0.1512 PD=2.76 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90007.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX32_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_ms__a22oi_4.pxi.spice"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 a_280_107# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=6.5505e+11p pd=6.27e+06u as=4.033e+11p ps=4.05e+06u
M1001 a_280_107# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=5.83425e+11p ps=4.82e+06u
M1002 VGND A2 a_280_107# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y B1 a_131_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.1872e+12p ps=1.108e+07u
M1004 a_131_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A2 a_131_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.72e+11p pd=5.68e+06u as=0p ps=0u
M1006 Y A1 a_280_107# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_131_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_131_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_131_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

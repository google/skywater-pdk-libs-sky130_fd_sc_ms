* File: sky130_fd_sc_ms__decap_4.pex.spice
* Created: Fri Aug 28 17:20:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DECAP_4%VGND 1 9 12 14 17 19 21 23 27 37
r25 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r26 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r27 31 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r28 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r29 28 33 6.71932 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=0.74 $Y=0 $X2=0.37
+ $Y2=0
r30 28 30 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=0.74 $Y=0 $X2=1.2
+ $Y2=0
r31 27 36 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.685
+ $Y2=0
r32 27 30 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.2
+ $Y2=0
r33 23 31 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r34 23 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.24
+ $Y2=0
r35 19 36 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=1.615 $Y=0.085
+ $X2=1.685 $Y2=0
r36 19 21 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=1.615 $Y=0.085
+ $X2=1.615 $Y2=0.64
r37 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.575
+ $Y=1.42 $X2=0.575 $Y2=1.42
r38 14 16 16.3674 $w=5.68e-07 $l=7.8e-07 $layer=LI1_cond $X=0.455 $Y=0.64
+ $X2=0.455 $Y2=1.42
r39 12 33 3.08726 $w=5.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.455 $Y=0.085
+ $X2=0.37 $Y2=0
r40 12 14 11.646 $w=5.68e-07 $l=5.55e-07 $layer=LI1_cond $X=0.455 $Y=0.085
+ $X2=0.455 $Y2=0.64
r41 10 17 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=0.575 $Y=1.83
+ $X2=0.575 $Y2=1.42
r42 9 10 57.2398 $w=1e-06 $l=6.3e-07 $layer=POLY_cond $X=0.91 $Y=2.46 $X2=0.91
+ $Y2=1.83
r43 1 21 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=1.475
+ $Y=0.425 $X2=1.615 $Y2=0.64
r44 1 14 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=1.475
+ $Y=0.425 $X2=0.335 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_MS__DECAP_4%VPWR 1 8 10 13 15 19 21 23 24 30 39
r26 39 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r27 38 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r28 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r29 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 30 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.2 $Y2=3.33
r31 30 36 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.24 $Y2=3.33
r32 27 29 14.8985 $w=5.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.43 $Y=2.105
+ $X2=1.43 $Y2=2.815
r33 23 27 14.4788 $w=5.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.43 $Y=1.415
+ $X2=1.43 $Y2=2.105
r34 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.31
+ $Y=1.415 $X2=1.31 $Y2=1.415
r35 21 38 3.19482 $w=5.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=1.43 $Y=3.245
+ $X2=1.532 $Y2=3.33
r36 21 29 9.02305 $w=5.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.43 $Y=3.245
+ $X2=1.43 $Y2=2.815
r37 20 35 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r38 19 38 6.61175 $w=1.7e-07 $l=3.87e-07 $layer=LI1_cond $X=1.145 $Y=3.33
+ $X2=1.532 $Y2=3.33
r39 19 20 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.145 $Y=3.33
+ $X2=0.425 $Y2=3.33
r40 15 18 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.26 $Y=2.105
+ $X2=0.26 $Y2=2.815
r41 13 35 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r42 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.815
r43 11 24 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=1.31 $Y=1.045
+ $X2=1.31 $Y2=1.415
r44 10 11 23.8477 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=1.31 $Y=0.64
+ $X2=1.31 $Y2=1.045
r45 8 10 21.2651 $w=8.1e-07 $l=3.35e-07 $layer=POLY_cond $X=0.975 $Y=0.64
+ $X2=1.31 $Y2=0.64
r46 1 29 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.96 $X2=1.55 $Y2=2.815
r47 1 27 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.96 $X2=1.55 $Y2=2.105
r48 1 18 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.96 $X2=0.26 $Y2=2.815
r49 1 15 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.96 $X2=0.26 $Y2=2.105
.ends


* File: sky130_fd_sc_ms__o21ai_1.pxi.spice
* Created: Fri Aug 28 17:54:29 2020
* 
x_PM_SKY130_FD_SC_MS__O21AI_1%A1 N_A1_c_39_n N_A1_M1005_g N_A1_M1001_g A1
+ N_A1_c_41_n N_A1_c_42_n PM_SKY130_FD_SC_MS__O21AI_1%A1
x_PM_SKY130_FD_SC_MS__O21AI_1%A2 N_A2_M1004_g N_A2_M1000_g A2 N_A2_c_70_n
+ N_A2_c_71_n PM_SKY130_FD_SC_MS__O21AI_1%A2
x_PM_SKY130_FD_SC_MS__O21AI_1%B1 N_B1_M1002_g N_B1_M1003_g B1 B1 N_B1_c_106_n
+ PM_SKY130_FD_SC_MS__O21AI_1%B1
x_PM_SKY130_FD_SC_MS__O21AI_1%VPWR N_VPWR_M1001_s N_VPWR_M1002_d N_VPWR_c_133_n
+ N_VPWR_c_134_n N_VPWR_c_135_n N_VPWR_c_136_n N_VPWR_c_137_n VPWR
+ N_VPWR_c_138_n N_VPWR_c_132_n PM_SKY130_FD_SC_MS__O21AI_1%VPWR
x_PM_SKY130_FD_SC_MS__O21AI_1%Y N_Y_M1003_d N_Y_M1004_d N_Y_c_159_n N_Y_c_160_n
+ N_Y_c_161_n Y Y N_Y_c_163_n N_Y_c_162_n PM_SKY130_FD_SC_MS__O21AI_1%Y
x_PM_SKY130_FD_SC_MS__O21AI_1%A_27_74# N_A_27_74#_M1005_s N_A_27_74#_M1000_d
+ N_A_27_74#_c_199_n N_A_27_74#_c_203_n N_A_27_74#_c_200_n N_A_27_74#_c_201_n
+ PM_SKY130_FD_SC_MS__O21AI_1%A_27_74#
x_PM_SKY130_FD_SC_MS__O21AI_1%VGND N_VGND_M1005_d VGND N_VGND_c_230_n
+ N_VGND_c_231_n N_VGND_c_232_n N_VGND_c_233_n PM_SKY130_FD_SC_MS__O21AI_1%VGND
cc_1 VNB N_A1_c_39_n 0.0240813f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_2 VNB N_A1_M1001_g 0.00857766f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=2.4
cc_3 VNB N_A1_c_41_n 0.0206951f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.385
cc_4 VNB N_A1_c_42_n 0.063848f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.385
cc_5 VNB N_A2_M1000_g 0.0268063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A2_c_70_n 0.00245973f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.385
cc_7 VNB N_A2_c_71_n 0.0322632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B1_M1003_g 0.0329453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB B1 0.01855f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.385
cc_10 VNB N_B1_c_106_n 0.0277039f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.385
cc_11 VNB N_VPWR_c_132_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_Y_c_159_n 0.0231532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_Y_c_160_n 7.88229e-19 $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.385
cc_14 VNB N_Y_c_161_n 0.0281704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_Y_c_162_n 0.00413149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_74#_c_199_n 0.0149177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_c_200_n 0.0139746f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.385
cc_18 VNB N_A_27_74#_c_201_n 0.00256335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_230_n 0.031602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_231_n 0.159013f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.385
cc_21 VNB N_VGND_c_232_n 0.0182531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_233_n 0.023075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VPB N_A1_M1001_g 0.0272611f $X=-0.19 $Y=1.66 $X2=0.735 $Y2=2.4
cc_24 VPB N_A2_M1004_g 0.0232039f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_25 VPB N_A2_c_70_n 0.00203745f $X=-0.19 $Y=1.66 $X2=0.735 $Y2=1.385
cc_26 VPB N_A2_c_71_n 0.008255f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_27 VPB N_B1_M1002_g 0.0276983f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_28 VPB B1 0.0175258f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.385
cc_29 VPB N_B1_c_106_n 0.00579202f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.385
cc_30 VPB N_VPWR_c_133_n 0.0151484f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_134_n 0.0147081f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_135_n 0.0484671f $X=-0.19 $Y=1.66 $X2=0.735 $Y2=1.385
cc_33 VPB N_VPWR_c_136_n 0.011849f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.365
cc_34 VPB N_VPWR_c_137_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_138_n 0.0352341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_132_n 0.0712219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_Y_c_163_n 0.0048658f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.365
cc_38 VPB N_Y_c_162_n 0.0012908f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 N_A1_M1001_g N_A2_M1004_g 0.0468731f $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_40 N_A1_c_42_n N_A2_M1000_g 0.00239f $X=0.735 $Y=1.385 $X2=0 $Y2=0
cc_41 N_A1_c_42_n N_A2_c_70_n 4.75213e-19 $X=0.735 $Y=1.385 $X2=0 $Y2=0
cc_42 N_A1_c_42_n N_A2_c_71_n 0.0468731f $X=0.735 $Y=1.385 $X2=0 $Y2=0
cc_43 N_A1_M1001_g N_VPWR_c_133_n 0.00935256f $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_44 N_A1_c_41_n N_VPWR_c_133_n 0.0149317f $X=0.39 $Y=1.385 $X2=0 $Y2=0
cc_45 N_A1_c_42_n N_VPWR_c_133_n 0.00593824f $X=0.735 $Y=1.385 $X2=0 $Y2=0
cc_46 N_A1_M1001_g N_VPWR_c_138_n 0.00441589f $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_47 N_A1_M1001_g N_VPWR_c_132_n 0.00730489f $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_48 N_A1_c_39_n N_Y_c_160_n 0.00710272f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_49 N_A1_M1001_g N_Y_c_163_n 0.0285831f $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_50 N_A1_c_39_n N_Y_c_162_n 7.57456e-19 $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_51 N_A1_M1001_g N_Y_c_162_n 0.0164193f $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_52 N_A1_c_41_n N_Y_c_162_n 0.0270948f $X=0.39 $Y=1.385 $X2=0 $Y2=0
cc_53 N_A1_c_42_n N_Y_c_162_n 0.0114711f $X=0.735 $Y=1.385 $X2=0 $Y2=0
cc_54 N_A1_c_39_n N_A_27_74#_c_199_n 4.59808e-19 $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_55 N_A1_c_39_n N_A_27_74#_c_203_n 0.0116592f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_56 N_A1_c_41_n N_A_27_74#_c_203_n 0.00452942f $X=0.39 $Y=1.385 $X2=0 $Y2=0
cc_57 N_A1_c_42_n N_A_27_74#_c_203_n 0.00456427f $X=0.735 $Y=1.385 $X2=0 $Y2=0
cc_58 N_A1_c_39_n N_A_27_74#_c_200_n 0.00905744f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_59 N_A1_c_41_n N_A_27_74#_c_200_n 0.0250699f $X=0.39 $Y=1.385 $X2=0 $Y2=0
cc_60 N_A1_c_42_n N_A_27_74#_c_200_n 0.0012195f $X=0.735 $Y=1.385 $X2=0 $Y2=0
cc_61 N_A1_c_39_n N_VGND_c_231_n 0.00429381f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_62 N_A1_c_39_n N_VGND_c_232_n 0.00329909f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_63 N_A1_c_39_n N_VGND_c_233_n 0.00816535f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_64 N_A2_M1004_g N_B1_M1002_g 0.018983f $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_65 N_A2_c_70_n N_B1_M1002_g 2.7523e-19 $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_66 N_A2_M1000_g N_B1_M1003_g 0.0331423f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_67 N_A2_M1004_g B1 3.15296e-19 $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_68 N_A2_c_70_n B1 0.036629f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_69 N_A2_c_71_n B1 0.00262232f $X=1.405 $Y=1.515 $X2=0 $Y2=0
cc_70 N_A2_c_70_n N_B1_c_106_n 2.75737e-19 $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_71 N_A2_c_71_n N_B1_c_106_n 0.0174845f $X=1.405 $Y=1.515 $X2=0 $Y2=0
cc_72 N_A2_M1004_g N_VPWR_c_135_n 8.05794e-19 $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_73 N_A2_M1004_g N_VPWR_c_138_n 0.00349816f $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_74 N_A2_M1004_g N_VPWR_c_132_n 0.00430952f $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_75 N_A2_M1000_g N_Y_c_159_n 0.0147665f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_76 N_A2_c_70_n N_Y_c_159_n 0.0250422f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_77 N_A2_c_71_n N_Y_c_159_n 0.00184421f $X=1.405 $Y=1.515 $X2=0 $Y2=0
cc_78 N_A2_M1004_g N_Y_c_163_n 0.0324826f $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_79 N_A2_c_70_n N_Y_c_163_n 0.0252628f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_80 N_A2_c_71_n N_Y_c_163_n 0.00450805f $X=1.405 $Y=1.515 $X2=0 $Y2=0
cc_81 N_A2_M1000_g N_Y_c_162_n 0.00317248f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_82 N_A2_c_70_n N_Y_c_162_n 0.0322798f $X=1.23 $Y=1.515 $X2=0 $Y2=0
cc_83 N_A2_c_71_n N_Y_c_162_n 0.00589856f $X=1.405 $Y=1.515 $X2=0 $Y2=0
cc_84 N_A2_M1000_g N_A_27_74#_c_203_n 0.01182f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_85 N_A2_M1000_g N_A_27_74#_c_201_n 5.92733e-19 $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_86 N_A2_M1000_g N_VGND_c_230_n 0.00329926f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_87 N_A2_M1000_g N_VGND_c_231_n 0.00425862f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_88 N_A2_M1000_g N_VGND_c_233_n 0.00816535f $X=1.405 $Y=0.74 $X2=0 $Y2=0
cc_89 N_B1_M1002_g N_VPWR_c_135_n 0.0216844f $X=1.81 $Y=2.4 $X2=0 $Y2=0
cc_90 B1 N_VPWR_c_135_n 0.0262242f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_91 N_B1_c_106_n N_VPWR_c_135_n 7.8095e-19 $X=1.885 $Y=1.515 $X2=0 $Y2=0
cc_92 N_B1_M1002_g N_VPWR_c_138_n 0.00460063f $X=1.81 $Y=2.4 $X2=0 $Y2=0
cc_93 N_B1_M1002_g N_VPWR_c_132_n 0.00910297f $X=1.81 $Y=2.4 $X2=0 $Y2=0
cc_94 N_B1_M1003_g N_Y_c_159_n 0.0158149f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_95 B1 N_Y_c_159_n 0.0584272f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_96 N_B1_c_106_n N_Y_c_159_n 0.00427424f $X=1.885 $Y=1.515 $X2=0 $Y2=0
cc_97 N_B1_M1003_g N_Y_c_161_n 0.0128452f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_98 N_B1_M1002_g N_Y_c_163_n 0.011193f $X=1.81 $Y=2.4 $X2=0 $Y2=0
cc_99 N_B1_M1003_g N_A_27_74#_c_203_n 0.00214696f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_100 N_B1_M1003_g N_A_27_74#_c_201_n 0.00475124f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_101 N_B1_M1003_g N_VGND_c_230_n 0.00434272f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_102 N_B1_M1003_g N_VGND_c_231_n 0.00825242f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_103 N_VPWR_c_135_n N_Y_c_163_n 0.0516097f $X=2.035 $Y=2.115 $X2=0 $Y2=0
cc_104 N_VPWR_c_138_n N_Y_c_163_n 0.0356472f $X=1.87 $Y=3.33 $X2=0 $Y2=0
cc_105 N_VPWR_c_132_n N_Y_c_163_n 0.0288601f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_106 N_VPWR_c_133_n N_Y_c_162_n 0.0922408f $X=0.47 $Y=1.985 $X2=0 $Y2=0
cc_107 A_165_368# N_Y_c_163_n 0.00509749f $X=0.825 $Y=1.84 $X2=1.38 $Y2=2.115
cc_108 A_165_368# N_Y_c_162_n 0.00126422f $X=0.825 $Y=1.84 $X2=1.135 $Y2=1.95
cc_109 N_Y_c_159_n N_A_27_74#_M1000_d 0.00176461f $X=1.955 $Y=1.095 $X2=0 $Y2=0
cc_110 N_Y_c_159_n N_A_27_74#_c_203_n 0.0525194f $X=1.955 $Y=1.095 $X2=0 $Y2=0
cc_111 N_Y_c_160_n N_A_27_74#_c_203_n 0.0138309f $X=0.895 $Y=1.095 $X2=0 $Y2=0
cc_112 N_Y_c_161_n N_A_27_74#_c_201_n 0.0126166f $X=2.12 $Y=0.515 $X2=0 $Y2=0
cc_113 N_Y_c_159_n N_VGND_M1005_d 0.00498687f $X=1.955 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_114 N_Y_c_160_n N_VGND_M1005_d 0.00350137f $X=0.895 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_115 N_Y_c_161_n N_VGND_c_230_n 0.0146357f $X=2.12 $Y=0.515 $X2=0 $Y2=0
cc_116 N_Y_c_161_n N_VGND_c_231_n 0.0121141f $X=2.12 $Y=0.515 $X2=0 $Y2=0
cc_117 N_A_27_74#_c_203_n N_VGND_M1005_d 0.0171612f $X=1.48 $Y=0.755 $X2=-0.19
+ $Y2=-0.245
cc_118 N_A_27_74#_c_203_n N_VGND_c_230_n 0.00255882f $X=1.48 $Y=0.755 $X2=0
+ $Y2=0
cc_119 N_A_27_74#_c_201_n N_VGND_c_230_n 0.0131355f $X=1.632 $Y=0.67 $X2=0 $Y2=0
cc_120 N_A_27_74#_c_199_n N_VGND_c_231_n 0.0111794f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_121 N_A_27_74#_c_203_n N_VGND_c_231_n 0.0111174f $X=1.48 $Y=0.755 $X2=0 $Y2=0
cc_122 N_A_27_74#_c_200_n N_VGND_c_231_n 5.83956e-19 $X=0.445 $Y=0.755 $X2=0
+ $Y2=0
cc_123 N_A_27_74#_c_201_n N_VGND_c_231_n 0.0109537f $X=1.632 $Y=0.67 $X2=0 $Y2=0
cc_124 N_A_27_74#_c_199_n N_VGND_c_232_n 0.0134907f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_125 N_A_27_74#_c_203_n N_VGND_c_232_n 0.00218193f $X=1.48 $Y=0.755 $X2=0
+ $Y2=0
cc_126 N_A_27_74#_c_200_n N_VGND_c_232_n 3.88305e-19 $X=0.445 $Y=0.755 $X2=0
+ $Y2=0
cc_127 N_A_27_74#_c_199_n N_VGND_c_233_n 0.00658978f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_128 N_A_27_74#_c_203_n N_VGND_c_233_n 0.0495128f $X=1.48 $Y=0.755 $X2=0 $Y2=0
cc_129 N_A_27_74#_c_201_n N_VGND_c_233_n 0.00309085f $X=1.632 $Y=0.67 $X2=0
+ $Y2=0

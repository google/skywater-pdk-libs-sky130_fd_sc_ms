* File: sky130_fd_sc_ms__o41a_1.pxi.spice
* Created: Fri Aug 28 18:04:34 2020
* 
x_PM_SKY130_FD_SC_MS__O41A_1%A_83_270# N_A_83_270#_M1004_s N_A_83_270#_M1002_d
+ N_A_83_270#_M1000_g N_A_83_270#_M1010_g N_A_83_270#_c_78_n N_A_83_270#_c_73_n
+ N_A_83_270#_c_74_n N_A_83_270#_c_75_n N_A_83_270#_c_80_n N_A_83_270#_c_118_p
+ N_A_83_270#_c_76_n N_A_83_270#_c_81_n PM_SKY130_FD_SC_MS__O41A_1%A_83_270#
x_PM_SKY130_FD_SC_MS__O41A_1%B1 N_B1_M1004_g N_B1_c_144_n N_B1_M1002_g B1
+ N_B1_c_145_n PM_SKY130_FD_SC_MS__O41A_1%B1
x_PM_SKY130_FD_SC_MS__O41A_1%A4 N_A4_M1001_g N_A4_c_181_n N_A4_M1003_g A4
+ N_A4_c_183_n PM_SKY130_FD_SC_MS__O41A_1%A4
x_PM_SKY130_FD_SC_MS__O41A_1%A3 N_A3_M1007_g N_A3_M1011_g A3 A3 A3 A3
+ N_A3_c_227_n N_A3_c_228_n PM_SKY130_FD_SC_MS__O41A_1%A3
x_PM_SKY130_FD_SC_MS__O41A_1%A2 N_A2_M1006_g N_A2_M1005_g A2 A2 A2 A2
+ N_A2_c_271_n N_A2_c_272_n PM_SKY130_FD_SC_MS__O41A_1%A2
x_PM_SKY130_FD_SC_MS__O41A_1%A1 N_A1_M1009_g N_A1_M1008_g A1 A1 N_A1_c_308_n
+ N_A1_c_309_n PM_SKY130_FD_SC_MS__O41A_1%A1
x_PM_SKY130_FD_SC_MS__O41A_1%X N_X_M1010_s N_X_M1000_s N_X_c_335_n N_X_c_336_n X
+ X N_X_c_337_n X PM_SKY130_FD_SC_MS__O41A_1%X
x_PM_SKY130_FD_SC_MS__O41A_1%VPWR N_VPWR_M1000_d N_VPWR_M1009_d N_VPWR_c_357_n
+ N_VPWR_c_358_n N_VPWR_c_359_n VPWR N_VPWR_c_360_n N_VPWR_c_361_n
+ N_VPWR_c_362_n N_VPWR_c_356_n PM_SKY130_FD_SC_MS__O41A_1%VPWR
x_PM_SKY130_FD_SC_MS__O41A_1%VGND N_VGND_M1010_d N_VGND_M1001_d N_VGND_M1006_d
+ N_VGND_c_403_n N_VGND_c_404_n N_VGND_c_405_n N_VGND_c_406_n N_VGND_c_407_n
+ VGND N_VGND_c_408_n N_VGND_c_409_n N_VGND_c_410_n N_VGND_c_411_n
+ N_VGND_c_412_n N_VGND_c_413_n PM_SKY130_FD_SC_MS__O41A_1%VGND
x_PM_SKY130_FD_SC_MS__O41A_1%A_326_74# N_A_326_74#_M1004_d N_A_326_74#_M1011_d
+ N_A_326_74#_M1008_d N_A_326_74#_c_459_n N_A_326_74#_c_460_n
+ N_A_326_74#_c_461_n N_A_326_74#_c_462_n N_A_326_74#_c_463_n
+ N_A_326_74#_c_464_n N_A_326_74#_c_465_n PM_SKY130_FD_SC_MS__O41A_1%A_326_74#
cc_1 VNB N_A_83_270#_M1010_g 0.0303327f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_83_270#_c_73_n 0.00593596f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.515
cc_3 VNB N_A_83_270#_c_74_n 0.033347f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.515
cc_4 VNB N_A_83_270#_c_75_n 0.0192328f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=1.195
cc_5 VNB N_A_83_270#_c_76_n 0.0111398f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=0.515
cc_6 VNB N_B1_M1004_g 0.042114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_B1_c_144_n 0.0229061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B1_c_145_n 0.00319006f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_9 VNB N_A4_M1001_g 0.0237112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A4_c_181_n 0.033205f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A4_M1003_g 0.0067955f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.68
cc_12 VNB N_A4_c_183_n 0.00660497f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_13 VNB N_A3_M1007_g 0.00587431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A3_M1011_g 0.0253751f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.68
cc_15 VNB N_A3_c_227_n 0.0328488f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.515
cc_16 VNB N_A3_c_228_n 0.00250171f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.515
cc_17 VNB N_A2_M1006_g 0.0309777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A2_M1005_g 0.00155616f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.68
cc_19 VNB N_A2_c_271_n 0.0313748f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.515
cc_20 VNB N_A2_c_272_n 0.00505659f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.515
cc_21 VNB N_A1_M1008_g 0.0464113f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.68
cc_22 VNB N_A1_c_308_n 0.0305237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A1_c_309_n 0.0184746f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.515
cc_24 VNB N_X_c_335_n 0.0264414f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_25 VNB N_X_c_336_n 0.00871852f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_26 VNB N_X_c_337_n 0.0247491f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=0.515
cc_27 VNB N_VPWR_c_356_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_403_n 0.0130175f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_29 VNB N_VGND_c_404_n 0.00900728f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.95
cc_30 VNB N_VGND_c_405_n 0.00814066f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=1.195
cc_31 VNB N_VGND_c_406_n 0.0339528f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=2.035
cc_32 VNB N_VGND_c_407_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.11
cc_33 VNB N_VGND_c_408_n 0.0173128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_409_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_410_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_411_n 0.255913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_412_n 0.00750435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_413_n 0.0100141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_326_74#_c_459_n 0.00280384f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_40 VNB N_A_326_74#_c_460_n 0.00829425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_326_74#_c_461_n 0.00864861f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.515
cc_42 VNB N_A_326_74#_c_462_n 0.00280333f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.515
cc_43 VNB N_A_326_74#_c_463_n 0.0225415f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=1.195
cc_44 VNB N_A_326_74#_c_464_n 0.0216332f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.11
cc_45 VNB N_A_326_74#_c_465_n 0.00898142f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=0.515
cc_46 VPB N_A_83_270#_M1000_g 0.0274339f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_47 VPB N_A_83_270#_c_78_n 0.0016796f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.95
cc_48 VPB N_A_83_270#_c_74_n 0.00718091f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.515
cc_49 VPB N_A_83_270#_c_80_n 0.0111243f $X=-0.19 $Y=1.66 $X2=1.75 $Y2=2.035
cc_50 VPB N_A_83_270#_c_81_n 3.36213e-19 $X=-0.19 $Y=1.66 $X2=1.915 $Y2=2.13
cc_51 VPB N_B1_c_144_n 0.0533774f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_B1_c_145_n 0.00256692f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_53 VPB N_A4_M1003_g 0.0239989f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.68
cc_54 VPB N_A4_c_183_n 0.00510077f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_55 VPB N_A3_M1007_g 0.0235268f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A3_c_228_n 0.00120077f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.515
cc_57 VPB N_A2_M1005_g 0.0241831f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.68
cc_58 VPB N_A2_c_272_n 0.00254494f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.515
cc_59 VPB N_A1_M1009_g 0.0262382f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A1_c_308_n 0.00601933f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A1_c_309_n 0.0202663f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.515
cc_62 VPB X 0.00626527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB X 0.0225276f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.515
cc_64 VPB N_X_c_337_n 0.024049f $X=-0.19 $Y=1.66 $X2=1.34 $Y2=0.515
cc_65 VPB N_VPWR_c_357_n 0.0156627f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_66 VPB N_VPWR_c_358_n 0.0142087f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_67 VPB N_VPWR_c_359_n 0.0370109f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_360_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.515
cc_69 VPB N_VPWR_c_361_n 0.0639218f $X=-0.19 $Y=1.66 $X2=0.785 $Y2=2.035
cc_70 VPB N_VPWR_c_362_n 0.0177663f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.195
cc_71 VPB N_VPWR_c_356_n 0.0864649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 N_A_83_270#_c_73_n N_B1_M1004_g 0.00186326f $X=0.62 $Y=1.515 $X2=0 $Y2=0
cc_73 N_A_83_270#_c_74_n N_B1_M1004_g 0.00112947f $X=0.62 $Y=1.515 $X2=0 $Y2=0
cc_74 N_A_83_270#_c_75_n N_B1_M1004_g 0.00743377f $X=1.175 $Y=1.195 $X2=0 $Y2=0
cc_75 N_A_83_270#_c_76_n N_B1_M1004_g 0.0111697f $X=1.34 $Y=0.515 $X2=0 $Y2=0
cc_76 N_A_83_270#_M1000_g N_B1_c_144_n 0.00277372f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_77 N_A_83_270#_c_78_n N_B1_c_144_n 0.00311571f $X=0.62 $Y=1.95 $X2=0 $Y2=0
cc_78 N_A_83_270#_c_74_n N_B1_c_144_n 0.00498282f $X=0.62 $Y=1.515 $X2=0 $Y2=0
cc_79 N_A_83_270#_c_75_n N_B1_c_144_n 0.00572457f $X=1.175 $Y=1.195 $X2=0 $Y2=0
cc_80 N_A_83_270#_c_80_n N_B1_c_144_n 0.0296595f $X=1.75 $Y=2.035 $X2=0 $Y2=0
cc_81 N_A_83_270#_c_81_n N_B1_c_144_n 0.00398164f $X=1.915 $Y=2.13 $X2=0 $Y2=0
cc_82 N_A_83_270#_M1000_g N_B1_c_145_n 3.34568e-19 $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_83 N_A_83_270#_c_78_n N_B1_c_145_n 0.0146046f $X=0.62 $Y=1.95 $X2=0 $Y2=0
cc_84 N_A_83_270#_c_73_n N_B1_c_145_n 0.00345372f $X=0.62 $Y=1.515 $X2=0 $Y2=0
cc_85 N_A_83_270#_c_74_n N_B1_c_145_n 0.0017264f $X=0.62 $Y=1.515 $X2=0 $Y2=0
cc_86 N_A_83_270#_c_75_n N_B1_c_145_n 0.0351249f $X=1.175 $Y=1.195 $X2=0 $Y2=0
cc_87 N_A_83_270#_c_80_n N_B1_c_145_n 0.0376375f $X=1.75 $Y=2.035 $X2=0 $Y2=0
cc_88 N_A_83_270#_c_75_n N_A4_M1001_g 3.72646e-19 $X=1.175 $Y=1.195 $X2=0 $Y2=0
cc_89 N_A_83_270#_c_76_n N_A4_M1001_g 5.94612e-19 $X=1.34 $Y=0.515 $X2=0 $Y2=0
cc_90 N_A_83_270#_c_75_n N_A4_c_181_n 2.73291e-19 $X=1.175 $Y=1.195 $X2=0 $Y2=0
cc_91 N_A_83_270#_c_80_n N_A4_c_181_n 6.87595e-19 $X=1.75 $Y=2.035 $X2=0 $Y2=0
cc_92 N_A_83_270#_c_80_n N_A4_M1003_g 0.00312576f $X=1.75 $Y=2.035 $X2=0 $Y2=0
cc_93 N_A_83_270#_c_81_n N_A4_M1003_g 0.013876f $X=1.915 $Y=2.13 $X2=0 $Y2=0
cc_94 N_A_83_270#_c_75_n N_A4_c_183_n 0.00393762f $X=1.175 $Y=1.195 $X2=0 $Y2=0
cc_95 N_A_83_270#_c_80_n N_A4_c_183_n 0.0161787f $X=1.75 $Y=2.035 $X2=0 $Y2=0
cc_96 N_A_83_270#_c_80_n N_A3_M1007_g 4.46427e-19 $X=1.75 $Y=2.035 $X2=0 $Y2=0
cc_97 N_A_83_270#_c_81_n N_A3_M1007_g 0.00190931f $X=1.915 $Y=2.13 $X2=0 $Y2=0
cc_98 N_A_83_270#_c_80_n N_A3_c_228_n 0.00693615f $X=1.75 $Y=2.035 $X2=0 $Y2=0
cc_99 N_A_83_270#_c_81_n N_A3_c_228_n 0.0278624f $X=1.915 $Y=2.13 $X2=0 $Y2=0
cc_100 N_A_83_270#_M1010_g N_X_c_335_n 0.00207706f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_101 N_A_83_270#_c_73_n N_X_c_336_n 0.00133215f $X=0.62 $Y=1.515 $X2=0 $Y2=0
cc_102 N_A_83_270#_M1000_g X 0.00339366f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_103 N_A_83_270#_M1000_g X 0.0068231f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_104 N_A_83_270#_M1010_g N_X_c_337_n 0.0047754f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A_83_270#_c_78_n N_X_c_337_n 0.0324341f $X=0.62 $Y=1.95 $X2=0 $Y2=0
cc_106 N_A_83_270#_c_73_n N_X_c_337_n 0.0237307f $X=0.62 $Y=1.515 $X2=0 $Y2=0
cc_107 N_A_83_270#_c_74_n N_X_c_337_n 0.0226927f $X=0.62 $Y=1.515 $X2=0 $Y2=0
cc_108 N_A_83_270#_c_118_p N_X_c_337_n 0.0133618f $X=0.785 $Y=2.035 $X2=0 $Y2=0
cc_109 N_A_83_270#_c_78_n N_VPWR_M1000_d 0.00278911f $X=0.62 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_110 N_A_83_270#_c_80_n N_VPWR_M1000_d 0.0125087f $X=1.75 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_111 N_A_83_270#_c_118_p N_VPWR_M1000_d 0.00155484f $X=0.785 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_112 N_A_83_270#_M1000_g N_VPWR_c_357_n 0.00689713f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_113 N_A_83_270#_c_74_n N_VPWR_c_357_n 4.9998e-19 $X=0.62 $Y=1.515 $X2=0 $Y2=0
cc_114 N_A_83_270#_c_80_n N_VPWR_c_357_n 0.0565039f $X=1.75 $Y=2.035 $X2=0 $Y2=0
cc_115 N_A_83_270#_c_118_p N_VPWR_c_357_n 0.0119464f $X=0.785 $Y=2.035 $X2=0
+ $Y2=0
cc_116 N_A_83_270#_c_81_n N_VPWR_c_357_n 0.0203312f $X=1.915 $Y=2.13 $X2=0 $Y2=0
cc_117 N_A_83_270#_M1000_g N_VPWR_c_360_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A_83_270#_c_81_n N_VPWR_c_361_n 0.00832525f $X=1.915 $Y=2.13 $X2=0
+ $Y2=0
cc_119 N_A_83_270#_M1000_g N_VPWR_c_356_n 0.00990469f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_120 N_A_83_270#_c_81_n N_VPWR_c_356_n 0.0109296f $X=1.915 $Y=2.13 $X2=0 $Y2=0
cc_121 N_A_83_270#_c_73_n N_VGND_M1010_d 0.00188126f $X=0.62 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_122 N_A_83_270#_M1010_g N_VGND_c_403_n 0.0148187f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_123 N_A_83_270#_c_73_n N_VGND_c_403_n 0.0166905f $X=0.62 $Y=1.515 $X2=0 $Y2=0
cc_124 N_A_83_270#_c_74_n N_VGND_c_403_n 7.62615e-19 $X=0.62 $Y=1.515 $X2=0
+ $Y2=0
cc_125 N_A_83_270#_c_75_n N_VGND_c_403_n 0.0131435f $X=1.175 $Y=1.195 $X2=0
+ $Y2=0
cc_126 N_A_83_270#_c_76_n N_VGND_c_403_n 0.0403642f $X=1.34 $Y=0.515 $X2=0 $Y2=0
cc_127 N_A_83_270#_c_76_n N_VGND_c_406_n 0.0145639f $X=1.34 $Y=0.515 $X2=0 $Y2=0
cc_128 N_A_83_270#_M1010_g N_VGND_c_408_n 0.00383152f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_129 N_A_83_270#_M1010_g N_VGND_c_411_n 0.00761198f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_130 N_A_83_270#_c_76_n N_VGND_c_411_n 0.0119984f $X=1.34 $Y=0.515 $X2=0 $Y2=0
cc_131 N_A_83_270#_c_76_n N_A_326_74#_c_459_n 0.0195517f $X=1.34 $Y=0.515 $X2=0
+ $Y2=0
cc_132 N_A_83_270#_c_76_n N_A_326_74#_c_461_n 0.00682867f $X=1.34 $Y=0.515 $X2=0
+ $Y2=0
cc_133 N_B1_M1004_g N_A4_M1001_g 0.0191404f $X=1.555 $Y=0.69 $X2=0 $Y2=0
cc_134 N_B1_M1004_g N_A4_c_181_n 0.0177663f $X=1.555 $Y=0.69 $X2=0 $Y2=0
cc_135 N_B1_c_145_n N_A4_c_181_n 2.39091e-19 $X=1.415 $Y=1.615 $X2=0 $Y2=0
cc_136 N_B1_c_144_n N_A4_M1003_g 0.0320004f $X=1.605 $Y=1.91 $X2=0 $Y2=0
cc_137 N_B1_c_145_n N_A4_M1003_g 2.41039e-19 $X=1.415 $Y=1.615 $X2=0 $Y2=0
cc_138 N_B1_M1004_g N_A4_c_183_n 0.00168307f $X=1.555 $Y=0.69 $X2=0 $Y2=0
cc_139 N_B1_c_144_n N_A4_c_183_n 0.00235244f $X=1.605 $Y=1.91 $X2=0 $Y2=0
cc_140 N_B1_c_145_n N_A4_c_183_n 0.0180089f $X=1.415 $Y=1.615 $X2=0 $Y2=0
cc_141 N_B1_c_144_n N_VPWR_c_357_n 0.0192112f $X=1.605 $Y=1.91 $X2=0 $Y2=0
cc_142 N_B1_c_144_n N_VPWR_c_361_n 0.00499552f $X=1.605 $Y=1.91 $X2=0 $Y2=0
cc_143 N_B1_c_144_n N_VPWR_c_356_n 0.00524041f $X=1.605 $Y=1.91 $X2=0 $Y2=0
cc_144 N_B1_M1004_g N_VGND_c_403_n 0.00391465f $X=1.555 $Y=0.69 $X2=0 $Y2=0
cc_145 N_B1_M1004_g N_VGND_c_406_n 0.00434272f $X=1.555 $Y=0.69 $X2=0 $Y2=0
cc_146 N_B1_M1004_g N_VGND_c_411_n 0.0082698f $X=1.555 $Y=0.69 $X2=0 $Y2=0
cc_147 N_B1_M1004_g N_A_326_74#_c_459_n 0.00266933f $X=1.555 $Y=0.69 $X2=0 $Y2=0
cc_148 N_B1_M1004_g N_A_326_74#_c_461_n 9.23518e-19 $X=1.555 $Y=0.69 $X2=0 $Y2=0
cc_149 N_A4_M1003_g N_A3_M1007_g 0.0441463f $X=2.14 $Y=2.4 $X2=0 $Y2=0
cc_150 N_A4_M1001_g N_A3_M1011_g 0.0230092f $X=2.055 $Y=0.69 $X2=0 $Y2=0
cc_151 N_A4_c_181_n N_A3_M1011_g 9.08436e-19 $X=2.14 $Y=1.52 $X2=0 $Y2=0
cc_152 N_A4_c_183_n N_A3_M1011_g 6.6431e-19 $X=2.035 $Y=1.355 $X2=0 $Y2=0
cc_153 N_A4_c_181_n N_A3_c_227_n 0.0509565f $X=2.14 $Y=1.52 $X2=0 $Y2=0
cc_154 N_A4_c_183_n N_A3_c_227_n 0.00342973f $X=2.035 $Y=1.355 $X2=0 $Y2=0
cc_155 N_A4_c_181_n N_A3_c_228_n 6.49186e-19 $X=2.14 $Y=1.52 $X2=0 $Y2=0
cc_156 N_A4_M1003_g N_A3_c_228_n 0.00466828f $X=2.14 $Y=2.4 $X2=0 $Y2=0
cc_157 N_A4_c_183_n N_A3_c_228_n 0.0406201f $X=2.035 $Y=1.355 $X2=0 $Y2=0
cc_158 N_A4_M1003_g N_VPWR_c_357_n 0.00452705f $X=2.14 $Y=2.4 $X2=0 $Y2=0
cc_159 N_A4_M1003_g N_VPWR_c_361_n 0.00524256f $X=2.14 $Y=2.4 $X2=0 $Y2=0
cc_160 N_A4_M1003_g N_VPWR_c_356_n 0.00992373f $X=2.14 $Y=2.4 $X2=0 $Y2=0
cc_161 N_A4_M1001_g N_VGND_c_404_n 0.00525427f $X=2.055 $Y=0.69 $X2=0 $Y2=0
cc_162 N_A4_M1001_g N_VGND_c_406_n 0.00434272f $X=2.055 $Y=0.69 $X2=0 $Y2=0
cc_163 N_A4_M1001_g N_VGND_c_411_n 0.00448875f $X=2.055 $Y=0.69 $X2=0 $Y2=0
cc_164 N_A4_M1001_g N_A_326_74#_c_459_n 0.00731128f $X=2.055 $Y=0.69 $X2=0 $Y2=0
cc_165 N_A4_M1001_g N_A_326_74#_c_460_n 0.00920125f $X=2.055 $Y=0.69 $X2=0 $Y2=0
cc_166 N_A4_c_181_n N_A_326_74#_c_460_n 6.2263e-19 $X=2.14 $Y=1.52 $X2=0 $Y2=0
cc_167 N_A4_c_183_n N_A_326_74#_c_460_n 0.0210835f $X=2.035 $Y=1.355 $X2=0 $Y2=0
cc_168 N_A4_M1001_g N_A_326_74#_c_461_n 8.39937e-19 $X=2.055 $Y=0.69 $X2=0 $Y2=0
cc_169 N_A4_c_181_n N_A_326_74#_c_461_n 8.57327e-19 $X=2.14 $Y=1.52 $X2=0 $Y2=0
cc_170 N_A4_c_183_n N_A_326_74#_c_461_n 0.0116993f $X=2.035 $Y=1.355 $X2=0 $Y2=0
cc_171 N_A4_M1001_g N_A_326_74#_c_462_n 5.97046e-19 $X=2.055 $Y=0.69 $X2=0 $Y2=0
cc_172 N_A3_M1011_g N_A2_M1006_g 0.0222036f $X=2.625 $Y=0.69 $X2=0 $Y2=0
cc_173 N_A3_c_227_n N_A2_M1006_g 0.0177025f $X=2.635 $Y=1.385 $X2=0 $Y2=0
cc_174 N_A3_c_228_n N_A2_M1006_g 5.15832e-19 $X=2.635 $Y=1.385 $X2=0 $Y2=0
cc_175 N_A3_M1007_g N_A2_c_271_n 0.0462577f $X=2.56 $Y=2.4 $X2=0 $Y2=0
cc_176 N_A3_c_228_n N_A2_c_271_n 0.00518295f $X=2.635 $Y=1.385 $X2=0 $Y2=0
cc_177 N_A3_M1007_g N_A2_c_272_n 0.00156648f $X=2.56 $Y=2.4 $X2=0 $Y2=0
cc_178 N_A3_c_227_n N_A2_c_272_n 0.00153722f $X=2.635 $Y=1.385 $X2=0 $Y2=0
cc_179 N_A3_c_228_n N_A2_c_272_n 0.0752928f $X=2.635 $Y=1.385 $X2=0 $Y2=0
cc_180 N_A3_M1007_g N_VPWR_c_361_n 0.00365007f $X=2.56 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A3_c_228_n N_VPWR_c_361_n 0.00925382f $X=2.635 $Y=1.385 $X2=0 $Y2=0
cc_182 N_A3_M1007_g N_VPWR_c_356_n 0.00444515f $X=2.56 $Y=2.4 $X2=0 $Y2=0
cc_183 N_A3_c_228_n N_VPWR_c_356_n 0.0105443f $X=2.635 $Y=1.385 $X2=0 $Y2=0
cc_184 N_A3_c_228_n A_530_368# 0.0111776f $X=2.635 $Y=1.385 $X2=-0.19 $Y2=-0.245
cc_185 N_A3_M1011_g N_VGND_c_404_n 0.00387235f $X=2.625 $Y=0.69 $X2=0 $Y2=0
cc_186 N_A3_M1011_g N_VGND_c_405_n 4.25277e-19 $X=2.625 $Y=0.69 $X2=0 $Y2=0
cc_187 N_A3_M1011_g N_VGND_c_409_n 0.00434272f $X=2.625 $Y=0.69 $X2=0 $Y2=0
cc_188 N_A3_M1011_g N_VGND_c_411_n 0.00448792f $X=2.625 $Y=0.69 $X2=0 $Y2=0
cc_189 N_A3_M1011_g N_A_326_74#_c_459_n 5.97046e-19 $X=2.625 $Y=0.69 $X2=0 $Y2=0
cc_190 N_A3_M1011_g N_A_326_74#_c_460_n 0.00935164f $X=2.625 $Y=0.69 $X2=0 $Y2=0
cc_191 N_A3_c_227_n N_A_326_74#_c_460_n 5.31095e-19 $X=2.635 $Y=1.385 $X2=0
+ $Y2=0
cc_192 N_A3_c_228_n N_A_326_74#_c_460_n 0.0139058f $X=2.635 $Y=1.385 $X2=0 $Y2=0
cc_193 N_A3_M1011_g N_A_326_74#_c_462_n 0.00730737f $X=2.625 $Y=0.69 $X2=0 $Y2=0
cc_194 N_A3_M1011_g N_A_326_74#_c_465_n 8.85434e-19 $X=2.625 $Y=0.69 $X2=0 $Y2=0
cc_195 N_A3_c_227_n N_A_326_74#_c_465_n 7.62276e-19 $X=2.635 $Y=1.385 $X2=0
+ $Y2=0
cc_196 N_A3_c_228_n N_A_326_74#_c_465_n 0.00964811f $X=2.635 $Y=1.385 $X2=0
+ $Y2=0
cc_197 N_A2_M1006_g N_A1_M1008_g 0.0200135f $X=3.115 $Y=0.69 $X2=0 $Y2=0
cc_198 N_A2_c_271_n N_A1_M1008_g 0.00172681f $X=3.205 $Y=1.465 $X2=0 $Y2=0
cc_199 N_A2_c_272_n N_A1_M1008_g 2.87867e-19 $X=3.205 $Y=1.465 $X2=0 $Y2=0
cc_200 N_A2_M1005_g N_A1_c_308_n 0.0398379f $X=3.13 $Y=2.4 $X2=0 $Y2=0
cc_201 N_A2_c_271_n N_A1_c_308_n 0.0144946f $X=3.205 $Y=1.465 $X2=0 $Y2=0
cc_202 N_A2_c_272_n N_A1_c_308_n 0.0138201f $X=3.205 $Y=1.465 $X2=0 $Y2=0
cc_203 N_A2_M1005_g N_A1_c_309_n 5.363e-19 $X=3.13 $Y=2.4 $X2=0 $Y2=0
cc_204 N_A2_c_271_n N_A1_c_309_n 0.00102824f $X=3.205 $Y=1.465 $X2=0 $Y2=0
cc_205 N_A2_c_272_n N_A1_c_309_n 0.0497024f $X=3.205 $Y=1.465 $X2=0 $Y2=0
cc_206 N_A2_M1005_g N_VPWR_c_359_n 0.00140744f $X=3.13 $Y=2.4 $X2=0 $Y2=0
cc_207 N_A2_c_272_n N_VPWR_c_359_n 0.0240626f $X=3.205 $Y=1.465 $X2=0 $Y2=0
cc_208 N_A2_M1005_g N_VPWR_c_361_n 0.00363952f $X=3.13 $Y=2.4 $X2=0 $Y2=0
cc_209 N_A2_c_272_n N_VPWR_c_361_n 0.00985991f $X=3.205 $Y=1.465 $X2=0 $Y2=0
cc_210 N_A2_M1005_g N_VPWR_c_356_n 0.00446867f $X=3.13 $Y=2.4 $X2=0 $Y2=0
cc_211 N_A2_c_272_n N_VPWR_c_356_n 0.0117596f $X=3.205 $Y=1.465 $X2=0 $Y2=0
cc_212 N_A2_c_272_n A_644_368# 0.0137905f $X=3.205 $Y=1.465 $X2=-0.19 $Y2=-0.245
cc_213 N_A2_M1006_g N_VGND_c_405_n 0.0136443f $X=3.115 $Y=0.69 $X2=0 $Y2=0
cc_214 N_A2_M1006_g N_VGND_c_409_n 0.00413917f $X=3.115 $Y=0.69 $X2=0 $Y2=0
cc_215 N_A2_M1006_g N_VGND_c_411_n 0.00417193f $X=3.115 $Y=0.69 $X2=0 $Y2=0
cc_216 N_A2_M1006_g N_A_326_74#_c_462_n 0.00265992f $X=3.115 $Y=0.69 $X2=0 $Y2=0
cc_217 N_A2_M1006_g N_A_326_74#_c_463_n 0.0138853f $X=3.115 $Y=0.69 $X2=0 $Y2=0
cc_218 N_A2_c_271_n N_A_326_74#_c_463_n 0.00113397f $X=3.205 $Y=1.465 $X2=0
+ $Y2=0
cc_219 N_A2_c_272_n N_A_326_74#_c_463_n 0.0195066f $X=3.205 $Y=1.465 $X2=0 $Y2=0
cc_220 N_A2_M1006_g N_A_326_74#_c_464_n 9.0724e-19 $X=3.115 $Y=0.69 $X2=0 $Y2=0
cc_221 N_A1_c_309_n N_VPWR_M1009_d 0.00726344f $X=3.775 $Y=1.515 $X2=0 $Y2=0
cc_222 N_A1_M1009_g N_VPWR_c_359_n 0.0178955f $X=3.7 $Y=2.4 $X2=0 $Y2=0
cc_223 N_A1_c_308_n N_VPWR_c_359_n 3.89265e-19 $X=3.775 $Y=1.515 $X2=0 $Y2=0
cc_224 N_A1_c_309_n N_VPWR_c_359_n 0.0337305f $X=3.775 $Y=1.515 $X2=0 $Y2=0
cc_225 N_A1_M1009_g N_VPWR_c_361_n 0.00460063f $X=3.7 $Y=2.4 $X2=0 $Y2=0
cc_226 N_A1_M1009_g N_VPWR_c_356_n 0.00909693f $X=3.7 $Y=2.4 $X2=0 $Y2=0
cc_227 N_A1_M1008_g N_VGND_c_405_n 0.00623438f $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_228 N_A1_M1008_g N_VGND_c_410_n 0.00434272f $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_229 N_A1_M1008_g N_VGND_c_411_n 0.00452716f $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_230 N_A1_M1008_g N_A_326_74#_c_463_n 0.0119089f $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_231 N_A1_c_308_n N_A_326_74#_c_463_n 0.00113236f $X=3.775 $Y=1.515 $X2=0
+ $Y2=0
cc_232 N_A1_c_309_n N_A_326_74#_c_463_n 0.0310954f $X=3.775 $Y=1.515 $X2=0 $Y2=0
cc_233 N_A1_M1008_g N_A_326_74#_c_464_n 0.00786806f $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_234 X N_VPWR_c_357_n 0.026735f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_235 X N_VPWR_c_360_n 0.0145564f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_236 X N_VPWR_c_356_n 0.0119772f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_237 N_X_c_335_n N_VGND_c_403_n 0.023562f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_238 N_X_c_335_n N_VGND_c_408_n 0.0115122f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_239 N_X_c_335_n N_VGND_c_411_n 0.0095288f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_240 N_VGND_c_404_n N_A_326_74#_c_459_n 0.0131729f $X=2.34 $Y=0.515 $X2=0
+ $Y2=0
cc_241 N_VGND_c_406_n N_A_326_74#_c_459_n 0.0145482f $X=2.175 $Y=0 $X2=0 $Y2=0
cc_242 N_VGND_c_411_n N_A_326_74#_c_459_n 0.0119922f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_243 N_VGND_M1001_d N_A_326_74#_c_460_n 0.00373913f $X=2.13 $Y=0.37 $X2=0
+ $Y2=0
cc_244 N_VGND_c_404_n N_A_326_74#_c_460_n 0.0243707f $X=2.34 $Y=0.515 $X2=0
+ $Y2=0
cc_245 N_VGND_c_411_n N_A_326_74#_c_460_n 0.0109408f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_246 N_VGND_c_404_n N_A_326_74#_c_462_n 0.0131729f $X=2.34 $Y=0.515 $X2=0
+ $Y2=0
cc_247 N_VGND_c_405_n N_A_326_74#_c_462_n 0.0141032f $X=3.44 $Y=0.515 $X2=0
+ $Y2=0
cc_248 N_VGND_c_409_n N_A_326_74#_c_462_n 0.0145482f $X=3.175 $Y=0 $X2=0 $Y2=0
cc_249 N_VGND_c_411_n N_A_326_74#_c_462_n 0.0119922f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_250 N_VGND_M1006_d N_A_326_74#_c_463_n 0.00644036f $X=3.19 $Y=0.37 $X2=0
+ $Y2=0
cc_251 N_VGND_c_405_n N_A_326_74#_c_463_n 0.0365648f $X=3.44 $Y=0.515 $X2=0
+ $Y2=0
cc_252 N_VGND_c_411_n N_A_326_74#_c_463_n 0.0114864f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_253 N_VGND_c_405_n N_A_326_74#_c_464_n 0.0132315f $X=3.44 $Y=0.515 $X2=0
+ $Y2=0
cc_254 N_VGND_c_410_n N_A_326_74#_c_464_n 0.0145639f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_255 N_VGND_c_411_n N_A_326_74#_c_464_n 0.0119984f $X=4.08 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__o32a_4.spice
* Created: Wed Sep  2 12:26:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o32a_4.pex.spice"
.subckt sky130_fd_sc_ms__o32a_4  VNB VPB B1 B2 A3 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1015 N_X_M1015_d N_A_83_256#_M1015_g N_VGND_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2543 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.3
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1020 N_X_M1015_d N_A_83_256#_M1020_g N_VGND_M1020_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.7
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1024 N_X_M1024_d N_A_83_256#_M1024_g N_VGND_M1020_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.14985 AS=0.1554 PD=1.145 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.3
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1027 N_X_M1024_d N_A_83_256#_M1027_g N_VGND_M1027_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.14985 AS=0.2109 PD=1.145 PS=2.05 NRD=20.268 NRS=0 M=1 R=4.93333
+ SA=75001.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_A_83_256#_M1010_d N_B1_M1010_g N_A_564_74#_M1010_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75004.7 A=0.096 P=1.58 MULT=1
MM1025 N_A_83_256#_M1010_d N_B1_M1025_g N_A_564_74#_M1025_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75000.6 SB=75004.3 A=0.096 P=1.58 MULT=1
MM1021 N_A_564_74#_M1025_s N_B2_M1021_g N_A_83_256#_M1021_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.112 AS=0.112 PD=0.99 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75001.1 SB=75003.8 A=0.096 P=1.58 MULT=1
MM1022 N_A_564_74#_M1022_d N_B2_M1022_g N_A_83_256#_M1021_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1216 AS=0.112 PD=1.02 PS=0.99 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75001.6 SB=75003.3 A=0.096 P=1.58 MULT=1
MM1002 N_A_564_74#_M1022_d N_A3_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1216 AS=0.1184 PD=1.02 PS=1.01 NRD=5.616 NRS=7.488 M=1 R=4.26667
+ SA=75002.2 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1012 N_A_564_74#_M1012_d N_A3_M1012_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.096 AS=0.1184 PD=0.94 PS=1.01 NRD=3.744 NRS=9.372 M=1 R=4.26667
+ SA=75002.7 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1004 N_A_564_74#_M1012_d N_A2_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.096 AS=0.112 PD=0.94 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75003.1
+ SB=75001.8 A=0.096 P=1.58 MULT=1
MM1007 N_A_564_74#_M1007_d N_A2_M1007_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75003.6
+ SB=75001.3 A=0.096 P=1.58 MULT=1
MM1005 N_VGND_M1005_d N_A1_M1005_g N_A_564_74#_M1007_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.152 AS=0.0896 PD=1.115 PS=0.92 NRD=17.808 NRS=0 M=1 R=4.26667 SA=75004.1
+ SB=75000.8 A=0.096 P=1.58 MULT=1
MM1014 N_VGND_M1005_d N_A1_M1014_g N_A_564_74#_M1014_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.152 AS=0.1824 PD=1.115 PS=1.85 NRD=18.744 NRS=0 M=1 R=4.26667 SA=75004.7
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1003 N_VPWR_M1003_d N_A_83_256#_M1003_g N_X_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003.6 A=0.2016 P=2.6 MULT=1
MM1006 N_VPWR_M1006_d N_A_83_256#_M1006_g N_X_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90003.1 A=0.2016 P=2.6 MULT=1
MM1008 N_VPWR_M1006_d N_A_83_256#_M1008_g N_X_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.2184 PD=1.44 PS=1.51 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.1
+ SB=90002.6 A=0.2016 P=2.6 MULT=1
MM1009 N_VPWR_M1009_d N_A_83_256#_M1009_g N_X_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.222204 AS=0.2184 PD=1.59547 PS=1.51 NRD=0 NRS=11.426 M=1 R=6.22222
+ SA=90001.7 SB=90002.1 A=0.2016 P=2.6 MULT=1
MM1018 N_A_537_388#_M1018_d N_B1_M1018_g N_VPWR_M1009_d VPB PSHORT L=0.18 W=1
+ AD=0.205 AS=0.198396 PD=1.41 PS=1.42453 NRD=12.7853 NRS=22.6353 M=1 R=5.55556
+ SA=90002.3 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1016 N_A_83_256#_M1016_d N_B2_M1016_g N_A_537_388#_M1018_d VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.205 PD=1.27 PS=1.41 NRD=0 NRS=12.7853 M=1 R=5.55556
+ SA=90002.9 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1019 N_A_83_256#_M1016_d N_B2_M1019_g N_A_537_388#_M1019_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90003.3
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1023 N_A_537_388#_M1019_s N_B1_M1023_g N_VPWR_M1023_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.33 PD=1.27 PS=2.66 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90003.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1000 N_A_961_392#_M1000_d N_A3_M1000_g N_A_83_256#_M1000_s VPB PSHORT L=0.18
+ W=1 AD=0.28 AS=0.145 PD=2.56 PS=1.29 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90002.7 A=0.18 P=2.36 MULT=1
MM1017 N_A_961_392#_M1017_d N_A3_M1017_g N_A_83_256#_M1000_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.145 PD=1.27 PS=1.29 NRD=0 NRS=2.9353 M=1 R=5.55556
+ SA=90000.7 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1001 N_A_1237_392#_M1001_d N_A2_M1001_g N_A_961_392#_M1017_d VPB PSHORT L=0.18
+ W=1 AD=0.23 AS=0.135 PD=1.46 PS=1.27 NRD=17.73 NRS=0 M=1 R=5.55556 SA=90001.1
+ SB=90001.7 A=0.18 P=2.36 MULT=1
MM1011 N_A_1237_392#_M1001_d N_A1_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1
+ AD=0.23 AS=0.145 PD=1.46 PS=1.29 NRD=17.73 NRS=0.9653 M=1 R=5.55556 SA=90001.7
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1026 N_A_1237_392#_M1026_d N_A1_M1026_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.145 PD=1.27 PS=1.29 NRD=0 NRS=0.9653 M=1 R=5.55556 SA=90002.2
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1013 N_A_1237_392#_M1026_d N_A2_M1013_g N_A_961_392#_M1013_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556 SA=90002.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_ms__o32a_4.pxi.spice"
*
.ends
*
*

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__o211ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__o211ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.350000 1.795000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.250400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 4.195000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.847200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 5.635000 1.780000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.847200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.870000 1.350000 7.075000 1.780000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.780800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.430000 1.950000 8.035000 2.120000 ;
        RECT 2.430000 2.120000 2.760000 2.735000 ;
        RECT 3.380000 2.120000 3.710000 2.735000 ;
        RECT 4.940000 2.120000 5.270000 2.980000 ;
        RECT 5.940000 2.120000 6.270000 2.980000 ;
        RECT 6.505000 0.595000 6.675000 1.010000 ;
        RECT 6.505000 1.010000 7.545000 1.180000 ;
        RECT 7.365000 0.595000 7.545000 1.010000 ;
        RECT 7.365000 1.180000 7.545000 1.550000 ;
        RECT 7.365000 1.550000 8.035000 1.950000 ;
        RECT 7.545000 2.120000 8.035000 2.890000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.115000  0.350000 0.445000 1.010000 ;
      RECT 0.115000  1.010000 5.765000 1.180000 ;
      RECT 0.130000  1.950000 2.260000 2.120000 ;
      RECT 0.130000  2.120000 0.460000 2.980000 ;
      RECT 0.615000  0.085000 0.945000 0.840000 ;
      RECT 0.660000  2.290000 0.830000 3.245000 ;
      RECT 1.030000  2.120000 1.360000 2.980000 ;
      RECT 1.125000  0.350000 1.375000 1.010000 ;
      RECT 1.545000  0.085000 1.875000 0.840000 ;
      RECT 1.560000  2.290000 1.730000 3.245000 ;
      RECT 1.930000  2.120000 2.260000 2.905000 ;
      RECT 1.930000  2.905000 4.210000 3.075000 ;
      RECT 2.055000  0.350000 2.225000 1.010000 ;
      RECT 2.405000  0.085000 2.735000 0.840000 ;
      RECT 2.915000  0.350000 3.085000 1.010000 ;
      RECT 2.960000  2.290000 3.210000 2.905000 ;
      RECT 3.265000  0.085000 3.595000 0.840000 ;
      RECT 3.795000  0.350000 3.965000 0.820000 ;
      RECT 3.795000  0.820000 4.905000 1.010000 ;
      RECT 3.880000  2.290000 4.210000 2.905000 ;
      RECT 4.145000  0.255000 8.045000 0.425000 ;
      RECT 4.145000  0.425000 5.255000 0.650000 ;
      RECT 4.440000  2.290000 4.770000 3.245000 ;
      RECT 5.085000  0.650000 5.255000 0.840000 ;
      RECT 5.435000  0.595000 5.765000 1.010000 ;
      RECT 5.440000  2.290000 5.770000 3.245000 ;
      RECT 5.995000  0.425000 6.325000 1.180000 ;
      RECT 6.440000  2.290000 7.290000 3.245000 ;
      RECT 6.855000  0.425000 7.185000 0.840000 ;
      RECT 7.715000  0.425000 8.045000 1.180000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_ms__o211ai_4
END LIBRARY

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR a_86_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 a_492_125# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X2 a_86_260# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X3 a_971_392# A2 a_699_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X4 VGND A3 a_492_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 a_699_392# A3 a_86_260# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X6 a_86_260# B1 a_492_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X7 a_699_392# A2 a_971_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X8 VPWR a_86_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X9 a_492_125# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X10 a_971_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X11 VGND a_86_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 a_492_125# B1 a_86_260# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 VGND A2 a_492_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X14 VPWR A1 a_971_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X15 VPWR B1 a_86_260# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X16 X a_86_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 VGND a_86_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 X a_86_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_86_260# A3 a_699_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X20 X a_86_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X21 X a_86_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X22 a_492_125# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X23 VGND A1 a_492_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends

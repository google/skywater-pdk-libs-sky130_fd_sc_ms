* File: sky130_fd_sc_ms__a22o_4.pxi.spice
* Created: Wed Sep  2 11:53:19 2020
* 
x_PM_SKY130_FD_SC_MS__A22O_4%A_95_306# N_A_95_306#_M1001_d N_A_95_306#_M1003_d
+ N_A_95_306#_M1008_d N_A_95_306#_M1014_s N_A_95_306#_M1009_g
+ N_A_95_306#_c_131_n N_A_95_306#_c_132_n N_A_95_306#_M1010_g
+ N_A_95_306#_c_133_n N_A_95_306#_M1005_g N_A_95_306#_M1011_g
+ N_A_95_306#_c_135_n N_A_95_306#_M1007_g N_A_95_306#_M1015_g
+ N_A_95_306#_c_136_n N_A_95_306#_M1017_g N_A_95_306#_c_137_n
+ N_A_95_306#_M1020_g N_A_95_306#_c_138_n N_A_95_306#_c_139_n
+ N_A_95_306#_c_221_p N_A_95_306#_c_140_n N_A_95_306#_c_157_n
+ N_A_95_306#_c_158_n N_A_95_306#_c_159_n N_A_95_306#_c_160_n
+ N_A_95_306#_c_161_n N_A_95_306#_c_141_n N_A_95_306#_c_142_n
+ N_A_95_306#_c_143_n N_A_95_306#_c_144_n N_A_95_306#_c_145_n
+ N_A_95_306#_c_146_n PM_SKY130_FD_SC_MS__A22O_4%A_95_306#
x_PM_SKY130_FD_SC_MS__A22O_4%B2 N_B2_M1008_g N_B2_M1000_g N_B2_M1019_g
+ N_B2_M1022_g N_B2_c_328_n N_B2_c_329_n N_B2_c_321_n N_B2_c_322_n N_B2_c_323_n
+ N_B2_c_324_n N_B2_c_325_n N_B2_c_358_n B2 B2 N_B2_c_334_n
+ PM_SKY130_FD_SC_MS__A22O_4%B2
x_PM_SKY130_FD_SC_MS__A22O_4%B1 N_B1_M1012_g N_B1_M1001_g N_B1_M1018_g
+ N_B1_M1014_g B1 N_B1_c_419_n PM_SKY130_FD_SC_MS__A22O_4%B1
x_PM_SKY130_FD_SC_MS__A22O_4%A1 N_A1_M1004_g N_A1_M1003_g N_A1_M1021_g
+ N_A1_M1013_g A1 A1 N_A1_c_471_n PM_SKY130_FD_SC_MS__A22O_4%A1
x_PM_SKY130_FD_SC_MS__A22O_4%A2 N_A2_M1006_g N_A2_M1002_g N_A2_c_520_n
+ N_A2_c_521_n N_A2_M1016_g N_A2_M1023_g N_A2_c_524_n A2 N_A2_c_526_n
+ PM_SKY130_FD_SC_MS__A22O_4%A2
x_PM_SKY130_FD_SC_MS__A22O_4%VPWR N_VPWR_M1009_s N_VPWR_M1010_s N_VPWR_M1015_s
+ N_VPWR_M1006_s N_VPWR_M1021_d N_VPWR_c_582_n N_VPWR_c_583_n N_VPWR_c_584_n
+ N_VPWR_c_585_n N_VPWR_c_586_n N_VPWR_c_587_n N_VPWR_c_588_n N_VPWR_c_589_n
+ VPWR N_VPWR_c_590_n N_VPWR_c_591_n N_VPWR_c_592_n N_VPWR_c_593_n
+ N_VPWR_c_581_n N_VPWR_c_595_n N_VPWR_c_596_n N_VPWR_c_597_n
+ PM_SKY130_FD_SC_MS__A22O_4%VPWR
x_PM_SKY130_FD_SC_MS__A22O_4%X N_X_M1005_d N_X_M1017_d N_X_M1009_d N_X_M1011_d
+ N_X_c_676_n N_X_c_671_n N_X_c_677_n N_X_c_692_n N_X_c_672_n N_X_c_673_n
+ N_X_c_704_n X X N_X_c_675_n PM_SKY130_FD_SC_MS__A22O_4%X
x_PM_SKY130_FD_SC_MS__A22O_4%A_555_392# N_A_555_392#_M1008_s
+ N_A_555_392#_M1012_d N_A_555_392#_M1019_s N_A_555_392#_M1004_s
+ N_A_555_392#_M1016_d N_A_555_392#_c_735_n N_A_555_392#_c_749_n
+ N_A_555_392#_c_736_n N_A_555_392#_c_791_n N_A_555_392#_c_737_n
+ N_A_555_392#_c_738_n N_A_555_392#_c_739_n N_A_555_392#_c_740_n
+ N_A_555_392#_c_741_n N_A_555_392#_c_754_n N_A_555_392#_c_742_n
+ N_A_555_392#_c_743_n PM_SKY130_FD_SC_MS__A22O_4%A_555_392#
x_PM_SKY130_FD_SC_MS__A22O_4%VGND N_VGND_M1005_s N_VGND_M1007_s N_VGND_M1020_s
+ N_VGND_M1022_s N_VGND_M1023_s N_VGND_c_809_n N_VGND_c_810_n N_VGND_c_811_n
+ N_VGND_c_812_n N_VGND_c_813_n N_VGND_c_814_n N_VGND_c_815_n N_VGND_c_816_n
+ N_VGND_c_817_n N_VGND_c_818_n N_VGND_c_819_n N_VGND_c_820_n N_VGND_c_821_n
+ N_VGND_c_822_n VGND N_VGND_c_823_n N_VGND_c_824_n N_VGND_c_825_n
+ PM_SKY130_FD_SC_MS__A22O_4%VGND
x_PM_SKY130_FD_SC_MS__A22O_4%A_645_120# N_A_645_120#_M1000_d
+ N_A_645_120#_M1018_s N_A_645_120#_c_897_n N_A_645_120#_c_898_n
+ PM_SKY130_FD_SC_MS__A22O_4%A_645_120#
x_PM_SKY130_FD_SC_MS__A22O_4%A_1064_123# N_A_1064_123#_M1002_d
+ N_A_1064_123#_M1013_s N_A_1064_123#_c_917_n N_A_1064_123#_c_914_n
+ N_A_1064_123#_c_915_n PM_SKY130_FD_SC_MS__A22O_4%A_1064_123#
cc_1 VNB N_A_95_306#_c_131_n 0.0111784f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.605
cc_2 VNB N_A_95_306#_c_132_n 0.0142618f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.605
cc_3 VNB N_A_95_306#_c_133_n 0.00733251f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=1.605
cc_4 VNB N_A_95_306#_M1005_g 0.0278837f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.87
cc_5 VNB N_A_95_306#_c_135_n 0.0153169f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.35
cc_6 VNB N_A_95_306#_c_136_n 0.0162201f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=1.35
cc_7 VNB N_A_95_306#_c_137_n 0.0172571f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.35
cc_8 VNB N_A_95_306#_c_138_n 0.00762043f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.605
cc_9 VNB N_A_95_306#_c_139_n 0.00479297f $X=-0.19 $Y=-0.245 $X2=1.417 $Y2=1.605
cc_10 VNB N_A_95_306#_c_140_n 0.00322996f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=1.68
cc_11 VNB N_A_95_306#_c_141_n 0.00618103f $X=-0.19 $Y=-0.245 $X2=3.63 $Y2=1.132
cc_12 VNB N_A_95_306#_c_142_n 0.00304687f $X=-0.19 $Y=-0.245 $X2=3.96 $Y2=1.132
cc_13 VNB N_A_95_306#_c_143_n 0.00229391f $X=-0.19 $Y=-0.245 $X2=5.89 $Y2=1.105
cc_14 VNB N_A_95_306#_c_144_n 0.0141457f $X=-0.19 $Y=-0.245 $X2=5.725 $Y2=1.145
cc_15 VNB N_A_95_306#_c_145_n 0.0039374f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.515
cc_16 VNB N_A_95_306#_c_146_n 0.0443893f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.515
cc_17 VNB N_B2_M1000_g 0.02243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B2_M1022_g 0.0230208f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.4
cc_19 VNB N_B2_c_321_n 7.59216e-19 $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=2.4
cc_20 VNB N_B2_c_322_n 0.0037501f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=1.605
cc_21 VNB N_B2_c_323_n 0.0165844f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=1.605
cc_22 VNB N_B2_c_324_n 0.0184476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B2_c_325_n 0.00181489f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=2.4
cc_24 VNB N_B1_M1001_g 0.0210564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B1_M1018_g 0.0217123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB B1 8.16208e-19 $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.605
cc_27 VNB N_B1_c_419_n 0.0252562f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.87
cc_28 VNB N_A1_M1003_g 0.0194032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A1_M1013_g 0.0193298f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=2.4
cc_30 VNB A1 0.00392757f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.605
cc_31 VNB N_A1_c_471_n 0.0266595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A2_M1006_g 0.0109566f $X=-0.19 $Y=-0.245 $X2=3.215 $Y2=1.96
cc_33 VNB N_A2_M1002_g 0.0114364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A2_c_520_n 0.0902248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A2_c_521_n 0.00932321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A2_M1016_g 0.0203142f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.68
cc_37 VNB N_A2_M1023_g 0.0330549f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.605
cc_38 VNB N_A2_c_524_n 0.0285318f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=2.4
cc_39 VNB A2 0.0131334f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=1.605
cc_40 VNB N_A2_c_526_n 0.0472248f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.87
cc_41 VNB N_VPWR_c_581_n 0.302998f $X=-0.19 $Y=-0.245 $X2=3.35 $Y2=2.867
cc_42 VNB N_X_c_671_n 0.00251264f $X=-0.19 $Y=-0.245 $X2=1.28 $Y2=1.605
cc_43 VNB N_X_c_672_n 0.00252589f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.35
cc_44 VNB N_X_c_673_n 0.00571544f $X=-0.19 $Y=-0.245 $X2=1.915 $Y2=1.68
cc_45 VNB X 0.0131314f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=0.87
cc_46 VNB N_X_c_675_n 0.0457248f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=0.87
cc_47 VNB N_VGND_c_809_n 0.0371369f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.605
cc_48 VNB N_VGND_c_810_n 0.00886349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_811_n 0.0176237f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.87
cc_50 VNB N_VGND_c_812_n 0.0172788f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=2.4
cc_51 VNB N_VGND_c_813_n 0.049564f $X=-0.19 $Y=-0.245 $X2=1.555 $Y2=1.605
cc_52 VNB N_VGND_c_814_n 0.0331697f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.87
cc_53 VNB N_VGND_c_815_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=1.915 $Y2=1.68
cc_54 VNB N_VGND_c_816_n 0.0178473f $X=-0.19 $Y=-0.245 $X2=1.915 $Y2=2.4
cc_55 VNB N_VGND_c_817_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_818_n 0.0178473f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=0.87
cc_57 VNB N_VGND_c_819_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=0.87
cc_58 VNB N_VGND_c_820_n 0.0112126f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.35
cc_59 VNB N_VGND_c_821_n 0.0480638f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=0.87
cc_60 VNB N_VGND_c_822_n 0.00528596f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=0.87
cc_61 VNB N_VGND_c_823_n 0.042264f $X=-0.19 $Y=-0.245 $X2=4.25 $Y2=2.78
cc_62 VNB N_VGND_c_824_n 0.442195f $X=-0.19 $Y=-0.245 $X2=3.795 $Y2=1.09
cc_63 VNB N_VGND_c_825_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=3.96 $Y2=1.132
cc_64 VNB N_A_645_120#_c_897_n 0.00288446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_645_120#_c_898_n 0.00740647f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.68
cc_66 VNB N_A_1064_123#_c_914_n 0.00186167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1064_123#_c_915_n 0.00325899f $X=-0.19 $Y=-0.245 $X2=0.565
+ $Y2=1.68
cc_68 VPB N_A_95_306#_M1009_g 0.027617f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=2.4
cc_69 VPB N_A_95_306#_c_131_n 0.00314639f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.605
cc_70 VPB N_A_95_306#_c_132_n 0.0014875f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.605
cc_71 VPB N_A_95_306#_M1010_g 0.0205586f $X=-0.19 $Y=1.66 $X2=1.015 $Y2=2.4
cc_72 VPB N_A_95_306#_c_133_n 0.00220943f $X=-0.19 $Y=1.66 $X2=1.28 $Y2=1.605
cc_73 VPB N_A_95_306#_M1011_g 0.0206261f $X=-0.19 $Y=1.66 $X2=1.465 $Y2=2.4
cc_74 VPB N_A_95_306#_M1015_g 0.0231187f $X=-0.19 $Y=1.66 $X2=1.915 $Y2=2.4
cc_75 VPB N_A_95_306#_c_138_n 3.82064e-19 $X=-0.19 $Y=1.66 $X2=1.015 $Y2=1.605
cc_76 VPB N_A_95_306#_c_139_n 7.12428e-19 $X=-0.19 $Y=1.66 $X2=1.417 $Y2=1.605
cc_77 VPB N_A_95_306#_c_140_n 0.00727707f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=1.68
cc_78 VPB N_A_95_306#_c_157_n 0.0252699f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=2.905
cc_79 VPB N_A_95_306#_c_158_n 0.00353271f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=2.99
cc_80 VPB N_A_95_306#_c_159_n 0.00457582f $X=-0.19 $Y=1.66 $X2=4.25 $Y2=2.78
cc_81 VPB N_A_95_306#_c_160_n 0.00834022f $X=-0.19 $Y=1.66 $X2=3.185 $Y2=2.867
cc_82 VPB N_A_95_306#_c_161_n 0.00195225f $X=-0.19 $Y=1.66 $X2=3.515 $Y2=2.867
cc_83 VPB N_A_95_306#_c_145_n 0.00215125f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.515
cc_84 VPB N_A_95_306#_c_146_n 0.0282315f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=1.515
cc_85 VPB N_B2_M1008_g 0.0254906f $X=-0.19 $Y=1.66 $X2=3.215 $Y2=1.96
cc_86 VPB N_B2_M1019_g 0.0243802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_B2_c_328_n 0.00175124f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.605
cc_88 VPB N_B2_c_329_n 0.00181541f $X=-0.19 $Y=1.66 $X2=1.015 $Y2=2.4
cc_89 VPB N_B2_c_322_n 0.0032539f $X=-0.19 $Y=1.66 $X2=1.28 $Y2=1.605
cc_90 VPB N_B2_c_323_n 0.0104799f $X=-0.19 $Y=1.66 $X2=1.105 $Y2=1.605
cc_91 VPB N_B2_c_324_n 0.0115696f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_B2_c_325_n 7.66814e-19 $X=-0.19 $Y=1.66 $X2=1.465 $Y2=2.4
cc_93 VPB N_B2_c_334_n 0.0056589f $X=-0.19 $Y=1.66 $X2=2.215 $Y2=0.87
cc_94 VPB N_B1_M1012_g 0.0226037f $X=-0.19 $Y=1.66 $X2=3.215 $Y2=1.96
cc_95 VPB N_B1_M1014_g 0.0222515f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=2.4
cc_96 VPB B1 6.39981e-19 $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.605
cc_97 VPB N_B1_c_419_n 0.0123219f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.87
cc_98 VPB N_A1_M1004_g 0.0249233f $X=-0.19 $Y=1.66 $X2=3.215 $Y2=1.96
cc_99 VPB N_A1_M1021_g 0.0219617f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB A1 0.00275828f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.605
cc_101 VPB N_A1_c_471_n 0.0156643f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A2_M1006_g 0.032509f $X=-0.19 $Y=1.66 $X2=3.215 $Y2=1.96
cc_103 VPB N_A2_M1016_g 0.0407804f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.68
cc_104 VPB N_VPWR_c_582_n 0.0139106f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_583_n 0.0508739f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.605
cc_106 VPB N_VPWR_c_584_n 0.00676446f $X=-0.19 $Y=1.66 $X2=1.105 $Y2=1.605
cc_107 VPB N_VPWR_c_585_n 0.0213173f $X=-0.19 $Y=1.66 $X2=1.465 $Y2=2.4
cc_108 VPB N_VPWR_c_586_n 0.00730495f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=0.87
cc_109 VPB N_VPWR_c_587_n 0.00335558f $X=-0.19 $Y=1.66 $X2=1.915 $Y2=2.4
cc_110 VPB N_VPWR_c_588_n 0.0175706f $X=-0.19 $Y=1.66 $X2=2.215 $Y2=0.87
cc_111 VPB N_VPWR_c_589_n 0.00601644f $X=-0.19 $Y=1.66 $X2=2.215 $Y2=0.87
cc_112 VPB N_VPWR_c_590_n 0.0164465f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=0.87
cc_113 VPB N_VPWR_c_591_n 0.0206041f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=1.68
cc_114 VPB N_VPWR_c_592_n 0.0676687f $X=-0.19 $Y=1.66 $X2=2.855 $Y2=1.18
cc_115 VPB N_VPWR_c_593_n 0.0235962f $X=-0.19 $Y=1.66 $X2=2.555 $Y2=1.515
cc_116 VPB N_VPWR_c_581_n 0.0952417f $X=-0.19 $Y=1.66 $X2=3.35 $Y2=2.867
cc_117 VPB N_VPWR_c_595_n 0.00458862f $X=-0.19 $Y=1.66 $X2=3.63 $Y2=1.132
cc_118 VPB N_VPWR_c_596_n 0.0047828f $X=-0.19 $Y=1.66 $X2=5.89 $Y2=1.105
cc_119 VPB N_VPWR_c_597_n 0.00893493f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=1.515
cc_120 VPB N_X_c_676_n 0.00453875f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=2.4
cc_121 VPB N_X_c_677_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.87
cc_122 VPB N_A_555_392#_c_735_n 0.00278896f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.605
cc_123 VPB N_A_555_392#_c_736_n 0.00408467f $X=-0.19 $Y=1.66 $X2=1.105 $Y2=1.605
cc_124 VPB N_A_555_392#_c_737_n 0.00754304f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_555_392#_c_738_n 0.00202354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_555_392#_c_739_n 0.00711489f $X=-0.19 $Y=1.66 $X2=1.555 $Y2=1.605
cc_127 VPB N_A_555_392#_c_740_n 0.0120216f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=0.87
cc_128 VPB N_A_555_392#_c_741_n 0.0345796f $X=-0.19 $Y=1.66 $X2=1.915 $Y2=1.68
cc_129 VPB N_A_555_392#_c_742_n 0.00252309f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=0.87
cc_130 VPB N_A_555_392#_c_743_n 0.00177335f $X=-0.19 $Y=1.66 $X2=1.417 $Y2=1.605
cc_131 N_A_95_306#_c_157_n N_B2_M1008_g 0.00665186f $X=2.56 $Y=2.905 $X2=0 $Y2=0
cc_132 N_A_95_306#_c_160_n N_B2_M1008_g 0.0102933f $X=3.185 $Y=2.867 $X2=0 $Y2=0
cc_133 N_A_95_306#_c_161_n N_B2_M1008_g 0.00678295f $X=3.515 $Y=2.867 $X2=0
+ $Y2=0
cc_134 N_A_95_306#_c_137_n N_B2_M1000_g 0.0233895f $X=2.645 $Y=1.35 $X2=0 $Y2=0
cc_135 N_A_95_306#_c_140_n N_B2_M1000_g 0.00398423f $X=2.56 $Y=1.68 $X2=0 $Y2=0
cc_136 N_A_95_306#_c_141_n N_B2_M1000_g 0.0145118f $X=3.63 $Y=1.132 $X2=0 $Y2=0
cc_137 N_A_95_306#_c_142_n N_B2_M1000_g 4.59187e-19 $X=3.96 $Y=1.132 $X2=0 $Y2=0
cc_138 N_A_95_306#_c_159_n N_B2_M1019_g 0.00472091f $X=4.25 $Y=2.78 $X2=0 $Y2=0
cc_139 N_A_95_306#_c_142_n N_B2_M1022_g 4.50172e-19 $X=3.96 $Y=1.132 $X2=0 $Y2=0
cc_140 N_A_95_306#_c_144_n N_B2_M1022_g 0.015625f $X=5.725 $Y=1.145 $X2=0 $Y2=0
cc_141 N_A_95_306#_c_157_n N_B2_c_328_n 0.00530716f $X=2.56 $Y=2.905 $X2=0 $Y2=0
cc_142 N_A_95_306#_M1014_s N_B2_c_329_n 0.00268337f $X=4.115 $Y=1.96 $X2=0 $Y2=0
cc_143 N_A_95_306#_c_144_n N_B2_c_321_n 0.0134773f $X=5.725 $Y=1.145 $X2=0 $Y2=0
cc_144 N_A_95_306#_c_144_n N_B2_c_322_n 0.0337589f $X=5.725 $Y=1.145 $X2=0 $Y2=0
cc_145 N_A_95_306#_c_144_n N_B2_c_323_n 0.00414034f $X=5.725 $Y=1.145 $X2=0
+ $Y2=0
cc_146 N_A_95_306#_c_140_n N_B2_c_324_n 0.00182761f $X=2.56 $Y=1.68 $X2=0 $Y2=0
cc_147 N_A_95_306#_c_157_n N_B2_c_324_n 0.00180383f $X=2.56 $Y=2.905 $X2=0 $Y2=0
cc_148 N_A_95_306#_c_141_n N_B2_c_324_n 0.00500757f $X=3.63 $Y=1.132 $X2=0 $Y2=0
cc_149 N_A_95_306#_c_146_n N_B2_c_324_n 0.0139355f $X=2.645 $Y=1.515 $X2=0 $Y2=0
cc_150 N_A_95_306#_c_140_n N_B2_c_325_n 0.0205422f $X=2.56 $Y=1.68 $X2=0 $Y2=0
cc_151 N_A_95_306#_c_157_n N_B2_c_325_n 0.00342481f $X=2.56 $Y=2.905 $X2=0 $Y2=0
cc_152 N_A_95_306#_c_141_n N_B2_c_325_n 0.0221918f $X=3.63 $Y=1.132 $X2=0 $Y2=0
cc_153 N_A_95_306#_c_146_n N_B2_c_325_n 2.0818e-19 $X=2.645 $Y=1.515 $X2=0 $Y2=0
cc_154 N_A_95_306#_M1008_d N_B2_c_358_n 5.66935e-19 $X=3.215 $Y=1.96 $X2=0 $Y2=0
cc_155 N_A_95_306#_M1008_d N_B2_c_334_n 0.00109482f $X=3.215 $Y=1.96 $X2=0 $Y2=0
cc_156 N_A_95_306#_c_141_n N_B2_c_334_n 0.0103076f $X=3.63 $Y=1.132 $X2=0 $Y2=0
cc_157 N_A_95_306#_c_159_n N_B1_M1012_g 0.0117137f $X=4.25 $Y=2.78 $X2=0 $Y2=0
cc_158 N_A_95_306#_c_161_n N_B1_M1012_g 0.00466343f $X=3.515 $Y=2.867 $X2=0
+ $Y2=0
cc_159 N_A_95_306#_c_141_n N_B1_M1001_g 0.0077677f $X=3.63 $Y=1.132 $X2=0 $Y2=0
cc_160 N_A_95_306#_c_142_n N_B1_M1001_g 0.00306707f $X=3.96 $Y=1.132 $X2=0 $Y2=0
cc_161 N_A_95_306#_c_142_n N_B1_M1018_g 0.00351834f $X=3.96 $Y=1.132 $X2=0 $Y2=0
cc_162 N_A_95_306#_c_144_n N_B1_M1018_g 0.00900647f $X=5.725 $Y=1.145 $X2=0
+ $Y2=0
cc_163 N_A_95_306#_c_159_n N_B1_M1014_g 0.013547f $X=4.25 $Y=2.78 $X2=0 $Y2=0
cc_164 N_A_95_306#_c_161_n N_B1_M1014_g 4.43424e-19 $X=3.515 $Y=2.867 $X2=0
+ $Y2=0
cc_165 N_A_95_306#_c_141_n B1 0.0246846f $X=3.63 $Y=1.132 $X2=0 $Y2=0
cc_166 N_A_95_306#_c_141_n N_B1_c_419_n 4.06731e-19 $X=3.63 $Y=1.132 $X2=0 $Y2=0
cc_167 N_A_95_306#_c_142_n N_B1_c_419_n 0.00116486f $X=3.96 $Y=1.132 $X2=0 $Y2=0
cc_168 N_A_95_306#_c_144_n N_B1_c_419_n 7.92241e-19 $X=5.725 $Y=1.145 $X2=0
+ $Y2=0
cc_169 N_A_95_306#_c_143_n N_A1_M1003_g 0.00290472f $X=5.89 $Y=1.105 $X2=0 $Y2=0
cc_170 N_A_95_306#_c_144_n N_A1_M1003_g 0.00778018f $X=5.725 $Y=1.145 $X2=0
+ $Y2=0
cc_171 N_A_95_306#_c_143_n N_A1_M1013_g 0.00358331f $X=5.89 $Y=1.105 $X2=0 $Y2=0
cc_172 N_A_95_306#_c_143_n A1 0.0248801f $X=5.89 $Y=1.105 $X2=0 $Y2=0
cc_173 N_A_95_306#_c_144_n A1 0.0225843f $X=5.725 $Y=1.145 $X2=0 $Y2=0
cc_174 N_A_95_306#_c_143_n N_A1_c_471_n 0.00245375f $X=5.89 $Y=1.105 $X2=0 $Y2=0
cc_175 N_A_95_306#_c_144_n N_A1_c_471_n 0.00182565f $X=5.725 $Y=1.145 $X2=0
+ $Y2=0
cc_176 N_A_95_306#_c_143_n N_A2_M1002_g 4.29877e-19 $X=5.89 $Y=1.105 $X2=0 $Y2=0
cc_177 N_A_95_306#_c_144_n N_A2_M1002_g 0.0172761f $X=5.725 $Y=1.145 $X2=0 $Y2=0
cc_178 N_A_95_306#_c_144_n N_A2_c_524_n 0.0131753f $X=5.725 $Y=1.145 $X2=0 $Y2=0
cc_179 N_A_95_306#_c_144_n A2 0.0099843f $X=5.725 $Y=1.145 $X2=0 $Y2=0
cc_180 N_A_95_306#_c_144_n N_A2_c_526_n 5.55026e-19 $X=5.725 $Y=1.145 $X2=0
+ $Y2=0
cc_181 N_A_95_306#_M1009_g N_VPWR_c_583_n 0.0197062f $X=0.565 $Y=2.4 $X2=0 $Y2=0
cc_182 N_A_95_306#_M1010_g N_VPWR_c_583_n 6.64525e-19 $X=1.015 $Y=2.4 $X2=0
+ $Y2=0
cc_183 N_A_95_306#_M1009_g N_VPWR_c_584_n 6.92757e-19 $X=0.565 $Y=2.4 $X2=0
+ $Y2=0
cc_184 N_A_95_306#_M1010_g N_VPWR_c_584_n 0.0186187f $X=1.015 $Y=2.4 $X2=0 $Y2=0
cc_185 N_A_95_306#_c_133_n N_VPWR_c_584_n 0.00188407f $X=1.28 $Y=1.605 $X2=0
+ $Y2=0
cc_186 N_A_95_306#_M1011_g N_VPWR_c_584_n 0.00334711f $X=1.465 $Y=2.4 $X2=0
+ $Y2=0
cc_187 N_A_95_306#_M1015_g N_VPWR_c_585_n 0.00542061f $X=1.915 $Y=2.4 $X2=0
+ $Y2=0
cc_188 N_A_95_306#_c_221_p N_VPWR_c_585_n 0.0202791f $X=2.475 $Y=1.515 $X2=0
+ $Y2=0
cc_189 N_A_95_306#_c_157_n N_VPWR_c_585_n 0.0817994f $X=2.56 $Y=2.905 $X2=0
+ $Y2=0
cc_190 N_A_95_306#_c_158_n N_VPWR_c_585_n 0.0147457f $X=2.645 $Y=2.99 $X2=0
+ $Y2=0
cc_191 N_A_95_306#_c_146_n N_VPWR_c_585_n 0.0067372f $X=2.645 $Y=1.515 $X2=0
+ $Y2=0
cc_192 N_A_95_306#_M1009_g N_VPWR_c_590_n 0.00460063f $X=0.565 $Y=2.4 $X2=0
+ $Y2=0
cc_193 N_A_95_306#_M1010_g N_VPWR_c_590_n 0.00460063f $X=1.015 $Y=2.4 $X2=0
+ $Y2=0
cc_194 N_A_95_306#_M1011_g N_VPWR_c_591_n 0.005209f $X=1.465 $Y=2.4 $X2=0 $Y2=0
cc_195 N_A_95_306#_M1015_g N_VPWR_c_591_n 0.005209f $X=1.915 $Y=2.4 $X2=0 $Y2=0
cc_196 N_A_95_306#_c_158_n N_VPWR_c_592_n 0.0121867f $X=2.645 $Y=2.99 $X2=0
+ $Y2=0
cc_197 N_A_95_306#_c_159_n N_VPWR_c_592_n 0.0369149f $X=4.25 $Y=2.78 $X2=0 $Y2=0
cc_198 N_A_95_306#_c_160_n N_VPWR_c_592_n 0.0567478f $X=3.185 $Y=2.867 $X2=0
+ $Y2=0
cc_199 N_A_95_306#_M1009_g N_VPWR_c_581_n 0.00908554f $X=0.565 $Y=2.4 $X2=0
+ $Y2=0
cc_200 N_A_95_306#_M1010_g N_VPWR_c_581_n 0.00908554f $X=1.015 $Y=2.4 $X2=0
+ $Y2=0
cc_201 N_A_95_306#_M1011_g N_VPWR_c_581_n 0.00982266f $X=1.465 $Y=2.4 $X2=0
+ $Y2=0
cc_202 N_A_95_306#_M1015_g N_VPWR_c_581_n 0.00987399f $X=1.915 $Y=2.4 $X2=0
+ $Y2=0
cc_203 N_A_95_306#_c_158_n N_VPWR_c_581_n 0.00660921f $X=2.645 $Y=2.99 $X2=0
+ $Y2=0
cc_204 N_A_95_306#_c_159_n N_VPWR_c_581_n 0.0306828f $X=4.25 $Y=2.78 $X2=0 $Y2=0
cc_205 N_A_95_306#_c_160_n N_VPWR_c_581_n 0.0320004f $X=3.185 $Y=2.867 $X2=0
+ $Y2=0
cc_206 N_A_95_306#_M1009_g N_X_c_676_n 0.00418763f $X=0.565 $Y=2.4 $X2=0 $Y2=0
cc_207 N_A_95_306#_c_131_n N_X_c_676_n 0.00457783f $X=0.925 $Y=1.605 $X2=0 $Y2=0
cc_208 N_A_95_306#_M1010_g N_X_c_676_n 0.00232604f $X=1.015 $Y=2.4 $X2=0 $Y2=0
cc_209 N_A_95_306#_M1005_g N_X_c_671_n 0.00813435f $X=1.355 $Y=0.87 $X2=0 $Y2=0
cc_210 N_A_95_306#_c_135_n N_X_c_671_n 3.97481e-19 $X=1.785 $Y=1.35 $X2=0 $Y2=0
cc_211 N_A_95_306#_c_139_n N_X_c_671_n 2.14997e-19 $X=1.417 $Y=1.605 $X2=0 $Y2=0
cc_212 N_A_95_306#_M1010_g N_X_c_677_n 8.23405e-19 $X=1.015 $Y=2.4 $X2=0 $Y2=0
cc_213 N_A_95_306#_M1011_g N_X_c_677_n 0.0195345f $X=1.465 $Y=2.4 $X2=0 $Y2=0
cc_214 N_A_95_306#_M1015_g N_X_c_677_n 0.0208717f $X=1.915 $Y=2.4 $X2=0 $Y2=0
cc_215 N_A_95_306#_c_139_n N_X_c_677_n 0.00101194f $X=1.417 $Y=1.605 $X2=0 $Y2=0
cc_216 N_A_95_306#_c_221_p N_X_c_677_n 0.00231492f $X=2.475 $Y=1.515 $X2=0 $Y2=0
cc_217 N_A_95_306#_c_157_n N_X_c_677_n 0.00474608f $X=2.56 $Y=2.905 $X2=0 $Y2=0
cc_218 N_A_95_306#_c_145_n N_X_c_677_n 0.00252337f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_219 N_A_95_306#_c_146_n N_X_c_677_n 0.00189656f $X=2.645 $Y=1.515 $X2=0 $Y2=0
cc_220 N_A_95_306#_c_135_n N_X_c_692_n 0.00202331f $X=1.785 $Y=1.35 $X2=0 $Y2=0
cc_221 N_A_95_306#_c_136_n N_X_c_692_n 0.01168f $X=2.215 $Y=1.35 $X2=0 $Y2=0
cc_222 N_A_95_306#_c_221_p N_X_c_692_n 0.0299782f $X=2.475 $Y=1.515 $X2=0 $Y2=0
cc_223 N_A_95_306#_c_140_n N_X_c_692_n 0.00341346f $X=2.56 $Y=1.68 $X2=0 $Y2=0
cc_224 N_A_95_306#_c_146_n N_X_c_692_n 0.00584539f $X=2.645 $Y=1.515 $X2=0 $Y2=0
cc_225 N_A_95_306#_c_135_n N_X_c_672_n 6.0186e-19 $X=1.785 $Y=1.35 $X2=0 $Y2=0
cc_226 N_A_95_306#_c_136_n N_X_c_672_n 0.00736569f $X=2.215 $Y=1.35 $X2=0 $Y2=0
cc_227 N_A_95_306#_c_131_n N_X_c_673_n 0.00397312f $X=0.925 $Y=1.605 $X2=0 $Y2=0
cc_228 N_A_95_306#_c_133_n N_X_c_673_n 0.00738952f $X=1.28 $Y=1.605 $X2=0 $Y2=0
cc_229 N_A_95_306#_M1005_g N_X_c_673_n 0.0199862f $X=1.355 $Y=0.87 $X2=0 $Y2=0
cc_230 N_A_95_306#_c_138_n N_X_c_673_n 0.0138583f $X=1.015 $Y=1.605 $X2=0 $Y2=0
cc_231 N_A_95_306#_c_139_n N_X_c_673_n 0.00599317f $X=1.417 $Y=1.605 $X2=0 $Y2=0
cc_232 N_A_95_306#_M1005_g N_X_c_704_n 0.0105486f $X=1.355 $Y=0.87 $X2=0 $Y2=0
cc_233 N_A_95_306#_c_135_n N_X_c_704_n 0.0148936f $X=1.785 $Y=1.35 $X2=0 $Y2=0
cc_234 N_A_95_306#_c_136_n N_X_c_704_n 0.00103837f $X=2.215 $Y=1.35 $X2=0 $Y2=0
cc_235 N_A_95_306#_c_139_n N_X_c_704_n 0.00880219f $X=1.417 $Y=1.605 $X2=0 $Y2=0
cc_236 N_A_95_306#_c_221_p N_X_c_704_n 0.025226f $X=2.475 $Y=1.515 $X2=0 $Y2=0
cc_237 N_A_95_306#_c_145_n N_X_c_704_n 0.00364852f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_238 N_A_95_306#_c_146_n N_X_c_704_n 0.0109931f $X=2.645 $Y=1.515 $X2=0 $Y2=0
cc_239 N_A_95_306#_c_131_n X 0.0110935f $X=0.925 $Y=1.605 $X2=0 $Y2=0
cc_240 N_A_95_306#_c_132_n N_X_c_675_n 0.0101126f $X=0.655 $Y=1.605 $X2=0 $Y2=0
cc_241 N_A_95_306#_c_160_n N_A_555_392#_M1008_s 0.00352558f $X=3.185 $Y=2.867
+ $X2=-0.19 $Y2=-0.245
cc_242 N_A_95_306#_c_159_n N_A_555_392#_M1012_d 0.00169505f $X=4.25 $Y=2.78
+ $X2=0 $Y2=0
cc_243 N_A_95_306#_c_140_n N_A_555_392#_c_735_n 0.0026803f $X=2.56 $Y=1.68 $X2=0
+ $Y2=0
cc_244 N_A_95_306#_c_157_n N_A_555_392#_c_735_n 0.0587925f $X=2.56 $Y=2.905
+ $X2=0 $Y2=0
cc_245 N_A_95_306#_c_141_n N_A_555_392#_c_735_n 0.00410878f $X=3.63 $Y=1.132
+ $X2=0 $Y2=0
cc_246 N_A_95_306#_M1008_d N_A_555_392#_c_749_n 0.00326883f $X=3.215 $Y=1.96
+ $X2=0 $Y2=0
cc_247 N_A_95_306#_M1014_s N_A_555_392#_c_749_n 0.00435499f $X=4.115 $Y=1.96
+ $X2=0 $Y2=0
cc_248 N_A_95_306#_c_160_n N_A_555_392#_c_749_n 0.00420217f $X=3.185 $Y=2.867
+ $X2=0 $Y2=0
cc_249 N_A_95_306#_c_161_n N_A_555_392#_c_749_n 0.0641284f $X=3.515 $Y=2.867
+ $X2=0 $Y2=0
cc_250 N_A_95_306#_c_144_n N_A_555_392#_c_736_n 0.00674632f $X=5.725 $Y=1.145
+ $X2=0 $Y2=0
cc_251 N_A_95_306#_c_160_n N_A_555_392#_c_754_n 0.0123303f $X=3.185 $Y=2.867
+ $X2=0 $Y2=0
cc_252 N_A_95_306#_c_159_n N_A_555_392#_c_742_n 0.0123955f $X=4.25 $Y=2.78 $X2=0
+ $Y2=0
cc_253 N_A_95_306#_c_140_n N_VGND_M1020_s 8.59214e-19 $X=2.56 $Y=1.68 $X2=0
+ $Y2=0
cc_254 N_A_95_306#_c_141_n N_VGND_M1020_s 0.00172209f $X=3.63 $Y=1.132 $X2=0
+ $Y2=0
cc_255 N_A_95_306#_c_144_n N_VGND_M1022_s 0.0128721f $X=5.725 $Y=1.145 $X2=0
+ $Y2=0
cc_256 N_A_95_306#_M1005_g N_VGND_c_809_n 0.00564714f $X=1.355 $Y=0.87 $X2=0
+ $Y2=0
cc_257 N_A_95_306#_c_138_n N_VGND_c_809_n 8.71085e-19 $X=1.015 $Y=1.605 $X2=0
+ $Y2=0
cc_258 N_A_95_306#_M1005_g N_VGND_c_810_n 4.52371e-19 $X=1.355 $Y=0.87 $X2=0
+ $Y2=0
cc_259 N_A_95_306#_c_135_n N_VGND_c_810_n 0.00782105f $X=1.785 $Y=1.35 $X2=0
+ $Y2=0
cc_260 N_A_95_306#_c_136_n N_VGND_c_810_n 0.00159705f $X=2.215 $Y=1.35 $X2=0
+ $Y2=0
cc_261 N_A_95_306#_c_136_n N_VGND_c_811_n 4.76302e-19 $X=2.215 $Y=1.35 $X2=0
+ $Y2=0
cc_262 N_A_95_306#_c_137_n N_VGND_c_811_n 0.0105834f $X=2.645 $Y=1.35 $X2=0
+ $Y2=0
cc_263 N_A_95_306#_c_140_n N_VGND_c_811_n 0.00892131f $X=2.56 $Y=1.68 $X2=0
+ $Y2=0
cc_264 N_A_95_306#_c_141_n N_VGND_c_811_n 0.013225f $X=3.63 $Y=1.132 $X2=0 $Y2=0
cc_265 N_A_95_306#_c_144_n N_VGND_c_812_n 0.015373f $X=5.725 $Y=1.145 $X2=0
+ $Y2=0
cc_266 N_A_95_306#_M1005_g N_VGND_c_816_n 0.00467453f $X=1.355 $Y=0.87 $X2=0
+ $Y2=0
cc_267 N_A_95_306#_c_135_n N_VGND_c_816_n 0.00405273f $X=1.785 $Y=1.35 $X2=0
+ $Y2=0
cc_268 N_A_95_306#_c_136_n N_VGND_c_818_n 0.00467453f $X=2.215 $Y=1.35 $X2=0
+ $Y2=0
cc_269 N_A_95_306#_c_137_n N_VGND_c_818_n 0.00405273f $X=2.645 $Y=1.35 $X2=0
+ $Y2=0
cc_270 N_A_95_306#_M1005_g N_VGND_c_824_n 0.00505379f $X=1.355 $Y=0.87 $X2=0
+ $Y2=0
cc_271 N_A_95_306#_c_135_n N_VGND_c_824_n 0.00424518f $X=1.785 $Y=1.35 $X2=0
+ $Y2=0
cc_272 N_A_95_306#_c_136_n N_VGND_c_824_n 0.00505379f $X=2.215 $Y=1.35 $X2=0
+ $Y2=0
cc_273 N_A_95_306#_c_137_n N_VGND_c_824_n 0.00424518f $X=2.645 $Y=1.35 $X2=0
+ $Y2=0
cc_274 N_A_95_306#_c_141_n N_A_645_120#_M1000_d 0.00216063f $X=3.63 $Y=1.132
+ $X2=-0.19 $Y2=-0.245
cc_275 N_A_95_306#_c_144_n N_A_645_120#_M1018_s 0.00224844f $X=5.725 $Y=1.145
+ $X2=0 $Y2=0
cc_276 N_A_95_306#_c_144_n N_A_645_120#_c_897_n 0.0161813f $X=5.725 $Y=1.145
+ $X2=0 $Y2=0
cc_277 N_A_95_306#_M1001_d N_A_645_120#_c_898_n 0.00169898f $X=3.655 $Y=0.6
+ $X2=0 $Y2=0
cc_278 N_A_95_306#_c_141_n N_A_645_120#_c_898_n 0.0162287f $X=3.63 $Y=1.132
+ $X2=0 $Y2=0
cc_279 N_A_95_306#_c_142_n N_A_645_120#_c_898_n 0.0163695f $X=3.96 $Y=1.132
+ $X2=0 $Y2=0
cc_280 N_A_95_306#_c_144_n N_A_645_120#_c_898_n 0.00607509f $X=5.725 $Y=1.145
+ $X2=0 $Y2=0
cc_281 N_A_95_306#_c_144_n N_A_1064_123#_M1002_d 0.00210096f $X=5.725 $Y=1.145
+ $X2=-0.19 $Y2=-0.245
cc_282 N_A_95_306#_M1003_d N_A_1064_123#_c_917_n 0.00408194f $X=5.75 $Y=0.615
+ $X2=0 $Y2=0
cc_283 N_A_95_306#_c_143_n N_A_1064_123#_c_917_n 0.0158841f $X=5.89 $Y=1.105
+ $X2=0 $Y2=0
cc_284 N_A_95_306#_c_144_n N_A_1064_123#_c_917_n 0.0164704f $X=5.725 $Y=1.145
+ $X2=0 $Y2=0
cc_285 N_A_95_306#_c_143_n N_A_1064_123#_c_915_n 0.0106625f $X=5.89 $Y=1.105
+ $X2=0 $Y2=0
cc_286 N_B2_M1008_g N_B1_M1012_g 0.0448754f $X=3.125 $Y=2.46 $X2=0 $Y2=0
cc_287 N_B2_c_328_n N_B1_M1012_g 0.00354307f $X=3.24 $Y=1.935 $X2=0 $Y2=0
cc_288 N_B2_c_329_n N_B1_M1012_g 8.82362e-19 $X=4.11 $Y=1.935 $X2=0 $Y2=0
cc_289 N_B2_c_334_n N_B1_M1012_g 0.0135008f $X=4.025 $Y=2.042 $X2=0 $Y2=0
cc_290 N_B2_M1000_g N_B1_M1001_g 0.0291033f $X=3.15 $Y=0.92 $X2=0 $Y2=0
cc_291 N_B2_M1022_g N_B1_M1018_g 0.0246028f $X=4.485 $Y=0.935 $X2=0 $Y2=0
cc_292 N_B2_M1019_g N_B1_M1014_g 0.0445324f $X=4.475 $Y=2.46 $X2=0 $Y2=0
cc_293 N_B2_c_329_n N_B1_M1014_g 0.00879217f $X=4.11 $Y=1.935 $X2=0 $Y2=0
cc_294 N_B2_c_334_n N_B1_M1014_g 0.00807945f $X=4.025 $Y=2.042 $X2=0 $Y2=0
cc_295 N_B2_c_321_n B1 0.0226234f $X=4.195 $Y=1.605 $X2=0 $Y2=0
cc_296 N_B2_c_324_n B1 3.6348e-19 $X=3.11 $Y=1.6 $X2=0 $Y2=0
cc_297 N_B2_c_325_n B1 0.0258902f $X=3.24 $Y=1.6 $X2=0 $Y2=0
cc_298 N_B2_c_334_n B1 0.0245722f $X=4.025 $Y=2.042 $X2=0 $Y2=0
cc_299 N_B2_M1022_g N_B1_c_419_n 2.32253e-19 $X=4.485 $Y=0.935 $X2=0 $Y2=0
cc_300 N_B2_c_321_n N_B1_c_419_n 0.0118645f $X=4.195 $Y=1.605 $X2=0 $Y2=0
cc_301 N_B2_c_323_n N_B1_c_419_n 0.021459f $X=4.49 $Y=1.605 $X2=0 $Y2=0
cc_302 N_B2_c_324_n N_B1_c_419_n 0.0216346f $X=3.11 $Y=1.6 $X2=0 $Y2=0
cc_303 N_B2_c_325_n N_B1_c_419_n 0.00203145f $X=3.24 $Y=1.6 $X2=0 $Y2=0
cc_304 N_B2_c_334_n N_B1_c_419_n 0.00107735f $X=4.025 $Y=2.042 $X2=0 $Y2=0
cc_305 N_B2_M1019_g N_A2_M1006_g 0.0139875f $X=4.475 $Y=2.46 $X2=0 $Y2=0
cc_306 N_B2_M1022_g N_A2_M1002_g 0.0108695f $X=4.485 $Y=0.935 $X2=0 $Y2=0
cc_307 N_B2_M1022_g N_A2_c_524_n 0.00562171f $X=4.485 $Y=0.935 $X2=0 $Y2=0
cc_308 N_B2_c_322_n N_A2_c_524_n 0.00222306f $X=4.49 $Y=1.605 $X2=0 $Y2=0
cc_309 N_B2_c_323_n N_A2_c_524_n 0.0200398f $X=4.49 $Y=1.605 $X2=0 $Y2=0
cc_310 N_B2_M1022_g A2 3.85498e-19 $X=4.485 $Y=0.935 $X2=0 $Y2=0
cc_311 N_B2_M1022_g N_A2_c_526_n 4.96786e-19 $X=4.485 $Y=0.935 $X2=0 $Y2=0
cc_312 N_B2_M1019_g N_VPWR_c_586_n 6.2684e-19 $X=4.475 $Y=2.46 $X2=0 $Y2=0
cc_313 N_B2_M1008_g N_VPWR_c_592_n 0.00333926f $X=3.125 $Y=2.46 $X2=0 $Y2=0
cc_314 N_B2_M1019_g N_VPWR_c_592_n 0.00519794f $X=4.475 $Y=2.46 $X2=0 $Y2=0
cc_315 N_B2_M1008_g N_VPWR_c_581_n 0.00427931f $X=3.125 $Y=2.46 $X2=0 $Y2=0
cc_316 N_B2_M1019_g N_VPWR_c_581_n 0.00535486f $X=4.475 $Y=2.46 $X2=0 $Y2=0
cc_317 N_B2_c_334_n N_A_555_392#_M1012_d 0.00167444f $X=4.025 $Y=2.042 $X2=0
+ $Y2=0
cc_318 N_B2_M1008_g N_A_555_392#_c_735_n 8.76298e-19 $X=3.125 $Y=2.46 $X2=0
+ $Y2=0
cc_319 N_B2_c_324_n N_A_555_392#_c_735_n 0.00117128f $X=3.11 $Y=1.6 $X2=0 $Y2=0
cc_320 N_B2_c_358_n N_A_555_392#_c_735_n 0.00956392f $X=3.325 $Y=2.042 $X2=0
+ $Y2=0
cc_321 N_B2_M1008_g N_A_555_392#_c_749_n 0.0132079f $X=3.125 $Y=2.46 $X2=0 $Y2=0
cc_322 N_B2_M1019_g N_A_555_392#_c_749_n 0.0132548f $X=4.475 $Y=2.46 $X2=0 $Y2=0
cc_323 N_B2_c_329_n N_A_555_392#_c_749_n 0.00875864f $X=4.11 $Y=1.935 $X2=0
+ $Y2=0
cc_324 N_B2_c_322_n N_A_555_392#_c_749_n 0.01086f $X=4.49 $Y=1.605 $X2=0 $Y2=0
cc_325 N_B2_c_323_n N_A_555_392#_c_749_n 8.25875e-19 $X=4.49 $Y=1.605 $X2=0
+ $Y2=0
cc_326 N_B2_c_325_n N_A_555_392#_c_749_n 0.00341618f $X=3.24 $Y=1.6 $X2=0 $Y2=0
cc_327 N_B2_c_358_n N_A_555_392#_c_749_n 0.00844548f $X=3.325 $Y=2.042 $X2=0
+ $Y2=0
cc_328 N_B2_c_334_n N_A_555_392#_c_749_n 0.0376457f $X=4.025 $Y=2.042 $X2=0
+ $Y2=0
cc_329 N_B2_M1019_g N_A_555_392#_c_736_n 2.39624e-19 $X=4.475 $Y=2.46 $X2=0
+ $Y2=0
cc_330 N_B2_c_329_n N_A_555_392#_c_736_n 0.00461309f $X=4.11 $Y=1.935 $X2=0
+ $Y2=0
cc_331 N_B2_c_322_n N_A_555_392#_c_736_n 0.00337333f $X=4.49 $Y=1.605 $X2=0
+ $Y2=0
cc_332 N_B2_c_323_n N_A_555_392#_c_736_n 9.31826e-19 $X=4.49 $Y=1.605 $X2=0
+ $Y2=0
cc_333 N_B2_M1000_g N_VGND_c_811_n 0.00499212f $X=3.15 $Y=0.92 $X2=0 $Y2=0
cc_334 N_B2_M1022_g N_VGND_c_812_n 0.008067f $X=4.485 $Y=0.935 $X2=0 $Y2=0
cc_335 N_B2_M1000_g N_VGND_c_823_n 0.00411835f $X=3.15 $Y=0.92 $X2=0 $Y2=0
cc_336 N_B2_M1022_g N_VGND_c_823_n 0.00349617f $X=4.485 $Y=0.935 $X2=0 $Y2=0
cc_337 N_B2_M1000_g N_VGND_c_824_n 0.00476395f $X=3.15 $Y=0.92 $X2=0 $Y2=0
cc_338 N_B2_M1022_g N_VGND_c_824_n 0.00396651f $X=4.485 $Y=0.935 $X2=0 $Y2=0
cc_339 N_B2_M1022_g N_A_645_120#_c_897_n 2.97537e-19 $X=4.485 $Y=0.935 $X2=0
+ $Y2=0
cc_340 N_B2_M1000_g N_A_645_120#_c_898_n 0.00359638f $X=3.15 $Y=0.92 $X2=0 $Y2=0
cc_341 N_B1_M1012_g N_VPWR_c_592_n 0.00347303f $X=3.575 $Y=2.46 $X2=0 $Y2=0
cc_342 N_B1_M1014_g N_VPWR_c_592_n 0.00349978f $X=4.025 $Y=2.46 $X2=0 $Y2=0
cc_343 N_B1_M1012_g N_VPWR_c_581_n 0.00428491f $X=3.575 $Y=2.46 $X2=0 $Y2=0
cc_344 N_B1_M1014_g N_VPWR_c_581_n 0.00429629f $X=4.025 $Y=2.46 $X2=0 $Y2=0
cc_345 N_B1_M1012_g N_A_555_392#_c_749_n 0.0096306f $X=3.575 $Y=2.46 $X2=0 $Y2=0
cc_346 N_B1_M1014_g N_A_555_392#_c_749_n 0.0096269f $X=4.025 $Y=2.46 $X2=0 $Y2=0
cc_347 N_B1_M1018_g N_VGND_c_812_n 9.3562e-19 $X=4.01 $Y=0.92 $X2=0 $Y2=0
cc_348 N_B1_M1001_g N_VGND_c_823_n 0.00327294f $X=3.58 $Y=0.92 $X2=0 $Y2=0
cc_349 N_B1_M1018_g N_VGND_c_823_n 0.00327294f $X=4.01 $Y=0.92 $X2=0 $Y2=0
cc_350 N_B1_M1001_g N_VGND_c_824_n 0.00476395f $X=3.58 $Y=0.92 $X2=0 $Y2=0
cc_351 N_B1_M1018_g N_VGND_c_824_n 0.00476395f $X=4.01 $Y=0.92 $X2=0 $Y2=0
cc_352 N_B1_M1001_g N_A_645_120#_c_898_n 0.0114295f $X=3.58 $Y=0.92 $X2=0 $Y2=0
cc_353 N_B1_M1018_g N_A_645_120#_c_898_n 0.0114847f $X=4.01 $Y=0.92 $X2=0 $Y2=0
cc_354 A1 N_A2_M1006_g 0.00707418f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_355 N_A1_c_471_n N_A2_M1006_g 0.0327512f $X=6.105 $Y=1.615 $X2=0 $Y2=0
cc_356 N_A1_M1003_g N_A2_c_520_n 0.00985192f $X=5.675 $Y=0.935 $X2=0 $Y2=0
cc_357 N_A1_M1013_g N_A2_c_520_n 0.00985192f $X=6.105 $Y=0.935 $X2=0 $Y2=0
cc_358 N_A1_M1013_g N_A2_c_521_n 0.0130116f $X=6.105 $Y=0.935 $X2=0 $Y2=0
cc_359 N_A1_M1021_g N_A2_M1016_g 0.0283677f $X=6.07 $Y=2.46 $X2=0 $Y2=0
cc_360 A1 N_A2_M1016_g 0.00184168f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_361 N_A1_c_471_n N_A2_M1016_g 0.0130116f $X=6.105 $Y=1.615 $X2=0 $Y2=0
cc_362 N_A1_M1013_g N_A2_M1023_g 0.00918444f $X=6.105 $Y=0.935 $X2=0 $Y2=0
cc_363 A1 N_A2_c_524_n 8.81484e-19 $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_364 N_A1_c_471_n N_A2_c_524_n 0.00192331f $X=6.105 $Y=1.615 $X2=0 $Y2=0
cc_365 N_A1_M1003_g N_A2_c_526_n 0.0301212f $X=5.675 $Y=0.935 $X2=0 $Y2=0
cc_366 N_A1_M1004_g N_VPWR_c_586_n 0.00728073f $X=5.62 $Y=2.46 $X2=0 $Y2=0
cc_367 N_A1_M1004_g N_VPWR_c_587_n 5.56271e-19 $X=5.62 $Y=2.46 $X2=0 $Y2=0
cc_368 N_A1_M1021_g N_VPWR_c_587_n 0.0134077f $X=6.07 $Y=2.46 $X2=0 $Y2=0
cc_369 N_A1_M1004_g N_VPWR_c_588_n 0.005209f $X=5.62 $Y=2.46 $X2=0 $Y2=0
cc_370 N_A1_M1021_g N_VPWR_c_588_n 0.00460063f $X=6.07 $Y=2.46 $X2=0 $Y2=0
cc_371 N_A1_M1004_g N_VPWR_c_581_n 0.00983402f $X=5.62 $Y=2.46 $X2=0 $Y2=0
cc_372 N_A1_M1021_g N_VPWR_c_581_n 0.00908554f $X=6.07 $Y=2.46 $X2=0 $Y2=0
cc_373 N_A1_M1004_g N_A_555_392#_c_737_n 0.0138961f $X=5.62 $Y=2.46 $X2=0 $Y2=0
cc_374 A1 N_A_555_392#_c_737_n 0.0205887f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_375 N_A1_M1004_g N_A_555_392#_c_738_n 0.0120462f $X=5.62 $Y=2.46 $X2=0 $Y2=0
cc_376 N_A1_M1021_g N_A_555_392#_c_739_n 0.015699f $X=6.07 $Y=2.46 $X2=0 $Y2=0
cc_377 A1 N_A_555_392#_c_739_n 0.0133617f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_378 N_A1_c_471_n N_A_555_392#_c_739_n 8.30124e-19 $X=6.105 $Y=1.615 $X2=0
+ $Y2=0
cc_379 N_A1_M1004_g N_A_555_392#_c_743_n 0.0010042f $X=5.62 $Y=2.46 $X2=0 $Y2=0
cc_380 A1 N_A_555_392#_c_743_n 0.0209507f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_381 N_A1_c_471_n N_A_555_392#_c_743_n 0.00225438f $X=6.105 $Y=1.615 $X2=0
+ $Y2=0
cc_382 N_A1_M1013_g N_VGND_c_813_n 5.60436e-19 $X=6.105 $Y=0.935 $X2=0 $Y2=0
cc_383 N_A1_M1003_g N_VGND_c_824_n 9.15321e-19 $X=5.675 $Y=0.935 $X2=0 $Y2=0
cc_384 N_A1_M1013_g N_VGND_c_824_n 9.15321e-19 $X=6.105 $Y=0.935 $X2=0 $Y2=0
cc_385 N_A1_M1003_g N_A_1064_123#_c_917_n 0.00924024f $X=5.675 $Y=0.935 $X2=0
+ $Y2=0
cc_386 N_A1_M1013_g N_A_1064_123#_c_917_n 0.0116768f $X=6.105 $Y=0.935 $X2=0
+ $Y2=0
cc_387 A1 N_A_1064_123#_c_917_n 0.00149839f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_388 N_A1_M1013_g N_A_1064_123#_c_914_n 4.59247e-19 $X=6.105 $Y=0.935 $X2=0
+ $Y2=0
cc_389 N_A2_M1006_g N_VPWR_c_586_n 0.0231023f $X=4.955 $Y=2.46 $X2=0 $Y2=0
cc_390 N_A2_M1016_g N_VPWR_c_587_n 0.0164336f $X=6.52 $Y=2.46 $X2=0 $Y2=0
cc_391 N_A2_M1006_g N_VPWR_c_592_n 0.00521592f $X=4.955 $Y=2.46 $X2=0 $Y2=0
cc_392 N_A2_M1016_g N_VPWR_c_593_n 0.00460063f $X=6.52 $Y=2.46 $X2=0 $Y2=0
cc_393 N_A2_M1006_g N_VPWR_c_581_n 0.0102937f $X=4.955 $Y=2.46 $X2=0 $Y2=0
cc_394 N_A2_M1016_g N_VPWR_c_581_n 0.00912769f $X=6.52 $Y=2.46 $X2=0 $Y2=0
cc_395 N_A2_M1006_g N_A_555_392#_c_736_n 3.87094e-19 $X=4.955 $Y=2.46 $X2=0
+ $Y2=0
cc_396 N_A2_M1006_g N_A_555_392#_c_737_n 0.0210065f $X=4.955 $Y=2.46 $X2=0 $Y2=0
cc_397 N_A2_c_524_n N_A_555_392#_c_737_n 0.00766307f $X=5.245 $Y=1.405 $X2=0
+ $Y2=0
cc_398 N_A2_M1006_g N_A_555_392#_c_738_n 0.00114485f $X=4.955 $Y=2.46 $X2=0
+ $Y2=0
cc_399 N_A2_M1016_g N_A_555_392#_c_739_n 0.019475f $X=6.52 $Y=2.46 $X2=0 $Y2=0
cc_400 N_A2_M1016_g N_A_555_392#_c_740_n 4.17659e-19 $X=6.52 $Y=2.46 $X2=0 $Y2=0
cc_401 N_A2_M1016_g N_A_555_392#_c_741_n 4.69176e-19 $X=6.52 $Y=2.46 $X2=0 $Y2=0
cc_402 A2 N_VGND_M1022_s 0.00292336f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_403 N_A2_M1002_g N_VGND_c_812_n 0.00341364f $X=5.245 $Y=0.935 $X2=0 $Y2=0
cc_404 A2 N_VGND_c_812_n 0.0333508f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_405 N_A2_c_526_n N_VGND_c_812_n 0.00545095f $X=5.155 $Y=0.2 $X2=0 $Y2=0
cc_406 N_A2_c_520_n N_VGND_c_813_n 0.00811888f $X=6.46 $Y=0.2 $X2=0 $Y2=0
cc_407 N_A2_M1023_g N_VGND_c_813_n 0.026056f $X=6.535 $Y=0.935 $X2=0 $Y2=0
cc_408 A2 N_VGND_c_821_n 0.0236953f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_409 N_A2_c_526_n N_VGND_c_821_n 0.0403962f $X=5.155 $Y=0.2 $X2=0 $Y2=0
cc_410 N_A2_c_520_n N_VGND_c_824_n 0.0406735f $X=6.46 $Y=0.2 $X2=0 $Y2=0
cc_411 A2 N_VGND_c_824_n 0.0124201f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_412 N_A2_c_526_n N_VGND_c_824_n 0.0100036f $X=5.155 $Y=0.2 $X2=0 $Y2=0
cc_413 N_A2_M1002_g N_A_1064_123#_c_917_n 0.00393563f $X=5.245 $Y=0.935 $X2=0
+ $Y2=0
cc_414 N_A2_c_520_n N_A_1064_123#_c_917_n 0.00827463f $X=6.46 $Y=0.2 $X2=0 $Y2=0
cc_415 A2 N_A_1064_123#_c_917_n 0.00164856f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_416 N_A2_c_520_n N_A_1064_123#_c_914_n 0.00275881f $X=6.46 $Y=0.2 $X2=0 $Y2=0
cc_417 N_VPWR_c_583_n N_X_c_676_n 0.0362185f $X=0.34 $Y=1.985 $X2=0 $Y2=0
cc_418 N_VPWR_c_584_n N_X_c_676_n 0.0378999f $X=1.24 $Y=1.985 $X2=0 $Y2=0
cc_419 N_VPWR_c_590_n N_X_c_676_n 0.00749631f $X=1.075 $Y=3.33 $X2=0 $Y2=0
cc_420 N_VPWR_c_581_n N_X_c_676_n 0.0062048f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_421 N_VPWR_c_584_n N_X_c_677_n 0.0395686f $X=1.24 $Y=1.985 $X2=0 $Y2=0
cc_422 N_VPWR_c_585_n N_X_c_677_n 0.0379043f $X=2.14 $Y=2.015 $X2=0 $Y2=0
cc_423 N_VPWR_c_591_n N_X_c_677_n 0.0144623f $X=2.055 $Y=3.33 $X2=0 $Y2=0
cc_424 N_VPWR_c_581_n N_X_c_677_n 0.0118344f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_425 N_VPWR_c_584_n N_X_c_673_n 0.0213492f $X=1.24 $Y=1.985 $X2=0 $Y2=0
cc_426 N_VPWR_c_583_n N_X_c_675_n 0.0118946f $X=0.34 $Y=1.985 $X2=0 $Y2=0
cc_427 N_VPWR_c_581_n N_A_555_392#_c_749_n 0.00792216f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_428 N_VPWR_c_586_n N_A_555_392#_c_791_n 0.00234701f $X=5.27 $Y=2.375 $X2=0
+ $Y2=0
cc_429 N_VPWR_M1006_s N_A_555_392#_c_737_n 0.00504389f $X=5.045 $Y=1.96 $X2=0
+ $Y2=0
cc_430 N_VPWR_c_586_n N_A_555_392#_c_737_n 0.0308696f $X=5.27 $Y=2.375 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_586_n N_A_555_392#_c_738_n 0.0256472f $X=5.27 $Y=2.375 $X2=0
+ $Y2=0
cc_432 N_VPWR_c_587_n N_A_555_392#_c_738_n 0.0234083f $X=6.295 $Y=2.375 $X2=0
+ $Y2=0
cc_433 N_VPWR_c_588_n N_A_555_392#_c_738_n 0.0109793f $X=6.13 $Y=3.33 $X2=0
+ $Y2=0
cc_434 N_VPWR_c_581_n N_A_555_392#_c_738_n 0.00901959f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_435 N_VPWR_M1021_d N_A_555_392#_c_739_n 0.00165831f $X=6.16 $Y=1.96 $X2=0
+ $Y2=0
cc_436 N_VPWR_c_587_n N_A_555_392#_c_739_n 0.0170259f $X=6.295 $Y=2.375 $X2=0
+ $Y2=0
cc_437 N_VPWR_c_587_n N_A_555_392#_c_741_n 0.0234083f $X=6.295 $Y=2.375 $X2=0
+ $Y2=0
cc_438 N_VPWR_c_593_n N_A_555_392#_c_741_n 0.011066f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_439 N_VPWR_c_581_n N_A_555_392#_c_741_n 0.00915947f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_440 N_VPWR_c_586_n N_A_555_392#_c_742_n 0.0536134f $X=5.27 $Y=2.375 $X2=0
+ $Y2=0
cc_441 N_VPWR_c_592_n N_A_555_392#_c_742_n 0.011066f $X=5.035 $Y=3.33 $X2=0
+ $Y2=0
cc_442 N_VPWR_c_581_n N_A_555_392#_c_742_n 0.00915947f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_443 N_X_c_673_n N_VGND_M1005_s 0.00275278f $X=1.405 $Y=1.33 $X2=-0.19
+ $Y2=-0.245
cc_444 N_X_c_692_n N_VGND_M1007_s 0.0044545f $X=2.265 $Y=1.095 $X2=0 $Y2=0
cc_445 N_X_c_671_n N_VGND_c_809_n 0.0175587f $X=1.57 $Y=0.645 $X2=0 $Y2=0
cc_446 N_X_c_673_n N_VGND_c_809_n 0.0218366f $X=1.405 $Y=1.33 $X2=0 $Y2=0
cc_447 N_X_c_671_n N_VGND_c_810_n 0.0130934f $X=1.57 $Y=0.645 $X2=0 $Y2=0
cc_448 N_X_c_672_n N_VGND_c_810_n 0.0130934f $X=2.43 $Y=0.645 $X2=0 $Y2=0
cc_449 N_X_c_704_n N_VGND_c_810_n 0.0154032f $X=1.855 $Y=1.33 $X2=0 $Y2=0
cc_450 N_X_c_672_n N_VGND_c_811_n 0.0166774f $X=2.43 $Y=0.645 $X2=0 $Y2=0
cc_451 N_X_c_671_n N_VGND_c_816_n 0.00704565f $X=1.57 $Y=0.645 $X2=0 $Y2=0
cc_452 N_X_c_672_n N_VGND_c_818_n 0.00718756f $X=2.43 $Y=0.645 $X2=0 $Y2=0
cc_453 N_X_c_671_n N_VGND_c_824_n 0.00830435f $X=1.57 $Y=0.645 $X2=0 $Y2=0
cc_454 N_X_c_672_n N_VGND_c_824_n 0.0083989f $X=2.43 $Y=0.645 $X2=0 $Y2=0
cc_455 N_A_555_392#_c_739_n N_VGND_c_813_n 0.0021668f $X=6.66 $Y=2.035 $X2=0
+ $Y2=0
cc_456 N_A_555_392#_c_740_n N_VGND_c_813_n 0.00898193f $X=6.785 $Y=2.12 $X2=0
+ $Y2=0
cc_457 N_A_555_392#_c_739_n N_A_1064_123#_c_915_n 0.00539705f $X=6.66 $Y=2.035
+ $X2=0 $Y2=0
cc_458 N_VGND_c_812_n N_A_645_120#_c_897_n 0.0133114f $X=4.7 $Y=0.76 $X2=0 $Y2=0
cc_459 N_VGND_c_811_n N_A_645_120#_c_898_n 0.0109419f $X=2.86 $Y=0.75 $X2=0
+ $Y2=0
cc_460 N_VGND_c_823_n N_A_645_120#_c_898_n 0.0238447f $X=4.535 $Y=0 $X2=0 $Y2=0
cc_461 N_VGND_c_824_n N_A_645_120#_c_898_n 0.0346781f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_462 N_VGND_c_812_n N_A_1064_123#_c_917_n 0.00574236f $X=4.7 $Y=0.76 $X2=0
+ $Y2=0
cc_463 N_VGND_c_821_n N_A_1064_123#_c_917_n 0.0122684f $X=6.585 $Y=0 $X2=0 $Y2=0
cc_464 N_VGND_c_824_n N_A_1064_123#_c_917_n 0.0214259f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_465 N_VGND_c_813_n N_A_1064_123#_c_914_n 0.0096909f $X=6.75 $Y=0.76 $X2=0
+ $Y2=0
cc_466 N_VGND_c_821_n N_A_1064_123#_c_914_n 0.00374365f $X=6.585 $Y=0 $X2=0
+ $Y2=0
cc_467 N_VGND_c_824_n N_A_1064_123#_c_914_n 0.00464028f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_468 N_VGND_c_813_n N_A_1064_123#_c_915_n 0.0160983f $X=6.75 $Y=0.76 $X2=0
+ $Y2=0

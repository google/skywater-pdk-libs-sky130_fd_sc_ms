* File: sky130_fd_sc_ms__o21ai_2.spice
* Created: Fri Aug 28 17:54:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o21ai_2.pex.spice"
.subckt sky130_fd_sc_ms__o21ai_2  VNB VPB A1 A2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1009 N_A_27_74#_M1009_d N_A1_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.2
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1007 N_A_27_74#_M1007_d N_A2_M1007_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10915 AS=0.1295 PD=1.035 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1011 N_A_27_74#_M1007_d N_A2_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10915 AS=0.12395 PD=1.035 PS=1.075 NRD=2.424 NRS=8.916 M=1 R=4.93333
+ SA=75001.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1010 N_A_27_74#_M1010_d N_A1_M1010_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.12025 AS=0.12395 PD=1.065 PS=1.075 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1005 N_Y_M1005_d N_B1_M1005_g N_A_27_74#_M1010_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.11655 AS=0.12025 PD=1.055 PS=1.065 NRD=4.86 NRS=7.296 M=1 R=4.93333
+ SA=75002.1 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1008 N_Y_M1005_d N_B1_M1008_g N_A_27_74#_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.11655 AS=0.2109 PD=1.055 PS=2.05 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75002.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g N_A_119_368#_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90002.5 A=0.2016 P=2.6 MULT=1
MM1001 N_A_119_368#_M1000_s N_A2_M1001_g N_Y_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.6
+ SB=90002.1 A=0.2016 P=2.6 MULT=1
MM1003 N_A_119_368#_M1003_d N_A2_M1003_g N_Y_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_119_368#_M1003_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.6
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1004_d N_B1_M1004_g N_VPWR_M1002_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.1
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1006 N_Y_M1004_d N_B1_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__o21ai_2.pxi.spice"
*
.ends
*
*

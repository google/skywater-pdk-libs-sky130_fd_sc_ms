* NGSPICE file created from sky130_fd_sc_ms__einvp_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__einvp_1 A TE VGND VNB VPB VPWR Z
M1000 a_313_392# a_44_549# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=3.115e+11p ps=2.71e+06u
M1001 a_318_74# TE VGND VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=2.276e+11p ps=2.16e+06u
M1002 Z A a_318_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1003 VGND TE a_44_549# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.604e+11p ps=2.08e+06u
M1004 Z A a_313_392# VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1005 VPWR TE a_44_549# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=2.583e+11p ps=2.07e+06u
.ends


* File: sky130_fd_sc_ms__a32oi_2.spice
* Created: Fri Aug 28 17:08:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a32oi_2.pex.spice"
.subckt sky130_fd_sc_ms__a32oi_2  VNB VPB B2 B1 A1 A2 A3 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1011 N_A_27_74#_M1011_d N_B2_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1221 PD=2.05 PS=1.07 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1017 N_A_27_74#_M1017_d N_B2_M1017_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1221 PD=1.02 PS=1.07 NRD=0 NRS=8.1 M=1 R=4.93333 SA=75000.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1007 N_Y_M1007_d N_B1_M1007_g N_A_27_74#_M1017_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1010 N_Y_M1007_d N_B1_M1010_g N_A_27_74#_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.6
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1008 N_Y_M1008_d N_A1_M1008_g N_A_507_74#_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1018 N_Y_M1008_d N_A1_M1018_g N_A_507_74#_M1018_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.11285 PD=1.02 PS=1.045 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1012 N_A_507_74#_M1018_s N_A2_M1012_g N_A_771_74#_M1012_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.11285 AS=0.14615 PD=1.045 PS=1.135 NRD=4.044 NRS=7.296 M=1
+ R=4.93333 SA=75001.1 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1014 N_A_507_74#_M1014_d N_A2_M1014_g N_A_771_74#_M1012_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.14615 PD=2.05 PS=1.135 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_A_771_74#_M1005_d N_A3_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1009 N_A_771_74#_M1005_d N_A3_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_B2_M1000_g N_A_27_368#_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1764 AS=0.3192 PD=1.435 PS=2.81 NRD=7.0329 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90005.2 A=0.2016 P=2.6 MULT=1
MM1006 N_Y_M1000_d N_B2_M1006_g N_A_27_368#_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1764 AS=0.1792 PD=1.435 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.7
+ SB=90004.7 A=0.2016 P=2.6 MULT=1
MM1001 N_A_27_368#_M1006_s N_B1_M1001_g N_Y_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.2
+ SB=90004.2 A=0.2016 P=2.6 MULT=1
MM1003 N_A_27_368#_M1003_d N_B1_M1003_g N_Y_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90001.7
+ SB=90003.7 A=0.2016 P=2.6 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_27_368#_M1003_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3696 AS=0.1792 PD=1.78 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.2
+ SB=90003.2 A=0.2016 P=2.6 MULT=1
MM1015 N_VPWR_M1002_d N_A1_M1015_g N_A_27_368#_M1015_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3696 AS=0.1512 PD=1.78 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003
+ SB=90002.3 A=0.2016 P=2.6 MULT=1
MM1004 N_A_27_368#_M1015_s N_A2_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1876 PD=1.39 PS=1.455 NRD=0 NRS=8.7862 M=1 R=6.22222 SA=90003.5
+ SB=90001.9 A=0.2016 P=2.6 MULT=1
MM1019 N_A_27_368#_M1019_d N_A2_M1019_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2492 AS=0.1876 PD=1.565 PS=1.455 NRD=15.2281 NRS=0.8668 M=1 R=6.22222
+ SA=90004 SB=90001.4 A=0.2016 P=2.6 MULT=1
MM1013 N_VPWR_M1013_d N_A3_M1013_g N_A_27_368#_M1019_d VPB PSHORT L=0.18 W=1.12
+ AD=0.2072 AS=0.2492 PD=1.49 PS=1.565 NRD=7.8997 NRS=13.7703 M=1 R=6.22222
+ SA=90004.6 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1016 N_VPWR_M1013_d N_A3_M1016_g N_A_27_368#_M1016_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2072 AS=0.3136 PD=1.49 PS=2.8 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90005.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX20_noxref VNB VPB NWDIODE A=12.3132 P=16.96
*
.include "sky130_fd_sc_ms__a32oi_2.pxi.spice"
*
.ends
*
*

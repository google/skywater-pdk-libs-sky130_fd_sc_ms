* File: sky130_fd_sc_ms__and4_1.pex.spice
* Created: Wed Sep  2 11:58:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__AND4_1%A 3 7 9 10 12 13 14 18 19
c37 3 0 8.64864e-20 $X=0.555 $Y=2.54
r38 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.285 $X2=0.59 $Y2=1.285
r39 13 14 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.62 $Y=1.295
+ $X2=0.62 $Y2=1.665
r40 13 19 0.295498 $w=3.88e-07 $l=1e-08 $layer=LI1_cond $X=0.62 $Y=1.295
+ $X2=0.62 $Y2=1.285
r41 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.59 $Y=1.625
+ $X2=0.59 $Y2=1.285
r42 11 12 36.5727 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.625
+ $X2=0.59 $Y2=1.79
r43 10 18 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=0.59 $Y=1.235 $X2=0.59
+ $Y2=1.285
r44 9 10 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.66 $Y=1.085
+ $X2=0.66 $Y2=1.235
r45 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.82 $Y=0.69 $X2=0.82
+ $Y2=1.085
r46 3 12 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=0.555 $Y=2.54
+ $X2=0.555 $Y2=1.79
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_1%B 3 7 9 10 11 12 18
c38 9 0 1.73901e-19 $X=1.2 $Y=0.555
r39 18 21 40.7727 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.64
+ $X2=1.14 $Y2=1.805
r40 18 20 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.64
+ $X2=1.14 $Y2=1.475
r41 12 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.64 $X2=1.15 $Y2=1.64
r42 11 12 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.15 $Y=1.295
+ $X2=1.15 $Y2=1.64
r43 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=0.925
+ $X2=1.15 $Y2=1.295
r44 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=0.555
+ $X2=1.15 $Y2=0.925
r45 7 20 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=1.21 $Y=0.69
+ $X2=1.21 $Y2=1.475
r46 3 21 285.702 $w=1.8e-07 $l=7.35e-07 $layer=POLY_cond $X=1.055 $Y=2.54
+ $X2=1.055 $Y2=1.805
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_1%C 3 6 9 10 11 12 13 14 15 21
c40 12 0 1.66221e-19 $X=1.68 $Y=0.555
c41 6 0 8.74143e-20 $X=1.765 $Y=2.54
r42 14 15 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.69 $Y=1.285
+ $X2=1.69 $Y2=1.665
r43 14 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.69
+ $Y=1.285 $X2=1.69 $Y2=1.285
r44 13 14 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.69 $Y=0.925
+ $X2=1.69 $Y2=1.285
r45 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.69 $Y=0.555
+ $X2=1.69 $Y2=0.925
r46 10 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.69 $Y=1.625
+ $X2=1.69 $Y2=1.285
r47 10 11 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.625
+ $X2=1.69 $Y2=1.79
r48 9 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.12
+ $X2=1.69 $Y2=1.285
r49 6 11 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=1.765 $Y=2.54
+ $X2=1.765 $Y2=1.79
r50 3 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.6 $Y=0.69 $X2=1.6
+ $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_1%D 3 7 9 12 13
c43 7 0 3.01287e-19 $X=2.265 $Y=2.54
r44 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.515
+ $X2=2.23 $Y2=1.68
r45 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.515
+ $X2=2.23 $Y2=1.35
r46 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=1.515 $X2=2.23 $Y2=1.515
r47 9 13 4.93904 $w=3.48e-07 $l=1.5e-07 $layer=LI1_cond $X=2.22 $Y=1.665
+ $X2=2.22 $Y2=1.515
r48 7 15 334.29 $w=1.8e-07 $l=8.6e-07 $layer=POLY_cond $X=2.265 $Y=2.54
+ $X2=2.265 $Y2=1.68
r49 3 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.17 $Y=0.69 $X2=2.17
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_1%A_96_74# 1 2 3 12 16 19 20 21 24 26 30 32 35
+ 39 41 42 46 52
r98 47 52 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=2.77 $Y=1.485 $X2=2.85
+ $Y2=1.485
r99 47 49 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.77 $Y=1.485 $X2=2.68
+ $Y2=1.485
r100 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.485 $X2=2.77 $Y2=1.485
r101 43 46 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.655 $Y=1.485
+ $X2=2.77 $Y2=1.485
r102 36 39 8.74444 $w=5.93e-07 $l=4.35e-07 $layer=LI1_cond $X=0.17 $Y=0.652
+ $X2=0.605 $Y2=0.652
r103 34 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=1.65
+ $X2=2.655 $Y2=1.485
r104 34 35 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.655 $Y=1.65
+ $X2=2.655 $Y2=1.96
r105 33 42 8.61065 $w=1.7e-07 $l=1.68464e-07 $layer=LI1_cond $X=2.205 $Y=2.045
+ $X2=2.04 $Y2=2.052
r106 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.57 $Y=2.045
+ $X2=2.655 $Y2=1.96
r107 32 33 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.57 $Y=2.045
+ $X2=2.205 $Y2=2.045
r108 28 42 0.89609 $w=3.3e-07 $l=9.3e-08 $layer=LI1_cond $X=2.04 $Y=2.145
+ $X2=2.04 $Y2=2.052
r109 28 30 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=2.04 $Y=2.145
+ $X2=2.04 $Y2=2.28
r110 27 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=2.06
+ $X2=0.78 $Y2=2.06
r111 26 42 8.61065 $w=1.7e-07 $l=1.68953e-07 $layer=LI1_cond $X=1.875 $Y=2.06
+ $X2=2.04 $Y2=2.052
r112 26 27 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=1.875 $Y=2.06
+ $X2=0.945 $Y2=2.06
r113 22 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=2.145
+ $X2=0.78 $Y2=2.06
r114 22 24 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.78 $Y=2.145
+ $X2=0.78 $Y2=2.28
r115 20 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=2.06
+ $X2=0.78 $Y2=2.06
r116 20 21 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.615 $Y=2.06
+ $X2=0.255 $Y2=2.06
r117 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=1.975
+ $X2=0.255 $Y2=2.06
r118 18 36 8.26286 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=0.17 $Y=0.95
+ $X2=0.17 $Y2=0.652
r119 18 19 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=0.17 $Y=0.95
+ $X2=0.17 $Y2=1.975
r120 14 52 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.85 $Y=1.65
+ $X2=2.85 $Y2=1.485
r121 14 16 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=2.85 $Y=1.65
+ $X2=2.85 $Y2=2.4
r122 10 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.32
+ $X2=2.68 $Y2=1.485
r123 10 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.68 $Y=1.32
+ $X2=2.68 $Y2=0.74
r124 3 30 300 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_PDIFF $count=2 $X=1.855
+ $Y=2.12 $X2=2.04 $Y2=2.28
r125 2 24 300 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=2 $X=0.645
+ $Y=2.12 $X2=0.78 $Y2=2.28
r126 1 39 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.48
+ $Y=0.37 $X2=0.605 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_1%VPWR 1 2 3 10 12 16 20 22 24 29 36 37 43 46
r49 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 37 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 34 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.74 $Y=3.33
+ $X2=2.575 $Y2=3.33
r55 34 36 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.74 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r58 30 43 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=1.705 $Y=3.33
+ $X2=1.41 $Y2=3.33
r59 30 32 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.705 $Y=3.33
+ $X2=2.16 $Y2=3.33
r60 29 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.41 $Y=3.33
+ $X2=2.575 $Y2=3.33
r61 29 32 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.41 $Y=3.33
+ $X2=2.16 $Y2=3.33
r62 28 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r63 28 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r64 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r65 25 40 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r66 25 27 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r67 24 43 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=1.41 $Y2=3.33
r68 24 27 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=0.72 $Y2=3.33
r69 22 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r70 22 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r71 18 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.575 $Y=3.245
+ $X2=2.575 $Y2=3.33
r72 18 20 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=2.575 $Y=3.245
+ $X2=2.575 $Y2=2.465
r73 14 43 2.48142 $w=5.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.41 $Y=3.245
+ $X2=1.41 $Y2=3.33
r74 14 16 16.4207 $w=5.88e-07 $l=8.1e-07 $layer=LI1_cond $X=1.41 $Y=3.245
+ $X2=1.41 $Y2=2.435
r75 10 40 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r76 10 12 28.2872 $w=3.28e-07 $l=8.1e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.435
r77 3 20 300 $w=1.7e-07 $l=4.41503e-07 $layer=licon1_PDIFF $count=2 $X=2.355
+ $Y=2.12 $X2=2.575 $Y2=2.465
r78 2 16 300 $w=1.7e-07 $l=4.27434e-07 $layer=licon1_PDIFF $count=2 $X=1.145
+ $Y=2.12 $X2=1.41 $Y2=2.435
r79 1 12 300 $w=1.7e-07 $l=3.80657e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_1%X 1 2 9 14 15 16 17 21
c24 14 0 1.35066e-19 $X=3.075 $Y=1.985
r25 17 27 10.6778 $w=5.43e-07 $l=2.05e-07 $layer=LI1_cond $X=3.002 $Y=0.925
+ $X2=3.002 $Y2=1.13
r26 16 17 8.12016 $w=5.43e-07 $l=3.7e-07 $layer=LI1_cond $X=3.002 $Y=0.555
+ $X2=3.002 $Y2=0.925
r27 16 21 0.877856 $w=5.43e-07 $l=4e-08 $layer=LI1_cond $X=3.002 $Y=0.555
+ $X2=3.002 $Y2=0.515
r28 15 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.19 $Y=1.82 $X2=3.19
+ $Y2=1.13
r29 14 15 8.52431 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=3.092 $Y=1.985
+ $X2=3.092 $Y2=1.82
r30 7 14 0.536754 $w=3.63e-07 $l=1.7e-08 $layer=LI1_cond $X=3.092 $Y=2.002
+ $X2=3.092 $Y2=1.985
r31 7 9 25.6695 $w=3.63e-07 $l=8.13e-07 $layer=LI1_cond $X=3.092 $Y=2.002
+ $X2=3.092 $Y2=2.815
r32 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=1.84 $X2=3.075 $Y2=1.985
r33 2 9 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=1.84 $X2=3.075 $Y2=2.815
r34 1 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.755
+ $Y=0.37 $X2=2.895 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__AND4_1%VGND 1 6 9 10 11 21 22
r30 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r31 19 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r32 18 19 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r33 14 18 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r34 14 15 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r35 11 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r36 11 15 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r37 9 18 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.16
+ $Y2=0
r38 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.385
+ $Y2=0
r39 8 21 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.55 $Y=0 $X2=3.12
+ $Y2=0
r40 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.55 $Y=0 $X2=2.385
+ $Y2=0
r41 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=0.085
+ $X2=2.385 $Y2=0
r42 4 6 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.385 $Y=0.085
+ $X2=2.385 $Y2=0.515
r43 1 6 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.245
+ $Y=0.37 $X2=2.385 $Y2=0.515
.ends


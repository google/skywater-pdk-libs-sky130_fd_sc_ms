* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfrbp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_27_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X1 VGND a_819_119# a_1037_119# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 a_1399_119# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 VGND a_1747_74# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VPWR RESET_B a_1235_119# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X5 a_413_90# SCE a_545_97# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X6 a_1235_119# a_1037_119# a_1321_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X7 a_819_119# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 a_1369_93# a_819_119# a_1747_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X9 VGND a_2513_424# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_545_97# SCD a_225_90# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X11 a_413_90# a_1037_119# a_1235_119# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X12 a_2008_48# a_1747_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X13 VPWR SCE a_341_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X14 VPWR a_819_119# a_1037_119# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 a_1235_119# a_819_119# a_1331_463# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X16 a_2513_424# a_1747_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X17 VGND RESET_B a_2124_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X18 a_413_90# a_819_119# a_1235_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X19 a_1966_74# a_2008_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X20 a_413_90# a_27_74# a_515_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X21 a_1321_119# a_1369_93# a_1399_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X22 a_312_90# D a_413_90# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X23 a_2513_424# a_1747_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X24 a_1331_463# a_1369_93# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X25 a_1747_74# a_819_119# a_1966_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X26 VPWR a_1235_119# a_1369_93# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X27 a_819_119# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X28 a_515_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X29 VPWR a_1747_74# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X30 VPWR RESET_B a_2008_48# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X31 a_2124_74# a_1747_74# a_2008_48# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X32 a_1369_93# a_1037_119# a_1747_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X33 a_225_90# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X34 VGND a_1235_119# a_1369_93# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X35 VPWR RESET_B a_413_90# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X36 a_225_90# a_27_74# a_312_90# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X37 a_341_464# D a_413_90# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X38 a_27_74# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X39 a_1747_74# a_1037_119# a_1972_489# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X40 a_1972_489# a_2008_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X41 VPWR a_2513_424# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
.ends

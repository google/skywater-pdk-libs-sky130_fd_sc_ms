* File: sky130_fd_sc_ms__clkinv_1.pxi.spice
* Created: Wed Sep  2 12:01:34 2020
* 
x_PM_SKY130_FD_SC_MS__CLKINV_1%A N_A_M1001_g N_A_M1000_g N_A_M1002_g A A
+ N_A_c_28_n N_A_c_29_n N_A_c_30_n PM_SKY130_FD_SC_MS__CLKINV_1%A
x_PM_SKY130_FD_SC_MS__CLKINV_1%VPWR N_VPWR_M1001_s N_VPWR_M1002_s N_VPWR_c_60_n
+ N_VPWR_c_61_n N_VPWR_c_62_n N_VPWR_c_63_n VPWR N_VPWR_c_64_n N_VPWR_c_59_n
+ PM_SKY130_FD_SC_MS__CLKINV_1%VPWR
x_PM_SKY130_FD_SC_MS__CLKINV_1%Y N_Y_M1000_d N_Y_M1001_d N_Y_c_84_n N_Y_c_79_n Y
+ Y Y Y Y N_Y_c_81_n Y N_Y_c_83_n PM_SKY130_FD_SC_MS__CLKINV_1%Y
x_PM_SKY130_FD_SC_MS__CLKINV_1%VGND N_VGND_M1000_s N_VGND_c_105_n N_VGND_c_106_n
+ VGND N_VGND_c_107_n N_VGND_c_108_n PM_SKY130_FD_SC_MS__CLKINV_1%VGND
cc_1 VNB N_A_M1000_g 0.027297f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.58
cc_2 VNB A 0.0282826f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_3 VNB N_A_c_28_n 0.0453666f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.425
cc_4 VNB N_A_c_29_n 0.0578814f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.085
cc_5 VNB N_A_c_30_n 0.00540078f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.765
cc_6 VNB N_VPWR_c_59_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.765
cc_7 VNB N_Y_c_79_n 0.00750462f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.54
cc_8 VNB Y 0.0520536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_Y_c_81_n 0.0160574f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.765
cc_10 VNB N_VGND_c_105_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_VGND_c_106_n 0.0282119f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.58
cc_12 VNB N_VGND_c_107_n 0.0282669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_VGND_c_108_n 0.11676f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_14 VPB N_A_M1001_g 0.0289261f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.54
cc_15 VPB N_A_M1002_g 0.0251919f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.54
cc_16 VPB A 0.0108313f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_17 VPB N_A_c_30_n 0.0388458f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.765
cc_18 VPB N_VPWR_c_60_n 0.0103331f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.58
cc_19 VPB N_VPWR_c_61_n 0.0473151f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.93
cc_20 VPB N_VPWR_c_62_n 0.0116777f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.54
cc_21 VPB N_VPWR_c_63_n 0.0237119f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_22 VPB N_VPWR_c_64_n 0.0183948f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.235
cc_23 VPB N_VPWR_c_59_n 0.0487345f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.765
cc_24 VPB Y 0.0230423f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_25 VPB N_Y_c_83_n 0.0211992f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_26 N_A_M1001_g N_VPWR_c_61_n 0.00751355f $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_27 A N_VPWR_c_61_n 0.0136621f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_28 N_A_M1001_g N_VPWR_c_63_n 3.98302e-19 $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_29 N_A_M1002_g N_VPWR_c_63_n 0.0102983f $X=0.945 $Y=2.54 $X2=0 $Y2=0
cc_30 N_A_M1001_g N_VPWR_c_64_n 0.00521549f $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_31 N_A_M1002_g N_VPWR_c_64_n 0.00460063f $X=0.945 $Y=2.54 $X2=0 $Y2=0
cc_32 N_A_M1001_g N_VPWR_c_59_n 0.00986531f $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_33 N_A_M1002_g N_VPWR_c_59_n 0.00908554f $X=0.945 $Y=2.54 $X2=0 $Y2=0
cc_34 N_A_M1001_g N_Y_c_84_n 0.00823914f $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_35 N_A_M1000_g N_Y_c_79_n 0.00458999f $X=0.565 $Y=0.58 $X2=0 $Y2=0
cc_36 A N_Y_c_79_n 0.00696579f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_37 N_A_c_29_n N_Y_c_79_n 0.0121436f $X=0.59 $Y=1.085 $X2=0 $Y2=0
cc_38 N_A_M1000_g Y 0.00534936f $X=0.565 $Y=0.58 $X2=0 $Y2=0
cc_39 A Y 0.0489624f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_40 N_A_c_29_n Y 0.0394859f $X=0.59 $Y=1.085 $X2=0 $Y2=0
cc_41 N_A_M1001_g N_Y_c_83_n 0.00492104f $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_42 N_A_M1002_g N_Y_c_83_n 0.0282018f $X=0.945 $Y=2.54 $X2=0 $Y2=0
cc_43 A N_Y_c_83_n 0.0166619f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_44 N_A_c_30_n N_Y_c_83_n 0.00102886f $X=0.59 $Y=1.765 $X2=0 $Y2=0
cc_45 N_A_M1000_g N_VGND_c_106_n 0.0124698f $X=0.565 $Y=0.58 $X2=0 $Y2=0
cc_46 A N_VGND_c_106_n 0.0151075f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_47 N_A_c_29_n N_VGND_c_106_n 7.38054e-19 $X=0.59 $Y=1.085 $X2=0 $Y2=0
cc_48 N_A_M1000_g N_VGND_c_107_n 0.00433162f $X=0.565 $Y=0.58 $X2=0 $Y2=0
cc_49 N_A_M1000_g N_VGND_c_108_n 0.00825282f $X=0.565 $Y=0.58 $X2=0 $Y2=0
cc_50 N_VPWR_c_64_n N_Y_c_84_n 0.00904111f $X=1.005 $Y=3.33 $X2=0 $Y2=0
cc_51 N_VPWR_c_59_n N_Y_c_84_n 0.00986687f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_52 N_VPWR_M1002_s N_Y_c_83_n 0.00385022f $X=1.035 $Y=2.12 $X2=0 $Y2=0
cc_53 N_VPWR_c_61_n N_Y_c_83_n 0.0127651f $X=0.27 $Y=2.265 $X2=0 $Y2=0
cc_54 N_VPWR_c_63_n N_Y_c_83_n 0.0221401f $X=1.17 $Y=2.79 $X2=0 $Y2=0
cc_55 N_Y_c_79_n N_VGND_c_106_n 0.0146598f $X=1.085 $Y=0.515 $X2=0 $Y2=0
cc_56 N_Y_c_79_n N_VGND_c_107_n 0.0197467f $X=1.085 $Y=0.515 $X2=0 $Y2=0
cc_57 N_Y_c_81_n N_VGND_c_107_n 0.010709f $X=1.205 $Y=0.68 $X2=0 $Y2=0
cc_58 N_Y_c_79_n N_VGND_c_108_n 0.0168182f $X=1.085 $Y=0.515 $X2=0 $Y2=0
cc_59 N_Y_c_81_n N_VGND_c_108_n 0.008864f $X=1.205 $Y=0.68 $X2=0 $Y2=0

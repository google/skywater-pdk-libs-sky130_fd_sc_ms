* File: sky130_fd_sc_ms__o22a_1.pxi.spice
* Created: Wed Sep  2 12:23:29 2020
* 
x_PM_SKY130_FD_SC_MS__O22A_1%A_83_260# N_A_83_260#_M1003_d N_A_83_260#_M1007_d
+ N_A_83_260#_M1002_g N_A_83_260#_M1009_g N_A_83_260#_c_63_n N_A_83_260#_c_108_p
+ N_A_83_260#_c_64_n N_A_83_260#_c_70_n N_A_83_260#_c_65_n N_A_83_260#_c_66_n
+ N_A_83_260#_c_67_n N_A_83_260#_c_75_p N_A_83_260#_c_77_p
+ PM_SKY130_FD_SC_MS__O22A_1%A_83_260#
x_PM_SKY130_FD_SC_MS__O22A_1%B1 N_B1_M1003_g N_B1_M1005_g B1 N_B1_c_139_n
+ N_B1_c_140_n PM_SKY130_FD_SC_MS__O22A_1%B1
x_PM_SKY130_FD_SC_MS__O22A_1%B2 N_B2_c_175_n N_B2_M1007_g N_B2_M1006_g
+ N_B2_c_178_n N_B2_c_179_n B2 N_B2_c_180_n PM_SKY130_FD_SC_MS__O22A_1%B2
x_PM_SKY130_FD_SC_MS__O22A_1%A2 N_A2_M1004_g N_A2_M1008_g A2 N_A2_c_222_n
+ N_A2_c_223_n PM_SKY130_FD_SC_MS__O22A_1%A2
x_PM_SKY130_FD_SC_MS__O22A_1%A1 N_A1_M1001_g N_A1_M1000_g A1 N_A1_c_263_n
+ PM_SKY130_FD_SC_MS__O22A_1%A1
x_PM_SKY130_FD_SC_MS__O22A_1%X N_X_M1009_s N_X_M1002_s N_X_c_288_n N_X_c_289_n X
+ X X X N_X_c_290_n PM_SKY130_FD_SC_MS__O22A_1%X
x_PM_SKY130_FD_SC_MS__O22A_1%VPWR N_VPWR_M1002_d N_VPWR_M1001_d N_VPWR_c_309_n
+ N_VPWR_c_310_n N_VPWR_c_311_n VPWR N_VPWR_c_312_n N_VPWR_c_313_n
+ N_VPWR_c_314_n N_VPWR_c_308_n PM_SKY130_FD_SC_MS__O22A_1%VPWR
x_PM_SKY130_FD_SC_MS__O22A_1%VGND N_VGND_M1009_d N_VGND_M1004_d N_VGND_c_349_n
+ N_VGND_c_350_n VGND N_VGND_c_351_n N_VGND_c_352_n N_VGND_c_353_n
+ N_VGND_c_354_n N_VGND_c_355_n N_VGND_c_356_n PM_SKY130_FD_SC_MS__O22A_1%VGND
x_PM_SKY130_FD_SC_MS__O22A_1%A_299_139# N_A_299_139#_M1003_s
+ N_A_299_139#_M1006_d N_A_299_139#_M1000_d N_A_299_139#_c_389_n
+ N_A_299_139#_c_405_n N_A_299_139#_c_396_n N_A_299_139#_c_390_n
+ N_A_299_139#_c_397_n N_A_299_139#_c_391_n
+ PM_SKY130_FD_SC_MS__O22A_1%A_299_139#
cc_1 VNB N_A_83_260#_M1002_g 0.00260026f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A_83_260#_M1009_g 0.0298754f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_3 VNB N_A_83_260#_c_63_n 0.0158547f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_4 VNB N_A_83_260#_c_64_n 0.00260369f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=1.97
cc_5 VNB N_A_83_260#_c_65_n 0.0107741f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=1.215
cc_6 VNB N_A_83_260#_c_66_n 0.0553097f $X=-0.19 $Y=-0.245 $X2=0.93 $Y2=1.465
cc_7 VNB N_A_83_260#_c_67_n 0.0173604f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.202
cc_8 VNB N_B1_M1003_g 0.0219239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B1_c_139_n 0.0384003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B1_c_140_n 0.00479522f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.465
cc_11 VNB N_B2_c_175_n 0.0055117f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=0.695
cc_12 VNB N_B2_M1007_g 0.00838156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B2_M1006_g 0.00974696f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_14 VNB N_B2_c_178_n 0.0230388f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_15 VNB N_B2_c_179_n 0.0422378f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_16 VNB N_B2_c_180_n 0.0123671f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=2.14
cc_17 VNB N_A2_M1004_g 0.0204256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A2_c_222_n 0.016352f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_19 VNB N_A2_c_223_n 0.0040305f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_20 VNB N_A1_M1000_g 0.0309121f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.63
cc_21 VNB A1 0.0101032f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_22 VNB N_A1_c_263_n 0.0186679f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_23 VNB N_X_c_288_n 0.027165f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_24 VNB N_X_c_289_n 0.0101198f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_25 VNB N_X_c_290_n 0.0250186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_308_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_349_n 0.0175259f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_28 VNB N_VGND_c_350_n 0.0272042f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_29 VNB N_VGND_c_351_n 0.0171566f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_30 VNB N_VGND_c_352_n 0.0498673f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=1.97
cc_31 VNB N_VGND_c_353_n 0.020239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_354_n 0.248297f $X=-0.19 $Y=-0.245 $X2=2.09 $Y2=1.202
cc_33 VNB N_VGND_c_355_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=2.26 $Y2=1.202
cc_34 VNB N_VGND_c_356_n 0.00653982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_299_139#_c_389_n 0.00337111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_299_139#_c_390_n 0.0152494f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_37 VNB N_A_299_139#_c_391_n 0.023023f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.215
cc_38 VPB N_A_83_260#_M1002_g 0.0347152f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_39 VPB N_A_83_260#_c_64_n 0.00228663f $X=-0.19 $Y=1.66 $X2=2.26 $Y2=1.97
cc_40 VPB N_A_83_260#_c_70_n 0.00231613f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=2.815
cc_41 VPB N_B1_M1005_g 0.0278485f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_42 VPB N_B1_c_139_n 0.031934f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_B1_c_140_n 0.00465035f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.465
cc_44 VPB N_B2_M1007_g 0.0270817f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A2_M1008_g 0.0232991f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.63
cc_46 VPB N_A2_c_222_n 0.0141338f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_47 VPB N_A2_c_223_n 0.00292555f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_48 VPB N_A1_M1001_g 0.0291537f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB A1 0.00778911f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_50 VPB N_A1_c_263_n 0.0141222f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_51 VPB X 0.0136968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB X 0.0415472f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=2.14
cc_53 VPB N_X_c_290_n 0.00769959f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_309_n 0.0160367f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_55 VPB N_VPWR_c_310_n 0.0123157f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_56 VPB N_VPWR_c_311_n 0.0477013f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_312_n 0.0189171f $X=-0.19 $Y=1.66 $X2=2.56 $Y2=2.815
cc_58 VPB N_VPWR_c_313_n 0.0459048f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=1.465
cc_59 VPB N_VPWR_c_314_n 0.0235395f $X=-0.19 $Y=1.66 $X2=2.26 $Y2=2.055
cc_60 VPB N_VPWR_c_308_n 0.07397f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 N_A_83_260#_c_64_n N_B1_M1003_g 0.00315367f $X=2.26 $Y=1.97 $X2=0 $Y2=0
cc_62 N_A_83_260#_c_65_n N_B1_M1003_g 0.0010886f $X=1.01 $Y=1.215 $X2=0 $Y2=0
cc_63 N_A_83_260#_c_66_n N_B1_M1003_g 0.00347063f $X=0.93 $Y=1.465 $X2=0 $Y2=0
cc_64 N_A_83_260#_c_67_n N_B1_M1003_g 0.00946308f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_65 N_A_83_260#_c_75_p N_B1_M1003_g 0.0021184f $X=2.26 $Y=1.202 $X2=0 $Y2=0
cc_66 N_A_83_260#_c_70_n N_B1_M1005_g 0.00238694f $X=2.56 $Y=2.815 $X2=0 $Y2=0
cc_67 N_A_83_260#_c_77_p N_B1_M1005_g 0.00162162f $X=2.56 $Y=2.135 $X2=0 $Y2=0
cc_68 N_A_83_260#_c_64_n N_B1_c_139_n 0.0055332f $X=2.26 $Y=1.97 $X2=0 $Y2=0
cc_69 N_A_83_260#_c_65_n N_B1_c_139_n 6.76009e-19 $X=1.01 $Y=1.215 $X2=0 $Y2=0
cc_70 N_A_83_260#_c_66_n N_B1_c_139_n 0.00922917f $X=0.93 $Y=1.465 $X2=0 $Y2=0
cc_71 N_A_83_260#_c_67_n N_B1_c_139_n 0.00300073f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_72 N_A_83_260#_c_75_p N_B1_c_139_n 3.91515e-19 $X=2.26 $Y=1.202 $X2=0 $Y2=0
cc_73 N_A_83_260#_c_64_n N_B1_c_140_n 0.0262171f $X=2.26 $Y=1.97 $X2=0 $Y2=0
cc_74 N_A_83_260#_c_65_n N_B1_c_140_n 0.00919512f $X=1.01 $Y=1.215 $X2=0 $Y2=0
cc_75 N_A_83_260#_c_66_n N_B1_c_140_n 6.74389e-19 $X=0.93 $Y=1.465 $X2=0 $Y2=0
cc_76 N_A_83_260#_c_67_n N_B1_c_140_n 0.0452308f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_77 N_A_83_260#_c_64_n N_B2_c_175_n 0.00243203f $X=2.26 $Y=1.97 $X2=-0.19
+ $Y2=-0.245
cc_78 N_A_83_260#_c_64_n N_B2_M1007_g 0.0110807f $X=2.26 $Y=1.97 $X2=0 $Y2=0
cc_79 N_A_83_260#_c_70_n N_B2_M1007_g 0.016214f $X=2.56 $Y=2.815 $X2=0 $Y2=0
cc_80 N_A_83_260#_c_77_p N_B2_M1007_g 0.0140685f $X=2.56 $Y=2.135 $X2=0 $Y2=0
cc_81 N_A_83_260#_c_64_n N_B2_M1006_g 0.00319876f $X=2.26 $Y=1.97 $X2=0 $Y2=0
cc_82 N_A_83_260#_c_75_p N_B2_M1006_g 0.00453123f $X=2.26 $Y=1.202 $X2=0 $Y2=0
cc_83 N_A_83_260#_c_67_n N_B2_c_178_n 0.00599251f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_84 N_A_83_260#_M1009_g N_B2_c_180_n 0.00103253f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_85 N_A_83_260#_c_65_n N_B2_c_180_n 3.962e-19 $X=1.01 $Y=1.215 $X2=0 $Y2=0
cc_86 N_A_83_260#_c_67_n N_B2_c_180_n 0.00852348f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_87 N_A_83_260#_c_64_n N_A2_M1004_g 9.40991e-19 $X=2.26 $Y=1.97 $X2=0 $Y2=0
cc_88 N_A_83_260#_c_64_n N_A2_M1008_g 9.07119e-19 $X=2.26 $Y=1.97 $X2=0 $Y2=0
cc_89 N_A_83_260#_c_70_n N_A2_M1008_g 0.0182387f $X=2.56 $Y=2.815 $X2=0 $Y2=0
cc_90 N_A_83_260#_c_77_p N_A2_M1008_g 0.0040238f $X=2.56 $Y=2.135 $X2=0 $Y2=0
cc_91 N_A_83_260#_c_64_n N_A2_c_222_n 2.87256e-19 $X=2.26 $Y=1.97 $X2=0 $Y2=0
cc_92 N_A_83_260#_c_64_n N_A2_c_223_n 0.0245237f $X=2.26 $Y=1.97 $X2=0 $Y2=0
cc_93 N_A_83_260#_c_77_p N_A2_c_223_n 0.0131668f $X=2.56 $Y=2.135 $X2=0 $Y2=0
cc_94 N_A_83_260#_c_70_n N_A1_M1001_g 0.00259267f $X=2.56 $Y=2.815 $X2=0 $Y2=0
cc_95 N_A_83_260#_c_77_p N_A1_M1001_g 5.17764e-19 $X=2.56 $Y=2.135 $X2=0 $Y2=0
cc_96 N_A_83_260#_M1009_g N_X_c_288_n 0.00239685f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_97 N_A_83_260#_M1002_g X 0.00871641f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_98 N_A_83_260#_c_108_p X 0.00138666f $X=0.925 $Y=1.465 $X2=0 $Y2=0
cc_99 N_A_83_260#_M1002_g X 0.0132074f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_100 N_A_83_260#_M1009_g N_X_c_290_n 0.00288366f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_101 N_A_83_260#_c_63_n N_X_c_290_n 0.0136309f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_102 N_A_83_260#_c_108_p N_X_c_290_n 0.0255805f $X=0.925 $Y=1.465 $X2=0 $Y2=0
cc_103 N_A_83_260#_c_65_n N_X_c_290_n 0.00347497f $X=1.01 $Y=1.215 $X2=0 $Y2=0
cc_104 N_A_83_260#_M1002_g N_VPWR_c_309_n 0.00585939f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_105 N_A_83_260#_c_108_p N_VPWR_c_309_n 0.0135501f $X=0.925 $Y=1.465 $X2=0
+ $Y2=0
cc_106 N_A_83_260#_c_70_n N_VPWR_c_309_n 0.0256466f $X=2.56 $Y=2.815 $X2=0 $Y2=0
cc_107 N_A_83_260#_c_65_n N_VPWR_c_309_n 0.00812676f $X=1.01 $Y=1.215 $X2=0
+ $Y2=0
cc_108 N_A_83_260#_c_66_n N_VPWR_c_309_n 0.00753152f $X=0.93 $Y=1.465 $X2=0
+ $Y2=0
cc_109 N_A_83_260#_c_77_p N_VPWR_c_309_n 0.00800091f $X=2.56 $Y=2.135 $X2=0
+ $Y2=0
cc_110 N_A_83_260#_c_70_n N_VPWR_c_311_n 0.0203083f $X=2.56 $Y=2.815 $X2=0 $Y2=0
cc_111 N_A_83_260#_c_77_p N_VPWR_c_311_n 0.00423395f $X=2.56 $Y=2.135 $X2=0
+ $Y2=0
cc_112 N_A_83_260#_M1002_g N_VPWR_c_312_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_113 N_A_83_260#_c_70_n N_VPWR_c_313_n 0.0144623f $X=2.56 $Y=2.815 $X2=0 $Y2=0
cc_114 N_A_83_260#_M1002_g N_VPWR_c_308_n 0.00990469f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_115 N_A_83_260#_c_70_n N_VPWR_c_308_n 0.0118344f $X=2.56 $Y=2.815 $X2=0 $Y2=0
cc_116 N_A_83_260#_c_77_p A_401_392# 0.0024232f $X=2.56 $Y=2.135 $X2=-0.19
+ $Y2=-0.245
cc_117 N_A_83_260#_M1009_g N_VGND_c_349_n 0.0149103f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_118 N_A_83_260#_c_63_n N_VGND_c_349_n 0.00622694f $X=0.505 $Y=1.465 $X2=0
+ $Y2=0
cc_119 N_A_83_260#_c_108_p N_VGND_c_349_n 0.014292f $X=0.925 $Y=1.465 $X2=0
+ $Y2=0
cc_120 N_A_83_260#_M1009_g N_VGND_c_351_n 0.00383152f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_121 N_A_83_260#_M1009_g N_VGND_c_354_n 0.00761198f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_122 N_A_83_260#_c_67_n N_A_299_139#_M1003_s 0.00440797f $X=1.905 $Y=1.202
+ $X2=-0.19 $Y2=-0.245
cc_123 N_A_83_260#_M1003_d N_A_299_139#_c_389_n 0.00421372f $X=1.93 $Y=0.695
+ $X2=0 $Y2=0
cc_124 N_A_83_260#_c_67_n N_A_299_139#_c_389_n 0.0240084f $X=1.905 $Y=1.202
+ $X2=0 $Y2=0
cc_125 N_A_83_260#_c_75_p N_A_299_139#_c_389_n 0.0233695f $X=2.26 $Y=1.202 $X2=0
+ $Y2=0
cc_126 N_A_83_260#_c_75_p N_A_299_139#_c_396_n 0.00163712f $X=2.26 $Y=1.202
+ $X2=0 $Y2=0
cc_127 N_A_83_260#_c_75_p N_A_299_139#_c_397_n 0.0135439f $X=2.26 $Y=1.202 $X2=0
+ $Y2=0
cc_128 N_B1_M1003_g N_B2_c_175_n 0.00209685f $X=1.855 $Y=1.015 $X2=-0.19
+ $Y2=-0.245
cc_129 N_B1_c_139_n N_B2_c_175_n 0.0418793f $X=1.84 $Y=1.635 $X2=-0.19
+ $Y2=-0.245
cc_130 N_B1_c_140_n N_B2_c_175_n 3.6513e-19 $X=1.84 $Y=1.635 $X2=-0.19
+ $Y2=-0.245
cc_131 N_B1_M1005_g N_B2_M1007_g 0.0418793f $X=1.915 $Y=2.46 $X2=0 $Y2=0
cc_132 N_B1_M1003_g N_B2_M1006_g 0.0194929f $X=1.855 $Y=1.015 $X2=0 $Y2=0
cc_133 N_B1_M1003_g N_B2_c_178_n 0.00604329f $X=1.855 $Y=1.015 $X2=0 $Y2=0
cc_134 N_B1_M1003_g N_B2_c_179_n 0.00129799f $X=1.855 $Y=1.015 $X2=0 $Y2=0
cc_135 N_B1_M1003_g N_B2_c_180_n 0.00215635f $X=1.855 $Y=1.015 $X2=0 $Y2=0
cc_136 N_B1_M1005_g N_VPWR_c_309_n 0.0236744f $X=1.915 $Y=2.46 $X2=0 $Y2=0
cc_137 N_B1_c_139_n N_VPWR_c_309_n 0.00363808f $X=1.84 $Y=1.635 $X2=0 $Y2=0
cc_138 N_B1_c_140_n N_VPWR_c_309_n 0.0373097f $X=1.84 $Y=1.635 $X2=0 $Y2=0
cc_139 N_B1_M1005_g N_VPWR_c_313_n 0.00475445f $X=1.915 $Y=2.46 $X2=0 $Y2=0
cc_140 N_B1_M1005_g N_VPWR_c_308_n 0.00938478f $X=1.915 $Y=2.46 $X2=0 $Y2=0
cc_141 N_B1_M1003_g N_VGND_c_352_n 4.64175e-19 $X=1.855 $Y=1.015 $X2=0 $Y2=0
cc_142 N_B1_M1003_g N_A_299_139#_c_389_n 0.00901709f $X=1.855 $Y=1.015 $X2=0
+ $Y2=0
cc_143 N_B2_c_175_n N_A2_M1004_g 0.00300985f $X=2.335 $Y=1.5 $X2=0 $Y2=0
cc_144 N_B2_M1006_g N_A2_M1004_g 0.0204823f $X=2.325 $Y=1.015 $X2=0 $Y2=0
cc_145 N_B2_c_179_n N_A2_M1004_g 0.00120024f $X=2.305 $Y=0.42 $X2=0 $Y2=0
cc_146 N_B2_M1007_g N_A2_M1008_g 0.0145683f $X=2.335 $Y=2.46 $X2=0 $Y2=0
cc_147 N_B2_c_175_n N_A2_c_222_n 0.0165024f $X=2.335 $Y=1.5 $X2=0 $Y2=0
cc_148 N_B2_c_175_n N_A2_c_223_n 0.00224417f $X=2.335 $Y=1.5 $X2=0 $Y2=0
cc_149 N_B2_M1007_g N_VPWR_c_309_n 0.00303026f $X=2.335 $Y=2.46 $X2=0 $Y2=0
cc_150 N_B2_M1007_g N_VPWR_c_313_n 0.005209f $X=2.335 $Y=2.46 $X2=0 $Y2=0
cc_151 N_B2_M1007_g N_VPWR_c_308_n 0.00983291f $X=2.335 $Y=2.46 $X2=0 $Y2=0
cc_152 N_B2_c_180_n N_VGND_c_349_n 0.0309525f $X=1.305 $Y=0.462 $X2=0 $Y2=0
cc_153 N_B2_c_178_n N_VGND_c_350_n 0.0141143f $X=2.305 $Y=0.42 $X2=0 $Y2=0
cc_154 N_B2_c_179_n N_VGND_c_350_n 0.00195451f $X=2.305 $Y=0.42 $X2=0 $Y2=0
cc_155 N_B2_c_179_n N_VGND_c_352_n 0.00783549f $X=2.305 $Y=0.42 $X2=0 $Y2=0
cc_156 N_B2_c_180_n N_VGND_c_352_n 0.0926586f $X=1.305 $Y=0.462 $X2=0 $Y2=0
cc_157 N_B2_c_179_n N_VGND_c_354_n 0.011167f $X=2.305 $Y=0.42 $X2=0 $Y2=0
cc_158 N_B2_c_180_n N_VGND_c_354_n 0.0526994f $X=1.305 $Y=0.462 $X2=0 $Y2=0
cc_159 N_B2_M1006_g N_A_299_139#_c_389_n 0.0105407f $X=2.325 $Y=1.015 $X2=0
+ $Y2=0
cc_160 N_B2_c_178_n N_A_299_139#_c_389_n 0.0649092f $X=2.305 $Y=0.42 $X2=0 $Y2=0
cc_161 N_B2_c_179_n N_A_299_139#_c_389_n 0.00378752f $X=2.305 $Y=0.42 $X2=0
+ $Y2=0
cc_162 N_B2_M1006_g N_A_299_139#_c_396_n 0.00344339f $X=2.325 $Y=1.015 $X2=0
+ $Y2=0
cc_163 N_B2_M1006_g N_A_299_139#_c_397_n 0.00124396f $X=2.325 $Y=1.015 $X2=0
+ $Y2=0
cc_164 N_A2_M1008_g N_A1_M1001_g 0.0426724f $X=2.785 $Y=2.46 $X2=0 $Y2=0
cc_165 N_A2_M1004_g N_A1_M1000_g 0.020765f $X=2.755 $Y=1.015 $X2=0 $Y2=0
cc_166 N_A2_c_222_n A1 4.18174e-19 $X=2.83 $Y=1.635 $X2=0 $Y2=0
cc_167 N_A2_c_223_n A1 0.0199019f $X=2.83 $Y=1.635 $X2=0 $Y2=0
cc_168 N_A2_c_222_n N_A1_c_263_n 0.0181729f $X=2.83 $Y=1.635 $X2=0 $Y2=0
cc_169 N_A2_c_223_n N_A1_c_263_n 4.18284e-19 $X=2.83 $Y=1.635 $X2=0 $Y2=0
cc_170 N_A2_M1008_g N_VPWR_c_311_n 0.00363663f $X=2.785 $Y=2.46 $X2=0 $Y2=0
cc_171 N_A2_M1008_g N_VPWR_c_313_n 0.005209f $X=2.785 $Y=2.46 $X2=0 $Y2=0
cc_172 N_A2_M1008_g N_VPWR_c_308_n 0.00984377f $X=2.785 $Y=2.46 $X2=0 $Y2=0
cc_173 N_A2_M1004_g N_VGND_c_350_n 0.00511389f $X=2.755 $Y=1.015 $X2=0 $Y2=0
cc_174 N_A2_M1004_g N_VGND_c_352_n 0.00367092f $X=2.755 $Y=1.015 $X2=0 $Y2=0
cc_175 N_A2_M1004_g N_VGND_c_354_n 0.0045051f $X=2.755 $Y=1.015 $X2=0 $Y2=0
cc_176 N_A2_c_223_n N_A_299_139#_c_389_n 3.28827e-19 $X=2.83 $Y=1.635 $X2=0
+ $Y2=0
cc_177 N_A2_M1004_g N_A_299_139#_c_405_n 0.00241154f $X=2.755 $Y=1.015 $X2=0
+ $Y2=0
cc_178 N_A2_M1004_g N_A_299_139#_c_396_n 0.00416793f $X=2.755 $Y=1.015 $X2=0
+ $Y2=0
cc_179 N_A2_M1004_g N_A_299_139#_c_390_n 0.011631f $X=2.755 $Y=1.015 $X2=0 $Y2=0
cc_180 N_A2_c_222_n N_A_299_139#_c_390_n 0.00375164f $X=2.83 $Y=1.635 $X2=0
+ $Y2=0
cc_181 N_A2_c_223_n N_A_299_139#_c_390_n 0.0190059f $X=2.83 $Y=1.635 $X2=0 $Y2=0
cc_182 N_A2_M1004_g N_A_299_139#_c_397_n 0.00199254f $X=2.755 $Y=1.015 $X2=0
+ $Y2=0
cc_183 N_A2_c_223_n N_A_299_139#_c_397_n 0.0117835f $X=2.83 $Y=1.635 $X2=0 $Y2=0
cc_184 N_A2_M1004_g N_A_299_139#_c_391_n 8.28157e-19 $X=2.755 $Y=1.015 $X2=0
+ $Y2=0
cc_185 N_A1_M1001_g N_VPWR_c_311_n 0.0270439f $X=3.325 $Y=2.46 $X2=0 $Y2=0
cc_186 A1 N_VPWR_c_311_n 0.0250523f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_187 N_A1_c_263_n N_VPWR_c_311_n 0.00334038f $X=3.4 $Y=1.635 $X2=0 $Y2=0
cc_188 N_A1_M1001_g N_VPWR_c_313_n 0.00460063f $X=3.325 $Y=2.46 $X2=0 $Y2=0
cc_189 N_A1_M1001_g N_VPWR_c_308_n 0.00909457f $X=3.325 $Y=2.46 $X2=0 $Y2=0
cc_190 N_A1_M1000_g N_VGND_c_350_n 0.00599119f $X=3.345 $Y=0.97 $X2=0 $Y2=0
cc_191 N_A1_M1000_g N_VGND_c_353_n 0.00387791f $X=3.345 $Y=0.97 $X2=0 $Y2=0
cc_192 N_A1_M1000_g N_VGND_c_354_n 0.00462577f $X=3.345 $Y=0.97 $X2=0 $Y2=0
cc_193 N_A1_M1000_g N_A_299_139#_c_396_n 7.76236e-19 $X=3.345 $Y=0.97 $X2=0
+ $Y2=0
cc_194 N_A1_M1000_g N_A_299_139#_c_390_n 0.0125821f $X=3.345 $Y=0.97 $X2=0 $Y2=0
cc_195 A1 N_A_299_139#_c_390_n 0.0389835f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_196 N_A1_c_263_n N_A_299_139#_c_390_n 0.00429329f $X=3.4 $Y=1.635 $X2=0 $Y2=0
cc_197 N_A1_M1000_g N_A_299_139#_c_391_n 0.00768327f $X=3.345 $Y=0.97 $X2=0
+ $Y2=0
cc_198 X N_VPWR_c_309_n 0.0386794f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_199 X N_VPWR_c_312_n 0.0158876f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_200 X N_VPWR_c_308_n 0.0130823f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_201 N_X_c_288_n N_VGND_c_349_n 0.0226038f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_202 N_X_c_288_n N_VGND_c_351_n 0.0124046f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_203 N_X_c_288_n N_VGND_c_354_n 0.0102675f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_204 N_VGND_c_349_n N_A_299_139#_c_389_n 0.00653306f $X=0.71 $Y=0.515 $X2=0
+ $Y2=0
cc_205 N_VGND_c_352_n N_A_299_139#_c_389_n 8.81826e-19 $X=2.885 $Y=0 $X2=0 $Y2=0
cc_206 N_VGND_c_354_n N_A_299_139#_c_389_n 0.00320664f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_207 N_VGND_c_352_n N_A_299_139#_c_405_n 0.00205276f $X=2.885 $Y=0 $X2=0 $Y2=0
cc_208 N_VGND_c_354_n N_A_299_139#_c_405_n 0.00462418f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_209 N_VGND_M1004_d N_A_299_139#_c_390_n 0.00832046f $X=2.83 $Y=0.695 $X2=0
+ $Y2=0
cc_210 N_VGND_c_350_n N_A_299_139#_c_390_n 0.0265229f $X=3.055 $Y=0.795 $X2=0
+ $Y2=0
cc_211 N_VGND_c_350_n N_A_299_139#_c_391_n 0.0131765f $X=3.055 $Y=0.795 $X2=0
+ $Y2=0
cc_212 N_VGND_c_353_n N_A_299_139#_c_391_n 0.00664851f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_213 N_VGND_c_354_n N_A_299_139#_c_391_n 0.00995444f $X=3.6 $Y=0 $X2=0 $Y2=0

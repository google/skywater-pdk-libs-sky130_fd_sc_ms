* File: sky130_fd_sc_ms__buf_1.spice
* Created: Fri Aug 28 17:15:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__buf_1.pex.spice"
.subckt sky130_fd_sc_ms__buf_1  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_M1002_g N_A_27_164#_M1002_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.129591 AS=0.24915 PD=0.997674 PS=2.37 NRD=18 NRS=0 M=1 R=3.66667
+ SA=75000.4 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1003 N_X_M1003_d N_A_27_164#_M1003_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_A_27_164#_M1001_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1632 AS=0.2352 PD=1.27714 PS=2.24 NRD=10.5395 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1000 N_X_M1000_d N_A_27_164#_M1000_g N_VPWR_M1001_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.2176 PD=2.8 PS=1.70286 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX4_noxref VNB VPB NWDIODE A=4.278 P=8.32
*
.include "sky130_fd_sc_ms__buf_1.pxi.spice"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlrtp_1 D GATE RESET_B VGND VNB VPB VPWR Q
X0 a_363_74# a_219_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X1 VPWR a_643_74# a_817_48# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X2 a_1045_74# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VPWR a_27_424# a_571_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X4 VPWR a_817_48# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 a_817_48# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X6 a_27_424# D VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X7 a_571_392# a_219_424# a_643_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X8 a_565_74# a_363_74# a_643_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 a_769_74# a_817_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X10 a_643_74# a_363_74# a_762_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X11 VGND GATE a_219_424# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VGND a_27_424# a_565_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 a_643_74# a_219_424# a_769_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X14 a_762_508# a_817_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X15 a_27_424# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X16 a_817_48# a_643_74# a_1045_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 VPWR GATE a_219_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X18 VGND a_817_48# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_363_74# a_219_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

* File: sky130_fd_sc_ms__or2b_2.spice
* Created: Fri Aug 28 18:06:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__or2b_2.pex.spice"
.subckt sky130_fd_sc_ms__or2b_2  VNB VPB B_N A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_B_N_M1002_g N_A_27_368#_M1002_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.107506 AS=0.15675 PD=0.937984 PS=1.67 NRD=17.448 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75002.3 A=0.0825 P=1.4 MULT=1
MM1004 N_X_M1004_d N_A_187_48#_M1004_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.10545 AS=0.144644 PD=1.025 PS=1.26202 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1005 N_X_M1004_d N_A_187_48#_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10545 AS=0.251922 PD=1.025 PS=1.53899 NRD=0.804 NRS=0 M=1 R=4.93333
+ SA=75001 SB=75001.4 A=0.111 P=1.78 MULT=1
MM1003 N_A_187_48#_M1003_d N_A_M1003_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1104 AS=0.217878 PD=0.985 PS=1.33101 NRD=12.18 NRS=0.936 M=1 R=4.26667
+ SA=75001.8 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1007 N_VGND_M1007_d N_A_27_368#_M1007_g N_A_187_48#_M1003_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.2336 AS=0.1104 PD=2.01 PS=0.985 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.3 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1001 N_VPWR_M1001_d N_B_N_M1001_g N_A_27_368#_M1001_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1614 AS=0.2352 PD=1.26429 PS=2.24 NRD=32.1504 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90002.5 A=0.1512 P=2.04 MULT=1
MM1008 N_VPWR_M1001_d N_A_187_48#_M1008_g N_X_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2152 AS=0.2716 PD=1.68571 PS=1.605 NRD=0 NRS=17.5724 M=1 R=6.22222
+ SA=90000.6 SB=90001.8 A=0.2016 P=2.6 MULT=1
MM1009 N_VPWR_M1009_d N_A_187_48#_M1009_g N_X_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.223789 AS=0.2716 PD=1.59547 PS=1.605 NRD=0 NRS=18.4589 M=1 R=6.22222
+ SA=90001.3 SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1006 A_473_368# N_A_M1006_g N_VPWR_M1009_d VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.199811 PD=1.24 PS=1.42453 NRD=12.7853 NRS=23.64 M=1 R=5.55556 SA=90001.9
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1000 N_A_187_48#_M1000_d N_A_27_368#_M1000_g A_473_368# VPB PSHORT L=0.18 W=1
+ AD=0.4 AS=0.12 PD=2.8 PS=1.24 NRD=22.6353 NRS=12.7853 M=1 R=5.55556 SA=90002.3
+ SB=90000.3 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__or2b_2.pxi.spice"
*
.ends
*
*

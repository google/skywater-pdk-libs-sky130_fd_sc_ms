# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__o32ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.765000 1.350000 10.915000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.350000 8.515000 1.780000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.430000 5.635000 1.780000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.430000 4.195000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.430000 1.795000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  2.287500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.595000 0.875000 1.090000 ;
        RECT 0.545000 1.090000 5.975000 1.260000 ;
        RECT 0.645000 1.950000 5.975000 2.120000 ;
        RECT 0.645000 2.120000 0.815000 2.735000 ;
        RECT 1.465000 2.120000 1.795000 2.735000 ;
        RECT 1.555000 0.595000 1.805000 1.090000 ;
        RECT 2.475000 0.595000 2.805000 1.090000 ;
        RECT 3.475000 0.595000 3.805000 1.090000 ;
        RECT 4.735000 2.120000 5.065000 2.735000 ;
        RECT 5.635000 2.120000 5.965000 2.735000 ;
        RECT 5.805000 1.260000 5.975000 1.950000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  3.245000 11.040000 3.415000 ;
      RECT  0.115000  0.255000  4.305000 0.425000 ;
      RECT  0.115000  0.425000  0.365000 1.130000 ;
      RECT  0.115000  1.950000  0.445000 2.905000 ;
      RECT  0.115000  2.905000  2.245000 3.075000 ;
      RECT  1.015000  2.290000  1.265000 2.905000 ;
      RECT  1.045000  0.425000  1.375000 0.920000 ;
      RECT  1.975000  0.425000  2.305000 0.920000 ;
      RECT  1.995000  2.290000  4.055000 2.460000 ;
      RECT  1.995000  2.460000  2.245000 2.905000 ;
      RECT  2.445000  2.630000  2.615000 3.245000 ;
      RECT  2.815000  2.460000  3.145000 2.980000 ;
      RECT  2.975000  0.425000  3.305000 0.920000 ;
      RECT  3.345000  2.630000  3.515000 3.245000 ;
      RECT  3.725000  2.460000  4.055000 2.980000 ;
      RECT  3.975000  0.425000  4.305000 0.750000 ;
      RECT  3.975000  0.750000  6.670000 0.920000 ;
      RECT  4.285000  2.290000  4.535000 2.905000 ;
      RECT  4.285000  2.905000  8.465000 3.075000 ;
      RECT  4.485000  0.085000  4.815000 0.580000 ;
      RECT  4.995000  0.330000  5.325000 0.750000 ;
      RECT  5.265000  2.290000  5.435000 2.905000 ;
      RECT  5.495000  0.085000  5.825000 0.580000 ;
      RECT  5.995000  0.330000  6.670000 0.750000 ;
      RECT  6.145000  1.950000  6.465000 2.905000 ;
      RECT  6.330000  0.920000  6.670000 1.010000 ;
      RECT  6.330000  1.010000 10.670000 1.180000 ;
      RECT  6.635000  1.950000 10.475000 2.120000 ;
      RECT  6.635000  2.120000  6.965000 2.735000 ;
      RECT  6.840000  0.085000  7.170000 0.840000 ;
      RECT  7.135000  2.290000  7.465000 2.905000 ;
      RECT  7.340000  0.350000  7.670000 1.010000 ;
      RECT  7.635000  2.120000  7.965000 2.735000 ;
      RECT  7.840000  0.085000  8.170000 0.840000 ;
      RECT  8.135000  2.290000  8.465000 2.905000 ;
      RECT  8.340000  0.350000  8.670000 1.010000 ;
      RECT  8.695000  2.290000  8.945000 3.245000 ;
      RECT  8.840000  0.085000  9.170000 0.840000 ;
      RECT  9.145000  2.120000  9.475000 2.980000 ;
      RECT  9.340000  0.350000  9.670000 1.010000 ;
      RECT  9.645000  2.290000  9.975000 3.245000 ;
      RECT  9.840000  0.085000 10.170000 0.840000 ;
      RECT 10.145000  2.120000 10.475000 2.980000 ;
      RECT 10.340000  0.350000 10.670000 1.010000 ;
      RECT 10.675000  1.950000 10.925000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
  END
END sky130_fd_sc_ms__o32ai_4

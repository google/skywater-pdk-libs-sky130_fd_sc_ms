* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 a_1013_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=1.06e+12p pd=1.012e+07u as=1.4248e+12p ps=1.338e+07u
M1001 a_137_260# A1 a_1210_74# VNB nlowvt w=640000u l=150000u
+  ad=7.168e+11p pd=7.36e+06u as=5.184e+11p ps=5.46e+06u
M1002 a_137_260# D1 a_549_392# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=7.9e+11p ps=7.58e+06u
M1003 VGND a_137_260# X VNB nlowvt w=740000u l=150000u
+  ad=1.3711e+12p pd=1.359e+07u as=4.144e+11p ps=4.08e+06u
M1004 VGND C1 a_137_260# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_549_392# D1 a_137_260# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_817_392# C1 a_549_392# VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=0p ps=0u
M1007 a_1210_74# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_549_392# C1 a_817_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B1 a_137_260# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_137_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_137_260# D1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_1210_74# A1 a_137_260# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_817_392# B1 a_1013_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_137_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1015 a_1013_392# B1 a_817_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_137_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A1 a_1013_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_137_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1013_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_137_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND D1 a_137_260# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_137_260# C1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR a_137_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 X a_137_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR A2 a_1013_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_137_260# B1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND A2 a_1210_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

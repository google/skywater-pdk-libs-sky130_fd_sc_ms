* File: sky130_fd_sc_ms__nand4bb_1.pxi.spice
* Created: Wed Sep  2 12:14:51 2020
* 
x_PM_SKY130_FD_SC_MS__NAND4BB_1%A_N N_A_N_c_74_n N_A_N_M1010_g N_A_N_M1002_g A_N
+ N_A_N_c_77_n N_A_N_c_78_n PM_SKY130_FD_SC_MS__NAND4BB_1%A_N
x_PM_SKY130_FD_SC_MS__NAND4BB_1%B_N N_B_N_M1006_g N_B_N_M1000_g B_N B_N
+ N_B_N_c_104_n PM_SKY130_FD_SC_MS__NAND4BB_1%B_N
x_PM_SKY130_FD_SC_MS__NAND4BB_1%A_27_398# N_A_27_398#_M1002_s
+ N_A_27_398#_M1010_s N_A_27_398#_M1004_g N_A_27_398#_c_137_n
+ N_A_27_398#_M1009_g N_A_27_398#_c_144_n N_A_27_398#_c_138_n
+ N_A_27_398#_c_139_n N_A_27_398#_c_140_n N_A_27_398#_c_141_n
+ N_A_27_398#_c_142_n PM_SKY130_FD_SC_MS__NAND4BB_1%A_27_398#
x_PM_SKY130_FD_SC_MS__NAND4BB_1%A_229_398# N_A_229_398#_M1000_d
+ N_A_229_398#_M1006_d N_A_229_398#_M1001_g N_A_229_398#_M1008_g
+ N_A_229_398#_c_209_n N_A_229_398#_c_201_n N_A_229_398#_c_202_n
+ N_A_229_398#_c_203_n N_A_229_398#_c_211_n N_A_229_398#_c_204_n
+ N_A_229_398#_c_205_n N_A_229_398#_c_206_n N_A_229_398#_c_207_n
+ PM_SKY130_FD_SC_MS__NAND4BB_1%A_229_398#
x_PM_SKY130_FD_SC_MS__NAND4BB_1%C N_C_M1011_g N_C_M1007_g C C N_C_c_279_n
+ N_C_c_280_n PM_SKY130_FD_SC_MS__NAND4BB_1%C
x_PM_SKY130_FD_SC_MS__NAND4BB_1%D N_D_M1003_g N_D_M1005_g D N_D_c_323_n
+ N_D_c_324_n PM_SKY130_FD_SC_MS__NAND4BB_1%D
x_PM_SKY130_FD_SC_MS__NAND4BB_1%VPWR N_VPWR_M1010_d N_VPWR_M1004_d
+ N_VPWR_M1007_d N_VPWR_c_363_n N_VPWR_c_364_n N_VPWR_c_365_n N_VPWR_c_366_n
+ N_VPWR_c_367_n N_VPWR_c_368_n N_VPWR_c_369_n VPWR N_VPWR_c_370_n
+ N_VPWR_c_371_n N_VPWR_c_362_n N_VPWR_c_373_n
+ PM_SKY130_FD_SC_MS__NAND4BB_1%VPWR
x_PM_SKY130_FD_SC_MS__NAND4BB_1%Y N_Y_M1009_s N_Y_M1004_s N_Y_M1008_d
+ N_Y_M1005_d N_Y_c_420_n N_Y_c_433_n N_Y_c_424_n N_Y_c_454_n N_Y_c_457_n
+ N_Y_c_421_n N_Y_c_422_n N_Y_c_425_n N_Y_c_423_n N_Y_c_427_n N_Y_c_428_n Y
+ N_Y_c_429_n PM_SKY130_FD_SC_MS__NAND4BB_1%Y
x_PM_SKY130_FD_SC_MS__NAND4BB_1%VGND N_VGND_M1002_d N_VGND_M1003_d
+ N_VGND_c_512_n N_VGND_c_513_n N_VGND_c_514_n VGND N_VGND_c_515_n
+ N_VGND_c_516_n N_VGND_c_517_n PM_SKY130_FD_SC_MS__NAND4BB_1%VGND
cc_1 VNB N_A_N_c_74_n 0.00668084f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_2 VNB N_A_N_M1010_g 0.0113864f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.41
cc_3 VNB N_A_N_M1002_g 0.0158898f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.97
cc_4 VNB N_A_N_c_77_n 0.0211239f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=0.42
cc_5 VNB N_A_N_c_78_n 0.0537695f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.42
cc_6 VNB N_B_N_M1000_g 0.0307295f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.97
cc_7 VNB B_N 0.00795483f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_8 VNB N_B_N_c_104_n 0.0181595f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=0.42
cc_9 VNB N_A_27_398#_M1004_g 0.0080765f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.375
cc_10 VNB N_A_27_398#_c_137_n 0.0213945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_398#_c_138_n 0.0145839f $X=-0.19 $Y=-0.245 $X2=0.302 $Y2=0.555
cc_12 VNB N_A_27_398#_c_139_n 0.0221586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_398#_c_140_n 0.017953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_398#_c_141_n 0.00769994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_398#_c_142_n 0.05015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_229_398#_M1008_g 0.00689193f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=0.42
cc_17 VNB N_A_229_398#_c_201_n 0.00835289f $X=-0.19 $Y=-0.245 $X2=0.302 $Y2=0.42
cc_18 VNB N_A_229_398#_c_202_n 0.0023091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_229_398#_c_203_n 0.00272739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_229_398#_c_204_n 0.00733291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_229_398#_c_205_n 0.00896425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_229_398#_c_206_n 0.0327686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_229_398#_c_207_n 0.0184894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_C_M1007_g 0.00654267f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.375
cc_25 VNB C 0.00268364f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.97
cc_26 VNB N_C_c_279_n 0.0326491f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=0.42
cc_27 VNB N_C_c_280_n 0.0193704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_D_M1003_g 0.0274698f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.41
cc_29 VNB N_D_c_323_n 0.027378f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=0.42
cc_30 VNB N_D_c_324_n 0.00476542f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=0.42
cc_31 VNB N_VPWR_c_362_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_420_n 0.0206563f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_421_n 0.0203676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_Y_c_422_n 0.00111978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_Y_c_423_n 0.0230393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_512_n 0.0252046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_513_n 0.0138117f $X=-0.19 $Y=-0.245 $X2=0.315 $Y2=0.42
cc_38 VNB N_VGND_c_514_n 0.0331513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_515_n 0.0738552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_516_n 0.0256348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_517_n 0.264832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VPB N_A_N_M1010_g 0.0367227f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.41
cc_43 VPB N_B_N_M1006_g 0.0306921f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.41
cc_44 VPB B_N 0.00758401f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.47
cc_45 VPB N_B_N_c_104_n 0.0147994f $X=-0.19 $Y=1.66 $X2=0.315 $Y2=0.42
cc_46 VPB N_A_27_398#_M1004_g 0.0313316f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.375
cc_47 VPB N_A_27_398#_c_144_n 0.0386754f $X=-0.19 $Y=1.66 $X2=0.302 $Y2=0.42
cc_48 VPB N_A_27_398#_c_140_n 0.014809f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_229_398#_M1008_g 0.0244775f $X=-0.19 $Y=1.66 $X2=0.315 $Y2=0.42
cc_50 VPB N_A_229_398#_c_209_n 0.0136975f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.42
cc_51 VPB N_A_229_398#_c_203_n 0.00384499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_229_398#_c_211_n 0.0144935f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_C_M1007_g 0.0249762f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.375
cc_54 VPB N_D_M1005_g 0.0274945f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.97
cc_55 VPB N_D_c_323_n 0.00573083f $X=-0.19 $Y=1.66 $X2=0.315 $Y2=0.42
cc_56 VPB N_D_c_324_n 0.00431084f $X=-0.19 $Y=1.66 $X2=0.315 $Y2=0.42
cc_57 VPB N_VPWR_c_363_n 0.0238061f $X=-0.19 $Y=1.66 $X2=0.315 $Y2=0.42
cc_58 VPB N_VPWR_c_364_n 0.00678741f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.42
cc_59 VPB N_VPWR_c_365_n 0.00899828f $X=-0.19 $Y=1.66 $X2=0.302 $Y2=0.555
cc_60 VPB N_VPWR_c_366_n 0.0345306f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_367_n 0.00785853f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_368_n 0.0185368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_369_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_370_n 0.0197293f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_371_n 0.0216364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_362_n 0.0778151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_373_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_Y_c_424_n 0.00275675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_Y_c_425_n 0.0418296f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_Y_c_423_n 0.0129607f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_Y_c_427_n 0.0100055f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_Y_c_428_n 0.00786683f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_Y_c_429_n 0.0108315f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 N_A_N_M1010_g N_B_N_M1006_g 0.0135499f $X=0.505 $Y=2.41 $X2=0 $Y2=0
cc_75 N_A_N_c_78_n N_B_N_M1000_g 0.02321f $X=0.52 $Y=0.42 $X2=0 $Y2=0
cc_76 N_A_N_M1010_g B_N 0.00387379f $X=0.505 $Y=2.41 $X2=0 $Y2=0
cc_77 N_A_N_M1010_g N_B_N_c_104_n 0.0155852f $X=0.505 $Y=2.41 $X2=0 $Y2=0
cc_78 N_A_N_M1010_g N_A_27_398#_c_144_n 0.015087f $X=0.505 $Y=2.41 $X2=0 $Y2=0
cc_79 N_A_N_M1002_g N_A_27_398#_c_138_n 0.0154613f $X=0.52 $Y=0.97 $X2=0 $Y2=0
cc_80 N_A_N_c_77_n N_A_27_398#_c_138_n 2.7753e-19 $X=0.315 $Y=0.42 $X2=0 $Y2=0
cc_81 N_A_N_c_74_n N_A_27_398#_c_139_n 0.00113738f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_82 N_A_N_M1002_g N_A_27_398#_c_139_n 0.00814439f $X=0.52 $Y=0.97 $X2=0 $Y2=0
cc_83 N_A_N_c_77_n N_A_27_398#_c_139_n 0.0263917f $X=0.315 $Y=0.42 $X2=0 $Y2=0
cc_84 N_A_N_c_78_n N_A_27_398#_c_139_n 0.0016705f $X=0.52 $Y=0.42 $X2=0 $Y2=0
cc_85 N_A_N_c_74_n N_A_27_398#_c_140_n 0.0171159f $X=0.505 $Y=1.465 $X2=0 $Y2=0
cc_86 N_A_N_M1002_g N_A_27_398#_c_140_n 0.00257859f $X=0.52 $Y=0.97 $X2=0 $Y2=0
cc_87 N_A_N_M1010_g N_VPWR_c_363_n 0.00460946f $X=0.505 $Y=2.41 $X2=0 $Y2=0
cc_88 N_A_N_M1010_g N_VPWR_c_370_n 0.00560776f $X=0.505 $Y=2.41 $X2=0 $Y2=0
cc_89 N_A_N_M1010_g N_VPWR_c_362_n 0.00606454f $X=0.505 $Y=2.41 $X2=0 $Y2=0
cc_90 N_A_N_c_77_n N_VGND_c_512_n 0.0329753f $X=0.315 $Y=0.42 $X2=0 $Y2=0
cc_91 N_A_N_c_78_n N_VGND_c_512_n 0.0111733f $X=0.52 $Y=0.42 $X2=0 $Y2=0
cc_92 N_A_N_c_77_n N_VGND_c_516_n 0.0233084f $X=0.315 $Y=0.42 $X2=0 $Y2=0
cc_93 N_A_N_c_78_n N_VGND_c_516_n 0.00654921f $X=0.52 $Y=0.42 $X2=0 $Y2=0
cc_94 N_A_N_c_77_n N_VGND_c_517_n 0.0133606f $X=0.315 $Y=0.42 $X2=0 $Y2=0
cc_95 N_A_N_c_78_n N_VGND_c_517_n 0.0041842f $X=0.52 $Y=0.42 $X2=0 $Y2=0
cc_96 B_N N_A_27_398#_M1004_g 0.00625965f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_97 N_B_N_M1000_g N_A_27_398#_c_138_n 0.0161954f $X=1.1 $Y=0.925 $X2=0 $Y2=0
cc_98 B_N N_A_27_398#_c_138_n 0.0543686f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_99 N_B_N_c_104_n N_A_27_398#_c_138_n 0.00427209f $X=1.01 $Y=1.635 $X2=0 $Y2=0
cc_100 N_B_N_M1000_g N_A_27_398#_c_139_n 7.96521e-19 $X=1.1 $Y=0.925 $X2=0 $Y2=0
cc_101 B_N N_A_27_398#_c_140_n 0.0178516f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_102 N_B_N_M1000_g N_A_27_398#_c_141_n 0.00116302f $X=1.1 $Y=0.925 $X2=0 $Y2=0
cc_103 B_N N_A_27_398#_c_141_n 0.00375077f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_104 N_B_N_M1000_g N_A_27_398#_c_142_n 0.00760094f $X=1.1 $Y=0.925 $X2=0 $Y2=0
cc_105 B_N N_A_27_398#_c_142_n 7.37692e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_106 N_B_N_M1006_g N_A_229_398#_c_211_n 0.0148701f $X=1.055 $Y=2.41 $X2=0
+ $Y2=0
cc_107 B_N N_A_229_398#_c_211_n 0.0173094f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_108 N_B_N_c_104_n N_A_229_398#_c_211_n 8.17195e-19 $X=1.01 $Y=1.635 $X2=0
+ $Y2=0
cc_109 N_B_N_M1000_g N_A_229_398#_c_204_n 0.00452024f $X=1.1 $Y=0.925 $X2=0
+ $Y2=0
cc_110 N_B_N_M1006_g N_VPWR_c_363_n 0.0046091f $X=1.055 $Y=2.41 $X2=0 $Y2=0
cc_111 B_N N_VPWR_c_363_n 0.0286067f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_112 N_B_N_c_104_n N_VPWR_c_363_n 0.00230627f $X=1.01 $Y=1.635 $X2=0 $Y2=0
cc_113 N_B_N_M1006_g N_VPWR_c_366_n 0.00560776f $X=1.055 $Y=2.41 $X2=0 $Y2=0
cc_114 N_B_N_M1006_g N_VPWR_c_362_n 0.00606454f $X=1.055 $Y=2.41 $X2=0 $Y2=0
cc_115 N_B_N_M1000_g N_Y_c_420_n 0.00275122f $X=1.1 $Y=0.925 $X2=0 $Y2=0
cc_116 N_B_N_M1006_g N_Y_c_427_n 0.00425204f $X=1.055 $Y=2.41 $X2=0 $Y2=0
cc_117 N_B_N_M1000_g N_VGND_c_512_n 0.00535347f $X=1.1 $Y=0.925 $X2=0 $Y2=0
cc_118 N_B_N_M1000_g N_VGND_c_515_n 0.00387193f $X=1.1 $Y=0.925 $X2=0 $Y2=0
cc_119 N_B_N_M1000_g N_VGND_c_517_n 0.00462577f $X=1.1 $Y=0.925 $X2=0 $Y2=0
cc_120 N_A_27_398#_c_138_n N_A_229_398#_M1000_d 0.00232397f $X=1.685 $Y=1.215
+ $X2=-0.19 $Y2=-0.245
cc_121 N_A_27_398#_M1004_g N_A_229_398#_M1008_g 0.032951f $X=2.065 $Y=2.4 $X2=0
+ $Y2=0
cc_122 N_A_27_398#_M1004_g N_A_229_398#_c_209_n 0.018376f $X=2.065 $Y=2.4 $X2=0
+ $Y2=0
cc_123 N_A_27_398#_c_138_n N_A_229_398#_c_209_n 0.00691896f $X=1.685 $Y=1.215
+ $X2=0 $Y2=0
cc_124 N_A_27_398#_c_141_n N_A_229_398#_c_209_n 0.0111546f $X=1.85 $Y=1.215
+ $X2=0 $Y2=0
cc_125 N_A_27_398#_c_142_n N_A_229_398#_c_209_n 0.00148395f $X=2.1 $Y=1.385
+ $X2=0 $Y2=0
cc_126 N_A_27_398#_c_137_n N_A_229_398#_c_201_n 0.0162635f $X=2.1 $Y=1.22 $X2=0
+ $Y2=0
cc_127 N_A_27_398#_c_141_n N_A_229_398#_c_201_n 0.0246367f $X=1.85 $Y=1.215
+ $X2=0 $Y2=0
cc_128 N_A_27_398#_c_142_n N_A_229_398#_c_201_n 0.00174013f $X=2.1 $Y=1.385
+ $X2=0 $Y2=0
cc_129 N_A_27_398#_c_137_n N_A_229_398#_c_202_n 0.00171321f $X=2.1 $Y=1.22 $X2=0
+ $Y2=0
cc_130 N_A_27_398#_c_141_n N_A_229_398#_c_202_n 0.00713039f $X=1.85 $Y=1.215
+ $X2=0 $Y2=0
cc_131 N_A_27_398#_M1004_g N_A_229_398#_c_203_n 0.00852058f $X=2.065 $Y=2.4
+ $X2=0 $Y2=0
cc_132 N_A_27_398#_M1004_g N_A_229_398#_c_211_n 0.00403553f $X=2.065 $Y=2.4
+ $X2=0 $Y2=0
cc_133 N_A_27_398#_c_138_n N_A_229_398#_c_211_n 0.00419957f $X=1.685 $Y=1.215
+ $X2=0 $Y2=0
cc_134 N_A_27_398#_c_137_n N_A_229_398#_c_204_n 0.00302206f $X=2.1 $Y=1.22 $X2=0
+ $Y2=0
cc_135 N_A_27_398#_c_138_n N_A_229_398#_c_204_n 0.0362968f $X=1.685 $Y=1.215
+ $X2=0 $Y2=0
cc_136 N_A_27_398#_c_141_n N_A_229_398#_c_205_n 0.0272167f $X=1.85 $Y=1.215
+ $X2=0 $Y2=0
cc_137 N_A_27_398#_c_142_n N_A_229_398#_c_205_n 0.00305474f $X=2.1 $Y=1.385
+ $X2=0 $Y2=0
cc_138 N_A_27_398#_c_141_n N_A_229_398#_c_206_n 2.21999e-19 $X=1.85 $Y=1.215
+ $X2=0 $Y2=0
cc_139 N_A_27_398#_c_142_n N_A_229_398#_c_206_n 0.0341467f $X=2.1 $Y=1.385 $X2=0
+ $Y2=0
cc_140 N_A_27_398#_c_137_n N_A_229_398#_c_207_n 0.0341467f $X=2.1 $Y=1.22 $X2=0
+ $Y2=0
cc_141 N_A_27_398#_c_144_n N_VPWR_c_363_n 0.0345631f $X=0.28 $Y=2.135 $X2=0
+ $Y2=0
cc_142 N_A_27_398#_M1004_g N_VPWR_c_364_n 0.00567957f $X=2.065 $Y=2.4 $X2=0
+ $Y2=0
cc_143 N_A_27_398#_M1004_g N_VPWR_c_366_n 0.005209f $X=2.065 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A_27_398#_c_144_n N_VPWR_c_370_n 0.00949319f $X=0.28 $Y=2.135 $X2=0
+ $Y2=0
cc_145 N_A_27_398#_M1004_g N_VPWR_c_362_n 0.00541161f $X=2.065 $Y=2.4 $X2=0
+ $Y2=0
cc_146 N_A_27_398#_c_144_n N_VPWR_c_362_n 0.0110977f $X=0.28 $Y=2.135 $X2=0
+ $Y2=0
cc_147 N_A_27_398#_c_137_n N_Y_c_420_n 0.0104202f $X=2.1 $Y=1.22 $X2=0 $Y2=0
cc_148 N_A_27_398#_M1004_g N_Y_c_433_n 0.0102408f $X=2.065 $Y=2.4 $X2=0 $Y2=0
cc_149 N_A_27_398#_M1004_g N_Y_c_427_n 0.00888366f $X=2.065 $Y=2.4 $X2=0 $Y2=0
cc_150 N_A_27_398#_c_138_n N_VGND_M1002_d 0.00380084f $X=1.685 $Y=1.215
+ $X2=-0.19 $Y2=-0.245
cc_151 N_A_27_398#_c_138_n N_VGND_c_512_n 0.0257093f $X=1.685 $Y=1.215 $X2=0
+ $Y2=0
cc_152 N_A_27_398#_c_137_n N_VGND_c_515_n 0.00291649f $X=2.1 $Y=1.22 $X2=0 $Y2=0
cc_153 N_A_27_398#_c_137_n N_VGND_c_517_n 0.0036383f $X=2.1 $Y=1.22 $X2=0 $Y2=0
cc_154 N_A_27_398#_c_139_n N_VGND_c_517_n 9.95189e-19 $X=0.47 $Y=1.07 $X2=0
+ $Y2=0
cc_155 N_A_229_398#_M1008_g N_C_M1007_g 0.0197143f $X=2.655 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A_229_398#_c_201_n C 0.00438395f $X=2.185 $Y=0.875 $X2=0 $Y2=0
cc_157 N_A_229_398#_c_202_n C 0.00690774f $X=2.27 $Y=1.22 $X2=0 $Y2=0
cc_158 N_A_229_398#_c_205_n C 0.0195437f $X=2.58 $Y=1.385 $X2=0 $Y2=0
cc_159 N_A_229_398#_c_206_n C 4.19484e-19 $X=2.58 $Y=1.385 $X2=0 $Y2=0
cc_160 N_A_229_398#_c_207_n C 0.00159237f $X=2.58 $Y=1.22 $X2=0 $Y2=0
cc_161 N_A_229_398#_c_205_n N_C_c_279_n 0.00120656f $X=2.58 $Y=1.385 $X2=0 $Y2=0
cc_162 N_A_229_398#_c_206_n N_C_c_279_n 0.0176384f $X=2.58 $Y=1.385 $X2=0 $Y2=0
cc_163 N_A_229_398#_c_207_n N_C_c_280_n 0.0275008f $X=2.58 $Y=1.22 $X2=0 $Y2=0
cc_164 N_A_229_398#_c_209_n N_VPWR_M1004_d 0.00325885f $X=2.185 $Y=2.055 $X2=0
+ $Y2=0
cc_165 N_A_229_398#_c_203_n N_VPWR_M1004_d 0.00123078f $X=2.27 $Y=1.97 $X2=0
+ $Y2=0
cc_166 N_A_229_398#_c_211_n N_VPWR_c_363_n 0.0353487f $X=1.28 $Y=2.135 $X2=0
+ $Y2=0
cc_167 N_A_229_398#_M1008_g N_VPWR_c_364_n 0.00885644f $X=2.655 $Y=2.4 $X2=0
+ $Y2=0
cc_168 N_A_229_398#_c_211_n N_VPWR_c_366_n 0.00949319f $X=1.28 $Y=2.135 $X2=0
+ $Y2=0
cc_169 N_A_229_398#_M1008_g N_VPWR_c_368_n 0.00460063f $X=2.655 $Y=2.4 $X2=0
+ $Y2=0
cc_170 N_A_229_398#_M1008_g N_VPWR_c_362_n 0.00463681f $X=2.655 $Y=2.4 $X2=0
+ $Y2=0
cc_171 N_A_229_398#_c_211_n N_VPWR_c_362_n 0.0110977f $X=1.28 $Y=2.135 $X2=0
+ $Y2=0
cc_172 N_A_229_398#_c_201_n N_Y_M1009_s 0.00433781f $X=2.185 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_173 N_A_229_398#_c_209_n N_Y_M1004_s 0.0063345f $X=2.185 $Y=2.055 $X2=0 $Y2=0
cc_174 N_A_229_398#_c_201_n N_Y_c_420_n 0.0380801f $X=2.185 $Y=0.875 $X2=0 $Y2=0
cc_175 N_A_229_398#_c_205_n N_Y_c_420_n 0.00927084f $X=2.58 $Y=1.385 $X2=0 $Y2=0
cc_176 N_A_229_398#_c_206_n N_Y_c_420_n 0.00321424f $X=2.58 $Y=1.385 $X2=0 $Y2=0
cc_177 N_A_229_398#_c_207_n N_Y_c_420_n 0.016417f $X=2.58 $Y=1.22 $X2=0 $Y2=0
cc_178 N_A_229_398#_c_209_n N_Y_c_433_n 0.0215898f $X=2.185 $Y=2.055 $X2=0 $Y2=0
cc_179 N_A_229_398#_M1008_g N_Y_c_424_n 3.04814e-19 $X=2.655 $Y=2.4 $X2=0 $Y2=0
cc_180 N_A_229_398#_M1008_g N_Y_c_427_n 7.61858e-19 $X=2.655 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A_229_398#_c_209_n N_Y_c_427_n 0.0220487f $X=2.185 $Y=2.055 $X2=0 $Y2=0
cc_182 N_A_229_398#_c_211_n N_Y_c_427_n 0.0370727f $X=1.28 $Y=2.135 $X2=0 $Y2=0
cc_183 N_A_229_398#_M1008_g N_Y_c_429_n 0.0240657f $X=2.655 $Y=2.4 $X2=0 $Y2=0
cc_184 N_A_229_398#_c_203_n N_Y_c_429_n 0.00629656f $X=2.27 $Y=1.97 $X2=0 $Y2=0
cc_185 N_A_229_398#_c_205_n N_Y_c_429_n 0.0122115f $X=2.58 $Y=1.385 $X2=0 $Y2=0
cc_186 N_A_229_398#_c_206_n N_Y_c_429_n 9.94418e-19 $X=2.58 $Y=1.385 $X2=0 $Y2=0
cc_187 N_A_229_398#_c_204_n N_VGND_c_512_n 0.0138983f $X=1.49 $Y=0.795 $X2=0
+ $Y2=0
cc_188 N_A_229_398#_c_204_n N_VGND_c_515_n 0.00651976f $X=1.49 $Y=0.795 $X2=0
+ $Y2=0
cc_189 N_A_229_398#_c_207_n N_VGND_c_515_n 0.00291649f $X=2.58 $Y=1.22 $X2=0
+ $Y2=0
cc_190 N_A_229_398#_c_201_n N_VGND_c_517_n 0.00894977f $X=2.185 $Y=0.875 $X2=0
+ $Y2=0
cc_191 N_A_229_398#_c_204_n N_VGND_c_517_n 0.00998901f $X=1.49 $Y=0.795 $X2=0
+ $Y2=0
cc_192 N_A_229_398#_c_207_n N_VGND_c_517_n 0.00360083f $X=2.58 $Y=1.22 $X2=0
+ $Y2=0
cc_193 N_A_229_398#_c_201_n A_435_74# 0.0037689f $X=2.185 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_194 N_A_229_398#_c_202_n A_435_74# 0.00207986f $X=2.27 $Y=1.22 $X2=-0.19
+ $Y2=-0.245
cc_195 C N_D_M1003_g 0.00297693f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_196 N_C_c_279_n N_D_M1003_g 0.0177788f $X=3.15 $Y=1.385 $X2=0 $Y2=0
cc_197 N_C_c_280_n N_D_M1003_g 0.0253098f $X=3.15 $Y=1.22 $X2=0 $Y2=0
cc_198 N_C_M1007_g N_D_M1005_g 0.0217308f $X=3.155 $Y=2.4 $X2=0 $Y2=0
cc_199 N_C_M1007_g N_D_c_323_n 0.00473123f $X=3.155 $Y=2.4 $X2=0 $Y2=0
cc_200 C N_D_c_323_n 2.21387e-19 $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_201 N_C_M1007_g N_D_c_324_n 0.00532322f $X=3.155 $Y=2.4 $X2=0 $Y2=0
cc_202 C N_D_c_324_n 0.0160735f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_203 N_C_c_279_n N_D_c_324_n 0.00123002f $X=3.15 $Y=1.385 $X2=0 $Y2=0
cc_204 N_C_M1007_g N_VPWR_c_364_n 4.26433e-19 $X=3.155 $Y=2.4 $X2=0 $Y2=0
cc_205 N_C_M1007_g N_VPWR_c_365_n 0.00203999f $X=3.155 $Y=2.4 $X2=0 $Y2=0
cc_206 N_C_M1007_g N_VPWR_c_368_n 0.005209f $X=3.155 $Y=2.4 $X2=0 $Y2=0
cc_207 N_C_M1007_g N_VPWR_c_362_n 0.00983143f $X=3.155 $Y=2.4 $X2=0 $Y2=0
cc_208 C N_Y_c_420_n 0.0193446f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_209 N_C_c_279_n N_Y_c_420_n 4.92145e-19 $X=3.15 $Y=1.385 $X2=0 $Y2=0
cc_210 N_C_c_280_n N_Y_c_420_n 0.01594f $X=3.15 $Y=1.22 $X2=0 $Y2=0
cc_211 N_C_M1007_g N_Y_c_424_n 0.00644808f $X=3.155 $Y=2.4 $X2=0 $Y2=0
cc_212 N_C_M1007_g N_Y_c_454_n 0.0152306f $X=3.155 $Y=2.4 $X2=0 $Y2=0
cc_213 C N_Y_c_454_n 0.00740674f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_214 N_C_c_279_n N_Y_c_454_n 2.26227e-19 $X=3.15 $Y=1.385 $X2=0 $Y2=0
cc_215 C N_Y_c_457_n 0.0152478f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_216 N_C_c_280_n N_Y_c_457_n 0.00381676f $X=3.15 $Y=1.22 $X2=0 $Y2=0
cc_217 C N_Y_c_422_n 0.0147075f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_218 N_C_c_280_n N_Y_c_422_n 4.96616e-19 $X=3.15 $Y=1.22 $X2=0 $Y2=0
cc_219 N_C_M1007_g N_Y_c_425_n 5.97851e-19 $X=3.155 $Y=2.4 $X2=0 $Y2=0
cc_220 N_C_M1007_g N_Y_c_429_n 0.010691f $X=3.155 $Y=2.4 $X2=0 $Y2=0
cc_221 C N_Y_c_429_n 0.00666519f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_222 N_C_c_279_n N_Y_c_429_n 5.85476e-19 $X=3.15 $Y=1.385 $X2=0 $Y2=0
cc_223 N_C_c_280_n N_VGND_c_515_n 0.00291649f $X=3.15 $Y=1.22 $X2=0 $Y2=0
cc_224 N_C_c_280_n N_VGND_c_517_n 0.00360678f $X=3.15 $Y=1.22 $X2=0 $Y2=0
cc_225 C A_627_74# 0.00402242f $X=3.035 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_226 N_D_M1005_g N_VPWR_c_365_n 0.00343717f $X=3.705 $Y=2.4 $X2=0 $Y2=0
cc_227 N_D_M1005_g N_VPWR_c_371_n 0.005209f $X=3.705 $Y=2.4 $X2=0 $Y2=0
cc_228 N_D_M1005_g N_VPWR_c_362_n 0.00986644f $X=3.705 $Y=2.4 $X2=0 $Y2=0
cc_229 N_D_M1003_g N_Y_c_420_n 0.00950424f $X=3.63 $Y=0.74 $X2=0 $Y2=0
cc_230 N_D_M1005_g N_Y_c_454_n 0.0134232f $X=3.705 $Y=2.4 $X2=0 $Y2=0
cc_231 N_D_c_323_n N_Y_c_454_n 2.19966e-19 $X=3.72 $Y=1.515 $X2=0 $Y2=0
cc_232 N_D_c_324_n N_Y_c_454_n 0.0192103f $X=3.72 $Y=1.515 $X2=0 $Y2=0
cc_233 N_D_M1003_g N_Y_c_457_n 0.0144061f $X=3.63 $Y=0.74 $X2=0 $Y2=0
cc_234 N_D_M1003_g N_Y_c_421_n 0.00742328f $X=3.63 $Y=0.74 $X2=0 $Y2=0
cc_235 N_D_c_323_n N_Y_c_421_n 0.00125338f $X=3.72 $Y=1.515 $X2=0 $Y2=0
cc_236 N_D_c_324_n N_Y_c_421_n 0.0174298f $X=3.72 $Y=1.515 $X2=0 $Y2=0
cc_237 N_D_M1003_g N_Y_c_422_n 0.0044161f $X=3.63 $Y=0.74 $X2=0 $Y2=0
cc_238 N_D_c_324_n N_Y_c_422_n 0.0144298f $X=3.72 $Y=1.515 $X2=0 $Y2=0
cc_239 N_D_M1005_g N_Y_c_425_n 0.0121146f $X=3.705 $Y=2.4 $X2=0 $Y2=0
cc_240 N_D_M1003_g N_Y_c_423_n 0.00477786f $X=3.63 $Y=0.74 $X2=0 $Y2=0
cc_241 N_D_M1005_g N_Y_c_423_n 0.00546002f $X=3.705 $Y=2.4 $X2=0 $Y2=0
cc_242 N_D_c_323_n N_Y_c_423_n 0.00739878f $X=3.72 $Y=1.515 $X2=0 $Y2=0
cc_243 N_D_c_324_n N_Y_c_423_n 0.0332222f $X=3.72 $Y=1.515 $X2=0 $Y2=0
cc_244 N_D_M1005_g N_Y_c_428_n 8.8334e-19 $X=3.705 $Y=2.4 $X2=0 $Y2=0
cc_245 N_D_c_323_n N_Y_c_428_n 4.052e-19 $X=3.72 $Y=1.515 $X2=0 $Y2=0
cc_246 N_D_c_324_n N_Y_c_428_n 0.00774613f $X=3.72 $Y=1.515 $X2=0 $Y2=0
cc_247 N_D_M1005_g N_Y_c_429_n 0.00127267f $X=3.705 $Y=2.4 $X2=0 $Y2=0
cc_248 N_D_M1003_g N_VGND_c_514_n 0.0143888f $X=3.63 $Y=0.74 $X2=0 $Y2=0
cc_249 N_D_M1003_g N_VGND_c_515_n 0.00348163f $X=3.63 $Y=0.74 $X2=0 $Y2=0
cc_250 N_D_M1003_g N_VGND_c_517_n 0.00547865f $X=3.63 $Y=0.74 $X2=0 $Y2=0
cc_251 N_VPWR_M1004_d N_Y_c_433_n 0.0109184f $X=2.155 $Y=1.84 $X2=0 $Y2=0
cc_252 N_VPWR_c_364_n N_Y_c_433_n 0.0235743f $X=2.385 $Y=2.815 $X2=0 $Y2=0
cc_253 N_VPWR_c_362_n N_Y_c_433_n 0.00587618f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_254 N_VPWR_c_364_n N_Y_c_424_n 0.0136383f $X=2.385 $Y=2.815 $X2=0 $Y2=0
cc_255 N_VPWR_c_368_n N_Y_c_424_n 0.014549f $X=3.265 $Y=3.33 $X2=0 $Y2=0
cc_256 N_VPWR_c_362_n N_Y_c_424_n 0.0119743f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_257 N_VPWR_M1007_d N_Y_c_454_n 0.0102689f $X=3.245 $Y=1.84 $X2=0 $Y2=0
cc_258 N_VPWR_c_365_n N_Y_c_454_n 0.0208278f $X=3.43 $Y=2.455 $X2=0 $Y2=0
cc_259 N_VPWR_c_365_n N_Y_c_425_n 0.0280302f $X=3.43 $Y=2.455 $X2=0 $Y2=0
cc_260 N_VPWR_c_371_n N_Y_c_425_n 0.0203497f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_261 N_VPWR_c_362_n N_Y_c_425_n 0.0167756f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_262 N_VPWR_c_364_n N_Y_c_427_n 0.0132022f $X=2.385 $Y=2.815 $X2=0 $Y2=0
cc_263 N_VPWR_c_366_n N_Y_c_427_n 0.0145333f $X=2.175 $Y=3.33 $X2=0 $Y2=0
cc_264 N_VPWR_c_362_n N_Y_c_427_n 0.0119681f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_265 N_VPWR_c_364_n N_Y_c_429_n 0.00235032f $X=2.385 $Y=2.815 $X2=0 $Y2=0
cc_266 N_VPWR_c_365_n N_Y_c_429_n 0.0272647f $X=3.43 $Y=2.455 $X2=0 $Y2=0
cc_267 N_VPWR_c_362_n N_Y_c_429_n 0.00570155f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_268 N_Y_c_421_n N_VGND_M1003_d 0.00419683f $X=4.055 $Y=1.095 $X2=0 $Y2=0
cc_269 N_Y_c_420_n N_VGND_c_514_n 0.0222791f $X=3.485 $Y=0.485 $X2=0 $Y2=0
cc_270 N_Y_c_457_n N_VGND_c_514_n 0.0162446f $X=3.57 $Y=1.01 $X2=0 $Y2=0
cc_271 N_Y_c_421_n N_VGND_c_514_n 0.0281795f $X=4.055 $Y=1.095 $X2=0 $Y2=0
cc_272 N_Y_c_420_n N_VGND_c_515_n 0.0795465f $X=3.485 $Y=0.485 $X2=0 $Y2=0
cc_273 N_Y_c_420_n N_VGND_c_517_n 0.0668803f $X=3.485 $Y=0.485 $X2=0 $Y2=0
cc_274 N_Y_c_420_n A_435_74# 0.0013155f $X=3.485 $Y=0.485 $X2=-0.19 $Y2=-0.245
cc_275 N_Y_c_420_n A_513_74# 0.0103574f $X=3.485 $Y=0.485 $X2=-0.19 $Y2=-0.245
cc_276 N_Y_c_420_n A_627_74# 0.00894458f $X=3.485 $Y=0.485 $X2=-0.19 $Y2=-0.245
cc_277 N_Y_c_457_n A_627_74# 0.00432805f $X=3.57 $Y=1.01 $X2=-0.19 $Y2=-0.245
cc_278 N_Y_c_422_n A_627_74# 9.34031e-19 $X=3.655 $Y=1.095 $X2=-0.19 $Y2=-0.245

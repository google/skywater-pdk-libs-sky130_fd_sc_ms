* File: sky130_fd_sc_ms__dlrtn_1.pex.spice
* Created: Fri Aug 28 17:27:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLRTN_1%D 3 7 9 12
r29 12 15 40.7387 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.592 $Y=1.615
+ $X2=0.592 $Y2=1.78
r30 12 14 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.592 $Y=1.615
+ $X2=0.592 $Y2=1.45
r31 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.615 $X2=0.6 $Y2=1.615
r32 9 13 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.72 $Y=1.615 $X2=0.6
+ $Y2=1.615
r33 7 15 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=0.51 $Y=2.39 $X2=0.51
+ $Y2=1.78
r34 3 14 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.495 $Y=0.955
+ $X2=0.495 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_1%GATE_N 3 7 9 12
r38 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.615
+ $X2=1.17 $Y2=1.78
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.615
+ $X2=1.17 $Y2=1.45
r40 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.615 $X2=1.17 $Y2=1.615
r41 7 15 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=1.13 $Y=2.39 $X2=1.13
+ $Y2=1.78
r42 3 14 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.085 $Y=0.86
+ $X2=1.085 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_1%A_232_98# 1 2 9 13 17 20 23 25 26 29 31 36
+ 37 39 40 43 44 47 48
c128 29 0 1.46239e-19 $X=3.875 $Y=1.805
r129 55 57 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.875 $Y=2.195
+ $X2=3.89 $Y2=2.195
r130 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.74
+ $Y=1.505 $X2=1.74 $Y2=1.505
r131 47 48 9.42615 $w=4.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.432 $Y=2.115
+ $X2=1.432 $Y2=1.95
r132 44 57 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=4.08 $Y=2.195
+ $X2=3.89 $Y2=2.195
r133 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.08
+ $Y=2.195 $X2=4.08 $Y2=2.195
r134 41 43 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.08 $Y=2.52
+ $X2=4.08 $Y2=2.195
r135 39 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.915 $Y=2.605
+ $X2=4.08 $Y2=2.52
r136 39 40 146.139 $w=1.68e-07 $l=2.24e-06 $layer=LI1_cond $X=3.915 $Y=2.605
+ $X2=1.675 $Y2=2.605
r137 37 51 9.11389 $w=2.71e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.59 $Y=1.67
+ $X2=1.675 $Y2=1.505
r138 37 48 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.59 $Y=1.67
+ $X2=1.59 $Y2=1.95
r139 36 40 9.10402 $w=1.7e-07 $l=2.82319e-07 $layer=LI1_cond $X=1.432 $Y=2.52
+ $X2=1.675 $Y2=2.605
r140 35 47 1.89893 $w=4.83e-07 $l=7.7e-08 $layer=LI1_cond $X=1.432 $Y=2.192
+ $X2=1.432 $Y2=2.115
r141 35 36 8.08894 $w=4.83e-07 $l=3.28e-07 $layer=LI1_cond $X=1.432 $Y=2.192
+ $X2=1.432 $Y2=2.52
r142 31 51 18.9077 $w=2.71e-07 $l=4.2e-07 $layer=LI1_cond $X=1.675 $Y=1.085
+ $X2=1.675 $Y2=1.505
r143 31 33 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.505 $Y=1.085
+ $X2=1.3 $Y2=1.085
r144 27 29 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=3.72 $Y=1.805
+ $X2=3.875 $Y2=1.805
r145 25 52 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=2.065 $Y=1.505
+ $X2=1.74 $Y2=1.505
r146 25 26 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.065 $Y=1.505
+ $X2=2.065 $Y2=1.34
r147 21 57 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.89 $Y=2.36
+ $X2=3.89 $Y2=2.195
r148 21 23 151.597 $w=1.8e-07 $l=3.9e-07 $layer=POLY_cond $X=3.89 $Y=2.36
+ $X2=3.89 $Y2=2.75
r149 20 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.875 $Y=2.03
+ $X2=3.875 $Y2=2.195
r150 19 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.875 $Y=1.88
+ $X2=3.875 $Y2=1.805
r151 19 20 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.875 $Y=1.88
+ $X2=3.875 $Y2=2.03
r152 15 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.72 $Y=1.73
+ $X2=3.72 $Y2=1.805
r153 15 17 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=3.72 $Y=1.73
+ $X2=3.72 $Y2=0.69
r154 11 26 34.7346 $w=1.65e-07 $l=1.6e-07 $layer=POLY_cond $X=2.225 $Y=1.34
+ $X2=2.065 $Y2=1.34
r155 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.225 $Y=1.34
+ $X2=2.225 $Y2=0.78
r156 7 26 34.7346 $w=1.65e-07 $l=3.7229e-07 $layer=POLY_cond $X=2.155 $Y=1.67
+ $X2=2.065 $Y2=1.34
r157 7 9 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=2.155 $Y=1.67
+ $X2=2.155 $Y2=2.38
r158 2 47 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.22
+ $Y=1.97 $X2=1.355 $Y2=2.115
r159 1 33 182 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.49 $X2=1.3 $Y2=1.035
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_1%A_27_136# 1 2 7 9 11 13 15 19 24 25 28 31 33
+ 34
c79 7 0 7.69973e-20 $X=2.775 $Y=1.59
r80 33 34 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.272 $Y=2.115
+ $X2=0.272 $Y2=1.95
r81 31 34 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.18 $Y=1.25 $X2=0.18
+ $Y2=1.95
r82 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.7
+ $Y=1.425 $X2=2.7 $Y2=1.425
r83 26 28 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.7 $Y=0.75 $X2=2.7
+ $Y2=1.425
r84 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.535 $Y=0.665
+ $X2=2.7 $Y2=0.75
r85 24 25 136.353 $w=1.68e-07 $l=2.09e-06 $layer=LI1_cond $X=2.535 $Y=0.665
+ $X2=0.445 $Y2=0.665
r86 17 31 8.81775 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=0.27 $Y=1.075
+ $X2=0.27 $Y2=1.25
r87 17 19 3.95123 $w=3.48e-07 $l=1.2e-07 $layer=LI1_cond $X=0.27 $Y=1.075
+ $X2=0.27 $Y2=0.955
r88 16 25 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=0.27 $Y=0.75
+ $X2=0.445 $Y2=0.665
r89 16 19 6.75002 $w=3.48e-07 $l=2.05e-07 $layer=LI1_cond $X=0.27 $Y=0.75
+ $X2=0.27 $Y2=0.955
r90 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.33 $Y=1.085
+ $X2=3.33 $Y2=0.69
r91 12 29 47.839 $w=2.67e-07 $l=3.37565e-07 $layer=POLY_cond $X=2.865 $Y=1.16
+ $X2=2.7 $Y2=1.425
r92 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.255 $Y=1.16
+ $X2=3.33 $Y2=1.085
r93 11 12 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.255 $Y=1.16
+ $X2=2.865 $Y2=1.16
r94 7 29 34.9261 $w=2.67e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.775 $Y=1.59
+ $X2=2.7 $Y2=1.425
r95 7 9 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=2.775 $Y=1.59
+ $X2=2.775 $Y2=2.46
r96 2 33 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.14
+ $Y=1.97 $X2=0.285 $Y2=2.115
r97 1 19 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.68 $X2=0.28 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_1%A_357_392# 1 2 9 13 16 17 22 23 24 26 27 32
+ 38
c97 32 0 7.69973e-20 $X=2.16 $Y=1.045
c98 26 0 1.0947e-19 $X=4.17 $Y=1.355
c99 17 0 1.46239e-19 $X=3.075 $Y=1.925
r100 37 38 7.70264 $w=5.08e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=2.095
+ $X2=2.245 $Y2=2.095
r101 35 37 5.39408 $w=5.08e-07 $l=2.3e-07 $layer=LI1_cond $X=1.93 $Y=2.095
+ $X2=2.16 $Y2=2.095
r102 30 32 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=2.01 $Y=1.045
+ $X2=2.16 $Y2=1.045
r103 27 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.17 $Y=1.355
+ $X2=4.17 $Y2=1.19
r104 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.17
+ $Y=1.355 $X2=4.17 $Y2=1.355
r105 24 26 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=3.405 $Y=1.355
+ $X2=4.17 $Y2=1.355
r106 23 41 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.24 $Y=1.61
+ $X2=3.24 $Y2=1.775
r107 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.24
+ $Y=1.61 $X2=3.24 $Y2=1.61
r108 20 22 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=3.24 $Y=1.84
+ $X2=3.24 $Y2=1.61
r109 19 24 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=3.24 $Y=1.52
+ $X2=3.405 $Y2=1.355
r110 19 22 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.24 $Y=1.52 $X2=3.24
+ $Y2=1.61
r111 17 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.075 $Y=1.925
+ $X2=3.24 $Y2=1.84
r112 17 38 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.075 $Y=1.925
+ $X2=2.245 $Y2=1.925
r113 16 37 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=2.16 $Y=1.84
+ $X2=2.16 $Y2=2.095
r114 15 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.16 $Y=1.17
+ $X2=2.16 $Y2=1.045
r115 15 16 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.16 $Y=1.17
+ $X2=2.16 $Y2=1.84
r116 13 43 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.195 $Y=0.58
+ $X2=4.195 $Y2=1.19
r117 9 41 266.266 $w=1.8e-07 $l=6.85e-07 $layer=POLY_cond $X=3.195 $Y=2.46
+ $X2=3.195 $Y2=1.775
r118 2 35 600 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=1.785
+ $Y=1.96 $X2=1.93 $Y2=2.145
r119 1 30 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=1.865
+ $Y=0.41 $X2=2.01 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_1%A_897_406# 1 2 9 13 16 19 23 26 27 30 34 40
+ 42 43 44 49 52 53
c122 53 0 1.72324e-19 $X=6.61 $Y=1.485
c123 44 0 4.25141e-20 $X=5.715 $Y=1.72
c124 43 0 1.67582e-19 $X=5.715 $Y=1.805
c125 40 0 1.20795e-19 $X=6.415 $Y=1.805
c126 27 0 1.83245e-19 $X=5.465 $Y=2.195
c127 16 0 1.0947e-19 $X=4.65 $Y=2.03
r128 53 59 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=6.615 $Y=1.485
+ $X2=6.615 $Y2=1.65
r129 53 58 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=6.615 $Y=1.485
+ $X2=6.615 $Y2=1.32
r130 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.61
+ $Y=1.485 $X2=6.61 $Y2=1.485
r131 47 49 3.46863 $w=4.98e-07 $l=1.45e-07 $layer=LI1_cond $X=5.715 $Y=2.195
+ $X2=5.715 $Y2=2.34
r132 46 47 5.02353 $w=4.98e-07 $l=2.1e-07 $layer=LI1_cond $X=5.715 $Y=1.985
+ $X2=5.715 $Y2=2.195
r133 43 46 4.30588 $w=4.98e-07 $l=1.8e-07 $layer=LI1_cond $X=5.715 $Y=1.805
+ $X2=5.715 $Y2=1.985
r134 43 44 7.60339 $w=4.98e-07 $l=8.5e-08 $layer=LI1_cond $X=5.715 $Y=1.805
+ $X2=5.715 $Y2=1.72
r135 42 44 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.55 $Y=1.13
+ $X2=5.55 $Y2=1.72
r136 41 43 7.15667 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=5.965 $Y=1.805
+ $X2=5.715 $Y2=1.805
r137 40 52 13.9429 $w=2.8e-07 $l=4e-07 $layer=LI1_cond $X=6.415 $Y=1.805
+ $X2=6.595 $Y2=1.485
r138 40 41 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=6.415 $Y=1.805
+ $X2=5.965 $Y2=1.805
r139 32 42 9.56083 $w=3.93e-07 $l=1.97e-07 $layer=LI1_cond $X=5.437 $Y=0.933
+ $X2=5.437 $Y2=1.13
r140 32 34 12.1955 $w=3.93e-07 $l=4.18e-07 $layer=LI1_cond $X=5.437 $Y=0.933
+ $X2=5.437 $Y2=0.515
r141 30 56 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.65 $Y=2.195
+ $X2=4.65 $Y2=2.36
r142 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.65
+ $Y=2.195 $X2=4.65 $Y2=2.195
r143 27 47 3.16914 $w=3.3e-07 $l=2.5e-07 $layer=LI1_cond $X=5.465 $Y=2.195
+ $X2=5.715 $Y2=2.195
r144 27 29 28.4618 $w=3.28e-07 $l=8.15e-07 $layer=LI1_cond $X=5.465 $Y=2.195
+ $X2=4.65 $Y2=2.195
r145 25 26 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=4.635 $Y=1.34
+ $X2=4.635 $Y2=1.49
r146 23 59 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=6.695 $Y=2.4
+ $X2=6.695 $Y2=1.65
r147 19 58 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.6 $Y=0.74 $X2=6.6
+ $Y2=1.32
r148 16 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.65 $Y=2.03
+ $X2=4.65 $Y2=2.195
r149 16 26 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=4.65 $Y=2.03
+ $X2=4.65 $Y2=1.49
r150 13 25 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=4.62 $Y=0.58
+ $X2=4.62 $Y2=1.34
r151 9 56 151.597 $w=1.8e-07 $l=3.9e-07 $layer=POLY_cond $X=4.575 $Y=2.75
+ $X2=4.575 $Y2=2.36
r152 2 49 300 $w=1.7e-07 $l=6e-07 $layer=licon1_PDIFF $count=2 $X=5.58 $Y=1.84
+ $X2=5.8 $Y2=2.34
r153 2 46 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=5.58
+ $Y=1.84 $X2=5.8 $Y2=1.985
r154 1 34 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.26
+ $Y=0.37 $X2=5.405 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_1%A_657_392# 1 2 7 8 9 11 12 14 21 26 27 28 31
+ 33 34 36 38 39
c104 9 0 2.88377e-19 $X=5.49 $Y=1.725
c105 8 0 1.70198e-19 $X=5.295 $Y=1.26
c106 7 0 1.83245e-19 $X=5.545 $Y=1.26
r107 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.13
+ $Y=1.465 $X2=5.13 $Y2=1.465
r108 36 38 8.97739 $w=3.02e-07 $l=2.13787e-07 $layer=LI1_cond $X=4.985 $Y=1.3
+ $X2=5.097 $Y2=1.465
r109 35 36 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.985 $Y=1.02
+ $X2=4.985 $Y2=1.3
r110 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.9 $Y=0.935
+ $X2=4.985 $Y2=1.02
r111 33 34 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4.9 $Y=0.935
+ $X2=4.145 $Y2=0.935
r112 29 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.98 $Y=0.85
+ $X2=4.145 $Y2=0.935
r113 29 31 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=3.98 $Y=0.85
+ $X2=3.98 $Y2=0.58
r114 27 38 12.5232 $w=3.02e-07 $l=3.96447e-07 $layer=LI1_cond $X=4.9 $Y=1.775
+ $X2=5.097 $Y2=1.465
r115 27 28 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=4.9 $Y=1.775
+ $X2=3.745 $Y2=1.775
r116 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.66 $Y=1.86
+ $X2=3.745 $Y2=1.775
r117 25 26 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.66 $Y=1.86
+ $X2=3.66 $Y2=2.18
r118 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.575 $Y=2.265
+ $X2=3.66 $Y2=2.18
r119 21 23 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.575 $Y=2.265
+ $X2=3.425 $Y2=2.265
r120 17 39 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=5.13 $Y=1.575
+ $X2=5.13 $Y2=1.465
r121 15 39 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=5.13 $Y=1.335
+ $X2=5.13 $Y2=1.465
r122 12 14 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.62 $Y=1.185
+ $X2=5.62 $Y2=0.74
r123 9 17 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=5.49 $Y=1.65
+ $X2=5.13 $Y2=1.65
r124 9 11 164.683 $w=1.8e-07 $l=6.15e-07 $layer=POLY_cond $X=5.49 $Y=1.725
+ $X2=5.49 $Y2=2.34
r125 8 15 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.295 $Y=1.26
+ $X2=5.13 $Y2=1.335
r126 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.545 $Y=1.26
+ $X2=5.62 $Y2=1.185
r127 7 8 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=5.545 $Y=1.26
+ $X2=5.295 $Y2=1.26
r128 2 23 600 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=1 $X=3.285
+ $Y=1.96 $X2=3.425 $Y2=2.265
r129 1 31 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=3.795
+ $Y=0.37 $X2=3.98 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_1%RESET_B 3 6 8 11 13
c41 13 0 4.25141e-20 $X=6.07 $Y=1.22
r42 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.07 $Y=1.385
+ $X2=6.07 $Y2=1.55
r43 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.07 $Y=1.385
+ $X2=6.07 $Y2=1.22
r44 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.07
+ $Y=1.385 $X2=6.07 $Y2=1.385
r45 8 12 2.96342 $w=3.48e-07 $l=9e-08 $layer=LI1_cond $X=6.06 $Y=1.295 $X2=6.06
+ $Y2=1.385
r46 6 14 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=6.11 $Y=2.34 $X2=6.11
+ $Y2=1.55
r47 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.01 $Y=0.74 $X2=6.01
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_1%VPWR 1 2 3 4 17 21 25 30 31 32 41 48 55 56
+ 59 62 69
r74 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r75 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r76 56 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r77 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r78 53 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.585 $Y=3.33
+ $X2=6.42 $Y2=3.33
r79 53 55 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.585 $Y=3.33
+ $X2=6.96 $Y2=3.33
r80 52 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r81 52 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.04
+ $Y2=3.33
r82 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r83 49 51 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.43 $Y=3.33 $X2=6
+ $Y2=3.33
r84 48 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.255 $Y=3.33
+ $X2=6.42 $Y2=3.33
r85 48 51 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.255 $Y=3.33 $X2=6
+ $Y2=3.33
r86 47 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r87 46 47 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r88 43 46 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.56 $Y2=3.33
r89 43 44 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r90 41 49 10.1669 $w=1.7e-07 $l=3.98e-07 $layer=LI1_cond $X=5.032 $Y=3.33
+ $X2=5.43 $Y2=3.33
r91 41 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r92 41 62 9.55358 $w=7.93e-07 $l=6.35e-07 $layer=LI1_cond $X=5.032 $Y=3.33
+ $X2=5.032 $Y2=2.695
r93 41 46 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.635 $Y=3.33
+ $X2=4.56 $Y2=3.33
r94 40 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r95 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r96 37 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r97 37 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r98 36 39 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r99 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r100 34 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=0.82 $Y2=3.33
r101 34 36 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=1.2 $Y2=3.33
r102 32 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r103 32 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r104 30 39 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.3 $Y=3.33
+ $X2=2.16 $Y2=3.33
r105 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.3 $Y=3.33
+ $X2=2.465 $Y2=3.33
r106 29 43 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=2.63 $Y=3.33
+ $X2=2.64 $Y2=3.33
r107 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.63 $Y=3.33
+ $X2=2.465 $Y2=3.33
r108 25 28 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.42 $Y=2.145
+ $X2=6.42 $Y2=2.825
r109 23 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=3.245
+ $X2=6.42 $Y2=3.33
r110 23 28 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=6.42 $Y=3.245
+ $X2=6.42 $Y2=2.825
r111 19 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=3.245
+ $X2=2.465 $Y2=3.33
r112 19 21 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=2.465 $Y=3.245
+ $X2=2.465 $Y2=2.945
r113 15 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=3.245
+ $X2=0.82 $Y2=3.33
r114 15 17 39.4624 $w=3.28e-07 $l=1.13e-06 $layer=LI1_cond $X=0.82 $Y=3.245
+ $X2=0.82 $Y2=2.115
r115 4 28 600 $w=1.7e-07 $l=1.08946e-06 $layer=licon1_PDIFF $count=1 $X=6.2
+ $Y=1.84 $X2=6.42 $Y2=2.825
r116 4 25 300 $w=1.7e-07 $l=4.00156e-07 $layer=licon1_PDIFF $count=2 $X=6.2
+ $Y=1.84 $X2=6.42 $Y2=2.145
r117 3 62 300 $w=1.7e-07 $l=6.73053e-07 $layer=licon1_PDIFF $count=2 $X=4.665
+ $Y=2.54 $X2=5.265 $Y2=2.695
r118 2 21 600 $w=1.7e-07 $l=1.08946e-06 $layer=licon1_PDIFF $count=1 $X=2.245
+ $Y=1.96 $X2=2.465 $Y2=2.945
r119 1 17 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=0.6
+ $Y=1.97 $X2=0.82 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_1%Q 1 2 9 13 14 15 16 23 32
r22 21 23 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=6.935 $Y=2 $X2=6.935
+ $Y2=2.035
r23 15 16 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=6.935 $Y=2.405
+ $X2=6.935 $Y2=2.775
r24 14 21 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=6.935 $Y=1.975
+ $X2=6.935 $Y2=2
r25 14 32 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=6.935 $Y=1.975
+ $X2=6.935 $Y2=1.82
r26 14 15 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=6.935 $Y=2.06
+ $X2=6.935 $Y2=2.405
r27 14 23 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=6.935 $Y=2.06
+ $X2=6.935 $Y2=2.035
r28 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.03 $Y=1.13 $X2=7.03
+ $Y2=1.82
r29 7 13 9.39714 $w=3.83e-07 $l=1.92e-07 $layer=LI1_cond $X=6.922 $Y=0.938
+ $X2=6.922 $Y2=1.13
r30 7 9 12.6619 $w=3.83e-07 $l=4.23e-07 $layer=LI1_cond $X=6.922 $Y=0.938
+ $X2=6.922 $Y2=0.515
r31 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.785
+ $Y=1.84 $X2=6.92 $Y2=1.985
r32 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.785
+ $Y=1.84 $X2=6.92 $Y2=2.815
r33 1 9 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=6.675
+ $Y=0.37 $X2=6.895 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRTN_1%VGND 1 2 3 4 15 19 22 23 25 26 27 29 53 54
+ 58 66 72
c67 19 0 1.72324e-19 $X=6.305 $Y=0.49
c68 15 0 1.70198e-19 $X=4.84 $Y=0.515
r69 70 72 7.43269 $w=4.93e-07 $l=8e-08 $layer=LI1_cond $X=3.12 $Y=0.162 $X2=3.2
+ $Y2=0.162
r70 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r71 68 70 2.05387 $w=4.93e-07 $l=8.5e-08 $layer=LI1_cond $X=3.035 $Y=0.162
+ $X2=3.12 $Y2=0.162
r72 65 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r73 64 68 9.54446 $w=4.93e-07 $l=3.95e-07 $layer=LI1_cond $X=2.64 $Y=0.162
+ $X2=3.035 $Y2=0.162
r74 64 66 12.3861 $w=4.93e-07 $l=2.85e-07 $layer=LI1_cond $X=2.64 $Y=0.162
+ $X2=2.355 $Y2=0.162
r75 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r76 58 61 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.79 $Y=0 $X2=0.79
+ $Y2=0.325
r77 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r78 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r79 51 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r80 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r81 48 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r82 47 50 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=6 $Y2=0
r83 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r84 45 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r85 44 72 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=3.2
+ $Y2=0
r86 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r87 41 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r88 40 66 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=2.355
+ $Y2=0
r89 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r90 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r91 38 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r92 37 40 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r93 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r94 35 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r95 35 37 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r96 32 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r97 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r98 29 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r99 29 31 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.24
+ $Y2=0
r100 27 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r101 27 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r102 25 50 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.14 $Y=0 $X2=6
+ $Y2=0
r103 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.14 $Y=0 $X2=6.305
+ $Y2=0
r104 24 53 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=6.47 $Y=0 $X2=6.96
+ $Y2=0
r105 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.47 $Y=0 $X2=6.305
+ $Y2=0
r106 22 44 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=4.67 $Y=0 $X2=4.56
+ $Y2=0
r107 22 23 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.67 $Y=0 $X2=4.84
+ $Y2=0
r108 21 47 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=5.01 $Y=0 $X2=5.04
+ $Y2=0
r109 21 23 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.01 $Y=0 $X2=4.84
+ $Y2=0
r110 17 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.305 $Y=0.085
+ $X2=6.305 $Y2=0
r111 17 19 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=6.305 $Y=0.085
+ $X2=6.305 $Y2=0.49
r112 13 23 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.84 $Y=0.085
+ $X2=4.84 $Y2=0
r113 13 15 14.575 $w=3.38e-07 $l=4.3e-07 $layer=LI1_cond $X=4.84 $Y=0.085
+ $X2=4.84 $Y2=0.515
r114 4 19 91 $w=1.7e-07 $l=2.73496e-07 $layer=licon1_NDIFF $count=2 $X=6.085
+ $Y=0.37 $X2=6.305 $Y2=0.49
r115 3 15 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=4.695
+ $Y=0.37 $X2=4.84 $Y2=0.515
r116 2 68 91 $w=1.7e-07 $l=7.76338e-07 $layer=licon1_NDIFF $count=2 $X=2.3
+ $Y=0.41 $X2=3.035 $Y2=0.325
r117 1 61 182 $w=1.7e-07 $l=4.51802e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.68 $X2=0.79 $Y2=0.325
.ends


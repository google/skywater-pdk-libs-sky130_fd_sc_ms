* File: sky130_fd_sc_ms__a32oi_2.pxi.spice
* Created: Fri Aug 28 17:08:47 2020
* 
x_PM_SKY130_FD_SC_MS__A32OI_2%B2 N_B2_M1011_g N_B2_M1000_g N_B2_M1017_g
+ N_B2_M1006_g N_B2_c_107_n B2 N_B2_c_108_n N_B2_c_109_n
+ PM_SKY130_FD_SC_MS__A32OI_2%B2
x_PM_SKY130_FD_SC_MS__A32OI_2%B1 N_B1_c_151_n N_B1_M1007_g N_B1_M1001_g
+ N_B1_c_153_n N_B1_M1010_g N_B1_M1003_g B1 B1 N_B1_c_156_n
+ PM_SKY130_FD_SC_MS__A32OI_2%B1
x_PM_SKY130_FD_SC_MS__A32OI_2%A1 N_A1_M1002_g N_A1_c_208_n N_A1_M1008_g
+ N_A1_c_209_n N_A1_M1018_g N_A1_M1015_g A1 N_A1_c_212_n
+ PM_SKY130_FD_SC_MS__A32OI_2%A1
x_PM_SKY130_FD_SC_MS__A32OI_2%A2 N_A2_M1012_g N_A2_M1004_g N_A2_M1019_g
+ N_A2_M1014_g N_A2_c_266_n N_A2_c_267_n N_A2_c_268_n A2 A2 N_A2_c_269_n
+ PM_SKY130_FD_SC_MS__A32OI_2%A2
x_PM_SKY130_FD_SC_MS__A32OI_2%A3 N_A3_M1013_g N_A3_c_322_n N_A3_M1005_g
+ N_A3_M1016_g N_A3_c_324_n N_A3_M1009_g A3 N_A3_c_326_n
+ PM_SKY130_FD_SC_MS__A32OI_2%A3
x_PM_SKY130_FD_SC_MS__A32OI_2%A_27_368# N_A_27_368#_M1000_s N_A_27_368#_M1006_s
+ N_A_27_368#_M1003_d N_A_27_368#_M1015_s N_A_27_368#_M1019_d
+ N_A_27_368#_M1016_s N_A_27_368#_c_362_n N_A_27_368#_c_363_n
+ N_A_27_368#_c_364_n N_A_27_368#_c_379_n N_A_27_368#_c_365_n
+ N_A_27_368#_c_416_p N_A_27_368#_c_385_n N_A_27_368#_c_366_n
+ N_A_27_368#_c_390_n N_A_27_368#_c_367_n N_A_27_368#_c_368_n
+ N_A_27_368#_c_369_n N_A_27_368#_c_370_n N_A_27_368#_c_371_n
+ N_A_27_368#_c_388_n PM_SKY130_FD_SC_MS__A32OI_2%A_27_368#
x_PM_SKY130_FD_SC_MS__A32OI_2%Y N_Y_M1007_d N_Y_M1008_d N_Y_M1000_d N_Y_M1001_s
+ N_Y_c_450_n N_Y_c_460_n N_Y_c_451_n N_Y_c_467_n N_Y_c_447_n N_Y_c_452_n
+ N_Y_c_523_p N_Y_c_474_n N_Y_c_453_n N_Y_c_489_n N_Y_c_448_n Y N_Y_c_455_n Y
+ PM_SKY130_FD_SC_MS__A32OI_2%Y
x_PM_SKY130_FD_SC_MS__A32OI_2%VPWR N_VPWR_M1002_d N_VPWR_M1004_s N_VPWR_M1013_d
+ N_VPWR_c_528_n N_VPWR_c_529_n N_VPWR_c_530_n N_VPWR_c_531_n N_VPWR_c_532_n
+ VPWR N_VPWR_c_533_n N_VPWR_c_534_n N_VPWR_c_535_n N_VPWR_c_527_n
+ N_VPWR_c_537_n N_VPWR_c_538_n PM_SKY130_FD_SC_MS__A32OI_2%VPWR
x_PM_SKY130_FD_SC_MS__A32OI_2%A_27_74# N_A_27_74#_M1011_d N_A_27_74#_M1017_d
+ N_A_27_74#_M1010_s N_A_27_74#_c_595_n N_A_27_74#_c_596_n N_A_27_74#_c_597_n
+ N_A_27_74#_c_598_n N_A_27_74#_c_599_n N_A_27_74#_c_600_n
+ PM_SKY130_FD_SC_MS__A32OI_2%A_27_74#
x_PM_SKY130_FD_SC_MS__A32OI_2%VGND N_VGND_M1011_s N_VGND_M1005_s N_VGND_M1009_s
+ N_VGND_c_632_n N_VGND_c_633_n N_VGND_c_634_n N_VGND_c_635_n VGND
+ N_VGND_c_636_n N_VGND_c_637_n N_VGND_c_638_n N_VGND_c_639_n N_VGND_c_640_n
+ N_VGND_c_641_n PM_SKY130_FD_SC_MS__A32OI_2%VGND
x_PM_SKY130_FD_SC_MS__A32OI_2%A_507_74# N_A_507_74#_M1008_s N_A_507_74#_M1018_s
+ N_A_507_74#_M1014_d N_A_507_74#_c_699_n N_A_507_74#_c_700_n
+ N_A_507_74#_c_701_n N_A_507_74#_c_702_n N_A_507_74#_c_703_n
+ N_A_507_74#_c_704_n PM_SKY130_FD_SC_MS__A32OI_2%A_507_74#
x_PM_SKY130_FD_SC_MS__A32OI_2%A_771_74# N_A_771_74#_M1012_s N_A_771_74#_M1005_d
+ N_A_771_74#_c_766_n N_A_771_74#_c_743_n N_A_771_74#_c_744_n
+ N_A_771_74#_c_745_n PM_SKY130_FD_SC_MS__A32OI_2%A_771_74#
cc_1 VNB N_B2_M1011_g 0.0296069f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_B2_M1000_g 0.00173149f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_3 VNB N_B2_M1017_g 0.0221212f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.74
cc_4 VNB N_B2_M1006_g 0.00170288f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_5 VNB N_B2_c_107_n 0.00135493f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_6 VNB N_B2_c_108_n 0.0480139f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.465
cc_7 VNB N_B2_c_109_n 0.0184277f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=1.54
cc_8 VNB N_B1_c_151_n 0.0164156f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_9 VNB N_B1_M1001_g 0.00641195f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_10 VNB N_B1_c_153_n 0.0207512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B1_M1003_g 0.00642584f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.63
cc_12 VNB B1 0.00940302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B1_c_156_n 0.0571794f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_14 VNB N_A1_M1002_g 0.00752125f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_15 VNB N_A1_c_208_n 0.0205288f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.63
cc_16 VNB N_A1_c_209_n 0.0164898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_M1015_g 0.00714313f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.63
cc_18 VNB A1 0.00441958f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_19 VNB N_A1_c_212_n 0.0762351f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_20 VNB N_A2_M1012_g 0.0249505f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_21 VNB N_A2_M1014_g 0.0289552f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_22 VNB N_A2_c_266_n 0.00990425f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_23 VNB N_A2_c_267_n 0.0162689f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_24 VNB N_A2_c_268_n 0.0139879f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_25 VNB N_A2_c_269_n 0.00476662f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_26 VNB N_A3_M1013_g 0.00707227f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_27 VNB N_A3_c_322_n 0.0192891f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.63
cc_28 VNB N_A3_M1016_g 0.00959774f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.74
cc_29 VNB N_A3_c_324_n 0.0209684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB A3 0.0140818f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_31 VNB N_A3_c_326_n 0.111366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_447_n 0.0117593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_448_n 0.00184708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB Y 0.00206864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VPWR_c_527_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_27_74#_c_595_n 0.0247745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_74#_c_596_n 0.00666543f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_38 VNB N_A_27_74#_c_597_n 0.00978809f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_39 VNB N_A_27_74#_c_598_n 0.00302115f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_40 VNB N_A_27_74#_c_599_n 0.00217191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_74#_c_600_n 0.00716337f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_42 VNB N_VGND_c_632_n 0.00615265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_633_n 0.0123645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_634_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_45 VNB N_VGND_c_635_n 0.0341338f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_46 VNB N_VGND_c_636_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_47 VNB N_VGND_c_637_n 0.0965919f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.465
cc_48 VNB N_VGND_c_638_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_639_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_640_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_641_n 0.353339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_507_74#_c_699_n 0.00199363f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.74
cc_53 VNB N_A_507_74#_c_700_n 0.00487422f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_54 VNB N_A_507_74#_c_701_n 0.00713963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_507_74#_c_702_n 0.00384069f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_56 VNB N_A_507_74#_c_703_n 0.00655402f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_57 VNB N_A_507_74#_c_704_n 0.0022203f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.465
cc_58 VNB N_A_771_74#_c_743_n 0.0275552f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=0.74
cc_59 VNB N_A_771_74#_c_744_n 0.00341417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_771_74#_c_745_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_61 VPB N_B2_M1000_g 0.0267736f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_62 VPB N_B2_M1006_g 0.0226216f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_63 VPB N_B2_c_109_n 0.00802605f $X=-0.19 $Y=1.66 $X2=0.355 $Y2=1.54
cc_64 VPB N_B1_M1001_g 0.0226555f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_65 VPB N_B1_M1003_g 0.0219049f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.63
cc_66 VPB N_A1_M1002_g 0.0249875f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_67 VPB N_A1_M1015_g 0.0256655f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.63
cc_68 VPB N_A2_M1004_g 0.0215337f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_69 VPB N_A2_M1019_g 0.0232282f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=0.74
cc_70 VPB N_A2_c_266_n 6.39815e-19 $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.465
cc_71 VPB N_A2_c_267_n 0.00513808f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.465
cc_72 VPB N_A2_c_268_n 9.02447e-19 $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.465
cc_73 VPB N_A2_c_269_n 0.00613664f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.465
cc_74 VPB N_A3_M1013_g 0.0247016f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_75 VPB N_A3_M1016_g 0.029935f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=0.74
cc_76 VPB N_A_27_368#_c_362_n 0.0366851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_27_368#_c_363_n 0.00237811f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_27_368#_c_364_n 0.00971634f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.465
cc_79 VPB N_A_27_368#_c_365_n 0.00565218f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.54
cc_80 VPB N_A_27_368#_c_366_n 0.00233694f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_27_368#_c_367_n 0.00611944f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_27_368#_c_368_n 0.00392211f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_27_368#_c_369_n 0.0147997f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_27_368#_c_370_n 0.0439896f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_27_368#_c_371_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_Y_c_450_n 0.00292147f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.63
cc_87 VPB N_Y_c_451_n 0.00613428f $X=-0.19 $Y=1.66 $X2=0.355 $Y2=1.465
cc_88 VPB N_Y_c_452_n 0.0107069f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.465
cc_89 VPB N_Y_c_453_n 0.00321801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB Y 0.00110955f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_Y_c_455_n 0.00194701f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_528_n 0.00652507f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_529_n 0.00573348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_530_n 0.00969617f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.465
cc_95 VPB N_VPWR_c_531_n 0.021538f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_532_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.465
cc_97 VPB N_VPWR_c_533_n 0.0616651f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.465
cc_98 VPB N_VPWR_c_534_n 0.0174563f $X=-0.19 $Y=1.66 $X2=0.355 $Y2=1.54
cc_99 VPB N_VPWR_c_535_n 0.027107f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_527_n 0.0794224f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_537_n 0.0132517f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_538_n 0.00641592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 N_B2_M1017_g N_B1_c_151_n 0.0167802f $X=0.975 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_104 N_B2_M1006_g N_B1_M1001_g 0.019567f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_105 N_B2_M1017_g B1 3.50863e-19 $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_106 N_B2_c_107_n B1 0.0101592f $X=0.925 $Y=1.465 $X2=0 $Y2=0
cc_107 N_B2_c_108_n B1 9.46057e-19 $X=1.005 $Y=1.465 $X2=0 $Y2=0
cc_108 N_B2_c_107_n N_B1_c_156_n 0.00166231f $X=0.925 $Y=1.465 $X2=0 $Y2=0
cc_109 N_B2_c_108_n N_B1_c_156_n 0.0238956f $X=1.005 $Y=1.465 $X2=0 $Y2=0
cc_110 N_B2_M1000_g N_A_27_368#_c_362_n 0.0124992f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_111 N_B2_M1006_g N_A_27_368#_c_362_n 2.81906e-19 $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_112 N_B2_c_107_n N_A_27_368#_c_362_n 0.00307517f $X=0.925 $Y=1.465 $X2=0
+ $Y2=0
cc_113 N_B2_c_109_n N_A_27_368#_c_362_n 0.0205168f $X=0.355 $Y=1.54 $X2=0 $Y2=0
cc_114 N_B2_M1000_g N_A_27_368#_c_363_n 0.012228f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_115 N_B2_M1006_g N_A_27_368#_c_363_n 0.0144568f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_116 N_B2_M1000_g N_A_27_368#_c_364_n 0.00282152f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_117 N_B2_M1000_g N_Y_c_450_n 0.00132973f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_118 N_B2_M1006_g N_Y_c_450_n 0.00133968f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_119 N_B2_c_107_n N_Y_c_450_n 0.027698f $X=0.925 $Y=1.465 $X2=0 $Y2=0
cc_120 N_B2_c_108_n N_Y_c_450_n 0.00320408f $X=1.005 $Y=1.465 $X2=0 $Y2=0
cc_121 N_B2_M1006_g N_Y_c_460_n 0.0106396f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_122 N_B2_M1006_g N_Y_c_451_n 0.0132394f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_123 N_B2_c_107_n N_Y_c_451_n 0.0103209f $X=0.925 $Y=1.465 $X2=0 $Y2=0
cc_124 N_B2_M1000_g N_VPWR_c_533_n 0.00333901f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_125 N_B2_M1006_g N_VPWR_c_533_n 0.00333926f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_126 N_B2_M1000_g N_VPWR_c_527_n 0.00426886f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_127 N_B2_M1006_g N_VPWR_c_527_n 0.00423695f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_128 N_B2_M1011_g N_A_27_74#_c_595_n 0.00159319f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_129 N_B2_M1011_g N_A_27_74#_c_596_n 0.0128698f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_130 N_B2_M1017_g N_A_27_74#_c_596_n 0.0134606f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_131 N_B2_c_107_n N_A_27_74#_c_596_n 0.0535577f $X=0.925 $Y=1.465 $X2=0 $Y2=0
cc_132 N_B2_c_108_n N_A_27_74#_c_596_n 0.00469212f $X=1.005 $Y=1.465 $X2=0 $Y2=0
cc_133 N_B2_c_109_n N_A_27_74#_c_597_n 0.0217492f $X=0.355 $Y=1.54 $X2=0 $Y2=0
cc_134 N_B2_M1017_g N_A_27_74#_c_599_n 0.00106427f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_135 N_B2_M1011_g N_VGND_c_632_n 0.0125039f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_136 N_B2_M1017_g N_VGND_c_632_n 0.00182553f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_137 N_B2_M1011_g N_VGND_c_636_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_138 N_B2_M1017_g N_VGND_c_637_n 0.00461464f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_139 N_B2_M1011_g N_VGND_c_641_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_140 N_B2_M1017_g N_VGND_c_641_n 0.00908237f $X=0.975 $Y=0.74 $X2=0 $Y2=0
cc_141 N_B1_M1003_g N_A1_M1002_g 0.0212603f $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_142 B1 A1 0.0311944f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_143 N_B1_c_156_n A1 3.24246e-19 $X=2.005 $Y=1.385 $X2=0 $Y2=0
cc_144 B1 N_A1_c_212_n 0.00251916f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_145 N_B1_c_156_n N_A1_c_212_n 0.0184231f $X=2.005 $Y=1.385 $X2=0 $Y2=0
cc_146 N_B1_M1001_g N_A_27_368#_c_379_n 0.0124108f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_147 N_B1_M1003_g N_A_27_368#_c_379_n 2.72638e-19 $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_148 N_B1_M1001_g N_A_27_368#_c_365_n 0.0119307f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_149 N_B1_M1003_g N_A_27_368#_c_365_n 0.0142975f $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_150 N_B1_M1001_g N_A_27_368#_c_371_n 0.00211007f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_151 N_B1_M1001_g N_Y_c_460_n 5.83856e-19 $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_152 N_B1_M1001_g N_Y_c_451_n 0.018058f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_153 B1 N_Y_c_451_n 0.00587472f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_154 N_B1_c_156_n N_Y_c_451_n 0.00268119f $X=2.005 $Y=1.385 $X2=0 $Y2=0
cc_155 N_B1_M1003_g N_Y_c_467_n 0.00974982f $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_156 N_B1_c_153_n N_Y_c_447_n 0.0114763f $X=1.835 $Y=1.22 $X2=0 $Y2=0
cc_157 B1 N_Y_c_447_n 0.03567f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_158 N_B1_c_156_n N_Y_c_447_n 0.00154259f $X=2.005 $Y=1.385 $X2=0 $Y2=0
cc_159 N_B1_M1003_g N_Y_c_452_n 0.0131783f $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_160 B1 N_Y_c_452_n 0.0248442f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_161 N_B1_c_156_n N_Y_c_452_n 0.00179364f $X=2.005 $Y=1.385 $X2=0 $Y2=0
cc_162 N_B1_c_151_n N_Y_c_474_n 0.00608134f $X=1.405 $Y=1.22 $X2=0 $Y2=0
cc_163 N_B1_c_153_n N_Y_c_474_n 0.0100827f $X=1.835 $Y=1.22 $X2=0 $Y2=0
cc_164 B1 N_Y_c_474_n 0.01963f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_165 N_B1_c_156_n N_Y_c_474_n 6.70031e-19 $X=2.005 $Y=1.385 $X2=0 $Y2=0
cc_166 N_B1_M1001_g N_Y_c_453_n 0.00270544f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_167 N_B1_M1003_g N_Y_c_453_n 0.00404913f $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_168 B1 N_Y_c_453_n 0.0279177f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_169 N_B1_c_156_n N_Y_c_453_n 0.00381358f $X=2.005 $Y=1.385 $X2=0 $Y2=0
cc_170 N_B1_M1001_g N_VPWR_c_533_n 0.00333896f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_171 N_B1_M1003_g N_VPWR_c_533_n 0.00333926f $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_172 N_B1_M1001_g N_VPWR_c_527_n 0.0042374f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_173 N_B1_M1003_g N_VPWR_c_527_n 0.00423742f $X=2.005 $Y=2.4 $X2=0 $Y2=0
cc_174 N_B1_c_151_n N_A_27_74#_c_596_n 6.05444e-19 $X=1.405 $Y=1.22 $X2=0 $Y2=0
cc_175 N_B1_c_151_n N_A_27_74#_c_598_n 0.0119575f $X=1.405 $Y=1.22 $X2=0 $Y2=0
cc_176 N_B1_c_153_n N_A_27_74#_c_598_n 0.0107047f $X=1.835 $Y=1.22 $X2=0 $Y2=0
cc_177 N_B1_c_153_n N_A_27_74#_c_600_n 0.00165289f $X=1.835 $Y=1.22 $X2=0 $Y2=0
cc_178 N_B1_c_151_n N_VGND_c_637_n 0.00278271f $X=1.405 $Y=1.22 $X2=0 $Y2=0
cc_179 N_B1_c_153_n N_VGND_c_637_n 0.00278271f $X=1.835 $Y=1.22 $X2=0 $Y2=0
cc_180 N_B1_c_151_n N_VGND_c_641_n 0.00353526f $X=1.405 $Y=1.22 $X2=0 $Y2=0
cc_181 N_B1_c_153_n N_VGND_c_641_n 0.00357518f $X=1.835 $Y=1.22 $X2=0 $Y2=0
cc_182 N_A1_c_209_n N_A2_M1012_g 0.0117174f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_183 N_A1_c_212_n N_A2_M1012_g 0.0196099f $X=3.345 $Y=1.385 $X2=0 $Y2=0
cc_184 N_A1_M1015_g N_A2_c_266_n 0.0196099f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_185 N_A1_c_212_n N_A2_c_269_n 0.00452181f $X=3.345 $Y=1.385 $X2=0 $Y2=0
cc_186 N_A1_M1002_g N_A_27_368#_c_365_n 0.00109676f $X=2.505 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A1_M1002_g N_A_27_368#_c_385_n 0.0159392f $X=2.505 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A1_M1015_g N_A_27_368#_c_385_n 0.0188795f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_189 N_A1_c_212_n N_A_27_368#_c_385_n 8.27888e-19 $X=3.345 $Y=1.385 $X2=0
+ $Y2=0
cc_190 N_A1_M1015_g N_A_27_368#_c_388_n 0.00849992f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_191 N_A1_c_208_n N_Y_c_447_n 0.0162888f $X=2.895 $Y=1.22 $X2=0 $Y2=0
cc_192 A1 N_Y_c_447_n 0.0256443f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_193 N_A1_c_212_n N_Y_c_447_n 0.00325816f $X=3.345 $Y=1.385 $X2=0 $Y2=0
cc_194 N_A1_M1002_g N_Y_c_452_n 0.0141827f $X=2.505 $Y=2.4 $X2=0 $Y2=0
cc_195 A1 N_Y_c_452_n 0.0244344f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_196 N_A1_c_212_n N_Y_c_452_n 0.0100168f $X=3.345 $Y=1.385 $X2=0 $Y2=0
cc_197 N_A1_M1002_g N_Y_c_453_n 3.25485e-19 $X=2.505 $Y=2.4 $X2=0 $Y2=0
cc_198 N_A1_c_212_n N_Y_c_489_n 0.0077643f $X=3.345 $Y=1.385 $X2=0 $Y2=0
cc_199 N_A1_c_208_n N_Y_c_448_n 0.00251469f $X=2.895 $Y=1.22 $X2=0 $Y2=0
cc_200 N_A1_c_209_n N_Y_c_448_n 0.00224552f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_201 A1 N_Y_c_448_n 0.0214567f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_202 N_A1_c_212_n N_Y_c_448_n 0.00306807f $X=3.345 $Y=1.385 $X2=0 $Y2=0
cc_203 N_A1_M1002_g Y 0.00323021f $X=2.505 $Y=2.4 $X2=0 $Y2=0
cc_204 N_A1_M1015_g Y 0.00236283f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_205 N_A1_c_212_n Y 0.0131017f $X=3.345 $Y=1.385 $X2=0 $Y2=0
cc_206 N_A1_M1015_g N_Y_c_455_n 0.00366775f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_207 N_A1_M1002_g N_VPWR_c_528_n 0.0111752f $X=2.505 $Y=2.4 $X2=0 $Y2=0
cc_208 N_A1_M1015_g N_VPWR_c_528_n 0.0119253f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_209 N_A1_M1002_g N_VPWR_c_533_n 0.00475445f $X=2.505 $Y=2.4 $X2=0 $Y2=0
cc_210 N_A1_M1015_g N_VPWR_c_534_n 0.00475445f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_211 N_A1_M1002_g N_VPWR_c_527_n 0.00939227f $X=2.505 $Y=2.4 $X2=0 $Y2=0
cc_212 N_A1_M1015_g N_VPWR_c_527_n 0.00938771f $X=3.345 $Y=2.4 $X2=0 $Y2=0
cc_213 N_A1_c_208_n N_A_27_74#_c_600_n 9.7204e-19 $X=2.895 $Y=1.22 $X2=0 $Y2=0
cc_214 N_A1_c_208_n N_VGND_c_637_n 0.00279469f $X=2.895 $Y=1.22 $X2=0 $Y2=0
cc_215 N_A1_c_209_n N_VGND_c_637_n 0.00278247f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_216 N_A1_c_208_n N_VGND_c_641_n 0.00357517f $X=2.895 $Y=1.22 $X2=0 $Y2=0
cc_217 N_A1_c_209_n N_VGND_c_641_n 0.00353752f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_218 N_A1_c_208_n N_A_507_74#_c_699_n 0.0079299f $X=2.895 $Y=1.22 $X2=0 $Y2=0
cc_219 N_A1_c_209_n N_A_507_74#_c_699_n 0.0100711f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_220 N_A1_c_208_n N_A_507_74#_c_700_n 6.12241e-19 $X=2.895 $Y=1.22 $X2=0 $Y2=0
cc_221 N_A1_c_209_n N_A_507_74#_c_700_n 0.010463f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_222 N_A1_c_212_n N_A_507_74#_c_700_n 0.00184747f $X=3.345 $Y=1.385 $X2=0
+ $Y2=0
cc_223 N_A1_c_208_n N_A_507_74#_c_703_n 0.00735466f $X=2.895 $Y=1.22 $X2=0 $Y2=0
cc_224 N_A1_c_209_n N_A_507_74#_c_703_n 5.3819e-19 $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_225 N_A1_c_209_n N_A_507_74#_c_704_n 0.00194567f $X=3.325 $Y=1.22 $X2=0 $Y2=0
cc_226 N_A2_c_268_n N_A3_M1013_g 0.0180084f $X=4.31 $Y=1.515 $X2=0 $Y2=0
cc_227 N_A2_M1014_g N_A3_c_326_n 0.0180084f $X=4.325 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A2_c_269_n N_A3_c_326_n 0.0022179f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_229 N_A2_M1004_g N_A_27_368#_c_366_n 0.00942379f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_230 N_A2_M1004_g N_A_27_368#_c_390_n 0.0138797f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_231 N_A2_M1019_g N_A_27_368#_c_390_n 0.0182336f $X=4.31 $Y=2.4 $X2=0 $Y2=0
cc_232 N_A2_c_267_n N_A_27_368#_c_390_n 8.4521e-19 $X=4.22 $Y=1.515 $X2=0 $Y2=0
cc_233 N_A2_c_269_n N_A_27_368#_c_390_n 0.0447968f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_234 N_A2_M1019_g N_A_27_368#_c_367_n 0.00545254f $X=4.31 $Y=2.4 $X2=0 $Y2=0
cc_235 N_A2_c_269_n N_A_27_368#_c_367_n 0.00525994f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_236 N_A2_M1019_g N_A_27_368#_c_368_n 9.79037e-19 $X=4.31 $Y=2.4 $X2=0 $Y2=0
cc_237 N_A2_M1004_g N_A_27_368#_c_388_n 0.00359078f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_238 N_A2_M1019_g N_A_27_368#_c_388_n 6.12264e-19 $X=4.31 $Y=2.4 $X2=0 $Y2=0
cc_239 N_A2_c_269_n N_A_27_368#_c_388_n 0.018893f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_240 N_A2_M1012_g N_Y_c_489_n 4.94418e-19 $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_241 N_A2_c_269_n Y 0.0234231f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_242 N_A2_c_269_n N_Y_c_455_n 0.00420638f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_243 N_A2_M1004_g N_VPWR_c_528_n 4.86935e-19 $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_244 N_A2_M1004_g N_VPWR_c_529_n 0.00220607f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_245 N_A2_M1019_g N_VPWR_c_529_n 0.0134365f $X=4.31 $Y=2.4 $X2=0 $Y2=0
cc_246 N_A2_M1019_g N_VPWR_c_531_n 0.00460063f $X=4.31 $Y=2.4 $X2=0 $Y2=0
cc_247 N_A2_M1004_g N_VPWR_c_534_n 0.005209f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_248 N_A2_M1004_g N_VPWR_c_527_n 0.0098233f $X=3.795 $Y=2.4 $X2=0 $Y2=0
cc_249 N_A2_M1019_g N_VPWR_c_527_n 0.00910094f $X=4.31 $Y=2.4 $X2=0 $Y2=0
cc_250 N_A2_M1014_g N_VGND_c_633_n 0.00177115f $X=4.325 $Y=0.74 $X2=0 $Y2=0
cc_251 N_A2_M1012_g N_VGND_c_637_n 0.00278271f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A2_M1014_g N_VGND_c_637_n 0.00278247f $X=4.325 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A2_M1012_g N_VGND_c_641_n 0.00354791f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A2_M1014_g N_VGND_c_641_n 0.00359462f $X=4.325 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A2_M1012_g N_A_507_74#_c_700_n 4.70861e-19 $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A2_c_269_n N_A_507_74#_c_700_n 0.0164713f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_257 N_A2_M1012_g N_A_507_74#_c_701_n 0.0123067f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_258 N_A2_M1014_g N_A_507_74#_c_701_n 0.0124893f $X=4.325 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A2_M1012_g N_A_507_74#_c_702_n 5.11757e-19 $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A2_M1014_g N_A_507_74#_c_702_n 0.00736432f $X=4.325 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A2_M1012_g N_A_507_74#_c_704_n 0.00142735f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A2_M1014_g N_A_771_74#_c_743_n 0.015265f $X=4.325 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A2_c_269_n N_A_771_74#_c_743_n 0.0124962f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_264 N_A2_M1012_g N_A_771_74#_c_744_n 0.00177175f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_265 N_A2_c_267_n N_A_771_74#_c_744_n 0.00521491f $X=4.22 $Y=1.515 $X2=0 $Y2=0
cc_266 N_A2_c_269_n N_A_771_74#_c_744_n 0.0279649f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_267 N_A3_M1013_g N_A_27_368#_c_367_n 0.00710408f $X=4.935 $Y=2.4 $X2=0 $Y2=0
cc_268 N_A3_M1016_g N_A_27_368#_c_367_n 2.99728e-19 $X=5.485 $Y=2.4 $X2=0 $Y2=0
cc_269 N_A3_M1013_g N_A_27_368#_c_368_n 0.0223921f $X=4.935 $Y=2.4 $X2=0 $Y2=0
cc_270 N_A3_M1013_g N_A_27_368#_c_369_n 0.0149409f $X=4.935 $Y=2.4 $X2=0 $Y2=0
cc_271 N_A3_M1016_g N_A_27_368#_c_369_n 0.0187109f $X=5.485 $Y=2.4 $X2=0 $Y2=0
cc_272 A3 N_A_27_368#_c_369_n 0.00760155f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_273 N_A3_c_326_n N_A_27_368#_c_369_n 0.0155008f $X=5.95 $Y=1.385 $X2=0 $Y2=0
cc_274 N_A3_M1013_g N_A_27_368#_c_370_n 4.81831e-19 $X=4.935 $Y=2.4 $X2=0 $Y2=0
cc_275 N_A3_M1016_g N_A_27_368#_c_370_n 0.0156993f $X=5.485 $Y=2.4 $X2=0 $Y2=0
cc_276 N_A3_M1013_g N_VPWR_c_529_n 9.14446e-19 $X=4.935 $Y=2.4 $X2=0 $Y2=0
cc_277 N_A3_M1013_g N_VPWR_c_530_n 0.00343717f $X=4.935 $Y=2.4 $X2=0 $Y2=0
cc_278 N_A3_M1016_g N_VPWR_c_530_n 0.00343717f $X=5.485 $Y=2.4 $X2=0 $Y2=0
cc_279 N_A3_M1013_g N_VPWR_c_531_n 0.005209f $X=4.935 $Y=2.4 $X2=0 $Y2=0
cc_280 N_A3_M1016_g N_VPWR_c_535_n 0.005209f $X=5.485 $Y=2.4 $X2=0 $Y2=0
cc_281 N_A3_M1013_g N_VPWR_c_527_n 0.00984066f $X=4.935 $Y=2.4 $X2=0 $Y2=0
cc_282 N_A3_M1016_g N_VPWR_c_527_n 0.00986878f $X=5.485 $Y=2.4 $X2=0 $Y2=0
cc_283 N_A3_c_322_n N_VGND_c_633_n 0.00562548f $X=5.315 $Y=1.22 $X2=0 $Y2=0
cc_284 N_A3_c_322_n N_VGND_c_635_n 5.69925e-19 $X=5.315 $Y=1.22 $X2=0 $Y2=0
cc_285 N_A3_c_324_n N_VGND_c_635_n 0.0122959f $X=5.745 $Y=1.22 $X2=0 $Y2=0
cc_286 A3 N_VGND_c_635_n 0.0251682f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_287 N_A3_c_326_n N_VGND_c_635_n 0.00192797f $X=5.95 $Y=1.385 $X2=0 $Y2=0
cc_288 N_A3_c_322_n N_VGND_c_638_n 0.00434272f $X=5.315 $Y=1.22 $X2=0 $Y2=0
cc_289 N_A3_c_324_n N_VGND_c_638_n 0.00383152f $X=5.745 $Y=1.22 $X2=0 $Y2=0
cc_290 N_A3_c_322_n N_VGND_c_641_n 0.00825283f $X=5.315 $Y=1.22 $X2=0 $Y2=0
cc_291 N_A3_c_324_n N_VGND_c_641_n 0.0075754f $X=5.745 $Y=1.22 $X2=0 $Y2=0
cc_292 N_A3_c_322_n N_A_771_74#_c_743_n 0.0161504f $X=5.315 $Y=1.22 $X2=0 $Y2=0
cc_293 N_A3_c_324_n N_A_771_74#_c_743_n 0.00218762f $X=5.745 $Y=1.22 $X2=0 $Y2=0
cc_294 N_A3_c_326_n N_A_771_74#_c_743_n 0.0173251f $X=5.95 $Y=1.385 $X2=0 $Y2=0
cc_295 N_A3_c_322_n N_A_771_74#_c_745_n 0.013408f $X=5.315 $Y=1.22 $X2=0 $Y2=0
cc_296 N_A3_c_324_n N_A_771_74#_c_745_n 3.97481e-19 $X=5.745 $Y=1.22 $X2=0 $Y2=0
cc_297 N_A_27_368#_c_363_n N_Y_M1000_d 0.00213667f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_298 N_A_27_368#_c_365_n N_Y_M1001_s 0.00218982f $X=2.115 $Y=2.99 $X2=0 $Y2=0
cc_299 N_A_27_368#_c_363_n N_Y_c_460_n 0.0173278f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_300 N_A_27_368#_M1006_s N_Y_c_451_n 0.00218982f $X=1.095 $Y=1.84 $X2=0 $Y2=0
cc_301 N_A_27_368#_c_379_n N_Y_c_451_n 0.0189268f $X=1.28 $Y=2.27 $X2=0 $Y2=0
cc_302 N_A_27_368#_c_365_n N_Y_c_467_n 0.0177084f $X=2.115 $Y=2.99 $X2=0 $Y2=0
cc_303 N_A_27_368#_M1003_d N_Y_c_452_n 0.00218982f $X=2.095 $Y=1.84 $X2=0 $Y2=0
cc_304 N_A_27_368#_c_416_p N_Y_c_452_n 0.0167599f $X=2.257 $Y=2.23 $X2=0 $Y2=0
cc_305 N_A_27_368#_c_385_n N_Y_c_452_n 0.0377698f $X=3.405 $Y=2.145 $X2=0 $Y2=0
cc_306 N_A_27_368#_c_385_n N_Y_c_455_n 0.0157022f $X=3.405 $Y=2.145 $X2=0 $Y2=0
cc_307 N_A_27_368#_c_385_n N_VPWR_M1002_d 0.0138433f $X=3.405 $Y=2.145 $X2=-0.19
+ $Y2=1.66
cc_308 N_A_27_368#_c_390_n N_VPWR_M1004_s 0.0043996f $X=4.42 $Y=2.035 $X2=0
+ $Y2=0
cc_309 N_A_27_368#_c_369_n N_VPWR_M1013_d 0.00274845f $X=5.545 $Y=1.805 $X2=0
+ $Y2=0
cc_310 N_A_27_368#_c_365_n N_VPWR_c_528_n 0.0125197f $X=2.115 $Y=2.99 $X2=0
+ $Y2=0
cc_311 N_A_27_368#_c_385_n N_VPWR_c_528_n 0.0479939f $X=3.405 $Y=2.145 $X2=0
+ $Y2=0
cc_312 N_A_27_368#_c_366_n N_VPWR_c_528_n 0.0252394f $X=3.57 $Y=2.465 $X2=0
+ $Y2=0
cc_313 N_A_27_368#_c_366_n N_VPWR_c_529_n 0.0261113f $X=3.57 $Y=2.465 $X2=0
+ $Y2=0
cc_314 N_A_27_368#_c_390_n N_VPWR_c_529_n 0.0201472f $X=4.42 $Y=2.035 $X2=0
+ $Y2=0
cc_315 N_A_27_368#_c_368_n N_VPWR_c_529_n 0.026897f $X=4.585 $Y=2.4 $X2=0 $Y2=0
cc_316 N_A_27_368#_c_368_n N_VPWR_c_530_n 0.0346454f $X=4.585 $Y=2.4 $X2=0 $Y2=0
cc_317 N_A_27_368#_c_369_n N_VPWR_c_530_n 0.0208278f $X=5.545 $Y=1.805 $X2=0
+ $Y2=0
cc_318 N_A_27_368#_c_370_n N_VPWR_c_530_n 0.0353111f $X=5.71 $Y=1.985 $X2=0
+ $Y2=0
cc_319 N_A_27_368#_c_368_n N_VPWR_c_531_n 0.0201266f $X=4.585 $Y=2.4 $X2=0 $Y2=0
cc_320 N_A_27_368#_c_363_n N_VPWR_c_533_n 0.0421297f $X=1.115 $Y=2.99 $X2=0
+ $Y2=0
cc_321 N_A_27_368#_c_364_n N_VPWR_c_533_n 0.0235688f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_322 N_A_27_368#_c_365_n N_VPWR_c_533_n 0.062575f $X=2.115 $Y=2.99 $X2=0 $Y2=0
cc_323 N_A_27_368#_c_371_n N_VPWR_c_533_n 0.0235512f $X=1.28 $Y=2.99 $X2=0 $Y2=0
cc_324 N_A_27_368#_c_366_n N_VPWR_c_534_n 0.012541f $X=3.57 $Y=2.465 $X2=0 $Y2=0
cc_325 N_A_27_368#_c_370_n N_VPWR_c_535_n 0.014549f $X=5.71 $Y=1.985 $X2=0 $Y2=0
cc_326 N_A_27_368#_c_363_n N_VPWR_c_527_n 0.0236586f $X=1.115 $Y=2.99 $X2=0
+ $Y2=0
cc_327 N_A_27_368#_c_364_n N_VPWR_c_527_n 0.0127152f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_328 N_A_27_368#_c_365_n N_VPWR_c_527_n 0.0347615f $X=2.115 $Y=2.99 $X2=0
+ $Y2=0
cc_329 N_A_27_368#_c_366_n N_VPWR_c_527_n 0.0103123f $X=3.57 $Y=2.465 $X2=0
+ $Y2=0
cc_330 N_A_27_368#_c_368_n N_VPWR_c_527_n 0.0165909f $X=4.585 $Y=2.4 $X2=0 $Y2=0
cc_331 N_A_27_368#_c_370_n N_VPWR_c_527_n 0.0119743f $X=5.71 $Y=1.985 $X2=0
+ $Y2=0
cc_332 N_A_27_368#_c_371_n N_VPWR_c_527_n 0.0126924f $X=1.28 $Y=2.99 $X2=0 $Y2=0
cc_333 N_A_27_368#_c_367_n N_A_771_74#_c_743_n 0.0123321f $X=4.647 $Y=2.12 $X2=0
+ $Y2=0
cc_334 N_A_27_368#_c_369_n N_A_771_74#_c_743_n 0.0242613f $X=5.545 $Y=1.805
+ $X2=0 $Y2=0
cc_335 N_Y_c_452_n N_VPWR_M1002_d 0.00437204f $X=3.005 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_336 N_Y_c_455_n N_VPWR_M1002_d 0.0026139f $X=3.12 $Y=1.72 $X2=-0.19
+ $Y2=-0.245
cc_337 N_Y_c_447_n N_A_27_74#_M1010_s 0.00747698f $X=3.005 $Y=0.925 $X2=0 $Y2=0
cc_338 N_Y_c_451_n N_A_27_74#_c_596_n 0.00589106f $X=1.615 $Y=1.885 $X2=0 $Y2=0
cc_339 N_Y_M1007_d N_A_27_74#_c_598_n 0.00176461f $X=1.48 $Y=0.37 $X2=0 $Y2=0
cc_340 N_Y_c_447_n N_A_27_74#_c_598_n 0.00352531f $X=3.005 $Y=0.925 $X2=0 $Y2=0
cc_341 N_Y_c_474_n N_A_27_74#_c_598_n 0.0154609f $X=1.62 $Y=0.8 $X2=0 $Y2=0
cc_342 N_Y_c_447_n N_A_27_74#_c_600_n 0.0242753f $X=3.005 $Y=0.925 $X2=0 $Y2=0
cc_343 N_Y_c_447_n N_VGND_c_641_n 0.00986599f $X=3.005 $Y=0.925 $X2=0 $Y2=0
cc_344 N_Y_c_447_n N_A_507_74#_M1008_s 0.0052985f $X=3.005 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_345 N_Y_M1008_d N_A_507_74#_c_699_n 0.00176461f $X=2.97 $Y=0.37 $X2=0 $Y2=0
cc_346 N_Y_c_447_n N_A_507_74#_c_699_n 0.0035136f $X=3.005 $Y=0.925 $X2=0 $Y2=0
cc_347 N_Y_c_523_p N_A_507_74#_c_699_n 0.0126348f $X=3.105 $Y=1.01 $X2=0 $Y2=0
cc_348 N_Y_c_448_n N_A_507_74#_c_700_n 0.00523541f $X=3.12 $Y=1.235 $X2=0 $Y2=0
cc_349 N_Y_c_447_n N_A_507_74#_c_703_n 0.0206029f $X=3.005 $Y=0.925 $X2=0 $Y2=0
cc_350 N_Y_c_448_n N_A_771_74#_c_744_n 0.00159757f $X=3.12 $Y=1.235 $X2=0 $Y2=0
cc_351 N_A_27_74#_c_596_n N_VGND_M1011_s 0.00229612f $X=1.105 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_352 N_A_27_74#_c_595_n N_VGND_c_632_n 0.0164982f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_353 N_A_27_74#_c_596_n N_VGND_c_632_n 0.0193595f $X=1.105 $Y=1.045 $X2=0
+ $Y2=0
cc_354 N_A_27_74#_c_599_n N_VGND_c_632_n 0.00814404f $X=1.275 $Y=0.34 $X2=0
+ $Y2=0
cc_355 N_A_27_74#_c_595_n N_VGND_c_636_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_356 N_A_27_74#_c_598_n N_VGND_c_637_n 0.042902f $X=1.955 $Y=0.34 $X2=0 $Y2=0
cc_357 N_A_27_74#_c_599_n N_VGND_c_637_n 0.0121867f $X=1.275 $Y=0.34 $X2=0 $Y2=0
cc_358 N_A_27_74#_c_600_n N_VGND_c_637_n 0.0226635f $X=2.12 $Y=0.34 $X2=0 $Y2=0
cc_359 N_A_27_74#_c_595_n N_VGND_c_641_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_360 N_A_27_74#_c_598_n N_VGND_c_641_n 0.0241973f $X=1.955 $Y=0.34 $X2=0 $Y2=0
cc_361 N_A_27_74#_c_599_n N_VGND_c_641_n 0.00660921f $X=1.275 $Y=0.34 $X2=0
+ $Y2=0
cc_362 N_A_27_74#_c_600_n N_VGND_c_641_n 0.0125932f $X=2.12 $Y=0.34 $X2=0 $Y2=0
cc_363 N_A_27_74#_c_600_n N_A_507_74#_c_703_n 0.0279789f $X=2.12 $Y=0.34 $X2=0
+ $Y2=0
cc_364 N_VGND_c_637_n N_A_507_74#_c_699_n 0.0333877f $X=4.935 $Y=0 $X2=0 $Y2=0
cc_365 N_VGND_c_641_n N_A_507_74#_c_699_n 0.0187857f $X=6 $Y=0 $X2=0 $Y2=0
cc_366 N_VGND_c_633_n N_A_507_74#_c_701_n 0.011925f $X=5.1 $Y=0.675 $X2=0 $Y2=0
cc_367 N_VGND_c_637_n N_A_507_74#_c_701_n 0.065612f $X=4.935 $Y=0 $X2=0 $Y2=0
cc_368 N_VGND_c_641_n N_A_507_74#_c_701_n 0.0365975f $X=6 $Y=0 $X2=0 $Y2=0
cc_369 N_VGND_c_633_n N_A_507_74#_c_702_n 0.0273691f $X=5.1 $Y=0.675 $X2=0 $Y2=0
cc_370 N_VGND_c_637_n N_A_507_74#_c_703_n 0.0225845f $X=4.935 $Y=0 $X2=0 $Y2=0
cc_371 N_VGND_c_641_n N_A_507_74#_c_703_n 0.0124836f $X=6 $Y=0 $X2=0 $Y2=0
cc_372 N_VGND_c_637_n N_A_507_74#_c_704_n 0.0235688f $X=4.935 $Y=0 $X2=0 $Y2=0
cc_373 N_VGND_c_641_n N_A_507_74#_c_704_n 0.0127152f $X=6 $Y=0 $X2=0 $Y2=0
cc_374 N_VGND_M1005_s N_A_771_74#_c_743_n 0.00299905f $X=4.955 $Y=0.37 $X2=0
+ $Y2=0
cc_375 N_VGND_c_633_n N_A_771_74#_c_743_n 0.0201544f $X=5.1 $Y=0.675 $X2=0 $Y2=0
cc_376 N_VGND_c_633_n N_A_771_74#_c_745_n 0.0175587f $X=5.1 $Y=0.675 $X2=0 $Y2=0
cc_377 N_VGND_c_635_n N_A_771_74#_c_745_n 0.0243832f $X=5.96 $Y=0.515 $X2=0
+ $Y2=0
cc_378 N_VGND_c_638_n N_A_771_74#_c_745_n 0.0109942f $X=5.795 $Y=0 $X2=0 $Y2=0
cc_379 N_VGND_c_641_n N_A_771_74#_c_745_n 0.00904371f $X=6 $Y=0 $X2=0 $Y2=0
cc_380 N_A_507_74#_c_701_n N_A_771_74#_M1012_s 0.0030917f $X=4.375 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_381 N_A_507_74#_c_701_n N_A_771_74#_c_766_n 0.0211419f $X=4.375 $Y=0.34 $X2=0
+ $Y2=0
cc_382 N_A_507_74#_M1014_d N_A_771_74#_c_743_n 0.00299905f $X=4.4 $Y=0.37 $X2=0
+ $Y2=0
cc_383 N_A_507_74#_c_701_n N_A_771_74#_c_743_n 0.00304353f $X=4.375 $Y=0.34
+ $X2=0 $Y2=0
cc_384 N_A_507_74#_c_702_n N_A_771_74#_c_743_n 0.021673f $X=4.54 $Y=0.675 $X2=0
+ $Y2=0
cc_385 N_A_507_74#_c_700_n N_A_771_74#_c_744_n 0.00585736f $X=3.54 $Y=0.515
+ $X2=0 $Y2=0

* File: sky130_fd_sc_ms__sdlclkp_2.spice
* Created: Wed Sep  2 12:32:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdlclkp_2.pex.spice"
.subckt sky130_fd_sc_ms__sdlclkp_2  VNB VPB SCE GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1015 N_A_114_112#_M1015_d N_SCE_M1015_g N_VGND_M1015_s VNB NLOWVT L=0.15
+ W=0.55 AD=0.077 AS=0.15675 PD=0.83 PS=1.67 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.2 A=0.0825 P=1.4 MULT=1
MM1014 N_VGND_M1014_d N_GATE_M1014_g N_A_114_112#_M1015_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.161184 AS=0.077 PD=1.20233 PS=0.83 NRD=51.936 NRS=0 M=1 R=3.66667
+ SA=75000.6 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1006 N_A_318_74#_M1006_d N_A_288_48#_M1006_g N_VGND_M1014_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.216866 PD=2.05 PS=1.61767 NRD=0 NRS=38.604 M=1 R=4.93333
+ SA=75001 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1023 N_A_580_74#_M1023_d N_A_288_48#_M1023_g N_A_114_112#_M1023_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.110425 AS=0.33275 PD=1.04897 PS=2.31 NRD=2.172 NRS=69.816
+ M=1 R=3.66667 SA=75000.5 SB=75001.4 A=0.0825 P=1.4 MULT=1
MM1018 A_685_81# N_A_318_74#_M1018_g N_A_580_74#_M1023_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0843247 PD=0.66 PS=0.801031 NRD=18.564 NRS=24.276 M=1
+ R=2.8 SA=75001.1 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_706_317#_M1019_g A_685_81# VNB NLOWVT L=0.15 W=0.42
+ AD=0.109562 AS=0.0504 PD=0.919655 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75001.4 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1004 N_A_706_317#_M1004_d N_A_580_74#_M1004_g N_VGND_M1019_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.193038 PD=2.05 PS=1.62034 NRD=0 NRS=40.536 M=1 R=4.93333
+ SA=75001.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_CLK_M1002_g N_A_288_48#_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.13135 AS=0.2109 PD=1.095 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1016 A_1198_74# N_CLK_M1016_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.0777 AS=0.13135 PD=0.95 PS=1.095 NRD=8.1 NRS=0.804 M=1 R=4.93333
+ SA=75000.7 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1011 N_A_1198_374#_M1011_d N_A_706_317#_M1011_g A_1198_74# VNB NLOWVT L=0.15
+ W=0.74 AD=0.2035 AS=0.0777 PD=2.03 PS=0.95 NRD=0 NRS=8.1 M=1 R=4.93333
+ SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_GCLK_M1009_d N_A_1198_374#_M1009_g N_VGND_M1009_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2035 PD=1.02 PS=2.03 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1017 N_GCLK_M1009_d N_A_1198_374#_M1017_g N_VGND_M1017_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2035 PD=1.02 PS=2.03 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1022 A_117_424# N_SCE_M1022_g N_VPWR_M1022_s VPB PSHORT L=0.18 W=0.84
+ AD=0.0882 AS=0.2268 PD=1.05 PS=2.22 NRD=11.7215 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.6 A=0.1512 P=2.04 MULT=1
MM1008 N_A_114_112#_M1008_d N_GATE_M1008_g A_117_424# VPB PSHORT L=0.18 W=0.84
+ AD=0.2268 AS=0.0882 PD=2.22 PS=1.05 NRD=0 NRS=11.7215 M=1 R=4.66667 SA=90000.6
+ SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1012 N_A_318_74#_M1012_d N_A_288_48#_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18
+ W=0.84 AD=0.2268 AS=0.3681 PD=2.22 PS=2.95 NRD=0 NRS=89.8714 M=1 R=4.66667
+ SA=90000.3 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1005 N_A_580_74#_M1005_d N_A_318_74#_M1005_g N_A_114_112#_M1005_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1722 AS=0.2268 PD=1.58 PS=2.22 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90000.9 A=0.1512 P=2.04 MULT=1
MM1013 A_711_451# N_A_288_48#_M1013_g N_A_580_74#_M1005_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0441 AS=0.0861 PD=0.63 PS=0.79 NRD=23.443 NRS=32.8202 M=1
+ R=2.33333 SA=90000.7 SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1007 N_VPWR_M1007_d N_A_706_317#_M1007_g A_711_451# VPB PSHORT L=0.18 W=0.42
+ AD=0.0910636 AS=0.0441 PD=0.799091 PS=0.63 NRD=35.1645 NRS=23.443 M=1
+ R=2.33333 SA=90001.1 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1000 N_A_706_317#_M1000_d N_A_580_74#_M1000_g N_VPWR_M1007_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3024 AS=0.242836 PD=2.78 PS=2.13091 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.7 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1010 N_VPWR_M1010_d N_CLK_M1010_g N_A_288_48#_M1010_s VPB PSHORT L=0.18 W=0.84
+ AD=0.16469 AS=0.2268 PD=1.3513 PS=2.22 NRD=33.0763 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90002.1 A=0.1512 P=2.04 MULT=1
MM1021 N_A_1198_374#_M1021_d N_CLK_M1021_g N_VPWR_M1010_d VPB PSHORT L=0.18 W=1
+ AD=0.2425 AS=0.19606 PD=1.485 PS=1.6087 NRD=41.3503 NRS=0 M=1 R=5.55556
+ SA=90000.6 SB=90001.9 A=0.18 P=2.36 MULT=1
MM1020 N_VPWR_M1020_d N_A_706_317#_M1020_g N_A_1198_374#_M1021_d VPB PSHORT
+ L=0.18 W=1 AD=0.208585 AS=0.2425 PD=1.43868 PS=1.485 NRD=16.2328 NRS=0 M=1
+ R=5.55556 SA=90001.2 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1001 N_GCLK_M1001_d N_A_1198_374#_M1001_g N_VPWR_M1020_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.233615 PD=1.39 PS=1.61132 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90001.6 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1003 N_GCLK_M1001_d N_A_1198_374#_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX24_noxref VNB VPB NWDIODE A=16.0894 P=21
*
.include "sky130_fd_sc_ms__sdlclkp_2.pxi.spice"
*
.ends
*
*

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__o41a_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__o41a_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.297600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.610000 1.350000 4.195000 2.150000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.297600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.300000 3.370000 2.890000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.297600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.470000 1.220000 2.800000 2.890000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.297600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.870000 1.190000 2.275000 1.780000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.247200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.450000 1.580000 1.780000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  0.524500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.350000 0.375000 1.130000 ;
        RECT 0.115000 1.130000 0.285000 2.290000 ;
        RECT 0.115000 2.290000 0.445000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.455000  1.350000 0.785000 1.950000 ;
      RECT 0.455000  1.950000 2.080000 2.120000 ;
      RECT 0.545000  0.085000 0.945000 0.940000 ;
      RECT 0.615000  1.110000 1.505000 1.280000 ;
      RECT 0.615000  1.280000 0.785000 1.350000 ;
      RECT 0.615000  2.290000 1.540000 3.245000 ;
      RECT 1.175000  0.350000 1.505000 1.110000 ;
      RECT 1.675000  0.350000 2.005000 0.850000 ;
      RECT 1.675000  0.850000 4.205000 1.020000 ;
      RECT 1.750000  2.120000 2.080000 2.845000 ;
      RECT 2.175000  0.085000 2.505000 0.680000 ;
      RECT 2.675000  0.350000 3.005000 0.850000 ;
      RECT 3.175000  0.085000 3.705000 0.680000 ;
      RECT 3.760000  2.320000 4.205000 3.245000 ;
      RECT 3.875000  0.350000 4.205000 0.850000 ;
      RECT 3.875000  1.020000 4.205000 1.030000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_ms__o41a_1
END LIBRARY

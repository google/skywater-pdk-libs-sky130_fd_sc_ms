* File: sky130_fd_sc_ms__a2111o_1.pex.spice
* Created: Wed Sep  2 11:49:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A2111O_1%A1 1 3 8 10 11 15 16 19
r37 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.675 $Y=0.405
+ $X2=0.675 $Y2=0.57
r38 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.675
+ $Y=0.405 $X2=0.675 $Y2=0.405
r39 11 16 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.675 $Y=0.555
+ $X2=0.675 $Y2=0.405
r40 11 19 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.675 $Y=0.555
+ $X2=0.51 $Y2=0.555
r41 10 19 13.5287 $w=2.28e-07 $l=2.7e-07 $layer=LI1_cond $X=0.24 $Y=0.555
+ $X2=0.51 $Y2=0.555
r42 8 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.765 $Y=1 $X2=0.765
+ $Y2=1.395
r43 8 18 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.765 $Y=1 $X2=0.765
+ $Y2=0.57
r44 1 9 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.75 $Y=1.485 $X2=0.75
+ $Y2=1.395
r45 1 3 378.992 $w=1.8e-07 $l=9.75e-07 $layer=POLY_cond $X=0.75 $Y=1.485
+ $X2=0.75 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A2111O_1%A2 3 7 9 10 11 16
c41 7 0 1.41057e-19 $X=1.24 $Y=2.46
c42 3 0 1.36987e-19 $X=1.125 $Y=1
r43 16 19 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.215 $Y=1.635
+ $X2=1.215 $Y2=1.8
r44 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.215 $Y=1.635
+ $X2=1.215 $Y2=1.47
r45 10 11 18.4391 $w=2.98e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.65
+ $X2=2.16 $Y2=1.65
r46 9 10 18.4391 $w=2.98e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.65 $X2=1.68
+ $Y2=1.65
r47 9 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.215
+ $Y=1.635 $X2=1.215 $Y2=1.635
r48 7 19 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.24 $Y=2.46 $X2=1.24
+ $Y2=1.8
r49 3 18 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.125 $Y=1 $X2=1.125
+ $Y2=1.47
.ends

.subckt PM_SKY130_FD_SC_MS__A2111O_1%B1 4 7 10 11 14
c41 11 0 1.36987e-19 $X=1.68 $Y=0.555
c42 4 0 3.01101e-20 $X=1.665 $Y=1
r43 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.6 $Y=0.37 $X2=1.6
+ $Y2=0.535
r44 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=0.37 $X2=1.6 $Y2=0.37
r45 11 15 7.78276 $w=2.9e-07 $l=1.85e-07 $layer=LI1_cond $X=1.615 $Y=0.555
+ $X2=1.615 $Y2=0.37
r46 9 10 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=1.685 $Y=1.395
+ $X2=1.685 $Y2=1.545
r47 7 10 355.669 $w=1.8e-07 $l=9.15e-07 $layer=POLY_cond $X=1.69 $Y=2.46
+ $X2=1.69 $Y2=1.545
r48 4 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.665 $Y=1 $X2=1.665
+ $Y2=1.395
r49 4 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.665 $Y=1 $X2=1.665
+ $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_MS__A2111O_1%C1 1 3 8 10 13
c42 10 0 3.31031e-20 $X=2.16 $Y=0.555
c43 8 0 3.01101e-20 $X=2.095 $Y=1
r44 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=0.37
+ $X2=2.17 $Y2=0.535
r45 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.17
+ $Y=0.37 $X2=2.17 $Y2=0.37
r46 10 14 7.78276 $w=2.9e-07 $l=1.85e-07 $layer=LI1_cond $X=2.17 $Y=0.555
+ $X2=2.17 $Y2=0.37
r47 8 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.095 $Y=1 $X2=2.095
+ $Y2=1.395
r48 8 16 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.095 $Y=1 $X2=2.095
+ $Y2=0.535
r49 1 9 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.08 $Y=1.485 $X2=2.08
+ $Y2=1.395
r50 1 3 378.992 $w=1.8e-07 $l=9.75e-07 $layer=POLY_cond $X=2.08 $Y=1.485
+ $X2=2.08 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A2111O_1%D1 3 7 9 16
c33 9 0 1.05647e-19 $X=2.64 $Y=1.665
r34 14 16 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=2.61 $Y=1.635
+ $X2=2.715 $Y2=1.635
r35 11 14 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=2.47 $Y=1.635
+ $X2=2.61 $Y2=1.635
r36 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.635 $X2=2.61 $Y2=1.635
r37 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.715 $Y=1.47
+ $X2=2.715 $Y2=1.635
r38 5 7 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.715 $Y=1.47 $X2=2.715
+ $Y2=1
r39 1 11 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.47 $Y=1.8 $X2=2.47
+ $Y2=1.635
r40 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.47 $Y=1.8 $X2=2.47
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A2111O_1%A_85_136# 1 2 3 4 15 19 21 22 23 25 29 33
+ 36 39 43 48 55 57
c95 33 0 3.31031e-20 $X=2.93 $Y=0.825
c96 25 0 3.01101e-20 $X=2.845 $Y=1.245
c97 23 0 3.01101e-20 $X=1.715 $Y=1.245
c98 21 0 1.05647e-19 $X=3.71 $Y=1.485
r99 53 55 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.695 $Y=2.055
+ $X2=3.03 $Y2=2.055
r100 48 50 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.88 $Y=1.085
+ $X2=1.88 $Y2=1.245
r101 43 45 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=0.55 $Y=1.09
+ $X2=0.55 $Y2=1.245
r102 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.525
+ $Y=1.485 $X2=3.525 $Y2=1.485
r103 37 57 2.66945 $w=3.3e-07 $l=4.39744e-07 $layer=LI1_cond $X=3.115 $Y=1.485
+ $X2=2.845 $Y2=1.16
r104 37 39 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.115 $Y=1.485
+ $X2=3.525 $Y2=1.485
r105 36 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=1.97
+ $X2=3.03 $Y2=2.055
r106 35 57 3.44865 $w=1.7e-07 $l=5.75109e-07 $layer=LI1_cond $X=3.03 $Y=1.65
+ $X2=2.845 $Y2=1.16
r107 35 36 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.03 $Y=1.65
+ $X2=3.03 $Y2=1.97
r108 31 57 3.44865 $w=2.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.98 $Y=1.16
+ $X2=2.845 $Y2=1.16
r109 31 33 14.2988 $w=2.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.98 $Y=1.16
+ $X2=2.98 $Y2=0.825
r110 29 53 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.695 $Y=2.815
+ $X2=2.695 $Y2=2.14
r111 26 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.045 $Y=1.245
+ $X2=1.88 $Y2=1.245
r112 25 57 2.66945 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.845 $Y=1.245
+ $X2=2.845 $Y2=1.16
r113 25 26 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=2.845 $Y=1.245
+ $X2=2.045 $Y2=1.245
r114 24 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.715 $Y=1.245
+ $X2=0.55 $Y2=1.245
r115 23 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.715 $Y=1.245
+ $X2=1.88 $Y2=1.245
r116 23 24 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=1.715 $Y=1.245
+ $X2=0.715 $Y2=1.245
r117 21 40 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=3.71 $Y=1.485
+ $X2=3.525 $Y2=1.485
r118 21 22 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.71 $Y=1.485 $X2=3.8
+ $Y2=1.485
r119 17 22 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=3.815 $Y=1.32
+ $X2=3.8 $Y2=1.485
r120 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.815 $Y=1.32
+ $X2=3.815 $Y2=0.76
r121 13 22 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=3.8 $Y=1.65
+ $X2=3.8 $Y2=1.485
r122 13 15 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=3.8 $Y=1.65 $X2=3.8
+ $Y2=2.4
r123 4 53 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.56
+ $Y=1.96 $X2=2.695 $Y2=2.135
r124 4 29 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.56
+ $Y=1.96 $X2=2.695 $Y2=2.815
r125 3 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.79
+ $Y=0.68 $X2=2.93 $Y2=0.825
r126 2 48 182 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_NDIFF $count=1 $X=1.74
+ $Y=0.68 $X2=1.88 $Y2=1.085
r127 1 43 182 $w=1.7e-07 $l=4.68348e-07 $layer=licon1_NDIFF $count=1 $X=0.425
+ $Y=0.68 $X2=0.55 $Y2=1.09
.ends

.subckt PM_SKY130_FD_SC_MS__A2111O_1%A_80_392# 1 2 7 9 11 13 15
c29 7 0 1.41057e-19 $X=0.525 $Y=2.14
r30 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.465 $Y=2.14
+ $X2=1.465 $Y2=2.055
r31 13 15 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.465 $Y=2.14
+ $X2=1.465 $Y2=2.815
r32 12 18 4.99254 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.69 $Y=2.055
+ $X2=0.525 $Y2=2.04
r33 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.3 $Y=2.055
+ $X2=1.465 $Y2=2.055
r34 11 12 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.3 $Y=2.055
+ $X2=0.69 $Y2=2.055
r35 7 18 2.77363 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=0.525 $Y=2.14 $X2=0.525
+ $Y2=2.04
r36 7 9 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.525 $Y=2.14
+ $X2=0.525 $Y2=2.815
r37 2 20 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.33
+ $Y=1.96 $X2=1.465 $Y2=2.135
r38 2 15 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.33
+ $Y=1.96 $X2=1.465 $Y2=2.815
r39 1 18 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.4
+ $Y=1.96 $X2=0.525 $Y2=2.105
r40 1 9 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.4
+ $Y=1.96 $X2=0.525 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__A2111O_1%VPWR 1 2 9 13 18 19 21 22 23 36 37
r42 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r43 34 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r44 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 30 33 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 27 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 23 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r50 23 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r51 21 33 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.41 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 21 22 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.41 $Y=3.33
+ $X2=3.535 $Y2=3.33
r53 20 36 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.66 $Y=3.33
+ $X2=4.08 $Y2=3.33
r54 20 22 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.66 $Y=3.33
+ $X2=3.535 $Y2=3.33
r55 18 26 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.89 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 18 19 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.89 $Y=3.33
+ $X2=0.995 $Y2=3.33
r57 17 30 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=1.1 $Y=3.33 $X2=1.2
+ $Y2=3.33
r58 17 19 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.1 $Y=3.33
+ $X2=0.995 $Y2=3.33
r59 13 16 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=3.535 $Y=1.985
+ $X2=3.535 $Y2=2.815
r60 11 22 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=3.245
+ $X2=3.535 $Y2=3.33
r61 11 16 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=3.535 $Y=3.245
+ $X2=3.535 $Y2=2.815
r62 7 19 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.995 $Y=3.245
+ $X2=0.995 $Y2=3.33
r63 7 9 40.6667 $w=2.08e-07 $l=7.7e-07 $layer=LI1_cond $X=0.995 $Y=3.245
+ $X2=0.995 $Y2=2.475
r64 2 16 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=3.45
+ $Y=1.84 $X2=3.575 $Y2=2.815
r65 2 13 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.45
+ $Y=1.84 $X2=3.575 $Y2=1.985
r66 1 9 300 $w=1.7e-07 $l=5.8741e-07 $layer=licon1_PDIFF $count=2 $X=0.84
+ $Y=1.96 $X2=0.995 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_MS__A2111O_1%X 1 2 7 8 9 10 11 12 13
r12 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=4.027 $Y=2.405
+ $X2=4.027 $Y2=2.775
r13 11 12 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=4.027 $Y=1.985
+ $X2=4.027 $Y2=2.405
r14 10 11 11.0084 $w=3.33e-07 $l=3.2e-07 $layer=LI1_cond $X=4.027 $Y=1.665
+ $X2=4.027 $Y2=1.985
r15 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=4.027 $Y=1.295
+ $X2=4.027 $Y2=1.665
r16 8 9 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=4.027 $Y=0.925
+ $X2=4.027 $Y2=1.295
r17 7 8 13.4165 $w=3.33e-07 $l=3.9e-07 $layer=LI1_cond $X=4.027 $Y=0.535
+ $X2=4.027 $Y2=0.925
r18 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.84 $X2=4.025 $Y2=2.815
r19 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.84 $X2=4.025 $Y2=1.985
r20 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.89
+ $Y=0.39 $X2=4.03 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_MS__A2111O_1%VGND 1 2 3 11 13 16 21 26 29 30 31 33 42 48
+ 49 52 55
r71 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r72 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r73 49 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r74 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r75 46 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.56
+ $Y2=0
r76 46 48 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.685 $Y=0 $X2=4.08
+ $Y2=0
r77 45 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r78 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r79 42 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.435 $Y=0 $X2=3.56
+ $Y2=0
r80 42 44 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.435 $Y=0 $X2=3.12
+ $Y2=0
r81 38 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.18
+ $Y2=0
r82 38 40 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=2.16
+ $Y2=0
r83 36 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r84 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r85 33 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=0 $X2=1.18
+ $Y2=0
r86 33 35 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.095 $Y=0 $X2=0.72
+ $Y2=0
r87 31 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r88 31 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r89 31 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r90 29 40 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.505 $Y=0 $X2=2.16
+ $Y2=0
r91 29 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=0 $X2=2.59
+ $Y2=0
r92 28 44 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.675 $Y=0 $X2=3.12
+ $Y2=0
r93 28 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.59
+ $Y2=0
r94 24 26 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.5 $Y=0.825 $X2=2.59
+ $Y2=0.825
r95 18 21 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.18 $Y=0.825
+ $X2=1.34 $Y2=0.825
r96 14 55 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.56 $Y=0.085
+ $X2=3.56 $Y2=0
r97 14 16 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=3.56 $Y=0.085
+ $X2=3.56 $Y2=0.535
r98 13 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.59 $Y=0.66
+ $X2=2.59 $Y2=0.825
r99 12 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=0.085
+ $X2=2.59 $Y2=0
r100 12 13 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.59 $Y=0.085
+ $X2=2.59 $Y2=0.66
r101 11 18 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.18 $Y=0.66
+ $X2=1.18 $Y2=0.825
r102 10 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.18 $Y2=0
r103 10 11 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.18 $Y2=0.66
r104 3 16 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=3.475
+ $Y=0.39 $X2=3.6 $Y2=0.535
r105 2 24 182 $w=1.7e-07 $l=3.95917e-07 $layer=licon1_NDIFF $count=1 $X=2.17
+ $Y=0.68 $X2=2.5 $Y2=0.825
r106 1 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.2
+ $Y=0.68 $X2=1.34 $Y2=0.825
.ends


* NGSPICE file created from sky130_fd_sc_ms__dlrtn_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__dlrtn_1 D GATE_N RESET_B VGND VNB VPB VPWR Q
M1000 a_232_98# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=1.64835e+12p ps=1.063e+07u
M1001 VGND a_897_406# a_854_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
M1002 Q a_897_406# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=1.70685e+12p ps=1.247e+07u
M1003 a_854_74# a_357_392# a_657_392# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.915e+11p ps=1.93e+06u
M1004 a_573_392# a_27_136# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1005 a_232_98# GATE_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1006 a_796_508# a_232_98# a_657_392# VPB pshort w=420000u l=180000u
+  ad=2.121e+11p pd=1.85e+06u as=3.816e+11p ps=3.03e+06u
M1007 VPWR a_897_406# a_796_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND RESET_B a_1139_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1009 VPWR a_232_98# a_357_392# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1010 a_681_74# a_27_136# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1011 VPWR RESET_B a_897_406# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=4.4e+11p ps=2.88e+06u
M1012 VPWR D a_27_136# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1013 VGND D a_27_136# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1014 a_1139_74# a_657_392# a_897_406# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1015 Q a_897_406# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.701e+11p pd=2.21e+06u as=0p ps=0u
M1016 VGND a_232_98# a_357_392# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1017 a_657_392# a_232_98# a_681_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_657_392# a_357_392# a_573_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_897_406# a_657_392# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


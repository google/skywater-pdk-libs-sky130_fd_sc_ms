* File: sky130_fd_sc_ms__dfrtn_1.spice
* Created: Wed Sep  2 12:02:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dfrtn_1.pex.spice"
.subckt sky130_fd_sc_ms__dfrtn_1  VNB VPB D CLK_N RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* CLK_N	CLK_N
* D	D
* VPB	VPB
* VNB	VNB
MM1028 A_120_74# N_D_M1028_g N_A_33_74#_M1028_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_RESET_B_M1024_g A_120_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0504 PD=1.37 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_CLK_N_M1013_g N_A_300_347#_M1013_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.14615 AS=0.2442 PD=1.135 PS=2.14 NRD=8.916 NRS=3.24 M=1 R=4.93333
+ SA=75000.3 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1011 N_A_510_74#_M1011_d N_A_300_347#_M1011_g N_VGND_M1013_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2257 AS=0.14615 PD=2.09 PS=1.135 NRD=6.48 NRS=9.72 M=1 R=4.93333
+ SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_A_714_119#_M1006_d N_A_510_74#_M1006_g N_A_33_74#_M1006_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1113 PD=0.95 PS=1.37 NRD=71.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75005.7 A=0.063 P=1.14 MULT=1
MM1019 A_850_119# N_A_300_347#_M1019_g N_A_714_119#_M1006_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=0.95 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75005 A=0.063 P=1.14 MULT=1
MM1016 A_922_119# N_A_856_294#_M1016_g A_850_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75001.2
+ SB=75004.7 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_RESET_B_M1009_g A_922_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.167584 AS=0.0441 PD=1.2419 PS=0.63 NRD=24.276 NRS=14.28 M=1 R=2.8
+ SA=75001.6 SB=75004.3 A=0.063 P=1.14 MULT=1
MM1020 N_A_856_294#_M1020_d N_A_714_119#_M1020_g N_VGND_M1009_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1073 AS=0.295266 PD=1.03 PS=2.1881 NRD=0 NRS=55.776 M=1
+ R=4.93333 SA=75001.5 SB=75002.2 A=0.111 P=1.78 MULT=1
MM1007 N_A_1266_119#_M1007_d N_A_300_347#_M1007_g N_A_856_294#_M1020_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.391307 AS=0.1073 PD=2.56448 PS=1.03 NRD=51.888
+ NRS=1.62 M=1 R=4.93333 SA=75001.9 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1022 A_1550_119# N_A_510_74#_M1022_g N_A_1266_119#_M1007_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.222093 PD=0.66 PS=1.45552 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75004.4 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_1598_93#_M1002_g A_1550_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0504 PD=0.81 PS=0.66 NRD=15.708 NRS=18.564 M=1 R=2.8 SA=75004.8
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1010 A_1736_119# N_RESET_B_M1010_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0819 PD=0.66 PS=0.81 NRD=18.564 NRS=15.708 M=1 R=2.8 SA=75005.3
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_A_1598_93#_M1004_d N_A_1266_119#_M1004_g A_1736_119# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75005.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_A_1266_119#_M1021_g N_A_1934_94#_M1021_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.107506 AS=0.15675 PD=0.937984 PS=1.67 NRD=18 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1027 N_Q_M1027_d N_A_1934_94#_M1027_g N_VGND_M1021_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2146 AS=0.144644 PD=2.06 PS=1.26202 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1030 N_A_33_74#_M1030_d N_D_M1030_g N_VPWR_M1030_s VPB PSHORT L=0.18 W=0.42
+ AD=0.0567 AS=0.1155 PD=0.69 PS=1.39 NRD=0 NRS=0 M=1 R=2.33333 SA=90000.2
+ SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1031 N_VPWR_M1031_d N_RESET_B_M1031_g N_A_33_74#_M1030_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1113 AS=0.0567 PD=1.37 PS=0.69 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1017 N_VPWR_M1017_d N_CLK_N_M1017_g N_A_300_347#_M1017_s VPB PSHORT L=0.18 W=1
+ AD=0.210787 AS=0.29575 PD=1.47 PS=2.65 NRD=12.7853 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1003 N_A_510_74#_M1003_d N_A_300_347#_M1003_g N_VPWR_M1017_d VPB PSHORT L=0.18
+ W=1 AD=0.265 AS=0.210787 PD=2.53 PS=1.47 NRD=0 NRS=11.8003 M=1 R=5.55556
+ SA=90000.8 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1012 N_A_714_119#_M1012_d N_A_300_347#_M1012_g N_A_33_74#_M1012_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0567 AS=0.1176 PD=0.69 PS=1.4 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90001.5 A=0.0756 P=1.2 MULT=1
MM1014 A_820_457# N_A_510_74#_M1014_g N_A_714_119#_M1012_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0441 AS=0.0567 PD=0.63 PS=0.69 NRD=23.443 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1005 N_VPWR_M1005_d N_A_856_294#_M1005_g A_820_457# VPB PSHORT L=0.18 W=0.42
+ AD=0.0693 AS=0.0441 PD=0.75 PS=0.63 NRD=11.7215 NRS=23.443 M=1 R=2.33333
+ SA=90001 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1018 N_A_714_119#_M1018_d N_RESET_B_M1018_g N_VPWR_M1005_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1092 AS=0.0693 PD=1.36 PS=0.75 NRD=0 NRS=11.7215 M=1 R=2.33333
+ SA=90001.5 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1000 N_A_856_294#_M1000_d N_A_714_119#_M1000_g N_VPWR_M1000_s VPB PSHORT
+ L=0.18 W=1 AD=0.375 AS=0.26 PD=1.75 PS=2.52 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90002 A=0.18 P=2.36 MULT=1
MM1001 N_A_1266_119#_M1001_d N_A_510_74#_M1001_g N_A_856_294#_M1000_d VPB PSHORT
+ L=0.18 W=1 AD=0.300282 AS=0.375 PD=2.35211 PS=1.75 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90001.1 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1029 A_1550_508# N_A_300_347#_M1029_g N_A_1266_119#_M1001_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.126118 PD=0.66 PS=0.987887 NRD=30.4759 NRS=0 M=1
+ R=2.33333 SA=90001.9 SB=90001.6 A=0.0756 P=1.2 MULT=1
MM1008 N_VPWR_M1008_d N_A_1598_93#_M1008_g A_1550_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.0756 AS=0.0504 PD=0.78 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.33333 SA=90002.4
+ SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1015 N_A_1598_93#_M1015_d N_RESET_B_M1015_g N_VPWR_M1008_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0567 AS=0.0756 PD=0.69 PS=0.78 NRD=0 NRS=39.8531 M=1 R=2.33333
+ SA=90002.9 SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1023 N_VPWR_M1023_d N_A_1266_119#_M1023_g N_A_1598_93#_M1015_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90003.4 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1025 N_VPWR_M1025_d N_A_1266_119#_M1025_g N_A_1934_94#_M1025_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.147 AS=0.2184 PD=1.23857 PS=2.2 NRD=10.5395 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1026 N_Q_M1026_d N_A_1934_94#_M1026_g N_VPWR_M1025_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3024 AS=0.196 PD=2.78 PS=1.65143 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX32_noxref VNB VPB NWDIODE A=21.3751 P=26.8
c_118 VNB 0 4.82778e-19 $X=0 $Y=0
c_231 VPB 0 1.58987e-19 $X=0 $Y=3.085
c_1630 A_120_74# 0 1.52323e-19 $X=0.6 $Y=0.37
*
.include "sky130_fd_sc_ms__dfrtn_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__sdfrbp_2.spice
* Created: Fri Aug 28 18:11:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdfrbp_2.pex.spice"
.subckt sky130_fd_sc_ms__sdfrbp_2  VNB VPB SCE D SCD CLK RESET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1030 N_VGND_M1030_d N_SCE_M1030_g N_A_27_79#_M1030_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1155 AS=0.1197 PD=1.39 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 noxref_26 N_A_27_79#_M1012_g N_noxref_25_M1012_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1026 N_A_388_79#_M1026_d N_D_M1026_g noxref_26 VNB NLOWVT L=0.15 W=0.42
+ AD=0.13545 AS=0.0504 PD=1.065 PS=0.66 NRD=101.424 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1031 noxref_27 N_SCE_M1031_g N_A_388_79#_M1026_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.13545 PD=0.66 PS=1.065 NRD=18.564 NRS=2.856 M=1 R=2.8
+ SA=75001.4 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1013 N_noxref_25_M1013_d N_SCD_M1013_g noxref_27 VNB NLOWVT L=0.15 W=0.42
+ AD=0.0777 AS=0.0504 PD=0.79 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.8
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_RESET_B_M1003_g N_noxref_25_M1013_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.1281 AS=0.0777 PD=1.45 PS=0.79 NRD=5.712 NRS=25.704 M=1 R=2.8
+ SA=75002.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_CLK_M1021_g N_A_852_119#_M1021_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.195675 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1033 N_A_1025_119#_M1033_d N_A_852_119#_M1033_g N_VGND_M1021_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1014 N_A_1223_119#_M1014_d N_A_852_119#_M1014_g N_A_388_79#_M1014_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004 A=0.063 P=1.14 MULT=1
MM1015 A_1323_119# N_A_1025_119#_M1015_g N_A_1223_119#_M1014_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1043 A_1401_119# N_A_1370_290#_M1043_g A_1323_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75003.1 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_RESET_B_M1011_g A_1401_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.279132 AS=0.0504 PD=1.43434 PS=0.66 NRD=174.168 NRS=18.564 M=1 R=2.8
+ SA=75001.5 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1007 N_A_1370_290#_M1007_d N_A_1223_119#_M1007_g N_VGND_M1011_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.425343 PD=0.92 PS=2.18566 NRD=0 NRS=114.288 M=1
+ R=4.26667 SA=75002 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1017 N_A_1790_74#_M1017_d N_A_1025_119#_M1017_g N_A_1370_290#_M1007_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.261434 AS=0.0896 PD=1.85962 PS=0.92 NRD=105.936
+ NRS=0 M=1 R=4.26667 SA=75002.4 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1002 A_2000_74# N_A_852_119#_M1002_g N_A_1790_74#_M1017_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0441 AS=0.171566 PD=0.63 PS=1.22038 NRD=14.28 NRS=15.708 M=1 R=2.8
+ SA=75003.1 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1045 N_VGND_M1045_d N_A_2006_373#_M1045_g A_2000_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.5
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1024 A_2158_74# N_RESET_B_M1024_g N_VGND_M1045_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75003.9
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1016 N_A_2006_373#_M1016_d N_A_1790_74#_M1016_g A_2158_74# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75004.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1025 N_Q_N_M1025_d N_A_1790_74#_M1025_g N_VGND_M1025_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.27675 PD=1.02 PS=2.42 NRD=0 NRS=10.536 M=1 R=4.93333
+ SA=75000.2 SB=75001 A=0.111 P=1.78 MULT=1
MM1037 N_Q_N_M1025_d N_A_1790_74#_M1037_g N_VGND_M1037_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.124942 PD=1.02 PS=1.14217 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1010 N_A_2607_392#_M1010_d N_A_1790_74#_M1010_g N_VGND_M1037_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.108058 PD=1.81 PS=0.987826 NRD=0 NRS=8.436 M=1
+ R=4.26667 SA=75001.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1018 N_Q_M1018_d N_A_2607_392#_M1018_g N_VGND_M1018_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2183 PD=1.02 PS=2.07 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1038 N_Q_M1018_d N_A_2607_392#_M1038_g N_VGND_M1038_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1998 PD=1.02 PS=2.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_VPWR_M1009_d N_SCE_M1009_g N_A_27_79#_M1009_s VPB PSHORT L=0.18 W=0.64
+ AD=0.248 AS=0.1792 PD=1.415 PS=1.84 NRD=13.8491 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90003.1 A=0.1152 P=1.64 MULT=1
MM1039 A_310_464# N_SCE_M1039_g N_VPWR_M1009_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.248 PD=0.88 PS=1.415 NRD=19.9955 NRS=0 M=1 R=3.55556 SA=90001.1
+ SB=90002.1 A=0.1152 P=1.64 MULT=1
MM1006 N_A_388_79#_M1006_d N_D_M1006_g A_310_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.196837 AS=0.0768 PD=1.29 PS=0.88 NRD=41.5473 NRS=19.9955 M=1 R=3.55556
+ SA=90001.6 SB=90001.7 A=0.1152 P=1.64 MULT=1
MM1027 A_541_483# N_A_27_79#_M1027_g N_A_388_79#_M1006_d VPB PSHORT L=0.18
+ W=0.64 AD=0.0768 AS=0.196837 PD=0.88 PS=1.29 NRD=19.9955 NRS=43.0839 M=1
+ R=3.55556 SA=90002 SB=90001.2 A=0.1152 P=1.64 MULT=1
MM1041 N_VPWR_M1041_d N_SCD_M1041_g A_541_483# VPB PSHORT L=0.18 W=0.64
+ AD=0.1184 AS=0.0768 PD=1.01 PS=0.88 NRD=4.6098 NRS=19.9955 M=1 R=3.55556
+ SA=90002.4 SB=90000.8 A=0.1152 P=1.64 MULT=1
MM1035 N_A_388_79#_M1035_d N_RESET_B_M1035_g N_VPWR_M1041_d VPB PSHORT L=0.18
+ W=0.64 AD=0.192 AS=0.1184 PD=1.88 PS=1.01 NRD=4.6098 NRS=23.0687 M=1 R=3.55556
+ SA=90003 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1019 N_VPWR_M1019_d N_CLK_M1019_g N_A_852_119#_M1019_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1036 N_A_1025_119#_M1036_d N_A_852_119#_M1036_g N_VPWR_M1019_d VPB PSHORT
+ L=0.18 W=1.12 AD=0.2912 AS=0.1512 PD=2.76 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1032 N_A_1223_119#_M1032_d N_A_1025_119#_M1032_g N_A_388_79#_M1032_s VPB
+ PSHORT L=0.18 W=0.42 AD=0.0567 AS=0.1113 PD=0.69 PS=1.37 NRD=0 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90001.6 A=0.0756 P=1.2 MULT=1
MM1040 A_1328_457# N_A_852_119#_M1040_g N_A_1223_119#_M1032_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0441 AS=0.0567 PD=0.63 PS=0.69 NRD=23.443 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1020 N_VPWR_M1020_d N_A_1370_290#_M1020_g A_1328_457# VPB PSHORT L=0.18 W=0.42
+ AD=0.121387 AS=0.0441 PD=1.11 PS=0.63 NRD=109.749 NRS=23.443 M=1 R=2.33333
+ SA=90001 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1034 N_A_1223_119#_M1034_d N_RESET_B_M1034_g N_VPWR_M1020_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1113 AS=0.121387 PD=1.37 PS=1.11 NRD=0 NRS=109.749 M=1 R=2.33333
+ SA=90001.6 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1000 N_A_1370_290#_M1000_d N_A_1223_119#_M1000_g N_VPWR_M1000_s VPB PSHORT
+ L=0.18 W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1004 N_A_1790_74#_M1004_d N_A_852_119#_M1004_g N_A_1370_290#_M1000_d VPB
+ PSHORT L=0.18 W=1 AD=0.268732 AS=0.135 PD=2.26761 PS=1.27 NRD=37.4103 NRS=0
+ M=1 R=5.55556 SA=90000.6 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1042 A_1958_471# N_A_1025_119#_M1042_g N_A_1790_74#_M1004_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.112868 PD=0.66 PS=0.952394 NRD=30.4759 NRS=46.886 M=1
+ R=2.33333 SA=90001.3 SB=90003.4 A=0.0756 P=1.2 MULT=1
MM1022 N_VPWR_M1022_d N_A_2006_373#_M1022_g A_1958_471# VPB PSHORT L=0.18 W=0.42
+ AD=0.202162 AS=0.0504 PD=1.32 PS=0.66 NRD=100.844 NRS=30.4759 M=1 R=2.33333
+ SA=90001.7 SB=90003 A=0.0756 P=1.2 MULT=1
MM1023 N_A_2006_373#_M1023_d N_RESET_B_M1023_g N_VPWR_M1022_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0567 AS=0.202162 PD=0.69 PS=1.32 NRD=0 NRS=199.955 M=1 R=2.33333
+ SA=90002.6 SB=90002.1 A=0.0756 P=1.2 MULT=1
MM1028 N_VPWR_M1028_d N_A_1790_74#_M1028_g N_A_2006_373#_M1023_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.0903 AS=0.0567 PD=0.804545 PS=0.69 NRD=105.533 NRS=0 M=1
+ R=2.33333 SA=90003 SB=90001.7 A=0.0756 P=1.2 MULT=1
MM1005 N_Q_N_M1005_d N_A_1790_74#_M1005_g N_VPWR_M1028_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2408 PD=1.39 PS=2.14545 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.4 SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1008 N_Q_N_M1005_d N_A_1790_74#_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.187547 PD=1.39 PS=1.52679 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.9 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1029 N_A_2607_392#_M1029_d N_A_1790_74#_M1029_g N_VPWR_M1008_s VPB PSHORT
+ L=0.18 W=1 AD=0.26 AS=0.167453 PD=2.52 PS=1.36321 NRD=0 NRS=9.8303 M=1
+ R=5.55556 SA=90002.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A_2607_392#_M1001_g N_Q_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1044 N_VPWR_M1044_d N_A_2607_392#_M1044_g N_Q_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3024 AS=0.1512 PD=2.78 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX46_noxref VNB VPB NWDIODE A=28.7103 P=34.48
c_156 VNB 0 1.52826e-19 $X=0 $Y=0
c_2043 A_1958_471# 0 1.02173e-19 $X=9.79 $Y=2.355
*
.include "sky130_fd_sc_ms__sdfrbp_2.pxi.spice"
*
.ends
*
*

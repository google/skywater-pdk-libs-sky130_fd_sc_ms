* NGSPICE file created from sky130_fd_sc_ms__a211o_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 VGND a_81_264# X VNB nlowvt w=740000u l=150000u
+  ad=5.3685e+11p pd=4.68e+06u as=1.961e+11p ps=2.01e+06u
M1001 a_81_264# C1 a_553_392# VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=2.1e+11p ps=2.42e+06u
M1002 a_279_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.3e+11p pd=5.06e+06u as=5.912e+11p ps=5.36e+06u
M1003 VGND B1 a_81_264# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=3.488e+11p ps=3.65e+06u
M1004 a_81_264# C1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_553_392# B1 a_279_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_366_136# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=2.08e+11p pd=1.93e+06u as=0p ps=0u
M1007 VPWR a_81_264# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.912e+11p ps=2.76e+06u
M1008 a_81_264# A1 a_366_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A2 a_279_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__inv_4.spice
* Created: Fri Aug 28 17:38:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__inv_4.pex.spice"
.subckt sky130_fd_sc_ms__inv_4  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_M1002_g N_Y_M1002_s VNB NLOWVT L=0.15 W=0.74 AD=0.2331
+ AS=0.1184 PD=2.11 PS=1.06 NRD=4.86 NRS=6.48 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g N_Y_M1002_s VNB NLOWVT L=0.15 W=0.74 AD=0.1221
+ AS=0.1184 PD=1.07 PS=1.06 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7 SB=75001.1
+ A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1003_d N_A_M1004_g N_Y_M1004_s VNB NLOWVT L=0.15 W=0.74 AD=0.1221
+ AS=0.1036 PD=1.07 PS=1.02 NRD=8.1 NRS=0 M=1 R=4.93333 SA=75001.2 SB=75000.6
+ A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_A_M1005_g N_Y_M1004_s VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2 SB=90001.5
+ A=0.2016 P=2.6 MULT=1
MM1001 N_Y_M1000_d N_A_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6 SB=90001.1
+ A=0.2016 P=2.6 MULT=1
MM1006 N_Y_M1006_d N_A_M1006_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1 SB=90000.6
+ A=0.2016 P=2.6 MULT=1
MM1007 N_Y_M1006_d N_A_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.1708 P=9.28
*
.include "sky130_fd_sc_ms__inv_4.pxi.spice"
*
.ends
*
*

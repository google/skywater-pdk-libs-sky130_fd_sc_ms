* File: sky130_fd_sc_ms__and4_1.spice
* Created: Wed Sep  2 11:58:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__and4_1.pex.spice"
.subckt sky130_fd_sc_ms__and4_1  VNB VPB A B C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1009 A_179_74# N_A_M1009_g N_A_96_74#_M1009_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1696 PD=0.88 PS=1.81 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1007 A_257_74# N_B_M1007_g A_179_74# VNB NLOWVT L=0.15 W=0.64 AD=0.0768
+ AS=0.0768 PD=0.88 PS=0.88 NRD=12.18 NRS=12.18 M=1 R=4.26667 SA=75000.6
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1008 A_335_74# N_C_M1008_g A_257_74# VNB NLOWVT L=0.15 W=0.64 AD=0.1344
+ AS=0.0768 PD=1.06 PS=0.88 NRD=29.052 NRS=12.18 M=1 R=4.26667 SA=75001
+ SB=75001.3 A=0.096 P=1.58 MULT=1
MM1003 N_VGND_M1003_d N_D_M1003_g A_335_74# VNB NLOWVT L=0.15 W=0.64 AD=0.118446
+ AS=0.1344 PD=1.02029 PS=1.06 NRD=0 NRS=29.052 M=1 R=4.26667 SA=75001.5
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1005 N_X_M1005_d N_A_96_74#_M1005_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.136954 PD=2.05 PS=1.17971 NRD=0 NRS=12.972 M=1 R=4.93333
+ SA=75001.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_A_96_74#_M1004_d N_A_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1344 AS=0.2772 PD=1.16 PS=2.34 NRD=0 NRS=10.5395 M=1 R=4.66667 SA=90000.2
+ SB=90002.5 A=0.1512 P=2.04 MULT=1
MM1000 N_VPWR_M1000_d N_B_M1000_g N_A_96_74#_M1004_d VPB PSHORT L=0.18 W=0.84
+ AD=0.2226 AS=0.1344 PD=1.37 PS=1.16 NRD=29.3136 NRS=10.5395 M=1 R=4.66667
+ SA=90000.7 SB=90002 A=0.1512 P=2.04 MULT=1
MM1002 N_A_96_74#_M1002_d N_C_M1002_g N_VPWR_M1000_d VPB PSHORT L=0.18 W=0.84
+ AD=0.1344 AS=0.2226 PD=1.16 PS=1.37 NRD=10.5395 NRS=29.3136 M=1 R=4.66667
+ SA=90001.4 SB=90001.3 A=0.1512 P=2.04 MULT=1
MM1001 N_VPWR_M1001_d N_D_M1001_g N_A_96_74#_M1002_d VPB PSHORT L=0.18 W=0.84
+ AD=0.1758 AS=0.1344 PD=1.30714 PS=1.16 NRD=18.7544 NRS=0 M=1 R=4.66667
+ SA=90001.9 SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1006 N_X_M1006_d N_A_96_74#_M1006_g N_VPWR_M1001_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.2344 PD=2.8 PS=1.74286 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90001.9 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__and4_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__clkinv_1.pex.spice
* Created: Fri Aug 28 17:19:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__CLKINV_1%A 3 7 11 13 14 20 23 27
r33 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.765 $X2=0.59 $Y2=1.765
r34 23 25 50.3829 $w=6.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.72 $Y=1.085
+ $X2=0.72 $Y2=0.92
r35 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.085 $X2=0.59 $Y2=1.085
r36 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.425 $X2=0.59 $Y2=1.425
r37 18 27 12.7388 $w=6.3e-07 $l=4.5873e-08 $layer=POLY_cond $X=0.72 $Y=1.765
+ $X2=0.72 $Y2=1.765
r38 18 20 16.1358 $w=6.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.72 $Y=1.765
+ $X2=0.72 $Y2=1.425
r39 17 23 12.7388 $w=6.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.72 $Y=1.235
+ $X2=0.72 $Y2=1.085
r40 17 20 16.1358 $w=6.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.72 $Y=1.235
+ $X2=0.72 $Y2=1.425
r41 14 28 2.40157 $w=5.08e-07 $l=1e-07 $layer=LI1_cond $X=0.44 $Y=1.665 $X2=0.44
+ $Y2=1.765
r42 14 21 5.76378 $w=5.08e-07 $l=2.4e-07 $layer=LI1_cond $X=0.44 $Y=1.665
+ $X2=0.44 $Y2=1.425
r43 13 21 3.12205 $w=5.08e-07 $l=1.3e-07 $layer=LI1_cond $X=0.44 $Y=1.295
+ $X2=0.44 $Y2=1.425
r44 13 24 5.04331 $w=5.08e-07 $l=2.1e-07 $layer=LI1_cond $X=0.44 $Y=1.295
+ $X2=0.44 $Y2=1.085
r45 9 27 27.1783 $w=3.15e-07 $l=2.96226e-07 $layer=POLY_cond $X=0.945 $Y=1.93
+ $X2=0.72 $Y2=1.765
r46 9 11 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=0.945 $Y=1.93
+ $X2=0.945 $Y2=2.54
r47 7 25 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.565 $Y=0.58
+ $X2=0.565 $Y2=0.92
r48 1 27 27.1783 $w=3.15e-07 $l=2.96226e-07 $layer=POLY_cond $X=0.495 $Y=1.93
+ $X2=0.72 $Y2=1.765
r49 1 3 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.93
+ $X2=0.495 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_MS__CLKINV_1%VPWR 1 2 7 9 11 13 15 17 27
r20 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r21 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r22 18 23 4.02368 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.177 $Y2=3.33
r23 18 20 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.72 $Y2=3.33
r24 17 26 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.222 $Y2=3.33
r25 17 20 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.72 $Y2=3.33
r26 15 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r27 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r28 15 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r29 11 26 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.222 $Y2=3.33
r30 11 13 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=2.79
r31 7 23 3.11948 $w=2.5e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.23 $Y=3.245
+ $X2=0.177 $Y2=3.33
r32 7 9 45.1758 $w=2.48e-07 $l=9.8e-07 $layer=LI1_cond $X=0.23 $Y=3.245 $X2=0.23
+ $Y2=2.265
r33 2 13 600 $w=1.7e-07 $l=7.34405e-07 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=2.12 $X2=1.17 $Y2=2.79
r34 1 9 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.27 $Y2=2.265
.ends

.subckt PM_SKY130_FD_SC_MS__CLKINV_1%Y 1 2 9 11 15 16 17 18 19 26 36 45
r26 40 43 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.695 $Y=2.265
+ $X2=0.72 $Y2=2.265
r27 27 45 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=1.205 $Y=2.1
+ $X2=1.205 $Y2=2.265
r28 27 36 3.1212 $w=2.38e-07 $l=6.5e-08 $layer=LI1_cond $X=1.205 $Y=2.1
+ $X2=1.205 $Y2=2.035
r29 19 45 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.2 $Y=2.265
+ $X2=1.205 $Y2=2.265
r30 19 43 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=2.265
+ $X2=0.72 $Y2=2.265
r31 19 36 0.480185 $w=2.38e-07 $l=1e-08 $layer=LI1_cond $X=1.205 $Y=2.025
+ $X2=1.205 $Y2=2.035
r32 18 19 17.2866 $w=2.38e-07 $l=3.6e-07 $layer=LI1_cond $X=1.205 $Y=1.665
+ $X2=1.205 $Y2=2.025
r33 17 18 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.205 $Y=1.295
+ $X2=1.205 $Y2=1.665
r34 16 17 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.205 $Y=0.925
+ $X2=1.205 $Y2=1.295
r35 16 26 11.7645 $w=2.38e-07 $l=2.45e-07 $layer=LI1_cond $X=1.205 $Y=0.925
+ $X2=1.205 $Y2=0.68
r36 15 26 4.07572 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=1.205 $Y=0.515
+ $X2=1.205 $Y2=0.68
r37 11 15 2.96416 $w=3.3e-07 $l=1.2e-07 $layer=LI1_cond $X=1.085 $Y=0.515
+ $X2=1.205 $Y2=0.515
r38 11 13 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.085 $Y=0.515
+ $X2=0.78 $Y2=0.515
r39 7 40 1.70047 $w=2.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.695 $Y=2.43
+ $X2=0.695 $Y2=2.265
r40 7 9 14.8171 $w=2.78e-07 $l=3.6e-07 $layer=LI1_cond $X=0.695 $Y=2.43
+ $X2=0.695 $Y2=2.79
r41 2 43 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.12 $X2=0.72 $Y2=2.265
r42 2 9 600 $w=1.7e-07 $l=7.34405e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.12 $X2=0.72 $Y2=2.79
r43 1 15 182 $w=1.7e-07 $l=5.88048e-07 $layer=licon1_NDIFF $count=1 $X=0.64
+ $Y=0.37 $X2=1.16 $Y2=0.515
r44 1 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.64
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__CLKINV_1%VGND 1 4 6 8 12 13
r14 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r15 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r16 10 16 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r17 10 12 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=1.2
+ $Y2=0
r18 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r19 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r20 4 16 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r21 4 6 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.28 $Y=0.085 $X2=0.28
+ $Y2=0.55
r22 1 6 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.55
.ends


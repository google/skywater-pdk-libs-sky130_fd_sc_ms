* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__ebufn_1 A TE_B VGND VNB VPB VPWR Z
X0 VGND A a_229_74# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X1 VPWR A a_229_74# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X2 VPWR TE_B a_569_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 a_569_368# a_229_74# Z VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X4 a_27_404# TE_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X5 a_27_404# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X6 a_569_74# a_229_74# Z VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VGND a_27_404# a_569_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

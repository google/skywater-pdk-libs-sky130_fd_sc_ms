* File: sky130_fd_sc_ms__nand4_1.spice
* Created: Fri Aug 28 17:44:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nand4_1.pex.spice"
.subckt sky130_fd_sc_ms__nand4_1  VNB VPB D C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1000 A_181_74# N_D_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.2923 PD=0.98 PS=2.72 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.3 SB=75001.7
+ A=0.111 P=1.78 MULT=1
MM1003 A_259_74# N_C_M1003_g A_181_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.0888 PD=1.16 PS=0.98 NRD=25.128 NRS=10.536 M=1 R=4.93333 SA=75000.7
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1006 A_373_74# N_B_M1006_g A_259_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.1554 PD=1.16 PS=1.16 NRD=25.128 NRS=25.128 M=1 R=4.93333 SA=75001.3
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1007 N_Y_M1007_d N_A_M1007_g A_373_74# VNB NLOWVT L=0.15 W=0.74 AD=0.2085
+ AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=25.128 M=1 R=4.93333 SA=75001.8 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_D_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.2 SB=90001.8
+ A=0.2016 P=2.6 MULT=1
MM1002 N_VPWR_M1002_d N_C_M1002_g N_Y_M1001_d VPB PSHORT L=0.18 W=1.12 AD=0.2408
+ AS=0.1512 PD=1.55 PS=1.39 NRD=12.2928 NRS=0 M=1 R=6.22222 SA=90000.7
+ SB=90001.3 A=0.2016 P=2.6 MULT=1
MM1005 N_Y_M1005_d N_B_M1005_g N_VPWR_M1002_d VPB PSHORT L=0.18 W=1.12 AD=0.1792
+ AS=0.2408 PD=1.44 PS=1.55 NRD=0 NRS=14.0658 M=1 R=6.22222 SA=90001.3
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g N_Y_M1005_d VPB PSHORT L=0.18 W=1.12 AD=0.3136
+ AS=0.1792 PD=2.8 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.8 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ms__nand4_1.pxi.spice"
*
.ends
*
*

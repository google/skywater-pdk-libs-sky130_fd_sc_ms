* File: sky130_fd_sc_ms__sdfrtp_4.pxi.spice
* Created: Fri Aug 28 18:12:28 2020
* 
x_PM_SKY130_FD_SC_MS__SDFRTP_4%A_27_74# N_A_27_74#_M1042_s N_A_27_74#_M1004_s
+ N_A_27_74#_c_294_n N_A_27_74#_c_295_n N_A_27_74#_M1007_g N_A_27_74#_M1024_g
+ N_A_27_74#_c_296_n N_A_27_74#_c_297_n N_A_27_74#_c_303_n N_A_27_74#_c_298_n
+ N_A_27_74#_c_304_n N_A_27_74#_c_299_n N_A_27_74#_c_305_n N_A_27_74#_c_306_n
+ N_A_27_74#_c_307_n N_A_27_74#_c_300_n PM_SKY130_FD_SC_MS__SDFRTP_4%A_27_74#
x_PM_SKY130_FD_SC_MS__SDFRTP_4%SCE N_SCE_M1004_g N_SCE_M1042_g N_SCE_M1039_g
+ N_SCE_c_374_n N_SCE_M1025_g N_SCE_c_376_n N_SCE_c_377_n N_SCE_c_378_n
+ N_SCE_c_379_n SCE SCE SCE N_SCE_c_380_n SCE N_SCE_c_381_n
+ PM_SKY130_FD_SC_MS__SDFRTP_4%SCE
x_PM_SKY130_FD_SC_MS__SDFRTP_4%D N_D_M1008_g N_D_M1021_g D N_D_c_452_n
+ N_D_c_453_n N_D_c_454_n PM_SKY130_FD_SC_MS__SDFRTP_4%D
x_PM_SKY130_FD_SC_MS__SDFRTP_4%SCD N_SCD_M1043_g N_SCD_M1005_g N_SCD_c_494_n
+ N_SCD_c_498_n SCD SCD N_SCD_c_496_n PM_SKY130_FD_SC_MS__SDFRTP_4%SCD
x_PM_SKY130_FD_SC_MS__SDFRTP_4%CLK N_CLK_c_534_n N_CLK_M1038_g N_CLK_M1026_g CLK
+ PM_SKY130_FD_SC_MS__SDFRTP_4%CLK
x_PM_SKY130_FD_SC_MS__SDFRTP_4%A_1037_387# N_A_1037_387#_M1041_d
+ N_A_1037_387#_M1040_d N_A_1037_387#_M1016_g N_A_1037_387#_c_587_n
+ N_A_1037_387#_M1017_g N_A_1037_387#_c_589_n N_A_1037_387#_M1006_g
+ N_A_1037_387#_c_590_n N_A_1037_387#_c_591_n N_A_1037_387#_M1014_g
+ N_A_1037_387#_c_592_n N_A_1037_387#_c_593_n N_A_1037_387#_c_594_n
+ N_A_1037_387#_c_595_n N_A_1037_387#_c_596_n N_A_1037_387#_c_597_n
+ N_A_1037_387#_c_598_n N_A_1037_387#_c_651_p N_A_1037_387#_c_599_n
+ N_A_1037_387#_c_600_n N_A_1037_387#_c_601_n N_A_1037_387#_c_602_n
+ N_A_1037_387#_c_637_p N_A_1037_387#_c_614_n N_A_1037_387#_c_615_n
+ N_A_1037_387#_c_603_n N_A_1037_387#_c_604_n N_A_1037_387#_c_605_n
+ N_A_1037_387#_c_606_n N_A_1037_387#_c_607_n
+ PM_SKY130_FD_SC_MS__SDFRTP_4%A_1037_387#
x_PM_SKY130_FD_SC_MS__SDFRTP_4%A_1367_112# N_A_1367_112#_M1028_d
+ N_A_1367_112#_M1018_d N_A_1367_112#_M1000_g N_A_1367_112#_M1002_g
+ N_A_1367_112#_c_814_n N_A_1367_112#_c_815_n N_A_1367_112#_c_831_n
+ N_A_1367_112#_c_816_n N_A_1367_112#_c_817_n N_A_1367_112#_c_822_n
+ N_A_1367_112#_c_843_n N_A_1367_112#_c_845_n
+ PM_SKY130_FD_SC_MS__SDFRTP_4%A_1367_112#
x_PM_SKY130_FD_SC_MS__SDFRTP_4%RESET_B N_RESET_B_M1013_g N_RESET_B_M1035_g
+ N_RESET_B_c_917_n N_RESET_B_c_918_n N_RESET_B_c_925_n N_RESET_B_c_926_n
+ N_RESET_B_M1034_g N_RESET_B_c_920_n N_RESET_B_c_921_n N_RESET_B_c_922_n
+ N_RESET_B_M1003_g N_RESET_B_M1045_g N_RESET_B_M1031_g N_RESET_B_c_931_n
+ N_RESET_B_c_932_n N_RESET_B_c_933_n N_RESET_B_c_934_n N_RESET_B_c_935_n
+ N_RESET_B_c_936_n RESET_B N_RESET_B_c_938_n N_RESET_B_c_939_n
+ N_RESET_B_c_940_n N_RESET_B_c_941_n PM_SKY130_FD_SC_MS__SDFRTP_4%RESET_B
x_PM_SKY130_FD_SC_MS__SDFRTP_4%A_1233_138# N_A_1233_138#_M1027_d
+ N_A_1233_138#_M1016_d N_A_1233_138#_M1003_d N_A_1233_138#_M1028_g
+ N_A_1233_138#_c_1132_n N_A_1233_138#_M1018_g N_A_1233_138#_c_1141_n
+ N_A_1233_138#_c_1154_n N_A_1233_138#_c_1133_n N_A_1233_138#_c_1177_n
+ N_A_1233_138#_c_1134_n N_A_1233_138#_c_1135_n N_A_1233_138#_c_1136_n
+ N_A_1233_138#_c_1137_n N_A_1233_138#_c_1138_n N_A_1233_138#_c_1145_n
+ PM_SKY130_FD_SC_MS__SDFRTP_4%A_1233_138#
x_PM_SKY130_FD_SC_MS__SDFRTP_4%A_834_93# N_A_834_93#_M1038_s N_A_834_93#_M1026_s
+ N_A_834_93#_M1040_g N_A_834_93#_M1041_g N_A_834_93#_c_1261_n
+ N_A_834_93#_c_1262_n N_A_834_93#_c_1263_n N_A_834_93#_c_1276_n
+ N_A_834_93#_c_1277_n N_A_834_93#_c_1264_n N_A_834_93#_c_1265_n
+ N_A_834_93#_M1027_g N_A_834_93#_M1012_g N_A_834_93#_c_1279_n
+ N_A_834_93#_M1022_g N_A_834_93#_c_1266_n N_A_834_93#_c_1267_n
+ N_A_834_93#_M1036_g N_A_834_93#_c_1283_n N_A_834_93#_c_1289_n
+ N_A_834_93#_c_1290_n N_A_834_93#_c_1292_n N_A_834_93#_c_1269_n
+ N_A_834_93#_c_1284_n N_A_834_93#_c_1270_n N_A_834_93#_c_1299_n
+ N_A_834_93#_c_1271_n N_A_834_93#_c_1272_n N_A_834_93#_c_1273_n
+ PM_SKY130_FD_SC_MS__SDFRTP_4%A_834_93#
x_PM_SKY130_FD_SC_MS__SDFRTP_4%A_2003_48# N_A_2003_48#_M1030_d
+ N_A_2003_48#_M1031_d N_A_2003_48#_M1032_g N_A_2003_48#_M1010_g
+ N_A_2003_48#_c_1452_n N_A_2003_48#_c_1453_n N_A_2003_48#_c_1454_n
+ N_A_2003_48#_c_1455_n N_A_2003_48#_c_1456_n N_A_2003_48#_c_1460_n
+ N_A_2003_48#_c_1457_n N_A_2003_48#_c_1458_n
+ PM_SKY130_FD_SC_MS__SDFRTP_4%A_2003_48#
x_PM_SKY130_FD_SC_MS__SDFRTP_4%A_1745_74# N_A_1745_74#_M1006_d
+ N_A_1745_74#_M1022_d N_A_1745_74#_c_1535_n N_A_1745_74#_M1030_g
+ N_A_1745_74#_c_1536_n N_A_1745_74#_M1044_g N_A_1745_74#_c_1537_n
+ N_A_1745_74#_c_1552_n N_A_1745_74#_M1001_g N_A_1745_74#_c_1538_n
+ N_A_1745_74#_M1011_g N_A_1745_74#_c_1539_n N_A_1745_74#_c_1540_n
+ N_A_1745_74#_c_1554_n N_A_1745_74#_M1046_g N_A_1745_74#_c_1541_n
+ N_A_1745_74#_c_1542_n N_A_1745_74#_c_1543_n N_A_1745_74#_c_1567_n
+ N_A_1745_74#_c_1556_n N_A_1745_74#_c_1544_n N_A_1745_74#_c_1545_n
+ N_A_1745_74#_c_1546_n N_A_1745_74#_c_1558_n N_A_1745_74#_c_1559_n
+ N_A_1745_74#_c_1560_n N_A_1745_74#_c_1547_n N_A_1745_74#_c_1548_n
+ N_A_1745_74#_c_1549_n PM_SKY130_FD_SC_MS__SDFRTP_4%A_1745_74#
x_PM_SKY130_FD_SC_MS__SDFRTP_4%A_2339_74# N_A_2339_74#_M1011_s
+ N_A_2339_74#_M1001_s N_A_2339_74#_c_1693_n N_A_2339_74#_M1009_g
+ N_A_2339_74#_c_1694_n N_A_2339_74#_c_1695_n N_A_2339_74#_c_1696_n
+ N_A_2339_74#_M1020_g N_A_2339_74#_M1015_g N_A_2339_74#_M1019_g
+ N_A_2339_74#_M1023_g N_A_2339_74#_c_1700_n N_A_2339_74#_M1033_g
+ N_A_2339_74#_M1029_g N_A_2339_74#_c_1702_n N_A_2339_74#_M1037_g
+ N_A_2339_74#_c_1703_n N_A_2339_74#_c_1704_n N_A_2339_74#_c_1705_n
+ N_A_2339_74#_c_1706_n N_A_2339_74#_c_1707_n
+ PM_SKY130_FD_SC_MS__SDFRTP_4%A_2339_74#
x_PM_SKY130_FD_SC_MS__SDFRTP_4%VPWR N_VPWR_M1004_d N_VPWR_M1043_d N_VPWR_M1026_d
+ N_VPWR_M1002_d N_VPWR_M1018_s N_VPWR_M1010_d N_VPWR_M1044_d N_VPWR_M1046_d
+ N_VPWR_M1019_s N_VPWR_M1029_s N_VPWR_c_1814_n N_VPWR_c_1815_n N_VPWR_c_1816_n
+ N_VPWR_c_1817_n N_VPWR_c_1818_n N_VPWR_c_1819_n N_VPWR_c_1820_n
+ N_VPWR_c_1821_n N_VPWR_c_1822_n N_VPWR_c_1823_n N_VPWR_c_1824_n
+ N_VPWR_c_1825_n N_VPWR_c_1826_n N_VPWR_c_1827_n N_VPWR_c_1828_n
+ N_VPWR_c_1829_n VPWR N_VPWR_c_1830_n N_VPWR_c_1831_n N_VPWR_c_1832_n
+ N_VPWR_c_1833_n N_VPWR_c_1834_n N_VPWR_c_1835_n N_VPWR_c_1836_n
+ N_VPWR_c_1837_n N_VPWR_c_1838_n N_VPWR_c_1839_n N_VPWR_c_1840_n
+ N_VPWR_c_1841_n N_VPWR_c_1842_n N_VPWR_c_1813_n
+ PM_SKY130_FD_SC_MS__SDFRTP_4%VPWR
x_PM_SKY130_FD_SC_MS__SDFRTP_4%A_415_81# N_A_415_81#_M1008_d N_A_415_81#_M1027_s
+ N_A_415_81#_M1021_d N_A_415_81#_M1035_d N_A_415_81#_M1016_s
+ N_A_415_81#_c_2019_n N_A_415_81#_c_2004_n N_A_415_81#_c_2005_n
+ N_A_415_81#_c_2012_n N_A_415_81#_c_2006_n N_A_415_81#_c_2013_n
+ N_A_415_81#_c_2007_n N_A_415_81#_c_2008_n N_A_415_81#_c_2014_n
+ N_A_415_81#_c_2015_n N_A_415_81#_c_2009_n N_A_415_81#_c_2017_n
+ N_A_415_81#_c_2010_n N_A_415_81#_c_2018_n
+ PM_SKY130_FD_SC_MS__SDFRTP_4%A_415_81#
x_PM_SKY130_FD_SC_MS__SDFRTP_4%Q N_Q_M1009_s N_Q_M1033_s N_Q_M1015_d N_Q_M1023_d
+ N_Q_c_2150_n N_Q_c_2161_n N_Q_c_2165_n N_Q_c_2154_n N_Q_c_2155_n N_Q_c_2156_n
+ N_Q_c_2157_n N_Q_c_2151_n N_Q_c_2152_n Q PM_SKY130_FD_SC_MS__SDFRTP_4%Q
x_PM_SKY130_FD_SC_MS__SDFRTP_4%VGND N_VGND_M1042_d N_VGND_M1013_d N_VGND_M1038_d
+ N_VGND_M1034_d N_VGND_M1032_d N_VGND_M1011_d N_VGND_M1020_d N_VGND_M1037_d
+ N_VGND_c_2218_n N_VGND_c_2219_n N_VGND_c_2220_n N_VGND_c_2221_n
+ N_VGND_c_2222_n N_VGND_c_2223_n N_VGND_c_2224_n N_VGND_c_2225_n
+ N_VGND_c_2226_n N_VGND_c_2227_n N_VGND_c_2228_n VGND N_VGND_c_2229_n
+ N_VGND_c_2230_n N_VGND_c_2231_n N_VGND_c_2232_n N_VGND_c_2233_n
+ N_VGND_c_2234_n N_VGND_c_2235_n N_VGND_c_2236_n N_VGND_c_2237_n
+ N_VGND_c_2238_n N_VGND_c_2239_n N_VGND_c_2240_n
+ PM_SKY130_FD_SC_MS__SDFRTP_4%VGND
x_PM_SKY130_FD_SC_MS__SDFRTP_4%noxref_24 N_noxref_24_M1007_s N_noxref_24_M1005_d
+ N_noxref_24_c_2363_n N_noxref_24_c_2364_n N_noxref_24_c_2365_n
+ PM_SKY130_FD_SC_MS__SDFRTP_4%noxref_24
cc_1 VNB N_A_27_74#_c_294_n 0.0258189f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_2 VNB N_A_27_74#_c_295_n 0.0213547f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.935
cc_3 VNB N_A_27_74#_c_296_n 0.0257773f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_4 VNB N_A_27_74#_c_297_n 0.0190417f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.005
cc_5 VNB N_A_27_74#_c_298_n 0.00987534f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_6 VNB N_A_27_74#_c_299_n 0.018224f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_7 VNB N_A_27_74#_c_300_n 0.0395906f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.01
cc_8 VNB N_SCE_M1042_g 0.0668709f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_9 VNB N_SCE_c_374_n 0.0481513f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.64
cc_10 VNB N_SCE_M1025_g 0.0214295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_SCE_c_376_n 0.00775502f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_12 VNB N_SCE_c_377_n 0.0420954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_SCE_c_378_n 0.0133027f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.265
cc_14 VNB N_SCE_c_379_n 0.00565867f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.465
cc_15 VNB N_SCE_c_380_n 0.0106235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_SCE_c_381_n 0.00168276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_D_M1021_g 0.0274525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_D_c_452_n 0.0376278f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_19 VNB N_D_c_453_n 0.00724067f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.16
cc_20 VNB N_D_c_454_n 0.0170107f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.64
cc_21 VNB N_SCD_M1005_g 0.0409572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_SCD_c_494_n 0.00372888f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_23 VNB SCD 0.00358506f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.16
cc_24 VNB N_SCD_c_496_n 0.0156486f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_25 VNB N_CLK_c_534_n 0.0847518f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=0.37
cc_26 VNB CLK 0.0181649f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.01
cc_27 VNB N_A_1037_387#_c_587_n 0.00940815f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.615
cc_28 VNB N_A_1037_387#_M1017_g 0.0358586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_1037_387#_c_589_n 0.0168538f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_30 VNB N_A_1037_387#_c_590_n 0.0237434f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.265
cc_31 VNB N_A_1037_387#_c_591_n 0.00657402f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.005
cc_32 VNB N_A_1037_387#_c_592_n 0.00949995f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_33 VNB N_A_1037_387#_c_593_n 6.4492e-19 $X=-0.19 $Y=-0.245 $X2=2.375 $Y2=2.09
cc_34 VNB N_A_1037_387#_c_594_n 0.037314f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=2.09
cc_35 VNB N_A_1037_387#_c_595_n 0.00479168f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_36 VNB N_A_1037_387#_c_596_n 4.85147e-19 $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.09
cc_37 VNB N_A_1037_387#_c_597_n 0.00173551f $X=-0.19 $Y=-0.245 $X2=2.53
+ $Y2=1.995
cc_38 VNB N_A_1037_387#_c_598_n 0.00102705f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=2.09
cc_39 VNB N_A_1037_387#_c_599_n 0.00657839f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_40 VNB N_A_1037_387#_c_600_n 0.00209509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_1037_387#_c_601_n 0.00144678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1037_387#_c_602_n 0.005194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1037_387#_c_603_n 0.00108143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1037_387#_c_604_n 0.00756725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1037_387#_c_605_n 0.0332641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_1037_387#_c_606_n 0.00593212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1037_387#_c_607_n 0.00976988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1367_112#_M1000_g 0.035113f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.935
cc_49 VNB N_A_1367_112#_c_814_n 0.00471142f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_50 VNB N_A_1367_112#_c_815_n 0.014438f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_51 VNB N_A_1367_112#_c_816_n 0.00556937f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.465
cc_52 VNB N_A_1367_112#_c_817_n 0.00450848f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.465
cc_53 VNB N_RESET_B_M1013_g 0.052812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_RESET_B_c_917_n 0.267629f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.01
cc_55 VNB N_RESET_B_c_918_n 0.012806f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.935
cc_56 VNB N_RESET_B_M1034_g 0.0336923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_RESET_B_c_920_n 0.0235284f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.935
cc_58 VNB N_RESET_B_c_921_n 0.00691999f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_59 VNB N_RESET_B_c_922_n 0.0186961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_RESET_B_M1045_g 0.0569134f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.1
cc_61 VNB N_A_1233_138#_M1028_g 0.0225417f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.16
cc_62 VNB N_A_1233_138#_c_1132_n 0.0164104f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.64
cc_63 VNB N_A_1233_138#_c_1133_n 0.00369363f $X=-0.19 $Y=-0.245 $X2=0.975
+ $Y2=1.1
cc_64 VNB N_A_1233_138#_c_1134_n 5.47792e-19 $X=-0.19 $Y=-0.245 $X2=2.375
+ $Y2=2.09
cc_65 VNB N_A_1233_138#_c_1135_n 0.00176601f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=2.09
cc_66 VNB N_A_1233_138#_c_1136_n 0.00526285f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.09
cc_67 VNB N_A_1233_138#_c_1137_n 0.0281158f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_68 VNB N_A_1233_138#_c_1138_n 0.00176618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_834_93#_c_1261_n 0.0166468f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.64
cc_70 VNB N_A_834_93#_c_1262_n 0.0243897f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.935
cc_71 VNB N_A_834_93#_c_1263_n 0.00295443f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_72 VNB N_A_834_93#_c_1264_n 0.0277159f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.265
cc_73 VNB N_A_834_93#_c_1265_n 0.0172456f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.175
cc_74 VNB N_A_834_93#_c_1266_n 0.0193702f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=1.995
cc_75 VNB N_A_834_93#_c_1267_n 0.00478428f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=1.995
cc_76 VNB N_A_834_93#_M1036_g 0.0510568f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=2.09
cc_77 VNB N_A_834_93#_c_1269_n 0.00169001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_834_93#_c_1270_n 0.00323883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_834_93#_c_1271_n 0.00181774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_834_93#_c_1272_n 0.0194018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_834_93#_c_1273_n 0.0154198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_2003_48#_M1032_g 0.0340019f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.935
cc_83 VNB N_A_2003_48#_M1010_g 0.0060931f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.64
cc_84 VNB N_A_2003_48#_c_1452_n 0.0178026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_2003_48#_c_1453_n 0.00567377f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_86 VNB N_A_2003_48#_c_1454_n 0.00480935f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.465
cc_87 VNB N_A_2003_48#_c_1455_n 0.00289977f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.1
cc_88 VNB N_A_2003_48#_c_1456_n 0.031198f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_89 VNB N_A_2003_48#_c_1457_n 0.00270148f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_90 VNB N_A_2003_48#_c_1458_n 0.00662489f $X=-0.19 $Y=-0.245 $X2=2.53
+ $Y2=1.995
cc_91 VNB N_A_1745_74#_c_1535_n 0.021255f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_92 VNB N_A_1745_74#_c_1536_n 0.00668157f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.16
cc_93 VNB N_A_1745_74#_c_1537_n 0.0250522f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.935
cc_94 VNB N_A_1745_74#_c_1538_n 0.0185474f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.005
cc_95 VNB N_A_1745_74#_c_1539_n 0.0159493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1745_74#_c_1540_n 0.0140662f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.1
cc_97 VNB N_A_1745_74#_c_1541_n 0.0143997f $X=-0.19 $Y=-0.245 $X2=2.375 $Y2=2.09
cc_98 VNB N_A_1745_74#_c_1542_n 0.00257119f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=2.09
cc_99 VNB N_A_1745_74#_c_1543_n 0.00496366f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_100 VNB N_A_1745_74#_c_1544_n 0.00146437f $X=-0.19 $Y=-0.245 $X2=0.975
+ $Y2=1.1
cc_101 VNB N_A_1745_74#_c_1545_n 0.00359384f $X=-0.19 $Y=-0.245 $X2=2.53
+ $Y2=1.995
cc_102 VNB N_A_1745_74#_c_1546_n 0.0291774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1745_74#_c_1547_n 0.00123798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1745_74#_c_1548_n 0.00179963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1745_74#_c_1549_n 0.0646681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_2339_74#_c_1693_n 0.0177259f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_107 VNB N_A_2339_74#_c_1694_n 0.0142247f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.615
cc_108 VNB N_A_2339_74#_c_1695_n 0.00638412f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.615
cc_109 VNB N_A_2339_74#_c_1696_n 0.021315f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.16
cc_110 VNB N_A_2339_74#_M1015_g 0.00352464f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_111 VNB N_A_2339_74#_M1019_g 0.00313742f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.005
cc_112 VNB N_A_2339_74#_M1023_g 0.00312223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_2339_74#_c_1700_n 0.0221017f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_114 VNB N_A_2339_74#_M1029_g 0.003575f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=2.09
cc_115 VNB N_A_2339_74#_c_1702_n 0.0216728f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.09
cc_116 VNB N_A_2339_74#_c_1703_n 0.00311192f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=2.09
cc_117 VNB N_A_2339_74#_c_1704_n 0.00104691f $X=-0.19 $Y=-0.245 $X2=0.975
+ $Y2=1.1
cc_118 VNB N_A_2339_74#_c_1705_n 0.00999107f $X=-0.19 $Y=-0.245 $X2=2.53
+ $Y2=1.995
cc_119 VNB N_A_2339_74#_c_1706_n 0.00570341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_2339_74#_c_1707_n 0.11445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VPWR_c_1813_n 0.621437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_415_81#_c_2004_n 0.0200812f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.265
cc_123 VNB N_A_415_81#_c_2005_n 0.00510274f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.465
cc_124 VNB N_A_415_81#_c_2006_n 0.00334006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_415_81#_c_2007_n 0.00530091f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.09
cc_126 VNB N_A_415_81#_c_2008_n 0.00155689f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_127 VNB N_A_415_81#_c_2009_n 0.00251617f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=2.09
cc_128 VNB N_A_415_81#_c_2010_n 0.00503812f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_129 VNB N_Q_c_2150_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_Q_c_2151_n 0.00178889f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=1.995
cc_131 VNB N_Q_c_2152_n 0.00200996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB Q 0.0195094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2218_n 0.0110567f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_134 VNB N_VGND_c_2219_n 0.0124691f $X=-0.19 $Y=-0.245 $X2=2.375 $Y2=2.09
cc_135 VNB N_VGND_c_2220_n 0.0146422f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=1.995
cc_136 VNB N_VGND_c_2221_n 0.00428891f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=2.09
cc_137 VNB N_VGND_c_2222_n 0.00497485f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_138 VNB N_VGND_c_2223_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=1.995
cc_139 VNB N_VGND_c_2224_n 0.0413125f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=2.16
cc_140 VNB N_VGND_c_2225_n 0.0646059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2226_n 0.00399507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2227_n 0.0198576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2228_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2229_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2230_n 0.0577219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2231_n 0.0602754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2232_n 0.0428668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2233_n 0.0151727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2234_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2235_n 0.0142666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2236_n 0.00808418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2237_n 0.00481148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2238_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2239_n 0.0272142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2240_n 0.76539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_noxref_24_c_2363_n 0.0135787f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_157 VNB N_noxref_24_c_2364_n 0.00655627f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.935
cc_158 VNB N_noxref_24_c_2365_n 0.00264023f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.64
cc_159 VPB N_A_27_74#_M1024_g 0.0231566f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.64
cc_160 VPB N_A_27_74#_c_297_n 0.016494f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.005
cc_161 VPB N_A_27_74#_c_303_n 0.0337004f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_162 VPB N_A_27_74#_c_304_n 0.0349952f $X=-0.19 $Y=1.66 $X2=2.375 $Y2=2.09
cc_163 VPB N_A_27_74#_c_305_n 0.0129728f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_164 VPB N_A_27_74#_c_306_n 0.00593531f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.995
cc_165 VPB N_A_27_74#_c_307_n 0.0278636f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.995
cc_166 VPB N_SCE_M1004_g 0.0591491f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_SCE_M1039_g 0.0511293f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_168 VPB N_SCE_c_376_n 0.00782879f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_169 VPB N_SCE_c_377_n 0.0410982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_SCE_c_379_n 0.00298426f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_171 VPB N_SCE_c_381_n 0.00270951f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_D_M1021_g 0.0522201f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_SCD_c_494_n 0.032149f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_174 VPB N_SCD_c_498_n 0.0333828f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_175 VPB SCD 0.00339002f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.16
cc_176 VPB N_CLK_c_534_n 0.0171168f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=0.37
cc_177 VPB N_CLK_M1026_g 0.0260261f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB CLK 0.00168095f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=1.01
cc_179 VPB N_A_1037_387#_M1016_g 0.0346011f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.935
cc_180 VPB N_A_1037_387#_c_587_n 0.0139705f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_181 VPB N_A_1037_387#_M1014_g 0.0245981f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_182 VPB N_A_1037_387#_c_596_n 0.0027361f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_183 VPB N_A_1037_387#_c_597_n 0.00201099f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.995
cc_184 VPB N_A_1037_387#_c_602_n 0.00112302f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_1037_387#_c_614_n 0.00501177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_1037_387#_c_615_n 0.0331884f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_1037_387#_c_607_n 0.0200155f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_1367_112#_M1002_g 0.0350694f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.64
cc_189 VPB N_A_1367_112#_c_814_n 0.00199812f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.58
cc_190 VPB N_A_1367_112#_c_815_n 0.0359063f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_191 VPB N_A_1367_112#_c_817_n 7.08723e-19 $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_192 VPB N_A_1367_112#_c_822_n 0.00313252f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_193 VPB N_RESET_B_M1013_g 0.00651144f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_RESET_B_c_925_n 0.0391944f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_195 VPB N_RESET_B_c_926_n 0.0258864f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_196 VPB N_RESET_B_c_922_n 0.010912f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_RESET_B_M1003_g 0.024019f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.175
cc_198 VPB N_RESET_B_M1045_g 0.00996849f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_199 VPB N_RESET_B_M1031_g 0.0406275f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_RESET_B_c_931_n 0.021365f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_201 VPB N_RESET_B_c_932_n 0.0204556f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=1.995
cc_202 VPB N_RESET_B_c_933_n 0.00174228f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.995
cc_203 VPB N_RESET_B_c_934_n 0.0213442f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.995
cc_204 VPB N_RESET_B_c_935_n 0.00238517f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_RESET_B_c_936_n 0.00203191f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.995
cc_206 VPB RESET_B 0.00336207f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_RESET_B_c_938_n 0.00300368f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_RESET_B_c_939_n 0.054615f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_RESET_B_c_940_n 0.00478311f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_RESET_B_c_941_n 0.0461414f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_1233_138#_c_1132_n 0.00954671f $X=-0.19 $Y=1.66 $X2=2.495
+ $Y2=2.64
cc_212 VPB N_A_1233_138#_M1018_g 0.0217885f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_213 VPB N_A_1233_138#_c_1141_n 0.00303721f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.265
cc_214 VPB N_A_1233_138#_c_1133_n 0.00622911f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_215 VPB N_A_1233_138#_c_1134_n 0.0120245f $X=-0.19 $Y=1.66 $X2=2.375 $Y2=2.09
cc_216 VPB N_A_1233_138#_c_1137_n 0.00783535f $X=-0.19 $Y=1.66 $X2=2.54
+ $Y2=1.995
cc_217 VPB N_A_1233_138#_c_1145_n 0.00179594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_834_93#_M1040_g 0.0212731f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.935
cc_219 VPB N_A_834_93#_c_1263_n 0.0781447f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.58
cc_220 VPB N_A_834_93#_c_1276_n 0.0582987f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_221 VPB N_A_834_93#_c_1277_n 0.0106868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_834_93#_M1012_g 0.0391803f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_223 VPB N_A_834_93#_c_1279_n 0.185027f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_224 VPB N_A_834_93#_M1022_g 0.027891f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_225 VPB N_A_834_93#_c_1266_n 0.0188847f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=1.995
cc_226 VPB N_A_834_93#_c_1267_n 0.00334601f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.995
cc_227 VPB N_A_834_93#_c_1283_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_228 VPB N_A_834_93#_c_1284_n 0.00283353f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_834_93#_c_1271_n 0.00241584f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_834_93#_c_1272_n 0.0103893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_2003_48#_M1010_g 0.0649017f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.64
cc_232 VPB N_A_2003_48#_c_1460_n 0.00804843f $X=-0.19 $Y=1.66 $X2=0.445 $Y2=2.09
cc_233 VPB N_A_2003_48#_c_1457_n 0.0184686f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.1
cc_234 VPB N_A_1745_74#_c_1536_n 3.48694e-19 $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.16
cc_235 VPB N_A_1745_74#_M1044_g 0.0693498f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.64
cc_236 VPB N_A_1745_74#_c_1552_n 0.0169346f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_237 VPB N_A_1745_74#_c_1540_n 0.00996836f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_238 VPB N_A_1745_74#_c_1554_n 0.0169548f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_239 VPB N_A_1745_74#_c_1542_n 0.00426118f $X=-0.19 $Y=1.66 $X2=0.445 $Y2=2.09
cc_240 VPB N_A_1745_74#_c_1556_n 0.00176039f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_A_1745_74#_c_1545_n 0.00118387f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.995
cc_242 VPB N_A_1745_74#_c_1558_n 0.0080022f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_1745_74#_c_1559_n 0.00236595f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_A_1745_74#_c_1560_n 0.00699846f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_2339_74#_M1015_g 0.0237135f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.58
cc_246 VPB N_A_2339_74#_M1019_g 0.0217889f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.005
cc_247 VPB N_A_2339_74#_M1023_g 0.0211609f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_A_2339_74#_M1029_g 0.024499f $X=-0.19 $Y=1.66 $X2=0.445 $Y2=2.09
cc_249 VPB N_A_2339_74#_c_1704_n 0.0035517f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_250 VPB N_VPWR_c_1814_n 0.00611419f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.1
cc_251 VPB N_VPWR_c_1815_n 0.00151893f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.995
cc_252 VPB N_VPWR_c_1816_n 0.0138296f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.01
cc_253 VPB N_VPWR_c_1817_n 0.0230775f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_254 VPB N_VPWR_c_1818_n 0.0142406f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=2.16
cc_255 VPB N_VPWR_c_1819_n 0.01372f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1820_n 0.0277625f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1821_n 0.0213687f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1822_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1823_n 0.00492117f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1824_n 0.0115177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1825_n 0.0443855f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1826_n 0.0328326f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1827_n 0.00485379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1828_n 0.0520927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1829_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1830_n 0.0191816f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1831_n 0.0457766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1832_n 0.0586031f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1833_n 0.0245819f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1834_n 0.0218508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1835_n 0.0173155f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1836_n 0.031111f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1837_n 0.00655093f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1838_n 0.00463502f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1839_n 0.00223798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1840_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1841_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1842_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_1813_n 0.126958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_A_415_81#_c_2005_n 0.00473919f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_281 VPB N_A_415_81#_c_2012_n 0.0113046f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_282 VPB N_A_415_81#_c_2013_n 5.29111e-19 $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.1
cc_283 VPB N_A_415_81#_c_2014_n 0.00625148f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.995
cc_284 VPB N_A_415_81#_c_2015_n 0.00190509f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.995
cc_285 VPB N_A_415_81#_c_2009_n 0.00578945f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=2.09
cc_286 VPB N_A_415_81#_c_2017_n 0.00231322f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.01
cc_287 VPB N_A_415_81#_c_2018_n 0.0113014f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_288 VPB N_Q_c_2154_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.005
cc_289 VPB N_Q_c_2155_n 0.00293927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_290 VPB N_Q_c_2156_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_291 VPB N_Q_c_2157_n 0.00221223f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_292 VPB Q 0.0137493f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_293 N_A_27_74#_c_303_n N_SCE_M1004_g 0.0184741f $X=0.28 $Y=2.465 $X2=0 $Y2=0
cc_294 N_A_27_74#_c_304_n N_SCE_M1004_g 0.0195433f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_295 N_A_27_74#_c_305_n N_SCE_M1004_g 0.00544367f $X=0.28 $Y=2.09 $X2=0 $Y2=0
cc_296 N_A_27_74#_c_296_n N_SCE_M1042_g 0.00686809f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_297 N_A_27_74#_c_297_n N_SCE_M1042_g 0.00830473f $X=0.2 $Y=2.005 $X2=0 $Y2=0
cc_298 N_A_27_74#_c_298_n N_SCE_M1042_g 0.0281157f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_299 N_A_27_74#_c_300_n N_SCE_M1042_g 0.0181297f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_300 N_A_27_74#_c_304_n N_SCE_M1039_g 0.018168f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_301 N_A_27_74#_c_306_n N_SCE_c_374_n 3.50012e-19 $X=2.53 $Y=1.995 $X2=0 $Y2=0
cc_302 N_A_27_74#_c_307_n N_SCE_c_374_n 0.0181978f $X=2.53 $Y=1.995 $X2=0 $Y2=0
cc_303 N_A_27_74#_c_297_n N_SCE_c_376_n 0.0158921f $X=0.2 $Y=2.005 $X2=0 $Y2=0
cc_304 N_A_27_74#_c_298_n N_SCE_c_376_n 0.00162366f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_305 N_A_27_74#_c_294_n N_SCE_c_377_n 0.0106974f $X=1.41 $Y=1.01 $X2=0 $Y2=0
cc_306 N_A_27_74#_c_298_n N_SCE_c_377_n 0.00180358f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_307 N_A_27_74#_c_304_n N_SCE_c_377_n 0.0170396f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_308 N_A_27_74#_c_300_n N_SCE_c_377_n 0.0175645f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_309 N_A_27_74#_c_304_n N_SCE_c_378_n 0.0253169f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_310 N_A_27_74#_c_306_n N_SCE_c_378_n 0.00219771f $X=2.53 $Y=1.995 $X2=0 $Y2=0
cc_311 N_A_27_74#_c_306_n N_SCE_c_379_n 0.0242979f $X=2.53 $Y=1.995 $X2=0 $Y2=0
cc_312 N_A_27_74#_c_307_n N_SCE_c_379_n 0.00100601f $X=2.53 $Y=1.995 $X2=0 $Y2=0
cc_313 N_A_27_74#_c_294_n N_SCE_c_380_n 0.00818136f $X=1.41 $Y=1.01 $X2=0 $Y2=0
cc_314 N_A_27_74#_c_297_n N_SCE_c_380_n 0.0170838f $X=0.2 $Y=2.005 $X2=0 $Y2=0
cc_315 N_A_27_74#_c_298_n N_SCE_c_380_n 0.0353374f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_316 N_A_27_74#_c_304_n N_SCE_c_380_n 0.0893268f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_317 N_A_27_74#_c_300_n N_SCE_c_380_n 0.00202099f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_318 N_A_27_74#_M1024_g N_D_M1021_g 0.0153877f $X=2.495 $Y=2.64 $X2=0 $Y2=0
cc_319 N_A_27_74#_c_304_n N_D_M1021_g 0.0168703f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_320 N_A_27_74#_c_306_n N_D_M1021_g 0.00124829f $X=2.53 $Y=1.995 $X2=0 $Y2=0
cc_321 N_A_27_74#_c_307_n N_D_M1021_g 0.0193155f $X=2.53 $Y=1.995 $X2=0 $Y2=0
cc_322 N_A_27_74#_c_294_n N_D_c_452_n 0.00979811f $X=1.41 $Y=1.01 $X2=0 $Y2=0
cc_323 N_A_27_74#_c_298_n N_D_c_452_n 2.46751e-19 $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_324 N_A_27_74#_c_300_n N_D_c_452_n 0.00223479f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_325 N_A_27_74#_c_295_n N_D_c_453_n 0.00580814f $X=1.485 $Y=0.935 $X2=0 $Y2=0
cc_326 N_A_27_74#_c_298_n N_D_c_453_n 0.0143876f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_327 N_A_27_74#_c_300_n N_D_c_453_n 8.79717e-19 $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_328 N_A_27_74#_c_295_n N_D_c_454_n 0.0224455f $X=1.485 $Y=0.935 $X2=0 $Y2=0
cc_329 N_A_27_74#_c_306_n N_SCD_c_494_n 0.00256419f $X=2.53 $Y=1.995 $X2=0 $Y2=0
cc_330 N_A_27_74#_c_307_n N_SCD_c_494_n 0.0206967f $X=2.53 $Y=1.995 $X2=0 $Y2=0
cc_331 N_A_27_74#_M1024_g N_SCD_c_498_n 0.0312525f $X=2.495 $Y=2.64 $X2=0 $Y2=0
cc_332 N_A_27_74#_c_306_n SCD 0.0195527f $X=2.53 $Y=1.995 $X2=0 $Y2=0
cc_333 N_A_27_74#_c_307_n SCD 3.7256e-19 $X=2.53 $Y=1.995 $X2=0 $Y2=0
cc_334 N_A_27_74#_M1024_g N_VPWR_c_1814_n 0.00145742f $X=2.495 $Y=2.64 $X2=0
+ $Y2=0
cc_335 N_A_27_74#_c_303_n N_VPWR_c_1830_n 0.014549f $X=0.28 $Y=2.465 $X2=0 $Y2=0
cc_336 N_A_27_74#_M1024_g N_VPWR_c_1831_n 0.005209f $X=2.495 $Y=2.64 $X2=0 $Y2=0
cc_337 N_A_27_74#_c_303_n N_VPWR_c_1836_n 0.0247088f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_338 N_A_27_74#_c_304_n N_VPWR_c_1836_n 0.0739847f $X=2.375 $Y=2.09 $X2=0
+ $Y2=0
cc_339 N_A_27_74#_M1024_g N_VPWR_c_1813_n 0.00528953f $X=2.495 $Y=2.64 $X2=0
+ $Y2=0
cc_340 N_A_27_74#_c_303_n N_VPWR_c_1813_n 0.0119743f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_341 N_A_27_74#_M1024_g N_A_415_81#_c_2019_n 0.010236f $X=2.495 $Y=2.64 $X2=0
+ $Y2=0
cc_342 N_A_27_74#_c_306_n N_A_415_81#_c_2019_n 0.018047f $X=2.53 $Y=1.995 $X2=0
+ $Y2=0
cc_343 N_A_27_74#_c_307_n N_A_415_81#_c_2019_n 6.21636e-19 $X=2.53 $Y=1.995
+ $X2=0 $Y2=0
cc_344 N_A_27_74#_M1024_g N_A_415_81#_c_2017_n 0.0110942f $X=2.495 $Y=2.64 $X2=0
+ $Y2=0
cc_345 N_A_27_74#_c_304_n N_A_415_81#_c_2017_n 0.0182356f $X=2.375 $Y=2.09 $X2=0
+ $Y2=0
cc_346 N_A_27_74#_c_306_n N_A_415_81#_c_2017_n 0.00358719f $X=2.53 $Y=1.995
+ $X2=0 $Y2=0
cc_347 N_A_27_74#_c_295_n N_VGND_c_2218_n 0.00287309f $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_348 N_A_27_74#_c_296_n N_VGND_c_2218_n 0.0156021f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_349 N_A_27_74#_c_298_n N_VGND_c_2218_n 0.0254818f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_350 N_A_27_74#_c_300_n N_VGND_c_2218_n 0.00149092f $X=0.975 $Y=1.01 $X2=0
+ $Y2=0
cc_351 N_A_27_74#_c_295_n N_VGND_c_2225_n 9.09582e-19 $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_352 N_A_27_74#_c_296_n N_VGND_c_2229_n 0.011066f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_353 N_A_27_74#_c_296_n N_VGND_c_2240_n 0.00915947f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_354 N_A_27_74#_c_295_n N_noxref_24_c_2363_n 0.011495f $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_355 N_A_27_74#_c_295_n N_noxref_24_c_2364_n 0.00899724f $X=1.485 $Y=0.935
+ $X2=0 $Y2=0
cc_356 N_A_27_74#_c_298_n N_noxref_24_c_2364_n 0.00178881f $X=0.975 $Y=1.1 $X2=0
+ $Y2=0
cc_357 N_A_27_74#_c_300_n N_noxref_24_c_2364_n 0.00859402f $X=0.975 $Y=1.01
+ $X2=0 $Y2=0
cc_358 N_SCE_c_377_n N_D_M1021_g 0.0847159f $X=1.535 $Y=1.67 $X2=0 $Y2=0
cc_359 N_SCE_c_378_n N_D_M1021_g 0.0144881f $X=2.405 $Y=1.575 $X2=0 $Y2=0
cc_360 N_SCE_c_379_n N_D_M1021_g 3.12323e-19 $X=2.53 $Y=1.425 $X2=0 $Y2=0
cc_361 N_SCE_c_381_n N_D_M1021_g 0.00479409f $X=1.795 $Y=1.662 $X2=0 $Y2=0
cc_362 N_SCE_c_374_n N_D_c_452_n 0.0261857f $X=2.7 $Y=1.05 $X2=0 $Y2=0
cc_363 N_SCE_M1025_g N_D_c_452_n 0.00235321f $X=2.7 $Y=0.615 $X2=0 $Y2=0
cc_364 N_SCE_c_379_n N_D_c_452_n 0.00139763f $X=2.53 $Y=1.425 $X2=0 $Y2=0
cc_365 N_SCE_c_381_n N_D_c_452_n 0.00411836f $X=1.795 $Y=1.662 $X2=0 $Y2=0
cc_366 N_SCE_c_374_n N_D_c_453_n 0.001089f $X=2.7 $Y=1.05 $X2=0 $Y2=0
cc_367 N_SCE_M1025_g N_D_c_453_n 5.59487e-19 $X=2.7 $Y=0.615 $X2=0 $Y2=0
cc_368 N_SCE_c_377_n N_D_c_453_n 0.00106377f $X=1.535 $Y=1.67 $X2=0 $Y2=0
cc_369 N_SCE_c_380_n N_D_c_453_n 0.0344941f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_370 N_SCE_M1025_g N_D_c_454_n 0.00891111f $X=2.7 $Y=0.615 $X2=0 $Y2=0
cc_371 N_SCE_c_374_n N_SCD_M1005_g 0.0100532f $X=2.7 $Y=1.05 $X2=0 $Y2=0
cc_372 N_SCE_M1025_g N_SCD_M1005_g 0.0572711f $X=2.7 $Y=0.615 $X2=0 $Y2=0
cc_373 N_SCE_c_379_n N_SCD_M1005_g 0.00386588f $X=2.53 $Y=1.425 $X2=0 $Y2=0
cc_374 N_SCE_c_379_n SCD 0.0148328f $X=2.53 $Y=1.425 $X2=0 $Y2=0
cc_375 N_SCE_c_374_n N_SCD_c_496_n 0.00937702f $X=2.7 $Y=1.05 $X2=0 $Y2=0
cc_376 N_SCE_c_379_n N_SCD_c_496_n 0.00253998f $X=2.53 $Y=1.425 $X2=0 $Y2=0
cc_377 N_SCE_M1004_g N_VPWR_c_1830_n 0.005209f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_378 N_SCE_M1039_g N_VPWR_c_1831_n 0.00461464f $X=1.625 $Y=2.64 $X2=0 $Y2=0
cc_379 N_SCE_M1004_g N_VPWR_c_1836_n 0.00585939f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_380 N_SCE_M1039_g N_VPWR_c_1836_n 0.0181112f $X=1.625 $Y=2.64 $X2=0 $Y2=0
cc_381 N_SCE_M1004_g N_VPWR_c_1813_n 0.00990469f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_382 N_SCE_M1039_g N_VPWR_c_1813_n 0.00908371f $X=1.625 $Y=2.64 $X2=0 $Y2=0
cc_383 N_SCE_c_374_n N_A_415_81#_c_2004_n 0.00197359f $X=2.7 $Y=1.05 $X2=0 $Y2=0
cc_384 N_SCE_M1025_g N_A_415_81#_c_2004_n 0.00257713f $X=2.7 $Y=0.615 $X2=0
+ $Y2=0
cc_385 N_SCE_M1039_g N_A_415_81#_c_2017_n 0.00179756f $X=1.625 $Y=2.64 $X2=0
+ $Y2=0
cc_386 N_SCE_c_374_n N_A_415_81#_c_2010_n 0.00682628f $X=2.7 $Y=1.05 $X2=0 $Y2=0
cc_387 N_SCE_M1025_g N_A_415_81#_c_2010_n 0.0122867f $X=2.7 $Y=0.615 $X2=0 $Y2=0
cc_388 N_SCE_c_378_n N_A_415_81#_c_2010_n 0.00245612f $X=2.405 $Y=1.575 $X2=0
+ $Y2=0
cc_389 N_SCE_c_379_n N_A_415_81#_c_2010_n 0.0200193f $X=2.53 $Y=1.425 $X2=0
+ $Y2=0
cc_390 N_SCE_M1042_g N_VGND_c_2218_n 0.0129468f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_391 N_SCE_M1025_g N_VGND_c_2225_n 9.15902e-19 $X=2.7 $Y=0.615 $X2=0 $Y2=0
cc_392 N_SCE_M1042_g N_VGND_c_2229_n 0.00383152f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_393 N_SCE_M1042_g N_VGND_c_2240_n 0.00761198f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_394 N_SCE_M1025_g N_noxref_24_c_2363_n 0.0108161f $X=2.7 $Y=0.615 $X2=0 $Y2=0
cc_395 N_SCE_M1042_g N_noxref_24_c_2364_n 9.19966e-19 $X=0.495 $Y=0.58 $X2=0
+ $Y2=0
cc_396 N_D_M1021_g N_VPWR_c_1831_n 0.005209f $X=2.045 $Y=2.64 $X2=0 $Y2=0
cc_397 N_D_M1021_g N_VPWR_c_1836_n 0.00232995f $X=2.045 $Y=2.64 $X2=0 $Y2=0
cc_398 N_D_M1021_g N_VPWR_c_1813_n 0.00983291f $X=2.045 $Y=2.64 $X2=0 $Y2=0
cc_399 N_D_M1021_g N_A_415_81#_c_2017_n 0.0126578f $X=2.045 $Y=2.64 $X2=0 $Y2=0
cc_400 N_D_c_452_n N_A_415_81#_c_2010_n 0.00118317f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_401 N_D_c_453_n N_A_415_81#_c_2010_n 0.0118953f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_402 N_D_c_454_n N_A_415_81#_c_2010_n 0.00586479f $X=1.952 $Y=0.935 $X2=0
+ $Y2=0
cc_403 N_D_c_454_n N_VGND_c_2225_n 9.15902e-19 $X=1.952 $Y=0.935 $X2=0 $Y2=0
cc_404 N_D_c_452_n N_noxref_24_c_2363_n 0.00121903f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_405 N_D_c_453_n N_noxref_24_c_2363_n 0.014028f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_406 N_D_c_454_n N_noxref_24_c_2363_n 0.0123477f $X=1.952 $Y=0.935 $X2=0 $Y2=0
cc_407 N_D_c_454_n N_noxref_24_c_2364_n 0.00108287f $X=1.952 $Y=0.935 $X2=0
+ $Y2=0
cc_408 N_D_c_453_n noxref_25 0.00395662f $X=1.935 $Y=1.1 $X2=-0.19 $Y2=-0.245
cc_409 N_SCD_M1005_g N_RESET_B_M1013_g 0.0296618f $X=3.06 $Y=0.615 $X2=0 $Y2=0
cc_410 SCD N_RESET_B_M1013_g 0.00226841f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_411 N_SCD_c_496_n N_RESET_B_M1013_g 0.0232039f $X=3.07 $Y=1.605 $X2=0 $Y2=0
cc_412 N_SCD_c_494_n N_RESET_B_c_926_n 0.0232039f $X=3.07 $Y=2.08 $X2=0 $Y2=0
cc_413 N_SCD_c_498_n N_RESET_B_c_931_n 0.0183524f $X=3.07 $Y=2.245 $X2=0 $Y2=0
cc_414 N_SCD_c_498_n N_VPWR_c_1814_n 0.0123606f $X=3.07 $Y=2.245 $X2=0 $Y2=0
cc_415 N_SCD_c_498_n N_VPWR_c_1831_n 0.00398535f $X=3.07 $Y=2.245 $X2=0 $Y2=0
cc_416 N_SCD_c_498_n N_VPWR_c_1813_n 0.0039465f $X=3.07 $Y=2.245 $X2=0 $Y2=0
cc_417 N_SCD_c_498_n N_A_415_81#_c_2019_n 0.0181987f $X=3.07 $Y=2.245 $X2=0
+ $Y2=0
cc_418 SCD N_A_415_81#_c_2019_n 0.020493f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_419 N_SCD_M1005_g N_A_415_81#_c_2004_n 0.0128507f $X=3.06 $Y=0.615 $X2=0
+ $Y2=0
cc_420 SCD N_A_415_81#_c_2004_n 0.0148869f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_421 N_SCD_c_496_n N_A_415_81#_c_2004_n 0.0022356f $X=3.07 $Y=1.605 $X2=0
+ $Y2=0
cc_422 N_SCD_M1005_g N_A_415_81#_c_2005_n 0.00624809f $X=3.06 $Y=0.615 $X2=0
+ $Y2=0
cc_423 N_SCD_c_498_n N_A_415_81#_c_2005_n 0.0037275f $X=3.07 $Y=2.245 $X2=0
+ $Y2=0
cc_424 SCD N_A_415_81#_c_2005_n 0.0562728f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_425 N_SCD_c_496_n N_A_415_81#_c_2005_n 0.00192445f $X=3.07 $Y=1.605 $X2=0
+ $Y2=0
cc_426 N_SCD_c_498_n N_A_415_81#_c_2017_n 0.00169232f $X=3.07 $Y=2.245 $X2=0
+ $Y2=0
cc_427 N_SCD_M1005_g N_A_415_81#_c_2010_n 0.00152614f $X=3.06 $Y=0.615 $X2=0
+ $Y2=0
cc_428 N_SCD_c_498_n N_A_415_81#_c_2018_n 4.73014e-19 $X=3.07 $Y=2.245 $X2=0
+ $Y2=0
cc_429 N_SCD_M1005_g N_VGND_c_2225_n 9.15902e-19 $X=3.06 $Y=0.615 $X2=0 $Y2=0
cc_430 N_SCD_M1005_g N_noxref_24_c_2363_n 0.00977032f $X=3.06 $Y=0.615 $X2=0
+ $Y2=0
cc_431 N_SCD_M1005_g N_noxref_24_c_2365_n 8.58945e-19 $X=3.06 $Y=0.615 $X2=0
+ $Y2=0
cc_432 N_CLK_c_534_n N_A_1037_387#_c_592_n 6.88559e-19 $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_433 N_CLK_M1026_g N_A_1037_387#_c_596_n 4.98055e-19 $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_434 N_CLK_c_534_n N_RESET_B_M1013_g 0.0215051f $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_435 CLK N_RESET_B_M1013_g 0.00739527f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_436 N_CLK_c_534_n N_RESET_B_c_917_n 0.0100723f $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_437 CLK N_RESET_B_c_917_n 0.0053784f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_438 N_CLK_c_534_n N_RESET_B_c_925_n 0.0169757f $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_439 N_CLK_M1026_g N_RESET_B_c_925_n 0.00513254f $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_440 CLK N_RESET_B_c_925_n 0.0026948f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_441 N_CLK_c_534_n N_RESET_B_c_932_n 5.9655e-19 $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_442 CLK N_RESET_B_c_932_n 0.00697481f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_443 N_CLK_M1026_g N_RESET_B_c_933_n 3.38591e-19 $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_444 CLK N_RESET_B_c_933_n 0.00449924f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_445 N_CLK_c_534_n N_RESET_B_c_938_n 6.89102e-19 $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_446 N_CLK_M1026_g N_RESET_B_c_938_n 9.54548e-19 $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_447 CLK N_RESET_B_c_938_n 0.0306648f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_448 CLK N_A_834_93#_M1038_s 0.00635712f $X=3.995 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_449 N_CLK_M1026_g N_A_834_93#_M1040_g 0.0488079f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_450 N_CLK_c_534_n N_A_834_93#_c_1289_n 0.00635441f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_451 N_CLK_c_534_n N_A_834_93#_c_1290_n 0.0113122f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_452 CLK N_A_834_93#_c_1290_n 0.00778119f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_453 N_CLK_c_534_n N_A_834_93#_c_1292_n 0.00409648f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_454 CLK N_A_834_93#_c_1292_n 0.0241453f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_455 N_CLK_c_534_n N_A_834_93#_c_1269_n 0.00342876f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_456 CLK N_A_834_93#_c_1269_n 0.0201012f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_457 N_CLK_M1026_g N_A_834_93#_c_1284_n 0.00211906f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_458 N_CLK_c_534_n N_A_834_93#_c_1270_n 0.00885609f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_459 CLK N_A_834_93#_c_1270_n 0.0113164f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_460 N_CLK_c_534_n N_A_834_93#_c_1299_n 0.00148522f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_461 N_CLK_M1026_g N_A_834_93#_c_1299_n 0.0165761f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_462 CLK N_A_834_93#_c_1299_n 0.0198685f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_463 N_CLK_c_534_n N_A_834_93#_c_1271_n 0.00334124f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_464 CLK N_A_834_93#_c_1271_n 0.0279371f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_465 N_CLK_c_534_n N_A_834_93#_c_1272_n 0.0198175f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_466 CLK N_A_834_93#_c_1272_n 2.931e-19 $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_467 N_CLK_c_534_n N_A_834_93#_c_1273_n 0.0210807f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_468 N_CLK_M1026_g N_VPWR_c_1815_n 0.017461f $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_469 N_CLK_M1026_g N_VPWR_c_1826_n 0.00401239f $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_470 N_CLK_M1026_g N_VPWR_c_1813_n 0.00589267f $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_471 CLK N_A_415_81#_c_2004_n 0.0145731f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_472 N_CLK_c_534_n N_A_415_81#_c_2005_n 0.00106344f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_473 CLK N_A_415_81#_c_2005_n 0.045375f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_474 N_CLK_M1026_g N_A_415_81#_c_2012_n 0.0159379f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_475 N_CLK_M1026_g N_A_415_81#_c_2018_n 0.0144989f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_476 N_CLK_c_534_n N_VGND_c_2219_n 0.0021241f $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_477 CLK N_VGND_c_2219_n 0.0142261f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_478 N_CLK_c_534_n N_VGND_c_2220_n 0.0028517f $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_479 N_CLK_c_534_n N_VGND_c_2240_n 9.39239e-19 $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_480 N_A_1037_387#_c_599_n N_A_1367_112#_M1028_d 0.00224844f $X=8.825 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_481 N_A_1037_387#_M1017_g N_A_1367_112#_M1000_g 0.030435f $X=6.52 $Y=0.9
+ $X2=0 $Y2=0
cc_482 N_A_1037_387#_c_594_n N_A_1367_112#_M1000_g 0.00321205f $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_483 N_A_1037_387#_c_604_n N_A_1367_112#_M1000_g 0.00342215f $X=7.14 $Y=0.415
+ $X2=0 $Y2=0
cc_484 N_A_1037_387#_M1016_g N_A_1367_112#_M1002_g 0.00285501f $X=6.135 $Y=2.525
+ $X2=0 $Y2=0
cc_485 N_A_1037_387#_M1016_g N_A_1367_112#_c_815_n 3.5795e-19 $X=6.135 $Y=2.525
+ $X2=0 $Y2=0
cc_486 N_A_1037_387#_c_587_n N_A_1367_112#_c_815_n 0.030435f $X=6.445 $Y=1.66
+ $X2=0 $Y2=0
cc_487 N_A_1037_387#_c_607_n N_A_1367_112#_c_815_n 0.0023084f $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_488 N_A_1037_387#_c_598_n N_A_1367_112#_c_831_n 0.00761753f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_489 N_A_1037_387#_c_604_n N_A_1367_112#_c_831_n 0.00974988f $X=7.14 $Y=0.415
+ $X2=0 $Y2=0
cc_490 N_A_1037_387#_c_591_n N_A_1367_112#_c_816_n 0.00476106f $X=8.725 $Y=1.16
+ $X2=0 $Y2=0
cc_491 N_A_1037_387#_c_602_n N_A_1367_112#_c_816_n 0.00539231f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_492 N_A_1037_387#_c_606_n N_A_1367_112#_c_816_n 0.0108396f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_493 N_A_1037_387#_c_591_n N_A_1367_112#_c_817_n 0.00855892f $X=8.725 $Y=1.16
+ $X2=0 $Y2=0
cc_494 N_A_1037_387#_c_602_n N_A_1367_112#_c_817_n 0.0129187f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_495 N_A_1037_387#_c_606_n N_A_1367_112#_c_817_n 0.0180376f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_496 N_A_1037_387#_M1014_g N_A_1367_112#_c_822_n 8.42394e-19 $X=9.835 $Y=2.75
+ $X2=0 $Y2=0
cc_497 N_A_1037_387#_c_602_n N_A_1367_112#_c_822_n 0.0240786f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_498 N_A_1037_387#_c_637_p N_A_1367_112#_c_822_n 0.0118335f $X=9.415 $Y=2.222
+ $X2=0 $Y2=0
cc_499 N_A_1037_387#_c_615_n N_A_1367_112#_c_822_n 2.16541e-19 $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_500 N_A_1037_387#_c_598_n N_A_1367_112#_c_843_n 0.0484504f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_501 N_A_1037_387#_c_599_n N_A_1367_112#_c_843_n 0.00422751f $X=8.825 $Y=0.34
+ $X2=0 $Y2=0
cc_502 N_A_1037_387#_c_589_n N_A_1367_112#_c_845_n 0.00932475f $X=8.65 $Y=1.085
+ $X2=0 $Y2=0
cc_503 N_A_1037_387#_c_591_n N_A_1367_112#_c_845_n 2.66567e-19 $X=8.725 $Y=1.16
+ $X2=0 $Y2=0
cc_504 N_A_1037_387#_c_599_n N_A_1367_112#_c_845_n 0.02112f $X=8.825 $Y=0.34
+ $X2=0 $Y2=0
cc_505 N_A_1037_387#_c_601_n N_A_1367_112#_c_845_n 0.0232075f $X=8.91 $Y=0.905
+ $X2=0 $Y2=0
cc_506 N_A_1037_387#_c_606_n N_A_1367_112#_c_845_n 0.0158476f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_507 N_A_1037_387#_M1017_g N_RESET_B_c_917_n 0.00526413f $X=6.52 $Y=0.9 $X2=0
+ $Y2=0
cc_508 N_A_1037_387#_c_594_n N_RESET_B_c_917_n 0.0257323f $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_509 N_A_1037_387#_c_595_n N_RESET_B_c_917_n 0.00969117f $X=5.62 $Y=0.415
+ $X2=0 $Y2=0
cc_510 N_A_1037_387#_c_604_n N_RESET_B_c_917_n 0.00184232f $X=7.14 $Y=0.415
+ $X2=0 $Y2=0
cc_511 N_A_1037_387#_c_598_n N_RESET_B_M1034_g 0.0116325f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_512 N_A_1037_387#_c_651_p N_RESET_B_M1034_g 0.0035287f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_513 N_A_1037_387#_c_600_n N_RESET_B_M1034_g 6.46496e-19 $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_514 N_A_1037_387#_c_604_n N_RESET_B_M1034_g 0.0104865f $X=7.14 $Y=0.415 $X2=0
+ $Y2=0
cc_515 N_A_1037_387#_M1040_d N_RESET_B_c_932_n 0.00355841f $X=5.185 $Y=1.935
+ $X2=0 $Y2=0
cc_516 N_A_1037_387#_M1016_g N_RESET_B_c_932_n 0.00393395f $X=6.135 $Y=2.525
+ $X2=0 $Y2=0
cc_517 N_A_1037_387#_c_587_n N_RESET_B_c_932_n 0.00374625f $X=6.445 $Y=1.66
+ $X2=0 $Y2=0
cc_518 N_A_1037_387#_c_596_n N_RESET_B_c_932_n 0.030298f $X=5.655 $Y=1.75 $X2=0
+ $Y2=0
cc_519 N_A_1037_387#_c_597_n N_RESET_B_c_932_n 0.016446f $X=6.065 $Y=1.75 $X2=0
+ $Y2=0
cc_520 N_A_1037_387#_c_607_n N_RESET_B_c_932_n 0.00388711f $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_521 N_A_1037_387#_c_602_n N_RESET_B_c_934_n 0.0104861f $X=9.33 $Y=2.065 $X2=0
+ $Y2=0
cc_522 N_A_1037_387#_c_637_p N_RESET_B_c_934_n 0.00467739f $X=9.415 $Y=2.222
+ $X2=0 $Y2=0
cc_523 N_A_1037_387#_c_614_n N_RESET_B_c_934_n 0.0172592f $X=9.79 $Y=2.215 $X2=0
+ $Y2=0
cc_524 N_A_1037_387#_c_615_n N_RESET_B_c_934_n 0.00245602f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_525 N_A_1037_387#_c_589_n N_A_1233_138#_M1028_g 0.0216734f $X=8.65 $Y=1.085
+ $X2=0 $Y2=0
cc_526 N_A_1037_387#_c_598_n N_A_1233_138#_M1028_g 0.00459622f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_527 N_A_1037_387#_c_599_n N_A_1233_138#_M1028_g 0.00898149f $X=8.825 $Y=0.34
+ $X2=0 $Y2=0
cc_528 N_A_1037_387#_c_600_n N_A_1233_138#_M1028_g 0.00298755f $X=8.1 $Y=0.34
+ $X2=0 $Y2=0
cc_529 N_A_1037_387#_c_591_n N_A_1233_138#_c_1132_n 0.0122034f $X=8.725 $Y=1.16
+ $X2=0 $Y2=0
cc_530 N_A_1037_387#_c_602_n N_A_1233_138#_c_1132_n 3.24172e-19 $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_531 N_A_1037_387#_M1016_g N_A_1233_138#_c_1141_n 6.00433e-19 $X=6.135
+ $Y=2.525 $X2=0 $Y2=0
cc_532 N_A_1037_387#_c_587_n N_A_1233_138#_c_1141_n 7.27569e-19 $X=6.445 $Y=1.66
+ $X2=0 $Y2=0
cc_533 N_A_1037_387#_M1017_g N_A_1233_138#_c_1154_n 0.0095662f $X=6.52 $Y=0.9
+ $X2=0 $Y2=0
cc_534 N_A_1037_387#_c_594_n N_A_1233_138#_c_1154_n 0.0143871f $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_535 N_A_1037_387#_M1016_g N_A_1233_138#_c_1133_n 5.84645e-19 $X=6.135
+ $Y=2.525 $X2=0 $Y2=0
cc_536 N_A_1037_387#_M1017_g N_A_1233_138#_c_1133_n 0.00659846f $X=6.52 $Y=0.9
+ $X2=0 $Y2=0
cc_537 N_A_1037_387#_c_587_n N_A_1233_138#_c_1138_n 4.04338e-19 $X=6.445 $Y=1.66
+ $X2=0 $Y2=0
cc_538 N_A_1037_387#_M1017_g N_A_1233_138#_c_1138_n 0.00592263f $X=6.52 $Y=0.9
+ $X2=0 $Y2=0
cc_539 N_A_1037_387#_c_594_n N_A_1233_138#_c_1138_n 0.0250786f $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_540 N_A_1037_387#_c_604_n N_A_1233_138#_c_1138_n 0.00225536f $X=7.14 $Y=0.415
+ $X2=0 $Y2=0
cc_541 N_A_1037_387#_M1016_g N_A_1233_138#_c_1145_n 2.41348e-19 $X=6.135
+ $Y=2.525 $X2=0 $Y2=0
cc_542 N_A_1037_387#_c_596_n N_A_834_93#_M1040_g 0.00606819f $X=5.655 $Y=1.75
+ $X2=0 $Y2=0
cc_543 N_A_1037_387#_c_593_n N_A_834_93#_c_1261_n 0.00625478f $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_544 N_A_1037_387#_c_596_n N_A_834_93#_c_1261_n 0.00587978f $X=5.655 $Y=1.75
+ $X2=0 $Y2=0
cc_545 N_A_1037_387#_c_593_n N_A_834_93#_c_1262_n 0.0114875f $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_546 N_A_1037_387#_c_596_n N_A_834_93#_c_1262_n 0.00177607f $X=5.655 $Y=1.75
+ $X2=0 $Y2=0
cc_547 N_A_1037_387#_c_597_n N_A_834_93#_c_1262_n 0.00264594f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_548 N_A_1037_387#_c_603_n N_A_834_93#_c_1262_n 0.00329714f $X=5.412 $Y=1.275
+ $X2=0 $Y2=0
cc_549 N_A_1037_387#_c_607_n N_A_834_93#_c_1262_n 0.0213581f $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_550 N_A_1037_387#_M1016_g N_A_834_93#_c_1263_n 0.0248664f $X=6.135 $Y=2.525
+ $X2=0 $Y2=0
cc_551 N_A_1037_387#_c_596_n N_A_834_93#_c_1263_n 0.0195374f $X=5.655 $Y=1.75
+ $X2=0 $Y2=0
cc_552 N_A_1037_387#_c_597_n N_A_834_93#_c_1263_n 0.00465901f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_553 N_A_1037_387#_M1016_g N_A_834_93#_c_1276_n 0.0123638f $X=6.135 $Y=2.525
+ $X2=0 $Y2=0
cc_554 N_A_1037_387#_c_597_n N_A_834_93#_c_1264_n 0.00369435f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_555 N_A_1037_387#_c_607_n N_A_834_93#_c_1264_n 0.0169891f $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_556 N_A_1037_387#_M1017_g N_A_834_93#_c_1265_n 0.0201381f $X=6.52 $Y=0.9
+ $X2=0 $Y2=0
cc_557 N_A_1037_387#_c_592_n N_A_834_93#_c_1265_n 0.00428521f $X=5.355 $Y=0.74
+ $X2=0 $Y2=0
cc_558 N_A_1037_387#_c_594_n N_A_834_93#_c_1265_n 0.00349197f $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_559 N_A_1037_387#_M1016_g N_A_834_93#_M1012_g 0.0134907f $X=6.135 $Y=2.525
+ $X2=0 $Y2=0
cc_560 N_A_1037_387#_c_587_n N_A_834_93#_M1012_g 0.00158155f $X=6.445 $Y=1.66
+ $X2=0 $Y2=0
cc_561 N_A_1037_387#_M1014_g N_A_834_93#_M1022_g 0.0153622f $X=9.835 $Y=2.75
+ $X2=0 $Y2=0
cc_562 N_A_1037_387#_c_602_n N_A_834_93#_M1022_g 0.0081799f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_563 N_A_1037_387#_c_637_p N_A_834_93#_M1022_g 0.00204696f $X=9.415 $Y=2.222
+ $X2=0 $Y2=0
cc_564 N_A_1037_387#_c_615_n N_A_834_93#_M1022_g 0.00816612f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_565 N_A_1037_387#_c_602_n N_A_834_93#_c_1266_n 0.0123734f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_566 N_A_1037_387#_c_614_n N_A_834_93#_c_1266_n 0.00422095f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_567 N_A_1037_387#_c_615_n N_A_834_93#_c_1266_n 0.00483559f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_568 N_A_1037_387#_c_605_n N_A_834_93#_c_1266_n 0.00926704f $X=9.25 $Y=1.07
+ $X2=0 $Y2=0
cc_569 N_A_1037_387#_c_590_n N_A_834_93#_c_1267_n 0.00926704f $X=9.085 $Y=1.16
+ $X2=0 $Y2=0
cc_570 N_A_1037_387#_c_606_n N_A_834_93#_c_1267_n 0.0013375f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_571 N_A_1037_387#_c_599_n N_A_834_93#_M1036_g 0.0039082f $X=8.825 $Y=0.34
+ $X2=0 $Y2=0
cc_572 N_A_1037_387#_c_601_n N_A_834_93#_M1036_g 0.00172497f $X=8.91 $Y=0.905
+ $X2=0 $Y2=0
cc_573 N_A_1037_387#_c_602_n N_A_834_93#_M1036_g 0.00175577f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_574 N_A_1037_387#_c_605_n N_A_834_93#_M1036_g 0.0213739f $X=9.25 $Y=1.07
+ $X2=0 $Y2=0
cc_575 N_A_1037_387#_c_606_n N_A_834_93#_M1036_g 3.81838e-19 $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_576 N_A_1037_387#_c_592_n N_A_834_93#_c_1289_n 0.00391727f $X=5.355 $Y=0.74
+ $X2=0 $Y2=0
cc_577 N_A_1037_387#_c_593_n N_A_834_93#_c_1269_n 0.00520535f $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_578 N_A_1037_387#_c_596_n N_A_834_93#_c_1284_n 0.00567735f $X=5.655 $Y=1.75
+ $X2=0 $Y2=0
cc_579 N_A_1037_387#_c_596_n N_A_834_93#_c_1299_n 0.0127334f $X=5.655 $Y=1.75
+ $X2=0 $Y2=0
cc_580 N_A_1037_387#_c_593_n N_A_834_93#_c_1271_n 0.0102343f $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_581 N_A_1037_387#_c_596_n N_A_834_93#_c_1271_n 0.0261924f $X=5.655 $Y=1.75
+ $X2=0 $Y2=0
cc_582 N_A_1037_387#_c_603_n N_A_834_93#_c_1271_n 0.00350345f $X=5.412 $Y=1.275
+ $X2=0 $Y2=0
cc_583 N_A_1037_387#_c_596_n N_A_834_93#_c_1272_n 0.00261646f $X=5.655 $Y=1.75
+ $X2=0 $Y2=0
cc_584 N_A_1037_387#_c_603_n N_A_834_93#_c_1272_n 0.0087648f $X=5.412 $Y=1.275
+ $X2=0 $Y2=0
cc_585 N_A_1037_387#_c_592_n N_A_834_93#_c_1273_n 0.00916871f $X=5.355 $Y=0.74
+ $X2=0 $Y2=0
cc_586 N_A_1037_387#_c_593_n N_A_834_93#_c_1273_n 9.57894e-19 $X=5.535 $Y=1.585
+ $X2=0 $Y2=0
cc_587 N_A_1037_387#_c_595_n N_A_834_93#_c_1273_n 0.00126334f $X=5.62 $Y=0.415
+ $X2=0 $Y2=0
cc_588 N_A_1037_387#_c_603_n N_A_834_93#_c_1273_n 0.00224086f $X=5.412 $Y=1.275
+ $X2=0 $Y2=0
cc_589 N_A_1037_387#_M1014_g N_A_2003_48#_M1010_g 0.0385164f $X=9.835 $Y=2.75
+ $X2=0 $Y2=0
cc_590 N_A_1037_387#_c_614_n N_A_2003_48#_M1010_g 3.87491e-19 $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_591 N_A_1037_387#_c_615_n N_A_2003_48#_M1010_g 0.0213989f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_592 N_A_1037_387#_c_599_n N_A_1745_74#_M1006_d 0.00191611f $X=8.825 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_593 N_A_1037_387#_c_601_n N_A_1745_74#_M1006_d 0.0113939f $X=8.91 $Y=0.905
+ $X2=-0.19 $Y2=-0.245
cc_594 N_A_1037_387#_c_606_n N_A_1745_74#_M1006_d 0.00132295f $X=9.33 $Y=1.07
+ $X2=-0.19 $Y2=-0.245
cc_595 N_A_1037_387#_c_602_n N_A_1745_74#_M1022_d 0.00781907f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_596 N_A_1037_387#_c_637_p N_A_1745_74#_M1022_d 0.00406853f $X=9.415 $Y=2.222
+ $X2=0 $Y2=0
cc_597 N_A_1037_387#_c_614_n N_A_1745_74#_M1022_d 0.0018712f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_598 N_A_1037_387#_c_589_n N_A_1745_74#_c_1567_n 6.35408e-19 $X=8.65 $Y=1.085
+ $X2=0 $Y2=0
cc_599 N_A_1037_387#_c_599_n N_A_1745_74#_c_1567_n 0.00169523f $X=8.825 $Y=0.34
+ $X2=0 $Y2=0
cc_600 N_A_1037_387#_c_601_n N_A_1745_74#_c_1567_n 0.0248143f $X=8.91 $Y=0.905
+ $X2=0 $Y2=0
cc_601 N_A_1037_387#_c_605_n N_A_1745_74#_c_1567_n 0.00569557f $X=9.25 $Y=1.07
+ $X2=0 $Y2=0
cc_602 N_A_1037_387#_c_606_n N_A_1745_74#_c_1567_n 0.0194065f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_603 N_A_1037_387#_M1014_g N_A_1745_74#_c_1556_n 0.0196588f $X=9.835 $Y=2.75
+ $X2=0 $Y2=0
cc_604 N_A_1037_387#_c_637_p N_A_1745_74#_c_1556_n 0.0116449f $X=9.415 $Y=2.222
+ $X2=0 $Y2=0
cc_605 N_A_1037_387#_c_614_n N_A_1745_74#_c_1556_n 0.0370403f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_606 N_A_1037_387#_c_615_n N_A_1745_74#_c_1556_n 0.0025882f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_607 N_A_1037_387#_c_601_n N_A_1745_74#_c_1544_n 0.00376918f $X=8.91 $Y=0.905
+ $X2=0 $Y2=0
cc_608 N_A_1037_387#_c_602_n N_A_1745_74#_c_1545_n 0.0357282f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_609 N_A_1037_387#_c_605_n N_A_1745_74#_c_1545_n 5.18898e-19 $X=9.25 $Y=1.07
+ $X2=0 $Y2=0
cc_610 N_A_1037_387#_c_606_n N_A_1745_74#_c_1545_n 0.014106f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_611 N_A_1037_387#_c_614_n N_A_1745_74#_c_1558_n 0.0123723f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_612 N_A_1037_387#_c_615_n N_A_1745_74#_c_1558_n 0.00350931f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_613 N_A_1037_387#_c_602_n N_A_1745_74#_c_1559_n 0.0141964f $X=9.33 $Y=2.065
+ $X2=0 $Y2=0
cc_614 N_A_1037_387#_c_614_n N_A_1745_74#_c_1559_n 0.0119213f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_615 N_A_1037_387#_c_615_n N_A_1745_74#_c_1559_n 9.43042e-19 $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_616 N_A_1037_387#_M1014_g N_A_1745_74#_c_1560_n 0.00315218f $X=9.835 $Y=2.75
+ $X2=0 $Y2=0
cc_617 N_A_1037_387#_c_614_n N_A_1745_74#_c_1560_n 0.0246458f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_618 N_A_1037_387#_c_615_n N_A_1745_74#_c_1560_n 0.00115119f $X=9.79 $Y=2.215
+ $X2=0 $Y2=0
cc_619 N_A_1037_387#_c_601_n N_A_1745_74#_c_1547_n 7.09256e-19 $X=8.91 $Y=0.905
+ $X2=0 $Y2=0
cc_620 N_A_1037_387#_c_605_n N_A_1745_74#_c_1547_n 5.62433e-19 $X=9.25 $Y=1.07
+ $X2=0 $Y2=0
cc_621 N_A_1037_387#_c_606_n N_A_1745_74#_c_1547_n 0.0131492f $X=9.33 $Y=1.07
+ $X2=0 $Y2=0
cc_622 N_A_1037_387#_M1014_g N_VPWR_c_1828_n 0.00365611f $X=9.835 $Y=2.75 $X2=0
+ $Y2=0
cc_623 N_A_1037_387#_M1016_g N_VPWR_c_1813_n 0.00112709f $X=6.135 $Y=2.525 $X2=0
+ $Y2=0
cc_624 N_A_1037_387#_M1014_g N_VPWR_c_1813_n 0.00448813f $X=9.835 $Y=2.75 $X2=0
+ $Y2=0
cc_625 N_A_1037_387#_M1040_d N_A_415_81#_c_2012_n 0.00645689f $X=5.185 $Y=1.935
+ $X2=0 $Y2=0
cc_626 N_A_1037_387#_c_596_n N_A_415_81#_c_2012_n 0.0308419f $X=5.655 $Y=1.75
+ $X2=0 $Y2=0
cc_627 N_A_1037_387#_c_597_n N_A_415_81#_c_2012_n 0.00244303f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_628 N_A_1037_387#_c_592_n N_A_415_81#_c_2006_n 0.0456345f $X=5.355 $Y=0.74
+ $X2=0 $Y2=0
cc_629 N_A_1037_387#_c_594_n N_A_415_81#_c_2006_n 0.013474f $X=7.055 $Y=0.415
+ $X2=0 $Y2=0
cc_630 N_A_1037_387#_M1016_g N_A_415_81#_c_2013_n 0.00810306f $X=6.135 $Y=2.525
+ $X2=0 $Y2=0
cc_631 N_A_1037_387#_c_596_n N_A_415_81#_c_2013_n 0.00156525f $X=5.655 $Y=1.75
+ $X2=0 $Y2=0
cc_632 N_A_1037_387#_M1017_g N_A_415_81#_c_2007_n 0.00647406f $X=6.52 $Y=0.9
+ $X2=0 $Y2=0
cc_633 N_A_1037_387#_c_597_n N_A_415_81#_c_2007_n 0.0178348f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_634 N_A_1037_387#_c_607_n N_A_415_81#_c_2007_n 0.00642584f $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_635 N_A_1037_387#_c_597_n N_A_415_81#_c_2008_n 0.0143281f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_636 N_A_1037_387#_c_603_n N_A_415_81#_c_2008_n 0.0132455f $X=5.412 $Y=1.275
+ $X2=0 $Y2=0
cc_637 N_A_1037_387#_c_607_n N_A_415_81#_c_2008_n 3.67954e-19 $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_638 N_A_1037_387#_M1016_g N_A_415_81#_c_2014_n 0.0126608f $X=6.135 $Y=2.525
+ $X2=0 $Y2=0
cc_639 N_A_1037_387#_c_587_n N_A_415_81#_c_2014_n 0.00252722f $X=6.445 $Y=1.66
+ $X2=0 $Y2=0
cc_640 N_A_1037_387#_c_597_n N_A_415_81#_c_2014_n 0.00797914f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_641 N_A_1037_387#_M1016_g N_A_415_81#_c_2015_n 0.00250688f $X=6.135 $Y=2.525
+ $X2=0 $Y2=0
cc_642 N_A_1037_387#_c_596_n N_A_415_81#_c_2015_n 0.0145535f $X=5.655 $Y=1.75
+ $X2=0 $Y2=0
cc_643 N_A_1037_387#_c_597_n N_A_415_81#_c_2015_n 0.0167177f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_644 N_A_1037_387#_c_607_n N_A_415_81#_c_2015_n 0.00323027f $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_645 N_A_1037_387#_M1016_g N_A_415_81#_c_2009_n 0.00366894f $X=6.135 $Y=2.525
+ $X2=0 $Y2=0
cc_646 N_A_1037_387#_c_587_n N_A_415_81#_c_2009_n 0.0104145f $X=6.445 $Y=1.66
+ $X2=0 $Y2=0
cc_647 N_A_1037_387#_M1017_g N_A_415_81#_c_2009_n 0.00514657f $X=6.52 $Y=0.9
+ $X2=0 $Y2=0
cc_648 N_A_1037_387#_c_597_n N_A_415_81#_c_2009_n 0.0256546f $X=6.065 $Y=1.75
+ $X2=0 $Y2=0
cc_649 N_A_1037_387#_c_607_n N_A_415_81#_c_2009_n 0.00187233f $X=6.065 $Y=1.66
+ $X2=0 $Y2=0
cc_650 N_A_1037_387#_c_598_n N_VGND_M1034_d 0.0162233f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_651 N_A_1037_387#_c_651_p N_VGND_M1034_d 0.00247125f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_652 N_A_1037_387#_c_600_n N_VGND_M1034_d 6.8704e-19 $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_653 N_A_1037_387#_c_592_n N_VGND_c_2220_n 0.0135874f $X=5.355 $Y=0.74 $X2=0
+ $Y2=0
cc_654 N_A_1037_387#_c_595_n N_VGND_c_2220_n 0.0148789f $X=5.62 $Y=0.415 $X2=0
+ $Y2=0
cc_655 N_A_1037_387#_c_594_n N_VGND_c_2230_n 0.0628116f $X=7.055 $Y=0.415 $X2=0
+ $Y2=0
cc_656 N_A_1037_387#_c_595_n N_VGND_c_2230_n 0.0201144f $X=5.62 $Y=0.415 $X2=0
+ $Y2=0
cc_657 N_A_1037_387#_c_598_n N_VGND_c_2230_n 0.00392706f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_658 N_A_1037_387#_c_604_n N_VGND_c_2230_n 0.00786741f $X=7.14 $Y=0.415 $X2=0
+ $Y2=0
cc_659 N_A_1037_387#_c_589_n N_VGND_c_2231_n 0.00278271f $X=8.65 $Y=1.085 $X2=0
+ $Y2=0
cc_660 N_A_1037_387#_c_598_n N_VGND_c_2231_n 0.00335833f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_661 N_A_1037_387#_c_599_n N_VGND_c_2231_n 0.0579202f $X=8.825 $Y=0.34 $X2=0
+ $Y2=0
cc_662 N_A_1037_387#_c_600_n N_VGND_c_2231_n 0.0118998f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_663 N_A_1037_387#_c_598_n N_VGND_c_2235_n 0.0246013f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_664 N_A_1037_387#_c_600_n N_VGND_c_2235_n 0.0135791f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_665 N_A_1037_387#_c_604_n N_VGND_c_2235_n 0.00555628f $X=7.14 $Y=0.415 $X2=0
+ $Y2=0
cc_666 N_A_1037_387#_c_589_n N_VGND_c_2240_n 0.00358928f $X=8.65 $Y=1.085 $X2=0
+ $Y2=0
cc_667 N_A_1037_387#_c_594_n N_VGND_c_2240_n 0.0456845f $X=7.055 $Y=0.415 $X2=0
+ $Y2=0
cc_668 N_A_1037_387#_c_595_n N_VGND_c_2240_n 0.0138463f $X=5.62 $Y=0.415 $X2=0
+ $Y2=0
cc_669 N_A_1037_387#_c_598_n N_VGND_c_2240_n 0.012145f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_670 N_A_1037_387#_c_599_n N_VGND_c_2240_n 0.0324872f $X=8.825 $Y=0.34 $X2=0
+ $Y2=0
cc_671 N_A_1037_387#_c_600_n N_VGND_c_2240_n 0.00655543f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_672 N_A_1037_387#_c_604_n N_VGND_c_2240_n 0.0055105f $X=7.14 $Y=0.415 $X2=0
+ $Y2=0
cc_673 N_A_1037_387#_c_604_n A_1397_138# 0.00203667f $X=7.14 $Y=0.415 $X2=-0.19
+ $Y2=-0.245
cc_674 N_A_1367_112#_M1000_g N_RESET_B_c_917_n 0.00526413f $X=6.91 $Y=0.9 $X2=0
+ $Y2=0
cc_675 N_A_1367_112#_M1000_g N_RESET_B_M1034_g 0.0394201f $X=6.91 $Y=0.9 $X2=0
+ $Y2=0
cc_676 N_A_1367_112#_c_814_n N_RESET_B_M1034_g 0.00515512f $X=7.19 $Y=1.78 $X2=0
+ $Y2=0
cc_677 N_A_1367_112#_c_831_n N_RESET_B_M1034_g 0.00422682f $X=7.325 $Y=1.005
+ $X2=0 $Y2=0
cc_678 N_A_1367_112#_c_843_n N_RESET_B_M1034_g 0.0067801f $X=8.27 $Y=0.842 $X2=0
+ $Y2=0
cc_679 N_A_1367_112#_c_843_n N_RESET_B_c_920_n 0.00990883f $X=8.27 $Y=0.842
+ $X2=0 $Y2=0
cc_680 N_A_1367_112#_c_814_n N_RESET_B_c_921_n 0.00753567f $X=7.19 $Y=1.78 $X2=0
+ $Y2=0
cc_681 N_A_1367_112#_c_815_n N_RESET_B_c_921_n 0.00620241f $X=7.19 $Y=1.78 $X2=0
+ $Y2=0
cc_682 N_A_1367_112#_M1000_g N_RESET_B_c_922_n 0.00348214f $X=6.91 $Y=0.9 $X2=0
+ $Y2=0
cc_683 N_A_1367_112#_c_814_n N_RESET_B_c_922_n 0.00130495f $X=7.19 $Y=1.78 $X2=0
+ $Y2=0
cc_684 N_A_1367_112#_c_815_n N_RESET_B_c_922_n 0.0199625f $X=7.19 $Y=1.78 $X2=0
+ $Y2=0
cc_685 N_A_1367_112#_M1002_g N_RESET_B_c_932_n 0.0105594f $X=7.025 $Y=2.525
+ $X2=0 $Y2=0
cc_686 N_A_1367_112#_c_814_n N_RESET_B_c_932_n 0.009228f $X=7.19 $Y=1.78 $X2=0
+ $Y2=0
cc_687 N_A_1367_112#_c_815_n N_RESET_B_c_932_n 0.00237054f $X=7.19 $Y=1.78 $X2=0
+ $Y2=0
cc_688 N_A_1367_112#_c_817_n N_RESET_B_c_934_n 0.00719097f $X=8.9 $Y=1.575 $X2=0
+ $Y2=0
cc_689 N_A_1367_112#_c_822_n N_RESET_B_c_934_n 0.030687f $X=8.9 $Y=1.88 $X2=0
+ $Y2=0
cc_690 N_A_1367_112#_M1002_g N_RESET_B_c_939_n 0.0198547f $X=7.025 $Y=2.525
+ $X2=0 $Y2=0
cc_691 N_A_1367_112#_c_816_n N_A_1233_138#_M1028_g 0.00313626f $X=8.57 $Y=1.405
+ $X2=0 $Y2=0
cc_692 N_A_1367_112#_c_843_n N_A_1233_138#_M1028_g 0.0131882f $X=8.27 $Y=0.842
+ $X2=0 $Y2=0
cc_693 N_A_1367_112#_c_816_n N_A_1233_138#_c_1132_n 0.00107424f $X=8.57 $Y=1.405
+ $X2=0 $Y2=0
cc_694 N_A_1367_112#_c_817_n N_A_1233_138#_c_1132_n 0.0132267f $X=8.9 $Y=1.575
+ $X2=0 $Y2=0
cc_695 N_A_1367_112#_c_822_n N_A_1233_138#_c_1132_n 0.00132806f $X=8.9 $Y=1.88
+ $X2=0 $Y2=0
cc_696 N_A_1367_112#_c_845_n N_A_1233_138#_c_1132_n 0.00405015f $X=8.57 $Y=0.842
+ $X2=0 $Y2=0
cc_697 N_A_1367_112#_c_822_n N_A_1233_138#_M1018_g 0.0207862f $X=8.9 $Y=1.88
+ $X2=0 $Y2=0
cc_698 N_A_1367_112#_M1000_g N_A_1233_138#_c_1154_n 0.00473706f $X=6.91 $Y=0.9
+ $X2=0 $Y2=0
cc_699 N_A_1367_112#_c_831_n N_A_1233_138#_c_1154_n 0.0130756f $X=7.325 $Y=1.005
+ $X2=0 $Y2=0
cc_700 N_A_1367_112#_M1000_g N_A_1233_138#_c_1133_n 0.00952502f $X=6.91 $Y=0.9
+ $X2=0 $Y2=0
cc_701 N_A_1367_112#_M1002_g N_A_1233_138#_c_1133_n 0.00540451f $X=7.025
+ $Y=2.525 $X2=0 $Y2=0
cc_702 N_A_1367_112#_c_814_n N_A_1233_138#_c_1133_n 0.062072f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_703 N_A_1367_112#_c_815_n N_A_1233_138#_c_1133_n 0.010397f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_704 N_A_1367_112#_c_831_n N_A_1233_138#_c_1133_n 0.00114989f $X=7.325
+ $Y=1.005 $X2=0 $Y2=0
cc_705 N_A_1367_112#_M1002_g N_A_1233_138#_c_1177_n 0.0121428f $X=7.025 $Y=2.525
+ $X2=0 $Y2=0
cc_706 N_A_1367_112#_c_814_n N_A_1233_138#_c_1177_n 0.00524316f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_707 N_A_1367_112#_c_815_n N_A_1233_138#_c_1177_n 0.00200238f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_708 N_A_1367_112#_M1002_g N_A_1233_138#_c_1134_n 0.00347134f $X=7.025
+ $Y=2.525 $X2=0 $Y2=0
cc_709 N_A_1367_112#_c_814_n N_A_1233_138#_c_1134_n 0.0274324f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_710 N_A_1367_112#_c_815_n N_A_1233_138#_c_1134_n 0.00201777f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_711 N_A_1367_112#_c_814_n N_A_1233_138#_c_1135_n 0.0268294f $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_712 N_A_1367_112#_c_843_n N_A_1233_138#_c_1135_n 0.0133196f $X=8.27 $Y=0.842
+ $X2=0 $Y2=0
cc_713 N_A_1367_112#_c_816_n N_A_1233_138#_c_1136_n 0.0115079f $X=8.57 $Y=1.405
+ $X2=0 $Y2=0
cc_714 N_A_1367_112#_c_817_n N_A_1233_138#_c_1136_n 0.0142233f $X=8.9 $Y=1.575
+ $X2=0 $Y2=0
cc_715 N_A_1367_112#_c_843_n N_A_1233_138#_c_1136_n 0.0443118f $X=8.27 $Y=0.842
+ $X2=0 $Y2=0
cc_716 N_A_1367_112#_c_816_n N_A_1233_138#_c_1137_n 0.00161618f $X=8.57 $Y=1.405
+ $X2=0 $Y2=0
cc_717 N_A_1367_112#_c_817_n N_A_1233_138#_c_1137_n 3.02987e-19 $X=8.9 $Y=1.575
+ $X2=0 $Y2=0
cc_718 N_A_1367_112#_c_843_n N_A_1233_138#_c_1137_n 0.00252719f $X=8.27 $Y=0.842
+ $X2=0 $Y2=0
cc_719 N_A_1367_112#_c_845_n N_A_1233_138#_c_1137_n 0.00137742f $X=8.57 $Y=0.842
+ $X2=0 $Y2=0
cc_720 N_A_1367_112#_M1000_g N_A_1233_138#_c_1138_n 0.00108413f $X=6.91 $Y=0.9
+ $X2=0 $Y2=0
cc_721 N_A_1367_112#_M1002_g N_A_1233_138#_c_1145_n 0.00102488f $X=7.025
+ $Y=2.525 $X2=0 $Y2=0
cc_722 N_A_1367_112#_M1002_g N_A_834_93#_M1012_g 0.0415994f $X=7.025 $Y=2.525
+ $X2=0 $Y2=0
cc_723 N_A_1367_112#_M1002_g N_A_834_93#_c_1279_n 0.0120603f $X=7.025 $Y=2.525
+ $X2=0 $Y2=0
cc_724 N_A_1367_112#_c_822_n N_A_834_93#_c_1279_n 0.00373896f $X=8.9 $Y=1.88
+ $X2=0 $Y2=0
cc_725 N_A_1367_112#_c_822_n N_A_834_93#_M1022_g 0.0161095f $X=8.9 $Y=1.88 $X2=0
+ $Y2=0
cc_726 N_A_1367_112#_c_817_n N_A_834_93#_c_1267_n 0.0021457f $X=8.9 $Y=1.575
+ $X2=0 $Y2=0
cc_727 N_A_1367_112#_c_822_n N_A_834_93#_c_1267_n 0.00253734f $X=8.9 $Y=1.88
+ $X2=0 $Y2=0
cc_728 N_A_1367_112#_c_822_n N_A_1745_74#_c_1556_n 0.00739135f $X=8.9 $Y=1.88
+ $X2=0 $Y2=0
cc_729 N_A_1367_112#_M1002_g N_VPWR_c_1816_n 0.004022f $X=7.025 $Y=2.525 $X2=0
+ $Y2=0
cc_730 N_A_1367_112#_c_817_n N_VPWR_c_1818_n 0.00342759f $X=8.9 $Y=1.575 $X2=0
+ $Y2=0
cc_731 N_A_1367_112#_c_822_n N_VPWR_c_1818_n 0.0352169f $X=8.9 $Y=1.88 $X2=0
+ $Y2=0
cc_732 N_A_1367_112#_c_845_n N_VPWR_c_1818_n 0.00374786f $X=8.57 $Y=0.842 $X2=0
+ $Y2=0
cc_733 N_A_1367_112#_c_822_n N_VPWR_c_1828_n 0.00741793f $X=8.9 $Y=1.88 $X2=0
+ $Y2=0
cc_734 N_A_1367_112#_M1002_g N_VPWR_c_1813_n 0.00112709f $X=7.025 $Y=2.525 $X2=0
+ $Y2=0
cc_735 N_A_1367_112#_c_822_n N_VPWR_c_1813_n 0.00901294f $X=8.9 $Y=1.88 $X2=0
+ $Y2=0
cc_736 N_A_1367_112#_M1000_g N_A_415_81#_c_2009_n 3.0177e-19 $X=6.91 $Y=0.9
+ $X2=0 $Y2=0
cc_737 N_A_1367_112#_c_815_n N_A_415_81#_c_2009_n 6.15582e-19 $X=7.19 $Y=1.78
+ $X2=0 $Y2=0
cc_738 N_A_1367_112#_c_843_n N_VGND_M1034_d 0.0155117f $X=8.27 $Y=0.842 $X2=0
+ $Y2=0
cc_739 N_A_1367_112#_c_831_n A_1397_138# 0.00260878f $X=7.325 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_740 N_RESET_B_c_920_n N_A_1233_138#_M1028_g 0.00269339f $X=7.575 $Y=1.26
+ $X2=0 $Y2=0
cc_741 N_RESET_B_c_934_n N_A_1233_138#_M1018_g 0.00776847f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_742 N_RESET_B_c_932_n N_A_1233_138#_c_1141_n 0.00814681f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_743 N_RESET_B_M1034_g N_A_1233_138#_c_1154_n 2.03434e-19 $X=7.3 $Y=0.9 $X2=0
+ $Y2=0
cc_744 N_RESET_B_M1034_g N_A_1233_138#_c_1133_n 2.11405e-19 $X=7.3 $Y=0.9 $X2=0
+ $Y2=0
cc_745 N_RESET_B_c_932_n N_A_1233_138#_c_1133_n 0.0238647f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_746 N_RESET_B_c_932_n N_A_1233_138#_c_1177_n 0.0208177f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_747 N_RESET_B_c_922_n N_A_1233_138#_c_1134_n 0.0119425f $X=7.66 $Y=1.82 $X2=0
+ $Y2=0
cc_748 N_RESET_B_M1003_g N_A_1233_138#_c_1134_n 0.0243684f $X=7.665 $Y=2.525
+ $X2=0 $Y2=0
cc_749 N_RESET_B_c_932_n N_A_1233_138#_c_1134_n 0.0261145f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_750 N_RESET_B_c_935_n N_A_1233_138#_c_1134_n 0.0106292f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_751 N_RESET_B_c_936_n N_A_1233_138#_c_1134_n 0.0363198f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_752 N_RESET_B_c_939_n N_A_1233_138#_c_1134_n 0.0143305f $X=7.98 $Y=1.985
+ $X2=0 $Y2=0
cc_753 N_RESET_B_c_920_n N_A_1233_138#_c_1135_n 0.00533024f $X=7.575 $Y=1.26
+ $X2=0 $Y2=0
cc_754 N_RESET_B_c_922_n N_A_1233_138#_c_1135_n 0.00463689f $X=7.66 $Y=1.82
+ $X2=0 $Y2=0
cc_755 N_RESET_B_c_920_n N_A_1233_138#_c_1136_n 0.00188178f $X=7.575 $Y=1.26
+ $X2=0 $Y2=0
cc_756 N_RESET_B_c_922_n N_A_1233_138#_c_1136_n 0.00587638f $X=7.66 $Y=1.82
+ $X2=0 $Y2=0
cc_757 N_RESET_B_c_932_n N_A_1233_138#_c_1136_n 0.00357593f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_758 N_RESET_B_c_934_n N_A_1233_138#_c_1136_n 0.00641796f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_759 N_RESET_B_c_935_n N_A_1233_138#_c_1136_n 0.00373314f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_760 N_RESET_B_c_936_n N_A_1233_138#_c_1136_n 0.0158779f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_761 N_RESET_B_c_939_n N_A_1233_138#_c_1136_n 0.00718951f $X=7.98 $Y=1.985
+ $X2=0 $Y2=0
cc_762 N_RESET_B_c_920_n N_A_1233_138#_c_1137_n 0.0194898f $X=7.575 $Y=1.26
+ $X2=0 $Y2=0
cc_763 N_RESET_B_c_934_n N_A_1233_138#_c_1137_n 0.00588371f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_764 N_RESET_B_c_936_n N_A_1233_138#_c_1137_n 6.12607e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_765 N_RESET_B_c_939_n N_A_1233_138#_c_1137_n 0.00918526f $X=7.98 $Y=1.985
+ $X2=0 $Y2=0
cc_766 N_RESET_B_c_932_n N_A_834_93#_M1026_s 0.00114543f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_767 N_RESET_B_c_932_n N_A_834_93#_M1040_g 0.00406718f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_768 N_RESET_B_c_932_n N_A_834_93#_c_1261_n 0.00281312f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_769 N_RESET_B_c_932_n N_A_834_93#_c_1263_n 0.00174208f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_770 N_RESET_B_c_917_n N_A_834_93#_c_1265_n 0.00526413f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_771 N_RESET_B_c_932_n N_A_834_93#_M1012_g 0.00440273f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_772 N_RESET_B_M1003_g N_A_834_93#_c_1279_n 0.0119874f $X=7.665 $Y=2.525 $X2=0
+ $Y2=0
cc_773 N_RESET_B_c_934_n N_A_834_93#_M1022_g 0.013655f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_774 N_RESET_B_c_934_n N_A_834_93#_c_1266_n 0.00393672f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_775 N_RESET_B_c_917_n N_A_834_93#_c_1290_n 0.00125026f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_776 N_RESET_B_c_933_n N_A_834_93#_c_1284_n 5.48045e-19 $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_777 N_RESET_B_c_938_n N_A_834_93#_c_1284_n 0.003169f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_778 N_RESET_B_c_917_n N_A_834_93#_c_1270_n 0.00782328f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_779 N_RESET_B_c_925_n N_A_834_93#_c_1299_n 6.92995e-19 $X=3.93 $Y=1.995 $X2=0
+ $Y2=0
cc_780 N_RESET_B_c_926_n N_A_834_93#_c_1299_n 0.00296415f $X=3.715 $Y=1.995
+ $X2=0 $Y2=0
cc_781 N_RESET_B_c_932_n N_A_834_93#_c_1299_n 0.0341168f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_782 N_RESET_B_c_933_n N_A_834_93#_c_1299_n 0.00205234f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_783 N_RESET_B_c_938_n N_A_834_93#_c_1299_n 0.0156062f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_784 N_RESET_B_c_932_n N_A_834_93#_c_1271_n 0.0089475f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_785 N_RESET_B_c_932_n N_A_834_93#_c_1272_n 6.06994e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_786 N_RESET_B_c_917_n N_A_834_93#_c_1273_n 0.0102563f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_787 N_RESET_B_M1045_g N_A_2003_48#_M1032_g 0.0216011f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_788 N_RESET_B_M1031_g N_A_2003_48#_M1010_g 0.0177072f $X=10.94 $Y=2.75 $X2=0
+ $Y2=0
cc_789 N_RESET_B_c_934_n N_A_2003_48#_M1010_g 0.0033828f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_790 N_RESET_B_c_940_n N_A_2003_48#_M1010_g 0.00106389f $X=10.75 $Y=1.985
+ $X2=0 $Y2=0
cc_791 N_RESET_B_c_941_n N_A_2003_48#_M1010_g 0.029932f $X=10.94 $Y=1.985 $X2=0
+ $Y2=0
cc_792 N_RESET_B_M1045_g N_A_2003_48#_c_1452_n 0.0128807f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_793 N_RESET_B_c_934_n N_A_2003_48#_c_1452_n 0.00879069f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_794 RESET_B N_A_2003_48#_c_1452_n 0.00259932f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_795 N_RESET_B_c_940_n N_A_2003_48#_c_1452_n 0.0152297f $X=10.75 $Y=1.985
+ $X2=0 $Y2=0
cc_796 N_RESET_B_c_941_n N_A_2003_48#_c_1452_n 0.00391556f $X=10.94 $Y=1.985
+ $X2=0 $Y2=0
cc_797 N_RESET_B_M1045_g N_A_2003_48#_c_1453_n 9.6789e-19 $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_798 N_RESET_B_M1045_g N_A_2003_48#_c_1455_n 0.00118187f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_799 N_RESET_B_c_934_n N_A_2003_48#_c_1455_n 0.00250381f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_800 N_RESET_B_M1045_g N_A_2003_48#_c_1456_n 0.029932f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_801 N_RESET_B_M1031_g N_A_2003_48#_c_1460_n 0.00826031f $X=10.94 $Y=2.75
+ $X2=0 $Y2=0
cc_802 N_RESET_B_M1045_g N_A_2003_48#_c_1457_n 0.00453304f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_803 RESET_B N_A_2003_48#_c_1457_n 0.00621393f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_804 N_RESET_B_c_940_n N_A_2003_48#_c_1457_n 0.0154382f $X=10.75 $Y=1.985
+ $X2=0 $Y2=0
cc_805 N_RESET_B_c_941_n N_A_2003_48#_c_1457_n 0.0113972f $X=10.94 $Y=1.985
+ $X2=0 $Y2=0
cc_806 N_RESET_B_c_934_n N_A_1745_74#_M1022_d 0.00241396f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_807 N_RESET_B_M1045_g N_A_1745_74#_c_1535_n 0.0694909f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_808 N_RESET_B_c_941_n N_A_1745_74#_M1044_g 0.0292624f $X=10.94 $Y=1.985 $X2=0
+ $Y2=0
cc_809 N_RESET_B_M1045_g N_A_1745_74#_c_1541_n 0.00550286f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_810 N_RESET_B_c_934_n N_A_1745_74#_c_1556_n 0.00707715f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_811 N_RESET_B_M1045_g N_A_1745_74#_c_1546_n 0.0150978f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_812 N_RESET_B_M1045_g N_A_1745_74#_c_1558_n 8.1654e-19 $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_813 N_RESET_B_c_934_n N_A_1745_74#_c_1558_n 0.0117357f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_814 N_RESET_B_c_940_n N_A_1745_74#_c_1558_n 0.00391217f $X=10.75 $Y=1.985
+ $X2=0 $Y2=0
cc_815 N_RESET_B_c_934_n N_A_1745_74#_c_1559_n 0.00499654f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_816 N_RESET_B_M1031_g N_A_1745_74#_c_1560_n 0.00187713f $X=10.94 $Y=2.75
+ $X2=0 $Y2=0
cc_817 N_RESET_B_c_934_n N_A_1745_74#_c_1560_n 0.0200435f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_818 RESET_B N_A_1745_74#_c_1560_n 4.97327e-19 $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_819 N_RESET_B_c_940_n N_A_1745_74#_c_1560_n 0.00972451f $X=10.75 $Y=1.985
+ $X2=0 $Y2=0
cc_820 N_RESET_B_c_941_n N_A_1745_74#_c_1560_n 8.72425e-19 $X=10.94 $Y=1.985
+ $X2=0 $Y2=0
cc_821 N_RESET_B_M1045_g N_A_1745_74#_c_1548_n 0.00118187f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_822 N_RESET_B_c_941_n N_A_1745_74#_c_1549_n 0.00231899f $X=10.94 $Y=1.985
+ $X2=0 $Y2=0
cc_823 N_RESET_B_c_932_n N_VPWR_M1026_d 4.24275e-19 $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_824 N_RESET_B_c_934_n N_VPWR_M1018_s 0.00559626f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_825 N_RESET_B_c_931_n N_VPWR_c_1814_n 0.00408327f $X=3.59 $Y=2.245 $X2=0
+ $Y2=0
cc_826 N_RESET_B_M1003_g N_VPWR_c_1816_n 0.00399686f $X=7.665 $Y=2.525 $X2=0
+ $Y2=0
cc_827 N_RESET_B_c_932_n N_VPWR_c_1816_n 7.4258e-19 $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_828 N_RESET_B_c_922_n N_VPWR_c_1818_n 0.00162316f $X=7.66 $Y=1.82 $X2=0 $Y2=0
cc_829 N_RESET_B_M1003_g N_VPWR_c_1818_n 0.00702856f $X=7.665 $Y=2.525 $X2=0
+ $Y2=0
cc_830 N_RESET_B_c_934_n N_VPWR_c_1818_n 0.0183856f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_831 N_RESET_B_c_935_n N_VPWR_c_1818_n 5.40997e-19 $X=8.065 $Y=2.035 $X2=0
+ $Y2=0
cc_832 N_RESET_B_c_936_n N_VPWR_c_1818_n 0.0179605f $X=7.92 $Y=2.035 $X2=0 $Y2=0
cc_833 N_RESET_B_c_939_n N_VPWR_c_1818_n 0.00111758f $X=7.98 $Y=1.985 $X2=0
+ $Y2=0
cc_834 N_RESET_B_M1031_g N_VPWR_c_1819_n 0.00674123f $X=10.94 $Y=2.75 $X2=0
+ $Y2=0
cc_835 N_RESET_B_c_934_n N_VPWR_c_1819_n 0.00540169f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_836 RESET_B N_VPWR_c_1819_n 0.00113612f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_837 N_RESET_B_c_940_n N_VPWR_c_1819_n 0.00684931f $X=10.75 $Y=1.985 $X2=0
+ $Y2=0
cc_838 N_RESET_B_c_941_n N_VPWR_c_1819_n 0.00269311f $X=10.94 $Y=1.985 $X2=0
+ $Y2=0
cc_839 N_RESET_B_c_931_n N_VPWR_c_1826_n 0.00440684f $X=3.59 $Y=2.245 $X2=0
+ $Y2=0
cc_840 N_RESET_B_M1031_g N_VPWR_c_1833_n 0.005209f $X=10.94 $Y=2.75 $X2=0 $Y2=0
cc_841 N_RESET_B_M1003_g N_VPWR_c_1813_n 0.00112709f $X=7.665 $Y=2.525 $X2=0
+ $Y2=0
cc_842 N_RESET_B_M1031_g N_VPWR_c_1813_n 0.00985174f $X=10.94 $Y=2.75 $X2=0
+ $Y2=0
cc_843 N_RESET_B_c_931_n N_VPWR_c_1813_n 0.00487308f $X=3.59 $Y=2.245 $X2=0
+ $Y2=0
cc_844 N_RESET_B_M1013_g N_A_415_81#_c_2004_n 0.0122453f $X=3.54 $Y=0.615 $X2=0
+ $Y2=0
cc_845 N_RESET_B_M1013_g N_A_415_81#_c_2005_n 0.0204261f $X=3.54 $Y=0.615 $X2=0
+ $Y2=0
cc_846 N_RESET_B_c_926_n N_A_415_81#_c_2005_n 0.0157764f $X=3.715 $Y=1.995 $X2=0
+ $Y2=0
cc_847 N_RESET_B_c_931_n N_A_415_81#_c_2005_n 0.00522456f $X=3.59 $Y=2.245 $X2=0
+ $Y2=0
cc_848 N_RESET_B_c_933_n N_A_415_81#_c_2005_n 0.00108729f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_849 N_RESET_B_c_938_n N_A_415_81#_c_2005_n 0.0228135f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_850 N_RESET_B_c_925_n N_A_415_81#_c_2012_n 0.00194418f $X=3.93 $Y=1.995 $X2=0
+ $Y2=0
cc_851 N_RESET_B_c_932_n N_A_415_81#_c_2012_n 0.0181319f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_852 N_RESET_B_c_933_n N_A_415_81#_c_2012_n 0.00350898f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_853 N_RESET_B_c_938_n N_A_415_81#_c_2012_n 0.00625123f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_854 N_RESET_B_c_932_n N_A_415_81#_c_2007_n 0.00381691f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_855 N_RESET_B_c_932_n N_A_415_81#_c_2014_n 0.0160834f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_856 N_RESET_B_c_932_n N_A_415_81#_c_2015_n 0.0155324f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_857 N_RESET_B_c_932_n N_A_415_81#_c_2009_n 0.011933f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_858 N_RESET_B_c_925_n N_A_415_81#_c_2018_n 0.00709459f $X=3.93 $Y=1.995 $X2=0
+ $Y2=0
cc_859 N_RESET_B_c_931_n N_A_415_81#_c_2018_n 0.0253011f $X=3.59 $Y=2.245 $X2=0
+ $Y2=0
cc_860 N_RESET_B_c_933_n N_A_415_81#_c_2018_n 7.08105e-19 $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_861 N_RESET_B_c_938_n N_A_415_81#_c_2018_n 0.017495f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_862 N_RESET_B_M1013_g N_VGND_c_2219_n 0.00138718f $X=3.54 $Y=0.615 $X2=0
+ $Y2=0
cc_863 N_RESET_B_c_917_n N_VGND_c_2219_n 0.0219402f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_864 N_RESET_B_c_917_n N_VGND_c_2220_n 0.02563f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_865 N_RESET_B_M1045_g N_VGND_c_2221_n 0.0101056f $X=10.63 $Y=0.58 $X2=0 $Y2=0
cc_866 N_RESET_B_c_918_n N_VGND_c_2225_n 0.00672974f $X=3.615 $Y=0.18 $X2=0
+ $Y2=0
cc_867 N_RESET_B_c_917_n N_VGND_c_2227_n 0.0221273f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_868 N_RESET_B_c_917_n N_VGND_c_2230_n 0.0531974f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_869 N_RESET_B_M1045_g N_VGND_c_2232_n 0.00383152f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_870 N_RESET_B_c_917_n N_VGND_c_2235_n 0.0108145f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_871 N_RESET_B_c_917_n N_VGND_c_2240_n 0.0880414f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_872 N_RESET_B_c_918_n N_VGND_c_2240_n 0.0112172f $X=3.615 $Y=0.18 $X2=0 $Y2=0
cc_873 N_RESET_B_M1045_g N_VGND_c_2240_n 0.0075694f $X=10.63 $Y=0.58 $X2=0 $Y2=0
cc_874 N_RESET_B_M1013_g N_noxref_24_c_2365_n 0.00696122f $X=3.54 $Y=0.615 $X2=0
+ $Y2=0
cc_875 N_A_1233_138#_c_1141_n N_A_834_93#_c_1276_n 0.00405916f $X=6.715 $Y=2.59
+ $X2=0 $Y2=0
cc_876 N_A_1233_138#_c_1138_n N_A_834_93#_c_1265_n 0.00525257f $X=6.305 $Y=0.87
+ $X2=0 $Y2=0
cc_877 N_A_1233_138#_c_1141_n N_A_834_93#_M1012_g 0.011473f $X=6.715 $Y=2.59
+ $X2=0 $Y2=0
cc_878 N_A_1233_138#_c_1133_n N_A_834_93#_M1012_g 0.00319744f $X=6.8 $Y=2.32
+ $X2=0 $Y2=0
cc_879 N_A_1233_138#_c_1145_n N_A_834_93#_M1012_g 0.00561127f $X=6.8 $Y=2.537
+ $X2=0 $Y2=0
cc_880 N_A_1233_138#_M1018_g N_A_834_93#_c_1279_n 0.0123594f $X=8.675 $Y=2.235
+ $X2=0 $Y2=0
cc_881 N_A_1233_138#_c_1177_n N_A_834_93#_c_1279_n 0.00156425f $X=7.495 $Y=2.405
+ $X2=0 $Y2=0
cc_882 N_A_1233_138#_c_1134_n N_A_834_93#_c_1279_n 0.00654552f $X=7.58 $Y=2.32
+ $X2=0 $Y2=0
cc_883 N_A_1233_138#_c_1145_n N_A_834_93#_c_1279_n 0.00142193f $X=6.8 $Y=2.537
+ $X2=0 $Y2=0
cc_884 N_A_1233_138#_M1018_g N_A_834_93#_M1022_g 0.0083082f $X=8.675 $Y=2.235
+ $X2=0 $Y2=0
cc_885 N_A_1233_138#_c_1132_n N_A_834_93#_c_1267_n 0.0083082f $X=8.585 $Y=1.52
+ $X2=0 $Y2=0
cc_886 N_A_1233_138#_c_1177_n N_VPWR_M1002_d 0.00774864f $X=7.495 $Y=2.405 $X2=0
+ $Y2=0
cc_887 N_A_1233_138#_c_1134_n N_VPWR_M1002_d 2.18741e-19 $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_888 N_A_1233_138#_c_1177_n N_VPWR_c_1816_n 0.0248409f $X=7.495 $Y=2.405 $X2=0
+ $Y2=0
cc_889 N_A_1233_138#_c_1134_n N_VPWR_c_1816_n 0.00570779f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_890 N_A_1233_138#_c_1145_n N_VPWR_c_1816_n 0.00116897f $X=6.8 $Y=2.537 $X2=0
+ $Y2=0
cc_891 N_A_1233_138#_c_1134_n N_VPWR_c_1817_n 0.00728415f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_892 N_A_1233_138#_c_1132_n N_VPWR_c_1818_n 0.004245f $X=8.585 $Y=1.52 $X2=0
+ $Y2=0
cc_893 N_A_1233_138#_M1018_g N_VPWR_c_1818_n 0.00504062f $X=8.675 $Y=2.235 $X2=0
+ $Y2=0
cc_894 N_A_1233_138#_c_1134_n N_VPWR_c_1818_n 0.0227301f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_895 N_A_1233_138#_c_1141_n N_VPWR_c_1832_n 0.00986974f $X=6.715 $Y=2.59 $X2=0
+ $Y2=0
cc_896 N_A_1233_138#_c_1145_n N_VPWR_c_1832_n 0.00388446f $X=6.8 $Y=2.537 $X2=0
+ $Y2=0
cc_897 N_A_1233_138#_M1018_g N_VPWR_c_1813_n 0.00112709f $X=8.675 $Y=2.235 $X2=0
+ $Y2=0
cc_898 N_A_1233_138#_c_1141_n N_VPWR_c_1813_n 0.0123602f $X=6.715 $Y=2.59 $X2=0
+ $Y2=0
cc_899 N_A_1233_138#_c_1177_n N_VPWR_c_1813_n 0.00921351f $X=7.495 $Y=2.405
+ $X2=0 $Y2=0
cc_900 N_A_1233_138#_c_1134_n N_VPWR_c_1813_n 0.0155036f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_901 N_A_1233_138#_c_1145_n N_VPWR_c_1813_n 0.00467845f $X=6.8 $Y=2.537 $X2=0
+ $Y2=0
cc_902 N_A_1233_138#_c_1138_n N_A_415_81#_c_2006_n 0.0152023f $X=6.305 $Y=0.87
+ $X2=0 $Y2=0
cc_903 N_A_1233_138#_c_1133_n N_A_415_81#_c_2013_n 0.0014826f $X=6.8 $Y=2.32
+ $X2=0 $Y2=0
cc_904 N_A_1233_138#_c_1145_n N_A_415_81#_c_2013_n 0.0027162f $X=6.8 $Y=2.537
+ $X2=0 $Y2=0
cc_905 N_A_1233_138#_c_1154_n N_A_415_81#_c_2007_n 0.00571315f $X=6.715 $Y=0.99
+ $X2=0 $Y2=0
cc_906 N_A_1233_138#_c_1133_n N_A_415_81#_c_2007_n 0.0135849f $X=6.8 $Y=2.32
+ $X2=0 $Y2=0
cc_907 N_A_1233_138#_c_1138_n N_A_415_81#_c_2007_n 0.021789f $X=6.305 $Y=0.87
+ $X2=0 $Y2=0
cc_908 N_A_1233_138#_c_1141_n N_A_415_81#_c_2014_n 0.0200051f $X=6.715 $Y=2.59
+ $X2=0 $Y2=0
cc_909 N_A_1233_138#_c_1133_n N_A_415_81#_c_2014_n 0.013599f $X=6.8 $Y=2.32
+ $X2=0 $Y2=0
cc_910 N_A_1233_138#_c_1133_n N_A_415_81#_c_2009_n 0.048566f $X=6.8 $Y=2.32
+ $X2=0 $Y2=0
cc_911 N_A_1233_138#_M1028_g N_VGND_c_2231_n 0.00278271f $X=8.175 $Y=0.74 $X2=0
+ $Y2=0
cc_912 N_A_1233_138#_M1028_g N_VGND_c_2235_n 0.00118431f $X=8.175 $Y=0.74 $X2=0
+ $Y2=0
cc_913 N_A_1233_138#_M1028_g N_VGND_c_2240_n 0.00358928f $X=8.175 $Y=0.74 $X2=0
+ $Y2=0
cc_914 N_A_1233_138#_c_1154_n A_1319_138# 0.00422251f $X=6.715 $Y=0.99 $X2=-0.19
+ $Y2=-0.245
cc_915 N_A_1233_138#_c_1133_n A_1319_138# 3.82916e-19 $X=6.8 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_916 N_A_834_93#_M1036_g N_A_2003_48#_M1032_g 0.0336121f $X=9.7 $Y=0.58 $X2=0
+ $Y2=0
cc_917 N_A_834_93#_c_1266_n N_A_2003_48#_M1010_g 0.00387806f $X=9.625 $Y=1.585
+ $X2=0 $Y2=0
cc_918 N_A_834_93#_M1036_g N_A_2003_48#_c_1455_n 0.00111235f $X=9.7 $Y=0.58
+ $X2=0 $Y2=0
cc_919 N_A_834_93#_c_1266_n N_A_2003_48#_c_1456_n 0.0336121f $X=9.625 $Y=1.585
+ $X2=0 $Y2=0
cc_920 N_A_834_93#_M1036_g N_A_1745_74#_c_1567_n 0.0163048f $X=9.7 $Y=0.58 $X2=0
+ $Y2=0
cc_921 N_A_834_93#_M1022_g N_A_1745_74#_c_1556_n 0.00594721f $X=9.125 $Y=2.235
+ $X2=0 $Y2=0
cc_922 N_A_834_93#_M1036_g N_A_1745_74#_c_1544_n 0.00585097f $X=9.7 $Y=0.58
+ $X2=0 $Y2=0
cc_923 N_A_834_93#_c_1266_n N_A_1745_74#_c_1545_n 0.00934901f $X=9.625 $Y=1.585
+ $X2=0 $Y2=0
cc_924 N_A_834_93#_M1036_g N_A_1745_74#_c_1545_n 0.0140808f $X=9.7 $Y=0.58 $X2=0
+ $Y2=0
cc_925 N_A_834_93#_M1036_g N_A_1745_74#_c_1546_n 0.00333053f $X=9.7 $Y=0.58
+ $X2=0 $Y2=0
cc_926 N_A_834_93#_c_1266_n N_A_1745_74#_c_1558_n 3.21304e-19 $X=9.625 $Y=1.585
+ $X2=0 $Y2=0
cc_927 N_A_834_93#_M1036_g N_A_1745_74#_c_1547_n 0.00274755f $X=9.7 $Y=0.58
+ $X2=0 $Y2=0
cc_928 N_A_834_93#_c_1299_n N_VPWR_M1026_d 0.00319612f $X=4.42 $Y=2.12 $X2=0
+ $Y2=0
cc_929 N_A_834_93#_M1040_g N_VPWR_c_1815_n 0.0105673f $X=5.095 $Y=2.495 $X2=0
+ $Y2=0
cc_930 N_A_834_93#_c_1263_n N_VPWR_c_1815_n 0.00201199f $X=5.615 $Y=3.075 $X2=0
+ $Y2=0
cc_931 N_A_834_93#_c_1277_n N_VPWR_c_1815_n 6.90101e-19 $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_932 N_A_834_93#_M1012_g N_VPWR_c_1816_n 0.00614938f $X=6.635 $Y=2.525 $X2=0
+ $Y2=0
cc_933 N_A_834_93#_c_1279_n N_VPWR_c_1816_n 0.0264476f $X=9.035 $Y=3.15 $X2=0
+ $Y2=0
cc_934 N_A_834_93#_c_1279_n N_VPWR_c_1817_n 0.0260616f $X=9.035 $Y=3.15 $X2=0
+ $Y2=0
cc_935 N_A_834_93#_c_1279_n N_VPWR_c_1818_n 0.0170937f $X=9.035 $Y=3.15 $X2=0
+ $Y2=0
cc_936 N_A_834_93#_M1022_g N_VPWR_c_1818_n 0.00538421f $X=9.125 $Y=2.235 $X2=0
+ $Y2=0
cc_937 N_A_834_93#_c_1279_n N_VPWR_c_1828_n 0.0212627f $X=9.035 $Y=3.15 $X2=0
+ $Y2=0
cc_938 N_A_834_93#_M1040_g N_VPWR_c_1832_n 0.00401239f $X=5.095 $Y=2.495 $X2=0
+ $Y2=0
cc_939 N_A_834_93#_c_1277_n N_VPWR_c_1832_n 0.0468577f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_940 N_A_834_93#_M1040_g N_VPWR_c_1813_n 0.00502672f $X=5.095 $Y=2.495 $X2=0
+ $Y2=0
cc_941 N_A_834_93#_c_1276_n N_VPWR_c_1813_n 0.0243879f $X=6.545 $Y=3.15 $X2=0
+ $Y2=0
cc_942 N_A_834_93#_c_1277_n N_VPWR_c_1813_n 0.00590281f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_943 N_A_834_93#_c_1279_n N_VPWR_c_1813_n 0.0712383f $X=9.035 $Y=3.15 $X2=0
+ $Y2=0
cc_944 N_A_834_93#_c_1283_n N_VPWR_c_1813_n 0.00500351f $X=6.635 $Y=3.15 $X2=0
+ $Y2=0
cc_945 N_A_834_93#_M1026_s N_A_415_81#_c_2012_n 0.00756295f $X=4.275 $Y=1.935
+ $X2=0 $Y2=0
cc_946 N_A_834_93#_M1040_g N_A_415_81#_c_2012_n 0.0156657f $X=5.095 $Y=2.495
+ $X2=0 $Y2=0
cc_947 N_A_834_93#_c_1263_n N_A_415_81#_c_2012_n 0.0133305f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_948 N_A_834_93#_c_1276_n N_A_415_81#_c_2012_n 7.47264e-19 $X=6.545 $Y=3.15
+ $X2=0 $Y2=0
cc_949 N_A_834_93#_c_1299_n N_A_415_81#_c_2012_n 0.0269661f $X=4.42 $Y=2.12
+ $X2=0 $Y2=0
cc_950 N_A_834_93#_c_1271_n N_A_415_81#_c_2012_n 0.00151294f $X=5.14 $Y=1.61
+ $X2=0 $Y2=0
cc_951 N_A_834_93#_c_1264_n N_A_415_81#_c_2006_n 0.00472055f $X=6.015 $Y=1.3
+ $X2=0 $Y2=0
cc_952 N_A_834_93#_c_1265_n N_A_415_81#_c_2006_n 0.00543791f $X=6.09 $Y=1.225
+ $X2=0 $Y2=0
cc_953 N_A_834_93#_c_1263_n N_A_415_81#_c_2013_n 0.00686866f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_954 N_A_834_93#_c_1276_n N_A_415_81#_c_2013_n 0.00408184f $X=6.545 $Y=3.15
+ $X2=0 $Y2=0
cc_955 N_A_834_93#_M1012_g N_A_415_81#_c_2013_n 4.5269e-19 $X=6.635 $Y=2.525
+ $X2=0 $Y2=0
cc_956 N_A_834_93#_c_1264_n N_A_415_81#_c_2007_n 0.0123495f $X=6.015 $Y=1.3
+ $X2=0 $Y2=0
cc_957 N_A_834_93#_c_1262_n N_A_415_81#_c_2008_n 9.57758e-19 $X=5.615 $Y=1.595
+ $X2=0 $Y2=0
cc_958 N_A_834_93#_c_1264_n N_A_415_81#_c_2008_n 0.00567123f $X=6.015 $Y=1.3
+ $X2=0 $Y2=0
cc_959 N_A_834_93#_M1012_g N_A_415_81#_c_2014_n 6.92003e-19 $X=6.635 $Y=2.525
+ $X2=0 $Y2=0
cc_960 N_A_834_93#_c_1263_n N_A_415_81#_c_2015_n 0.001267f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_961 N_A_834_93#_c_1262_n N_A_415_81#_c_2009_n 0.00422551f $X=5.615 $Y=1.595
+ $X2=0 $Y2=0
cc_962 N_A_834_93#_c_1290_n N_VGND_M1038_d 0.00733039f $X=4.81 $Y=1.005 $X2=0
+ $Y2=0
cc_963 N_A_834_93#_c_1269_n N_VGND_M1038_d 0.00428317f $X=4.915 $Y=1.445 $X2=0
+ $Y2=0
cc_964 N_A_834_93#_c_1270_n N_VGND_c_2219_n 0.0189707f $X=4.45 $Y=0.625 $X2=0
+ $Y2=0
cc_965 N_A_834_93#_c_1290_n N_VGND_c_2220_n 0.0246763f $X=4.81 $Y=1.005 $X2=0
+ $Y2=0
cc_966 N_A_834_93#_c_1270_n N_VGND_c_2220_n 0.0135218f $X=4.45 $Y=0.625 $X2=0
+ $Y2=0
cc_967 N_A_834_93#_c_1273_n N_VGND_c_2220_n 0.00213166f $X=5.14 $Y=1.41 $X2=0
+ $Y2=0
cc_968 N_A_834_93#_M1036_g N_VGND_c_2221_n 0.00156589f $X=9.7 $Y=0.58 $X2=0
+ $Y2=0
cc_969 N_A_834_93#_c_1270_n N_VGND_c_2227_n 0.00999994f $X=4.45 $Y=0.625 $X2=0
+ $Y2=0
cc_970 N_A_834_93#_M1036_g N_VGND_c_2231_n 0.00320499f $X=9.7 $Y=0.58 $X2=0
+ $Y2=0
cc_971 N_A_834_93#_M1036_g N_VGND_c_2240_n 0.00443186f $X=9.7 $Y=0.58 $X2=0
+ $Y2=0
cc_972 N_A_834_93#_c_1270_n N_VGND_c_2240_n 0.0112422f $X=4.45 $Y=0.625 $X2=0
+ $Y2=0
cc_973 N_A_834_93#_c_1273_n N_VGND_c_2240_n 8.45315e-19 $X=5.14 $Y=1.41 $X2=0
+ $Y2=0
cc_974 N_A_2003_48#_c_1453_n N_A_1745_74#_c_1535_n 0.00593167f $X=11.415 $Y=0.55
+ $X2=0 $Y2=0
cc_975 N_A_2003_48#_c_1454_n N_A_1745_74#_c_1535_n 0.00443992f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_976 N_A_2003_48#_c_1460_n N_A_1745_74#_c_1536_n 0.00843187f $X=11.165 $Y=2.75
+ $X2=0 $Y2=0
cc_977 N_A_2003_48#_c_1458_n N_A_1745_74#_c_1536_n 0.00146716f $X=11.5 $Y=1.47
+ $X2=0 $Y2=0
cc_978 N_A_2003_48#_c_1454_n N_A_1745_74#_c_1537_n 0.00271488f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_979 N_A_2003_48#_c_1458_n N_A_1745_74#_c_1539_n 4.51356e-19 $X=11.5 $Y=1.47
+ $X2=0 $Y2=0
cc_980 N_A_2003_48#_c_1454_n N_A_1745_74#_c_1541_n 0.00311356f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_981 N_A_2003_48#_c_1457_n N_A_1745_74#_c_1541_n 0.00843187f $X=11.165 $Y=2.52
+ $X2=0 $Y2=0
cc_982 N_A_2003_48#_c_1458_n N_A_1745_74#_c_1541_n 0.0149058f $X=11.5 $Y=1.47
+ $X2=0 $Y2=0
cc_983 N_A_2003_48#_M1032_g N_A_1745_74#_c_1567_n 0.00125881f $X=10.09 $Y=0.58
+ $X2=0 $Y2=0
cc_984 N_A_2003_48#_M1010_g N_A_1745_74#_c_1556_n 0.0112947f $X=10.255 $Y=2.75
+ $X2=0 $Y2=0
cc_985 N_A_2003_48#_M1032_g N_A_1745_74#_c_1544_n 9.29499e-19 $X=10.09 $Y=0.58
+ $X2=0 $Y2=0
cc_986 N_A_2003_48#_M1032_g N_A_1745_74#_c_1545_n 0.00223708f $X=10.09 $Y=0.58
+ $X2=0 $Y2=0
cc_987 N_A_2003_48#_M1010_g N_A_1745_74#_c_1545_n 0.00234903f $X=10.255 $Y=2.75
+ $X2=0 $Y2=0
cc_988 N_A_2003_48#_c_1455_n N_A_1745_74#_c_1545_n 0.0167585f $X=10.18 $Y=1.39
+ $X2=0 $Y2=0
cc_989 N_A_2003_48#_M1032_g N_A_1745_74#_c_1546_n 0.0143799f $X=10.09 $Y=0.58
+ $X2=0 $Y2=0
cc_990 N_A_2003_48#_c_1452_n N_A_1745_74#_c_1546_n 0.0259611f $X=11.16 $Y=1.47
+ $X2=0 $Y2=0
cc_991 N_A_2003_48#_c_1455_n N_A_1745_74#_c_1546_n 0.0242156f $X=10.18 $Y=1.39
+ $X2=0 $Y2=0
cc_992 N_A_2003_48#_c_1456_n N_A_1745_74#_c_1546_n 0.001245f $X=10.18 $Y=1.39
+ $X2=0 $Y2=0
cc_993 N_A_2003_48#_M1010_g N_A_1745_74#_c_1558_n 0.00995549f $X=10.255 $Y=2.75
+ $X2=0 $Y2=0
cc_994 N_A_2003_48#_c_1455_n N_A_1745_74#_c_1558_n 0.0210104f $X=10.18 $Y=1.39
+ $X2=0 $Y2=0
cc_995 N_A_2003_48#_c_1456_n N_A_1745_74#_c_1558_n 0.00106876f $X=10.18 $Y=1.39
+ $X2=0 $Y2=0
cc_996 N_A_2003_48#_M1010_g N_A_1745_74#_c_1560_n 0.0194047f $X=10.255 $Y=2.75
+ $X2=0 $Y2=0
cc_997 N_A_2003_48#_c_1452_n N_A_1745_74#_c_1548_n 0.0247317f $X=11.16 $Y=1.47
+ $X2=0 $Y2=0
cc_998 N_A_2003_48#_c_1453_n N_A_1745_74#_c_1548_n 0.014253f $X=11.415 $Y=0.55
+ $X2=0 $Y2=0
cc_999 N_A_2003_48#_c_1454_n N_A_1745_74#_c_1548_n 0.0236842f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_1000 N_A_2003_48#_c_1452_n N_A_1745_74#_c_1549_n 0.0121221f $X=11.16 $Y=1.47
+ $X2=0 $Y2=0
cc_1001 N_A_2003_48#_c_1453_n N_A_1745_74#_c_1549_n 0.00619797f $X=11.415
+ $Y=0.55 $X2=0 $Y2=0
cc_1002 N_A_2003_48#_c_1454_n N_A_1745_74#_c_1549_n 0.0191241f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_1003 N_A_2003_48#_c_1453_n N_A_2339_74#_c_1703_n 0.026931f $X=11.415 $Y=0.55
+ $X2=0 $Y2=0
cc_1004 N_A_2003_48#_c_1454_n N_A_2339_74#_c_1703_n 0.0405862f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_1005 N_A_2003_48#_c_1454_n N_A_2339_74#_c_1705_n 0.00909743f $X=11.5 $Y=1.385
+ $X2=0 $Y2=0
cc_1006 N_A_2003_48#_c_1457_n N_A_2339_74#_c_1705_n 0.00195796f $X=11.165
+ $Y=2.52 $X2=0 $Y2=0
cc_1007 N_A_2003_48#_c_1458_n N_A_2339_74#_c_1705_n 0.0157384f $X=11.5 $Y=1.47
+ $X2=0 $Y2=0
cc_1008 N_A_2003_48#_M1010_g N_VPWR_c_1819_n 0.00907747f $X=10.255 $Y=2.75 $X2=0
+ $Y2=0
cc_1009 N_A_2003_48#_c_1460_n N_VPWR_c_1819_n 0.016245f $X=11.165 $Y=2.75 $X2=0
+ $Y2=0
cc_1010 N_A_2003_48#_c_1457_n N_VPWR_c_1820_n 0.0470961f $X=11.165 $Y=2.52 $X2=0
+ $Y2=0
cc_1011 N_A_2003_48#_M1010_g N_VPWR_c_1828_n 0.00417766f $X=10.255 $Y=2.75 $X2=0
+ $Y2=0
cc_1012 N_A_2003_48#_c_1460_n N_VPWR_c_1833_n 0.0143566f $X=11.165 $Y=2.75 $X2=0
+ $Y2=0
cc_1013 N_A_2003_48#_M1010_g N_VPWR_c_1813_n 0.00627075f $X=10.255 $Y=2.75 $X2=0
+ $Y2=0
cc_1014 N_A_2003_48#_c_1460_n N_VPWR_c_1813_n 0.011899f $X=11.165 $Y=2.75 $X2=0
+ $Y2=0
cc_1015 N_A_2003_48#_M1032_g N_VGND_c_2221_n 0.00986387f $X=10.09 $Y=0.58 $X2=0
+ $Y2=0
cc_1016 N_A_2003_48#_c_1453_n N_VGND_c_2221_n 0.0104724f $X=11.415 $Y=0.55 $X2=0
+ $Y2=0
cc_1017 N_A_2003_48#_M1032_g N_VGND_c_2231_n 0.00383152f $X=10.09 $Y=0.58 $X2=0
+ $Y2=0
cc_1018 N_A_2003_48#_c_1453_n N_VGND_c_2232_n 0.0191719f $X=11.415 $Y=0.55 $X2=0
+ $Y2=0
cc_1019 N_A_2003_48#_M1032_g N_VGND_c_2240_n 0.0075725f $X=10.09 $Y=0.58 $X2=0
+ $Y2=0
cc_1020 N_A_2003_48#_c_1453_n N_VGND_c_2240_n 0.0192149f $X=11.415 $Y=0.55 $X2=0
+ $Y2=0
cc_1021 N_A_1745_74#_c_1538_n N_A_2339_74#_c_1693_n 0.00970941f $X=12.055
+ $Y=1.185 $X2=0 $Y2=0
cc_1022 N_A_1745_74#_c_1540_n N_A_2339_74#_c_1695_n 0.00936026f $X=12.4 $Y=1.69
+ $X2=0 $Y2=0
cc_1023 N_A_1745_74#_c_1543_n N_A_2339_74#_c_1695_n 0.00970941f $X=12.055
+ $Y=1.26 $X2=0 $Y2=0
cc_1024 N_A_1745_74#_c_1540_n N_A_2339_74#_M1015_g 0.021381f $X=12.4 $Y=1.69
+ $X2=0 $Y2=0
cc_1025 N_A_1745_74#_c_1535_n N_A_2339_74#_c_1703_n 5.54394e-19 $X=10.99 $Y=0.9
+ $X2=0 $Y2=0
cc_1026 N_A_1745_74#_c_1537_n N_A_2339_74#_c_1703_n 0.00765913f $X=11.98 $Y=1.26
+ $X2=0 $Y2=0
cc_1027 N_A_1745_74#_c_1538_n N_A_2339_74#_c_1703_n 0.0035045f $X=12.055
+ $Y=1.185 $X2=0 $Y2=0
cc_1028 N_A_1745_74#_c_1549_n N_A_2339_74#_c_1703_n 8.98164e-19 $X=11.535
+ $Y=1.117 $X2=0 $Y2=0
cc_1029 N_A_1745_74#_c_1536_n N_A_2339_74#_c_1704_n 0.00120599f $X=11.475
+ $Y=1.665 $X2=0 $Y2=0
cc_1030 N_A_1745_74#_c_1552_n N_A_2339_74#_c_1704_n 0.0151739f $X=12.04 $Y=1.765
+ $X2=0 $Y2=0
cc_1031 N_A_1745_74#_c_1539_n N_A_2339_74#_c_1704_n 6.63362e-19 $X=12.055
+ $Y=1.615 $X2=0 $Y2=0
cc_1032 N_A_1745_74#_c_1540_n N_A_2339_74#_c_1704_n 0.0129929f $X=12.4 $Y=1.69
+ $X2=0 $Y2=0
cc_1033 N_A_1745_74#_c_1554_n N_A_2339_74#_c_1704_n 0.0151665f $X=12.49 $Y=1.765
+ $X2=0 $Y2=0
cc_1034 N_A_1745_74#_c_1542_n N_A_2339_74#_c_1704_n 0.00313656f $X=12.04 $Y=1.69
+ $X2=0 $Y2=0
cc_1035 N_A_1745_74#_c_1536_n N_A_2339_74#_c_1705_n 2.72834e-19 $X=11.475
+ $Y=1.665 $X2=0 $Y2=0
cc_1036 N_A_1745_74#_c_1537_n N_A_2339_74#_c_1705_n 0.00807224f $X=11.98 $Y=1.26
+ $X2=0 $Y2=0
cc_1037 N_A_1745_74#_c_1539_n N_A_2339_74#_c_1705_n 0.0179017f $X=12.055
+ $Y=1.615 $X2=0 $Y2=0
cc_1038 N_A_1745_74#_c_1540_n N_A_2339_74#_c_1705_n 0.00884608f $X=12.4 $Y=1.69
+ $X2=0 $Y2=0
cc_1039 N_A_1745_74#_c_1541_n N_A_2339_74#_c_1705_n 0.00110135f $X=11.475
+ $Y=1.575 $X2=0 $Y2=0
cc_1040 N_A_1745_74#_c_1542_n N_A_2339_74#_c_1705_n 0.00157693f $X=12.04 $Y=1.69
+ $X2=0 $Y2=0
cc_1041 N_A_1745_74#_c_1543_n N_A_2339_74#_c_1705_n 0.00802343f $X=12.055
+ $Y=1.26 $X2=0 $Y2=0
cc_1042 N_A_1745_74#_c_1539_n N_A_2339_74#_c_1707_n 0.00212764f $X=12.055
+ $Y=1.615 $X2=0 $Y2=0
cc_1043 N_A_1745_74#_c_1556_n N_VPWR_c_1819_n 0.0271932f $X=10.125 $Y=2.715
+ $X2=0 $Y2=0
cc_1044 N_A_1745_74#_c_1560_n N_VPWR_c_1819_n 0.00221607f $X=10.21 $Y=2.55 $X2=0
+ $Y2=0
cc_1045 N_A_1745_74#_M1044_g N_VPWR_c_1820_n 0.0188578f $X=11.475 $Y=2.75 $X2=0
+ $Y2=0
cc_1046 N_A_1745_74#_c_1537_n N_VPWR_c_1820_n 0.00368592f $X=11.98 $Y=1.26 $X2=0
+ $Y2=0
cc_1047 N_A_1745_74#_c_1552_n N_VPWR_c_1820_n 0.00431879f $X=12.04 $Y=1.765
+ $X2=0 $Y2=0
cc_1048 N_A_1745_74#_c_1554_n N_VPWR_c_1821_n 0.00783519f $X=12.49 $Y=1.765
+ $X2=0 $Y2=0
cc_1049 N_A_1745_74#_c_1556_n N_VPWR_c_1828_n 0.02744f $X=10.125 $Y=2.715 $X2=0
+ $Y2=0
cc_1050 N_A_1745_74#_M1044_g N_VPWR_c_1833_n 0.00553757f $X=11.475 $Y=2.75 $X2=0
+ $Y2=0
cc_1051 N_A_1745_74#_c_1552_n N_VPWR_c_1834_n 0.00465228f $X=12.04 $Y=1.765
+ $X2=0 $Y2=0
cc_1052 N_A_1745_74#_c_1554_n N_VPWR_c_1834_n 0.00465228f $X=12.49 $Y=1.765
+ $X2=0 $Y2=0
cc_1053 N_A_1745_74#_M1044_g N_VPWR_c_1813_n 0.0109544f $X=11.475 $Y=2.75 $X2=0
+ $Y2=0
cc_1054 N_A_1745_74#_c_1552_n N_VPWR_c_1813_n 0.00555093f $X=12.04 $Y=1.765
+ $X2=0 $Y2=0
cc_1055 N_A_1745_74#_c_1554_n N_VPWR_c_1813_n 0.00555093f $X=12.49 $Y=1.765
+ $X2=0 $Y2=0
cc_1056 N_A_1745_74#_c_1556_n N_VPWR_c_1813_n 0.0331166f $X=10.125 $Y=2.715
+ $X2=0 $Y2=0
cc_1057 N_A_1745_74#_c_1556_n A_1985_508# 0.00402894f $X=10.125 $Y=2.715
+ $X2=-0.19 $Y2=-0.245
cc_1058 N_A_1745_74#_c_1535_n N_VGND_c_2221_n 0.00154514f $X=10.99 $Y=0.9 $X2=0
+ $Y2=0
cc_1059 N_A_1745_74#_c_1567_n N_VGND_c_2221_n 0.011455f $X=9.585 $Y=0.57 $X2=0
+ $Y2=0
cc_1060 N_A_1745_74#_c_1546_n N_VGND_c_2221_n 0.0267689f $X=10.915 $Y=0.97 $X2=0
+ $Y2=0
cc_1061 N_A_1745_74#_c_1538_n N_VGND_c_2222_n 0.0149682f $X=12.055 $Y=1.185
+ $X2=0 $Y2=0
cc_1062 N_A_1745_74#_c_1567_n N_VGND_c_2231_n 0.0190071f $X=9.585 $Y=0.57 $X2=0
+ $Y2=0
cc_1063 N_A_1745_74#_c_1535_n N_VGND_c_2232_n 0.00433941f $X=10.99 $Y=0.9 $X2=0
+ $Y2=0
cc_1064 N_A_1745_74#_c_1538_n N_VGND_c_2232_n 0.00383152f $X=12.055 $Y=1.185
+ $X2=0 $Y2=0
cc_1065 N_A_1745_74#_c_1535_n N_VGND_c_2240_n 0.00822721f $X=10.99 $Y=0.9 $X2=0
+ $Y2=0
cc_1066 N_A_1745_74#_c_1538_n N_VGND_c_2240_n 0.00762539f $X=12.055 $Y=1.185
+ $X2=0 $Y2=0
cc_1067 N_A_1745_74#_c_1567_n N_VGND_c_2240_n 0.0200126f $X=9.585 $Y=0.57 $X2=0
+ $Y2=0
cc_1068 N_A_2339_74#_c_1704_n N_VPWR_c_1820_n 0.030344f $X=12.265 $Y=1.985 $X2=0
+ $Y2=0
cc_1069 N_A_2339_74#_c_1705_n N_VPWR_c_1820_n 0.0106252f $X=12.43 $Y=1.435 $X2=0
+ $Y2=0
cc_1070 N_A_2339_74#_c_1694_n N_VPWR_c_1821_n 9.84896e-19 $X=12.84 $Y=1.3 $X2=0
+ $Y2=0
cc_1071 N_A_2339_74#_M1015_g N_VPWR_c_1821_n 0.00546744f $X=13.025 $Y=2.4 $X2=0
+ $Y2=0
cc_1072 N_A_2339_74#_c_1704_n N_VPWR_c_1821_n 0.0297549f $X=12.265 $Y=1.985
+ $X2=0 $Y2=0
cc_1073 N_A_2339_74#_c_1706_n N_VPWR_c_1821_n 0.0181117f $X=13.685 $Y=1.435
+ $X2=0 $Y2=0
cc_1074 N_A_2339_74#_c_1707_n N_VPWR_c_1821_n 0.00116289f $X=14.375 $Y=1.412
+ $X2=0 $Y2=0
cc_1075 N_A_2339_74#_M1015_g N_VPWR_c_1822_n 0.005209f $X=13.025 $Y=2.4 $X2=0
+ $Y2=0
cc_1076 N_A_2339_74#_M1019_g N_VPWR_c_1822_n 0.005209f $X=13.475 $Y=2.4 $X2=0
+ $Y2=0
cc_1077 N_A_2339_74#_M1019_g N_VPWR_c_1823_n 0.00362296f $X=13.475 $Y=2.4 $X2=0
+ $Y2=0
cc_1078 N_A_2339_74#_M1023_g N_VPWR_c_1823_n 0.0159323f $X=13.925 $Y=2.4 $X2=0
+ $Y2=0
cc_1079 N_A_2339_74#_M1029_g N_VPWR_c_1823_n 6.05118e-19 $X=14.375 $Y=2.4 $X2=0
+ $Y2=0
cc_1080 N_A_2339_74#_M1029_g N_VPWR_c_1825_n 0.00708612f $X=14.375 $Y=2.4 $X2=0
+ $Y2=0
cc_1081 N_A_2339_74#_c_1704_n N_VPWR_c_1834_n 0.00657675f $X=12.265 $Y=1.985
+ $X2=0 $Y2=0
cc_1082 N_A_2339_74#_M1023_g N_VPWR_c_1835_n 0.00460063f $X=13.925 $Y=2.4 $X2=0
+ $Y2=0
cc_1083 N_A_2339_74#_M1029_g N_VPWR_c_1835_n 0.00553757f $X=14.375 $Y=2.4 $X2=0
+ $Y2=0
cc_1084 N_A_2339_74#_M1015_g N_VPWR_c_1813_n 0.00987399f $X=13.025 $Y=2.4 $X2=0
+ $Y2=0
cc_1085 N_A_2339_74#_M1019_g N_VPWR_c_1813_n 0.00982266f $X=13.475 $Y=2.4 $X2=0
+ $Y2=0
cc_1086 N_A_2339_74#_M1023_g N_VPWR_c_1813_n 0.00908554f $X=13.925 $Y=2.4 $X2=0
+ $Y2=0
cc_1087 N_A_2339_74#_M1029_g N_VPWR_c_1813_n 0.0109139f $X=14.375 $Y=2.4 $X2=0
+ $Y2=0
cc_1088 N_A_2339_74#_c_1704_n N_VPWR_c_1813_n 0.00992028f $X=12.265 $Y=1.985
+ $X2=0 $Y2=0
cc_1089 N_A_2339_74#_c_1693_n N_Q_c_2150_n 0.00667713f $X=12.485 $Y=1.225 $X2=0
+ $Y2=0
cc_1090 N_A_2339_74#_c_1696_n N_Q_c_2150_n 0.0125407f $X=12.915 $Y=1.225 $X2=0
+ $Y2=0
cc_1091 N_A_2339_74#_c_1696_n N_Q_c_2161_n 0.0131906f $X=12.915 $Y=1.225 $X2=0
+ $Y2=0
cc_1092 N_A_2339_74#_c_1700_n N_Q_c_2161_n 0.0164669f $X=13.955 $Y=1.225 $X2=0
+ $Y2=0
cc_1093 N_A_2339_74#_c_1706_n N_Q_c_2161_n 0.0693421f $X=13.685 $Y=1.435 $X2=0
+ $Y2=0
cc_1094 N_A_2339_74#_c_1707_n N_Q_c_2161_n 0.0190905f $X=14.375 $Y=1.412 $X2=0
+ $Y2=0
cc_1095 N_A_2339_74#_c_1693_n N_Q_c_2165_n 0.00205797f $X=12.485 $Y=1.225 $X2=0
+ $Y2=0
cc_1096 N_A_2339_74#_c_1694_n N_Q_c_2165_n 0.00210982f $X=12.84 $Y=1.3 $X2=0
+ $Y2=0
cc_1097 N_A_2339_74#_c_1696_n N_Q_c_2165_n 7.32094e-19 $X=12.915 $Y=1.225 $X2=0
+ $Y2=0
cc_1098 N_A_2339_74#_c_1706_n N_Q_c_2165_n 0.0218379f $X=13.685 $Y=1.435 $X2=0
+ $Y2=0
cc_1099 N_A_2339_74#_M1015_g N_Q_c_2154_n 0.0136771f $X=13.025 $Y=2.4 $X2=0
+ $Y2=0
cc_1100 N_A_2339_74#_M1019_g N_Q_c_2154_n 0.0148573f $X=13.475 $Y=2.4 $X2=0
+ $Y2=0
cc_1101 N_A_2339_74#_M1023_g N_Q_c_2154_n 7.9417e-19 $X=13.925 $Y=2.4 $X2=0
+ $Y2=0
cc_1102 N_A_2339_74#_M1019_g N_Q_c_2155_n 0.012931f $X=13.475 $Y=2.4 $X2=0 $Y2=0
cc_1103 N_A_2339_74#_M1023_g N_Q_c_2155_n 0.0174957f $X=13.925 $Y=2.4 $X2=0
+ $Y2=0
cc_1104 N_A_2339_74#_c_1706_n N_Q_c_2155_n 0.0320444f $X=13.685 $Y=1.435 $X2=0
+ $Y2=0
cc_1105 N_A_2339_74#_c_1707_n N_Q_c_2155_n 0.00207172f $X=14.375 $Y=1.412 $X2=0
+ $Y2=0
cc_1106 N_A_2339_74#_M1015_g N_Q_c_2156_n 0.00373763f $X=13.025 $Y=2.4 $X2=0
+ $Y2=0
cc_1107 N_A_2339_74#_M1019_g N_Q_c_2156_n 0.00170419f $X=13.475 $Y=2.4 $X2=0
+ $Y2=0
cc_1108 N_A_2339_74#_c_1704_n N_Q_c_2156_n 0.00129088f $X=12.265 $Y=1.985 $X2=0
+ $Y2=0
cc_1109 N_A_2339_74#_c_1706_n N_Q_c_2156_n 0.0275631f $X=13.685 $Y=1.435 $X2=0
+ $Y2=0
cc_1110 N_A_2339_74#_c_1707_n N_Q_c_2156_n 0.00215053f $X=14.375 $Y=1.412 $X2=0
+ $Y2=0
cc_1111 N_A_2339_74#_M1023_g N_Q_c_2157_n 3.6581e-19 $X=13.925 $Y=2.4 $X2=0
+ $Y2=0
cc_1112 N_A_2339_74#_M1029_g N_Q_c_2157_n 3.99037e-19 $X=14.375 $Y=2.4 $X2=0
+ $Y2=0
cc_1113 N_A_2339_74#_c_1700_n N_Q_c_2151_n 3.92031e-19 $X=13.955 $Y=1.225 $X2=0
+ $Y2=0
cc_1114 N_A_2339_74#_c_1702_n N_Q_c_2151_n 3.92313e-19 $X=14.385 $Y=1.225 $X2=0
+ $Y2=0
cc_1115 N_A_2339_74#_c_1700_n N_Q_c_2152_n 0.00272065f $X=13.955 $Y=1.225 $X2=0
+ $Y2=0
cc_1116 N_A_2339_74#_c_1702_n N_Q_c_2152_n 0.00240279f $X=14.385 $Y=1.225 $X2=0
+ $Y2=0
cc_1117 N_A_2339_74#_c_1706_n N_Q_c_2152_n 0.00167694f $X=13.685 $Y=1.435 $X2=0
+ $Y2=0
cc_1118 N_A_2339_74#_c_1707_n N_Q_c_2152_n 0.00902935f $X=14.375 $Y=1.412 $X2=0
+ $Y2=0
cc_1119 N_A_2339_74#_M1023_g Q 0.00520905f $X=13.925 $Y=2.4 $X2=0 $Y2=0
cc_1120 N_A_2339_74#_M1029_g Q 0.0239402f $X=14.375 $Y=2.4 $X2=0 $Y2=0
cc_1121 N_A_2339_74#_c_1706_n Q 0.0194661f $X=13.685 $Y=1.435 $X2=0 $Y2=0
cc_1122 N_A_2339_74#_c_1707_n Q 0.0338078f $X=14.375 $Y=1.412 $X2=0 $Y2=0
cc_1123 N_A_2339_74#_c_1693_n N_VGND_c_2222_n 0.00182441f $X=12.485 $Y=1.225
+ $X2=0 $Y2=0
cc_1124 N_A_2339_74#_c_1703_n N_VGND_c_2222_n 0.0266033f $X=11.84 $Y=0.515 $X2=0
+ $Y2=0
cc_1125 N_A_2339_74#_c_1705_n N_VGND_c_2222_n 0.0191073f $X=12.43 $Y=1.435 $X2=0
+ $Y2=0
cc_1126 N_A_2339_74#_c_1700_n N_VGND_c_2224_n 4.98647e-19 $X=13.955 $Y=1.225
+ $X2=0 $Y2=0
cc_1127 N_A_2339_74#_c_1702_n N_VGND_c_2224_n 0.0149937f $X=14.385 $Y=1.225
+ $X2=0 $Y2=0
cc_1128 N_A_2339_74#_c_1703_n N_VGND_c_2232_n 0.00749631f $X=11.84 $Y=0.515
+ $X2=0 $Y2=0
cc_1129 N_A_2339_74#_c_1700_n N_VGND_c_2233_n 0.00383152f $X=13.955 $Y=1.225
+ $X2=0 $Y2=0
cc_1130 N_A_2339_74#_c_1702_n N_VGND_c_2233_n 0.00383152f $X=14.385 $Y=1.225
+ $X2=0 $Y2=0
cc_1131 N_A_2339_74#_c_1693_n N_VGND_c_2238_n 0.00434272f $X=12.485 $Y=1.225
+ $X2=0 $Y2=0
cc_1132 N_A_2339_74#_c_1696_n N_VGND_c_2238_n 0.00434272f $X=12.915 $Y=1.225
+ $X2=0 $Y2=0
cc_1133 N_A_2339_74#_c_1696_n N_VGND_c_2239_n 0.00452683f $X=12.915 $Y=1.225
+ $X2=0 $Y2=0
cc_1134 N_A_2339_74#_c_1700_n N_VGND_c_2239_n 0.0108787f $X=13.955 $Y=1.225
+ $X2=0 $Y2=0
cc_1135 N_A_2339_74#_c_1702_n N_VGND_c_2239_n 4.44374e-19 $X=14.385 $Y=1.225
+ $X2=0 $Y2=0
cc_1136 N_A_2339_74#_c_1693_n N_VGND_c_2240_n 0.00820158f $X=12.485 $Y=1.225
+ $X2=0 $Y2=0
cc_1137 N_A_2339_74#_c_1696_n N_VGND_c_2240_n 0.00825037f $X=12.915 $Y=1.225
+ $X2=0 $Y2=0
cc_1138 N_A_2339_74#_c_1700_n N_VGND_c_2240_n 0.00752925f $X=13.955 $Y=1.225
+ $X2=0 $Y2=0
cc_1139 N_A_2339_74#_c_1702_n N_VGND_c_2240_n 0.0075754f $X=14.385 $Y=1.225
+ $X2=0 $Y2=0
cc_1140 N_A_2339_74#_c_1703_n N_VGND_c_2240_n 0.0062048f $X=11.84 $Y=0.515 $X2=0
+ $Y2=0
cc_1141 N_VPWR_M1043_d N_A_415_81#_c_2019_n 0.00992117f $X=3.145 $Y=2.32 $X2=0
+ $Y2=0
cc_1142 N_VPWR_c_1814_n N_A_415_81#_c_2019_n 0.0223155f $X=3.285 $Y=2.79 $X2=0
+ $Y2=0
cc_1143 N_VPWR_c_1813_n N_A_415_81#_c_2019_n 0.0224686f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1144 N_VPWR_M1043_d N_A_415_81#_c_2005_n 3.08638e-19 $X=3.145 $Y=2.32 $X2=0
+ $Y2=0
cc_1145 N_VPWR_M1026_d N_A_415_81#_c_2012_n 0.00357274f $X=4.735 $Y=1.935 $X2=0
+ $Y2=0
cc_1146 N_VPWR_c_1815_n N_A_415_81#_c_2012_n 0.0162809f $X=4.87 $Y=2.88 $X2=0
+ $Y2=0
cc_1147 N_VPWR_c_1826_n N_A_415_81#_c_2012_n 0.0099286f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1148 N_VPWR_c_1832_n N_A_415_81#_c_2012_n 0.0112649f $X=7.17 $Y=3.33 $X2=0
+ $Y2=0
cc_1149 N_VPWR_c_1813_n N_A_415_81#_c_2012_n 0.0384554f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1150 N_VPWR_c_1832_n N_A_415_81#_c_2013_n 0.00451006f $X=7.17 $Y=3.33 $X2=0
+ $Y2=0
cc_1151 N_VPWR_c_1813_n N_A_415_81#_c_2013_n 0.00670405f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1152 N_VPWR_c_1814_n N_A_415_81#_c_2017_n 0.00705091f $X=3.285 $Y=2.79 $X2=0
+ $Y2=0
cc_1153 N_VPWR_c_1831_n N_A_415_81#_c_2017_n 0.0143725f $X=3.095 $Y=3.33 $X2=0
+ $Y2=0
cc_1154 N_VPWR_c_1836_n N_A_415_81#_c_2017_n 0.0198328f $X=1.4 $Y=2.465 $X2=0
+ $Y2=0
cc_1155 N_VPWR_c_1813_n N_A_415_81#_c_2017_n 0.0118007f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1156 N_VPWR_M1043_d N_A_415_81#_c_2018_n 6.73969e-19 $X=3.145 $Y=2.32 $X2=0
+ $Y2=0
cc_1157 N_VPWR_c_1814_n N_A_415_81#_c_2018_n 0.0290477f $X=3.285 $Y=2.79 $X2=0
+ $Y2=0
cc_1158 N_VPWR_c_1826_n N_A_415_81#_c_2018_n 0.0250854f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1159 N_VPWR_c_1813_n N_A_415_81#_c_2018_n 0.0211025f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1160 N_VPWR_c_1821_n N_Q_c_2154_n 0.0349062f $X=12.8 $Y=1.985 $X2=0 $Y2=0
cc_1161 N_VPWR_c_1822_n N_Q_c_2154_n 0.0144623f $X=13.615 $Y=3.33 $X2=0 $Y2=0
cc_1162 N_VPWR_c_1823_n N_Q_c_2154_n 0.0293385f $X=13.7 $Y=2.275 $X2=0 $Y2=0
cc_1163 N_VPWR_c_1813_n N_Q_c_2154_n 0.0118344f $X=14.64 $Y=3.33 $X2=0 $Y2=0
cc_1164 N_VPWR_M1019_s N_Q_c_2155_n 0.00165831f $X=13.565 $Y=1.84 $X2=0 $Y2=0
cc_1165 N_VPWR_c_1823_n N_Q_c_2155_n 0.0148589f $X=13.7 $Y=2.275 $X2=0 $Y2=0
cc_1166 N_VPWR_c_1821_n N_Q_c_2156_n 0.00511344f $X=12.8 $Y=1.985 $X2=0 $Y2=0
cc_1167 N_VPWR_c_1823_n N_Q_c_2157_n 0.0281293f $X=13.7 $Y=2.275 $X2=0 $Y2=0
cc_1168 N_VPWR_c_1825_n N_Q_c_2157_n 0.00140346f $X=14.6 $Y=2.275 $X2=0 $Y2=0
cc_1169 N_VPWR_c_1835_n N_Q_c_2157_n 0.00950426f $X=14.47 $Y=3.33 $X2=0 $Y2=0
cc_1170 N_VPWR_c_1813_n N_Q_c_2157_n 0.0078668f $X=14.64 $Y=3.33 $X2=0 $Y2=0
cc_1171 N_VPWR_M1029_s Q 0.00301672f $X=14.465 $Y=1.84 $X2=0 $Y2=0
cc_1172 N_VPWR_c_1825_n Q 0.0209488f $X=14.6 $Y=2.275 $X2=0 $Y2=0
cc_1173 N_A_415_81#_c_2019_n A_517_464# 0.0136292f $X=3.445 $Y=2.43 $X2=-0.19
+ $Y2=-0.245
cc_1174 N_A_415_81#_M1008_d N_noxref_24_c_2363_n 0.00984601f $X=2.075 $Y=0.405
+ $X2=0 $Y2=0
cc_1175 N_A_415_81#_c_2004_n N_noxref_24_c_2363_n 0.0108077f $X=3.445 $Y=1.005
+ $X2=0 $Y2=0
cc_1176 N_A_415_81#_c_2010_n N_noxref_24_c_2363_n 0.0251405f $X=2.485 $Y=0.68
+ $X2=0 $Y2=0
cc_1177 N_A_415_81#_c_2004_n N_noxref_24_c_2365_n 0.0219315f $X=3.445 $Y=1.005
+ $X2=0 $Y2=0
cc_1178 N_Q_c_2161_n N_VGND_M1020_d 0.019527f $X=14.085 $Y=1.015 $X2=0 $Y2=0
cc_1179 N_Q_c_2150_n N_VGND_c_2222_n 0.0224879f $X=12.7 $Y=0.515 $X2=0 $Y2=0
cc_1180 N_Q_c_2151_n N_VGND_c_2224_n 0.0214745f $X=14.17 $Y=0.515 $X2=0 $Y2=0
cc_1181 N_Q_c_2152_n N_VGND_c_2224_n 0.00176181f $X=14.17 $Y=1.3 $X2=0 $Y2=0
cc_1182 Q N_VGND_c_2224_n 0.0295377f $X=14.555 $Y=1.58 $X2=0 $Y2=0
cc_1183 N_Q_c_2151_n N_VGND_c_2233_n 0.00749631f $X=14.17 $Y=0.515 $X2=0 $Y2=0
cc_1184 N_Q_c_2150_n N_VGND_c_2238_n 0.0144922f $X=12.7 $Y=0.515 $X2=0 $Y2=0
cc_1185 N_Q_c_2150_n N_VGND_c_2239_n 0.0163053f $X=12.7 $Y=0.515 $X2=0 $Y2=0
cc_1186 N_Q_c_2161_n N_VGND_c_2239_n 0.0647108f $X=14.085 $Y=1.015 $X2=0 $Y2=0
cc_1187 N_Q_c_2151_n N_VGND_c_2239_n 0.0171417f $X=14.17 $Y=0.515 $X2=0 $Y2=0
cc_1188 N_Q_c_2150_n N_VGND_c_2240_n 0.0118826f $X=12.7 $Y=0.515 $X2=0 $Y2=0
cc_1189 N_Q_c_2151_n N_VGND_c_2240_n 0.0062048f $X=14.17 $Y=0.515 $X2=0 $Y2=0
cc_1190 N_VGND_c_2225_n N_noxref_24_c_2363_n 0.109833f $X=3.64 $Y=0 $X2=0 $Y2=0
cc_1191 N_VGND_c_2240_n N_noxref_24_c_2363_n 0.0641043f $X=14.64 $Y=0 $X2=0
+ $Y2=0
cc_1192 N_VGND_c_2218_n N_noxref_24_c_2364_n 0.0259561f $X=0.71 $Y=0.555 $X2=0
+ $Y2=0
cc_1193 N_VGND_c_2225_n N_noxref_24_c_2364_n 0.0225398f $X=3.64 $Y=0 $X2=0 $Y2=0
cc_1194 N_VGND_c_2240_n N_noxref_24_c_2364_n 0.0125704f $X=14.64 $Y=0 $X2=0
+ $Y2=0
cc_1195 N_VGND_c_2219_n N_noxref_24_c_2365_n 0.024649f $X=3.775 $Y=0.585 $X2=0
+ $Y2=0
cc_1196 N_VGND_c_2225_n N_noxref_24_c_2365_n 0.0229461f $X=3.64 $Y=0 $X2=0 $Y2=0
cc_1197 N_VGND_c_2240_n N_noxref_24_c_2365_n 0.0126298f $X=14.64 $Y=0 $X2=0
+ $Y2=0
cc_1198 N_noxref_24_c_2363_n noxref_25 0.00373495f $X=3.14 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1199 N_noxref_24_c_2363_n noxref_26 0.0017247f $X=3.14 $Y=0.34 $X2=-0.19
+ $Y2=-0.245

* File: sky130_fd_sc_ms__clkbuf_1.pxi.spice
* Created: Fri Aug 28 17:17:23 2020
* 
x_PM_SKY130_FD_SC_MS__CLKBUF_1%A N_A_M1003_g N_A_M1001_g A A N_A_c_41_n
+ PM_SKY130_FD_SC_MS__CLKBUF_1%A
x_PM_SKY130_FD_SC_MS__CLKBUF_1%A_27_74# N_A_27_74#_M1003_s N_A_27_74#_M1001_s
+ N_A_27_74#_c_73_n N_A_27_74#_M1000_g N_A_27_74#_M1002_g N_A_27_74#_c_76_n
+ N_A_27_74#_c_77_n N_A_27_74#_c_86_n N_A_27_74#_c_87_n N_A_27_74#_c_78_n
+ N_A_27_74#_c_79_n N_A_27_74#_c_103_n N_A_27_74#_c_80_n N_A_27_74#_c_81_n
+ N_A_27_74#_c_82_n N_A_27_74#_c_83_n N_A_27_74#_c_84_n
+ PM_SKY130_FD_SC_MS__CLKBUF_1%A_27_74#
x_PM_SKY130_FD_SC_MS__CLKBUF_1%VPWR N_VPWR_M1001_d N_VPWR_c_143_n N_VPWR_c_144_n
+ N_VPWR_c_145_n VPWR N_VPWR_c_146_n N_VPWR_c_142_n
+ PM_SKY130_FD_SC_MS__CLKBUF_1%VPWR
x_PM_SKY130_FD_SC_MS__CLKBUF_1%X N_X_M1002_d N_X_M1000_d X X X X X X X
+ N_X_c_168_n X PM_SKY130_FD_SC_MS__CLKBUF_1%X
x_PM_SKY130_FD_SC_MS__CLKBUF_1%VGND N_VGND_M1003_d VGND N_VGND_c_188_n
+ N_VGND_c_189_n N_VGND_c_190_n N_VGND_c_191_n PM_SKY130_FD_SC_MS__CLKBUF_1%VGND
cc_1 VNB N_A_M1003_g 0.0571724f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_2 VNB N_A_M1001_g 0.00186696f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=2.4
cc_3 VNB A 0.0173576f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_A_c_41_n 0.0635892f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.465
cc_5 VNB N_A_27_74#_c_73_n 0.0201001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_27_74#_M1000_g 0.00185623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_74#_M1002_g 0.029877f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.465
cc_8 VNB N_A_27_74#_c_76_n 0.0247105f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.465
cc_9 VNB N_A_27_74#_c_77_n 0.0264663f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.54
cc_10 VNB N_A_27_74#_c_78_n 0.0140881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_74#_c_79_n 0.00998406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_c_80_n 0.00523802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_81_n 0.00307467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_74#_c_82_n 3.97508e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_74#_c_83_n 0.0276446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_74#_c_84_n 0.0021899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_VPWR_c_142_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB X 0.0197233f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=2.4
cc_19 VNB X 0.0435818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_188_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_21 VNB N_VGND_c_189_n 0.137744f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_190_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_191_n 0.0270139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VPB N_A_M1001_g 0.0302784f $X=-0.19 $Y=1.66 $X2=0.735 $Y2=2.4
cc_25 VPB A 0.017159f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_26 VPB N_A_27_74#_M1000_g 0.0287814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_27 VPB N_A_27_74#_c_86_n 0.00718233f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_28 VPB N_A_27_74#_c_87_n 0.0352562f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.54
cc_29 VPB N_A_27_74#_c_82_n 0.00282165f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_143_n 0.00969617f $X=-0.19 $Y=1.66 $X2=0.735 $Y2=2.4
cc_31 VPB N_VPWR_c_144_n 0.0264706f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_32 VPB N_VPWR_c_145_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_33 VPB N_VPWR_c_146_n 0.0222728f $X=-0.19 $Y=1.66 $X2=0.735 $Y2=1.465
cc_34 VPB N_VPWR_c_142_n 0.0623715f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB X 0.00835129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB X 0.0449323f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_X_c_168_n 0.01426f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 A N_A_27_74#_c_73_n 0.00110703f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_39 N_A_c_41_n N_A_27_74#_c_73_n 0.018224f $X=0.735 $Y=1.465 $X2=0 $Y2=0
cc_40 N_A_M1001_g N_A_27_74#_M1000_g 0.0202386f $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_41 N_A_M1003_g N_A_27_74#_c_77_n 0.0203098f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_42 N_A_M1001_g N_A_27_74#_c_86_n 8.84614e-19 $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_43 A N_A_27_74#_c_86_n 0.0266342f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_44 N_A_c_41_n N_A_27_74#_c_86_n 0.00152012f $X=0.735 $Y=1.465 $X2=0 $Y2=0
cc_45 N_A_M1001_g N_A_27_74#_c_87_n 0.0120821f $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_46 N_A_M1003_g N_A_27_74#_c_78_n 0.0120783f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_47 A N_A_27_74#_c_78_n 0.0297157f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_48 N_A_c_41_n N_A_27_74#_c_78_n 0.00642643f $X=0.735 $Y=1.465 $X2=0 $Y2=0
cc_49 N_A_M1003_g N_A_27_74#_c_79_n 0.00419718f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_50 A N_A_27_74#_c_79_n 0.0277157f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_51 N_A_c_41_n N_A_27_74#_c_79_n 0.00617335f $X=0.735 $Y=1.465 $X2=0 $Y2=0
cc_52 N_A_M1001_g N_A_27_74#_c_103_n 0.0131848f $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_53 A N_A_27_74#_c_103_n 0.0114506f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_54 N_A_M1003_g N_A_27_74#_c_81_n 0.003256f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_55 A N_A_27_74#_c_81_n 0.0420921f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_56 N_A_c_41_n N_A_27_74#_c_81_n 8.01114e-19 $X=0.735 $Y=1.465 $X2=0 $Y2=0
cc_57 N_A_M1001_g N_A_27_74#_c_82_n 0.00366213f $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_58 N_A_M1003_g N_A_27_74#_c_83_n 0.00658075f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_59 N_A_M1001_g N_A_27_74#_c_84_n 8.01114e-19 $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_60 N_A_M1001_g N_VPWR_c_143_n 0.00343717f $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_61 N_A_M1001_g N_VPWR_c_144_n 0.005209f $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_62 N_A_M1001_g N_VPWR_c_142_n 0.00986895f $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_63 N_A_M1001_g X 6.0115e-19 $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_64 N_A_M1003_g N_VGND_c_189_n 0.00828694f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_65 N_A_M1003_g N_VGND_c_190_n 0.00434272f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_66 N_A_M1003_g N_VGND_c_191_n 0.0115577f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_67 N_A_27_74#_c_103_n N_VPWR_M1001_d 0.00866408f $X=1.005 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_68 N_A_27_74#_c_82_n N_VPWR_M1001_d 0.00206918f $X=1.09 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_69 N_A_27_74#_M1000_g N_VPWR_c_143_n 0.00343717f $X=1.285 $Y=2.4 $X2=0 $Y2=0
cc_70 N_A_27_74#_c_76_n N_VPWR_c_143_n 2.80311e-19 $X=1.282 $Y=1.63 $X2=0 $Y2=0
cc_71 N_A_27_74#_c_87_n N_VPWR_c_143_n 0.0266809f $X=0.51 $Y=2.815 $X2=0 $Y2=0
cc_72 N_A_27_74#_c_103_n N_VPWR_c_143_n 0.0219171f $X=1.005 $Y=2.035 $X2=0 $Y2=0
cc_73 N_A_27_74#_c_87_n N_VPWR_c_144_n 0.014549f $X=0.51 $Y=2.815 $X2=0 $Y2=0
cc_74 N_A_27_74#_M1000_g N_VPWR_c_146_n 0.005209f $X=1.285 $Y=2.4 $X2=0 $Y2=0
cc_75 N_A_27_74#_M1000_g N_VPWR_c_142_n 0.00986692f $X=1.285 $Y=2.4 $X2=0 $Y2=0
cc_76 N_A_27_74#_c_87_n N_VPWR_c_142_n 0.0119743f $X=0.51 $Y=2.815 $X2=0 $Y2=0
cc_77 N_A_27_74#_M1002_g X 0.010743f $X=1.425 $Y=0.58 $X2=0 $Y2=0
cc_78 N_A_27_74#_M1000_g X 0.00416426f $X=1.285 $Y=2.4 $X2=0 $Y2=0
cc_79 N_A_27_74#_M1002_g X 0.0248648f $X=1.425 $Y=0.58 $X2=0 $Y2=0
cc_80 N_A_27_74#_c_80_n X 0.0139294f $X=1.2 $Y=1.13 $X2=0 $Y2=0
cc_81 N_A_27_74#_c_81_n X 0.0389168f $X=1.2 $Y=1.435 $X2=0 $Y2=0
cc_82 N_A_27_74#_c_82_n X 0.00819752f $X=1.09 $Y=1.95 $X2=0 $Y2=0
cc_83 N_A_27_74#_M1000_g X 0.0140042f $X=1.285 $Y=2.4 $X2=0 $Y2=0
cc_84 N_A_27_74#_c_87_n X 0.00414522f $X=0.51 $Y=2.815 $X2=0 $Y2=0
cc_85 N_A_27_74#_M1000_g N_X_c_168_n 0.0034591f $X=1.285 $Y=2.4 $X2=0 $Y2=0
cc_86 N_A_27_74#_c_76_n N_X_c_168_n 0.00516595f $X=1.282 $Y=1.63 $X2=0 $Y2=0
cc_87 N_A_27_74#_c_82_n N_X_c_168_n 0.00584696f $X=1.09 $Y=1.95 $X2=0 $Y2=0
cc_88 N_A_27_74#_c_84_n N_X_c_168_n 0.00379591f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_89 N_A_27_74#_M1002_g N_VGND_c_188_n 0.00434272f $X=1.425 $Y=0.58 $X2=0 $Y2=0
cc_90 N_A_27_74#_M1002_g N_VGND_c_189_n 0.00828694f $X=1.425 $Y=0.58 $X2=0 $Y2=0
cc_91 N_A_27_74#_c_77_n N_VGND_c_189_n 0.0119984f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_92 N_A_27_74#_c_77_n N_VGND_c_190_n 0.0145639f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_93 N_A_27_74#_M1002_g N_VGND_c_191_n 0.0115577f $X=1.425 $Y=0.58 $X2=0 $Y2=0
cc_94 N_A_27_74#_c_77_n N_VGND_c_191_n 0.0132912f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_95 N_A_27_74#_c_78_n N_VGND_c_191_n 0.0220577f $X=1.005 $Y=1.045 $X2=0 $Y2=0
cc_96 N_A_27_74#_c_80_n N_VGND_c_191_n 0.0176776f $X=1.2 $Y=1.13 $X2=0 $Y2=0
cc_97 N_A_27_74#_c_83_n N_VGND_c_191_n 0.00172432f $X=1.23 $Y=1.125 $X2=0 $Y2=0
cc_98 N_VPWR_c_143_n X 0.0280302f $X=1.01 $Y=2.455 $X2=0 $Y2=0
cc_99 N_VPWR_c_146_n X 0.0203497f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_100 N_VPWR_c_142_n X 0.0167756f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_101 X N_VGND_c_188_n 0.0144458f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_102 X N_VGND_c_189_n 0.0119518f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_103 X N_VGND_c_191_n 0.0132912f $X=1.595 $Y=0.47 $X2=0 $Y2=0

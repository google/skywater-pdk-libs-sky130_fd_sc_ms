* File: sky130_fd_sc_ms__sdfstp_1.spice
* Created: Fri Aug 28 18:13:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdfstp_1.pex.spice"
.subckt sky130_fd_sc_ms__sdfstp_1  VNB VPB SCE D SCD CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1025 N_VGND_M1025_d N_SCE_M1025_g N_A_27_464#_M1025_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0819 AS=0.1197 PD=0.81 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1003 A_238_74# N_A_27_464#_M1003_g N_VGND_M1025_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0819 PD=0.66 PS=0.81 NRD=18.564 NRS=11.424 M=1 R=2.8 SA=75000.7
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1034 N_A_292_464#_M1034_d N_D_M1034_g A_238_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1005 A_402_74# N_SCE_M1005_g N_A_292_464#_M1034_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_SCD_M1004_g A_402_74# VNB NLOWVT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_CLK_M1006_g N_A_599_74#_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.2109 PD=1.16 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1015 N_A_800_74#_M1015_d N_A_599_74#_M1015_g N_VGND_M1006_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1014 N_A_998_81#_M1014_d N_A_599_74#_M1014_g N_A_292_464#_M1014_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1281 AS=0.1197 PD=1.03 PS=1.41 NRD=94.284 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1011 A_1150_81# N_A_800_74#_M1011_g N_A_998_81#_M1014_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.1281 PD=0.66 PS=1.03 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_1198_55#_M1009_g A_1150_81# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1032 A_1426_118# N_A_998_81#_M1032_g N_A_1198_55#_M1032_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_SET_B_M1012_g A_1426_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.186187 AS=0.0504 PD=1.10943 PS=0.66 NRD=12.132 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1000 A_1686_74# N_A_998_81#_M1000_g N_VGND_M1012_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.283713 PD=0.88 PS=1.69057 NRD=12.18 NRS=0 M=1 R=4.26667
+ SA=75001.2 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1001 N_A_1764_74#_M1001_d N_A_800_74#_M1001_g A_1686_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.214158 AS=0.0768 PD=1.47321 PS=0.88 NRD=20.616 NRS=12.18 M=1
+ R=4.26667 SA=75001.6 SB=75002 A=0.096 P=1.58 MULT=1
MM1037 A_1910_74# N_A_599_74#_M1037_g N_A_1764_74#_M1001_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.140542 PD=0.66 PS=0.966792 NRD=18.564 NRS=54.996 M=1
+ R=2.8 SA=75002.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1008 A_1988_74# N_A_1958_48#_M1008_g A_1910_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1596 AS=0.0504 PD=1.18 PS=0.66 NRD=92.856 NRS=18.564 M=1 R=2.8 SA=75002.5
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_SET_B_M1022_g A_1988_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0882 AS=0.1596 PD=0.84 PS=1.18 NRD=0 NRS=92.856 M=1 R=2.8 SA=75003.5
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1039 N_A_1958_48#_M1039_d N_A_1764_74#_M1039_g N_VGND_M1022_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1197 AS=0.0882 PD=1.41 PS=0.84 NRD=0 NRS=39.996 M=1 R=2.8
+ SA=75004 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1036 N_VGND_M1036_d N_A_1764_74#_M1036_g N_A_2395_112#_M1036_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.129591 AS=0.385 PD=0.997674 PS=2.5 NRD=18 NRS=140.724 M=1
+ R=3.66667 SA=75000.6 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1023 N_Q_M1023_d N_A_2395_112#_M1023_g N_VGND_M1036_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1017 N_VPWR_M1017_d N_SCE_M1017_g N_A_27_464#_M1017_s VPB PSHORT L=0.18 W=0.64
+ AD=0.0864 AS=0.176 PD=0.91 PS=1.83 NRD=0 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90002.2 A=0.1152 P=1.64 MULT=1
MM1018 A_208_464# N_SCE_M1018_g N_VPWR_M1017_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.0864 PD=0.88 PS=0.91 NRD=19.9955 NRS=0 M=1 R=3.55556 SA=90000.6
+ SB=90001.7 A=0.1152 P=1.64 MULT=1
MM1028 N_A_292_464#_M1028_d N_D_M1028_g A_208_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.144 AS=0.0768 PD=1.09 PS=0.88 NRD=26.1616 NRS=19.9955 M=1 R=3.55556
+ SA=90001.1 SB=90001.3 A=0.1152 P=1.64 MULT=1
MM1013 A_418_464# N_A_27_464#_M1013_g N_A_292_464#_M1028_d VPB PSHORT L=0.18
+ W=0.64 AD=0.0768 AS=0.144 PD=0.88 PS=1.09 NRD=19.9955 NRS=26.1616 M=1
+ R=3.55556 SA=90001.7 SB=90000.7 A=0.1152 P=1.64 MULT=1
MM1019 N_VPWR_M1019_d N_SCD_M1019_g A_418_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.2858 AS=0.0768 PD=2.37 PS=0.88 NRD=26.1616 NRS=19.9955 M=1 R=3.55556
+ SA=90002.1 SB=90000.3 A=0.1152 P=1.64 MULT=1
MM1029 N_VPWR_M1029_d N_CLK_M1029_g N_A_599_74#_M1029_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1033 N_A_800_74#_M1033_d N_A_599_74#_M1033_g N_VPWR_M1029_d VPB PSHORT L=0.18
+ W=1.12 AD=0.2908 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1002 N_A_998_81#_M1002_d N_A_800_74#_M1002_g N_A_292_464#_M1002_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0672 AS=0.1176 PD=0.74 PS=1.4 NRD=21.0987 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90003.1 A=0.0756 P=1.2 MULT=1
MM1010 A_1131_457# N_A_599_74#_M1010_g N_A_998_81#_M1002_d VPB PSHORT L=0.18
+ W=0.42 AD=0.07035 AS=0.0672 PD=0.755 PS=0.74 NRD=52.7566 NRS=0 M=1 R=2.33333
+ SA=90000.7 SB=90002.6 A=0.0756 P=1.2 MULT=1
MM1020 N_VPWR_M1020_d N_A_1198_55#_M1020_g A_1131_457# VPB PSHORT L=0.18 W=0.42
+ AD=0.1586 AS=0.07035 PD=1.265 PS=0.755 NRD=151.316 NRS=52.7566 M=1 R=2.33333
+ SA=90001.2 SB=90002.1 A=0.0756 P=1.2 MULT=1
MM1030 N_A_1198_55#_M1030_d N_A_998_81#_M1030_g N_VPWR_M1020_d VPB PSHORT L=0.18
+ W=0.42 AD=0.063 AS=0.1586 PD=0.72 PS=1.265 NRD=11.7215 NRS=151.316 M=1
+ R=2.33333 SA=90001.9 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1024 N_VPWR_M1024_d N_SET_B_M1024_g N_A_1198_55#_M1030_d VPB PSHORT L=0.18
+ W=0.42 AD=0.105 AS=0.063 PD=0.887324 PS=0.72 NRD=105.533 NRS=0 M=1 R=2.33333
+ SA=90002.4 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1007 N_A_1613_341#_M1007_d N_A_998_81#_M1007_g N_VPWR_M1024_d VPB PSHORT
+ L=0.18 W=1 AD=0.27 AS=0.25 PD=2.54 PS=2.11268 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90001.4 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1038 N_A_1764_74#_M1038_d N_A_800_74#_M1038_g N_A_1721_374#_M1038_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.090093 AS=0.2521 PD=0.816338 PS=3.04 NRD=46.886 NRS=255.726
+ M=1 R=2.33333 SA=90000.2 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1016 N_A_1613_341#_M1016_d N_A_599_74#_M1016_g N_A_1764_74#_M1038_d VPB PSHORT
+ L=0.18 W=1 AD=0.265 AS=0.214507 PD=2.53 PS=1.94366 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.4 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1026 N_VPWR_M1026_d N_A_1958_48#_M1026_g N_A_1721_374#_M1026_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0567 AS=0.1134 PD=0.69 PS=1.38 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1031 N_A_1764_74#_M1031_d N_SET_B_M1031_g N_VPWR_M1026_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1134 AS=0.0567 PD=1.38 PS=0.69 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1035 N_VPWR_M1035_d N_A_1764_74#_M1035_g N_A_1958_48#_M1035_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.1134 AS=0.1134 PD=1.38 PS=1.38 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1027 N_VPWR_M1027_d N_A_1764_74#_M1027_g N_A_2395_112#_M1027_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.147 AS=0.2268 PD=1.23857 PS=2.22 NRD=10.5395 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1021 N_Q_M1021_d N_A_2395_112#_M1021_g N_VPWR_M1027_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3024 AS=0.196 PD=2.78 PS=1.65143 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX40_noxref VNB VPB NWDIODE A=26.7411 P=32.59
*
.include "sky130_fd_sc_ms__sdfstp_1.pxi.spice"
*
.ends
*
*

* NGSPICE file created from sky130_fd_sc_ms__o211a_4.ext - technology: sky130A

.subckt sky130_fd_sc_ms__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 VPWR C1 a_91_48# VPB pshort w=840000u l=180000u
+  ad=2.3588e+12p pd=1.71e+07u as=7.736e+11p ps=7.08e+06u
M1001 a_971_391# A2 a_91_48# VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=0p ps=0u
M1002 VGND a_91_48# X VNB nlowvt w=740000u l=150000u
+  ad=1.1032e+12p pd=1.016e+07u as=4.144e+11p ps=4.08e+06u
M1003 a_91_48# A2 a_971_391# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_91_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1005 VPWR A1 a_971_391# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_91_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_91_48# C1 VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_91_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_91_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR B1 a_91_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_510_125# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=8.089e+11p pd=7.65e+06u as=0p ps=0u
M1012 VGND A1 a_510_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_91_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_510_125# B1 a_597_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.032e+11p ps=3.82e+06u
M1015 a_597_125# C1 a_91_48# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1016 X a_91_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_91_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_971_391# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_597_125# B1 a_510_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_91_48# C1 a_597_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND A2 a_510_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_510_125# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_91_48# B1 VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


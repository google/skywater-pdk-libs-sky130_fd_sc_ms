* File: sky130_fd_sc_ms__nand3b_1.pxi.spice
* Created: Wed Sep  2 12:13:50 2020
* 
x_PM_SKY130_FD_SC_MS__NAND3B_1%A_N N_A_N_M1004_g N_A_N_M1005_g A_N N_A_N_c_52_n
+ N_A_N_c_53_n PM_SKY130_FD_SC_MS__NAND3B_1%A_N
x_PM_SKY130_FD_SC_MS__NAND3B_1%C N_C_M1001_g N_C_M1006_g C N_C_c_83_n N_C_c_84_n
+ PM_SKY130_FD_SC_MS__NAND3B_1%C
x_PM_SKY130_FD_SC_MS__NAND3B_1%B N_B_M1007_g N_B_M1003_g B N_B_c_119_n
+ N_B_c_120_n PM_SKY130_FD_SC_MS__NAND3B_1%B
x_PM_SKY130_FD_SC_MS__NAND3B_1%A_27_116# N_A_27_116#_M1004_s N_A_27_116#_M1005_s
+ N_A_27_116#_M1002_g N_A_27_116#_M1000_g N_A_27_116#_c_161_n
+ N_A_27_116#_c_162_n N_A_27_116#_c_163_n N_A_27_116#_c_164_n
+ N_A_27_116#_c_169_n N_A_27_116#_c_165_n N_A_27_116#_c_166_n
+ N_A_27_116#_c_167_n PM_SKY130_FD_SC_MS__NAND3B_1%A_27_116#
x_PM_SKY130_FD_SC_MS__NAND3B_1%VPWR N_VPWR_M1005_d N_VPWR_M1003_d N_VPWR_c_229_n
+ N_VPWR_c_230_n N_VPWR_c_231_n N_VPWR_c_232_n N_VPWR_c_233_n N_VPWR_c_234_n
+ VPWR N_VPWR_c_235_n N_VPWR_c_228_n PM_SKY130_FD_SC_MS__NAND3B_1%VPWR
x_PM_SKY130_FD_SC_MS__NAND3B_1%Y N_Y_M1002_d N_Y_M1001_d N_Y_M1000_d N_Y_c_270_n
+ N_Y_c_266_n N_Y_c_276_n N_Y_c_264_n Y Y Y N_Y_c_268_n N_Y_c_265_n
+ PM_SKY130_FD_SC_MS__NAND3B_1%Y
x_PM_SKY130_FD_SC_MS__NAND3B_1%VGND N_VGND_M1004_d N_VGND_c_308_n VGND
+ N_VGND_c_309_n N_VGND_c_310_n N_VGND_c_311_n N_VGND_c_312_n
+ PM_SKY130_FD_SC_MS__NAND3B_1%VGND
cc_1 VNB N_A_N_M1004_g 0.0310639f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.855
cc_2 VNB N_A_N_c_52_n 0.0285727f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.515
cc_3 VNB N_A_N_c_53_n 0.00453475f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.515
cc_4 VNB N_C_M1006_g 0.0255815f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.26
cc_5 VNB N_C_c_83_n 0.0270197f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.515
cc_6 VNB N_C_c_84_n 0.00176544f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.515
cc_7 VNB N_B_M1007_g 0.0233178f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.855
cc_8 VNB N_B_c_119_n 0.0247038f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.515
cc_9 VNB N_B_c_120_n 0.00404949f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.515
cc_10 VNB N_A_27_116#_M1002_g 0.0267595f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_11 VNB N_A_27_116#_M1000_g 5.51373e-19 $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.515
cc_12 VNB N_A_27_116#_c_161_n 0.0191713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_116#_c_162_n 0.0257611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_116#_c_163_n 0.00199818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_116#_c_164_n 0.0111529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_116#_c_165_n 0.0238989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_116#_c_166_n 0.00579502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_116#_c_167_n 0.0337966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_228_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_264_n 0.03984f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.515
cc_21 VNB N_Y_c_265_n 0.0239082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_308_n 0.0174336f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.26
cc_23 VNB N_VGND_c_309_n 0.0181018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_310_n 0.0508477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_311_n 0.21221f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.665
cc_26 VNB N_VGND_c_312_n 0.0129456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VPB N_A_N_M1005_g 0.0275135f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=2.26
cc_28 VPB N_A_N_c_52_n 0.00644565f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.515
cc_29 VPB N_A_N_c_53_n 0.0052982f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.515
cc_30 VPB N_C_M1001_g 0.0223871f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.855
cc_31 VPB N_C_c_83_n 0.00564388f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.515
cc_32 VPB N_C_c_84_n 0.0033292f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.515
cc_33 VPB N_B_M1003_g 0.0221693f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=2.26
cc_34 VPB N_B_c_119_n 0.00555109f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.515
cc_35 VPB N_B_c_120_n 0.00348571f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.515
cc_36 VPB N_A_27_116#_M1000_g 0.0301849f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.515
cc_37 VPB N_A_27_116#_c_169_n 0.0412197f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_A_27_116#_c_165_n 0.0140111f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_229_n 0.0195668f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_40 VPB N_VPWR_c_230_n 0.00899828f $X=-0.19 $Y=1.66 $X2=0.597 $Y2=1.68
cc_41 VPB N_VPWR_c_231_n 0.0255433f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_42 VPB N_VPWR_c_232_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_233_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_234_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_235_n 0.0220385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_228_n 0.0625687f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_Y_c_266_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.515
cc_48 VPB Y 0.0432986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_Y_c_268_n 0.0170713f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_Y_c_265_n 0.0078721f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 N_A_N_M1005_g N_C_M1001_g 0.0161897f $X=0.66 $Y=2.26 $X2=0 $Y2=0
cc_52 N_A_N_c_53_n N_C_M1001_g 2.8893e-19 $X=0.61 $Y=1.515 $X2=0 $Y2=0
cc_53 N_A_N_M1004_g N_C_M1006_g 0.00972195f $X=0.495 $Y=0.855 $X2=0 $Y2=0
cc_54 N_A_N_c_52_n N_C_c_83_n 0.0174241f $X=0.61 $Y=1.515 $X2=0 $Y2=0
cc_55 N_A_N_c_53_n N_C_c_83_n 0.00203135f $X=0.61 $Y=1.515 $X2=0 $Y2=0
cc_56 N_A_N_M1005_g N_C_c_84_n 3.17807e-19 $X=0.66 $Y=2.26 $X2=0 $Y2=0
cc_57 N_A_N_c_52_n N_C_c_84_n 3.73308e-19 $X=0.61 $Y=1.515 $X2=0 $Y2=0
cc_58 N_A_N_c_53_n N_C_c_84_n 0.0334549f $X=0.61 $Y=1.515 $X2=0 $Y2=0
cc_59 N_A_N_M1004_g N_A_27_116#_c_161_n 0.00199671f $X=0.495 $Y=0.855 $X2=0
+ $Y2=0
cc_60 N_A_N_M1004_g N_A_27_116#_c_162_n 0.0161994f $X=0.495 $Y=0.855 $X2=0 $Y2=0
cc_61 N_A_N_c_52_n N_A_27_116#_c_162_n 0.00138029f $X=0.61 $Y=1.515 $X2=0 $Y2=0
cc_62 N_A_N_c_53_n N_A_27_116#_c_162_n 0.0262311f $X=0.61 $Y=1.515 $X2=0 $Y2=0
cc_63 N_A_N_M1005_g N_A_27_116#_c_169_n 0.011136f $X=0.66 $Y=2.26 $X2=0 $Y2=0
cc_64 N_A_N_c_52_n N_A_27_116#_c_169_n 0.0017419f $X=0.61 $Y=1.515 $X2=0 $Y2=0
cc_65 N_A_N_c_53_n N_A_27_116#_c_169_n 0.0107727f $X=0.61 $Y=1.515 $X2=0 $Y2=0
cc_66 N_A_N_M1004_g N_A_27_116#_c_165_n 0.0129934f $X=0.495 $Y=0.855 $X2=0 $Y2=0
cc_67 N_A_N_M1005_g N_A_27_116#_c_165_n 0.00418724f $X=0.66 $Y=2.26 $X2=0 $Y2=0
cc_68 N_A_N_c_53_n N_A_27_116#_c_165_n 0.0331559f $X=0.61 $Y=1.515 $X2=0 $Y2=0
cc_69 N_A_N_M1005_g N_VPWR_c_229_n 0.00776968f $X=0.66 $Y=2.26 $X2=0 $Y2=0
cc_70 N_A_N_c_53_n N_VPWR_c_229_n 0.0024416f $X=0.61 $Y=1.515 $X2=0 $Y2=0
cc_71 N_A_N_M1005_g N_VPWR_c_231_n 0.00465228f $X=0.66 $Y=2.26 $X2=0 $Y2=0
cc_72 N_A_N_M1005_g N_VPWR_c_228_n 0.00555093f $X=0.66 $Y=2.26 $X2=0 $Y2=0
cc_73 N_A_N_M1004_g N_VGND_c_308_n 0.0112592f $X=0.495 $Y=0.855 $X2=0 $Y2=0
cc_74 N_A_N_M1004_g N_VGND_c_309_n 0.00365567f $X=0.495 $Y=0.855 $X2=0 $Y2=0
cc_75 N_A_N_M1004_g N_VGND_c_311_n 0.00404919f $X=0.495 $Y=0.855 $X2=0 $Y2=0
cc_76 N_C_M1006_g N_B_M1007_g 0.0388863f $X=1.27 $Y=0.76 $X2=0 $Y2=0
cc_77 N_C_M1001_g N_B_M1003_g 0.0181457f $X=1.245 $Y=2.4 $X2=0 $Y2=0
cc_78 N_C_c_84_n N_B_M1003_g 3.38586e-19 $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_79 N_C_c_83_n N_B_c_119_n 0.0388863f $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_80 N_C_c_84_n N_B_c_119_n 4.06701e-19 $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_81 N_C_M1001_g N_B_c_120_n 3.65824e-19 $X=1.245 $Y=2.4 $X2=0 $Y2=0
cc_82 N_C_c_83_n N_B_c_120_n 0.00202352f $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_83 N_C_c_84_n N_B_c_120_n 0.0286239f $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_84 N_C_M1006_g N_A_27_116#_c_162_n 0.0155047f $X=1.27 $Y=0.76 $X2=0 $Y2=0
cc_85 N_C_c_83_n N_A_27_116#_c_162_n 0.00121525f $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_86 N_C_c_84_n N_A_27_116#_c_162_n 0.021788f $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_87 N_C_M1001_g N_VPWR_c_229_n 0.00414244f $X=1.245 $Y=2.4 $X2=0 $Y2=0
cc_88 N_C_c_83_n N_VPWR_c_229_n 6.35946e-19 $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_89 N_C_c_84_n N_VPWR_c_229_n 0.00885662f $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_90 N_C_M1001_g N_VPWR_c_233_n 0.005209f $X=1.245 $Y=2.4 $X2=0 $Y2=0
cc_91 N_C_M1001_g N_VPWR_c_228_n 0.00986837f $X=1.245 $Y=2.4 $X2=0 $Y2=0
cc_92 N_C_M1001_g N_Y_c_270_n 0.00236361f $X=1.245 $Y=2.4 $X2=0 $Y2=0
cc_93 N_C_c_84_n N_Y_c_270_n 0.00280522f $X=1.18 $Y=1.515 $X2=0 $Y2=0
cc_94 N_C_M1001_g N_Y_c_266_n 0.0103488f $X=1.245 $Y=2.4 $X2=0 $Y2=0
cc_95 N_C_M1006_g N_VGND_c_308_n 0.01739f $X=1.27 $Y=0.76 $X2=0 $Y2=0
cc_96 N_C_M1006_g N_VGND_c_310_n 0.00468165f $X=1.27 $Y=0.76 $X2=0 $Y2=0
cc_97 N_C_M1006_g N_VGND_c_311_n 0.00453141f $X=1.27 $Y=0.76 $X2=0 $Y2=0
cc_98 N_B_M1007_g N_A_27_116#_M1002_g 0.0344152f $X=1.66 $Y=0.76 $X2=0 $Y2=0
cc_99 N_B_M1003_g N_A_27_116#_M1000_g 0.0217308f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_100 N_B_c_119_n N_A_27_116#_M1000_g 0.00167197f $X=1.75 $Y=1.515 $X2=0 $Y2=0
cc_101 N_B_c_120_n N_A_27_116#_M1000_g 0.0024834f $X=1.75 $Y=1.515 $X2=0 $Y2=0
cc_102 N_B_M1007_g N_A_27_116#_c_162_n 0.0154731f $X=1.66 $Y=0.76 $X2=0 $Y2=0
cc_103 N_B_c_119_n N_A_27_116#_c_162_n 0.00121439f $X=1.75 $Y=1.515 $X2=0 $Y2=0
cc_104 N_B_c_120_n N_A_27_116#_c_162_n 0.0232305f $X=1.75 $Y=1.515 $X2=0 $Y2=0
cc_105 N_B_M1007_g N_A_27_116#_c_163_n 0.00296442f $X=1.66 $Y=0.76 $X2=0 $Y2=0
cc_106 N_B_M1007_g N_A_27_116#_c_166_n 5.87559e-19 $X=1.66 $Y=0.76 $X2=0 $Y2=0
cc_107 N_B_c_119_n N_A_27_116#_c_166_n 0.00170526f $X=1.75 $Y=1.515 $X2=0 $Y2=0
cc_108 N_B_c_120_n N_A_27_116#_c_166_n 0.0240984f $X=1.75 $Y=1.515 $X2=0 $Y2=0
cc_109 N_B_c_119_n N_A_27_116#_c_167_n 0.018763f $X=1.75 $Y=1.515 $X2=0 $Y2=0
cc_110 N_B_c_120_n N_A_27_116#_c_167_n 3.43837e-19 $X=1.75 $Y=1.515 $X2=0 $Y2=0
cc_111 N_B_M1003_g N_VPWR_c_230_n 0.00203999f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_112 N_B_M1003_g N_VPWR_c_233_n 0.005209f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_113 N_B_M1003_g N_VPWR_c_228_n 0.00982687f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_114 N_B_M1003_g N_Y_c_270_n 8.8334e-19 $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_115 N_B_c_120_n N_Y_c_270_n 0.0041171f $X=1.75 $Y=1.515 $X2=0 $Y2=0
cc_116 N_B_M1003_g N_Y_c_266_n 0.0119155f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_117 N_B_M1003_g N_Y_c_276_n 0.0134232f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_118 N_B_c_119_n N_Y_c_276_n 5.99772e-19 $X=1.75 $Y=1.515 $X2=0 $Y2=0
cc_119 N_B_c_120_n N_Y_c_276_n 0.0192103f $X=1.75 $Y=1.515 $X2=0 $Y2=0
cc_120 N_B_M1007_g N_Y_c_264_n 0.00193784f $X=1.66 $Y=0.76 $X2=0 $Y2=0
cc_121 N_B_M1003_g N_Y_c_268_n 0.00127282f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_122 N_B_M1007_g N_VGND_c_308_n 0.00269744f $X=1.66 $Y=0.76 $X2=0 $Y2=0
cc_123 N_B_M1007_g N_VGND_c_310_n 0.00563421f $X=1.66 $Y=0.76 $X2=0 $Y2=0
cc_124 N_B_M1007_g N_VGND_c_311_n 0.00539454f $X=1.66 $Y=0.76 $X2=0 $Y2=0
cc_125 N_A_27_116#_c_169_n N_VPWR_c_229_n 0.0264352f $X=0.435 $Y=2.115 $X2=0
+ $Y2=0
cc_126 N_A_27_116#_M1000_g N_VPWR_c_230_n 0.00343717f $X=2.245 $Y=2.4 $X2=0
+ $Y2=0
cc_127 N_A_27_116#_c_169_n N_VPWR_c_231_n 0.0100209f $X=0.435 $Y=2.115 $X2=0
+ $Y2=0
cc_128 N_A_27_116#_M1000_g N_VPWR_c_235_n 0.005209f $X=2.245 $Y=2.4 $X2=0 $Y2=0
cc_129 N_A_27_116#_M1000_g N_VPWR_c_228_n 0.00986692f $X=2.245 $Y=2.4 $X2=0
+ $Y2=0
cc_130 N_A_27_116#_c_169_n N_VPWR_c_228_n 0.0149809f $X=0.435 $Y=2.115 $X2=0
+ $Y2=0
cc_131 N_A_27_116#_M1000_g N_Y_c_266_n 6.00071e-19 $X=2.245 $Y=2.4 $X2=0 $Y2=0
cc_132 N_A_27_116#_M1000_g N_Y_c_276_n 0.014772f $X=2.245 $Y=2.4 $X2=0 $Y2=0
cc_133 N_A_27_116#_c_166_n N_Y_c_276_n 0.00895052f $X=2.29 $Y=1.485 $X2=0 $Y2=0
cc_134 N_A_27_116#_M1002_g N_Y_c_264_n 0.0222284f $X=2.2 $Y=0.76 $X2=0 $Y2=0
cc_135 N_A_27_116#_c_162_n N_Y_c_264_n 0.0145858f $X=2.085 $Y=1.065 $X2=0 $Y2=0
cc_136 N_A_27_116#_c_166_n N_Y_c_264_n 0.00703632f $X=2.29 $Y=1.485 $X2=0 $Y2=0
cc_137 N_A_27_116#_c_167_n N_Y_c_264_n 0.00330893f $X=2.29 $Y=1.485 $X2=0 $Y2=0
cc_138 N_A_27_116#_M1000_g Y 0.0132321f $X=2.245 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A_27_116#_M1000_g N_Y_c_268_n 0.00461176f $X=2.245 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A_27_116#_c_166_n N_Y_c_268_n 0.0124349f $X=2.29 $Y=1.485 $X2=0 $Y2=0
cc_141 N_A_27_116#_c_167_n N_Y_c_268_n 0.00279548f $X=2.29 $Y=1.485 $X2=0 $Y2=0
cc_142 N_A_27_116#_M1002_g N_Y_c_265_n 0.00203887f $X=2.2 $Y=0.76 $X2=0 $Y2=0
cc_143 N_A_27_116#_M1000_g N_Y_c_265_n 0.00367386f $X=2.245 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A_27_116#_c_163_n N_Y_c_265_n 0.00479588f $X=2.17 $Y=1.32 $X2=0 $Y2=0
cc_145 N_A_27_116#_c_166_n N_Y_c_265_n 0.0249903f $X=2.29 $Y=1.485 $X2=0 $Y2=0
cc_146 N_A_27_116#_c_167_n N_Y_c_265_n 0.00231223f $X=2.29 $Y=1.485 $X2=0 $Y2=0
cc_147 N_A_27_116#_c_162_n N_VGND_M1004_d 0.00761754f $X=2.085 $Y=1.065
+ $X2=-0.19 $Y2=-0.245
cc_148 N_A_27_116#_c_161_n N_VGND_c_308_n 0.0112316f $X=0.28 $Y=0.855 $X2=0
+ $Y2=0
cc_149 N_A_27_116#_c_162_n N_VGND_c_308_n 0.0451464f $X=2.085 $Y=1.065 $X2=0
+ $Y2=0
cc_150 N_A_27_116#_c_161_n N_VGND_c_309_n 0.00637154f $X=0.28 $Y=0.855 $X2=0
+ $Y2=0
cc_151 N_A_27_116#_M1002_g N_VGND_c_310_n 0.0053639f $X=2.2 $Y=0.76 $X2=0 $Y2=0
cc_152 N_A_27_116#_M1002_g N_VGND_c_311_n 0.00539454f $X=2.2 $Y=0.76 $X2=0 $Y2=0
cc_153 N_A_27_116#_c_161_n N_VGND_c_311_n 0.00857079f $X=0.28 $Y=0.855 $X2=0
+ $Y2=0
cc_154 N_A_27_116#_c_162_n A_269_78# 0.0048076f $X=2.085 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_155 N_A_27_116#_c_162_n A_347_78# 0.0107783f $X=2.085 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_156 N_VPWR_c_229_n N_Y_c_266_n 0.0330222f $X=0.97 $Y=2.035 $X2=0 $Y2=0
cc_157 N_VPWR_c_230_n N_Y_c_266_n 0.0266809f $X=1.97 $Y=2.455 $X2=0 $Y2=0
cc_158 N_VPWR_c_233_n N_Y_c_266_n 0.0144623f $X=1.805 $Y=3.33 $X2=0 $Y2=0
cc_159 N_VPWR_c_228_n N_Y_c_266_n 0.0118344f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_160 N_VPWR_M1003_d N_Y_c_276_n 0.0101293f $X=1.785 $Y=1.84 $X2=0 $Y2=0
cc_161 N_VPWR_c_230_n N_Y_c_276_n 0.0208278f $X=1.97 $Y=2.455 $X2=0 $Y2=0
cc_162 N_VPWR_c_230_n Y 0.0282945f $X=1.97 $Y=2.455 $X2=0 $Y2=0
cc_163 N_VPWR_c_235_n Y 0.0216883f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_164 N_VPWR_c_228_n Y 0.0178836f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_165 N_Y_c_264_n N_VGND_c_310_n 0.0221969f $X=2.71 $Y=1.15 $X2=0 $Y2=0
cc_166 N_Y_c_264_n N_VGND_c_311_n 0.0197591f $X=2.71 $Y=1.15 $X2=0 $Y2=0

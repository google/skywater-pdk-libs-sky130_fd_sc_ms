* File: sky130_fd_sc_ms__nor3b_2.pex.spice
* Created: Fri Aug 28 17:48:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NOR3B_2%C_N 3 7 9 12
c34 12 0 1.05511e-19 $X=0.59 $Y=1.615
r35 12 15 40.7387 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.582 $Y=1.615
+ $X2=0.582 $Y2=1.78
r36 12 14 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.582 $Y=1.615
+ $X2=0.582 $Y2=1.45
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.615 $X2=0.59 $Y2=1.615
r38 9 13 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.72 $Y=1.615
+ $X2=0.59 $Y2=1.615
r39 7 14 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.5 $Y=0.69 $X2=0.5
+ $Y2=1.45
r40 3 15 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=0.5 $Y=2.46 $X2=0.5
+ $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3B_2%A_27_392# 1 2 7 9 12 14 16 19 23 27 29 33 35
+ 36 37 46
c79 37 0 1.05511e-19 $X=1.17 $Y=1.195
c80 19 0 1.87864e-19 $X=1.95 $Y=2.4
c81 14 0 1.49881e-19 $X=1.515 $Y=1.22
r82 45 46 2.25234 $w=3.21e-07 $l=1.5e-08 $layer=POLY_cond $X=1.5 $Y=1.385
+ $X2=1.515 $Y2=1.385
r83 41 45 49.5514 $w=3.21e-07 $l=3.3e-07 $layer=POLY_cond $X=1.17 $Y=1.385
+ $X2=1.5 $Y2=1.385
r84 41 43 15.0156 $w=3.21e-07 $l=1e-07 $layer=POLY_cond $X=1.17 $Y=1.385
+ $X2=1.07 $Y2=1.385
r85 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.385 $X2=1.17 $Y2=1.385
r86 37 40 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=1.17 $Y=1.195
+ $X2=1.17 $Y2=1.385
r87 34 35 3.01551 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.45 $Y=1.195
+ $X2=0.267 $Y2=1.195
r88 33 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=1.195
+ $X2=1.17 $Y2=1.195
r89 33 34 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.005 $Y=1.195
+ $X2=0.45 $Y2=1.195
r90 29 31 29.3349 $w=2.73e-07 $l=7e-07 $layer=LI1_cond $X=0.222 $Y=2.115
+ $X2=0.222 $Y2=2.815
r91 27 36 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=0.222 $Y=2.087
+ $X2=0.222 $Y2=1.95
r92 27 29 1.1734 $w=2.73e-07 $l=2.8e-08 $layer=LI1_cond $X=0.222 $Y=2.087
+ $X2=0.222 $Y2=2.115
r93 25 35 3.49088 $w=2.67e-07 $l=1.32868e-07 $layer=LI1_cond $X=0.17 $Y=1.28
+ $X2=0.267 $Y2=1.195
r94 25 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.17 $Y=1.28
+ $X2=0.17 $Y2=1.95
r95 21 35 3.49088 $w=2.67e-07 $l=8.5e-08 $layer=LI1_cond $X=0.267 $Y=1.11
+ $X2=0.267 $Y2=1.195
r96 21 23 18.7864 $w=3.63e-07 $l=5.95e-07 $layer=LI1_cond $X=0.267 $Y=1.11
+ $X2=0.267 $Y2=0.515
r97 17 46 65.3178 $w=3.21e-07 $l=4.35e-07 $layer=POLY_cond $X=1.95 $Y=1.385
+ $X2=1.515 $Y2=1.385
r98 17 19 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=1.95 $Y=1.53
+ $X2=1.95 $Y2=2.4
r99 14 46 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=1.22
+ $X2=1.515 $Y2=1.385
r100 14 16 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.515 $Y=1.22
+ $X2=1.515 $Y2=0.74
r101 10 45 16.2883 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.5 $Y=1.55
+ $X2=1.5 $Y2=1.385
r102 10 12 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.5 $Y=1.55 $X2=1.5
+ $Y2=2.4
r103 7 43 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.07 $Y=1.22
+ $X2=1.07 $Y2=1.385
r104 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.07 $Y=1.22 $X2=1.07
+ $Y2=0.74
r105 2 31 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.275 $Y2=2.815
r106 2 29 400 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.275 $Y2=2.115
r107 1 23 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.37 $X2=0.285 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3B_2%B 3 7 11 15 17 19 21
r52 30 31 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=2.815 $Y=1.515
+ $X2=2.85 $Y2=1.515
r53 28 30 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=2.77 $Y=1.515
+ $X2=2.815 $Y2=1.515
r54 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.515 $X2=2.77 $Y2=1.515
r55 26 28 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=2.4 $Y=1.515
+ $X2=2.77 $Y2=1.515
r56 24 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.385 $Y=1.515
+ $X2=2.4 $Y2=1.515
r57 22 29 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=3.11 $Y=1.565
+ $X2=2.77 $Y2=1.565
r58 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.11
+ $Y=1.515 $X2=3.11 $Y2=1.515
r59 19 31 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.94 $Y=1.515 $X2=2.85
+ $Y2=1.515
r60 19 21 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=2.94 $Y=1.515
+ $X2=3.11 $Y2=1.515
r61 17 22 0.26801 $w=4.28e-07 $l=1e-08 $layer=LI1_cond $X=3.12 $Y=1.565 $X2=3.11
+ $Y2=1.565
r62 13 31 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.85 $Y=1.68
+ $X2=2.85 $Y2=1.515
r63 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.85 $Y=1.68
+ $X2=2.85 $Y2=2.4
r64 9 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.815 $Y=1.35
+ $X2=2.815 $Y2=1.515
r65 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.815 $Y=1.35
+ $X2=2.815 $Y2=0.74
r66 5 26 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.4 $Y=1.68 $X2=2.4
+ $Y2=1.515
r67 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.4 $Y=1.68 $X2=2.4
+ $Y2=2.4
r68 1 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.385 $Y=1.35
+ $X2=2.385 $Y2=1.515
r69 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.385 $Y=1.35
+ $X2=2.385 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3B_2%A 3 7 11 15 17 18 19 30
c47 11 0 1.81748e-19 $X=4.285 $Y=0.74
r48 29 30 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.285 $Y=1.515
+ $X2=4.3 $Y2=1.515
r49 27 29 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.195 $Y=1.515
+ $X2=4.285 $Y2=1.515
r50 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.195
+ $Y=1.515 $X2=4.195 $Y2=1.515
r51 25 27 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=3.85 $Y=1.515
+ $X2=4.195 $Y2=1.515
r52 23 25 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=3.805 $Y=1.515
+ $X2=3.85 $Y2=1.515
r53 19 28 9.78236 $w=4.28e-07 $l=3.65e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.195 $Y2=1.565
r54 18 28 3.08211 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=4.195 $Y2=1.565
r55 17 18 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=4.08 $Y2=1.565
r56 13 30 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.3 $Y=1.68 $X2=4.3
+ $Y2=1.515
r57 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.3 $Y=1.68 $X2=4.3
+ $Y2=2.4
r58 9 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.285 $Y=1.35
+ $X2=4.285 $Y2=1.515
r59 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.285 $Y=1.35
+ $X2=4.285 $Y2=0.74
r60 5 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.85 $Y=1.68
+ $X2=3.85 $Y2=1.515
r61 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.85 $Y=1.68 $X2=3.85
+ $Y2=2.4
r62 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.805 $Y=1.35
+ $X2=3.805 $Y2=1.515
r63 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.805 $Y=1.35
+ $X2=3.805 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3B_2%VPWR 1 2 3 12 18 20 22 26 28 33 41 47 50 54
r56 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r57 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r58 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 45 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r60 45 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r61 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r62 42 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.79 $Y=3.33
+ $X2=3.625 $Y2=3.33
r63 42 44 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.79 $Y=3.33
+ $X2=4.08 $Y2=3.33
r64 41 53 4.14492 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.612 $Y2=3.33
r65 41 44 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.08 $Y2=3.33
r66 40 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r67 39 40 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r68 37 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r69 36 39 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r70 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r71 34 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=3.33
+ $X2=0.725 $Y2=3.33
r72 34 36 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.89 $Y=3.33 $X2=1.2
+ $Y2=3.33
r73 33 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.46 $Y=3.33
+ $X2=3.625 $Y2=3.33
r74 33 39 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.46 $Y=3.33
+ $X2=3.12 $Y2=3.33
r75 31 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r76 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r77 28 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.725 $Y2=3.33
r78 28 30 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33 $X2=0.24
+ $Y2=3.33
r79 26 40 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=3.12 $Y2=3.33
r80 26 37 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r81 22 25 30.4419 $w=2.63e-07 $l=7e-07 $layer=LI1_cond $X=4.557 $Y=2.115
+ $X2=4.557 $Y2=2.815
r82 20 53 3.10315 $w=2.65e-07 $l=1.09087e-07 $layer=LI1_cond $X=4.557 $Y=3.245
+ $X2=4.612 $Y2=3.33
r83 20 25 18.7 $w=2.63e-07 $l=4.3e-07 $layer=LI1_cond $X=4.557 $Y=3.245
+ $X2=4.557 $Y2=2.815
r84 16 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=3.245
+ $X2=3.625 $Y2=3.33
r85 16 18 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=3.625 $Y=3.245
+ $X2=3.625 $Y2=2.395
r86 12 15 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.725 $Y=2.115
+ $X2=0.725 $Y2=2.815
r87 10 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=3.33
r88 10 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=2.815
r89 3 25 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.39
+ $Y=1.84 $X2=4.525 $Y2=2.815
r90 3 22 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=4.39
+ $Y=1.84 $X2=4.525 $Y2=2.115
r91 2 18 300 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_PDIFF $count=2 $X=3.485
+ $Y=1.84 $X2=3.625 $Y2=2.395
r92 1 15 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.96 $X2=0.725 $Y2=2.815
r93 1 12 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.96 $X2=0.725 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3B_2%A_227_368# 1 2 3 12 16 17 20 24 28 30
r44 26 28 19.2074 $w=2.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.105 $Y=2.905
+ $X2=3.105 $Y2=2.455
r45 25 30 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.29 $Y=2.99 $X2=2.15
+ $Y2=2.99
r46 24 26 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.97 $Y=2.99
+ $X2=3.105 $Y2=2.905
r47 24 25 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.97 $Y=2.99
+ $X2=2.29 $Y2=2.99
r48 20 23 34.1617 $w=2.78e-07 $l=8.3e-07 $layer=LI1_cond $X=2.15 $Y=1.985
+ $X2=2.15 $Y2=2.815
r49 18 30 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=2.905
+ $X2=2.15 $Y2=2.99
r50 18 23 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=2.15 $Y=2.905 $X2=2.15
+ $Y2=2.815
r51 16 30 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.01 $Y=2.99 $X2=2.15
+ $Y2=2.99
r52 16 17 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.01 $Y=2.99
+ $X2=1.44 $Y2=2.99
r53 12 15 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.275 $Y=1.985
+ $X2=1.275 $Y2=2.815
r54 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.275 $Y=2.905
+ $X2=1.44 $Y2=2.99
r55 10 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.275 $Y=2.905
+ $X2=1.275 $Y2=2.815
r56 3 28 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=2.94
+ $Y=1.84 $X2=3.075 $Y2=2.455
r57 2 23 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.04
+ $Y=1.84 $X2=2.175 $Y2=2.815
r58 2 20 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.04
+ $Y=1.84 $X2=2.175 $Y2=1.985
r59 1 15 400 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=1 $X=1.135
+ $Y=1.84 $X2=1.275 $Y2=2.815
r60 1 12 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.135
+ $Y=1.84 $X2=1.275 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3B_2%Y 1 2 3 4 15 19 23 25 29 31 33 34 35 38
c59 25 0 1.81748e-19 $X=3.925 $Y=1.045
c60 15 0 1.49881e-19 $X=1.285 $Y=0.515
r61 38 45 4.30525 $w=3.6e-07 $l=8.9861e-08 $layer=LI1_cond $X=1.81 $Y=0.95
+ $X2=1.725 $Y2=0.94
r62 35 38 11.2043 $w=3.58e-07 $l=3.5e-07 $layer=LI1_cond $X=2.16 $Y=0.95
+ $X2=1.81 $Y2=0.95
r63 34 45 2.31646 $w=2.37e-07 $l=4.5e-08 $layer=LI1_cond $X=1.68 $Y=0.94
+ $X2=1.725 $Y2=0.94
r64 31 35 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=2.505 $Y=0.95
+ $X2=2.16 $Y2=0.95
r65 31 33 3.88469 $w=2.65e-07 $l=9.5e-08 $layer=LI1_cond $X=2.505 $Y=0.95
+ $X2=2.6 $Y2=0.95
r66 27 29 19.7245 $w=2.58e-07 $l=4.45e-07 $layer=LI1_cond $X=4.055 $Y=0.96
+ $X2=4.055 $Y2=0.515
r67 26 33 3.88469 $w=2.65e-07 $l=1.3435e-07 $layer=LI1_cond $X=2.695 $Y=1.045
+ $X2=2.6 $Y2=0.95
r68 25 27 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.925 $Y=1.045
+ $X2=4.055 $Y2=0.96
r69 25 26 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=3.925 $Y=1.045
+ $X2=2.695 $Y2=1.045
r70 21 33 2.5638 $w=1.9e-07 $l=1.8e-07 $layer=LI1_cond $X=2.6 $Y=0.77 $X2=2.6
+ $Y2=0.95
r71 21 23 14.8852 $w=1.88e-07 $l=2.55e-07 $layer=LI1_cond $X=2.6 $Y=0.77 $X2=2.6
+ $Y2=0.515
r72 17 45 2.684 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.725 $Y=1.13 $X2=1.725
+ $Y2=0.94
r73 17 19 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=1.725 $Y=1.13
+ $X2=1.725 $Y2=1.985
r74 13 34 21.7747 $w=2.37e-07 $l=4.23e-07 $layer=LI1_cond $X=1.257 $Y=0.94
+ $X2=1.68 $Y2=0.94
r75 13 15 10.6863 $w=2.73e-07 $l=2.55e-07 $layer=LI1_cond $X=1.257 $Y=0.77
+ $X2=1.257 $Y2=0.515
r76 4 19 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.59
+ $Y=1.84 $X2=1.725 $Y2=1.985
r77 3 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.88
+ $Y=0.37 $X2=4.02 $Y2=0.515
r78 2 33 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=2.46
+ $Y=0.37 $X2=2.6 $Y2=0.965
r79 2 23 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.46
+ $Y=0.37 $X2=2.6 $Y2=0.515
r80 1 13 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=1.145
+ $Y=0.37 $X2=1.285 $Y2=0.855
r81 1 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.145
+ $Y=0.37 $X2=1.285 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3B_2%A_498_368# 1 2 9 11 13 16
c27 16 0 1.87864e-19 $X=2.625 $Y=2.035
r28 11 18 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.115 $Y=2.12
+ $X2=4.115 $Y2=2.035
r29 11 13 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=4.115 $Y=2.12
+ $X2=4.115 $Y2=2.44
r30 10 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.79 $Y=2.035
+ $X2=2.625 $Y2=2.035
r31 9 18 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.99 $Y=2.035
+ $X2=4.115 $Y2=2.035
r32 9 10 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=3.99 $Y=2.035
+ $X2=2.79 $Y2=2.035
r33 2 18 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=3.94
+ $Y=1.84 $X2=4.075 $Y2=2.035
r34 2 13 300 $w=1.7e-07 $l=6.64078e-07 $layer=licon1_PDIFF $count=2 $X=3.94
+ $Y=1.84 $X2=4.075 $Y2=2.44
r35 1 16 300 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=2 $X=2.49
+ $Y=1.84 $X2=2.625 $Y2=2.035
.ends

.subckt PM_SKY130_FD_SC_MS__NOR3B_2%VGND 1 2 3 4 15 17 19 21 23 38 44 49 55 58
+ 62 65
r65 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r66 60 62 11.8599 $w=8.53e-07 $l=1.55e-07 $layer=LI1_cond $X=3.6 $Y=0.342
+ $X2=3.755 $Y2=0.342
r67 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r68 57 60 0.14269 $w=8.53e-07 $l=1e-08 $layer=LI1_cond $X=3.59 $Y=0.342 $X2=3.6
+ $Y2=0.342
r69 57 58 19.9932 $w=8.53e-07 $l=7.25e-07 $layer=LI1_cond $X=3.59 $Y=0.342
+ $X2=2.865 $Y2=0.342
r70 54 55 10.7086 $w=6.83e-07 $l=1.65e-07 $layer=LI1_cond $X=2.17 $Y=0.257
+ $X2=2.335 $Y2=0.257
r71 51 54 0.17461 $w=6.83e-07 $l=1e-08 $layer=LI1_cond $X=2.16 $Y=0.257 $X2=2.17
+ $Y2=0.257
r72 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r73 48 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r74 47 51 8.38128 $w=6.83e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=0.257
+ $X2=2.16 $Y2=0.257
r75 47 49 9.83558 $w=6.83e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=0.257
+ $X2=1.565 $Y2=0.257
r76 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r77 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r78 42 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r79 42 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r80 41 62 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=3.755
+ $Y2=0
r81 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r82 38 64 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.577
+ $Y2=0
r83 38 41 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.08
+ $Y2=0
r84 37 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r85 36 58 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=2.865
+ $Y2=0
r86 36 55 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=2.335
+ $Y2=0
r87 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r88 32 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r89 32 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r90 31 49 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.565
+ $Y2=0
r91 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r92 29 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.785
+ $Y2=0
r93 29 31 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.2
+ $Y2=0
r94 26 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r95 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r96 23 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.785
+ $Y2=0
r97 23 25 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.24
+ $Y2=0
r98 21 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r99 21 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r100 17 64 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.52 $Y=0.085
+ $X2=4.577 $Y2=0
r101 17 19 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.52 $Y=0.085
+ $X2=4.52 $Y2=0.515
r102 13 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0
r103 13 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0.515
r104 4 19 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=4.36
+ $Y=0.37 $X2=4.52 $Y2=0.515
r105 3 57 91 $w=1.7e-07 $l=8.09012e-07 $layer=licon1_NDIFF $count=2 $X=2.89
+ $Y=0.37 $X2=3.59 $Y2=0.605
r106 2 54 91 $w=1.7e-07 $l=6.4846e-07 $layer=licon1_NDIFF $count=2 $X=1.59
+ $Y=0.37 $X2=2.17 $Y2=0.515
r107 1 15 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=0.575
+ $Y=0.37 $X2=0.785 $Y2=0.515
.ends


* File: sky130_fd_sc_ms__sdfstp_2.pxi.spice
* Created: Wed Sep  2 12:31:14 2020
* 
x_PM_SKY130_FD_SC_MS__SDFSTP_2%SCE N_SCE_c_320_n N_SCE_M1015_g N_SCE_M1043_g
+ N_SCE_c_322_n N_SCE_M1016_g N_SCE_M1039_g N_SCE_c_315_n N_SCE_c_316_n
+ N_SCE_c_317_n N_SCE_c_318_n SCE N_SCE_c_319_n PM_SKY130_FD_SC_MS__SDFSTP_2%SCE
x_PM_SKY130_FD_SC_MS__SDFSTP_2%A_27_74# N_A_27_74#_M1043_s N_A_27_74#_M1015_s
+ N_A_27_74#_M1038_g N_A_27_74#_M1005_g N_A_27_74#_c_391_n N_A_27_74#_c_392_n
+ N_A_27_74#_c_407_n N_A_27_74#_c_393_n N_A_27_74#_c_394_n N_A_27_74#_c_399_n
+ N_A_27_74#_c_400_n N_A_27_74#_c_395_n N_A_27_74#_c_401_n N_A_27_74#_c_396_n
+ PM_SKY130_FD_SC_MS__SDFSTP_2%A_27_74#
x_PM_SKY130_FD_SC_MS__SDFSTP_2%D N_D_M1023_g N_D_M1028_g D N_D_c_473_n
+ N_D_c_474_n PM_SKY130_FD_SC_MS__SDFSTP_2%D
x_PM_SKY130_FD_SC_MS__SDFSTP_2%SCD N_SCD_M1035_g N_SCD_c_515_n N_SCD_M1017_g SCD
+ SCD SCD N_SCD_c_517_n N_SCD_c_521_n PM_SKY130_FD_SC_MS__SDFSTP_2%SCD
x_PM_SKY130_FD_SC_MS__SDFSTP_2%CLK N_CLK_M1012_g N_CLK_M1032_g CLK N_CLK_c_560_n
+ N_CLK_c_561_n PM_SKY130_FD_SC_MS__SDFSTP_2%CLK
x_PM_SKY130_FD_SC_MS__SDFSTP_2%A_795_74# N_A_795_74#_M1006_d N_A_795_74#_M1040_d
+ N_A_795_74#_M1034_g N_A_795_74#_c_596_n N_A_795_74#_c_597_n
+ N_A_795_74#_M1031_g N_A_795_74#_c_599_n N_A_795_74#_c_600_n
+ N_A_795_74#_c_601_n N_A_795_74#_M1001_g N_A_795_74#_c_602_n
+ N_A_795_74#_c_603_n N_A_795_74#_M1036_g N_A_795_74#_M1019_g
+ N_A_795_74#_c_604_n N_A_795_74#_c_605_n N_A_795_74#_c_621_n
+ N_A_795_74#_c_606_n N_A_795_74#_c_607_n N_A_795_74#_c_622_n
+ N_A_795_74#_c_623_n N_A_795_74#_c_608_n N_A_795_74#_c_609_n
+ N_A_795_74#_c_625_n N_A_795_74#_c_626_n N_A_795_74#_c_627_n
+ N_A_795_74#_c_628_n N_A_795_74#_c_629_n N_A_795_74#_c_630_n
+ N_A_795_74#_c_631_n N_A_795_74#_c_632_n N_A_795_74#_c_610_n
+ N_A_795_74#_c_611_n N_A_795_74#_c_635_n N_A_795_74#_c_636_n
+ N_A_795_74#_c_612_n N_A_795_74#_c_637_n N_A_795_74#_c_613_n
+ N_A_795_74#_c_614_n N_A_795_74#_c_615_n N_A_795_74#_c_616_n
+ N_A_795_74#_c_617_n PM_SKY130_FD_SC_MS__SDFSTP_2%A_795_74#
x_PM_SKY130_FD_SC_MS__SDFSTP_2%A_1185_55# N_A_1185_55#_M1026_s
+ N_A_1185_55#_M1011_d N_A_1185_55#_c_874_n N_A_1185_55#_M1020_g
+ N_A_1185_55#_M1042_g N_A_1185_55#_c_875_n N_A_1185_55#_c_876_n
+ N_A_1185_55#_c_882_n N_A_1185_55#_c_877_n N_A_1185_55#_c_896_n
+ N_A_1185_55#_c_883_n N_A_1185_55#_c_878_n N_A_1185_55#_c_885_n
+ N_A_1185_55#_c_879_n N_A_1185_55#_c_880_n
+ PM_SKY130_FD_SC_MS__SDFSTP_2%A_1185_55#
x_PM_SKY130_FD_SC_MS__SDFSTP_2%A_991_81# N_A_991_81#_M1024_d N_A_991_81#_M1034_d
+ N_A_991_81#_c_970_n N_A_991_81#_M1011_g N_A_991_81#_c_972_n
+ N_A_991_81#_M1026_g N_A_991_81#_M1000_g N_A_991_81#_c_974_n
+ N_A_991_81#_M1029_g N_A_991_81#_M1007_g N_A_991_81#_c_976_n
+ N_A_991_81#_M1033_g N_A_991_81#_c_977_n N_A_991_81#_c_991_n
+ N_A_991_81#_c_992_n N_A_991_81#_c_978_n N_A_991_81#_c_979_n
+ N_A_991_81#_c_980_n N_A_991_81#_c_1064_n N_A_991_81#_c_981_n
+ N_A_991_81#_c_982_n N_A_991_81#_c_983_n N_A_991_81#_c_984_n
+ N_A_991_81#_c_985_n N_A_991_81#_c_986_n N_A_991_81#_c_987_n
+ PM_SKY130_FD_SC_MS__SDFSTP_2%A_991_81#
x_PM_SKY130_FD_SC_MS__SDFSTP_2%SET_B N_SET_B_M1021_g N_SET_B_M1027_g
+ N_SET_B_M1013_g N_SET_B_M1025_g N_SET_B_c_1155_n N_SET_B_c_1156_n
+ N_SET_B_c_1157_n SET_B N_SET_B_c_1159_n N_SET_B_c_1160_n N_SET_B_c_1161_n
+ PM_SKY130_FD_SC_MS__SDFSTP_2%SET_B
x_PM_SKY130_FD_SC_MS__SDFSTP_2%A_608_74# N_A_608_74#_M1012_s N_A_608_74#_M1032_s
+ N_A_608_74#_M1006_g N_A_608_74#_M1040_g N_A_608_74#_c_1285_n
+ N_A_608_74#_c_1299_n N_A_608_74#_c_1286_n N_A_608_74#_c_1287_n
+ N_A_608_74#_c_1300_n N_A_608_74#_c_1301_n N_A_608_74#_M1024_g
+ N_A_608_74#_M1018_g N_A_608_74#_c_1303_n N_A_608_74#_M1003_g
+ N_A_608_74#_c_1290_n N_A_608_74#_c_1291_n N_A_608_74#_c_1305_n
+ N_A_608_74#_c_1306_n N_A_608_74#_M1010_g N_A_608_74#_M1044_g
+ N_A_608_74#_c_1307_n N_A_608_74#_c_1308_n N_A_608_74#_c_1309_n
+ N_A_608_74#_c_1310_n N_A_608_74#_c_1293_n N_A_608_74#_c_1294_n
+ N_A_608_74#_c_1312_n N_A_608_74#_c_1313_n N_A_608_74#_c_1295_n
+ N_A_608_74#_c_1296_n N_A_608_74#_c_1297_n
+ PM_SKY130_FD_SC_MS__SDFSTP_2%A_608_74#
x_PM_SKY130_FD_SC_MS__SDFSTP_2%A_2186_367# N_A_2186_367#_M1030_d
+ N_A_2186_367#_M1009_s N_A_2186_367#_c_1490_n N_A_2186_367#_M1008_g
+ N_A_2186_367#_M1041_g N_A_2186_367#_c_1482_n N_A_2186_367#_c_1483_n
+ N_A_2186_367#_c_1493_n N_A_2186_367#_c_1494_n N_A_2186_367#_c_1495_n
+ N_A_2186_367#_c_1484_n N_A_2186_367#_c_1485_n N_A_2186_367#_c_1486_n
+ N_A_2186_367#_c_1487_n N_A_2186_367#_c_1488_n N_A_2186_367#_c_1489_n
+ PM_SKY130_FD_SC_MS__SDFSTP_2%A_2186_367#
x_PM_SKY130_FD_SC_MS__SDFSTP_2%A_1804_424# N_A_1804_424#_M1001_d
+ N_A_1804_424#_M1036_d N_A_1804_424#_M1003_s N_A_1804_424#_M1010_s
+ N_A_1804_424#_M1013_d N_A_1804_424#_M1030_g N_A_1804_424#_M1009_g
+ N_A_1804_424#_c_1587_n N_A_1804_424#_c_1588_n N_A_1804_424#_M1022_g
+ N_A_1804_424#_M1002_g N_A_1804_424#_c_1602_n N_A_1804_424#_c_1590_n
+ N_A_1804_424#_c_1603_n N_A_1804_424#_c_1604_n N_A_1804_424#_c_1605_n
+ N_A_1804_424#_c_1591_n N_A_1804_424#_c_1606_n N_A_1804_424#_c_1670_n
+ N_A_1804_424#_c_1592_n N_A_1804_424#_c_1607_n N_A_1804_424#_c_1593_n
+ N_A_1804_424#_c_1594_n N_A_1804_424#_c_1595_n N_A_1804_424#_c_1609_n
+ N_A_1804_424#_c_1610_n N_A_1804_424#_c_1611_n N_A_1804_424#_c_1596_n
+ N_A_1804_424#_c_1597_n N_A_1804_424#_c_1598_n N_A_1804_424#_c_1657_n
+ N_A_1804_424#_c_1612_n N_A_1804_424#_c_1613_n N_A_1804_424#_c_1599_n
+ PM_SKY130_FD_SC_MS__SDFSTP_2%A_1804_424#
x_PM_SKY130_FD_SC_MS__SDFSTP_2%A_2611_98# N_A_2611_98#_M1022_s
+ N_A_2611_98#_M1002_s N_A_2611_98#_M1004_g N_A_2611_98#_M1014_g
+ N_A_2611_98#_c_1780_n N_A_2611_98#_M1037_g N_A_2611_98#_M1045_g
+ N_A_2611_98#_c_1782_n N_A_2611_98#_c_1788_n N_A_2611_98#_c_1783_n
+ N_A_2611_98#_c_1784_n N_A_2611_98#_c_1785_n
+ PM_SKY130_FD_SC_MS__SDFSTP_2%A_2611_98#
x_PM_SKY130_FD_SC_MS__SDFSTP_2%VPWR N_VPWR_M1015_d N_VPWR_M1017_d N_VPWR_M1032_d
+ N_VPWR_M1042_d N_VPWR_M1021_d N_VPWR_M1007_s N_VPWR_M1008_d N_VPWR_M1009_d
+ N_VPWR_M1002_d N_VPWR_M1045_d N_VPWR_c_1856_n N_VPWR_c_1857_n N_VPWR_c_1858_n
+ N_VPWR_c_1859_n N_VPWR_c_1860_n N_VPWR_c_1861_n N_VPWR_c_1862_n
+ N_VPWR_c_1863_n N_VPWR_c_1864_n N_VPWR_c_1865_n N_VPWR_c_1866_n
+ N_VPWR_c_1867_n N_VPWR_c_1868_n N_VPWR_c_1869_n N_VPWR_c_1870_n
+ N_VPWR_c_1871_n N_VPWR_c_1872_n N_VPWR_c_1873_n VPWR N_VPWR_c_1874_n
+ N_VPWR_c_1875_n N_VPWR_c_1876_n N_VPWR_c_1877_n N_VPWR_c_1878_n
+ N_VPWR_c_1879_n N_VPWR_c_1880_n N_VPWR_c_1881_n N_VPWR_c_1882_n
+ N_VPWR_c_1883_n N_VPWR_c_1884_n N_VPWR_c_1885_n N_VPWR_c_1855_n
+ PM_SKY130_FD_SC_MS__SDFSTP_2%VPWR
x_PM_SKY130_FD_SC_MS__SDFSTP_2%A_293_464# N_A_293_464#_M1028_d
+ N_A_293_464#_M1024_s N_A_293_464#_M1023_d N_A_293_464#_M1034_s
+ N_A_293_464#_c_2052_n N_A_293_464#_c_2038_n N_A_293_464#_c_2039_n
+ N_A_293_464#_c_2040_n N_A_293_464#_c_2041_n N_A_293_464#_c_2045_n
+ N_A_293_464#_c_2046_n N_A_293_464#_c_2047_n N_A_293_464#_c_2075_n
+ N_A_293_464#_c_2048_n N_A_293_464#_c_2042_n N_A_293_464#_c_2043_n
+ N_A_293_464#_c_2050_n N_A_293_464#_c_2051_n
+ PM_SKY130_FD_SC_MS__SDFSTP_2%A_293_464#
x_PM_SKY130_FD_SC_MS__SDFSTP_2%A_1587_379# N_A_1587_379#_M1000_d
+ N_A_1587_379#_M1003_d N_A_1587_379#_c_2177_n N_A_1587_379#_c_2174_n
+ N_A_1587_379#_c_2190_n N_A_1587_379#_c_2175_n N_A_1587_379#_c_2176_n
+ PM_SKY130_FD_SC_MS__SDFSTP_2%A_1587_379#
x_PM_SKY130_FD_SC_MS__SDFSTP_2%Q N_Q_M1014_d N_Q_M1004_s N_Q_c_2208_n
+ N_Q_c_2213_n N_Q_c_2209_n N_Q_c_2210_n N_Q_c_2211_n Q Q
+ PM_SKY130_FD_SC_MS__SDFSTP_2%Q
x_PM_SKY130_FD_SC_MS__SDFSTP_2%VGND N_VGND_M1043_d N_VGND_M1035_d N_VGND_M1012_d
+ N_VGND_M1020_d N_VGND_M1027_d N_VGND_M1033_s N_VGND_M1025_d N_VGND_M1022_d
+ N_VGND_M1037_s N_VGND_c_2249_n N_VGND_c_2250_n N_VGND_c_2251_n N_VGND_c_2252_n
+ N_VGND_c_2253_n N_VGND_c_2254_n N_VGND_c_2255_n N_VGND_c_2256_n
+ N_VGND_c_2257_n N_VGND_c_2258_n N_VGND_c_2259_n VGND N_VGND_c_2260_n
+ N_VGND_c_2261_n N_VGND_c_2262_n N_VGND_c_2263_n N_VGND_c_2264_n
+ N_VGND_c_2265_n N_VGND_c_2266_n N_VGND_c_2267_n N_VGND_c_2268_n
+ N_VGND_c_2269_n N_VGND_c_2270_n N_VGND_c_2271_n N_VGND_c_2272_n
+ N_VGND_c_2273_n N_VGND_c_2274_n PM_SKY130_FD_SC_MS__SDFSTP_2%VGND
x_PM_SKY130_FD_SC_MS__SDFSTP_2%A_1641_74# N_A_1641_74#_M1029_d
+ N_A_1641_74#_M1001_s N_A_1641_74#_c_2411_n N_A_1641_74#_c_2412_n
+ N_A_1641_74#_c_2413_n N_A_1641_74#_c_2414_n
+ PM_SKY130_FD_SC_MS__SDFSTP_2%A_1641_74#
cc_1 VNB N_SCE_M1043_g 0.0625566f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_2 VNB N_SCE_M1039_g 0.0349556f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.58
cc_3 VNB N_SCE_c_315_n 0.0286809f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.495
cc_4 VNB N_SCE_c_316_n 0.00225026f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.495
cc_5 VNB N_SCE_c_317_n 0.00268133f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.415
cc_6 VNB N_SCE_c_318_n 0.0306519f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.415
cc_7 VNB N_SCE_c_319_n 0.0242476f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.635
cc_8 VNB N_A_27_74#_c_391_n 0.023955f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.58
cc_9 VNB N_A_27_74#_c_392_n 0.0203201f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.065
cc_10 VNB N_A_27_74#_c_393_n 0.0100668f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.415
cc_11 VNB N_A_27_74#_c_394_n 0.0334307f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.415
cc_12 VNB N_A_27_74#_c_395_n 0.0203203f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.58
cc_13 VNB N_A_27_74#_c_396_n 0.0182373f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.47
cc_14 VNB N_D_M1028_g 0.0618257f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.47
cc_15 VNB N_SCD_M1035_g 0.0344632f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.14
cc_16 VNB N_SCD_c_515_n 0.0255215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB SCD 0.00297672f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.14
cc_18 VNB N_SCD_c_517_n 0.0333042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_CLK_M1032_g 0.0070466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB CLK 0.00842451f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_21 VNB N_CLK_c_560_n 0.0323076f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.14
cc_22 VNB N_CLK_c_561_n 0.0200244f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.64
cc_23 VNB N_A_795_74#_c_596_n 0.0120986f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.14
cc_24 VNB N_A_795_74#_c_597_n 0.00683373f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.64
cc_25 VNB N_A_795_74#_M1031_g 0.0362022f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.58
cc_26 VNB N_A_795_74#_c_599_n 0.0279309f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.065
cc_27 VNB N_A_795_74#_c_600_n 0.00949433f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.065
cc_28 VNB N_A_795_74#_c_601_n 0.0175524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_795_74#_c_602_n 0.0168332f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.415
cc_30 VNB N_A_795_74#_c_603_n 0.0148787f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.415
cc_31 VNB N_A_795_74#_c_604_n 0.00400906f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.635
cc_32 VNB N_A_795_74#_c_605_n 0.00168954f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.415
cc_33 VNB N_A_795_74#_c_606_n 0.0170808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_795_74#_c_607_n 0.00264685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_795_74#_c_608_n 0.00341946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_795_74#_c_609_n 0.00339844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_795_74#_c_610_n 0.00752699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_795_74#_c_611_n 0.0169131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_795_74#_c_612_n 0.0051925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_795_74#_c_613_n 2.60503e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_795_74#_c_614_n 0.0241397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_795_74#_c_615_n 0.00785969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_795_74#_c_616_n 0.0126071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_795_74#_c_617_n 0.0186057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1185_55#_c_874_n 0.0173208f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.47
cc_46 VNB N_A_1185_55#_c_875_n 0.0362711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1185_55#_c_876_n 0.00116198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1185_55#_c_877_n 0.00722463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1185_55#_c_878_n 0.00471537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1185_55#_c_879_n 0.0061097f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.635
cc_51 VNB N_A_1185_55#_c_880_n 0.0204767f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.25
cc_52 VNB N_A_991_81#_c_970_n 0.0149666f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.47
cc_53 VNB N_A_991_81#_M1011_g 0.00584511f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_54 VNB N_A_991_81#_c_972_n 0.0180022f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.14
cc_55 VNB N_A_991_81#_M1000_g 0.00637895f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.58
cc_56 VNB N_A_991_81#_c_974_n 0.0168452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_991_81#_M1007_g 0.00566411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_991_81#_c_976_n 0.0170434f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.495
cc_59 VNB N_A_991_81#_c_977_n 0.031795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_991_81#_c_978_n 0.00798345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_991_81#_c_979_n 0.0235266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_991_81#_c_980_n 0.0101867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_991_81#_c_981_n 0.0296742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_991_81#_c_982_n 0.0240823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_991_81#_c_983_n 0.00126724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_991_81#_c_984_n 0.00103134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_991_81#_c_985_n 0.00183906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_991_81#_c_986_n 0.00325464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_991_81#_c_987_n 0.0727754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_SET_B_M1021_g 0.00671558f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.14
cc_71 VNB N_SET_B_M1027_g 0.0373019f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.47
cc_72 VNB N_SET_B_M1025_g 0.0515369f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=1.25
cc_73 VNB N_SET_B_c_1155_n 0.0389494f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.58
cc_74 VNB N_SET_B_c_1156_n 0.00220503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_SET_B_c_1157_n 0.00540182f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.065
cc_76 VNB SET_B 0.0040711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_SET_B_c_1159_n 0.0378364f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.495
cc_78 VNB N_SET_B_c_1160_n 0.0220211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_SET_B_c_1161_n 0.00779184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_608_74#_M1006_g 0.0255853f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_81 VNB N_A_608_74#_c_1285_n 0.0103779f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.58
cc_82 VNB N_A_608_74#_c_1286_n 0.0292071f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.065
cc_83 VNB N_A_608_74#_c_1287_n 0.0103124f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.065
cc_84 VNB N_A_608_74#_M1024_g 0.0272072f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.415
cc_85 VNB N_A_608_74#_M1003_g 0.00187228f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.47
cc_86 VNB N_A_608_74#_c_1290_n 0.0686567f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.415
cc_87 VNB N_A_608_74#_c_1291_n 0.00767386f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.25
cc_88 VNB N_A_608_74#_M1044_g 0.0455489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_608_74#_c_1293_n 0.00838246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_608_74#_c_1294_n 0.0120978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_608_74#_c_1295_n 0.00199494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_608_74#_c_1296_n 0.00302852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_608_74#_c_1297_n 0.0385409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_2186_367#_c_1482_n 0.0218664f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.58
cc_95 VNB N_A_2186_367#_c_1483_n 0.0255406f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.58
cc_96 VNB N_A_2186_367#_c_1484_n 0.00775159f $X=-0.19 $Y=-0.245 $X2=1.96
+ $Y2=1.415
cc_97 VNB N_A_2186_367#_c_1485_n 0.00617016f $X=-0.19 $Y=-0.245 $X2=1.92
+ $Y2=1.495
cc_98 VNB N_A_2186_367#_c_1486_n 0.00238188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_2186_367#_c_1487_n 0.0330841f $X=-0.19 $Y=-0.245 $X2=0.61
+ $Y2=1.635
cc_100 VNB N_A_2186_367#_c_1488_n 0.00377829f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.635
cc_101 VNB N_A_2186_367#_c_1489_n 0.0181222f $X=-0.19 $Y=-0.245 $X2=1.96
+ $Y2=1.415
cc_102 VNB N_A_1804_424#_M1030_g 0.0396191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1804_424#_c_1587_n 0.0812455f $X=-0.19 $Y=-0.245 $X2=1.795
+ $Y2=1.495
cc_104 VNB N_A_1804_424#_c_1588_n 0.0177817f $X=-0.19 $Y=-0.245 $X2=1.92
+ $Y2=1.415
cc_105 VNB N_A_1804_424#_M1002_g 0.00783058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1804_424#_c_1590_n 0.0124338f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.635
cc_107 VNB N_A_1804_424#_c_1591_n 0.00515896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_1804_424#_c_1592_n 0.00497081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_1804_424#_c_1593_n 0.00847186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_1804_424#_c_1594_n 0.0018227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_1804_424#_c_1595_n 0.00246574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_1804_424#_c_1596_n 0.00200957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_1804_424#_c_1597_n 0.0340509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_1804_424#_c_1598_n 0.00765385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_1804_424#_c_1599_n 0.0115341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_2611_98#_M1004_g 5.12161e-19 $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=0.58
cc_117 VNB N_A_2611_98#_M1014_g 0.0212563f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.64
cc_118 VNB N_A_2611_98#_c_1780_n 0.0160455f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=1.25
cc_119 VNB N_A_2611_98#_M1045_g 5.83046e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_2611_98#_c_1782_n 0.00961135f $X=-0.19 $Y=-0.245 $X2=1.795
+ $Y2=1.495
cc_121 VNB N_A_2611_98#_c_1783_n 0.00549082f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=1.58
cc_122 VNB N_A_2611_98#_c_1784_n 0.00102441f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.635
cc_123 VNB N_A_2611_98#_c_1785_n 0.0627395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VPWR_c_1855_n 0.621437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_293_464#_c_2038_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.065
cc_126 VNB N_A_293_464#_c_2039_n 0.0157325f $X=-0.19 $Y=-0.245 $X2=0.61
+ $Y2=2.065
cc_127 VNB N_A_293_464#_c_2040_n 0.00298819f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.065
cc_128 VNB N_A_293_464#_c_2041_n 0.00472436f $X=-0.19 $Y=-0.245 $X2=1.795
+ $Y2=1.495
cc_129 VNB N_A_293_464#_c_2042_n 0.00614445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_A_293_464#_c_2043_n 0.00705683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_Q_c_2208_n 0.00248472f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_132 VNB N_Q_c_2209_n 0.0019936f $X=-0.19 $Y=-0.245 $X2=1.94 $Y2=0.58
cc_133 VNB N_Q_c_2210_n 0.0016018f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.065
cc_134 VNB N_Q_c_2211_n 0.0112378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB Q 0.00712458f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.065
cc_136 VNB N_VGND_c_2249_n 0.00778079f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.495
cc_137 VNB N_VGND_c_2250_n 0.0101978f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.58
cc_138 VNB N_VGND_c_2251_n 0.0201354f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.635
cc_139 VNB N_VGND_c_2252_n 0.00641543f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.25
cc_140 VNB N_VGND_c_2253_n 0.00826914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2254_n 0.0130607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2255_n 0.0163952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2256_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2257_n 0.0444854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2258_n 0.0152199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2259_n 0.0590232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2260_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2261_n 0.0412906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2262_n 0.0293898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2263_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2264_n 0.0345145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2265_n 0.0198784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2266_n 0.00856226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2267_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2268_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2269_n 0.00942782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_2270_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2271_n 0.0702539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_2272_n 0.0234846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_2273_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_VGND_c_2274_n 0.827876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VNB N_A_1641_74#_c_2411_n 0.0024035f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=0.58
cc_163 VNB N_A_1641_74#_c_2412_n 0.017548f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.14
cc_164 VNB N_A_1641_74#_c_2413_n 0.00262272f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.64
cc_165 VNB N_A_1641_74#_c_2414_n 0.00193131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VPB N_SCE_c_320_n 0.0301327f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.99
cc_167 VPB N_SCE_M1015_g 0.0260819f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_168 VPB N_SCE_c_322_n 0.0263646f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.14
cc_169 VPB N_SCE_M1016_g 0.0218933f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_170 VPB SCE 8.61801e-19 $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_171 VPB N_SCE_c_319_n 4.81492e-19 $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.635
cc_172 VPB N_A_27_74#_M1005_g 0.0229139f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_173 VPB N_A_27_74#_c_392_n 0.0305464f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.065
cc_174 VPB N_A_27_74#_c_399_n 0.00362328f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_27_74#_c_400_n 0.0313416f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_176 VPB N_A_27_74#_c_401_n 0.0311143f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.635
cc_177 VPB N_D_M1023_g 0.0244166f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.14
cc_178 VPB N_D_M1028_g 0.0121448f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.47
cc_179 VPB N_D_c_473_n 0.0286108f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_180 VPB N_D_c_474_n 0.00778097f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_181 VPB N_SCD_c_515_n 0.0250802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_SCD_M1017_g 0.0253519f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_183 VPB SCD 0.0027614f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.14
cc_184 VPB N_SCD_c_521_n 0.0315846f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.065
cc_185 VPB N_CLK_M1032_g 0.0252927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_795_74#_M1034_g 0.0432042f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_187 VPB N_A_795_74#_c_596_n 0.00688565f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.14
cc_188 VPB N_A_795_74#_M1019_g 0.0376538f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_795_74#_c_621_n 0.00313813f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_795_74#_c_622_n 0.0228678f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_795_74#_c_623_n 0.00295859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_795_74#_c_608_n 0.00115773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_795_74#_c_625_n 0.00574112f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_795_74#_c_626_n 0.00140676f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_795_74#_c_627_n 0.0230817f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_795_74#_c_628_n 0.00242474f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_795_74#_c_629_n 0.0137064f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_795_74#_c_630_n 0.00177503f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_795_74#_c_631_n 0.00538502f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_795_74#_c_632_n 3.46324e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_795_74#_c_610_n 0.0228475f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_795_74#_c_611_n 0.0174517f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_795_74#_c_635_n 0.00570704f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_795_74#_c_636_n 0.0320872f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_795_74#_c_637_n 0.0182982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_795_74#_c_613_n 0.00399799f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_795_74#_c_614_n 0.00859831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_795_74#_c_615_n 0.0310447f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_1185_55#_M1042_g 0.0330476f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_210 VPB N_A_1185_55#_c_882_n 0.0155588f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=2.065
cc_211 VPB N_A_1185_55#_c_883_n 0.00757992f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.415
cc_212 VPB N_A_1185_55#_c_878_n 0.0246878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_1185_55#_c_885_n 0.00167294f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_991_81#_M1011_g 0.0486719f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_215 VPB N_A_991_81#_M1000_g 0.0234661f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=0.58
cc_216 VPB N_A_991_81#_M1007_g 0.0234586f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_991_81#_c_991_n 0.00407701f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.58
cc_218 VPB N_A_991_81#_c_992_n 6.35236e-19 $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.635
cc_219 VPB N_A_991_81#_c_984_n 0.00962111f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_SET_B_M1021_g 0.04856f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.14
cc_221 VPB N_SET_B_M1013_g 0.0615729f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.14
cc_222 VPB N_SET_B_c_1160_n 0.0169762f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_SET_B_c_1161_n 0.00397329f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_608_74#_M1040_g 0.020919f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_225 VPB N_A_608_74#_c_1299_n 0.0555956f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_608_74#_c_1300_n 0.05851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_608_74#_c_1301_n 0.0123683f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.495
cc_228 VPB N_A_608_74#_M1018_g 0.0294856f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_608_74#_c_1303_n 0.286876f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_608_74#_M1003_g 0.0384813f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.47
cc_231 VPB N_A_608_74#_c_1305_n 0.0292545f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_608_74#_c_1306_n 0.0183198f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_608_74#_c_1307_n 0.0146072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_608_74#_c_1308_n 0.0100299f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_608_74#_c_1309_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_608_74#_c_1310_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_A_608_74#_c_1294_n 0.00356464f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_A_608_74#_c_1312_n 0.011513f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_A_608_74#_c_1313_n 0.00459351f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_A_608_74#_c_1295_n 8.82238e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_A_608_74#_c_1297_n 0.00682341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_A_2186_367#_c_1490_n 0.00507685f $X=-0.19 $Y=1.66 $X2=0.495
+ $Y2=1.47
cc_243 VPB N_A_2186_367#_M1008_g 0.03914f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_244 VPB N_A_2186_367#_c_1482_n 0.0105007f $X=-0.19 $Y=1.66 $X2=1.94 $Y2=0.58
cc_245 VPB N_A_2186_367#_c_1493_n 0.00755624f $X=-0.19 $Y=1.66 $X2=0.61
+ $Y2=2.065
cc_246 VPB N_A_2186_367#_c_1494_n 0.00863008f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_2186_367#_c_1495_n 0.0037727f $X=-0.19 $Y=1.66 $X2=1.795
+ $Y2=1.495
cc_248 VPB N_A_2186_367#_c_1485_n 0.0126613f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.495
cc_249 VPB N_A_1804_424#_M1009_g 0.0466238f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.065
cc_250 VPB N_A_1804_424#_M1002_g 0.035459f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_A_1804_424#_c_1602_n 0.0213618f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.635
cc_252 VPB N_A_1804_424#_c_1603_n 0.0067705f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.415
cc_253 VPB N_A_1804_424#_c_1604_n 0.00739359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_A_1804_424#_c_1605_n 0.00279745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_A_1804_424#_c_1606_n 9.49732e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_A_1804_424#_c_1607_n 0.0025529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_A_1804_424#_c_1595_n 0.00611054f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_A_1804_424#_c_1609_n 0.0080375f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_A_1804_424#_c_1610_n 0.0165649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_A_1804_424#_c_1611_n 0.00210961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_A_1804_424#_c_1612_n 0.0111974f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_A_1804_424#_c_1613_n 0.021011f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_A_1804_424#_c_1599_n 0.0294988f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_A_2611_98#_M1004_g 0.0234586f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_265 VPB N_A_2611_98#_M1045_g 0.0257815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_A_2611_98#_c_1788_n 0.0167354f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.415
cc_267 VPB N_VPWR_c_1856_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1857_n 0.00963743f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.635
cc_269 VPB N_VPWR_c_1858_n 0.0196669f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.415
cc_270 VPB N_VPWR_c_1859_n 0.00339692f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1860_n 0.00554482f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1861_n 0.0125407f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1862_n 0.017862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1863_n 0.00554449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1864_n 0.0110131f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1865_n 0.0119849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1866_n 0.0116777f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1867_n 0.0347252f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_1868_n 0.0541194f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_VPWR_c_1869_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_VPWR_c_1870_n 0.027717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_VPWR_c_1871_n 0.00223798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_283 VPB N_VPWR_c_1872_n 0.019428f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_284 VPB N_VPWR_c_1873_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 VPB N_VPWR_c_1874_n 0.0180274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_286 VPB N_VPWR_c_1875_n 0.0455708f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_287 VPB N_VPWR_c_1876_n 0.0611503f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_288 VPB N_VPWR_c_1877_n 0.0328287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_289 VPB N_VPWR_c_1878_n 0.0196104f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_290 VPB N_VPWR_c_1879_n 0.0173363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_291 VPB N_VPWR_c_1880_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_292 VPB N_VPWR_c_1881_n 0.00631651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_293 VPB N_VPWR_c_1882_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_294 VPB N_VPWR_c_1883_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_295 VPB N_VPWR_c_1884_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_296 VPB N_VPWR_c_1885_n 0.00545601f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_297 VPB N_VPWR_c_1855_n 0.112692f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_298 VPB N_A_293_464#_c_2041_n 0.00529078f $X=-0.19 $Y=1.66 $X2=1.795
+ $Y2=1.495
cc_299 VPB N_A_293_464#_c_2045_n 0.00531638f $X=-0.19 $Y=1.66 $X2=0.805
+ $Y2=1.495
cc_300 VPB N_A_293_464#_c_2046_n 0.006234f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.415
cc_301 VPB N_A_293_464#_c_2047_n 0.00165521f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_302 VPB N_A_293_464#_c_2048_n 0.0123075f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.635
cc_303 VPB N_A_293_464#_c_2043_n 0.00207118f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_304 VPB N_A_293_464#_c_2050_n 0.00658745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_305 VPB N_A_293_464#_c_2051_n 0.00494889f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_306 VPB N_A_1587_379#_c_2174_n 0.0171101f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.14
cc_307 VPB N_A_1587_379#_c_2175_n 0.00219713f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_308 VPB N_A_1587_379#_c_2176_n 0.00693087f $X=-0.19 $Y=1.66 $X2=0.505
+ $Y2=2.065
cc_309 VPB N_Q_c_2213_n 0.00229053f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_310 VPB Q 0.00754175f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=2.065
cc_311 VPB Q 0.0173729f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.065
cc_312 N_SCE_M1043_g N_A_27_74#_c_391_n 0.0115261f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_313 N_SCE_M1043_g N_A_27_74#_c_392_n 0.00757393f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_314 N_SCE_c_316_n N_A_27_74#_c_392_n 0.0124456f $X=0.805 $Y=1.495 $X2=0 $Y2=0
cc_315 SCE N_A_27_74#_c_392_n 0.0386025f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_316 N_SCE_c_319_n N_A_27_74#_c_392_n 0.0229708f $X=0.64 $Y=1.635 $X2=0 $Y2=0
cc_317 N_SCE_M1015_g N_A_27_74#_c_407_n 0.0129619f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_318 N_SCE_c_322_n N_A_27_74#_c_407_n 6.1916e-19 $X=0.955 $Y=2.14 $X2=0 $Y2=0
cc_319 N_SCE_M1016_g N_A_27_74#_c_407_n 0.01765f $X=0.955 $Y=2.64 $X2=0 $Y2=0
cc_320 SCE N_A_27_74#_c_407_n 0.0223758f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_321 N_SCE_M1043_g N_A_27_74#_c_393_n 0.0166195f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_322 N_SCE_c_315_n N_A_27_74#_c_393_n 0.030574f $X=1.795 $Y=1.495 $X2=0 $Y2=0
cc_323 N_SCE_c_316_n N_A_27_74#_c_393_n 0.0272015f $X=0.805 $Y=1.495 $X2=0 $Y2=0
cc_324 N_SCE_c_319_n N_A_27_74#_c_393_n 0.00145805f $X=0.64 $Y=1.635 $X2=0 $Y2=0
cc_325 N_SCE_M1043_g N_A_27_74#_c_394_n 0.0123124f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_326 N_SCE_c_315_n N_A_27_74#_c_394_n 0.00793591f $X=1.795 $Y=1.495 $X2=0
+ $Y2=0
cc_327 N_SCE_c_317_n N_A_27_74#_c_399_n 0.0145428f $X=1.96 $Y=1.415 $X2=0 $Y2=0
cc_328 N_SCE_c_318_n N_A_27_74#_c_399_n 3.1381e-19 $X=1.96 $Y=1.415 $X2=0 $Y2=0
cc_329 N_SCE_c_317_n N_A_27_74#_c_400_n 3.16809e-19 $X=1.96 $Y=1.415 $X2=0 $Y2=0
cc_330 N_SCE_c_318_n N_A_27_74#_c_400_n 0.0184304f $X=1.96 $Y=1.415 $X2=0 $Y2=0
cc_331 N_SCE_M1043_g N_A_27_74#_c_395_n 0.00874187f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_332 N_SCE_c_319_n N_A_27_74#_c_395_n 2.24402e-19 $X=0.64 $Y=1.635 $X2=0 $Y2=0
cc_333 N_SCE_M1015_g N_A_27_74#_c_401_n 8.45069e-19 $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_334 N_SCE_M1043_g N_A_27_74#_c_396_n 0.0139046f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_335 N_SCE_M1016_g N_D_M1023_g 0.0522348f $X=0.955 $Y=2.64 $X2=0 $Y2=0
cc_336 N_SCE_M1039_g N_D_M1028_g 0.0284734f $X=1.94 $Y=0.58 $X2=0 $Y2=0
cc_337 N_SCE_c_315_n N_D_M1028_g 0.015938f $X=1.795 $Y=1.495 $X2=0 $Y2=0
cc_338 N_SCE_c_317_n N_D_M1028_g 0.00118673f $X=1.96 $Y=1.415 $X2=0 $Y2=0
cc_339 N_SCE_c_318_n N_D_M1028_g 0.0212609f $X=1.96 $Y=1.415 $X2=0 $Y2=0
cc_340 SCE N_D_M1028_g 0.00116396f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_341 N_SCE_c_319_n N_D_M1028_g 0.00639795f $X=0.64 $Y=1.635 $X2=0 $Y2=0
cc_342 N_SCE_c_320_n N_D_c_473_n 0.00384203f $X=0.61 $Y=1.99 $X2=0 $Y2=0
cc_343 N_SCE_c_322_n N_D_c_473_n 0.0102797f $X=0.955 $Y=2.14 $X2=0 $Y2=0
cc_344 N_SCE_c_315_n N_D_c_473_n 0.00439769f $X=1.795 $Y=1.495 $X2=0 $Y2=0
cc_345 SCE N_D_c_473_n 2.74008e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_346 N_SCE_c_320_n N_D_c_474_n 0.00146537f $X=0.61 $Y=1.99 $X2=0 $Y2=0
cc_347 N_SCE_c_322_n N_D_c_474_n 0.00182065f $X=0.955 $Y=2.14 $X2=0 $Y2=0
cc_348 N_SCE_c_315_n N_D_c_474_n 0.0291812f $X=1.795 $Y=1.495 $X2=0 $Y2=0
cc_349 SCE N_D_c_474_n 0.0180473f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_350 N_SCE_M1039_g N_SCD_M1035_g 0.0368573f $X=1.94 $Y=0.58 $X2=0 $Y2=0
cc_351 N_SCE_c_317_n N_SCD_c_517_n 2.87119e-19 $X=1.96 $Y=1.415 $X2=0 $Y2=0
cc_352 N_SCE_c_318_n N_SCD_c_517_n 0.0204387f $X=1.96 $Y=1.415 $X2=0 $Y2=0
cc_353 N_SCE_M1015_g N_VPWR_c_1856_n 0.0112582f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_354 N_SCE_M1016_g N_VPWR_c_1856_n 0.0104907f $X=0.955 $Y=2.64 $X2=0 $Y2=0
cc_355 N_SCE_M1015_g N_VPWR_c_1874_n 0.00460063f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_356 N_SCE_M1016_g N_VPWR_c_1875_n 0.00460063f $X=0.955 $Y=2.64 $X2=0 $Y2=0
cc_357 N_SCE_M1015_g N_VPWR_c_1855_n 0.00464602f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_358 N_SCE_M1016_g N_VPWR_c_1855_n 0.00460677f $X=0.955 $Y=2.64 $X2=0 $Y2=0
cc_359 N_SCE_M1016_g N_A_293_464#_c_2052_n 7.0025e-19 $X=0.955 $Y=2.64 $X2=0
+ $Y2=0
cc_360 N_SCE_M1039_g N_A_293_464#_c_2038_n 0.0125369f $X=1.94 $Y=0.58 $X2=0
+ $Y2=0
cc_361 N_SCE_M1039_g N_A_293_464#_c_2039_n 0.0111573f $X=1.94 $Y=0.58 $X2=0
+ $Y2=0
cc_362 N_SCE_c_317_n N_A_293_464#_c_2039_n 0.0111296f $X=1.96 $Y=1.415 $X2=0
+ $Y2=0
cc_363 N_SCE_c_318_n N_A_293_464#_c_2039_n 0.0032473f $X=1.96 $Y=1.415 $X2=0
+ $Y2=0
cc_364 N_SCE_M1039_g N_A_293_464#_c_2040_n 0.00274486f $X=1.94 $Y=0.58 $X2=0
+ $Y2=0
cc_365 N_SCE_c_315_n N_A_293_464#_c_2040_n 0.0123012f $X=1.795 $Y=1.495 $X2=0
+ $Y2=0
cc_366 N_SCE_c_317_n N_A_293_464#_c_2040_n 0.00785342f $X=1.96 $Y=1.415 $X2=0
+ $Y2=0
cc_367 N_SCE_c_318_n N_A_293_464#_c_2040_n 5.46117e-19 $X=1.96 $Y=1.415 $X2=0
+ $Y2=0
cc_368 N_SCE_M1039_g N_A_293_464#_c_2041_n 0.00343685f $X=1.94 $Y=0.58 $X2=0
+ $Y2=0
cc_369 N_SCE_c_317_n N_A_293_464#_c_2041_n 0.0242834f $X=1.96 $Y=1.415 $X2=0
+ $Y2=0
cc_370 N_SCE_c_318_n N_A_293_464#_c_2041_n 0.00204642f $X=1.96 $Y=1.415 $X2=0
+ $Y2=0
cc_371 N_SCE_M1043_g N_VGND_c_2249_n 0.00572943f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_372 N_SCE_M1039_g N_VGND_c_2250_n 0.00172001f $X=1.94 $Y=0.58 $X2=0 $Y2=0
cc_373 N_SCE_M1043_g N_VGND_c_2260_n 0.00434272f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_374 N_SCE_M1039_g N_VGND_c_2261_n 0.00434272f $X=1.94 $Y=0.58 $X2=0 $Y2=0
cc_375 N_SCE_M1043_g N_VGND_c_2274_n 0.00825349f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_376 N_SCE_M1039_g N_VGND_c_2274_n 0.00821825f $X=1.94 $Y=0.58 $X2=0 $Y2=0
cc_377 N_A_27_74#_M1005_g N_D_M1023_g 0.0250203f $X=2.005 $Y=2.64 $X2=0 $Y2=0
cc_378 N_A_27_74#_c_407_n N_D_M1023_g 0.0136825f $X=1.795 $Y=2.405 $X2=0 $Y2=0
cc_379 N_A_27_74#_c_399_n N_D_M1023_g 0.00322627f $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_380 N_A_27_74#_c_400_n N_D_M1023_g 3.90461e-19 $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_381 N_A_27_74#_c_393_n N_D_M1028_g 0.00157925f $X=1.06 $Y=1.065 $X2=0 $Y2=0
cc_382 N_A_27_74#_c_394_n N_D_M1028_g 0.0196496f $X=1.06 $Y=1.065 $X2=0 $Y2=0
cc_383 N_A_27_74#_c_396_n N_D_M1028_g 0.0336314f $X=1.06 $Y=0.9 $X2=0 $Y2=0
cc_384 N_A_27_74#_c_407_n N_D_c_473_n 0.00303821f $X=1.795 $Y=2.405 $X2=0 $Y2=0
cc_385 N_A_27_74#_c_399_n N_D_c_473_n 4.04344e-19 $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_386 N_A_27_74#_c_400_n N_D_c_473_n 0.0201404f $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_387 N_A_27_74#_c_407_n N_D_c_474_n 0.0324243f $X=1.795 $Y=2.405 $X2=0 $Y2=0
cc_388 N_A_27_74#_c_399_n N_D_c_474_n 0.0205429f $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_389 N_A_27_74#_c_400_n N_D_c_474_n 0.00111057f $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_390 N_A_27_74#_c_399_n N_SCD_c_515_n 4.37507e-19 $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_391 N_A_27_74#_c_400_n N_SCD_c_515_n 0.0204031f $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_392 N_A_27_74#_M1005_g N_SCD_M1017_g 0.048695f $X=2.005 $Y=2.64 $X2=0 $Y2=0
cc_393 N_A_27_74#_c_407_n N_VPWR_M1015_d 0.00308156f $X=1.795 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_394 N_A_27_74#_c_407_n N_VPWR_c_1856_n 0.0166513f $X=1.795 $Y=2.405 $X2=0
+ $Y2=0
cc_395 N_A_27_74#_c_401_n N_VPWR_c_1856_n 0.0112185f $X=0.28 $Y=2.475 $X2=0
+ $Y2=0
cc_396 N_A_27_74#_c_401_n N_VPWR_c_1874_n 0.0110622f $X=0.28 $Y=2.475 $X2=0
+ $Y2=0
cc_397 N_A_27_74#_M1005_g N_VPWR_c_1875_n 0.00361052f $X=2.005 $Y=2.64 $X2=0
+ $Y2=0
cc_398 N_A_27_74#_M1005_g N_VPWR_c_1855_n 0.00442185f $X=2.005 $Y=2.64 $X2=0
+ $Y2=0
cc_399 N_A_27_74#_c_407_n N_VPWR_c_1855_n 0.0238901f $X=1.795 $Y=2.405 $X2=0
+ $Y2=0
cc_400 N_A_27_74#_c_401_n N_VPWR_c_1855_n 0.00915799f $X=0.28 $Y=2.475 $X2=0
+ $Y2=0
cc_401 N_A_27_74#_c_407_n A_209_464# 0.00387589f $X=1.795 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_402 N_A_27_74#_c_407_n N_A_293_464#_M1023_d 0.0127809f $X=1.795 $Y=2.405
+ $X2=0 $Y2=0
cc_403 N_A_27_74#_M1005_g N_A_293_464#_c_2052_n 0.0161913f $X=2.005 $Y=2.64
+ $X2=0 $Y2=0
cc_404 N_A_27_74#_c_407_n N_A_293_464#_c_2052_n 0.0368886f $X=1.795 $Y=2.405
+ $X2=0 $Y2=0
cc_405 N_A_27_74#_c_400_n N_A_293_464#_c_2052_n 3.51567e-19 $X=1.96 $Y=1.995
+ $X2=0 $Y2=0
cc_406 N_A_27_74#_c_393_n N_A_293_464#_c_2038_n 3.9435e-19 $X=1.06 $Y=1.065
+ $X2=0 $Y2=0
cc_407 N_A_27_74#_c_396_n N_A_293_464#_c_2038_n 0.00202258f $X=1.06 $Y=0.9 $X2=0
+ $Y2=0
cc_408 N_A_27_74#_c_393_n N_A_293_464#_c_2040_n 0.00831735f $X=1.06 $Y=1.065
+ $X2=0 $Y2=0
cc_409 N_A_27_74#_M1005_g N_A_293_464#_c_2041_n 0.0056003f $X=2.005 $Y=2.64
+ $X2=0 $Y2=0
cc_410 N_A_27_74#_c_407_n N_A_293_464#_c_2041_n 0.0133253f $X=1.795 $Y=2.405
+ $X2=0 $Y2=0
cc_411 N_A_27_74#_c_399_n N_A_293_464#_c_2041_n 0.0359857f $X=1.96 $Y=1.995
+ $X2=0 $Y2=0
cc_412 N_A_27_74#_c_400_n N_A_293_464#_c_2041_n 0.00204642f $X=1.96 $Y=1.995
+ $X2=0 $Y2=0
cc_413 N_A_27_74#_M1005_g N_A_293_464#_c_2075_n 2.71809e-19 $X=2.005 $Y=2.64
+ $X2=0 $Y2=0
cc_414 N_A_27_74#_c_391_n N_VGND_c_2249_n 0.0132122f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_415 N_A_27_74#_c_393_n N_VGND_c_2249_n 0.0292604f $X=1.06 $Y=1.065 $X2=0
+ $Y2=0
cc_416 N_A_27_74#_c_394_n N_VGND_c_2249_n 0.00320405f $X=1.06 $Y=1.065 $X2=0
+ $Y2=0
cc_417 N_A_27_74#_c_396_n N_VGND_c_2249_n 0.015423f $X=1.06 $Y=0.9 $X2=0 $Y2=0
cc_418 N_A_27_74#_c_391_n N_VGND_c_2260_n 0.0145639f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_419 N_A_27_74#_c_396_n N_VGND_c_2261_n 0.00383152f $X=1.06 $Y=0.9 $X2=0 $Y2=0
cc_420 N_A_27_74#_c_391_n N_VGND_c_2274_n 0.0119984f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_421 N_A_27_74#_c_396_n N_VGND_c_2274_n 0.0075725f $X=1.06 $Y=0.9 $X2=0 $Y2=0
cc_422 N_D_M1023_g N_VPWR_c_1856_n 0.00159211f $X=1.375 $Y=2.64 $X2=0 $Y2=0
cc_423 N_D_M1023_g N_VPWR_c_1875_n 0.00521639f $X=1.375 $Y=2.64 $X2=0 $Y2=0
cc_424 N_D_M1023_g N_VPWR_c_1855_n 0.00538257f $X=1.375 $Y=2.64 $X2=0 $Y2=0
cc_425 N_D_M1023_g N_A_293_464#_c_2052_n 0.00954817f $X=1.375 $Y=2.64 $X2=0
+ $Y2=0
cc_426 N_D_M1028_g N_A_293_464#_c_2038_n 0.0116998f $X=1.51 $Y=0.58 $X2=0 $Y2=0
cc_427 N_D_M1028_g N_A_293_464#_c_2040_n 0.00483064f $X=1.51 $Y=0.58 $X2=0 $Y2=0
cc_428 N_D_M1028_g N_A_293_464#_c_2041_n 0.00511872f $X=1.51 $Y=0.58 $X2=0 $Y2=0
cc_429 N_D_c_474_n N_A_293_464#_c_2041_n 2.57555e-19 $X=1.42 $Y=1.985 $X2=0
+ $Y2=0
cc_430 N_D_M1028_g N_VGND_c_2249_n 0.00149152f $X=1.51 $Y=0.58 $X2=0 $Y2=0
cc_431 N_D_M1028_g N_VGND_c_2261_n 0.00434272f $X=1.51 $Y=0.58 $X2=0 $Y2=0
cc_432 N_D_M1028_g N_VGND_c_2274_n 0.00821077f $X=1.51 $Y=0.58 $X2=0 $Y2=0
cc_433 N_SCD_c_515_n N_CLK_M1032_g 0.00697845f $X=2.582 $Y=1.903 $X2=0 $Y2=0
cc_434 N_SCD_c_517_n N_CLK_c_560_n 0.00730373f $X=2.665 $Y=1.305 $X2=0 $Y2=0
cc_435 N_SCD_c_517_n N_CLK_c_561_n 0.00140608f $X=2.665 $Y=1.305 $X2=0 $Y2=0
cc_436 N_SCD_M1035_g N_A_608_74#_c_1293_n 0.00901831f $X=2.41 $Y=0.58 $X2=0
+ $Y2=0
cc_437 SCD N_A_608_74#_c_1294_n 0.0474887f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_438 N_SCD_c_517_n N_A_608_74#_c_1294_n 0.00687498f $X=2.665 $Y=1.305 $X2=0
+ $Y2=0
cc_439 N_SCD_c_515_n N_A_608_74#_c_1313_n 0.00301067f $X=2.582 $Y=1.903 $X2=0
+ $Y2=0
cc_440 SCD N_A_608_74#_c_1313_n 0.0196463f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_441 N_SCD_M1017_g N_VPWR_c_1857_n 0.00819721f $X=2.425 $Y=2.64 $X2=0 $Y2=0
cc_442 N_SCD_M1017_g N_VPWR_c_1875_n 0.00387257f $X=2.425 $Y=2.64 $X2=0 $Y2=0
cc_443 N_SCD_M1017_g N_VPWR_c_1855_n 0.00490016f $X=2.425 $Y=2.64 $X2=0 $Y2=0
cc_444 N_SCD_M1017_g N_A_293_464#_c_2052_n 2.74757e-19 $X=2.425 $Y=2.64 $X2=0
+ $Y2=0
cc_445 N_SCD_M1035_g N_A_293_464#_c_2038_n 0.00199239f $X=2.41 $Y=0.58 $X2=0
+ $Y2=0
cc_446 N_SCD_M1035_g N_A_293_464#_c_2039_n 0.00850446f $X=2.41 $Y=0.58 $X2=0
+ $Y2=0
cc_447 N_SCD_M1035_g N_A_293_464#_c_2041_n 0.00172798f $X=2.41 $Y=0.58 $X2=0
+ $Y2=0
cc_448 N_SCD_c_515_n N_A_293_464#_c_2041_n 0.0148573f $X=2.582 $Y=1.903 $X2=0
+ $Y2=0
cc_449 N_SCD_M1017_g N_A_293_464#_c_2041_n 0.0113817f $X=2.425 $Y=2.64 $X2=0
+ $Y2=0
cc_450 SCD N_A_293_464#_c_2041_n 0.069827f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_451 N_SCD_c_517_n N_A_293_464#_c_2041_n 0.0060148f $X=2.665 $Y=1.305 $X2=0
+ $Y2=0
cc_452 N_SCD_c_521_n N_A_293_464#_c_2041_n 0.00572276f $X=2.665 $Y=1.985 $X2=0
+ $Y2=0
cc_453 N_SCD_M1017_g N_A_293_464#_c_2045_n 0.0149256f $X=2.425 $Y=2.64 $X2=0
+ $Y2=0
cc_454 SCD N_A_293_464#_c_2045_n 0.00990286f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_455 N_SCD_c_521_n N_A_293_464#_c_2045_n 0.00306015f $X=2.665 $Y=1.985 $X2=0
+ $Y2=0
cc_456 N_SCD_M1017_g N_A_293_464#_c_2075_n 0.0126663f $X=2.425 $Y=2.64 $X2=0
+ $Y2=0
cc_457 N_SCD_M1017_g N_A_293_464#_c_2048_n 0.00476293f $X=2.425 $Y=2.64 $X2=0
+ $Y2=0
cc_458 N_SCD_M1035_g N_VGND_c_2250_n 0.0135277f $X=2.41 $Y=0.58 $X2=0 $Y2=0
cc_459 SCD N_VGND_c_2250_n 0.0100559f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_460 N_SCD_c_517_n N_VGND_c_2250_n 0.00355058f $X=2.665 $Y=1.305 $X2=0 $Y2=0
cc_461 N_SCD_M1035_g N_VGND_c_2261_n 0.00383152f $X=2.41 $Y=0.58 $X2=0 $Y2=0
cc_462 N_SCD_M1035_g N_VGND_c_2274_n 0.00757998f $X=2.41 $Y=0.58 $X2=0 $Y2=0
cc_463 CLK N_A_608_74#_M1006_g 0.00597538f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_464 N_CLK_c_560_n N_A_608_74#_M1006_g 0.0174253f $X=3.42 $Y=1.385 $X2=0 $Y2=0
cc_465 N_CLK_c_561_n N_A_608_74#_M1006_g 0.0175799f $X=3.42 $Y=1.22 $X2=0 $Y2=0
cc_466 N_CLK_M1032_g N_A_608_74#_M1040_g 0.0512489f $X=3.485 $Y=2.4 $X2=0 $Y2=0
cc_467 N_CLK_c_561_n N_A_608_74#_c_1293_n 0.00580215f $X=3.42 $Y=1.22 $X2=0
+ $Y2=0
cc_468 N_CLK_M1032_g N_A_608_74#_c_1294_n 0.00564264f $X=3.485 $Y=2.4 $X2=0
+ $Y2=0
cc_469 CLK N_A_608_74#_c_1294_n 0.0284508f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_470 N_CLK_c_560_n N_A_608_74#_c_1294_n 0.00287216f $X=3.42 $Y=1.385 $X2=0
+ $Y2=0
cc_471 N_CLK_c_561_n N_A_608_74#_c_1294_n 0.00371193f $X=3.42 $Y=1.22 $X2=0
+ $Y2=0
cc_472 N_CLK_M1032_g N_A_608_74#_c_1312_n 0.0130096f $X=3.485 $Y=2.4 $X2=0 $Y2=0
cc_473 CLK N_A_608_74#_c_1312_n 0.0227845f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_474 N_CLK_c_560_n N_A_608_74#_c_1312_n 0.00405624f $X=3.42 $Y=1.385 $X2=0
+ $Y2=0
cc_475 N_CLK_M1032_g N_A_608_74#_c_1295_n 0.00156138f $X=3.485 $Y=2.4 $X2=0
+ $Y2=0
cc_476 CLK N_A_608_74#_c_1295_n 0.0161169f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_477 CLK N_A_608_74#_c_1296_n 0.00294872f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_478 N_CLK_c_560_n N_A_608_74#_c_1296_n 0.00116809f $X=3.42 $Y=1.385 $X2=0
+ $Y2=0
cc_479 N_CLK_c_561_n N_A_608_74#_c_1296_n 0.00232554f $X=3.42 $Y=1.22 $X2=0
+ $Y2=0
cc_480 N_CLK_M1032_g N_A_608_74#_c_1297_n 0.00717734f $X=3.485 $Y=2.4 $X2=0
+ $Y2=0
cc_481 N_CLK_M1032_g N_VPWR_c_1857_n 0.0043823f $X=3.485 $Y=2.4 $X2=0 $Y2=0
cc_482 N_CLK_M1032_g N_VPWR_c_1858_n 0.00460063f $X=3.485 $Y=2.4 $X2=0 $Y2=0
cc_483 N_CLK_M1032_g N_VPWR_c_1859_n 0.0174569f $X=3.485 $Y=2.4 $X2=0 $Y2=0
cc_484 N_CLK_M1032_g N_VPWR_c_1855_n 0.00913687f $X=3.485 $Y=2.4 $X2=0 $Y2=0
cc_485 N_CLK_M1032_g N_A_293_464#_c_2046_n 0.0176054f $X=3.485 $Y=2.4 $X2=0
+ $Y2=0
cc_486 N_CLK_M1032_g N_A_293_464#_c_2048_n 0.00754259f $X=3.485 $Y=2.4 $X2=0
+ $Y2=0
cc_487 N_CLK_c_561_n N_VGND_c_2250_n 0.00333233f $X=3.42 $Y=1.22 $X2=0 $Y2=0
cc_488 N_CLK_c_561_n N_VGND_c_2251_n 0.00434272f $X=3.42 $Y=1.22 $X2=0 $Y2=0
cc_489 CLK N_VGND_c_2252_n 0.0164658f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_490 N_CLK_c_560_n N_VGND_c_2252_n 4.19963e-19 $X=3.42 $Y=1.385 $X2=0 $Y2=0
cc_491 N_CLK_c_561_n N_VGND_c_2252_n 0.00659657f $X=3.42 $Y=1.22 $X2=0 $Y2=0
cc_492 N_CLK_c_561_n N_VGND_c_2274_n 0.00825771f $X=3.42 $Y=1.22 $X2=0 $Y2=0
cc_493 N_A_795_74#_M1031_g N_A_1185_55#_c_874_n 0.0474535f $X=5.64 $Y=0.615
+ $X2=0 $Y2=0
cc_494 N_A_795_74#_c_625_n N_A_1185_55#_M1042_g 0.00134246f $X=5.645 $Y=2.255
+ $X2=0 $Y2=0
cc_495 N_A_795_74#_c_626_n N_A_1185_55#_M1042_g 0.00730577f $X=5.645 $Y=2.895
+ $X2=0 $Y2=0
cc_496 N_A_795_74#_c_627_n N_A_1185_55#_M1042_g 0.0188198f $X=6.515 $Y=2.17
+ $X2=0 $Y2=0
cc_497 N_A_795_74#_c_628_n N_A_1185_55#_M1042_g 0.00358158f $X=6.6 $Y=2.905
+ $X2=0 $Y2=0
cc_498 N_A_795_74#_M1031_g N_A_1185_55#_c_875_n 0.0118644f $X=5.64 $Y=0.615
+ $X2=0 $Y2=0
cc_499 N_A_795_74#_M1031_g N_A_1185_55#_c_876_n 0.00159877f $X=5.64 $Y=0.615
+ $X2=0 $Y2=0
cc_500 N_A_795_74#_c_627_n N_A_1185_55#_c_882_n 0.0138611f $X=6.515 $Y=2.17
+ $X2=0 $Y2=0
cc_501 N_A_795_74#_c_631_n N_A_1185_55#_c_882_n 0.00157945f $X=7.28 $Y=2.905
+ $X2=0 $Y2=0
cc_502 N_A_795_74#_c_632_n N_A_1185_55#_c_882_n 0.0133719f $X=7.365 $Y=1.81
+ $X2=0 $Y2=0
cc_503 N_A_795_74#_M1031_g N_A_1185_55#_c_896_n 5.16138e-19 $X=5.64 $Y=0.615
+ $X2=0 $Y2=0
cc_504 N_A_795_74#_c_627_n N_A_1185_55#_c_883_n 0.0135839f $X=6.515 $Y=2.17
+ $X2=0 $Y2=0
cc_505 N_A_795_74#_c_628_n N_A_1185_55#_c_883_n 0.0184532f $X=6.6 $Y=2.905 $X2=0
+ $Y2=0
cc_506 N_A_795_74#_c_629_n N_A_1185_55#_c_883_n 0.0127728f $X=7.195 $Y=2.99
+ $X2=0 $Y2=0
cc_507 N_A_795_74#_c_631_n N_A_1185_55#_c_883_n 0.0580551f $X=7.28 $Y=2.905
+ $X2=0 $Y2=0
cc_508 N_A_795_74#_c_625_n N_A_1185_55#_c_878_n 0.00116556f $X=5.645 $Y=2.255
+ $X2=0 $Y2=0
cc_509 N_A_795_74#_c_627_n N_A_1185_55#_c_878_n 0.00367368f $X=6.515 $Y=2.17
+ $X2=0 $Y2=0
cc_510 N_A_795_74#_c_615_n N_A_1185_55#_c_878_n 0.0259356f $X=5.565 $Y=1.655
+ $X2=0 $Y2=0
cc_511 N_A_795_74#_c_625_n N_A_1185_55#_c_885_n 0.0130405f $X=5.645 $Y=2.255
+ $X2=0 $Y2=0
cc_512 N_A_795_74#_c_627_n N_A_1185_55#_c_885_n 0.0415848f $X=6.515 $Y=2.17
+ $X2=0 $Y2=0
cc_513 N_A_795_74#_c_615_n N_A_1185_55#_c_885_n 2.48241e-19 $X=5.565 $Y=1.655
+ $X2=0 $Y2=0
cc_514 N_A_795_74#_c_597_n N_A_1185_55#_c_880_n 0.0118644f $X=5.625 $Y=1.35
+ $X2=0 $Y2=0
cc_515 N_A_795_74#_c_615_n N_A_1185_55#_c_880_n 0.00426508f $X=5.565 $Y=1.655
+ $X2=0 $Y2=0
cc_516 N_A_795_74#_c_606_n N_A_991_81#_M1024_d 2.28826e-19 $X=5 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_517 N_A_795_74#_c_609_n N_A_991_81#_M1024_d 0.00589878f $X=5.085 $Y=1.015
+ $X2=-0.19 $Y2=-0.245
cc_518 N_A_795_74#_c_627_n N_A_991_81#_M1011_g 0.00617207f $X=6.515 $Y=2.17
+ $X2=0 $Y2=0
cc_519 N_A_795_74#_c_628_n N_A_991_81#_M1011_g 0.0160819f $X=6.6 $Y=2.905 $X2=0
+ $Y2=0
cc_520 N_A_795_74#_c_629_n N_A_991_81#_M1011_g 0.00295426f $X=7.195 $Y=2.99
+ $X2=0 $Y2=0
cc_521 N_A_795_74#_c_631_n N_A_991_81#_M1011_g 7.02825e-19 $X=7.28 $Y=2.905
+ $X2=0 $Y2=0
cc_522 N_A_795_74#_c_632_n N_A_991_81#_M1011_g 2.30351e-19 $X=7.365 $Y=1.81
+ $X2=0 $Y2=0
cc_523 N_A_795_74#_c_631_n N_A_991_81#_M1000_g 0.00397697f $X=7.28 $Y=2.905
+ $X2=0 $Y2=0
cc_524 N_A_795_74#_c_637_n N_A_991_81#_M1000_g 0.0170236f $X=8.255 $Y=1.685
+ $X2=0 $Y2=0
cc_525 N_A_795_74#_c_613_n N_A_991_81#_M1000_g 9.68097e-19 $X=8.425 $Y=1.685
+ $X2=0 $Y2=0
cc_526 N_A_795_74#_c_637_n N_A_991_81#_M1007_g 0.0047106f $X=8.255 $Y=1.685
+ $X2=0 $Y2=0
cc_527 N_A_795_74#_c_613_n N_A_991_81#_M1007_g 0.0139563f $X=8.425 $Y=1.685
+ $X2=0 $Y2=0
cc_528 N_A_795_74#_M1034_g N_A_991_81#_c_991_n 8.08997e-19 $X=4.975 $Y=2.495
+ $X2=0 $Y2=0
cc_529 N_A_795_74#_c_626_n N_A_991_81#_c_991_n 0.0194049f $X=5.645 $Y=2.895
+ $X2=0 $Y2=0
cc_530 N_A_795_74#_c_622_n N_A_991_81#_c_992_n 0.0191167f $X=5.56 $Y=2.98 $X2=0
+ $Y2=0
cc_531 N_A_795_74#_c_597_n N_A_991_81#_c_978_n 0.00423998f $X=5.625 $Y=1.35
+ $X2=0 $Y2=0
cc_532 N_A_795_74#_M1031_g N_A_991_81#_c_978_n 0.0209349f $X=5.64 $Y=0.615 $X2=0
+ $Y2=0
cc_533 N_A_795_74#_c_606_n N_A_991_81#_c_978_n 0.00340526f $X=5 $Y=0.34 $X2=0
+ $Y2=0
cc_534 N_A_795_74#_c_608_n N_A_991_81#_c_978_n 0.00865059f $X=4.875 $Y=1.565
+ $X2=0 $Y2=0
cc_535 N_A_795_74#_c_609_n N_A_991_81#_c_978_n 0.0446184f $X=5.085 $Y=1.015
+ $X2=0 $Y2=0
cc_536 N_A_795_74#_c_612_n N_A_991_81#_c_978_n 0.0139975f $X=5.085 $Y=1.1 $X2=0
+ $Y2=0
cc_537 N_A_795_74#_c_616_n N_A_991_81#_c_978_n 0.0010998f $X=5.565 $Y=1.58 $X2=0
+ $Y2=0
cc_538 N_A_795_74#_c_627_n N_A_991_81#_c_979_n 0.00708192f $X=6.515 $Y=2.17
+ $X2=0 $Y2=0
cc_539 N_A_795_74#_c_615_n N_A_991_81#_c_979_n 4.23483e-19 $X=5.565 $Y=1.655
+ $X2=0 $Y2=0
cc_540 N_A_795_74#_c_616_n N_A_991_81#_c_979_n 0.011013f $X=5.565 $Y=1.58 $X2=0
+ $Y2=0
cc_541 N_A_795_74#_c_596_n N_A_991_81#_c_980_n 0.0114893f $X=5.4 $Y=1.655 $X2=0
+ $Y2=0
cc_542 N_A_795_74#_c_608_n N_A_991_81#_c_980_n 0.0138133f $X=4.875 $Y=1.565
+ $X2=0 $Y2=0
cc_543 N_A_795_74#_c_625_n N_A_991_81#_c_980_n 0.0192633f $X=5.645 $Y=2.255
+ $X2=0 $Y2=0
cc_544 N_A_795_74#_c_612_n N_A_991_81#_c_980_n 0.00243713f $X=5.085 $Y=1.1 $X2=0
+ $Y2=0
cc_545 N_A_795_74#_c_614_n N_A_991_81#_c_980_n 0.00165075f $X=5.065 $Y=1.565
+ $X2=0 $Y2=0
cc_546 N_A_795_74#_c_616_n N_A_991_81#_c_980_n 0.00452136f $X=5.565 $Y=1.58
+ $X2=0 $Y2=0
cc_547 N_A_795_74#_M1034_g N_A_991_81#_c_984_n 0.00836786f $X=4.975 $Y=2.495
+ $X2=0 $Y2=0
cc_548 N_A_795_74#_c_596_n N_A_991_81#_c_984_n 0.0132701f $X=5.4 $Y=1.655 $X2=0
+ $Y2=0
cc_549 N_A_795_74#_c_608_n N_A_991_81#_c_984_n 0.0128533f $X=4.875 $Y=1.565
+ $X2=0 $Y2=0
cc_550 N_A_795_74#_c_625_n N_A_991_81#_c_984_n 0.0374763f $X=5.645 $Y=2.255
+ $X2=0 $Y2=0
cc_551 N_A_795_74#_c_626_n N_A_991_81#_c_984_n 5.11006e-19 $X=5.645 $Y=2.895
+ $X2=0 $Y2=0
cc_552 N_A_795_74#_c_614_n N_A_991_81#_c_984_n 3.64028e-19 $X=5.065 $Y=1.565
+ $X2=0 $Y2=0
cc_553 N_A_795_74#_c_615_n N_A_991_81#_c_984_n 0.00251116f $X=5.565 $Y=1.655
+ $X2=0 $Y2=0
cc_554 N_A_795_74#_c_616_n N_A_991_81#_c_984_n 7.34463e-19 $X=5.565 $Y=1.58
+ $X2=0 $Y2=0
cc_555 N_A_795_74#_c_637_n N_A_991_81#_c_985_n 0.0235309f $X=8.255 $Y=1.685
+ $X2=0 $Y2=0
cc_556 N_A_795_74#_c_613_n N_A_991_81#_c_985_n 0.00630615f $X=8.425 $Y=1.685
+ $X2=0 $Y2=0
cc_557 N_A_795_74#_c_600_n N_A_991_81#_c_987_n 0.00756279f $X=9.14 $Y=1.16 $X2=0
+ $Y2=0
cc_558 N_A_795_74#_c_611_n N_A_991_81#_c_987_n 0.0083803f $X=8.975 $Y=1.64 $X2=0
+ $Y2=0
cc_559 N_A_795_74#_c_637_n N_A_991_81#_c_987_n 0.00169988f $X=8.255 $Y=1.685
+ $X2=0 $Y2=0
cc_560 N_A_795_74#_c_613_n N_A_991_81#_c_987_n 0.0106947f $X=8.425 $Y=1.685
+ $X2=0 $Y2=0
cc_561 N_A_795_74#_c_617_n N_A_991_81#_c_987_n 0.00558876f $X=8.975 $Y=1.475
+ $X2=0 $Y2=0
cc_562 N_A_795_74#_c_628_n N_SET_B_M1021_g 5.29289e-19 $X=6.6 $Y=2.905 $X2=0
+ $Y2=0
cc_563 N_A_795_74#_c_629_n N_SET_B_M1021_g 0.00183892f $X=7.195 $Y=2.99 $X2=0
+ $Y2=0
cc_564 N_A_795_74#_c_631_n N_SET_B_M1021_g 0.0260089f $X=7.28 $Y=2.905 $X2=0
+ $Y2=0
cc_565 N_A_795_74#_c_632_n N_SET_B_M1021_g 0.00772828f $X=7.365 $Y=1.81 $X2=0
+ $Y2=0
cc_566 N_A_795_74#_c_599_n N_SET_B_c_1155_n 0.00630186f $X=9.625 $Y=1.16 $X2=0
+ $Y2=0
cc_567 N_A_795_74#_c_600_n N_SET_B_c_1155_n 0.00131559f $X=9.14 $Y=1.16 $X2=0
+ $Y2=0
cc_568 N_A_795_74#_c_602_n N_SET_B_c_1155_n 0.00829517f $X=10.055 $Y=1.16 $X2=0
+ $Y2=0
cc_569 N_A_795_74#_c_604_n N_SET_B_c_1155_n 0.00149277f $X=9.7 $Y=1.16 $X2=0
+ $Y2=0
cc_570 N_A_795_74#_c_610_n N_SET_B_c_1155_n 0.00715649f $X=10 $Y=1.64 $X2=0
+ $Y2=0
cc_571 N_A_795_74#_c_611_n N_SET_B_c_1155_n 0.0045015f $X=8.975 $Y=1.64 $X2=0
+ $Y2=0
cc_572 N_A_795_74#_c_635_n N_SET_B_c_1155_n 0.0100687f $X=10.555 $Y=1.97 $X2=0
+ $Y2=0
cc_573 N_A_795_74#_c_637_n N_SET_B_c_1155_n 0.012825f $X=8.255 $Y=1.685 $X2=0
+ $Y2=0
cc_574 N_A_795_74#_c_613_n N_SET_B_c_1155_n 0.0535919f $X=8.425 $Y=1.685 $X2=0
+ $Y2=0
cc_575 N_A_795_74#_c_617_n N_SET_B_c_1155_n 0.0054977f $X=8.975 $Y=1.475 $X2=0
+ $Y2=0
cc_576 N_A_795_74#_c_632_n N_SET_B_c_1156_n 4.20079e-19 $X=7.365 $Y=1.81 $X2=0
+ $Y2=0
cc_577 N_A_795_74#_c_637_n N_SET_B_c_1156_n 0.0022884f $X=8.255 $Y=1.685 $X2=0
+ $Y2=0
cc_578 N_A_795_74#_c_632_n N_SET_B_c_1157_n 0.0126733f $X=7.365 $Y=1.81 $X2=0
+ $Y2=0
cc_579 N_A_795_74#_c_637_n N_SET_B_c_1157_n 0.0134421f $X=8.255 $Y=1.685 $X2=0
+ $Y2=0
cc_580 N_A_795_74#_c_632_n N_SET_B_c_1159_n 5.14458e-19 $X=7.365 $Y=1.81 $X2=0
+ $Y2=0
cc_581 N_A_795_74#_c_637_n N_SET_B_c_1159_n 0.00118211f $X=8.255 $Y=1.685 $X2=0
+ $Y2=0
cc_582 N_A_795_74#_c_605_n N_A_608_74#_M1006_g 0.00163108f $X=4.115 $Y=0.515
+ $X2=0 $Y2=0
cc_583 N_A_795_74#_c_607_n N_A_608_74#_M1006_g 0.00266901f $X=4.2 $Y=0.34 $X2=0
+ $Y2=0
cc_584 N_A_795_74#_c_623_n N_A_608_74#_M1040_g 0.00104356f $X=4.325 $Y=2.98
+ $X2=0 $Y2=0
cc_585 N_A_795_74#_c_608_n N_A_608_74#_c_1285_n 0.00118998f $X=4.875 $Y=1.565
+ $X2=0 $Y2=0
cc_586 N_A_795_74#_c_621_n N_A_608_74#_c_1299_n 0.00590439f $X=4.16 $Y=2.78
+ $X2=0 $Y2=0
cc_587 N_A_795_74#_c_622_n N_A_608_74#_c_1299_n 0.0134696f $X=5.56 $Y=2.98 $X2=0
+ $Y2=0
cc_588 N_A_795_74#_c_608_n N_A_608_74#_c_1286_n 0.0025543f $X=4.875 $Y=1.565
+ $X2=0 $Y2=0
cc_589 N_A_795_74#_c_612_n N_A_608_74#_c_1286_n 0.007948f $X=5.085 $Y=1.1 $X2=0
+ $Y2=0
cc_590 N_A_795_74#_c_614_n N_A_608_74#_c_1286_n 0.0160256f $X=5.065 $Y=1.565
+ $X2=0 $Y2=0
cc_591 N_A_795_74#_c_605_n N_A_608_74#_c_1287_n 8.15047e-19 $X=4.115 $Y=0.515
+ $X2=0 $Y2=0
cc_592 N_A_795_74#_c_606_n N_A_608_74#_c_1287_n 0.00184816f $X=5 $Y=0.34 $X2=0
+ $Y2=0
cc_593 N_A_795_74#_M1034_g N_A_608_74#_c_1300_n 0.0088468f $X=4.975 $Y=2.495
+ $X2=0 $Y2=0
cc_594 N_A_795_74#_c_622_n N_A_608_74#_c_1300_n 0.0136847f $X=5.56 $Y=2.98 $X2=0
+ $Y2=0
cc_595 N_A_795_74#_M1031_g N_A_608_74#_M1024_g 0.00858665f $X=5.64 $Y=0.615
+ $X2=0 $Y2=0
cc_596 N_A_795_74#_c_605_n N_A_608_74#_M1024_g 0.00311369f $X=4.115 $Y=0.515
+ $X2=0 $Y2=0
cc_597 N_A_795_74#_c_606_n N_A_608_74#_M1024_g 0.0136298f $X=5 $Y=0.34 $X2=0
+ $Y2=0
cc_598 N_A_795_74#_c_609_n N_A_608_74#_M1024_g 0.00592452f $X=5.085 $Y=1.015
+ $X2=0 $Y2=0
cc_599 N_A_795_74#_c_612_n N_A_608_74#_M1024_g 0.00464804f $X=5.085 $Y=1.1 $X2=0
+ $Y2=0
cc_600 N_A_795_74#_M1034_g N_A_608_74#_M1018_g 0.0102622f $X=4.975 $Y=2.495
+ $X2=0 $Y2=0
cc_601 N_A_795_74#_c_622_n N_A_608_74#_M1018_g 0.0173074f $X=5.56 $Y=2.98 $X2=0
+ $Y2=0
cc_602 N_A_795_74#_c_625_n N_A_608_74#_M1018_g 6.45027e-19 $X=5.645 $Y=2.255
+ $X2=0 $Y2=0
cc_603 N_A_795_74#_c_626_n N_A_608_74#_M1018_g 0.0159101f $X=5.645 $Y=2.895
+ $X2=0 $Y2=0
cc_604 N_A_795_74#_c_615_n N_A_608_74#_M1018_g 0.010993f $X=5.565 $Y=1.655 $X2=0
+ $Y2=0
cc_605 N_A_795_74#_c_622_n N_A_608_74#_c_1303_n 9.85337e-19 $X=5.56 $Y=2.98
+ $X2=0 $Y2=0
cc_606 N_A_795_74#_c_629_n N_A_608_74#_c_1303_n 0.0111624f $X=7.195 $Y=2.99
+ $X2=0 $Y2=0
cc_607 N_A_795_74#_c_630_n N_A_608_74#_c_1303_n 0.00320029f $X=6.685 $Y=2.99
+ $X2=0 $Y2=0
cc_608 N_A_795_74#_c_610_n N_A_608_74#_M1003_g 0.0153479f $X=10 $Y=1.64 $X2=0
+ $Y2=0
cc_609 N_A_795_74#_c_611_n N_A_608_74#_M1003_g 0.0118206f $X=8.975 $Y=1.64 $X2=0
+ $Y2=0
cc_610 N_A_795_74#_c_604_n N_A_608_74#_c_1290_n 0.0283403f $X=9.7 $Y=1.16 $X2=0
+ $Y2=0
cc_611 N_A_795_74#_c_610_n N_A_608_74#_c_1290_n 0.0272908f $X=10 $Y=1.64 $X2=0
+ $Y2=0
cc_612 N_A_795_74#_c_635_n N_A_608_74#_c_1290_n 0.00901037f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_613 N_A_795_74#_c_636_n N_A_608_74#_c_1290_n 0.0200004f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_614 N_A_795_74#_c_599_n N_A_608_74#_c_1291_n 0.0283403f $X=9.625 $Y=1.16
+ $X2=0 $Y2=0
cc_615 N_A_795_74#_c_610_n N_A_608_74#_c_1291_n 0.0048077f $X=10 $Y=1.64 $X2=0
+ $Y2=0
cc_616 N_A_795_74#_c_617_n N_A_608_74#_c_1291_n 0.0118206f $X=8.975 $Y=1.475
+ $X2=0 $Y2=0
cc_617 N_A_795_74#_M1019_g N_A_608_74#_c_1306_n 0.0152486f $X=10.63 $Y=2.75
+ $X2=0 $Y2=0
cc_618 N_A_795_74#_c_610_n N_A_608_74#_c_1306_n 0.00536301f $X=10 $Y=1.64 $X2=0
+ $Y2=0
cc_619 N_A_795_74#_c_636_n N_A_608_74#_c_1306_n 0.00341743f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_620 N_A_795_74#_c_603_n N_A_608_74#_M1044_g 0.024414f $X=10.13 $Y=1.085 $X2=0
+ $Y2=0
cc_621 N_A_795_74#_M1034_g N_A_608_74#_c_1307_n 0.00663995f $X=4.975 $Y=2.495
+ $X2=0 $Y2=0
cc_622 N_A_795_74#_M1034_g N_A_608_74#_c_1308_n 0.0204879f $X=4.975 $Y=2.495
+ $X2=0 $Y2=0
cc_623 N_A_795_74#_M1040_d N_A_608_74#_c_1312_n 0.00370981f $X=4.025 $Y=1.84
+ $X2=0 $Y2=0
cc_624 N_A_795_74#_c_605_n N_A_608_74#_c_1295_n 0.012379f $X=4.115 $Y=0.515
+ $X2=0 $Y2=0
cc_625 N_A_795_74#_c_605_n N_A_608_74#_c_1297_n 0.00102327f $X=4.115 $Y=0.515
+ $X2=0 $Y2=0
cc_626 N_A_795_74#_c_608_n N_A_608_74#_c_1297_n 3.17258e-19 $X=4.875 $Y=1.565
+ $X2=0 $Y2=0
cc_627 N_A_795_74#_c_614_n N_A_608_74#_c_1297_n 0.021129f $X=5.065 $Y=1.565
+ $X2=0 $Y2=0
cc_628 N_A_795_74#_c_636_n N_A_2186_367#_c_1490_n 0.0391129f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_629 N_A_795_74#_M1019_g N_A_2186_367#_M1008_g 0.0391129f $X=10.63 $Y=2.75
+ $X2=0 $Y2=0
cc_630 N_A_795_74#_c_636_n N_A_2186_367#_c_1482_n 0.00162157f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_631 N_A_795_74#_c_610_n N_A_1804_424#_M1010_s 0.00390815f $X=10 $Y=1.64 $X2=0
+ $Y2=0
cc_632 N_A_795_74#_c_635_n N_A_1804_424#_M1010_s 7.16004e-19 $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_633 N_A_795_74#_M1019_g N_A_1804_424#_c_1604_n 0.00305757f $X=10.63 $Y=2.75
+ $X2=0 $Y2=0
cc_634 N_A_795_74#_c_601_n N_A_1804_424#_c_1591_n 0.0109156f $X=9.7 $Y=1.085
+ $X2=0 $Y2=0
cc_635 N_A_795_74#_c_603_n N_A_1804_424#_c_1591_n 0.0133206f $X=10.13 $Y=1.085
+ $X2=0 $Y2=0
cc_636 N_A_795_74#_M1019_g N_A_1804_424#_c_1606_n 0.00906653f $X=10.63 $Y=2.75
+ $X2=0 $Y2=0
cc_637 N_A_795_74#_c_603_n N_A_1804_424#_c_1592_n 0.00571513f $X=10.13 $Y=1.085
+ $X2=0 $Y2=0
cc_638 N_A_795_74#_c_610_n N_A_1804_424#_c_1607_n 0.00575761f $X=10 $Y=1.64
+ $X2=0 $Y2=0
cc_639 N_A_795_74#_c_635_n N_A_1804_424#_c_1607_n 0.0230587f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_640 N_A_795_74#_c_636_n N_A_1804_424#_c_1607_n 0.0010483f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_641 N_A_795_74#_c_635_n N_A_1804_424#_c_1593_n 0.00705752f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_642 N_A_795_74#_c_636_n N_A_1804_424#_c_1593_n 8.63221e-19 $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_643 N_A_795_74#_c_610_n N_A_1804_424#_c_1594_n 0.00546536f $X=10 $Y=1.64
+ $X2=0 $Y2=0
cc_644 N_A_795_74#_c_635_n N_A_1804_424#_c_1594_n 0.00959246f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_645 N_A_795_74#_c_636_n N_A_1804_424#_c_1594_n 5.89689e-19 $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_646 N_A_795_74#_c_635_n N_A_1804_424#_c_1595_n 0.0128867f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_647 N_A_795_74#_c_636_n N_A_1804_424#_c_1595_n 4.82162e-19 $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_648 N_A_795_74#_c_601_n N_A_1804_424#_c_1598_n 0.00165289f $X=9.7 $Y=1.085
+ $X2=0 $Y2=0
cc_649 N_A_795_74#_M1019_g N_A_1804_424#_c_1612_n 0.013918f $X=10.63 $Y=2.75
+ $X2=0 $Y2=0
cc_650 N_A_795_74#_c_635_n N_A_1804_424#_c_1612_n 0.0207081f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_651 N_A_795_74#_c_636_n N_A_1804_424#_c_1612_n 0.00235196f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_652 N_A_795_74#_c_635_n N_A_1804_424#_c_1613_n 0.014313f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_653 N_A_795_74#_c_636_n N_A_1804_424#_c_1613_n 0.00520943f $X=10.555 $Y=1.97
+ $X2=0 $Y2=0
cc_654 N_A_795_74#_c_628_n N_VPWR_M1042_d 0.00437233f $X=6.6 $Y=2.905 $X2=0
+ $Y2=0
cc_655 N_A_795_74#_c_631_n N_VPWR_M1021_d 0.00382783f $X=7.28 $Y=2.905 $X2=0
+ $Y2=0
cc_656 N_A_795_74#_c_623_n N_VPWR_c_1859_n 0.00994466f $X=4.325 $Y=2.98 $X2=0
+ $Y2=0
cc_657 N_A_795_74#_c_622_n N_VPWR_c_1860_n 0.00867486f $X=5.56 $Y=2.98 $X2=0
+ $Y2=0
cc_658 N_A_795_74#_c_626_n N_VPWR_c_1860_n 0.0190638f $X=5.645 $Y=2.895 $X2=0
+ $Y2=0
cc_659 N_A_795_74#_c_627_n N_VPWR_c_1860_n 0.0177503f $X=6.515 $Y=2.17 $X2=0
+ $Y2=0
cc_660 N_A_795_74#_c_628_n N_VPWR_c_1860_n 0.0363339f $X=6.6 $Y=2.905 $X2=0
+ $Y2=0
cc_661 N_A_795_74#_c_630_n N_VPWR_c_1860_n 0.0147459f $X=6.685 $Y=2.99 $X2=0
+ $Y2=0
cc_662 N_A_795_74#_c_629_n N_VPWR_c_1861_n 0.0143583f $X=7.195 $Y=2.99 $X2=0
+ $Y2=0
cc_663 N_A_795_74#_c_631_n N_VPWR_c_1861_n 0.0617585f $X=7.28 $Y=2.905 $X2=0
+ $Y2=0
cc_664 N_A_795_74#_c_637_n N_VPWR_c_1861_n 0.0136226f $X=8.255 $Y=1.685 $X2=0
+ $Y2=0
cc_665 N_A_795_74#_M1019_g N_VPWR_c_1863_n 0.00134211f $X=10.63 $Y=2.75 $X2=0
+ $Y2=0
cc_666 N_A_795_74#_c_622_n N_VPWR_c_1868_n 0.085277f $X=5.56 $Y=2.98 $X2=0 $Y2=0
cc_667 N_A_795_74#_c_623_n N_VPWR_c_1868_n 0.0164393f $X=4.325 $Y=2.98 $X2=0
+ $Y2=0
cc_668 N_A_795_74#_c_629_n N_VPWR_c_1870_n 0.0443733f $X=7.195 $Y=2.99 $X2=0
+ $Y2=0
cc_669 N_A_795_74#_c_630_n N_VPWR_c_1870_n 0.0115893f $X=6.685 $Y=2.99 $X2=0
+ $Y2=0
cc_670 N_A_795_74#_M1019_g N_VPWR_c_1876_n 0.00553757f $X=10.63 $Y=2.75 $X2=0
+ $Y2=0
cc_671 N_A_795_74#_M1019_g N_VPWR_c_1855_n 0.00562325f $X=10.63 $Y=2.75 $X2=0
+ $Y2=0
cc_672 N_A_795_74#_c_622_n N_VPWR_c_1855_n 0.0470528f $X=5.56 $Y=2.98 $X2=0
+ $Y2=0
cc_673 N_A_795_74#_c_623_n N_VPWR_c_1855_n 0.00958732f $X=4.325 $Y=2.98 $X2=0
+ $Y2=0
cc_674 N_A_795_74#_c_629_n N_VPWR_c_1855_n 0.0229659f $X=7.195 $Y=2.99 $X2=0
+ $Y2=0
cc_675 N_A_795_74#_c_630_n N_VPWR_c_1855_n 0.00583135f $X=6.685 $Y=2.99 $X2=0
+ $Y2=0
cc_676 N_A_795_74#_c_606_n N_A_293_464#_M1024_s 0.00228614f $X=5 $Y=0.34 $X2=0
+ $Y2=0
cc_677 N_A_795_74#_M1040_d N_A_293_464#_c_2046_n 0.00465691f $X=4.025 $Y=1.84
+ $X2=0 $Y2=0
cc_678 N_A_795_74#_c_621_n N_A_293_464#_c_2046_n 0.019304f $X=4.16 $Y=2.78 $X2=0
+ $Y2=0
cc_679 N_A_795_74#_c_622_n N_A_293_464#_c_2046_n 0.00832577f $X=5.56 $Y=2.98
+ $X2=0 $Y2=0
cc_680 N_A_795_74#_M1034_g N_A_293_464#_c_2047_n 0.00422767f $X=4.975 $Y=2.495
+ $X2=0 $Y2=0
cc_681 N_A_795_74#_c_605_n N_A_293_464#_c_2042_n 0.0164119f $X=4.115 $Y=0.515
+ $X2=0 $Y2=0
cc_682 N_A_795_74#_c_606_n N_A_293_464#_c_2042_n 0.0249256f $X=5 $Y=0.34 $X2=0
+ $Y2=0
cc_683 N_A_795_74#_c_609_n N_A_293_464#_c_2042_n 0.0103527f $X=5.085 $Y=1.015
+ $X2=0 $Y2=0
cc_684 N_A_795_74#_c_612_n N_A_293_464#_c_2042_n 0.0052363f $X=5.085 $Y=1.1
+ $X2=0 $Y2=0
cc_685 N_A_795_74#_M1034_g N_A_293_464#_c_2043_n 0.00143241f $X=4.975 $Y=2.495
+ $X2=0 $Y2=0
cc_686 N_A_795_74#_c_605_n N_A_293_464#_c_2043_n 0.0171937f $X=4.115 $Y=0.515
+ $X2=0 $Y2=0
cc_687 N_A_795_74#_c_608_n N_A_293_464#_c_2043_n 0.0403116f $X=4.875 $Y=1.565
+ $X2=0 $Y2=0
cc_688 N_A_795_74#_c_609_n N_A_293_464#_c_2043_n 0.00693452f $X=5.085 $Y=1.015
+ $X2=0 $Y2=0
cc_689 N_A_795_74#_c_612_n N_A_293_464#_c_2043_n 0.0124645f $X=5.085 $Y=1.1
+ $X2=0 $Y2=0
cc_690 N_A_795_74#_c_614_n N_A_293_464#_c_2043_n 0.00203394f $X=5.065 $Y=1.565
+ $X2=0 $Y2=0
cc_691 N_A_795_74#_M1034_g N_A_293_464#_c_2050_n 0.00502684f $X=4.975 $Y=2.495
+ $X2=0 $Y2=0
cc_692 N_A_795_74#_c_608_n N_A_293_464#_c_2050_n 0.0132956f $X=4.875 $Y=1.565
+ $X2=0 $Y2=0
cc_693 N_A_795_74#_c_614_n N_A_293_464#_c_2050_n 0.00324793f $X=5.065 $Y=1.565
+ $X2=0 $Y2=0
cc_694 N_A_795_74#_M1034_g N_A_293_464#_c_2051_n 0.00722315f $X=4.975 $Y=2.495
+ $X2=0 $Y2=0
cc_695 N_A_795_74#_c_621_n N_A_293_464#_c_2051_n 0.00878202f $X=4.16 $Y=2.78
+ $X2=0 $Y2=0
cc_696 N_A_795_74#_c_622_n N_A_293_464#_c_2051_n 0.0258523f $X=5.56 $Y=2.98
+ $X2=0 $Y2=0
cc_697 N_A_795_74#_c_626_n A_1120_483# 0.00609261f $X=5.645 $Y=2.895 $X2=-0.19
+ $Y2=-0.245
cc_698 N_A_795_74#_c_610_n N_A_1587_379#_c_2177_n 0.00929881f $X=10 $Y=1.64
+ $X2=0 $Y2=0
cc_699 N_A_795_74#_c_637_n N_A_1587_379#_c_2177_n 0.012482f $X=8.255 $Y=1.685
+ $X2=0 $Y2=0
cc_700 N_A_795_74#_c_610_n N_A_1587_379#_c_2174_n 0.0948996f $X=10 $Y=1.64 $X2=0
+ $Y2=0
cc_701 N_A_795_74#_c_611_n N_A_1587_379#_c_2174_n 0.00798977f $X=8.975 $Y=1.64
+ $X2=0 $Y2=0
cc_702 N_A_795_74#_c_637_n N_A_1587_379#_c_2175_n 0.0217164f $X=8.255 $Y=1.685
+ $X2=0 $Y2=0
cc_703 N_A_795_74#_c_610_n N_A_1587_379#_c_2176_n 0.0134175f $X=10 $Y=1.64 $X2=0
+ $Y2=0
cc_704 N_A_795_74#_c_607_n N_VGND_c_2252_n 0.0112234f $X=4.2 $Y=0.34 $X2=0 $Y2=0
cc_705 N_A_795_74#_c_601_n N_VGND_c_2254_n 3.14208e-19 $X=9.7 $Y=1.085 $X2=0
+ $Y2=0
cc_706 N_A_795_74#_M1031_g N_VGND_c_2259_n 0.00527282f $X=5.64 $Y=0.615 $X2=0
+ $Y2=0
cc_707 N_A_795_74#_c_606_n N_VGND_c_2259_n 0.0636631f $X=5 $Y=0.34 $X2=0 $Y2=0
cc_708 N_A_795_74#_c_607_n N_VGND_c_2259_n 0.0121867f $X=4.2 $Y=0.34 $X2=0 $Y2=0
cc_709 N_A_795_74#_c_601_n N_VGND_c_2271_n 0.00278271f $X=9.7 $Y=1.085 $X2=0
+ $Y2=0
cc_710 N_A_795_74#_c_603_n N_VGND_c_2271_n 0.00278271f $X=10.13 $Y=1.085 $X2=0
+ $Y2=0
cc_711 N_A_795_74#_M1031_g N_VGND_c_2274_n 0.00534666f $X=5.64 $Y=0.615 $X2=0
+ $Y2=0
cc_712 N_A_795_74#_c_601_n N_VGND_c_2274_n 0.00358427f $X=9.7 $Y=1.085 $X2=0
+ $Y2=0
cc_713 N_A_795_74#_c_603_n N_VGND_c_2274_n 0.0035414f $X=10.13 $Y=1.085 $X2=0
+ $Y2=0
cc_714 N_A_795_74#_c_606_n N_VGND_c_2274_n 0.0366794f $X=5 $Y=0.34 $X2=0 $Y2=0
cc_715 N_A_795_74#_c_607_n N_VGND_c_2274_n 0.00660921f $X=4.2 $Y=0.34 $X2=0
+ $Y2=0
cc_716 N_A_795_74#_c_600_n N_A_1641_74#_c_2412_n 0.0178304f $X=9.14 $Y=1.16
+ $X2=0 $Y2=0
cc_717 N_A_795_74#_c_601_n N_A_1641_74#_c_2412_n 0.0116182f $X=9.7 $Y=1.085
+ $X2=0 $Y2=0
cc_718 N_A_795_74#_c_610_n N_A_1641_74#_c_2412_n 0.0233474f $X=10 $Y=1.64 $X2=0
+ $Y2=0
cc_719 N_A_795_74#_c_611_n N_A_1641_74#_c_2412_n 0.00335664f $X=8.975 $Y=1.64
+ $X2=0 $Y2=0
cc_720 N_A_795_74#_c_637_n N_A_1641_74#_c_2413_n 8.07173e-19 $X=8.255 $Y=1.685
+ $X2=0 $Y2=0
cc_721 N_A_795_74#_c_613_n N_A_1641_74#_c_2413_n 0.00555546f $X=8.425 $Y=1.685
+ $X2=0 $Y2=0
cc_722 N_A_795_74#_c_601_n N_A_1641_74#_c_2414_n 0.0110826f $X=9.7 $Y=1.085
+ $X2=0 $Y2=0
cc_723 N_A_795_74#_c_602_n N_A_1641_74#_c_2414_n 0.0027829f $X=10.055 $Y=1.16
+ $X2=0 $Y2=0
cc_724 N_A_795_74#_c_603_n N_A_1641_74#_c_2414_n 0.00708563f $X=10.13 $Y=1.085
+ $X2=0 $Y2=0
cc_725 N_A_795_74#_c_610_n N_A_1641_74#_c_2414_n 0.00654828f $X=10 $Y=1.64 $X2=0
+ $Y2=0
cc_726 N_A_1185_55#_c_882_n N_A_991_81#_c_970_n 0.00105699f $X=6.855 $Y=1.83
+ $X2=0 $Y2=0
cc_727 N_A_1185_55#_M1042_g N_A_991_81#_M1011_g 0.0146605f $X=6.03 $Y=2.525
+ $X2=0 $Y2=0
cc_728 N_A_1185_55#_c_882_n N_A_991_81#_M1011_g 0.0154789f $X=6.855 $Y=1.83
+ $X2=0 $Y2=0
cc_729 N_A_1185_55#_c_883_n N_A_991_81#_M1011_g 0.00609362f $X=6.94 $Y=2.515
+ $X2=0 $Y2=0
cc_730 N_A_1185_55#_c_878_n N_A_991_81#_M1011_g 0.0120011f $X=6.105 $Y=1.815
+ $X2=0 $Y2=0
cc_731 N_A_1185_55#_c_880_n N_A_991_81#_M1011_g 0.00242176f $X=6.105 $Y=1.65
+ $X2=0 $Y2=0
cc_732 N_A_1185_55#_c_876_n N_A_991_81#_c_972_n 0.00338254f $X=6.145 $Y=1.1
+ $X2=0 $Y2=0
cc_733 N_A_1185_55#_c_879_n N_A_991_81#_c_972_n 0.00677096f $X=6.855 $Y=0.525
+ $X2=0 $Y2=0
cc_734 N_A_1185_55#_c_874_n N_A_991_81#_c_977_n 0.00146983f $X=6 $Y=0.935 $X2=0
+ $Y2=0
cc_735 N_A_1185_55#_c_875_n N_A_991_81#_c_977_n 0.0177504f $X=6.055 $Y=1.265
+ $X2=0 $Y2=0
cc_736 N_A_1185_55#_c_876_n N_A_991_81#_c_977_n 5.30688e-19 $X=6.145 $Y=1.1
+ $X2=0 $Y2=0
cc_737 N_A_1185_55#_c_877_n N_A_991_81#_c_977_n 0.00370147f $X=6.69 $Y=0.615
+ $X2=0 $Y2=0
cc_738 N_A_1185_55#_c_879_n N_A_991_81#_c_977_n 0.00718643f $X=6.855 $Y=0.525
+ $X2=0 $Y2=0
cc_739 N_A_1185_55#_c_874_n N_A_991_81#_c_978_n 0.00224758f $X=6 $Y=0.935 $X2=0
+ $Y2=0
cc_740 N_A_1185_55#_c_875_n N_A_991_81#_c_978_n 0.00123351f $X=6.055 $Y=1.265
+ $X2=0 $Y2=0
cc_741 N_A_1185_55#_c_876_n N_A_991_81#_c_978_n 0.0189782f $X=6.145 $Y=1.1 $X2=0
+ $Y2=0
cc_742 N_A_1185_55#_c_896_n N_A_991_81#_c_978_n 0.00682346f $X=6.31 $Y=0.615
+ $X2=0 $Y2=0
cc_743 N_A_1185_55#_c_875_n N_A_991_81#_c_979_n 0.00359104f $X=6.055 $Y=1.265
+ $X2=0 $Y2=0
cc_744 N_A_1185_55#_c_876_n N_A_991_81#_c_979_n 0.0256385f $X=6.145 $Y=1.1 $X2=0
+ $Y2=0
cc_745 N_A_1185_55#_c_882_n N_A_991_81#_c_979_n 0.0441129f $X=6.855 $Y=1.83
+ $X2=0 $Y2=0
cc_746 N_A_1185_55#_c_877_n N_A_991_81#_c_979_n 0.0066704f $X=6.69 $Y=0.615
+ $X2=0 $Y2=0
cc_747 N_A_1185_55#_c_878_n N_A_991_81#_c_979_n 0.00168199f $X=6.105 $Y=1.815
+ $X2=0 $Y2=0
cc_748 N_A_1185_55#_c_885_n N_A_991_81#_c_979_n 0.0233235f $X=6.27 $Y=1.815
+ $X2=0 $Y2=0
cc_749 N_A_1185_55#_c_880_n N_A_991_81#_c_979_n 0.0111257f $X=6.105 $Y=1.65
+ $X2=0 $Y2=0
cc_750 N_A_1185_55#_c_875_n N_A_991_81#_c_1064_n 0.00103048f $X=6.055 $Y=1.265
+ $X2=0 $Y2=0
cc_751 N_A_1185_55#_c_876_n N_A_991_81#_c_1064_n 0.00937167f $X=6.145 $Y=1.1
+ $X2=0 $Y2=0
cc_752 N_A_1185_55#_c_880_n N_A_991_81#_c_1064_n 6.17268e-19 $X=6.105 $Y=1.65
+ $X2=0 $Y2=0
cc_753 N_A_1185_55#_c_876_n N_A_991_81#_c_981_n 6.07444e-19 $X=6.145 $Y=1.1
+ $X2=0 $Y2=0
cc_754 N_A_1185_55#_c_880_n N_A_991_81#_c_981_n 0.00843579f $X=6.105 $Y=1.65
+ $X2=0 $Y2=0
cc_755 N_A_1185_55#_c_879_n N_A_991_81#_c_982_n 0.00793363f $X=6.855 $Y=0.525
+ $X2=0 $Y2=0
cc_756 N_A_1185_55#_c_875_n N_A_991_81#_c_983_n 3.96639e-19 $X=6.055 $Y=1.265
+ $X2=0 $Y2=0
cc_757 N_A_1185_55#_c_876_n N_A_991_81#_c_983_n 0.0105303f $X=6.145 $Y=1.1 $X2=0
+ $Y2=0
cc_758 N_A_1185_55#_c_877_n N_A_991_81#_c_983_n 0.0112142f $X=6.69 $Y=0.615
+ $X2=0 $Y2=0
cc_759 N_A_1185_55#_c_879_n N_A_991_81#_c_983_n 0.0157846f $X=6.855 $Y=0.525
+ $X2=0 $Y2=0
cc_760 N_A_1185_55#_M1042_g N_A_991_81#_c_984_n 6.36414e-19 $X=6.03 $Y=2.525
+ $X2=0 $Y2=0
cc_761 N_A_1185_55#_c_878_n N_A_991_81#_c_984_n 2.0933e-19 $X=6.105 $Y=1.815
+ $X2=0 $Y2=0
cc_762 N_A_1185_55#_c_880_n N_A_991_81#_c_984_n 2.07566e-19 $X=6.105 $Y=1.65
+ $X2=0 $Y2=0
cc_763 N_A_1185_55#_c_882_n N_SET_B_M1021_g 0.00136415f $X=6.855 $Y=1.83 $X2=0
+ $Y2=0
cc_764 N_A_1185_55#_c_883_n N_SET_B_M1021_g 0.00402039f $X=6.94 $Y=2.515 $X2=0
+ $Y2=0
cc_765 N_A_1185_55#_c_879_n N_SET_B_M1027_g 0.00103321f $X=6.855 $Y=0.525 $X2=0
+ $Y2=0
cc_766 N_A_1185_55#_M1042_g N_A_608_74#_M1018_g 0.018444f $X=6.03 $Y=2.525 $X2=0
+ $Y2=0
cc_767 N_A_1185_55#_M1042_g N_A_608_74#_c_1303_n 0.0123939f $X=6.03 $Y=2.525
+ $X2=0 $Y2=0
cc_768 N_A_1185_55#_M1042_g N_VPWR_c_1860_n 0.00903974f $X=6.03 $Y=2.525 $X2=0
+ $Y2=0
cc_769 N_A_1185_55#_M1042_g N_VPWR_c_1855_n 9.76808e-19 $X=6.03 $Y=2.525 $X2=0
+ $Y2=0
cc_770 N_A_1185_55#_c_876_n N_VGND_M1020_d 0.00256846f $X=6.145 $Y=1.1 $X2=0
+ $Y2=0
cc_771 N_A_1185_55#_c_877_n N_VGND_M1020_d 0.00518446f $X=6.69 $Y=0.615 $X2=0
+ $Y2=0
cc_772 N_A_1185_55#_c_896_n N_VGND_M1020_d 0.00235471f $X=6.31 $Y=0.615 $X2=0
+ $Y2=0
cc_773 N_A_1185_55#_c_879_n N_VGND_c_2253_n 0.0107976f $X=6.855 $Y=0.525 $X2=0
+ $Y2=0
cc_774 N_A_1185_55#_c_874_n N_VGND_c_2258_n 0.00357449f $X=6 $Y=0.935 $X2=0
+ $Y2=0
cc_775 N_A_1185_55#_c_875_n N_VGND_c_2258_n 5.89315e-19 $X=6.055 $Y=1.265 $X2=0
+ $Y2=0
cc_776 N_A_1185_55#_c_877_n N_VGND_c_2258_n 0.0109664f $X=6.69 $Y=0.615 $X2=0
+ $Y2=0
cc_777 N_A_1185_55#_c_896_n N_VGND_c_2258_n 0.0144987f $X=6.31 $Y=0.615 $X2=0
+ $Y2=0
cc_778 N_A_1185_55#_c_879_n N_VGND_c_2258_n 6.74191e-19 $X=6.855 $Y=0.525 $X2=0
+ $Y2=0
cc_779 N_A_1185_55#_c_874_n N_VGND_c_2259_n 0.00463637f $X=6 $Y=0.935 $X2=0
+ $Y2=0
cc_780 N_A_1185_55#_c_896_n N_VGND_c_2259_n 0.00291775f $X=6.31 $Y=0.615 $X2=0
+ $Y2=0
cc_781 N_A_1185_55#_c_877_n N_VGND_c_2262_n 0.00533357f $X=6.69 $Y=0.615 $X2=0
+ $Y2=0
cc_782 N_A_1185_55#_c_879_n N_VGND_c_2262_n 0.0138937f $X=6.855 $Y=0.525 $X2=0
+ $Y2=0
cc_783 N_A_1185_55#_c_874_n N_VGND_c_2274_n 0.00534666f $X=6 $Y=0.935 $X2=0
+ $Y2=0
cc_784 N_A_1185_55#_c_877_n N_VGND_c_2274_n 0.00799229f $X=6.69 $Y=0.615 $X2=0
+ $Y2=0
cc_785 N_A_1185_55#_c_896_n N_VGND_c_2274_n 0.00597722f $X=6.31 $Y=0.615 $X2=0
+ $Y2=0
cc_786 N_A_1185_55#_c_879_n N_VGND_c_2274_n 0.0117406f $X=6.855 $Y=0.525 $X2=0
+ $Y2=0
cc_787 N_A_991_81#_c_970_n N_SET_B_M1021_g 0.00926619f $X=6.715 $Y=1.57 $X2=0
+ $Y2=0
cc_788 N_A_991_81#_M1011_g N_SET_B_M1021_g 0.0316695f $X=6.715 $Y=2.525 $X2=0
+ $Y2=0
cc_789 N_A_991_81#_M1000_g N_SET_B_M1021_g 0.0230815f $X=7.845 $Y=2.315 $X2=0
+ $Y2=0
cc_790 N_A_991_81#_c_972_n N_SET_B_M1027_g 0.040881f $X=7.07 $Y=0.865 $X2=0
+ $Y2=0
cc_791 N_A_991_81#_c_974_n N_SET_B_M1027_g 0.0171965f $X=8.13 $Y=1.085 $X2=0
+ $Y2=0
cc_792 N_A_991_81#_c_1064_n N_SET_B_M1027_g 8.84629e-19 $X=6.715 $Y=1.065 $X2=0
+ $Y2=0
cc_793 N_A_991_81#_c_981_n N_SET_B_M1027_g 0.00513936f $X=6.715 $Y=1.065 $X2=0
+ $Y2=0
cc_794 N_A_991_81#_c_982_n N_SET_B_M1027_g 0.0146456f $X=7.755 $Y=0.955 $X2=0
+ $Y2=0
cc_795 N_A_991_81#_c_986_n N_SET_B_M1027_g 0.00367161f $X=7.92 $Y=1.225 $X2=0
+ $Y2=0
cc_796 N_A_991_81#_c_982_n N_SET_B_c_1155_n 0.00755992f $X=7.755 $Y=0.955 $X2=0
+ $Y2=0
cc_797 N_A_991_81#_c_985_n N_SET_B_c_1155_n 0.0202042f $X=7.92 $Y=1.39 $X2=0
+ $Y2=0
cc_798 N_A_991_81#_c_987_n N_SET_B_c_1155_n 0.0182561f $X=8.295 $Y=1.32 $X2=0
+ $Y2=0
cc_799 N_A_991_81#_c_979_n N_SET_B_c_1156_n 2.14175e-19 $X=6.55 $Y=1.46 $X2=0
+ $Y2=0
cc_800 N_A_991_81#_c_1064_n N_SET_B_c_1156_n 0.0020303f $X=6.715 $Y=1.065 $X2=0
+ $Y2=0
cc_801 N_A_991_81#_c_981_n N_SET_B_c_1156_n 4.38236e-19 $X=6.715 $Y=1.065 $X2=0
+ $Y2=0
cc_802 N_A_991_81#_c_982_n N_SET_B_c_1156_n 0.00823128f $X=7.755 $Y=0.955 $X2=0
+ $Y2=0
cc_803 N_A_991_81#_c_985_n N_SET_B_c_1156_n 0.00130449f $X=7.92 $Y=1.39 $X2=0
+ $Y2=0
cc_804 N_A_991_81#_c_986_n N_SET_B_c_1156_n 0.00189718f $X=7.92 $Y=1.225 $X2=0
+ $Y2=0
cc_805 N_A_991_81#_c_987_n N_SET_B_c_1156_n 7.09844e-19 $X=8.295 $Y=1.32 $X2=0
+ $Y2=0
cc_806 N_A_991_81#_c_979_n N_SET_B_c_1157_n 0.0082709f $X=6.55 $Y=1.46 $X2=0
+ $Y2=0
cc_807 N_A_991_81#_c_1064_n N_SET_B_c_1157_n 0.00638026f $X=6.715 $Y=1.065 $X2=0
+ $Y2=0
cc_808 N_A_991_81#_c_981_n N_SET_B_c_1157_n 8.13904e-19 $X=6.715 $Y=1.065 $X2=0
+ $Y2=0
cc_809 N_A_991_81#_c_982_n N_SET_B_c_1157_n 0.0233965f $X=7.755 $Y=0.955 $X2=0
+ $Y2=0
cc_810 N_A_991_81#_c_986_n N_SET_B_c_1157_n 0.0216481f $X=7.92 $Y=1.225 $X2=0
+ $Y2=0
cc_811 N_A_991_81#_c_987_n N_SET_B_c_1157_n 0.00178299f $X=8.295 $Y=1.32 $X2=0
+ $Y2=0
cc_812 N_A_991_81#_c_977_n N_SET_B_c_1159_n 0.00166756f $X=7.07 $Y=0.94 $X2=0
+ $Y2=0
cc_813 N_A_991_81#_c_979_n N_SET_B_c_1159_n 8.22009e-19 $X=6.55 $Y=1.46 $X2=0
+ $Y2=0
cc_814 N_A_991_81#_c_1064_n N_SET_B_c_1159_n 6.05847e-19 $X=6.715 $Y=1.065 $X2=0
+ $Y2=0
cc_815 N_A_991_81#_c_981_n N_SET_B_c_1159_n 0.00926619f $X=6.715 $Y=1.065 $X2=0
+ $Y2=0
cc_816 N_A_991_81#_c_982_n N_SET_B_c_1159_n 0.00420665f $X=7.755 $Y=0.955 $X2=0
+ $Y2=0
cc_817 N_A_991_81#_c_985_n N_SET_B_c_1159_n 4.93533e-19 $X=7.92 $Y=1.39 $X2=0
+ $Y2=0
cc_818 N_A_991_81#_c_987_n N_SET_B_c_1159_n 0.0209248f $X=8.295 $Y=1.32 $X2=0
+ $Y2=0
cc_819 N_A_991_81#_c_978_n N_A_608_74#_M1024_g 0.00148512f $X=5.425 $Y=0.615
+ $X2=0 $Y2=0
cc_820 N_A_991_81#_c_991_n N_A_608_74#_M1018_g 0.00281166f $X=5.24 $Y=2.39 $X2=0
+ $Y2=0
cc_821 N_A_991_81#_M1011_g N_A_608_74#_c_1303_n 0.0109545f $X=6.715 $Y=2.525
+ $X2=0 $Y2=0
cc_822 N_A_991_81#_M1000_g N_A_608_74#_c_1303_n 0.0123594f $X=7.845 $Y=2.315
+ $X2=0 $Y2=0
cc_823 N_A_991_81#_M1007_g N_A_608_74#_c_1303_n 0.0123594f $X=8.295 $Y=2.315
+ $X2=0 $Y2=0
cc_824 N_A_991_81#_M1007_g N_A_1804_424#_c_1603_n 0.00285805f $X=8.295 $Y=2.315
+ $X2=0 $Y2=0
cc_825 N_A_991_81#_M1011_g N_VPWR_c_1860_n 0.00133128f $X=6.715 $Y=2.525 $X2=0
+ $Y2=0
cc_826 N_A_991_81#_M1000_g N_VPWR_c_1861_n 0.00310597f $X=7.845 $Y=2.315 $X2=0
+ $Y2=0
cc_827 N_A_991_81#_M1007_g N_VPWR_c_1862_n 0.00505401f $X=8.295 $Y=2.315 $X2=0
+ $Y2=0
cc_828 N_A_991_81#_M1000_g N_VPWR_c_1855_n 0.00112709f $X=7.845 $Y=2.315 $X2=0
+ $Y2=0
cc_829 N_A_991_81#_M1007_g N_VPWR_c_1855_n 0.00112709f $X=8.295 $Y=2.315 $X2=0
+ $Y2=0
cc_830 N_A_991_81#_c_984_n N_A_293_464#_c_2043_n 0.00564118f $X=5.24 $Y=2.265
+ $X2=0 $Y2=0
cc_831 N_A_991_81#_c_984_n N_A_293_464#_c_2050_n 0.0228445f $X=5.24 $Y=2.265
+ $X2=0 $Y2=0
cc_832 N_A_991_81#_c_991_n N_A_293_464#_c_2051_n 0.0165069f $X=5.24 $Y=2.39
+ $X2=0 $Y2=0
cc_833 N_A_991_81#_M1007_g N_A_1587_379#_c_2177_n 0.0138725f $X=8.295 $Y=2.315
+ $X2=0 $Y2=0
cc_834 N_A_991_81#_M1000_g N_A_1587_379#_c_2175_n 0.00939009f $X=7.845 $Y=2.315
+ $X2=0 $Y2=0
cc_835 N_A_991_81#_M1007_g N_A_1587_379#_c_2175_n 0.013314f $X=8.295 $Y=2.315
+ $X2=0 $Y2=0
cc_836 N_A_991_81#_M1007_g N_A_1587_379#_c_2176_n 0.00378019f $X=8.295 $Y=2.315
+ $X2=0 $Y2=0
cc_837 N_A_991_81#_c_982_n N_VGND_M1027_d 0.00373864f $X=7.755 $Y=0.955 $X2=0
+ $Y2=0
cc_838 N_A_991_81#_c_972_n N_VGND_c_2253_n 0.00149046f $X=7.07 $Y=0.865 $X2=0
+ $Y2=0
cc_839 N_A_991_81#_c_974_n N_VGND_c_2253_n 0.00600886f $X=8.13 $Y=1.085 $X2=0
+ $Y2=0
cc_840 N_A_991_81#_c_982_n N_VGND_c_2253_n 0.0290793f $X=7.755 $Y=0.955 $X2=0
+ $Y2=0
cc_841 N_A_991_81#_c_985_n N_VGND_c_2253_n 0.00136564f $X=7.92 $Y=1.39 $X2=0
+ $Y2=0
cc_842 N_A_991_81#_c_987_n N_VGND_c_2253_n 0.00113251f $X=8.295 $Y=1.32 $X2=0
+ $Y2=0
cc_843 N_A_991_81#_c_976_n N_VGND_c_2254_n 0.011645f $X=8.56 $Y=1.085 $X2=0
+ $Y2=0
cc_844 N_A_991_81#_c_972_n N_VGND_c_2258_n 0.00277351f $X=7.07 $Y=0.865 $X2=0
+ $Y2=0
cc_845 N_A_991_81#_c_978_n N_VGND_c_2259_n 0.00963155f $X=5.425 $Y=0.615 $X2=0
+ $Y2=0
cc_846 N_A_991_81#_c_972_n N_VGND_c_2262_n 0.00434272f $X=7.07 $Y=0.865 $X2=0
+ $Y2=0
cc_847 N_A_991_81#_c_974_n N_VGND_c_2263_n 0.00434272f $X=8.13 $Y=1.085 $X2=0
+ $Y2=0
cc_848 N_A_991_81#_c_976_n N_VGND_c_2263_n 0.00434272f $X=8.56 $Y=1.085 $X2=0
+ $Y2=0
cc_849 N_A_991_81#_c_972_n N_VGND_c_2274_n 0.00825979f $X=7.07 $Y=0.865 $X2=0
+ $Y2=0
cc_850 N_A_991_81#_c_974_n N_VGND_c_2274_n 0.00821975f $X=8.13 $Y=1.085 $X2=0
+ $Y2=0
cc_851 N_A_991_81#_c_976_n N_VGND_c_2274_n 0.00825283f $X=8.56 $Y=1.085 $X2=0
+ $Y2=0
cc_852 N_A_991_81#_c_978_n N_VGND_c_2274_n 0.00894247f $X=5.425 $Y=0.615 $X2=0
+ $Y2=0
cc_853 N_A_991_81#_c_974_n N_A_1641_74#_c_2411_n 0.00822305f $X=8.13 $Y=1.085
+ $X2=0 $Y2=0
cc_854 N_A_991_81#_c_976_n N_A_1641_74#_c_2411_n 0.0117724f $X=8.56 $Y=1.085
+ $X2=0 $Y2=0
cc_855 N_A_991_81#_c_982_n N_A_1641_74#_c_2411_n 8.79632e-19 $X=7.755 $Y=0.955
+ $X2=0 $Y2=0
cc_856 N_A_991_81#_c_976_n N_A_1641_74#_c_2412_n 0.0131495f $X=8.56 $Y=1.085
+ $X2=0 $Y2=0
cc_857 N_A_991_81#_c_974_n N_A_1641_74#_c_2413_n 0.00329746f $X=8.13 $Y=1.085
+ $X2=0 $Y2=0
cc_858 N_A_991_81#_c_976_n N_A_1641_74#_c_2413_n 0.00126919f $X=8.56 $Y=1.085
+ $X2=0 $Y2=0
cc_859 N_A_991_81#_c_982_n N_A_1641_74#_c_2413_n 0.00995113f $X=7.755 $Y=0.955
+ $X2=0 $Y2=0
cc_860 N_A_991_81#_c_986_n N_A_1641_74#_c_2413_n 8.54269e-19 $X=7.92 $Y=1.225
+ $X2=0 $Y2=0
cc_861 N_A_991_81#_c_987_n N_A_1641_74#_c_2413_n 0.00362919f $X=8.295 $Y=1.32
+ $X2=0 $Y2=0
cc_862 N_SET_B_M1021_g N_A_608_74#_c_1303_n 0.0112278f $X=7.21 $Y=2.525 $X2=0
+ $Y2=0
cc_863 N_SET_B_c_1155_n N_A_608_74#_c_1291_n 0.0158506f $X=11.615 $Y=1.295 $X2=0
+ $Y2=0
cc_864 N_SET_B_c_1155_n N_A_608_74#_M1044_g 0.00705218f $X=11.615 $Y=1.295 $X2=0
+ $Y2=0
cc_865 N_SET_B_M1013_g N_A_2186_367#_c_1490_n 0.0294304f $X=11.47 $Y=2.75 $X2=0
+ $Y2=0
cc_866 N_SET_B_M1025_g N_A_2186_367#_c_1482_n 0.00666993f $X=11.59 $Y=0.58 $X2=0
+ $Y2=0
cc_867 N_SET_B_c_1155_n N_A_2186_367#_c_1482_n 0.0036981f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_868 N_SET_B_c_1160_n N_A_2186_367#_c_1482_n 0.0294304f $X=11.61 $Y=1.635
+ $X2=0 $Y2=0
cc_869 N_SET_B_c_1161_n N_A_2186_367#_c_1482_n 0.00416418f $X=11.76 $Y=1.295
+ $X2=0 $Y2=0
cc_870 N_SET_B_M1025_g N_A_2186_367#_c_1483_n 0.0131197f $X=11.59 $Y=0.58 $X2=0
+ $Y2=0
cc_871 N_SET_B_c_1155_n N_A_2186_367#_c_1483_n 0.00814774f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_872 SET_B N_A_2186_367#_c_1483_n 0.00328346f $X=11.675 $Y=1.21 $X2=0 $Y2=0
cc_873 N_SET_B_c_1160_n N_A_2186_367#_c_1483_n 0.00258236f $X=11.61 $Y=1.635
+ $X2=0 $Y2=0
cc_874 N_SET_B_c_1161_n N_A_2186_367#_c_1483_n 0.0230245f $X=11.76 $Y=1.295
+ $X2=0 $Y2=0
cc_875 N_SET_B_M1013_g N_A_2186_367#_c_1493_n 0.00101182f $X=11.47 $Y=2.75 $X2=0
+ $Y2=0
cc_876 N_SET_B_M1013_g N_A_2186_367#_c_1495_n 7.16336e-19 $X=11.47 $Y=2.75 $X2=0
+ $Y2=0
cc_877 N_SET_B_M1025_g N_A_2186_367#_c_1486_n 0.00164729f $X=11.59 $Y=0.58 $X2=0
+ $Y2=0
cc_878 N_SET_B_c_1155_n N_A_2186_367#_c_1486_n 0.0202739f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_879 SET_B N_A_2186_367#_c_1486_n 2.21379e-19 $X=11.675 $Y=1.21 $X2=0 $Y2=0
cc_880 N_SET_B_c_1161_n N_A_2186_367#_c_1486_n 0.00377693f $X=11.76 $Y=1.295
+ $X2=0 $Y2=0
cc_881 N_SET_B_M1025_g N_A_2186_367#_c_1487_n 0.0182312f $X=11.59 $Y=0.58 $X2=0
+ $Y2=0
cc_882 N_SET_B_c_1155_n N_A_2186_367#_c_1487_n 0.00182071f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_883 N_SET_B_c_1161_n N_A_2186_367#_c_1487_n 3.01197e-19 $X=11.76 $Y=1.295
+ $X2=0 $Y2=0
cc_884 N_SET_B_M1025_g N_A_2186_367#_c_1489_n 0.0203492f $X=11.59 $Y=0.58 $X2=0
+ $Y2=0
cc_885 N_SET_B_M1025_g N_A_1804_424#_M1030_g 0.00849643f $X=11.59 $Y=0.58 $X2=0
+ $Y2=0
cc_886 N_SET_B_c_1155_n N_A_1804_424#_c_1592_n 0.0226921f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_887 N_SET_B_c_1155_n N_A_1804_424#_c_1593_n 0.0215392f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_888 N_SET_B_c_1160_n N_A_1804_424#_c_1593_n 3.78518e-19 $X=11.61 $Y=1.635
+ $X2=0 $Y2=0
cc_889 N_SET_B_c_1161_n N_A_1804_424#_c_1593_n 0.00736758f $X=11.76 $Y=1.295
+ $X2=0 $Y2=0
cc_890 N_SET_B_c_1160_n N_A_1804_424#_c_1595_n 0.00185705f $X=11.61 $Y=1.635
+ $X2=0 $Y2=0
cc_891 N_SET_B_c_1161_n N_A_1804_424#_c_1595_n 0.00867537f $X=11.76 $Y=1.295
+ $X2=0 $Y2=0
cc_892 N_SET_B_M1013_g N_A_1804_424#_c_1609_n 0.00992315f $X=11.47 $Y=2.75 $X2=0
+ $Y2=0
cc_893 SET_B N_A_1804_424#_c_1610_n 0.00102137f $X=11.675 $Y=1.21 $X2=0 $Y2=0
cc_894 N_SET_B_M1013_g N_A_1804_424#_c_1596_n 8.79832e-19 $X=11.47 $Y=2.75 $X2=0
+ $Y2=0
cc_895 N_SET_B_M1025_g N_A_1804_424#_c_1596_n 5.52256e-19 $X=11.59 $Y=0.58 $X2=0
+ $Y2=0
cc_896 SET_B N_A_1804_424#_c_1596_n 0.00702776f $X=11.675 $Y=1.21 $X2=0 $Y2=0
cc_897 N_SET_B_c_1160_n N_A_1804_424#_c_1596_n 3.63569e-19 $X=11.61 $Y=1.635
+ $X2=0 $Y2=0
cc_898 N_SET_B_c_1161_n N_A_1804_424#_c_1596_n 0.0327284f $X=11.76 $Y=1.295
+ $X2=0 $Y2=0
cc_899 N_SET_B_M1025_g N_A_1804_424#_c_1597_n 0.00770693f $X=11.59 $Y=0.58 $X2=0
+ $Y2=0
cc_900 SET_B N_A_1804_424#_c_1597_n 0.00460346f $X=11.675 $Y=1.21 $X2=0 $Y2=0
cc_901 N_SET_B_c_1160_n N_A_1804_424#_c_1597_n 0.0104335f $X=11.61 $Y=1.635
+ $X2=0 $Y2=0
cc_902 N_SET_B_c_1161_n N_A_1804_424#_c_1597_n 0.00510479f $X=11.76 $Y=1.295
+ $X2=0 $Y2=0
cc_903 N_SET_B_c_1155_n N_A_1804_424#_c_1657_n 0.00645725f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_904 N_SET_B_M1013_g N_A_1804_424#_c_1613_n 0.0316643f $X=11.47 $Y=2.75 $X2=0
+ $Y2=0
cc_905 N_SET_B_c_1155_n N_A_1804_424#_c_1613_n 0.0130421f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_906 SET_B N_A_1804_424#_c_1613_n 9.86625e-19 $X=11.675 $Y=1.21 $X2=0 $Y2=0
cc_907 N_SET_B_c_1160_n N_A_1804_424#_c_1613_n 0.00163909f $X=11.61 $Y=1.635
+ $X2=0 $Y2=0
cc_908 N_SET_B_c_1161_n N_A_1804_424#_c_1613_n 0.0357022f $X=11.76 $Y=1.295
+ $X2=0 $Y2=0
cc_909 N_SET_B_M1013_g N_A_1804_424#_c_1599_n 0.00647956f $X=11.47 $Y=2.75 $X2=0
+ $Y2=0
cc_910 N_SET_B_M1021_g N_VPWR_c_1861_n 0.00247204f $X=7.21 $Y=2.525 $X2=0 $Y2=0
cc_911 N_SET_B_M1013_g N_VPWR_c_1863_n 0.002979f $X=11.47 $Y=2.75 $X2=0 $Y2=0
cc_912 N_SET_B_M1013_g N_VPWR_c_1877_n 0.005209f $X=11.47 $Y=2.75 $X2=0 $Y2=0
cc_913 N_SET_B_M1013_g N_VPWR_c_1855_n 0.00543572f $X=11.47 $Y=2.75 $X2=0 $Y2=0
cc_914 N_SET_B_M1027_g N_VGND_c_2253_n 0.0159047f $X=7.46 $Y=0.58 $X2=0 $Y2=0
cc_915 N_SET_B_c_1155_n N_VGND_c_2253_n 0.00139039f $X=11.615 $Y=1.295 $X2=0
+ $Y2=0
cc_916 N_SET_B_M1027_g N_VGND_c_2262_n 0.00383152f $X=7.46 $Y=0.58 $X2=0 $Y2=0
cc_917 N_SET_B_M1025_g N_VGND_c_2271_n 0.00383152f $X=11.59 $Y=0.58 $X2=0 $Y2=0
cc_918 N_SET_B_M1025_g N_VGND_c_2272_n 0.0114386f $X=11.59 $Y=0.58 $X2=0 $Y2=0
cc_919 N_SET_B_M1027_g N_VGND_c_2274_n 0.0075725f $X=7.46 $Y=0.58 $X2=0 $Y2=0
cc_920 N_SET_B_M1025_g N_VGND_c_2274_n 0.00373161f $X=11.59 $Y=0.58 $X2=0 $Y2=0
cc_921 N_SET_B_M1027_g N_A_1641_74#_c_2411_n 0.00103176f $X=7.46 $Y=0.58 $X2=0
+ $Y2=0
cc_922 N_SET_B_c_1155_n N_A_1641_74#_c_2412_n 0.0321812f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_923 N_SET_B_c_1155_n N_A_1641_74#_c_2413_n 0.00922066f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_924 N_SET_B_c_1155_n N_A_1641_74#_c_2414_n 0.00864504f $X=11.615 $Y=1.295
+ $X2=0 $Y2=0
cc_925 N_A_608_74#_M1044_g N_A_2186_367#_c_1482_n 0.0191919f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_926 N_A_608_74#_M1044_g N_A_2186_367#_c_1486_n 0.00152879f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_927 N_A_608_74#_M1044_g N_A_2186_367#_c_1489_n 0.0512761f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_928 N_A_608_74#_M1003_g N_A_1804_424#_c_1604_n 0.0146934f $X=9.44 $Y=2.54
+ $X2=0 $Y2=0
cc_929 N_A_608_74#_c_1305_n N_A_1804_424#_c_1604_n 0.00211351f $X=9.8 $Y=3.15
+ $X2=0 $Y2=0
cc_930 N_A_608_74#_c_1306_n N_A_1804_424#_c_1604_n 0.0174109f $X=9.89 $Y=3.075
+ $X2=0 $Y2=0
cc_931 N_A_608_74#_c_1303_n N_A_1804_424#_c_1605_n 0.00909018f $X=9.35 $Y=3.15
+ $X2=0 $Y2=0
cc_932 N_A_608_74#_M1044_g N_A_1804_424#_c_1591_n 0.00520174f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_933 N_A_608_74#_c_1306_n N_A_1804_424#_c_1606_n 0.00763956f $X=9.89 $Y=3.075
+ $X2=0 $Y2=0
cc_934 N_A_608_74#_M1044_g N_A_1804_424#_c_1670_n 0.00385881f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_935 N_A_608_74#_M1044_g N_A_1804_424#_c_1592_n 0.0160324f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_936 N_A_608_74#_c_1306_n N_A_1804_424#_c_1607_n 0.00204088f $X=9.89 $Y=3.075
+ $X2=0 $Y2=0
cc_937 N_A_608_74#_c_1290_n N_A_1804_424#_c_1593_n 0.00361615f $X=10.555 $Y=1.52
+ $X2=0 $Y2=0
cc_938 N_A_608_74#_M1044_g N_A_1804_424#_c_1593_n 0.00274039f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_939 N_A_608_74#_c_1290_n N_A_1804_424#_c_1594_n 0.00972698f $X=10.555 $Y=1.52
+ $X2=0 $Y2=0
cc_940 N_A_608_74#_M1044_g N_A_1804_424#_c_1594_n 8.62813e-19 $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_941 N_A_608_74#_c_1290_n N_A_1804_424#_c_1595_n 5.16083e-19 $X=10.555 $Y=1.52
+ $X2=0 $Y2=0
cc_942 N_A_608_74#_c_1290_n N_A_1804_424#_c_1657_n 0.00374823f $X=10.555 $Y=1.52
+ $X2=0 $Y2=0
cc_943 N_A_608_74#_M1044_g N_A_1804_424#_c_1657_n 0.00327545f $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_944 N_A_608_74#_c_1312_n N_VPWR_M1032_d 0.00168223f $X=3.885 $Y=1.945 $X2=0
+ $Y2=0
cc_945 N_A_608_74#_M1040_g N_VPWR_c_1859_n 0.00887996f $X=3.935 $Y=2.4 $X2=0
+ $Y2=0
cc_946 N_A_608_74#_c_1299_n N_VPWR_c_1859_n 3.33864e-19 $X=4.455 $Y=3.075 $X2=0
+ $Y2=0
cc_947 N_A_608_74#_c_1301_n N_VPWR_c_1859_n 0.00232909f $X=4.53 $Y=3.15 $X2=0
+ $Y2=0
cc_948 N_A_608_74#_M1018_g N_VPWR_c_1860_n 0.00164269f $X=5.51 $Y=2.625 $X2=0
+ $Y2=0
cc_949 N_A_608_74#_c_1303_n N_VPWR_c_1860_n 0.0211465f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_950 N_A_608_74#_c_1303_n N_VPWR_c_1861_n 0.0170937f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_951 N_A_608_74#_c_1303_n N_VPWR_c_1862_n 0.0215219f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_952 N_A_608_74#_M1003_g N_VPWR_c_1862_n 4.91406e-19 $X=9.44 $Y=2.54 $X2=0
+ $Y2=0
cc_953 N_A_608_74#_M1040_g N_VPWR_c_1868_n 0.00460063f $X=3.935 $Y=2.4 $X2=0
+ $Y2=0
cc_954 N_A_608_74#_c_1301_n N_VPWR_c_1868_n 0.0424018f $X=4.53 $Y=3.15 $X2=0
+ $Y2=0
cc_955 N_A_608_74#_c_1303_n N_VPWR_c_1870_n 0.0290731f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_956 N_A_608_74#_c_1303_n N_VPWR_c_1872_n 0.0220248f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_957 N_A_608_74#_c_1303_n N_VPWR_c_1876_n 0.0331099f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_958 N_A_608_74#_M1040_g N_VPWR_c_1855_n 0.00909358f $X=3.935 $Y=2.4 $X2=0
+ $Y2=0
cc_959 N_A_608_74#_c_1300_n N_VPWR_c_1855_n 0.020954f $X=5.42 $Y=3.15 $X2=0
+ $Y2=0
cc_960 N_A_608_74#_c_1301_n N_VPWR_c_1855_n 0.00600101f $X=4.53 $Y=3.15 $X2=0
+ $Y2=0
cc_961 N_A_608_74#_c_1303_n N_VPWR_c_1855_n 0.105897f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_962 N_A_608_74#_c_1305_n N_VPWR_c_1855_n 0.0132544f $X=9.8 $Y=3.15 $X2=0
+ $Y2=0
cc_963 N_A_608_74#_c_1309_n N_VPWR_c_1855_n 0.00445211f $X=5.51 $Y=3.15 $X2=0
+ $Y2=0
cc_964 N_A_608_74#_c_1310_n N_VPWR_c_1855_n 0.00445015f $X=9.44 $Y=3.15 $X2=0
+ $Y2=0
cc_965 N_A_608_74#_c_1296_n N_A_293_464#_c_2039_n 0.00556071f $X=3.155 $Y=1.01
+ $X2=0 $Y2=0
cc_966 N_A_608_74#_c_1294_n N_A_293_464#_c_2041_n 0.00168773f $X=3.045 $Y=1.82
+ $X2=0 $Y2=0
cc_967 N_A_608_74#_M1032_s N_A_293_464#_c_2046_n 0.0111746f $X=3.125 $Y=1.84
+ $X2=0 $Y2=0
cc_968 N_A_608_74#_M1040_g N_A_293_464#_c_2046_n 0.0166424f $X=3.935 $Y=2.4
+ $X2=0 $Y2=0
cc_969 N_A_608_74#_c_1299_n N_A_293_464#_c_2046_n 0.0126173f $X=4.455 $Y=3.075
+ $X2=0 $Y2=0
cc_970 N_A_608_74#_c_1308_n N_A_293_464#_c_2046_n 0.0013146f $X=4.44 $Y=2.12
+ $X2=0 $Y2=0
cc_971 N_A_608_74#_c_1312_n N_A_293_464#_c_2046_n 0.0640258f $X=3.885 $Y=1.945
+ $X2=0 $Y2=0
cc_972 N_A_608_74#_c_1313_n N_A_293_464#_c_2046_n 8.29095e-19 $X=3.13 $Y=1.945
+ $X2=0 $Y2=0
cc_973 N_A_608_74#_c_1297_n N_A_293_464#_c_2046_n 0.00145017f $X=4.425 $Y=1.515
+ $X2=0 $Y2=0
cc_974 N_A_608_74#_c_1308_n N_A_293_464#_c_2047_n 0.00237977f $X=4.44 $Y=2.12
+ $X2=0 $Y2=0
cc_975 N_A_608_74#_c_1313_n N_A_293_464#_c_2048_n 0.0143305f $X=3.13 $Y=1.945
+ $X2=0 $Y2=0
cc_976 N_A_608_74#_c_1286_n N_A_293_464#_c_2042_n 0.00627096f $X=4.805 $Y=1.115
+ $X2=0 $Y2=0
cc_977 N_A_608_74#_c_1287_n N_A_293_464#_c_2042_n 7.52657e-19 $X=4.5 $Y=1.115
+ $X2=0 $Y2=0
cc_978 N_A_608_74#_M1024_g N_A_293_464#_c_2042_n 0.00370144f $X=4.88 $Y=0.615
+ $X2=0 $Y2=0
cc_979 N_A_608_74#_M1006_g N_A_293_464#_c_2043_n 0.00116188f $X=3.9 $Y=0.74
+ $X2=0 $Y2=0
cc_980 N_A_608_74#_M1040_g N_A_293_464#_c_2043_n 3.43045e-19 $X=3.935 $Y=2.4
+ $X2=0 $Y2=0
cc_981 N_A_608_74#_c_1285_n N_A_293_464#_c_2043_n 0.00609576f $X=4.425 $Y=1.35
+ $X2=0 $Y2=0
cc_982 N_A_608_74#_c_1286_n N_A_293_464#_c_2043_n 0.00700565f $X=4.805 $Y=1.115
+ $X2=0 $Y2=0
cc_983 N_A_608_74#_c_1287_n N_A_293_464#_c_2043_n 0.00416877f $X=4.5 $Y=1.115
+ $X2=0 $Y2=0
cc_984 N_A_608_74#_M1024_g N_A_293_464#_c_2043_n 0.0036657f $X=4.88 $Y=0.615
+ $X2=0 $Y2=0
cc_985 N_A_608_74#_c_1307_n N_A_293_464#_c_2043_n 0.0047582f $X=4.44 $Y=1.97
+ $X2=0 $Y2=0
cc_986 N_A_608_74#_c_1312_n N_A_293_464#_c_2043_n 0.0179403f $X=3.885 $Y=1.945
+ $X2=0 $Y2=0
cc_987 N_A_608_74#_c_1295_n N_A_293_464#_c_2043_n 0.0294141f $X=4.05 $Y=1.515
+ $X2=0 $Y2=0
cc_988 N_A_608_74#_c_1297_n N_A_293_464#_c_2043_n 0.0093602f $X=4.425 $Y=1.515
+ $X2=0 $Y2=0
cc_989 N_A_608_74#_c_1307_n N_A_293_464#_c_2050_n 0.00204597f $X=4.44 $Y=1.97
+ $X2=0 $Y2=0
cc_990 N_A_608_74#_c_1308_n N_A_293_464#_c_2050_n 0.00520632f $X=4.44 $Y=2.12
+ $X2=0 $Y2=0
cc_991 N_A_608_74#_c_1299_n N_A_293_464#_c_2051_n 0.00902539f $X=4.455 $Y=3.075
+ $X2=0 $Y2=0
cc_992 N_A_608_74#_M1003_g N_A_1587_379#_c_2174_n 0.0175812f $X=9.44 $Y=2.54
+ $X2=0 $Y2=0
cc_993 N_A_608_74#_c_1290_n N_A_1587_379#_c_2174_n 0.00141817f $X=10.555 $Y=1.52
+ $X2=0 $Y2=0
cc_994 N_A_608_74#_c_1306_n N_A_1587_379#_c_2174_n 0.00380755f $X=9.89 $Y=3.075
+ $X2=0 $Y2=0
cc_995 N_A_608_74#_M1003_g N_A_1587_379#_c_2190_n 0.0127899f $X=9.44 $Y=2.54
+ $X2=0 $Y2=0
cc_996 N_A_608_74#_c_1306_n N_A_1587_379#_c_2190_n 0.0136362f $X=9.89 $Y=3.075
+ $X2=0 $Y2=0
cc_997 N_A_608_74#_c_1303_n N_A_1587_379#_c_2175_n 0.00563439f $X=9.35 $Y=3.15
+ $X2=0 $Y2=0
cc_998 N_A_608_74#_M1003_g N_A_1587_379#_c_2176_n 0.00206087f $X=9.44 $Y=2.54
+ $X2=0 $Y2=0
cc_999 N_A_608_74#_c_1293_n N_VGND_c_2250_n 0.0328901f $X=3.185 $Y=0.515 $X2=0
+ $Y2=0
cc_1000 N_A_608_74#_c_1293_n N_VGND_c_2251_n 0.0172202f $X=3.185 $Y=0.515 $X2=0
+ $Y2=0
cc_1001 N_A_608_74#_M1006_g N_VGND_c_2252_n 0.0120099f $X=3.9 $Y=0.74 $X2=0
+ $Y2=0
cc_1002 N_A_608_74#_c_1293_n N_VGND_c_2252_n 0.026158f $X=3.185 $Y=0.515 $X2=0
+ $Y2=0
cc_1003 N_A_608_74#_M1006_g N_VGND_c_2259_n 0.00383152f $X=3.9 $Y=0.74 $X2=0
+ $Y2=0
cc_1004 N_A_608_74#_M1024_g N_VGND_c_2259_n 9.15902e-19 $X=4.88 $Y=0.615 $X2=0
+ $Y2=0
cc_1005 N_A_608_74#_M1044_g N_VGND_c_2271_n 0.00430908f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_1006 N_A_608_74#_M1006_g N_VGND_c_2274_n 0.00762539f $X=3.9 $Y=0.74 $X2=0
+ $Y2=0
cc_1007 N_A_608_74#_M1044_g N_VGND_c_2274_n 0.0081709f $X=10.63 $Y=0.58 $X2=0
+ $Y2=0
cc_1008 N_A_608_74#_c_1293_n N_VGND_c_2274_n 0.0142062f $X=3.185 $Y=0.515 $X2=0
+ $Y2=0
cc_1009 N_A_608_74#_c_1290_n N_A_1641_74#_c_2412_n 2.97622e-19 $X=10.555 $Y=1.52
+ $X2=0 $Y2=0
cc_1010 N_A_608_74#_c_1290_n N_A_1641_74#_c_2414_n 0.00134678f $X=10.555 $Y=1.52
+ $X2=0 $Y2=0
cc_1011 N_A_608_74#_M1044_g N_A_1641_74#_c_2414_n 2.88927e-19 $X=10.63 $Y=0.58
+ $X2=0 $Y2=0
cc_1012 N_A_2186_367#_c_1483_n N_A_1804_424#_M1030_g 0.012172f $X=12.5 $Y=0.875
+ $X2=0 $Y2=0
cc_1013 N_A_2186_367#_c_1484_n N_A_1804_424#_M1030_g 0.0010854f $X=12.64 $Y=0.58
+ $X2=0 $Y2=0
cc_1014 N_A_2186_367#_c_1485_n N_A_1804_424#_M1030_g 0.00600966f $X=12.72
+ $Y=2.31 $X2=0 $Y2=0
cc_1015 N_A_2186_367#_c_1488_n N_A_1804_424#_M1030_g 0.00339418f $X=12.652
+ $Y=0.875 $X2=0 $Y2=0
cc_1016 N_A_2186_367#_c_1493_n N_A_1804_424#_M1009_g 0.00352916f $X=12.225
+ $Y=2.75 $X2=0 $Y2=0
cc_1017 N_A_2186_367#_c_1494_n N_A_1804_424#_M1009_g 0.0180625f $X=12.635
+ $Y=2.395 $X2=0 $Y2=0
cc_1018 N_A_2186_367#_c_1485_n N_A_1804_424#_c_1587_n 0.0228379f $X=12.72
+ $Y=2.31 $X2=0 $Y2=0
cc_1019 N_A_2186_367#_c_1488_n N_A_1804_424#_c_1587_n 0.00532238f $X=12.652
+ $Y=0.875 $X2=0 $Y2=0
cc_1020 N_A_2186_367#_c_1484_n N_A_1804_424#_c_1588_n 0.00334701f $X=12.64
+ $Y=0.58 $X2=0 $Y2=0
cc_1021 N_A_2186_367#_c_1485_n N_A_1804_424#_c_1588_n 5.25537e-19 $X=12.72
+ $Y=2.31 $X2=0 $Y2=0
cc_1022 N_A_2186_367#_c_1485_n N_A_1804_424#_M1002_g 0.00212284f $X=12.72
+ $Y=2.31 $X2=0 $Y2=0
cc_1023 N_A_2186_367#_c_1494_n N_A_1804_424#_c_1602_n 3.45584e-19 $X=12.635
+ $Y=2.395 $X2=0 $Y2=0
cc_1024 N_A_2186_367#_c_1495_n N_A_1804_424#_c_1602_n 0.00135996f $X=12.31
+ $Y=2.395 $X2=0 $Y2=0
cc_1025 N_A_2186_367#_c_1485_n N_A_1804_424#_c_1602_n 0.0102395f $X=12.72
+ $Y=2.31 $X2=0 $Y2=0
cc_1026 N_A_2186_367#_c_1489_n N_A_1804_424#_c_1591_n 8.3456e-19 $X=11.11 $Y=0.9
+ $X2=0 $Y2=0
cc_1027 N_A_2186_367#_c_1489_n N_A_1804_424#_c_1670_n 0.00155017f $X=11.11
+ $Y=0.9 $X2=0 $Y2=0
cc_1028 N_A_2186_367#_c_1482_n N_A_1804_424#_c_1592_n 0.00119422f $X=11.02
+ $Y=1.835 $X2=0 $Y2=0
cc_1029 N_A_2186_367#_c_1482_n N_A_1804_424#_c_1593_n 0.00658133f $X=11.02
+ $Y=1.835 $X2=0 $Y2=0
cc_1030 N_A_2186_367#_c_1486_n N_A_1804_424#_c_1593_n 0.00748906f $X=11.11
+ $Y=0.875 $X2=0 $Y2=0
cc_1031 N_A_2186_367#_c_1490_n N_A_1804_424#_c_1595_n 0.00310124f $X=11.02
+ $Y=1.925 $X2=0 $Y2=0
cc_1032 N_A_2186_367#_M1008_g N_A_1804_424#_c_1595_n 0.00164141f $X=11.02
+ $Y=2.75 $X2=0 $Y2=0
cc_1033 N_A_2186_367#_c_1482_n N_A_1804_424#_c_1595_n 0.00880034f $X=11.02
+ $Y=1.835 $X2=0 $Y2=0
cc_1034 N_A_2186_367#_M1008_g N_A_1804_424#_c_1609_n 8.59873e-19 $X=11.02
+ $Y=2.75 $X2=0 $Y2=0
cc_1035 N_A_2186_367#_c_1493_n N_A_1804_424#_c_1609_n 0.036345f $X=12.225
+ $Y=2.75 $X2=0 $Y2=0
cc_1036 N_A_2186_367#_c_1495_n N_A_1804_424#_c_1609_n 3.9435e-19 $X=12.31
+ $Y=2.395 $X2=0 $Y2=0
cc_1037 N_A_2186_367#_c_1495_n N_A_1804_424#_c_1610_n 0.00628904f $X=12.31
+ $Y=2.395 $X2=0 $Y2=0
cc_1038 N_A_2186_367#_c_1494_n N_A_1804_424#_c_1611_n 0.0119564f $X=12.635
+ $Y=2.395 $X2=0 $Y2=0
cc_1039 N_A_2186_367#_c_1495_n N_A_1804_424#_c_1611_n 0.0155839f $X=12.31
+ $Y=2.395 $X2=0 $Y2=0
cc_1040 N_A_2186_367#_c_1485_n N_A_1804_424#_c_1611_n 0.0135424f $X=12.72
+ $Y=2.31 $X2=0 $Y2=0
cc_1041 N_A_2186_367#_c_1483_n N_A_1804_424#_c_1596_n 0.025786f $X=12.5 $Y=0.875
+ $X2=0 $Y2=0
cc_1042 N_A_2186_367#_c_1485_n N_A_1804_424#_c_1596_n 0.0618561f $X=12.72
+ $Y=2.31 $X2=0 $Y2=0
cc_1043 N_A_2186_367#_c_1483_n N_A_1804_424#_c_1597_n 0.00148844f $X=12.5
+ $Y=0.875 $X2=0 $Y2=0
cc_1044 N_A_2186_367#_c_1485_n N_A_1804_424#_c_1597_n 0.00182018f $X=12.72
+ $Y=2.31 $X2=0 $Y2=0
cc_1045 N_A_2186_367#_c_1488_n N_A_1804_424#_c_1597_n 4.75774e-19 $X=12.652
+ $Y=0.875 $X2=0 $Y2=0
cc_1046 N_A_2186_367#_c_1486_n N_A_1804_424#_c_1657_n 0.016946f $X=11.11
+ $Y=0.875 $X2=0 $Y2=0
cc_1047 N_A_2186_367#_c_1487_n N_A_1804_424#_c_1657_n 0.00155017f $X=11.11
+ $Y=1.065 $X2=0 $Y2=0
cc_1048 N_A_2186_367#_M1008_g N_A_1804_424#_c_1613_n 0.022796f $X=11.02 $Y=2.75
+ $X2=0 $Y2=0
cc_1049 N_A_2186_367#_c_1495_n N_A_1804_424#_c_1613_n 0.0136908f $X=12.31
+ $Y=2.395 $X2=0 $Y2=0
cc_1050 N_A_2186_367#_c_1485_n N_A_1804_424#_c_1599_n 0.0112411f $X=12.72
+ $Y=2.31 $X2=0 $Y2=0
cc_1051 N_A_2186_367#_c_1484_n N_A_2611_98#_c_1782_n 0.0214128f $X=12.64 $Y=0.58
+ $X2=0 $Y2=0
cc_1052 N_A_2186_367#_c_1485_n N_A_2611_98#_c_1782_n 0.0221171f $X=12.72 $Y=2.31
+ $X2=0 $Y2=0
cc_1053 N_A_2186_367#_c_1488_n N_A_2611_98#_c_1782_n 0.0121616f $X=12.652
+ $Y=0.875 $X2=0 $Y2=0
cc_1054 N_A_2186_367#_c_1494_n N_A_2611_98#_c_1788_n 0.0121746f $X=12.635
+ $Y=2.395 $X2=0 $Y2=0
cc_1055 N_A_2186_367#_c_1485_n N_A_2611_98#_c_1788_n 0.0423532f $X=12.72 $Y=2.31
+ $X2=0 $Y2=0
cc_1056 N_A_2186_367#_c_1485_n N_A_2611_98#_c_1784_n 0.0207869f $X=12.72 $Y=2.31
+ $X2=0 $Y2=0
cc_1057 N_A_2186_367#_M1008_g N_VPWR_c_1863_n 0.0109691f $X=11.02 $Y=2.75 $X2=0
+ $Y2=0
cc_1058 N_A_2186_367#_c_1493_n N_VPWR_c_1864_n 0.011548f $X=12.225 $Y=2.75 $X2=0
+ $Y2=0
cc_1059 N_A_2186_367#_c_1494_n N_VPWR_c_1864_n 0.0223822f $X=12.635 $Y=2.395
+ $X2=0 $Y2=0
cc_1060 N_A_2186_367#_M1008_g N_VPWR_c_1876_n 0.00460063f $X=11.02 $Y=2.75 $X2=0
+ $Y2=0
cc_1061 N_A_2186_367#_c_1493_n N_VPWR_c_1877_n 0.011054f $X=12.225 $Y=2.75 $X2=0
+ $Y2=0
cc_1062 N_A_2186_367#_M1008_g N_VPWR_c_1855_n 0.00464123f $X=11.02 $Y=2.75 $X2=0
+ $Y2=0
cc_1063 N_A_2186_367#_c_1493_n N_VPWR_c_1855_n 0.00915483f $X=12.225 $Y=2.75
+ $X2=0 $Y2=0
cc_1064 N_A_2186_367#_c_1494_n N_VPWR_c_1855_n 0.00677841f $X=12.635 $Y=2.395
+ $X2=0 $Y2=0
cc_1065 N_A_2186_367#_c_1484_n N_VGND_c_2264_n 0.013473f $X=12.64 $Y=0.58 $X2=0
+ $Y2=0
cc_1066 N_A_2186_367#_c_1489_n N_VGND_c_2271_n 0.00461464f $X=11.11 $Y=0.9 $X2=0
+ $Y2=0
cc_1067 N_A_2186_367#_c_1483_n N_VGND_c_2272_n 0.0458287f $X=12.5 $Y=0.875 $X2=0
+ $Y2=0
cc_1068 N_A_2186_367#_c_1484_n N_VGND_c_2272_n 0.0105067f $X=12.64 $Y=0.58 $X2=0
+ $Y2=0
cc_1069 N_A_2186_367#_c_1489_n N_VGND_c_2272_n 0.00163793f $X=11.11 $Y=0.9 $X2=0
+ $Y2=0
cc_1070 N_A_2186_367#_c_1483_n N_VGND_c_2274_n 0.0198116f $X=12.5 $Y=0.875 $X2=0
+ $Y2=0
cc_1071 N_A_2186_367#_c_1484_n N_VGND_c_2274_n 0.0111726f $X=12.64 $Y=0.58 $X2=0
+ $Y2=0
cc_1072 N_A_2186_367#_c_1486_n N_VGND_c_2274_n 0.0118158f $X=11.11 $Y=0.875
+ $X2=0 $Y2=0
cc_1073 N_A_2186_367#_c_1489_n N_VGND_c_2274_n 0.00451245f $X=11.11 $Y=0.9 $X2=0
+ $Y2=0
cc_1074 N_A_2186_367#_c_1486_n A_2219_74# 0.00386116f $X=11.11 $Y=0.875
+ $X2=-0.19 $Y2=-0.245
cc_1075 N_A_1804_424#_M1002_g N_A_2611_98#_M1004_g 0.0136985f $X=13.43 $Y=2.46
+ $X2=0 $Y2=0
cc_1076 N_A_1804_424#_c_1588_n N_A_2611_98#_M1014_g 0.0118486f $X=13.415
+ $Y=1.205 $X2=0 $Y2=0
cc_1077 N_A_1804_424#_c_1590_n N_A_2611_98#_M1014_g 0.00434128f $X=13.43
+ $Y=1.365 $X2=0 $Y2=0
cc_1078 N_A_1804_424#_M1030_g N_A_2611_98#_c_1782_n 6.58111e-19 $X=12.425
+ $Y=0.58 $X2=0 $Y2=0
cc_1079 N_A_1804_424#_c_1587_n N_A_2611_98#_c_1782_n 0.0126378f $X=13.34
+ $Y=1.365 $X2=0 $Y2=0
cc_1080 N_A_1804_424#_c_1588_n N_A_2611_98#_c_1782_n 0.0105297f $X=13.415
+ $Y=1.205 $X2=0 $Y2=0
cc_1081 N_A_1804_424#_c_1590_n N_A_2611_98#_c_1782_n 0.00227239f $X=13.43
+ $Y=1.365 $X2=0 $Y2=0
cc_1082 N_A_1804_424#_M1009_g N_A_2611_98#_c_1788_n 0.00610734f $X=12.45 $Y=2.75
+ $X2=0 $Y2=0
cc_1083 N_A_1804_424#_M1002_g N_A_2611_98#_c_1788_n 0.0233513f $X=13.43 $Y=2.46
+ $X2=0 $Y2=0
cc_1084 N_A_1804_424#_M1002_g N_A_2611_98#_c_1783_n 0.00994599f $X=13.43 $Y=2.46
+ $X2=0 $Y2=0
cc_1085 N_A_1804_424#_c_1590_n N_A_2611_98#_c_1783_n 0.0116487f $X=13.43
+ $Y=1.365 $X2=0 $Y2=0
cc_1086 N_A_1804_424#_c_1587_n N_A_2611_98#_c_1784_n 0.0146471f $X=13.34
+ $Y=1.365 $X2=0 $Y2=0
cc_1087 N_A_1804_424#_M1002_g N_A_2611_98#_c_1784_n 0.00285552f $X=13.43 $Y=2.46
+ $X2=0 $Y2=0
cc_1088 N_A_1804_424#_c_1590_n N_A_2611_98#_c_1784_n 8.38687e-19 $X=13.43
+ $Y=1.365 $X2=0 $Y2=0
cc_1089 N_A_1804_424#_c_1590_n N_A_2611_98#_c_1785_n 0.0215239f $X=13.43
+ $Y=1.365 $X2=0 $Y2=0
cc_1090 N_A_1804_424#_c_1603_n N_VPWR_c_1862_n 0.0265729f $X=9.165 $Y=2.4 $X2=0
+ $Y2=0
cc_1091 N_A_1804_424#_c_1605_n N_VPWR_c_1862_n 0.00960001f $X=9.33 $Y=2.99 $X2=0
+ $Y2=0
cc_1092 N_A_1804_424#_c_1604_n N_VPWR_c_1863_n 0.00498099f $X=10.105 $Y=2.99
+ $X2=0 $Y2=0
cc_1093 N_A_1804_424#_c_1606_n N_VPWR_c_1863_n 0.00685124f $X=10.27 $Y=2.745
+ $X2=0 $Y2=0
cc_1094 N_A_1804_424#_c_1609_n N_VPWR_c_1863_n 0.0117127f $X=11.695 $Y=2.75
+ $X2=0 $Y2=0
cc_1095 N_A_1804_424#_c_1613_n N_VPWR_c_1863_n 0.0186077f $X=11.86 $Y=2.222
+ $X2=0 $Y2=0
cc_1096 N_A_1804_424#_M1009_g N_VPWR_c_1864_n 0.0124849f $X=12.45 $Y=2.75 $X2=0
+ $Y2=0
cc_1097 N_A_1804_424#_M1002_g N_VPWR_c_1864_n 0.00345656f $X=13.43 $Y=2.46 $X2=0
+ $Y2=0
cc_1098 N_A_1804_424#_M1002_g N_VPWR_c_1865_n 0.00449062f $X=13.43 $Y=2.46 $X2=0
+ $Y2=0
cc_1099 N_A_1804_424#_c_1604_n N_VPWR_c_1876_n 0.0724435f $X=10.105 $Y=2.99
+ $X2=0 $Y2=0
cc_1100 N_A_1804_424#_c_1605_n N_VPWR_c_1876_n 0.0224969f $X=9.33 $Y=2.99 $X2=0
+ $Y2=0
cc_1101 N_A_1804_424#_M1009_g N_VPWR_c_1877_n 0.00460063f $X=12.45 $Y=2.75 $X2=0
+ $Y2=0
cc_1102 N_A_1804_424#_c_1609_n N_VPWR_c_1877_n 0.0142411f $X=11.695 $Y=2.75
+ $X2=0 $Y2=0
cc_1103 N_A_1804_424#_M1002_g N_VPWR_c_1878_n 0.005209f $X=13.43 $Y=2.46 $X2=0
+ $Y2=0
cc_1104 N_A_1804_424#_M1009_g N_VPWR_c_1855_n 0.00468499f $X=12.45 $Y=2.75 $X2=0
+ $Y2=0
cc_1105 N_A_1804_424#_M1002_g N_VPWR_c_1855_n 0.00987336f $X=13.43 $Y=2.46 $X2=0
+ $Y2=0
cc_1106 N_A_1804_424#_c_1604_n N_VPWR_c_1855_n 0.0390733f $X=10.105 $Y=2.99
+ $X2=0 $Y2=0
cc_1107 N_A_1804_424#_c_1605_n N_VPWR_c_1855_n 0.0113197f $X=9.33 $Y=2.99 $X2=0
+ $Y2=0
cc_1108 N_A_1804_424#_c_1609_n N_VPWR_c_1855_n 0.0118547f $X=11.695 $Y=2.75
+ $X2=0 $Y2=0
cc_1109 N_A_1804_424#_c_1612_n N_VPWR_c_1855_n 0.020251f $X=10.89 $Y=2.222 $X2=0
+ $Y2=0
cc_1110 N_A_1804_424#_c_1613_n N_VPWR_c_1855_n 0.00737176f $X=11.86 $Y=2.222
+ $X2=0 $Y2=0
cc_1111 N_A_1804_424#_c_1604_n N_A_1587_379#_M1003_d 0.00165831f $X=10.105
+ $Y=2.99 $X2=0 $Y2=0
cc_1112 N_A_1804_424#_M1003_s N_A_1587_379#_c_2174_n 0.0031013f $X=9.02 $Y=2.12
+ $X2=0 $Y2=0
cc_1113 N_A_1804_424#_c_1603_n N_A_1587_379#_c_2174_n 0.0238156f $X=9.165 $Y=2.4
+ $X2=0 $Y2=0
cc_1114 N_A_1804_424#_c_1604_n N_A_1587_379#_c_2190_n 0.0159318f $X=10.105
+ $Y=2.99 $X2=0 $Y2=0
cc_1115 N_A_1804_424#_c_1606_n N_A_1587_379#_c_2190_n 0.0139309f $X=10.27
+ $Y=2.745 $X2=0 $Y2=0
cc_1116 N_A_1804_424#_c_1607_n N_A_1587_379#_c_2190_n 0.00970031f $X=10.435
+ $Y=2.39 $X2=0 $Y2=0
cc_1117 N_A_1804_424#_c_1598_n N_VGND_c_2254_n 0.0310131f $X=9.415 $Y=0.34 $X2=0
+ $Y2=0
cc_1118 N_A_1804_424#_c_1588_n N_VGND_c_2255_n 0.00876736f $X=13.415 $Y=1.205
+ $X2=0 $Y2=0
cc_1119 N_A_1804_424#_M1030_g N_VGND_c_2264_n 0.00461464f $X=12.425 $Y=0.58
+ $X2=0 $Y2=0
cc_1120 N_A_1804_424#_c_1588_n N_VGND_c_2264_n 0.00473385f $X=13.415 $Y=1.205
+ $X2=0 $Y2=0
cc_1121 N_A_1804_424#_c_1591_n N_VGND_c_2271_n 0.0656534f $X=10.25 $Y=0.34 $X2=0
+ $Y2=0
cc_1122 N_A_1804_424#_c_1598_n N_VGND_c_2271_n 0.0228355f $X=9.415 $Y=0.34 $X2=0
+ $Y2=0
cc_1123 N_A_1804_424#_M1030_g N_VGND_c_2272_n 0.00435671f $X=12.425 $Y=0.58
+ $X2=0 $Y2=0
cc_1124 N_A_1804_424#_M1030_g N_VGND_c_2274_n 0.0045808f $X=12.425 $Y=0.58 $X2=0
+ $Y2=0
cc_1125 N_A_1804_424#_c_1588_n N_VGND_c_2274_n 0.00508379f $X=13.415 $Y=1.205
+ $X2=0 $Y2=0
cc_1126 N_A_1804_424#_c_1591_n N_VGND_c_2274_n 0.0365041f $X=10.25 $Y=0.34 $X2=0
+ $Y2=0
cc_1127 N_A_1804_424#_c_1598_n N_VGND_c_2274_n 0.0126251f $X=9.415 $Y=0.34 $X2=0
+ $Y2=0
cc_1128 N_A_1804_424#_c_1591_n N_A_1641_74#_M1001_s 0.00168754f $X=10.25 $Y=0.34
+ $X2=0 $Y2=0
cc_1129 N_A_1804_424#_M1001_d N_A_1641_74#_c_2412_n 0.0043689f $X=9.27 $Y=0.37
+ $X2=0 $Y2=0
cc_1130 N_A_1804_424#_c_1591_n N_A_1641_74#_c_2412_n 0.0037786f $X=10.25 $Y=0.34
+ $X2=0 $Y2=0
cc_1131 N_A_1804_424#_c_1598_n N_A_1641_74#_c_2412_n 0.024138f $X=9.415 $Y=0.34
+ $X2=0 $Y2=0
cc_1132 N_A_1804_424#_c_1591_n N_A_1641_74#_c_2414_n 0.0155812f $X=10.25 $Y=0.34
+ $X2=0 $Y2=0
cc_1133 N_A_1804_424#_c_1592_n N_A_1641_74#_c_2414_n 0.0109089f $X=10.495 $Y=1.4
+ $X2=0 $Y2=0
cc_1134 N_A_2611_98#_c_1788_n N_VPWR_c_1864_n 0.0249815f $X=13.205 $Y=2.105
+ $X2=0 $Y2=0
cc_1135 N_A_2611_98#_M1004_g N_VPWR_c_1865_n 0.00231368f $X=13.935 $Y=2.4 $X2=0
+ $Y2=0
cc_1136 N_A_2611_98#_c_1788_n N_VPWR_c_1865_n 0.0500555f $X=13.205 $Y=2.105
+ $X2=0 $Y2=0
cc_1137 N_A_2611_98#_c_1783_n N_VPWR_c_1865_n 0.0246466f $X=13.895 $Y=1.485
+ $X2=0 $Y2=0
cc_1138 N_A_2611_98#_c_1785_n N_VPWR_c_1865_n 0.00218979f $X=14.37 $Y=1.427
+ $X2=0 $Y2=0
cc_1139 N_A_2611_98#_M1004_g N_VPWR_c_1867_n 5.23753e-19 $X=13.935 $Y=2.4 $X2=0
+ $Y2=0
cc_1140 N_A_2611_98#_M1045_g N_VPWR_c_1867_n 0.0135584f $X=14.385 $Y=2.4 $X2=0
+ $Y2=0
cc_1141 N_A_2611_98#_c_1788_n N_VPWR_c_1878_n 0.0147721f $X=13.205 $Y=2.105
+ $X2=0 $Y2=0
cc_1142 N_A_2611_98#_M1004_g N_VPWR_c_1879_n 0.005209f $X=13.935 $Y=2.4 $X2=0
+ $Y2=0
cc_1143 N_A_2611_98#_M1045_g N_VPWR_c_1879_n 0.00460063f $X=14.385 $Y=2.4 $X2=0
+ $Y2=0
cc_1144 N_A_2611_98#_M1004_g N_VPWR_c_1855_n 0.00982203f $X=13.935 $Y=2.4 $X2=0
+ $Y2=0
cc_1145 N_A_2611_98#_M1045_g N_VPWR_c_1855_n 0.00908554f $X=14.385 $Y=2.4 $X2=0
+ $Y2=0
cc_1146 N_A_2611_98#_c_1788_n N_VPWR_c_1855_n 0.0121589f $X=13.205 $Y=2.105
+ $X2=0 $Y2=0
cc_1147 N_A_2611_98#_M1014_g N_Q_c_2208_n 0.00758611f $X=13.94 $Y=0.76 $X2=0
+ $Y2=0
cc_1148 N_A_2611_98#_c_1780_n N_Q_c_2208_n 0.00889128f $X=14.37 $Y=1.205 $X2=0
+ $Y2=0
cc_1149 N_A_2611_98#_M1004_g N_Q_c_2213_n 0.0103816f $X=13.935 $Y=2.4 $X2=0
+ $Y2=0
cc_1150 N_A_2611_98#_M1045_g N_Q_c_2213_n 3.83863e-19 $X=14.385 $Y=2.4 $X2=0
+ $Y2=0
cc_1151 N_A_2611_98#_M1014_g N_Q_c_2209_n 0.00253574f $X=13.94 $Y=0.76 $X2=0
+ $Y2=0
cc_1152 N_A_2611_98#_c_1780_n N_Q_c_2209_n 0.0024145f $X=14.37 $Y=1.205 $X2=0
+ $Y2=0
cc_1153 N_A_2611_98#_c_1783_n N_Q_c_2209_n 0.00111755f $X=13.895 $Y=1.485 $X2=0
+ $Y2=0
cc_1154 N_A_2611_98#_c_1785_n N_Q_c_2209_n 0.00215178f $X=14.37 $Y=1.427 $X2=0
+ $Y2=0
cc_1155 N_A_2611_98#_M1014_g N_Q_c_2210_n 0.00352031f $X=13.94 $Y=0.76 $X2=0
+ $Y2=0
cc_1156 N_A_2611_98#_c_1780_n N_Q_c_2210_n 0.0025985f $X=14.37 $Y=1.205 $X2=0
+ $Y2=0
cc_1157 N_A_2611_98#_c_1785_n N_Q_c_2210_n 0.0056321f $X=14.37 $Y=1.427 $X2=0
+ $Y2=0
cc_1158 N_A_2611_98#_c_1783_n N_Q_c_2211_n 0.0140641f $X=13.895 $Y=1.485 $X2=0
+ $Y2=0
cc_1159 N_A_2611_98#_c_1785_n N_Q_c_2211_n 0.0201262f $X=14.37 $Y=1.427 $X2=0
+ $Y2=0
cc_1160 N_A_2611_98#_M1004_g Q 0.0010146f $X=13.935 $Y=2.4 $X2=0 $Y2=0
cc_1161 N_A_2611_98#_M1045_g Q 0.00866136f $X=14.385 $Y=2.4 $X2=0 $Y2=0
cc_1162 N_A_2611_98#_c_1783_n Q 0.00775819f $X=13.895 $Y=1.485 $X2=0 $Y2=0
cc_1163 N_A_2611_98#_c_1785_n Q 0.00855109f $X=14.37 $Y=1.427 $X2=0 $Y2=0
cc_1164 N_A_2611_98#_M1004_g Q 0.00472141f $X=13.935 $Y=2.4 $X2=0 $Y2=0
cc_1165 N_A_2611_98#_M1045_g Q 0.020911f $X=14.385 $Y=2.4 $X2=0 $Y2=0
cc_1166 N_A_2611_98#_c_1783_n Q 7.50447e-19 $X=13.895 $Y=1.485 $X2=0 $Y2=0
cc_1167 N_A_2611_98#_c_1785_n Q 0.00247181f $X=14.37 $Y=1.427 $X2=0 $Y2=0
cc_1168 N_A_2611_98#_M1014_g N_VGND_c_2255_n 0.00737663f $X=13.94 $Y=0.76 $X2=0
+ $Y2=0
cc_1169 N_A_2611_98#_c_1782_n N_VGND_c_2255_n 0.0474865f $X=13.2 $Y=0.635 $X2=0
+ $Y2=0
cc_1170 N_A_2611_98#_c_1783_n N_VGND_c_2255_n 0.021633f $X=13.895 $Y=1.485 $X2=0
+ $Y2=0
cc_1171 N_A_2611_98#_c_1785_n N_VGND_c_2255_n 0.00172388f $X=14.37 $Y=1.427
+ $X2=0 $Y2=0
cc_1172 N_A_2611_98#_c_1780_n N_VGND_c_2257_n 0.00876453f $X=14.37 $Y=1.205
+ $X2=0 $Y2=0
cc_1173 N_A_2611_98#_c_1782_n N_VGND_c_2264_n 0.00977247f $X=13.2 $Y=0.635 $X2=0
+ $Y2=0
cc_1174 N_A_2611_98#_M1014_g N_VGND_c_2265_n 0.00537471f $X=13.94 $Y=0.76 $X2=0
+ $Y2=0
cc_1175 N_A_2611_98#_c_1780_n N_VGND_c_2265_n 0.0051044f $X=14.37 $Y=1.205 $X2=0
+ $Y2=0
cc_1176 N_A_2611_98#_M1014_g N_VGND_c_2274_n 0.00539454f $X=13.94 $Y=0.76 $X2=0
+ $Y2=0
cc_1177 N_A_2611_98#_c_1780_n N_VGND_c_2274_n 0.00539454f $X=14.37 $Y=1.205
+ $X2=0 $Y2=0
cc_1178 N_A_2611_98#_c_1782_n N_VGND_c_2274_n 0.0111804f $X=13.2 $Y=0.635 $X2=0
+ $Y2=0
cc_1179 N_VPWR_c_1856_n N_A_293_464#_c_2052_n 0.00764723f $X=0.73 $Y=2.78 $X2=0
+ $Y2=0
cc_1180 N_VPWR_c_1875_n N_A_293_464#_c_2052_n 0.0219007f $X=2.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1181 N_VPWR_c_1855_n N_A_293_464#_c_2052_n 0.0255415f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1182 N_VPWR_M1017_d N_A_293_464#_c_2045_n 0.00850355f $X=2.515 $Y=2.32 $X2=0
+ $Y2=0
cc_1183 N_VPWR_c_1857_n N_A_293_464#_c_2045_n 0.0245249f $X=2.725 $Y=2.995 $X2=0
+ $Y2=0
cc_1184 N_VPWR_c_1858_n N_A_293_464#_c_2045_n 0.00100823f $X=3.545 $Y=3.33 $X2=0
+ $Y2=0
cc_1185 N_VPWR_c_1875_n N_A_293_464#_c_2045_n 0.00235276f $X=2.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1186 N_VPWR_c_1855_n N_A_293_464#_c_2045_n 0.00734423f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1187 N_VPWR_M1032_d N_A_293_464#_c_2046_n 0.00332066f $X=3.575 $Y=1.84 $X2=0
+ $Y2=0
cc_1188 N_VPWR_c_1859_n N_A_293_464#_c_2046_n 0.0171101f $X=3.71 $Y=2.78 $X2=0
+ $Y2=0
cc_1189 N_VPWR_c_1875_n N_A_293_464#_c_2075_n 0.00468798f $X=2.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1190 N_VPWR_c_1855_n N_A_293_464#_c_2075_n 0.00569348f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1191 N_VPWR_c_1858_n N_A_293_464#_c_2048_n 0.00305321f $X=3.545 $Y=3.33 $X2=0
+ $Y2=0
cc_1192 N_VPWR_c_1859_n N_A_293_464#_c_2048_n 0.00302687f $X=3.71 $Y=2.78 $X2=0
+ $Y2=0
cc_1193 N_VPWR_c_1855_n N_A_293_464#_c_2048_n 0.00485809f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1194 N_VPWR_M1007_s N_A_1587_379#_c_2177_n 0.00437532f $X=8.385 $Y=1.895
+ $X2=0 $Y2=0
cc_1195 N_VPWR_c_1862_n N_A_1587_379#_c_2177_n 0.0124479f $X=8.52 $Y=2.58 $X2=0
+ $Y2=0
cc_1196 N_VPWR_c_1861_n N_A_1587_379#_c_2175_n 0.0177362f $X=7.62 $Y=2.23 $X2=0
+ $Y2=0
cc_1197 N_VPWR_c_1862_n N_A_1587_379#_c_2175_n 0.0122069f $X=8.52 $Y=2.58 $X2=0
+ $Y2=0
cc_1198 N_VPWR_c_1872_n N_A_1587_379#_c_2175_n 0.0074224f $X=8.435 $Y=3.33 $X2=0
+ $Y2=0
cc_1199 N_VPWR_c_1855_n N_A_1587_379#_c_2175_n 0.00904012f $X=14.64 $Y=3.33
+ $X2=0 $Y2=0
cc_1200 N_VPWR_M1007_s N_A_1587_379#_c_2176_n 0.00340727f $X=8.385 $Y=1.895
+ $X2=0 $Y2=0
cc_1201 N_VPWR_c_1862_n N_A_1587_379#_c_2176_n 0.00751656f $X=8.52 $Y=2.58 $X2=0
+ $Y2=0
cc_1202 N_VPWR_c_1865_n N_Q_c_2213_n 0.0311426f $X=13.705 $Y=2.085 $X2=0 $Y2=0
cc_1203 N_VPWR_c_1867_n N_Q_c_2213_n 0.0255358f $X=14.61 $Y=2.405 $X2=0 $Y2=0
cc_1204 N_VPWR_c_1879_n N_Q_c_2213_n 0.0123179f $X=14.445 $Y=3.33 $X2=0 $Y2=0
cc_1205 N_VPWR_c_1855_n N_Q_c_2213_n 0.0101276f $X=14.64 $Y=3.33 $X2=0 $Y2=0
cc_1206 N_VPWR_M1045_d Q 0.00385022f $X=14.475 $Y=1.84 $X2=0 $Y2=0
cc_1207 N_VPWR_c_1865_n Q 0.0145522f $X=13.705 $Y=2.085 $X2=0 $Y2=0
cc_1208 N_VPWR_c_1867_n Q 0.0212555f $X=14.61 $Y=2.405 $X2=0 $Y2=0
cc_1209 N_A_293_464#_c_2052_n A_419_464# 0.00393048f $X=2.215 $Y=2.785 $X2=-0.19
+ $Y2=-0.245
cc_1210 N_A_293_464#_c_2041_n A_419_464# 0.00139013f $X=2.3 $Y=2.49 $X2=-0.19
+ $Y2=-0.245
cc_1211 N_A_293_464#_c_2075_n A_419_464# 0.00335016f $X=2.3 $Y=2.575 $X2=-0.19
+ $Y2=-0.245
cc_1212 N_A_293_464#_c_2038_n N_VGND_c_2249_n 0.0107179f $X=1.725 $Y=0.58 $X2=0
+ $Y2=0
cc_1213 N_A_293_464#_c_2038_n N_VGND_c_2250_n 0.0108035f $X=1.725 $Y=0.58 $X2=0
+ $Y2=0
cc_1214 N_A_293_464#_c_2038_n N_VGND_c_2261_n 0.0144922f $X=1.725 $Y=0.58 $X2=0
+ $Y2=0
cc_1215 N_A_293_464#_c_2038_n N_VGND_c_2274_n 0.0118826f $X=1.725 $Y=0.58 $X2=0
+ $Y2=0
cc_1216 N_Q_c_2208_n N_VGND_c_2255_n 0.0558612f $X=14.155 $Y=0.535 $X2=0 $Y2=0
cc_1217 N_Q_c_2208_n N_VGND_c_2257_n 0.0596245f $X=14.155 $Y=0.535 $X2=0 $Y2=0
cc_1218 N_Q_c_2211_n N_VGND_c_2257_n 0.0217963f $X=14.465 $Y=1.49 $X2=0 $Y2=0
cc_1219 N_Q_c_2208_n N_VGND_c_2265_n 0.0143678f $X=14.155 $Y=0.535 $X2=0 $Y2=0
cc_1220 N_Q_c_2208_n N_VGND_c_2274_n 0.0128169f $X=14.155 $Y=0.535 $X2=0 $Y2=0
cc_1221 N_VGND_c_2253_n N_A_1641_74#_c_2411_n 0.0132241f $X=7.76 $Y=0.515 $X2=0
+ $Y2=0
cc_1222 N_VGND_c_2254_n N_A_1641_74#_c_2411_n 0.0138413f $X=8.855 $Y=0.53 $X2=0
+ $Y2=0
cc_1223 N_VGND_c_2263_n N_A_1641_74#_c_2411_n 0.0145302f $X=8.69 $Y=0 $X2=0
+ $Y2=0
cc_1224 N_VGND_c_2274_n N_A_1641_74#_c_2411_n 0.0118976f $X=14.64 $Y=0 $X2=0
+ $Y2=0
cc_1225 N_VGND_M1033_s N_A_1641_74#_c_2412_n 0.00454384f $X=8.635 $Y=0.37 $X2=0
+ $Y2=0
cc_1226 N_VGND_c_2254_n N_A_1641_74#_c_2412_n 0.0256711f $X=8.855 $Y=0.53 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__a2bb2oi_1.pxi.spice
* Created: Wed Sep  2 11:54:04 2020
* 
x_PM_SKY130_FD_SC_MS__A2BB2OI_1%A1_N N_A1_N_M1008_g N_A1_N_M1000_g A1_N
+ N_A1_N_c_66_n N_A1_N_c_67_n PM_SKY130_FD_SC_MS__A2BB2OI_1%A1_N
x_PM_SKY130_FD_SC_MS__A2BB2OI_1%A2_N N_A2_N_c_91_n N_A2_N_M1002_g N_A2_N_M1009_g
+ A2_N N_A2_N_c_93_n PM_SKY130_FD_SC_MS__A2BB2OI_1%A2_N
x_PM_SKY130_FD_SC_MS__A2BB2OI_1%A_126_112# N_A_126_112#_M1000_d
+ N_A_126_112#_M1002_d N_A_126_112#_M1004_g N_A_126_112#_c_134_n
+ N_A_126_112#_M1001_g N_A_126_112#_c_135_n N_A_126_112#_c_136_n
+ N_A_126_112#_c_137_n N_A_126_112#_c_138_n N_A_126_112#_c_139_n
+ N_A_126_112#_c_143_n N_A_126_112#_c_140_n N_A_126_112#_c_144_n
+ N_A_126_112#_c_141_n PM_SKY130_FD_SC_MS__A2BB2OI_1%A_126_112#
x_PM_SKY130_FD_SC_MS__A2BB2OI_1%B2 N_B2_M1006_g N_B2_M1007_g N_B2_c_208_n
+ N_B2_c_209_n B2 B2 N_B2_c_211_n PM_SKY130_FD_SC_MS__A2BB2OI_1%B2
x_PM_SKY130_FD_SC_MS__A2BB2OI_1%B1 N_B1_c_252_n N_B1_M1003_g N_B1_M1005_g B1
+ N_B1_c_255_n PM_SKY130_FD_SC_MS__A2BB2OI_1%B1
x_PM_SKY130_FD_SC_MS__A2BB2OI_1%VPWR N_VPWR_M1008_s N_VPWR_M1006_d
+ N_VPWR_c_282_n N_VPWR_c_283_n N_VPWR_c_284_n N_VPWR_c_285_n N_VPWR_c_286_n
+ N_VPWR_c_287_n VPWR N_VPWR_c_288_n N_VPWR_c_281_n
+ PM_SKY130_FD_SC_MS__A2BB2OI_1%VPWR
x_PM_SKY130_FD_SC_MS__A2BB2OI_1%Y N_Y_M1001_d N_Y_M1004_s N_Y_c_324_n
+ N_Y_c_336_n N_Y_c_325_n Y N_Y_c_328_n PM_SKY130_FD_SC_MS__A2BB2OI_1%Y
x_PM_SKY130_FD_SC_MS__A2BB2OI_1%A_402_368# N_A_402_368#_M1004_d
+ N_A_402_368#_M1005_d N_A_402_368#_c_371_n N_A_402_368#_c_378_n
+ N_A_402_368#_c_376_n N_A_402_368#_c_372_n N_A_402_368#_c_373_n
+ N_A_402_368#_c_374_n PM_SKY130_FD_SC_MS__A2BB2OI_1%A_402_368#
x_PM_SKY130_FD_SC_MS__A2BB2OI_1%VGND N_VGND_M1000_s N_VGND_M1009_d
+ N_VGND_M1003_d N_VGND_c_398_n N_VGND_c_399_n N_VGND_c_400_n N_VGND_c_401_n
+ VGND N_VGND_c_402_n N_VGND_c_403_n N_VGND_c_404_n N_VGND_c_405_n
+ PM_SKY130_FD_SC_MS__A2BB2OI_1%VGND
cc_1 VNB N_A1_N_M1008_g 0.00441374f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.46
cc_2 VNB N_A1_N_M1000_g 0.0237325f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.835
cc_3 VNB N_A1_N_c_66_n 0.00807592f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.425
cc_4 VNB N_A1_N_c_67_n 0.0633273f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.425
cc_5 VNB N_A2_N_c_91_n 0.0207996f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.59
cc_6 VNB N_A2_N_M1009_g 0.0306328f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.835
cc_7 VNB N_A2_N_c_93_n 0.0040235f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.425
cc_8 VNB N_A_126_112#_M1004_g 0.00676666f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_9 VNB N_A_126_112#_c_134_n 0.0192514f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.425
cc_10 VNB N_A_126_112#_c_135_n 0.0455804f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.425
cc_11 VNB N_A_126_112#_c_136_n 0.0106356f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.425
cc_12 VNB N_A_126_112#_c_137_n 0.00324684f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_13 VNB N_A_126_112#_c_138_n 0.00448426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_126_112#_c_139_n 0.00299965f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_126_112#_c_140_n 0.016101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_126_112#_c_141_n 0.00167709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B2_M1006_g 0.00625946f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.46
cc_18 VNB N_B2_c_208_n 0.0315615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B2_c_209_n 0.012229f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.425
cc_20 VNB B2 0.00266487f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.425
cc_21 VNB N_B2_c_211_n 0.0181973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B1_c_252_n 0.0214642f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.59
cc_23 VNB N_B1_M1005_g 0.00944953f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.835
cc_24 VNB B1 0.0113021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B1_c_255_n 0.0591523f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.425
cc_26 VNB N_VPWR_c_281_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_324_n 0.00408087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_325_n 0.00214178f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.425
cc_29 VNB N_VGND_c_398_n 0.0125919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_399_n 0.0476835f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.425
cc_31 VNB N_VGND_c_400_n 0.0129842f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.425
cc_32 VNB N_VGND_c_401_n 0.0350088f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.425
cc_33 VNB N_VGND_c_402_n 0.0198125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_403_n 0.029426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_404_n 0.037158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_405_n 0.220717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VPB N_A1_N_M1008_g 0.0366967f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.46
cc_38 VPB N_A1_N_c_66_n 0.00790246f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.425
cc_39 VPB N_A2_N_c_91_n 0.0180048f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.59
cc_40 VPB N_A2_N_M1002_g 0.0242051f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.46
cc_41 VPB N_A2_N_c_93_n 0.0084025f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.425
cc_42 VPB N_A_126_112#_M1004_g 0.027059f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_43 VPB N_A_126_112#_c_143_n 0.0111401f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A_126_112#_c_144_n 0.0139257f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A_126_112#_c_141_n 0.00590273f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_B2_M1006_g 0.0229798f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.46
cc_47 VPB B2 0.00409793f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=1.425
cc_48 VPB N_B1_M1005_g 0.0317187f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=0.835
cc_49 VPB N_VPWR_c_282_n 0.0121562f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=0.835
cc_50 VPB N_VPWR_c_283_n 0.051094f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_51 VPB N_VPWR_c_284_n 0.00540569f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.425
cc_52 VPB N_VPWR_c_285_n 0.00137138f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.665
cc_53 VPB N_VPWR_c_286_n 0.0561909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_287_n 0.00307912f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_288_n 0.0228467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_281_n 0.076547f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_Y_c_324_n 7.95989e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB Y 0.00641252f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_Y_c_328_n 0.00785683f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_402_368#_c_371_n 0.00201235f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_61 VPB N_A_402_368#_c_372_n 0.0234627f $X=-0.19 $Y=1.66 $X2=0.555 $Y2=1.425
cc_62 VPB N_A_402_368#_c_373_n 0.0180892f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_402_368#_c_374_n 0.00717518f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 N_A1_N_c_66_n N_A2_N_c_91_n 2.2065e-19 $X=0.27 $Y=1.425 $X2=-0.19
+ $Y2=-0.245
cc_65 N_A1_N_c_67_n N_A2_N_c_91_n 0.0510984f $X=0.51 $Y=1.425 $X2=-0.19
+ $Y2=-0.245
cc_66 N_A1_N_M1008_g N_A2_N_M1002_g 0.0470822f $X=0.51 $Y=2.46 $X2=0 $Y2=0
cc_67 N_A1_N_M1000_g N_A2_N_M1009_g 0.026924f $X=0.555 $Y=0.835 $X2=0 $Y2=0
cc_68 N_A1_N_c_66_n N_A2_N_M1009_g 8.21582e-19 $X=0.27 $Y=1.425 $X2=0 $Y2=0
cc_69 N_A1_N_c_67_n N_A2_N_M1009_g 0.00166236f $X=0.51 $Y=1.425 $X2=0 $Y2=0
cc_70 N_A1_N_c_66_n N_A2_N_c_93_n 0.026906f $X=0.27 $Y=1.425 $X2=0 $Y2=0
cc_71 N_A1_N_c_67_n N_A2_N_c_93_n 0.00355419f $X=0.51 $Y=1.425 $X2=0 $Y2=0
cc_72 N_A1_N_M1000_g N_A_126_112#_c_137_n 0.00609347f $X=0.555 $Y=0.835 $X2=0
+ $Y2=0
cc_73 N_A1_N_M1000_g N_A_126_112#_c_139_n 0.00485745f $X=0.555 $Y=0.835 $X2=0
+ $Y2=0
cc_74 N_A1_N_M1008_g N_A_126_112#_c_144_n 0.00280763f $X=0.51 $Y=2.46 $X2=0
+ $Y2=0
cc_75 N_A1_N_M1008_g N_VPWR_c_283_n 0.024801f $X=0.51 $Y=2.46 $X2=0 $Y2=0
cc_76 N_A1_N_c_66_n N_VPWR_c_283_n 0.0286221f $X=0.27 $Y=1.425 $X2=0 $Y2=0
cc_77 N_A1_N_c_67_n N_VPWR_c_283_n 0.00152171f $X=0.51 $Y=1.425 $X2=0 $Y2=0
cc_78 N_A1_N_M1008_g N_VPWR_c_286_n 0.00460063f $X=0.51 $Y=2.46 $X2=0 $Y2=0
cc_79 N_A1_N_M1008_g N_VPWR_c_281_n 0.00908061f $X=0.51 $Y=2.46 $X2=0 $Y2=0
cc_80 N_A1_N_M1000_g N_VGND_c_399_n 0.00759578f $X=0.555 $Y=0.835 $X2=0 $Y2=0
cc_81 N_A1_N_c_66_n N_VGND_c_399_n 0.0212796f $X=0.27 $Y=1.425 $X2=0 $Y2=0
cc_82 N_A1_N_c_67_n N_VGND_c_399_n 0.00195945f $X=0.51 $Y=1.425 $X2=0 $Y2=0
cc_83 N_A1_N_M1000_g N_VGND_c_402_n 0.0043356f $X=0.555 $Y=0.835 $X2=0 $Y2=0
cc_84 N_A1_N_M1000_g N_VGND_c_405_n 0.00487769f $X=0.555 $Y=0.835 $X2=0 $Y2=0
cc_85 N_A2_N_c_91_n N_A_126_112#_M1004_g 0.00303413f $X=0.9 $Y=1.83 $X2=0 $Y2=0
cc_86 N_A2_N_c_91_n N_A_126_112#_c_135_n 0.00622666f $X=0.9 $Y=1.83 $X2=0 $Y2=0
cc_87 N_A2_N_M1009_g N_A_126_112#_c_135_n 0.00790174f $X=0.985 $Y=0.835 $X2=0
+ $Y2=0
cc_88 N_A2_N_M1009_g N_A_126_112#_c_137_n 0.0115029f $X=0.985 $Y=0.835 $X2=0
+ $Y2=0
cc_89 N_A2_N_c_91_n N_A_126_112#_c_138_n 0.00310949f $X=0.9 $Y=1.83 $X2=0 $Y2=0
cc_90 N_A2_N_M1009_g N_A_126_112#_c_138_n 0.0131318f $X=0.985 $Y=0.835 $X2=0
+ $Y2=0
cc_91 N_A2_N_c_93_n N_A_126_112#_c_138_n 0.00723539f $X=1.005 $Y=1.615 $X2=0
+ $Y2=0
cc_92 N_A2_N_c_91_n N_A_126_112#_c_139_n 0.00189969f $X=0.9 $Y=1.83 $X2=0 $Y2=0
cc_93 N_A2_N_M1009_g N_A_126_112#_c_139_n 0.00204917f $X=0.985 $Y=0.835 $X2=0
+ $Y2=0
cc_94 N_A2_N_c_93_n N_A_126_112#_c_139_n 0.0179531f $X=1.005 $Y=1.615 $X2=0
+ $Y2=0
cc_95 N_A2_N_M1002_g N_A_126_112#_c_143_n 0.0160249f $X=0.9 $Y=2.46 $X2=0 $Y2=0
cc_96 N_A2_N_c_91_n N_A_126_112#_c_140_n 6.89529e-19 $X=0.9 $Y=1.83 $X2=0 $Y2=0
cc_97 N_A2_N_M1009_g N_A_126_112#_c_140_n 0.00852072f $X=0.985 $Y=0.835 $X2=0
+ $Y2=0
cc_98 N_A2_N_c_93_n N_A_126_112#_c_140_n 0.00833414f $X=1.005 $Y=1.615 $X2=0
+ $Y2=0
cc_99 N_A2_N_c_91_n N_A_126_112#_c_144_n 0.00637508f $X=0.9 $Y=1.83 $X2=0 $Y2=0
cc_100 N_A2_N_M1002_g N_A_126_112#_c_144_n 0.00365848f $X=0.9 $Y=2.46 $X2=0
+ $Y2=0
cc_101 N_A2_N_c_93_n N_A_126_112#_c_144_n 0.0115909f $X=1.005 $Y=1.615 $X2=0
+ $Y2=0
cc_102 N_A2_N_c_91_n N_A_126_112#_c_141_n 0.00419057f $X=0.9 $Y=1.83 $X2=0 $Y2=0
cc_103 N_A2_N_M1002_g N_A_126_112#_c_141_n 0.00369756f $X=0.9 $Y=2.46 $X2=0
+ $Y2=0
cc_104 N_A2_N_c_93_n N_A_126_112#_c_141_n 0.0178064f $X=1.005 $Y=1.615 $X2=0
+ $Y2=0
cc_105 N_A2_N_M1002_g N_VPWR_c_283_n 0.00335897f $X=0.9 $Y=2.46 $X2=0 $Y2=0
cc_106 N_A2_N_M1002_g N_VPWR_c_286_n 0.005209f $X=0.9 $Y=2.46 $X2=0 $Y2=0
cc_107 N_A2_N_M1002_g N_VPWR_c_281_n 0.00988003f $X=0.9 $Y=2.46 $X2=0 $Y2=0
cc_108 N_A2_N_M1002_g Y 6.07985e-19 $X=0.9 $Y=2.46 $X2=0 $Y2=0
cc_109 N_A2_N_M1002_g N_Y_c_328_n 9.90621e-19 $X=0.9 $Y=2.46 $X2=0 $Y2=0
cc_110 N_A2_N_M1009_g N_VGND_c_402_n 0.0043356f $X=0.985 $Y=0.835 $X2=0 $Y2=0
cc_111 N_A2_N_M1009_g N_VGND_c_404_n 0.0101051f $X=0.985 $Y=0.835 $X2=0 $Y2=0
cc_112 N_A2_N_M1009_g N_VGND_c_405_n 0.00487769f $X=0.985 $Y=0.835 $X2=0 $Y2=0
cc_113 N_A_126_112#_M1004_g N_B2_M1006_g 0.051661f $X=1.92 $Y=2.4 $X2=0 $Y2=0
cc_114 N_A_126_112#_c_136_n N_B2_c_208_n 0.0214626f $X=1.92 $Y=1.385 $X2=0 $Y2=0
cc_115 N_A_126_112#_c_136_n N_B2_c_209_n 3.62081e-19 $X=1.92 $Y=1.385 $X2=0
+ $Y2=0
cc_116 N_A_126_112#_c_134_n N_B2_c_211_n 0.0115596f $X=1.935 $Y=1.22 $X2=0 $Y2=0
cc_117 N_A_126_112#_c_144_n N_VPWR_c_283_n 0.0316443f $X=1.125 $Y=2.115 $X2=0
+ $Y2=0
cc_118 N_A_126_112#_M1004_g N_VPWR_c_284_n 5.40093e-19 $X=1.92 $Y=2.4 $X2=0
+ $Y2=0
cc_119 N_A_126_112#_M1004_g N_VPWR_c_286_n 0.005209f $X=1.92 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A_126_112#_c_143_n N_VPWR_c_286_n 0.014549f $X=1.125 $Y=2.815 $X2=0
+ $Y2=0
cc_121 N_A_126_112#_M1004_g N_VPWR_c_281_n 0.00988607f $X=1.92 $Y=2.4 $X2=0
+ $Y2=0
cc_122 N_A_126_112#_c_143_n N_VPWR_c_281_n 0.0119743f $X=1.125 $Y=2.815 $X2=0
+ $Y2=0
cc_123 N_A_126_112#_M1004_g N_Y_c_324_n 0.00581739f $X=1.92 $Y=2.4 $X2=0 $Y2=0
cc_124 N_A_126_112#_c_134_n N_Y_c_324_n 0.00510828f $X=1.935 $Y=1.22 $X2=0 $Y2=0
cc_125 N_A_126_112#_c_136_n N_Y_c_324_n 0.00931779f $X=1.92 $Y=1.385 $X2=0 $Y2=0
cc_126 N_A_126_112#_c_140_n N_Y_c_324_n 0.030479f $X=1.355 $Y=1.55 $X2=0 $Y2=0
cc_127 N_A_126_112#_c_141_n N_Y_c_324_n 0.00698697f $X=1.2 $Y=1.95 $X2=0 $Y2=0
cc_128 N_A_126_112#_c_134_n N_Y_c_336_n 0.0121303f $X=1.935 $Y=1.22 $X2=0 $Y2=0
cc_129 N_A_126_112#_c_140_n N_Y_c_336_n 0.00359949f $X=1.355 $Y=1.55 $X2=0 $Y2=0
cc_130 N_A_126_112#_M1004_g Y 0.023752f $X=1.92 $Y=2.4 $X2=0 $Y2=0
cc_131 N_A_126_112#_c_135_n Y 0.00581045f $X=1.83 $Y=1.385 $X2=0 $Y2=0
cc_132 N_A_126_112#_c_143_n Y 0.0170005f $X=1.125 $Y=2.815 $X2=0 $Y2=0
cc_133 N_A_126_112#_c_140_n Y 0.00749614f $X=1.355 $Y=1.55 $X2=0 $Y2=0
cc_134 N_A_126_112#_c_141_n Y 0.0312898f $X=1.2 $Y=1.95 $X2=0 $Y2=0
cc_135 N_A_126_112#_M1004_g N_Y_c_328_n 9.71144e-19 $X=1.92 $Y=2.4 $X2=0 $Y2=0
cc_136 N_A_126_112#_c_143_n N_Y_c_328_n 0.0361952f $X=1.125 $Y=2.815 $X2=0 $Y2=0
cc_137 N_A_126_112#_M1004_g N_A_402_368#_c_371_n 0.00640509f $X=1.92 $Y=2.4
+ $X2=0 $Y2=0
cc_138 N_A_126_112#_M1004_g N_A_402_368#_c_376_n 0.00369582f $X=1.92 $Y=2.4
+ $X2=0 $Y2=0
cc_139 N_A_126_112#_c_138_n N_VGND_M1009_d 0.0017426f $X=1.27 $Y=1.045 $X2=0
+ $Y2=0
cc_140 N_A_126_112#_c_140_n N_VGND_M1009_d 0.00480103f $X=1.355 $Y=1.55 $X2=0
+ $Y2=0
cc_141 N_A_126_112#_c_137_n N_VGND_c_399_n 0.0157455f $X=0.77 $Y=0.835 $X2=0
+ $Y2=0
cc_142 N_A_126_112#_c_137_n N_VGND_c_402_n 0.00800702f $X=0.77 $Y=0.835 $X2=0
+ $Y2=0
cc_143 N_A_126_112#_c_134_n N_VGND_c_403_n 0.00383152f $X=1.935 $Y=1.22 $X2=0
+ $Y2=0
cc_144 N_A_126_112#_c_134_n N_VGND_c_404_n 0.0120043f $X=1.935 $Y=1.22 $X2=0
+ $Y2=0
cc_145 N_A_126_112#_c_135_n N_VGND_c_404_n 0.00591277f $X=1.83 $Y=1.385 $X2=0
+ $Y2=0
cc_146 N_A_126_112#_c_137_n N_VGND_c_404_n 0.0103109f $X=0.77 $Y=0.835 $X2=0
+ $Y2=0
cc_147 N_A_126_112#_c_138_n N_VGND_c_404_n 0.0124114f $X=1.27 $Y=1.045 $X2=0
+ $Y2=0
cc_148 N_A_126_112#_c_140_n N_VGND_c_404_n 0.0262437f $X=1.355 $Y=1.55 $X2=0
+ $Y2=0
cc_149 N_A_126_112#_c_134_n N_VGND_c_405_n 0.00753023f $X=1.935 $Y=1.22 $X2=0
+ $Y2=0
cc_150 N_A_126_112#_c_137_n N_VGND_c_405_n 0.0105477f $X=0.77 $Y=0.835 $X2=0
+ $Y2=0
cc_151 N_B2_c_211_n N_B1_c_252_n 0.036204f $X=2.385 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_152 N_B2_M1006_g N_B1_M1005_g 0.0442613f $X=2.37 $Y=2.4 $X2=0 $Y2=0
cc_153 N_B2_c_208_n B1 2.21801e-19 $X=2.385 $Y=1.385 $X2=0 $Y2=0
cc_154 N_B2_c_209_n B1 0.0262884f $X=2.64 $Y=1.38 $X2=0 $Y2=0
cc_155 B2 B1 7.69126e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_156 N_B2_c_208_n N_B1_c_255_n 0.0209741f $X=2.385 $Y=1.385 $X2=0 $Y2=0
cc_157 N_B2_c_209_n N_B1_c_255_n 0.00279141f $X=2.64 $Y=1.38 $X2=0 $Y2=0
cc_158 B2 N_B1_c_255_n 0.00927777f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_159 B2 N_VPWR_M1006_d 0.00852692f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_160 N_B2_M1006_g N_VPWR_c_284_n 0.00351994f $X=2.37 $Y=2.4 $X2=0 $Y2=0
cc_161 N_B2_M1006_g N_VPWR_c_285_n 0.00367425f $X=2.37 $Y=2.4 $X2=0 $Y2=0
cc_162 N_B2_M1006_g N_VPWR_c_286_n 0.00460063f $X=2.37 $Y=2.4 $X2=0 $Y2=0
cc_163 N_B2_M1006_g N_VPWR_c_281_n 0.00443357f $X=2.37 $Y=2.4 $X2=0 $Y2=0
cc_164 N_B2_M1006_g N_Y_c_324_n 0.00156259f $X=2.37 $Y=2.4 $X2=0 $Y2=0
cc_165 N_B2_c_208_n N_Y_c_324_n 0.00103497f $X=2.385 $Y=1.385 $X2=0 $Y2=0
cc_166 N_B2_c_209_n N_Y_c_324_n 0.0249332f $X=2.64 $Y=1.38 $X2=0 $Y2=0
cc_167 B2 N_Y_c_324_n 0.00784186f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_168 N_B2_c_211_n N_Y_c_324_n 0.00215891f $X=2.385 $Y=1.22 $X2=0 $Y2=0
cc_169 N_B2_c_208_n N_Y_c_336_n 0.00148379f $X=2.385 $Y=1.385 $X2=0 $Y2=0
cc_170 N_B2_c_209_n N_Y_c_336_n 0.00483333f $X=2.64 $Y=1.38 $X2=0 $Y2=0
cc_171 N_B2_c_211_n N_Y_c_336_n 0.00359011f $X=2.385 $Y=1.22 $X2=0 $Y2=0
cc_172 N_B2_c_211_n N_Y_c_325_n 0.0101871f $X=2.385 $Y=1.22 $X2=0 $Y2=0
cc_173 N_B2_M1006_g Y 0.00104903f $X=2.37 $Y=2.4 $X2=0 $Y2=0
cc_174 N_B2_c_208_n Y 9.11254e-19 $X=2.385 $Y=1.385 $X2=0 $Y2=0
cc_175 N_B2_c_209_n Y 0.00114388f $X=2.64 $Y=1.38 $X2=0 $Y2=0
cc_176 B2 Y 0.00504648f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_177 N_B2_M1006_g N_A_402_368#_c_371_n 5.14662e-19 $X=2.37 $Y=2.4 $X2=0 $Y2=0
cc_178 N_B2_M1006_g N_A_402_368#_c_378_n 0.017603f $X=2.37 $Y=2.4 $X2=0 $Y2=0
cc_179 B2 N_A_402_368#_c_378_n 0.011053f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_180 B2 N_A_402_368#_c_372_n 0.00120069f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_181 N_B2_c_211_n N_VGND_c_401_n 0.00253877f $X=2.385 $Y=1.22 $X2=0 $Y2=0
cc_182 N_B2_c_211_n N_VGND_c_403_n 0.00434272f $X=2.385 $Y=1.22 $X2=0 $Y2=0
cc_183 N_B2_c_211_n N_VGND_c_404_n 6.57074e-19 $X=2.385 $Y=1.22 $X2=0 $Y2=0
cc_184 N_B2_c_211_n N_VGND_c_405_n 0.00821825f $X=2.385 $Y=1.22 $X2=0 $Y2=0
cc_185 N_B1_M1005_g N_VPWR_c_284_n 0.00232112f $X=2.85 $Y=2.4 $X2=0 $Y2=0
cc_186 N_B1_M1005_g N_VPWR_c_285_n 0.00404208f $X=2.85 $Y=2.4 $X2=0 $Y2=0
cc_187 N_B1_M1005_g N_VPWR_c_288_n 0.00519794f $X=2.85 $Y=2.4 $X2=0 $Y2=0
cc_188 N_B1_M1005_g N_VPWR_c_281_n 0.00521638f $X=2.85 $Y=2.4 $X2=0 $Y2=0
cc_189 N_B1_c_252_n N_Y_c_336_n 5.76856e-19 $X=2.835 $Y=1.22 $X2=0 $Y2=0
cc_190 N_B1_c_252_n N_Y_c_325_n 0.00160641f $X=2.835 $Y=1.22 $X2=0 $Y2=0
cc_191 N_B1_M1005_g N_A_402_368#_c_378_n 0.0164402f $X=2.85 $Y=2.4 $X2=0 $Y2=0
cc_192 N_B1_M1005_g N_A_402_368#_c_372_n 9.8167e-19 $X=2.85 $Y=2.4 $X2=0 $Y2=0
cc_193 B1 N_A_402_368#_c_372_n 0.0149782f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_194 N_B1_c_255_n N_A_402_368#_c_372_n 0.00185549f $X=3.09 $Y=1.385 $X2=0
+ $Y2=0
cc_195 N_B1_M1005_g N_A_402_368#_c_373_n 9.88899e-19 $X=2.85 $Y=2.4 $X2=0 $Y2=0
cc_196 N_B1_c_252_n N_VGND_c_401_n 0.0184513f $X=2.835 $Y=1.22 $X2=0 $Y2=0
cc_197 B1 N_VGND_c_401_n 0.0235157f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_198 N_B1_c_255_n N_VGND_c_401_n 0.001929f $X=3.09 $Y=1.385 $X2=0 $Y2=0
cc_199 N_B1_c_252_n N_VGND_c_403_n 0.00383152f $X=2.835 $Y=1.22 $X2=0 $Y2=0
cc_200 N_B1_c_252_n N_VGND_c_405_n 0.00757998f $X=2.835 $Y=1.22 $X2=0 $Y2=0
cc_201 N_VPWR_c_286_n N_Y_c_328_n 0.0110698f $X=2.43 $Y=3.33 $X2=0 $Y2=0
cc_202 N_VPWR_c_281_n N_Y_c_328_n 0.00916093f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_203 N_VPWR_c_285_n N_A_402_368#_c_371_n 0.00896295f $X=2.61 $Y=2.815 $X2=0
+ $Y2=0
cc_204 N_VPWR_c_286_n N_A_402_368#_c_371_n 0.0108673f $X=2.43 $Y=3.33 $X2=0
+ $Y2=0
cc_205 N_VPWR_c_281_n N_A_402_368#_c_371_n 0.00897581f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_206 N_VPWR_M1006_d N_A_402_368#_c_378_n 0.0044792f $X=2.46 $Y=1.84 $X2=0
+ $Y2=0
cc_207 N_VPWR_c_285_n N_A_402_368#_c_378_n 0.0174627f $X=2.61 $Y=2.815 $X2=0
+ $Y2=0
cc_208 N_VPWR_c_281_n N_A_402_368#_c_378_n 0.0127369f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_209 N_VPWR_c_285_n N_A_402_368#_c_373_n 0.00896295f $X=2.61 $Y=2.815 $X2=0
+ $Y2=0
cc_210 N_VPWR_c_288_n N_A_402_368#_c_373_n 0.011066f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_211 N_VPWR_c_281_n N_A_402_368#_c_373_n 0.00915947f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_212 Y N_A_402_368#_M1004_d 0.0084729f $X=2.075 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_213 N_Y_c_328_n N_A_402_368#_c_371_n 0.0139051f $X=1.695 $Y=1.985 $X2=0 $Y2=0
cc_214 Y N_A_402_368#_c_376_n 0.0156282f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_215 N_Y_c_336_n N_VGND_c_401_n 0.00365772f $X=2.185 $Y=0.88 $X2=0 $Y2=0
cc_216 N_Y_c_325_n N_VGND_c_401_n 0.0144183f $X=2.15 $Y=0.515 $X2=0 $Y2=0
cc_217 N_Y_c_325_n N_VGND_c_403_n 0.011237f $X=2.15 $Y=0.515 $X2=0 $Y2=0
cc_218 N_Y_c_336_n N_VGND_c_404_n 3.80876e-19 $X=2.185 $Y=0.88 $X2=0 $Y2=0
cc_219 N_Y_c_325_n N_VGND_c_404_n 0.0159304f $X=2.15 $Y=0.515 $X2=0 $Y2=0
cc_220 N_Y_c_325_n N_VGND_c_405_n 0.00933388f $X=2.15 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__dfxtp_2.spice
* Created: Fri Aug 28 17:25:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dfxtp_2.pex.spice"
.subckt sky130_fd_sc_ms__dfxtp_2  VNB VPB CLK D VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1024 N_VGND_M1024_d N_CLK_M1024_g N_A_27_74#_M1024_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1628 AS=0.2109 PD=1.18 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1025 N_A_209_368#_M1025_d N_A_27_74#_M1025_g N_VGND_M1024_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2775 AS=0.1628 PD=2.23 PS=1.18 NRD=14.592 NRS=25.944 M=1 R=4.93333
+ SA=75000.8 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1013 N_A_434_508#_M1013_d N_D_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.318675 PD=0.7 PS=2.49 NRD=0 NRS=201.06 M=1 R=2.8 SA=75000.5
+ SB=75003.1 A=0.063 P=1.14 MULT=1
MM1016 N_A_541_429#_M1016_d N_A_27_74#_M1016_g N_A_434_508#_M1013_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.076125 AS=0.0588 PD=0.835 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1015 A_708_101# N_A_209_368#_M1015_g N_A_541_429#_M1016_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.076125 PD=0.66 PS=0.835 NRD=18.564 NRS=7.14 M=1 R=2.8
+ SA=75001.1 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_695_459#_M1000_g A_708_101# VNB NLOWVT L=0.15 W=0.42
+ AD=0.180816 AS=0.0504 PD=1.2167 PS=0.66 NRD=107.28 NRS=18.564 M=1 R=2.8
+ SA=75001.5 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1003 N_A_695_459#_M1003_d N_A_541_429#_M1003_g N_VGND_M1000_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.236784 PD=0.83 PS=1.5933 NRD=0 NRS=73.08 M=1
+ R=3.66667 SA=75001.9 SB=75001.2 A=0.0825 P=1.4 MULT=1
MM1009 N_A_1022_424#_M1009_d N_A_209_368#_M1009_g N_A_695_459#_M1003_d VNB
+ NLOWVT L=0.15 W=0.55 AD=0.139229 AS=0.077 PD=1.33247 PS=0.83 NRD=32.724 NRS=0
+ M=1 R=3.66667 SA=75002.4 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1017 A_1172_124# N_A_27_74#_M1017_g N_A_1022_424#_M1009_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.106321 PD=0.66 PS=1.01753 NRD=18.564 NRS=22.848 M=1
+ R=2.8 SA=75002.7 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_1217_314#_M1001_g A_1172_124# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75003.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_1022_424#_M1020_g N_A_1217_314#_M1020_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.11405 AS=0.15675 PD=0.972093 PS=1.67 NRD=5.448 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75001.2 A=0.0825 P=1.4 MULT=1
MM1005 N_Q_M1005_d N_A_1217_314#_M1005_g N_VGND_M1020_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.15345 PD=1.02 PS=1.30791 NRD=0 NRS=15.396 M=1 R=4.93333
+ SA=75000.6 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1021 N_Q_M1005_d N_A_1217_314#_M1021_g N_VGND_M1021_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_VPWR_M1010_d N_CLK_M1010_g N_A_27_74#_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1011 N_A_209_368#_M1011_d N_A_27_74#_M1011_g N_VPWR_M1010_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1007 N_A_434_508#_M1007_d N_D_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=0.42
+ AD=0.109112 AS=0.2411 PD=1.17 PS=2.1 NRD=96.0375 NRS=243.453 M=1 R=2.33333
+ SA=90000.3 SB=90000.4 A=0.0756 P=1.2 MULT=1
MM1012 N_A_541_429#_M1012_d N_A_209_368#_M1012_g N_A_434_508#_M1007_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.106312 AS=0.109112 PD=1.145 PS=1.17 NRD=0 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90000.5 A=0.0756 P=1.2 MULT=1
MM1022 A_647_504# N_A_27_74#_M1022_g N_A_541_429#_M1012_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.106312 PD=0.66 PS=1.145 NRD=30.4759 NRS=92.9249 M=1
+ R=2.33333 SA=90000.3 SB=90003.2 A=0.0756 P=1.2 MULT=1
MM1002 N_VPWR_M1002_d N_A_695_459#_M1002_g A_647_504# VPB PSHORT L=0.18 W=0.42
+ AD=0.133583 AS=0.0504 PD=1.05 PS=0.66 NRD=123.381 NRS=30.4759 M=1 R=2.33333
+ SA=90000.7 SB=90002.7 A=0.0756 P=1.2 MULT=1
MM1004 N_A_695_459#_M1004_d N_A_541_429#_M1004_g N_VPWR_M1002_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2499 AS=0.267167 PD=1.435 PS=2.1 NRD=0 NRS=61.6807 M=1
+ R=4.66667 SA=90000.8 SB=90001.5 A=0.1512 P=2.04 MULT=1
MM1018 N_A_1022_424#_M1018_d N_A_27_74#_M1018_g N_A_695_459#_M1004_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.175 AS=0.2499 PD=1.58667 PS=1.435 NRD=0 NRS=73.8553 M=1
+ R=4.66667 SA=90001.5 SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1023 A_1128_508# N_A_209_368#_M1023_g N_A_1022_424#_M1018_d VPB PSHORT L=0.18
+ W=0.42 AD=0.09345 AS=0.0875 PD=0.865 PS=0.793333 NRD=78.5636 NRS=37.5088 M=1
+ R=2.33333 SA=90002.6 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1006 N_VPWR_M1006_d N_A_1217_314#_M1006_g A_1128_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.1155 AS=0.09345 PD=1.39 PS=0.865 NRD=0 NRS=78.5636 M=1 R=2.33333
+ SA=90003.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1019 N_VPWR_M1019_d N_A_1022_424#_M1019_g N_A_1217_314#_M1019_s VPB PSHORT
+ L=0.18 W=1 AD=0.167453 AS=0.28 PD=1.36321 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1008 N_Q_M1008_d N_A_1217_314#_M1008_g N_VPWR_M1019_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.187547 PD=1.39 PS=1.52679 NRD=0 NRS=8.7862 M=1 R=6.22222
+ SA=90000.6 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1014 N_Q_M1008_d N_A_1217_314#_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX26_noxref VNB VPB NWDIODE A=16.7772 P=21.76
c_1497 A_708_101# 0 4.2343e-20 $X=3.54 $Y=0.505
*
.include "sky130_fd_sc_ms__dfxtp_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__o32a_2.spice
* Created: Fri Aug 28 18:03:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o32a_2.pex.spice"
.subckt sky130_fd_sc_ms__o32a_2  VNB VPB A1 A2 A3 B2 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* B2	B2
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1010 N_X_M1010_d N_A_83_264#_M1010_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.3404 PD=1.02 PS=2.4 NRD=0 NRS=14.184 M=1 R=4.93333 SA=75000.4
+ SB=75003.8 A=0.111 P=1.78 MULT=1
MM1013 N_X_M1010_d N_A_83_264#_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.8
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1007 N_A_349_74#_M1007_d N_A1_M1007_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.4
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_A2_M1011_g N_A_349_74#_M1007_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.8
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1002 N_A_349_74#_M1002_d N_A3_M1002_g N_VGND_M1011_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1554 PD=1.09 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.4
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1001 N_A_83_264#_M1001_d N_B2_M1001_g N_A_349_74#_M1002_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.33855 AS=0.1295 PD=1.655 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75002.9 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1009 N_A_349_74#_M1009_d N_B1_M1009_g N_A_83_264#_M1001_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2627 AS=0.33855 PD=2.19 PS=1.655 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.9 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1004 N_X_M1004_d N_A_83_264#_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003.1 A=0.2016 P=2.6 MULT=1
MM1005 N_X_M1004_d N_A_83_264#_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.290566 PD=1.39 PS=1.73283 NRD=0 NRS=20.6653 M=1 R=6.22222
+ SA=90000.6 SB=90002.7 A=0.2016 P=2.6 MULT=1
MM1012 A_349_368# N_A1_M1012_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.259434 PD=1.24 PS=1.54717 NRD=12.7853 NRS=24.1128 M=1 R=5.55556
+ SA=90001.3 SB=90002.3 A=0.18 P=2.36 MULT=1
MM1000 A_433_368# N_A2_M1000_g A_349_368# VPB PSHORT L=0.18 W=1 AD=0.18 AS=0.12
+ PD=1.36 PS=1.24 NRD=24.6053 NRS=12.7853 M=1 R=5.55556 SA=90001.8 SB=90001.9
+ A=0.18 P=2.36 MULT=1
MM1006 N_A_83_264#_M1006_d N_A3_M1006_g A_433_368# VPB PSHORT L=0.18 W=1
+ AD=0.195 AS=0.18 PD=1.39 PS=1.36 NRD=10.8153 NRS=24.6053 M=1 R=5.55556
+ SA=90002.3 SB=90001.3 A=0.18 P=2.36 MULT=1
MM1003 A_655_368# N_B2_M1003_g N_A_83_264#_M1006_d VPB PSHORT L=0.18 W=1
+ AD=0.195 AS=0.195 PD=1.39 PS=1.39 NRD=27.5603 NRS=10.8153 M=1 R=5.55556
+ SA=90002.9 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_B1_M1008_g A_655_368# VPB PSHORT L=0.18 W=1 AD=0.28
+ AS=0.195 PD=2.56 PS=1.39 NRD=0 NRS=27.5603 M=1 R=5.55556 SA=90003.4 SB=90000.2
+ A=0.18 P=2.36 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_ms__o32a_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__a222oi_1.pex.spice
* Created: Wed Sep  2 11:52:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A222OI_1%C1 3 7 8 11 12 13
r30 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.43 $Y=1.285
+ $X2=0.43 $Y2=1.45
r31 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.43 $Y=1.285
+ $X2=0.43 $Y2=1.12
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.43
+ $Y=1.285 $X2=0.43 $Y2=1.285
r33 8 12 3.39186 $w=6.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.24 $Y=1.455
+ $X2=0.43 $Y2=1.455
r34 7 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.52 $Y=0.69 $X2=0.52
+ $Y2=1.12
r35 3 14 392.597 $w=1.8e-07 $l=1.01e-06 $layer=POLY_cond $X=0.505 $Y=2.46
+ $X2=0.505 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_MS__A222OI_1%C2 3 6 8 9 13 15
r35 13 16 78.1601 $w=4.8e-07 $l=5.05e-07 $layer=POLY_cond $X=1.075 $Y=1.285
+ $X2=1.075 $Y2=1.79
r36 13 15 45.9721 $w=4.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.075 $Y=1.285
+ $X2=1.075 $Y2=1.12
r37 8 9 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.15 $Y=1.285 $X2=1.15
+ $Y2=1.665
r38 8 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.15
+ $Y=1.285 $X2=1.15 $Y2=1.285
r39 6 16 260.435 $w=1.8e-07 $l=6.7e-07 $layer=POLY_cond $X=1.005 $Y=2.46
+ $X2=1.005 $Y2=1.79
r40 3 15 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.91 $Y=0.69 $X2=0.91
+ $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_MS__A222OI_1%B2 3 7 9 10 11 12 13 17
c39 11 0 8.91129e-20 $X=2.14 $Y=1.79
r40 12 13 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=2.14 $Y=1.285
+ $X2=2.14 $Y2=1.665
r41 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.14
+ $Y=1.285 $X2=2.14 $Y2=1.285
r42 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.14 $Y=1.625
+ $X2=2.14 $Y2=1.285
r43 10 11 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.14 $Y=1.625
+ $X2=2.14 $Y2=1.79
r44 9 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.14 $Y=1.12
+ $X2=2.14 $Y2=1.285
r45 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.23 $Y=0.69 $X2=2.23
+ $Y2=1.12
r46 3 11 260.435 $w=1.8e-07 $l=6.7e-07 $layer=POLY_cond $X=2.215 $Y=2.46
+ $X2=2.215 $Y2=1.79
.ends

.subckt PM_SKY130_FD_SC_MS__A222OI_1%B1 3 6 9 10 11 12 13 17
c40 6 0 1.71942e-19 $X=2.715 $Y=2.46
r41 12 13 12.5122 $w=3.48e-07 $l=3.8e-07 $layer=LI1_cond $X=2.7 $Y=1.285 $X2=2.7
+ $Y2=1.665
r42 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.71
+ $Y=1.285 $X2=2.71 $Y2=1.285
r43 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.71 $Y=1.625
+ $X2=2.71 $Y2=1.285
r44 10 11 34.9753 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.625
+ $X2=2.71 $Y2=1.79
r45 9 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.12
+ $X2=2.71 $Y2=1.285
r46 6 11 260.435 $w=1.8e-07 $l=6.7e-07 $layer=POLY_cond $X=2.715 $Y=2.46
+ $X2=2.715 $Y2=1.79
r47 3 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.62 $Y=0.69 $X2=2.62
+ $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_MS__A222OI_1%A1 2 5 9 10 11 12 16 17 18
r39 16 18 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=3.305 $Y=1.285
+ $X2=3.305 $Y2=1.12
r40 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.32
+ $Y=1.285 $X2=3.32 $Y2=1.285
r41 11 12 7.90266 $w=5.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.435 $Y=1.295
+ $X2=3.435 $Y2=1.665
r42 11 17 0.213585 $w=5.58e-07 $l=1e-08 $layer=LI1_cond $X=3.435 $Y=1.295
+ $X2=3.435 $Y2=1.285
r43 9 18 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.41 $Y=0.69 $X2=3.41
+ $Y2=1.12
r44 5 10 260.435 $w=1.8e-07 $l=6.7e-07 $layer=POLY_cond $X=3.215 $Y=2.46
+ $X2=3.215 $Y2=1.79
r45 2 10 43.2685 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=3.305 $Y=1.61
+ $X2=3.305 $Y2=1.79
r46 1 16 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=3.305 $Y=1.3
+ $X2=3.305 $Y2=1.285
r47 1 2 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=3.305 $Y=1.3 $X2=3.305
+ $Y2=1.61
.ends

.subckt PM_SKY130_FD_SC_MS__A222OI_1%A2 3 7 9 10 17
r28 15 17 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=3.815 $Y=1.345
+ $X2=4.05 $Y2=1.345
r29 13 15 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.8 $Y=1.345
+ $X2=3.815 $Y2=1.345
r30 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.05 $Y=1.295
+ $X2=4.05 $Y2=1.665
r31 9 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.05
+ $Y=1.345 $X2=4.05 $Y2=1.345
r32 5 15 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.815 $Y=1.51
+ $X2=3.815 $Y2=1.345
r33 5 7 369.274 $w=1.8e-07 $l=9.5e-07 $layer=POLY_cond $X=3.815 $Y=1.51
+ $X2=3.815 $Y2=2.46
r34 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.8 $Y=1.18 $X2=3.8
+ $Y2=1.345
r35 1 3 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=3.8 $Y=1.18 $X2=3.8
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__A222OI_1%Y 1 2 3 4 13 15 19 21 23 24 28 34 36 37 39
+ 40 41 56
c80 28 0 8.91129e-20 $X=1.57 $Y=1.96
r81 48 56 1.48702 $w=3.08e-07 $l=4e-08 $layer=LI1_cond $X=1.64 $Y=1.625 $X2=1.64
+ $Y2=1.665
r82 41 58 5.79065 $w=3.08e-07 $l=9.3e-08 $layer=LI1_cond $X=1.64 $Y=1.687
+ $X2=1.64 $Y2=1.78
r83 41 56 0.817863 $w=3.08e-07 $l=2.2e-08 $layer=LI1_cond $X=1.64 $Y=1.687
+ $X2=1.64 $Y2=1.665
r84 41 48 0.855038 $w=3.08e-07 $l=2.3e-08 $layer=LI1_cond $X=1.64 $Y=1.602
+ $X2=1.64 $Y2=1.625
r85 40 41 11.4129 $w=3.08e-07 $l=3.07e-07 $layer=LI1_cond $X=1.64 $Y=1.295
+ $X2=1.64 $Y2=1.602
r86 39 47 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=0.865
+ $X2=1.64 $Y2=0.95
r87 39 40 11.7103 $w=3.08e-07 $l=3.15e-07 $layer=LI1_cond $X=1.64 $Y=0.98
+ $X2=1.64 $Y2=1.295
r88 39 47 1.11527 $w=3.08e-07 $l=3e-08 $layer=LI1_cond $X=1.64 $Y=0.98 $X2=1.64
+ $Y2=0.95
r89 36 37 20.0288 $w=6.18e-07 $l=6.7e-07 $layer=LI1_cond $X=3.195 $Y=0.64
+ $X2=2.525 $Y2=0.64
r90 30 39 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.795 $Y=0.865
+ $X2=1.64 $Y2=0.865
r91 30 37 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.795 $Y=0.865
+ $X2=2.525 $Y2=0.865
r92 28 34 2.70057 $w=3.55e-07 $l=2.23495e-07 $layer=LI1_cond $X=1.57 $Y=1.96
+ $X2=1.385 $Y2=2.045
r93 28 58 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.57 $Y=1.96
+ $X2=1.57 $Y2=1.78
r94 23 39 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.485 $Y=0.865
+ $X2=1.64 $Y2=0.865
r95 23 24 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=1.485 $Y=0.865
+ $X2=0.47 $Y2=0.865
r96 22 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.045
+ $X2=0.28 $Y2=2.045
r97 21 34 4.08752 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=1.115 $Y=2.045
+ $X2=1.385 $Y2=2.045
r98 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=2.045
+ $X2=0.445 $Y2=2.045
r99 17 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.305 $Y=0.78
+ $X2=0.47 $Y2=0.865
r100 17 19 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.305 $Y=0.78
+ $X2=0.305 $Y2=0.515
r101 13 32 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.13 $X2=0.28
+ $Y2=2.045
r102 13 15 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=0.28 $Y=2.13
+ $X2=0.28 $Y2=2.815
r103 4 34 300 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_PDIFF $count=2 $X=1.095
+ $Y=1.96 $X2=1.28 $Y2=2.125
r104 3 32 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.125
r105 3 15 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r106 2 36 45.5 $w=1.7e-07 $l=5.59017e-07 $layer=licon1_NDIFF $count=4 $X=2.695
+ $Y=0.37 $X2=3.195 $Y2=0.495
r107 1 19 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.16
+ $Y=0.37 $X2=0.305 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A222OI_1%A_119_392# 1 2 9 11 12 15
r25 13 15 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=2.49 $Y=2.905
+ $X2=2.49 $Y2=2.465
r26 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.325 $Y=2.99
+ $X2=2.49 $Y2=2.905
r27 11 12 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.325 $Y=2.99
+ $X2=0.945 $Y2=2.99
r28 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.78 $Y=2.905
+ $X2=0.945 $Y2=2.99
r29 7 9 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.78 $Y=2.905 $X2=0.78
+ $Y2=2.465
r30 2 15 300 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_PDIFF $count=2 $X=2.305
+ $Y=1.96 $X2=2.49 $Y2=2.465
r31 1 9 300 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.96 $X2=0.78 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_MS__A222OI_1%A_369_392# 1 2 3 12 16 18 20 22 25 27
c42 16 0 1.71942e-19 $X=2.99 $Y=2.815
r43 20 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=2.13 $X2=4.04
+ $Y2=2.045
r44 20 22 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=4.04 $Y=2.13
+ $X2=4.04 $Y2=2.815
r45 19 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=2.045
+ $X2=2.99 $Y2=2.045
r46 18 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=2.045
+ $X2=4.04 $Y2=2.045
r47 18 19 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.875 $Y=2.045
+ $X2=3.155 $Y2=2.045
r48 14 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=2.13 $X2=2.99
+ $Y2=2.045
r49 14 16 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=2.99 $Y=2.13
+ $X2=2.99 $Y2=2.815
r50 13 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.155 $Y=2.045
+ $X2=1.99 $Y2=2.045
r51 12 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.825 $Y=2.045
+ $X2=2.99 $Y2=2.045
r52 12 13 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.825 $Y=2.045
+ $X2=2.155 $Y2=2.045
r53 3 29 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=1.96 $X2=4.04 $Y2=2.125
r54 3 22 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=1.96 $X2=4.04 $Y2=2.815
r55 2 27 400 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_PDIFF $count=1 $X=2.805
+ $Y=1.96 $X2=2.99 $Y2=2.125
r56 2 16 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=2.805
+ $Y=1.96 $X2=2.99 $Y2=2.815
r57 1 25 300 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=2 $X=1.845
+ $Y=1.96 $X2=1.99 $Y2=2.125
.ends

.subckt PM_SKY130_FD_SC_MS__A222OI_1%VPWR 1 6 9 10 11 21 22
r35 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r36 19 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r37 18 19 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 14 18 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 14 15 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 11 19 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 11 15 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=0.24 $Y2=3.33
r42 9 18 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.325 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.325 $Y=3.33
+ $X2=3.49 $Y2=3.33
r44 8 21 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.655 $Y=3.33
+ $X2=4.08 $Y2=3.33
r45 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.655 $Y=3.33
+ $X2=3.49 $Y2=3.33
r46 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.49 $Y=3.245 $X2=3.49
+ $Y2=3.33
r47 4 6 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=3.49 $Y=3.245 $X2=3.49
+ $Y2=2.465
r48 1 6 300 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_PDIFF $count=2 $X=3.305
+ $Y=1.96 $X2=3.49 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_MS__A222OI_1%VGND 1 2 7 9 11 18 25 37 40
r42 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r43 35 37 8.17678 $w=6.83e-07 $l=2e-08 $layer=LI1_cond $X=2.16 $Y=0.257 $X2=2.18
+ $Y2=0.257
r44 33 35 2.53184 $w=6.83e-07 $l=1.45e-07 $layer=LI1_cond $X=2.015 $Y=0.257
+ $X2=2.16 $Y2=0.257
r45 30 33 5.84943 $w=6.83e-07 $l=3.35e-07 $layer=LI1_cond $X=1.68 $Y=0.257
+ $X2=2.015 $Y2=0.257
r46 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r47 28 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r48 27 30 8.38128 $w=6.83e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=0.257
+ $X2=1.68 $Y2=0.257
r49 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r50 24 27 1.30957 $w=6.83e-07 $l=7.5e-08 $layer=LI1_cond $X=1.125 $Y=0.257
+ $X2=1.2 $Y2=0.257
r51 24 25 10.7086 $w=6.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.125 $Y=0.257
+ $X2=0.96 $Y2=0.257
r52 22 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r53 21 37 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=2.18
+ $Y2=0
r54 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r55 18 39 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.85 $Y=0 $X2=4.085
+ $Y2=0
r56 18 21 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.85 $Y=0 $X2=3.6
+ $Y2=0
r57 16 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r58 15 25 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=0.96
+ $Y2=0
r59 15 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r60 11 22 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r61 11 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r62 11 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r63 7 39 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=4.015 $Y=0.085
+ $X2=4.085 $Y2=0
r64 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.015 $Y=0.085
+ $X2=4.015 $Y2=0.515
r65 2 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.875
+ $Y=0.37 $X2=4.015 $Y2=0.515
r66 1 33 121.333 $w=1.7e-07 $l=1.10011e-06 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.37 $X2=2.015 $Y2=0.515
r67 1 24 121.333 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.37 $X2=1.125 $Y2=0.515
.ends


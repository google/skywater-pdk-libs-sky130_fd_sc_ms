* File: sky130_fd_sc_ms__and4bb_2.spice
* Created: Wed Sep  2 11:59:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__and4bb_2.pex.spice"
.subckt sky130_fd_sc_ms__and4bb_2  VNB VPB A_N C D B_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B_N	B_N
* D	D
* C	C
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1014 N_VGND_M1014_d N_A_N_M1014_g N_A_27_74#_M1014_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.15675 AS=0.15675 PD=1.67 PS=1.67 NRD=0 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1004 A_312_82# N_A_27_74#_M1004_g N_A_225_82#_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1002 A_390_82# N_A_354_252#_M1002_g A_312_82# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.0888 PD=1.13 PS=0.98 NRD=22.692 NRS=10.536 M=1 R=4.93333
+ SA=75000.6 SB=75003 A=0.111 P=1.78 MULT=1
MM1010 A_498_82# N_C_M1010_g A_390_82# VNB NLOWVT L=0.15 W=0.74 AD=0.1332
+ AS=0.1443 PD=1.1 PS=1.13 NRD=20.268 NRS=22.692 M=1 R=4.93333 SA=75001.1
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_D_M1011_g A_498_82# VNB NLOWVT L=0.15 W=0.74 AD=0.2553
+ AS=0.1332 PD=1.43 PS=1.1 NRD=0 NRS=20.268 M=1 R=4.93333 SA=75001.6 SB=75001.9
+ A=0.111 P=1.78 MULT=1
MM1003 N_X_M1003_d N_A_225_82#_M1003_g N_VGND_M1011_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2553 PD=1.02 PS=1.43 NRD=0 NRS=66.48 M=1 R=4.93333 SA=75002.5
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1007 N_X_M1003_d N_A_225_82#_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.216866 PD=1.02 PS=1.61767 NRD=0 NRS=38.604 M=1 R=4.93333
+ SA=75002.9 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1006 N_A_354_252#_M1006_d N_B_N_M1006_g N_VGND_M1007_s VNB NLOWVT L=0.15
+ W=0.55 AD=0.15675 AS=0.161184 PD=1.67 PS=1.20233 NRD=0 NRS=51.936 M=1
+ R=3.66667 SA=75003.5 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1015 N_VPWR_M1015_d N_A_N_M1015_g N_A_27_74#_M1015_s VPB PSHORT L=0.18 W=0.84
+ AD=0.170009 AS=0.2352 PD=1.26913 PS=2.24 NRD=27.5406 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90004.3 A=0.1512 P=2.04 MULT=1
MM1013 N_A_225_82#_M1013_d N_A_27_74#_M1013_g N_VPWR_M1015_d VPB PSHORT L=0.18
+ W=1 AD=0.27 AS=0.202391 PD=1.54 PS=1.51087 NRD=38.3953 NRS=0 M=1 R=5.55556
+ SA=90000.7 SB=90003.6 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_A_354_252#_M1012_g N_A_225_82#_M1013_d VPB PSHORT L=0.18
+ W=1 AD=0.24 AS=0.27 PD=1.48 PS=1.54 NRD=21.67 NRS=12.7853 M=1 R=5.55556
+ SA=90001.4 SB=90002.9 A=0.18 P=2.36 MULT=1
MM1000 N_A_225_82#_M1000_d N_C_M1000_g N_VPWR_M1012_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.24 PD=1.27 PS=1.48 NRD=0 NRS=17.73 M=1 R=5.55556 SA=90002
+ SB=90002.3 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_D_M1001_g N_A_225_82#_M1000_d VPB PSHORT L=0.18 W=1
+ AD=0.294811 AS=0.135 PD=1.61792 PS=1.27 NRD=26.5753 NRS=0 M=1 R=5.55556
+ SA=90002.5 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1008 N_X_M1008_d N_A_225_82#_M1008_g N_VPWR_M1001_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.330189 PD=1.39 PS=1.81208 NRD=0 NRS=31.6579 M=1 R=6.22222
+ SA=90002.9 SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1009 N_X_M1008_d N_A_225_82#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2152 PD=1.39 PS=1.68571 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.4
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1005 N_A_354_252#_M1005_d N_B_N_M1005_g N_VPWR_M1009_s VPB PSHORT L=0.18
+ W=0.84 AD=0.2478 AS=0.1614 PD=2.27 PS=1.26429 NRD=0 NRS=18.7544 M=1 R=4.66667
+ SA=90003.9 SB=90000.2 A=0.1512 P=2.04 MULT=1
DX16_noxref VNB VPB NWDIODE A=10.5276 P=15.04
c_48 VNB 0 1.18904e-19 $X=0 $Y=0
c_97 VPB 0 1.46091e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__and4bb_2.pxi.spice"
*
.ends
*
*

* NGSPICE file created from sky130_fd_sc_ms__a221o_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 VPWR A1 a_319_392# VPB pshort w=1e+06u l=180000u
+  ad=9.174e+11p pd=8.19e+06u as=5.4e+11p ps=5.08e+06u
M1001 a_89_260# A1 a_337_74# VNB nlowvt w=740000u l=150000u
+  ad=8.029e+11p pd=5.13e+06u as=1.554e+11p ps=1.9e+06u
M1002 X a_89_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=8.362e+11p ps=6.7e+06u
M1003 VGND a_89_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_319_392# B1 a_515_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=5.3e+11p ps=5.06e+06u
M1005 a_515_392# B2 a_319_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_89_260# C1 a_515_392# VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1007 a_337_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_603_74# B1 a_89_260# VNB nlowvt w=740000u l=150000u
+  ad=1.554e+11p pd=1.9e+06u as=0p ps=0u
M1009 VGND B2 a_603_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_89_260# C1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_89_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1012 VPWR a_89_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_319_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__o31a_4.pex.spice
* Created: Wed Sep  2 12:25:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O31A_4%A_86_260# 1 2 3 12 16 22 26 30 34 38 42 44 45
+ 56 59 61 63 67 71 73 75 77 84
c133 71 0 2.04502e-19 $X=2.465 $Y=1.3
c134 67 0 2.82748e-19 $X=3.105 $Y=0.77
c135 61 0 1.70893e-19 $X=2.94 $Y=1.215
c136 59 0 1.53462e-19 $X=2.63 $Y=2.815
c137 56 0 1.74626e-19 $X=2.63 $Y=2.105
c138 38 0 1.6164e-19 $X=1.83 $Y=0.74
r139 81 82 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=1.42 $Y=1.465
+ $X2=1.83 $Y2=1.465
r140 80 81 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.4 $Y=1.465 $X2=1.42
+ $Y2=1.465
r141 76 78 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.955 $Y=1.465
+ $X2=0.97 $Y2=1.465
r142 76 77 17.5095 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.955 $Y=1.465
+ $X2=0.88 $Y2=1.465
r143 65 67 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.105 $Y=1.13
+ $X2=3.105 $Y2=0.77
r144 64 73 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.715 $Y=2.46
+ $X2=2.59 $Y2=2.46
r145 63 75 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.925 $Y=2.46
+ $X2=4.09 $Y2=2.46
r146 63 64 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=3.925 $Y=2.46
+ $X2=2.715 $Y2=2.46
r147 62 71 5.16603 $w=2.5e-07 $l=2.89396e-07 $layer=LI1_cond $X=2.715 $Y=1.215
+ $X2=2.465 $Y2=1.3
r148 61 65 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.94 $Y=1.215
+ $X2=3.105 $Y2=1.13
r149 61 62 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.94 $Y=1.215
+ $X2=2.715 $Y2=1.215
r150 57 73 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=2.545
+ $X2=2.59 $Y2=2.46
r151 57 59 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=2.59 $Y=2.545
+ $X2=2.59 $Y2=2.815
r152 54 73 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=2.375
+ $X2=2.59 $Y2=2.46
r153 54 56 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=2.59 $Y=2.375
+ $X2=2.59 $Y2=2.105
r154 53 71 1.34256 $w=2.5e-07 $l=3.87492e-07 $layer=LI1_cond $X=2.59 $Y=1.63
+ $X2=2.465 $Y2=1.3
r155 53 56 21.8964 $w=2.48e-07 $l=4.75e-07 $layer=LI1_cond $X=2.59 $Y=1.63
+ $X2=2.59 $Y2=2.105
r156 52 84 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.85 $Y=1.465
+ $X2=1.87 $Y2=1.465
r157 52 82 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.85 $Y=1.465
+ $X2=1.83 $Y2=1.465
r158 51 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.85
+ $Y=1.465 $X2=1.85 $Y2=1.465
r159 48 80 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=1.17 $Y=1.465
+ $X2=1.4 $Y2=1.465
r160 48 78 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=1.17 $Y=1.465
+ $X2=0.97 $Y2=1.465
r161 47 51 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.17 $Y=1.465
+ $X2=1.85 $Y2=1.465
r162 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.465 $X2=1.17 $Y2=1.465
r163 45 71 5.16603 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=1.465
+ $X2=2.465 $Y2=1.3
r164 45 51 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.465 $Y=1.465
+ $X2=1.85 $Y2=1.465
r165 40 84 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.87 $Y=1.63
+ $X2=1.87 $Y2=1.465
r166 40 42 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.87 $Y=1.63
+ $X2=1.87 $Y2=2.4
r167 36 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.83 $Y=1.3
+ $X2=1.83 $Y2=1.465
r168 36 38 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.83 $Y=1.3
+ $X2=1.83 $Y2=0.74
r169 32 81 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=1.63
+ $X2=1.42 $Y2=1.465
r170 32 34 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.42 $Y=1.63
+ $X2=1.42 $Y2=2.4
r171 28 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.4 $Y=1.3 $X2=1.4
+ $Y2=1.465
r172 28 30 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.4 $Y=1.3 $X2=1.4
+ $Y2=0.74
r173 24 78 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.97 $Y=1.63
+ $X2=0.97 $Y2=1.465
r174 24 26 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.97 $Y=1.63
+ $X2=0.97 $Y2=2.4
r175 20 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.3
+ $X2=0.955 $Y2=1.465
r176 20 22 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.955 $Y=1.3
+ $X2=0.955 $Y2=0.74
r177 19 44 0.138649 $w=2.4e-07 $l=9e-08 $layer=POLY_cond $X=0.61 $Y=1.42
+ $X2=0.52 $Y2=1.42
r178 19 77 69.8776 $w=2.4e-07 $l=2.7e-07 $layer=POLY_cond $X=0.61 $Y=1.42
+ $X2=0.88 $Y2=1.42
r179 14 44 27.536 $w=1.65e-07 $l=1.22474e-07 $layer=POLY_cond $X=0.525 $Y=1.3
+ $X2=0.52 $Y2=1.42
r180 14 16 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.525 $Y=1.3
+ $X2=0.525 $Y2=0.74
r181 10 44 27.536 $w=1.65e-07 $l=1.2e-07 $layer=POLY_cond $X=0.52 $Y=1.54
+ $X2=0.52 $Y2=1.42
r182 10 12 334.29 $w=1.8e-07 $l=8.6e-07 $layer=POLY_cond $X=0.52 $Y=1.54
+ $X2=0.52 $Y2=2.4
r183 3 75 300 $w=1.7e-07 $l=5.63471e-07 $layer=licon1_PDIFF $count=2 $X=3.955
+ $Y=1.96 $X2=4.09 $Y2=2.46
r184 2 73 600 $w=1.7e-07 $l=5.63471e-07 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=1.96 $X2=2.63 $Y2=2.46
r185 2 59 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=1.96 $X2=2.63 $Y2=2.815
r186 2 56 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=1.96 $X2=2.63 $Y2=2.105
r187 1 67 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=2.915
+ $Y=0.625 $X2=3.105 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_4%B1 3 6 9 13 17 19 20 24 29
c58 29 0 1.00449e-19 $X=3.32 $Y=1.635
c59 13 0 1.53462e-19 $X=2.855 $Y=2.46
c60 9 0 3.30533e-19 $X=2.84 $Y=0.945
c61 3 0 2.02878e-19 $X=2.405 $Y=2.46
r62 27 29 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.07 $Y=1.635
+ $X2=3.32 $Y2=1.635
r63 25 27 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=2.855 $Y=1.635
+ $X2=3.07 $Y2=1.635
r64 23 25 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.84 $Y=1.635
+ $X2=2.855 $Y2=1.635
r65 23 24 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.84 $Y=1.635
+ $X2=2.765 $Y2=1.635
r66 19 20 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=3.07 $Y=1.635 $X2=3.07
+ $Y2=2.035
r67 19 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.07
+ $Y=1.635 $X2=3.07 $Y2=1.635
r68 15 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.32 $Y=1.47
+ $X2=3.32 $Y2=1.635
r69 15 17 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=3.32 $Y=1.47
+ $X2=3.32 $Y2=0.945
r70 11 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.855 $Y=1.8
+ $X2=2.855 $Y2=1.635
r71 11 13 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.855 $Y=1.8
+ $X2=2.855 $Y2=2.46
r72 7 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=1.47
+ $X2=2.84 $Y2=1.635
r73 7 9 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=2.84 $Y=1.47 $X2=2.84
+ $Y2=0.945
r74 6 24 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.495 $Y=1.545
+ $X2=2.765 $Y2=1.545
r75 1 6 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.405 $Y=1.62
+ $X2=2.495 $Y2=1.545
r76 1 3 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=2.405 $Y=1.62
+ $X2=2.405 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_4%A3 3 7 11 15 17 18 19 20 30
c54 11 0 1.51123e-19 $X=4.315 $Y=2.46
c55 7 0 2.84737e-19 $X=3.91 $Y=0.945
r56 30 31 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=4.315 $Y=1.62
+ $X2=4.34 $Y2=1.62
r57 28 30 11.055 $w=3.27e-07 $l=7.5e-08 $layer=POLY_cond $X=4.24 $Y=1.62
+ $X2=4.315 $Y2=1.62
r58 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.24
+ $Y=1.62 $X2=4.24 $Y2=1.62
r59 26 28 48.6422 $w=3.27e-07 $l=3.3e-07 $layer=POLY_cond $X=3.91 $Y=1.62
+ $X2=4.24 $Y2=1.62
r60 25 26 6.63303 $w=3.27e-07 $l=4.5e-08 $layer=POLY_cond $X=3.865 $Y=1.62
+ $X2=3.91 $Y2=1.62
r61 19 20 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.62
+ $X2=5.04 $Y2=1.62
r62 19 29 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=4.56 $Y=1.62
+ $X2=4.24 $Y2=1.62
r63 18 29 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.08 $Y=1.62 $X2=4.24
+ $Y2=1.62
r64 17 18 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.62 $X2=4.08
+ $Y2=1.62
r65 13 31 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.34 $Y=1.455
+ $X2=4.34 $Y2=1.62
r66 13 15 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.34 $Y=1.455
+ $X2=4.34 $Y2=0.945
r67 9 30 16.7191 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.315 $Y=1.785
+ $X2=4.315 $Y2=1.62
r68 9 11 262.379 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=4.315 $Y=1.785
+ $X2=4.315 $Y2=2.46
r69 5 26 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.91 $Y=1.455
+ $X2=3.91 $Y2=1.62
r70 5 7 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=3.91 $Y=1.455 $X2=3.91
+ $Y2=0.945
r71 1 25 16.7191 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.865 $Y=1.785
+ $X2=3.865 $Y2=1.62
r72 1 3 262.379 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.865 $Y=1.785
+ $X2=3.865 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_4%A1 3 7 11 15 17 25 26
c51 25 0 1.91258e-19 $X=5.71 $Y=1.62
c52 11 0 1.6294e-19 $X=5.7 $Y=0.945
r53 24 26 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=5.71 $Y=1.62
+ $X2=5.715 $Y2=1.62
r54 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.71
+ $Y=1.62 $X2=5.71 $Y2=1.62
r55 22 24 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=5.7 $Y=1.62 $X2=5.71
+ $Y2=1.62
r56 21 22 84.8077 $w=3.3e-07 $l=4.85e-07 $layer=POLY_cond $X=5.215 $Y=1.62
+ $X2=5.7 $Y2=1.62
r57 19 21 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.2 $Y=1.62
+ $X2=5.215 $Y2=1.62
r58 17 25 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=5.52 $Y=1.62
+ $X2=5.71 $Y2=1.62
r59 13 26 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.715 $Y=1.785
+ $X2=5.715 $Y2=1.62
r60 13 15 262.379 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=5.715 $Y=1.785
+ $X2=5.715 $Y2=2.46
r61 9 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.7 $Y=1.455 $X2=5.7
+ $Y2=1.62
r62 9 11 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=5.7 $Y=1.455 $X2=5.7
+ $Y2=0.945
r63 5 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.215 $Y=1.785
+ $X2=5.215 $Y2=1.62
r64 5 7 262.379 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=5.215 $Y=1.785
+ $X2=5.215 $Y2=2.46
r65 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.2 $Y=1.455 $X2=5.2
+ $Y2=1.62
r66 1 3 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=5.2 $Y=1.455 $X2=5.2
+ $Y2=0.945
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_4%A2 1 3 8 9 10 13 18 20 23
c60 8 0 1.44963e-19 $X=4.77 $Y=0.945
c61 3 0 3.42381e-19 $X=4.765 $Y=2.46
r62 23 26 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.28 $Y=1.62
+ $X2=6.28 $Y2=1.785
r63 23 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.28 $Y=1.62
+ $X2=6.28 $Y2=1.455
r64 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.28
+ $Y=1.62 $X2=6.28 $Y2=1.62
r65 20 24 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=6.48 $Y=1.62 $X2=6.28
+ $Y2=1.62
r66 18 25 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=6.2 $Y=0.945 $X2=6.2
+ $Y2=1.455
r67 15 18 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.2 $Y=0.255 $X2=6.2
+ $Y2=0.945
r68 13 26 262.379 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=6.205 $Y=2.46
+ $X2=6.205 $Y2=1.785
r69 9 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.125 $Y=0.18
+ $X2=6.2 $Y2=0.255
r70 9 10 656.34 $w=1.5e-07 $l=1.28e-06 $layer=POLY_cond $X=6.125 $Y=0.18
+ $X2=4.845 $Y2=0.18
r71 8 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.77 $Y=0.945
+ $X2=4.77 $Y2=1.34
r72 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.77 $Y=0.255
+ $X2=4.845 $Y2=0.18
r73 5 8 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.77 $Y=0.255 $X2=4.77
+ $Y2=0.945
r74 1 19 36.2738 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.765 $Y=1.43 $X2=4.765
+ $Y2=1.34
r75 1 3 400.371 $w=1.8e-07 $l=1.03e-06 $layer=POLY_cond $X=4.765 $Y=1.43
+ $X2=4.765 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_4%VPWR 1 2 3 4 5 16 18 24 28 34 38 41 42 43 49
+ 53 58 68 69 75 78 81
r90 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r91 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r92 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r93 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r94 69 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=5.52 $Y2=3.33
r95 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r96 66 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.605 $Y=3.33
+ $X2=5.44 $Y2=3.33
r97 66 68 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=5.605 $Y=3.33
+ $X2=6.48 $Y2=3.33
r98 65 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r99 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r100 62 65 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r101 61 64 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r102 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r103 59 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=3.33
+ $X2=3.08 $Y2=3.33
r104 59 61 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.245 $Y=3.33
+ $X2=3.6 $Y2=3.33
r105 58 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.275 $Y=3.33
+ $X2=5.44 $Y2=3.33
r106 58 64 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.275 $Y=3.33
+ $X2=5.04 $Y2=3.33
r107 57 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r108 57 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r109 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r110 54 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.26 $Y=3.33
+ $X2=2.135 $Y2=3.33
r111 54 56 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.26 $Y=3.33
+ $X2=2.64 $Y2=3.33
r112 53 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=3.08 $Y2=3.33
r113 53 56 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=2.64 $Y2=3.33
r114 52 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r115 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r116 49 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.01 $Y=3.33
+ $X2=2.135 $Y2=3.33
r117 49 51 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.01 $Y=3.33
+ $X2=1.68 $Y2=3.33
r118 48 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r119 48 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r120 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r121 45 72 3.99177 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.38 $Y=3.33
+ $X2=0.19 $Y2=3.33
r122 45 47 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.38 $Y=3.33
+ $X2=0.72 $Y2=3.33
r123 43 62 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.6 $Y2=3.33
r124 43 79 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r125 41 47 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.03 $Y=3.33
+ $X2=0.72 $Y2=3.33
r126 41 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.03 $Y=3.33
+ $X2=1.155 $Y2=3.33
r127 40 51 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.28 $Y=3.33 $X2=1.68
+ $Y2=3.33
r128 40 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.28 $Y=3.33
+ $X2=1.155 $Y2=3.33
r129 36 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.44 $Y=3.245
+ $X2=5.44 $Y2=3.33
r130 36 38 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=5.44 $Y=3.245
+ $X2=5.44 $Y2=2.8
r131 32 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.08 $Y2=3.33
r132 32 34 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.08 $Y2=2.805
r133 28 31 19.1306 $w=2.48e-07 $l=4.15e-07 $layer=LI1_cond $X=2.135 $Y=1.985
+ $X2=2.135 $Y2=2.4
r134 26 75 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.135 $Y=3.245
+ $X2=2.135 $Y2=3.33
r135 26 31 38.9526 $w=2.48e-07 $l=8.45e-07 $layer=LI1_cond $X=2.135 $Y=3.245
+ $X2=2.135 $Y2=2.4
r136 22 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=3.245
+ $X2=1.155 $Y2=3.33
r137 22 24 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=1.155 $Y=3.245
+ $X2=1.155 $Y2=2.305
r138 18 21 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.255 $Y=1.985
+ $X2=0.255 $Y2=2.815
r139 16 72 3.1514 $w=2.5e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.255 $Y=3.245
+ $X2=0.19 $Y2=3.33
r140 16 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.255 $Y=3.245
+ $X2=0.255 $Y2=2.815
r141 5 38 600 $w=1.7e-07 $l=9.04986e-07 $layer=licon1_PDIFF $count=1 $X=5.305
+ $Y=1.96 $X2=5.44 $Y2=2.8
r142 4 34 600 $w=1.7e-07 $l=9.1e-07 $layer=licon1_PDIFF $count=1 $X=2.945
+ $Y=1.96 $X2=3.08 $Y2=2.805
r143 3 31 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=1.96
+ $Y=1.84 $X2=2.095 $Y2=2.4
r144 3 28 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=1.84 $X2=2.095 $Y2=1.985
r145 2 24 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=1.06
+ $Y=1.84 $X2=1.195 $Y2=2.305
r146 1 21 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.84 $X2=0.295 $Y2=2.815
r147 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.84 $X2=0.295 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_4%X 1 2 3 4 13 15 19 23 27 28 29 30 31 32 33 50
+ 60
c64 15 0 1.6164e-19 $X=1.45 $Y=1.045
c65 13 0 9.88241e-20 $X=1.48 $Y=1.885
r66 57 60 0.664871 $w=2.58e-07 $l=1.5e-08 $layer=LI1_cond $X=0.705 $Y=1.97
+ $X2=0.705 $Y2=1.985
r67 43 50 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.74 $Y=0.96
+ $X2=0.74 $Y2=0.925
r68 32 33 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.705 $Y=2.405
+ $X2=0.705 $Y2=2.775
r69 31 52 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=1.885
+ $X2=0.705 $Y2=1.8
r70 31 57 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=1.885
+ $X2=0.705 $Y2=1.97
r71 31 32 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=0.705 $Y=2.045
+ $X2=0.705 $Y2=2.405
r72 31 60 2.65948 $w=2.58e-07 $l=6e-08 $layer=LI1_cond $X=0.705 $Y=2.045
+ $X2=0.705 $Y2=1.985
r73 30 52 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=1.8
r74 29 30 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.705 $Y=1.295
+ $X2=0.705 $Y2=1.665
r75 29 51 7.31358 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.705 $Y=1.295
+ $X2=0.705 $Y2=1.13
r76 28 43 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=1.045
+ $X2=0.74 $Y2=0.96
r77 28 51 3.19717 $w=2.95e-07 $l=1.00995e-07 $layer=LI1_cond $X=0.74 $Y=1.045
+ $X2=0.705 $Y2=1.13
r78 28 50 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.74 $Y=0.9
+ $X2=0.74 $Y2=0.925
r79 27 28 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.74 $Y=0.515
+ $X2=0.74 $Y2=0.9
r80 23 25 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.645 $Y=1.985
+ $X2=1.645 $Y2=2.815
r81 21 23 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.645 $Y=1.97
+ $X2=1.645 $Y2=1.985
r82 17 19 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=1.575 $Y=0.96
+ $X2=1.575 $Y2=0.515
r83 16 28 3.3845 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=1.045
+ $X2=0.74 $Y2=1.045
r84 15 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.45 $Y=1.045
+ $X2=1.575 $Y2=0.96
r85 15 16 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=1.45 $Y=1.045
+ $X2=0.905 $Y2=1.045
r86 14 31 2.90867 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.835 $Y=1.885
+ $X2=0.705 $Y2=1.885
r87 13 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.48 $Y=1.885
+ $X2=1.645 $Y2=1.97
r88 13 14 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.48 $Y=1.885
+ $X2=0.835 $Y2=1.885
r89 4 25 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.51
+ $Y=1.84 $X2=1.645 $Y2=2.815
r90 4 23 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.51
+ $Y=1.84 $X2=1.645 $Y2=1.985
r91 3 33 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.84 $X2=0.745 $Y2=2.815
r92 3 60 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.84 $X2=0.745 $Y2=1.985
r93 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.475
+ $Y=0.37 $X2=1.615 $Y2=0.515
r94 1 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.6
+ $Y=0.37 $X2=0.74 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_4%A_699_392# 1 2 3 10 16 18 20 22 25
c47 16 0 3.02247e-19 $X=4.54 $Y=2.475
r48 20 27 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.44 $Y=2.125 $X2=6.44
+ $Y2=2.04
r49 20 22 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=6.44 $Y=2.125
+ $X2=6.44 $Y2=2.815
r50 19 25 5.16603 $w=2.1e-07 $l=1.2339e-07 $layer=LI1_cond $X=4.645 $Y=2.04
+ $X2=4.54 $Y2=2.08
r51 18 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.275 $Y=2.04
+ $X2=6.44 $Y2=2.04
r52 18 19 106.342 $w=1.68e-07 $l=1.63e-06 $layer=LI1_cond $X=6.275 $Y=2.04
+ $X2=4.645 $Y2=2.04
r53 14 25 1.34256 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=4.54 $Y=2.205
+ $X2=4.54 $Y2=2.08
r54 14 16 14.2597 $w=2.08e-07 $l=2.7e-07 $layer=LI1_cond $X=4.54 $Y=2.205
+ $X2=4.54 $Y2=2.475
r55 10 25 5.16603 $w=2.1e-07 $l=1.05e-07 $layer=LI1_cond $X=4.435 $Y=2.08
+ $X2=4.54 $Y2=2.08
r56 10 12 36.6477 $w=2.48e-07 $l=7.95e-07 $layer=LI1_cond $X=4.435 $Y=2.08
+ $X2=3.64 $Y2=2.08
r57 3 27 400 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=1.96 $X2=6.44 $Y2=2.12
r58 3 22 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=1.96 $X2=6.44 $Y2=2.815
r59 2 25 600 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=1 $X=4.405
+ $Y=1.96 $X2=4.54 $Y2=2.12
r60 2 16 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=4.405
+ $Y=1.96 $X2=4.54 $Y2=2.475
r61 1 12 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=3.495
+ $Y=1.96 $X2=3.64 $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_4%A_971_392# 1 2 7 9 11 18
r25 12 16 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.075 $Y=2.38
+ $X2=4.95 $Y2=2.38
r26 11 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.775 $Y=2.38
+ $X2=5.94 $Y2=2.38
r27 11 12 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.775 $Y=2.38
+ $X2=5.075 $Y2=2.38
r28 7 16 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.95 $Y=2.465 $X2=4.95
+ $Y2=2.38
r29 7 9 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=4.95 $Y=2.465 $X2=4.95
+ $Y2=2.815
r30 2 18 300 $w=1.7e-07 $l=4.82804e-07 $layer=licon1_PDIFF $count=2 $X=5.805
+ $Y=1.96 $X2=5.94 $Y2=2.38
r31 1 16 600 $w=1.7e-07 $l=4.82804e-07 $layer=licon1_PDIFF $count=1 $X=4.855
+ $Y=1.96 $X2=4.99 $Y2=2.38
r32 1 9 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.855
+ $Y=1.96 $X2=4.99 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_4%VGND 1 2 3 4 5 6 19 21 25 29 33 37 41 44 45
+ 47 48 49 55 59 64 74 75 81 84 87
c96 59 0 1.61628e-19 $X=3.96 $Y=0
r97 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r98 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r99 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r100 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r101 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r102 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r103 72 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r104 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r105 69 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.15 $Y=0 $X2=4.985
+ $Y2=0
r106 69 71 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.15 $Y=0 $X2=5.52
+ $Y2=0
r107 68 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r108 68 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r109 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r110 65 84 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.085
+ $Y2=0
r111 65 67 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.56
+ $Y2=0
r112 64 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.82 $Y=0 $X2=4.985
+ $Y2=0
r113 64 67 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=4.82 $Y=0 $X2=4.56
+ $Y2=0
r114 63 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r115 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r116 60 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.045
+ $Y2=0
r117 60 62 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=2.21 $Y=0 $X2=3.6
+ $Y2=0
r118 59 84 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.96 $Y=0 $X2=4.085
+ $Y2=0
r119 59 62 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.96 $Y=0 $X2=3.6
+ $Y2=0
r120 58 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r121 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r122 55 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.88 $Y=0 $X2=2.045
+ $Y2=0
r123 55 57 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.88 $Y=0 $X2=1.68
+ $Y2=0
r124 54 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r125 54 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r126 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r127 51 78 3.97288 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0
+ $X2=0.197 $Y2=0
r128 51 53 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.395 $Y=0
+ $X2=0.72 $Y2=0
r129 49 63 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=3.6
+ $Y2=0
r130 49 82 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.36 $Y=0 $X2=2.16
+ $Y2=0
r131 47 71 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.75 $Y=0 $X2=5.52
+ $Y2=0
r132 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.75 $Y=0 $X2=5.915
+ $Y2=0
r133 46 74 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=6.08 $Y=0 $X2=6.48
+ $Y2=0
r134 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.08 $Y=0 $X2=5.915
+ $Y2=0
r135 44 53 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.085 $Y=0
+ $X2=0.72 $Y2=0
r136 44 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.085 $Y=0 $X2=1.17
+ $Y2=0
r137 43 57 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.255 $Y=0
+ $X2=1.68 $Y2=0
r138 43 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.17
+ $Y2=0
r139 39 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.915 $Y=0.085
+ $X2=5.915 $Y2=0
r140 39 41 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=5.915 $Y=0.085
+ $X2=5.915 $Y2=0.775
r141 35 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.985 $Y=0.085
+ $X2=4.985 $Y2=0
r142 35 37 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=4.985 $Y=0.085
+ $X2=4.985 $Y2=0.775
r143 31 84 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.085 $Y=0.085
+ $X2=4.085 $Y2=0
r144 31 33 31.8074 $w=2.48e-07 $l=6.9e-07 $layer=LI1_cond $X=4.085 $Y=0.085
+ $X2=4.085 $Y2=0.775
r145 27 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=0.085
+ $X2=2.045 $Y2=0
r146 27 29 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.045 $Y=0.085
+ $X2=2.045 $Y2=0.515
r147 23 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=0.085
+ $X2=1.17 $Y2=0
r148 23 25 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=1.17 $Y=0.085
+ $X2=1.17 $Y2=0.57
r149 19 78 3.17028 $w=2.5e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.197 $Y2=0
r150 19 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.27 $Y2=0.515
r151 6 41 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=5.775
+ $Y=0.625 $X2=5.915 $Y2=0.775
r152 5 37 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.625 $X2=4.985 $Y2=0.775
r153 4 33 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=3.985
+ $Y=0.625 $X2=4.125 $Y2=0.775
r154 3 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.905
+ $Y=0.37 $X2=2.045 $Y2=0.515
r155 2 25 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.37 $X2=1.17 $Y2=0.57
r156 1 21 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.165
+ $Y=0.37 $X2=0.31 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O31A_4%A_492_125# 1 2 3 4 5 18 20 21 25 26 27 30 32
+ 36 38 42 44 45
c86 36 0 1.6294e-19 $X=5.485 $Y=0.77
c87 30 0 1.44963e-19 $X=4.555 $Y=0.77
r88 40 42 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=6.415 $Y=1.115
+ $X2=6.415 $Y2=0.77
r89 39 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.57 $Y=1.2
+ $X2=5.445 $Y2=1.2
r90 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.25 $Y=1.2
+ $X2=6.415 $Y2=1.115
r91 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.25 $Y=1.2 $X2=5.57
+ $Y2=1.2
r92 34 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.445 $Y=1.115
+ $X2=5.445 $Y2=1.2
r93 34 36 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=5.445 $Y=1.115
+ $X2=5.445 $Y2=0.77
r94 33 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.64 $Y=1.2
+ $X2=4.515 $Y2=1.2
r95 32 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.32 $Y=1.2
+ $X2=5.445 $Y2=1.2
r96 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.32 $Y=1.2 $X2=4.64
+ $Y2=1.2
r97 28 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.515 $Y=1.115
+ $X2=4.515 $Y2=1.2
r98 28 30 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=4.515 $Y=1.115
+ $X2=4.515 $Y2=0.77
r99 26 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.39 $Y=1.2
+ $X2=4.515 $Y2=1.2
r100 26 27 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.39 $Y=1.2
+ $X2=3.78 $Y2=1.2
r101 23 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.615 $Y=1.115
+ $X2=3.78 $Y2=1.2
r102 23 25 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.615 $Y=1.115
+ $X2=3.615 $Y2=0.77
r103 22 25 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.615 $Y=0.435
+ $X2=3.615 $Y2=0.77
r104 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.45 $Y=0.35
+ $X2=3.615 $Y2=0.435
r105 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.45 $Y=0.35
+ $X2=2.77 $Y2=0.35
r106 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.605 $Y=0.435
+ $X2=2.77 $Y2=0.35
r107 16 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.605 $Y=0.435
+ $X2=2.605 $Y2=0.78
r108 5 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.275
+ $Y=0.625 $X2=6.415 $Y2=0.77
r109 4 36 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=5.275
+ $Y=0.625 $X2=5.485 $Y2=0.77
r110 3 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.415
+ $Y=0.625 $X2=4.555 $Y2=0.77
r111 2 25 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=3.395
+ $Y=0.625 $X2=3.615 $Y2=0.77
r112 1 18 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=2.46
+ $Y=0.625 $X2=2.605 $Y2=0.78
.ends


* File: sky130_fd_sc_ms__a22o_2.spice
* Created: Fri Aug 28 17:02:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a22o_2.pex.spice"
.subckt sky130_fd_sc_ms__a22o_2  VNB VPB A1 B1 B2 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* B2	B2
* B1	B1
* A1	A1
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_81_48#_M1002_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_81_48#_M1009_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_A_81_48#_M1008_d N_A1_M1008_g N_A_304_74#_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1006 A_491_74# N_B1_M1006_g N_A_81_48#_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.0925 AS=0.1295 PD=0.99 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1011_d N_B2_M1011_g A_491_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1443
+ AS=0.0925 PD=1.13 PS=0.99 NRD=6.48 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1004 N_A_304_74#_M1004_d N_A2_M1004_g N_VGND_M1011_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1443 PD=2.05 PS=1.13 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_X_M1005_d N_A_81_48#_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1007 N_X_M1005_d N_A_81_48#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.206038 PD=1.39 PS=1.56377 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90002 A=0.2016 P=2.6 MULT=1
MM1010 N_A_391_368#_M1010_d N_A1_M1010_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.183962 PD=1.27 PS=1.39623 NRD=0 NRS=16.7253 M=1 R=5.55556
+ SA=90001.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1003 N_A_81_48#_M1003_d N_B1_M1003_g N_A_391_368#_M1010_d VPB PSHORT L=0.18
+ W=1 AD=0.16 AS=0.135 PD=1.32 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.6
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1000 N_A_391_368#_M1000_d N_B2_M1000_g N_A_81_48#_M1003_d VPB PSHORT L=0.18
+ W=1 AD=0.17 AS=0.16 PD=1.34 PS=1.32 NRD=0.9653 NRS=8.8453 M=1 R=5.55556
+ SA=90002.1 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A2_M1001_g N_A_391_368#_M1000_d VPB PSHORT L=0.18 W=1
+ AD=0.26 AS=0.17 PD=2.52 PS=1.34 NRD=0 NRS=10.8153 M=1 R=5.55556 SA=90002.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
c_483 A_491_74# 0 1.11531e-19 $X=2.455 $Y=0.37
*
.include "sky130_fd_sc_ms__a22o_2.pxi.spice"
*
.ends
*
*

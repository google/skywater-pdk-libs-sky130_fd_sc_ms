* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or4_4 A B C D VGND VNB VPB VPWR X
X0 VGND C a_83_264# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_83_264# D a_965_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X2 VGND B a_83_264# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_83_264# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 X a_83_264# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 a_591_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X6 X a_83_264# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 a_83_264# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_965_392# D a_83_264# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X9 VGND a_83_264# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_591_392# B a_499_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X11 VGND a_83_264# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VPWR a_83_264# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X13 a_965_392# C a_499_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X14 a_499_392# B a_591_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X15 VPWR A a_591_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X16 a_499_392# C a_965_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X17 X a_83_264# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 VPWR a_83_264# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X19 X a_83_264# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

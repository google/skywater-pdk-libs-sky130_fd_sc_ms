* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__maj3_4 A B C VGND VNB VPB VPWR X
X0 VPWR a_222_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 a_504_392# B a_222_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X2 VPWR a_222_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 VGND A a_906_78# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 a_222_392# B a_122_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X5 VGND a_222_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VPWR A a_908_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X7 a_222_392# B a_114_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_222_392# B a_504_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X9 VPWR A a_122_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X10 a_908_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X11 a_504_125# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X12 X a_222_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_114_125# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X14 a_504_392# C VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X15 X a_222_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 VPWR C a_504_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X17 X a_222_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X18 a_906_78# C a_222_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X19 a_222_392# C a_906_78# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X20 a_122_392# B a_222_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X21 VGND a_222_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 X a_222_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X23 VGND A a_114_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X24 a_122_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X25 a_908_392# C a_222_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X26 VGND C a_504_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X27 a_114_125# B a_222_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X28 a_222_392# C a_908_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X29 a_222_392# B a_504_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X30 a_504_125# B a_222_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X31 a_906_78# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends

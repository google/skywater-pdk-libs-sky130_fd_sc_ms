* File: sky130_fd_sc_ms__fah_2.spice
* Created: Fri Aug 28 17:35:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__fah_2.pex.spice"
.subckt sky130_fd_sc_ms__fah_2  VNB VPB A B CI VPWR COUT SUM VGND
* 
* VGND	VGND
* SUM	SUM
* COUT	COUT
* VPWR	VPWR
* CI	CI
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1034 N_A_117_368#_M1034_d N_A_81_260#_M1034_g N_VGND_M1034_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1961 AS=0.222 PD=2.01 PS=2.08 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_A_M1012_g N_A_81_260#_M1012_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.2272 PD=0.92 PS=1.99 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75000.3
+ SB=75003.8 A=0.096 P=1.58 MULT=1
MM1000 N_A_416_392#_M1000_d N_A_M1000_g N_VGND_M1012_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.7
+ SB=75003.3 A=0.096 P=1.58 MULT=1
MM1003 N_A_517_424#_M1003_d N_B_M1003_g N_A_416_392#_M1000_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1952 AS=0.0896 PD=1.25 PS=0.92 NRD=61.872 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1005 N_A_117_368#_M1005_d N_A_481_379#_M1005_g N_A_517_424#_M1003_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.272 AS=0.1952 PD=1.49 PS=1.25 NRD=76.872 NRS=0 M=1
+ R=4.26667 SA=75001.9 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1004 N_A_852_424#_M1004_d N_B_M1004_g N_A_117_368#_M1005_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.2224 AS=0.272 PD=1.335 PS=1.49 NRD=50.616 NRS=29.988 M=1 R=4.26667
+ SA=75002.9 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1027 N_A_416_392#_M1027_d N_A_481_379#_M1027_g N_A_852_424#_M1004_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.2455 AS=0.2224 PD=2.38 PS=1.335 NRD=49.68 NRS=27.18 M=1
+ R=4.26667 SA=75003.7 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1033 N_A_481_379#_M1033_d N_B_M1033_g N_VGND_M1033_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.124942 AS=0.31405 PD=1.14217 PS=2.87 NRD=0 NRS=66.48 M=1 R=4.93333
+ SA=75000.3 SB=75004 A=0.111 P=1.78 MULT=1
MM1013 N_A_1454_424#_M1013_d N_A_852_424#_M1013_g N_A_481_379#_M1033_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.28 AS=0.108058 PD=1.515 PS=0.987826 NRD=88.116
+ NRS=8.436 M=1 R=4.26667 SA=75000.8 SB=75004.1 A=0.096 P=1.58 MULT=1
MM1015 N_A_1692_424#_M1015_d N_A_517_424#_M1015_g N_A_1454_424#_M1013_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.2176 AS=0.28 PD=1.32 PS=1.515 NRD=13.116 NRS=23.436
+ M=1 R=4.26667 SA=75001.9 SB=75003.1 A=0.096 P=1.58 MULT=1
MM1008 N_A_1898_424#_M1008_d N_A_852_424#_M1008_g N_A_1692_424#_M1015_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.23645 AS=0.2176 PD=1.45 PS=1.32 NRD=15.936
+ NRS=61.872 M=1 R=4.26667 SA=75002.7 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1028 N_A_2055_424#_M1028_d N_A_517_424#_M1028_g N_A_1898_424#_M1008_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.1344 AS=0.23645 PD=1.06 PS=1.45 NRD=1.872 NRS=60.936
+ M=1 R=4.26667 SA=75003.5 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1010 N_VGND_M1010_d N_A_1692_424#_M1010_g N_A_2055_424#_M1028_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1826 AS=0.1344 PD=1.32 PS=1.06 NRD=43.176 NRS=7.02 M=1
+ R=4.26667 SA=75004.1 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1017 N_A_1692_424#_M1017_d N_CI_M1017_g N_VGND_M1010_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.176 AS=0.1826 PD=1.83 PS=1.32 NRD=0 NRS=43.176 M=1 R=4.26667
+ SA=75004.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1011 N_COUT_M1011_d N_A_1454_424#_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2739 PD=1.02 PS=2.27 NRD=0 NRS=12.972 M=1 R=4.93333
+ SA=75000.3 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1035 N_COUT_M1011_d N_A_1454_424#_M1035_g N_VGND_M1035_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1035_s N_A_1898_424#_M1018_g N_SUM_M1018_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1073 PD=1.09 PS=1.03 NRD=11.34 NRS=0.804 M=1 R=4.93333
+ SA=75001.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1031 N_VGND_M1031_d N_A_1898_424#_M1031_g N_SUM_M1018_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1073 PD=2.05 PS=1.03 NRD=0 NRS=0.804 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1024 N_A_117_368#_M1024_d N_A_81_260#_M1024_g N_VPWR_M1024_s VPB PSHORT L=0.18
+ W=1.12 AD=0.2968 AS=0.3024 PD=2.77 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1029 N_VPWR_M1029_d N_A_M1029_g N_A_81_260#_M1029_s VPB PSHORT L=0.18 W=1
+ AD=0.165 AS=0.27 PD=1.33 PS=2.54 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90003.8 A=0.18 P=2.36 MULT=1
MM1019 N_A_416_392#_M1019_d N_A_M1019_g N_VPWR_M1029_d VPB PSHORT L=0.18 W=1
+ AD=0.170109 AS=0.165 PD=1.44022 PS=1.33 NRD=0 NRS=10.8153 M=1 R=5.55556
+ SA=90000.7 SB=90003.3 A=0.18 P=2.36 MULT=1
MM1030 N_A_517_424#_M1030_d N_A_481_379#_M1030_g N_A_416_392#_M1019_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.3717 AS=0.142891 PD=1.725 PS=1.20978 NRD=0 NRS=10.5395 M=1
+ R=4.66667 SA=90001.2 SB=90003.3 A=0.1512 P=2.04 MULT=1
MM1032 N_A_117_368#_M1032_d N_B_M1032_g N_A_517_424#_M1030_d VPB PSHORT L=0.18
+ W=0.84 AD=0.1806 AS=0.3717 PD=1.27 PS=1.725 NRD=17.5724 NRS=10.5395 M=1
+ R=4.66667 SA=90002.3 SB=90002.3 A=0.1512 P=2.04 MULT=1
MM1002 N_A_852_424#_M1002_d N_A_481_379#_M1002_g N_A_117_368#_M1032_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.5523 AS=0.1806 PD=2.155 PS=1.27 NRD=10.5395 NRS=17.5724 M=1
+ R=4.66667 SA=90002.9 SB=90001.7 A=0.1512 P=2.04 MULT=1
MM1014 N_A_416_392#_M1014_d N_B_M1014_g N_A_852_424#_M1002_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2268 AS=0.5523 PD=2.22 PS=2.155 NRD=0 NRS=90.2851 M=1 R=4.66667
+ SA=90004.4 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1025 N_A_481_379#_M1025_d N_B_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2088 AS=0.3024 PD=1.67429 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003.8 A=0.2016 P=2.6 MULT=1
MM1021 N_A_1454_424#_M1021_d N_A_517_424#_M1021_g N_A_481_379#_M1025_d VPB
+ PSHORT L=0.18 W=0.84 AD=0.4242 AS=0.1566 PD=1.85 PS=1.25571 NRD=72.693
+ NRS=30.8108 M=1 R=4.66667 SA=90000.7 SB=90004.5 A=0.1512 P=2.04 MULT=1
MM1026 N_A_1692_424#_M1026_d N_A_852_424#_M1026_g N_A_1454_424#_M1021_d VPB
+ PSHORT L=0.18 W=0.84 AD=0.357 AS=0.4242 PD=1.69 PS=1.85 NRD=110.222 NRS=0 M=1
+ R=4.66667 SA=90001.9 SB=90003.3 A=0.1512 P=2.04 MULT=1
MM1016 N_A_1898_424#_M1016_d N_A_517_424#_M1016_g N_A_1692_424#_M1026_d VPB
+ PSHORT L=0.18 W=0.84 AD=0.2541 AS=0.357 PD=1.445 PS=1.69 NRD=65.6601
+ NRS=23.443 M=1 R=4.66667 SA=90002.9 SB=90002.3 A=0.1512 P=2.04 MULT=1
MM1022 N_A_2055_424#_M1022_d N_A_852_424#_M1022_g N_A_1898_424#_M1016_d VPB
+ PSHORT L=0.18 W=0.84 AD=0.211917 AS=0.2541 PD=1.37413 PS=1.445 NRD=18.7544
+ NRS=10.5395 M=1 R=4.66667 SA=90003.7 SB=90001.5 A=0.1512 P=2.04 MULT=1
MM1020 N_VPWR_M1020_d N_A_1692_424#_M1020_g N_A_2055_424#_M1022_d VPB PSHORT
+ L=0.18 W=1 AD=0.2807 AS=0.252283 PD=1.7 PS=1.63587 NRD=44.4432 NRS=8.8453 M=1
+ R=5.55556 SA=90003.7 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1023 N_A_1692_424#_M1023_d N_CI_M1023_g N_VPWR_M1020_d VPB PSHORT L=0.18 W=1
+ AD=0.27 AS=0.2807 PD=2.54 PS=1.7 NRD=0 NRS=44.4432 M=1 R=5.55556 SA=90004.4
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1001 N_COUT_M1001_d N_A_1454_424#_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2862 PD=1.39 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1006 N_COUT_M1001_d N_A_1454_424#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1007 N_VPWR_M1006_s N_A_1898_424#_M1007_g N_SUM_M1007_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1568 PD=1.39 PS=1.4 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1009 N_VPWR_M1009_d N_A_1898_424#_M1009_g N_SUM_M1007_s VPB PSHORT L=0.18
+ W=1.12 AD=0.3192 AS=0.1568 PD=2.81 PS=1.4 NRD=1.7533 NRS=0 M=1 R=6.22222
+ SA=90001.5 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX36_noxref VNB VPB NWDIODE A=27.4908 P=33.28
c_152 VNB 0 7.1893e-20 $X=0 $Y=0
c_262 VPB 0 5.30342e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__fah_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__and3_2.pxi.spice
* Created: Wed Sep  2 11:57:44 2020
* 
x_PM_SKY130_FD_SC_MS__AND3_2%A N_A_c_57_n N_A_M1006_g N_A_c_59_n N_A_M1005_g A A
+ A N_A_c_62_n PM_SKY130_FD_SC_MS__AND3_2%A
x_PM_SKY130_FD_SC_MS__AND3_2%B N_B_M1007_g N_B_M1004_g B B N_B_c_92_n N_B_c_93_n
+ PM_SKY130_FD_SC_MS__AND3_2%B
x_PM_SKY130_FD_SC_MS__AND3_2%C N_C_M1003_g N_C_M1008_g C N_C_c_129_n N_C_c_130_n
+ PM_SKY130_FD_SC_MS__AND3_2%C
x_PM_SKY130_FD_SC_MS__AND3_2%A_41_384# N_A_41_384#_M1005_s N_A_41_384#_M1006_s
+ N_A_41_384#_M1007_d N_A_41_384#_M1000_g N_A_41_384#_M1001_g
+ N_A_41_384#_M1009_g N_A_41_384#_M1002_g N_A_41_384#_c_168_n
+ N_A_41_384#_c_182_n N_A_41_384#_c_202_n N_A_41_384#_c_175_n
+ N_A_41_384#_c_169_n N_A_41_384#_c_176_n N_A_41_384#_c_177_n
+ N_A_41_384#_c_170_n N_A_41_384#_c_171_n PM_SKY130_FD_SC_MS__AND3_2%A_41_384#
x_PM_SKY130_FD_SC_MS__AND3_2%VPWR N_VPWR_M1006_d N_VPWR_M1008_d N_VPWR_M1002_s
+ N_VPWR_c_262_n N_VPWR_c_263_n N_VPWR_c_264_n N_VPWR_c_265_n N_VPWR_c_266_n
+ N_VPWR_c_267_n VPWR N_VPWR_c_268_n N_VPWR_c_269_n N_VPWR_c_261_n
+ PM_SKY130_FD_SC_MS__AND3_2%VPWR
x_PM_SKY130_FD_SC_MS__AND3_2%X N_X_M1000_d N_X_M1001_d N_X_c_304_n N_X_c_307_n
+ N_X_c_308_n N_X_c_305_n X PM_SKY130_FD_SC_MS__AND3_2%X
x_PM_SKY130_FD_SC_MS__AND3_2%VGND N_VGND_M1003_d N_VGND_M1009_s N_VGND_c_345_n
+ N_VGND_c_346_n N_VGND_c_347_n VGND N_VGND_c_348_n N_VGND_c_349_n
+ N_VGND_c_350_n N_VGND_c_351_n PM_SKY130_FD_SC_MS__AND3_2%VGND
cc_1 VNB N_A_c_57_n 0.00691804f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.485
cc_2 VNB N_A_M1006_g 0.0113576f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.34
cc_3 VNB N_A_c_59_n 0.0324727f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.57
cc_4 VNB N_A_M1005_g 0.0117117f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1
cc_5 VNB A 0.045212f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=0.47
cc_6 VNB N_A_c_62_n 0.0476697f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.405
cc_7 VNB B 0.0034927f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1
cc_8 VNB N_B_c_92_n 0.0199635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B_c_93_n 0.0152038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB C 0.00354858f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1
cc_11 VNB N_C_c_129_n 0.0217853f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_12 VNB N_C_c_130_n 0.0185142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_41_384#_M1000_g 0.0222518f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=0.47
cc_14 VNB N_A_41_384#_M1009_g 0.0231292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_41_384#_c_168_n 0.0137129f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.462
cc_16 VNB N_A_41_384#_c_169_n 0.0199411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_41_384#_c_170_n 0.00344604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_41_384#_c_171_n 0.0587856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_261_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_X_c_304_n 0.00296545f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.395
cc_21 VNB N_X_c_305_n 0.00598001f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.405
cc_22 VNB X 0.00379924f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_345_n 0.0199076f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.395
cc_24 VNB N_VGND_c_346_n 0.0451591f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_25 VNB N_VGND_c_347_n 0.0275707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_348_n 0.0441425f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=0.405
cc_27 VNB N_VGND_c_349_n 0.0188369f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.405
cc_28 VNB N_VGND_c_350_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.462
cc_29 VNB N_VGND_c_351_n 0.214004f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VPB N_A_M1006_g 0.0344283f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=2.34
cc_31 VPB N_B_M1007_g 0.022585f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=2.34
cc_32 VPB B 0.00303485f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1
cc_33 VPB N_B_c_92_n 0.0107152f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_C_M1008_g 0.0237731f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.395
cc_35 VPB C 0.00165062f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1
cc_36 VPB N_C_c_129_n 0.0122147f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=0.47
cc_37 VPB N_A_41_384#_M1001_g 0.0237842f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=0.405
cc_38 VPB N_A_41_384#_M1002_g 0.0265313f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.462
cc_39 VPB N_A_41_384#_c_168_n 0.0119354f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.462
cc_40 VPB N_A_41_384#_c_175_n 0.00271444f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_A_41_384#_c_176_n 0.0356746f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A_41_384#_c_177_n 0.00318593f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A_41_384#_c_171_n 0.00931597f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_262_n 0.0268219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_263_n 0.0173426f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.405
cc_46 VPB N_VPWR_c_264_n 0.0128289f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_265_n 0.063207f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=0.405
cc_48 VPB N_VPWR_c_266_n 0.025575f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.462
cc_49 VPB N_VPWR_c_267_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=0.462
cc_50 VPB N_VPWR_c_268_n 0.019175f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_269_n 0.0285346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_261_n 0.0784136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_X_c_307_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_X_c_308_n 0.00103829f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.405
cc_55 VPB N_X_c_305_n 0.00128906f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=0.405
cc_56 N_A_M1006_g N_B_M1007_g 0.0247281f $X=0.575 $Y=2.34 $X2=0 $Y2=0
cc_57 N_A_c_57_n B 0.00119477f $X=0.575 $Y=1.485 $X2=0 $Y2=0
cc_58 N_A_M1005_g B 0.00223423f $X=0.59 $Y=1 $X2=0 $Y2=0
cc_59 A B 0.01291f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_60 N_A_c_57_n N_B_c_92_n 0.0168712f $X=0.575 $Y=1.485 $X2=0 $Y2=0
cc_61 N_A_c_59_n N_B_c_93_n 8.67721e-19 $X=0.59 $Y=0.57 $X2=0 $Y2=0
cc_62 N_A_M1005_g N_B_c_93_n 0.0245557f $X=0.59 $Y=1 $X2=0 $Y2=0
cc_63 A N_B_c_93_n 0.0109386f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_64 A N_C_c_130_n 0.00108821f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_65 N_A_c_57_n N_A_41_384#_c_168_n 0.00393408f $X=0.575 $Y=1.485 $X2=0 $Y2=0
cc_66 N_A_M1006_g N_A_41_384#_c_168_n 0.0169565f $X=0.575 $Y=2.34 $X2=0 $Y2=0
cc_67 N_A_M1005_g N_A_41_384#_c_168_n 0.0015053f $X=0.59 $Y=1 $X2=0 $Y2=0
cc_68 N_A_M1006_g N_A_41_384#_c_182_n 0.0176738f $X=0.575 $Y=2.34 $X2=0 $Y2=0
cc_69 N_A_M1005_g N_A_41_384#_c_169_n 0.012609f $X=0.59 $Y=1 $X2=0 $Y2=0
cc_70 A N_A_41_384#_c_169_n 0.0277772f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_71 N_A_c_62_n N_A_41_384#_c_169_n 0.00188139f $X=0.515 $Y=0.405 $X2=0 $Y2=0
cc_72 N_A_M1006_g N_A_41_384#_c_176_n 0.0136089f $X=0.575 $Y=2.34 $X2=0 $Y2=0
cc_73 N_A_M1006_g N_A_41_384#_c_177_n 8.07074e-19 $X=0.575 $Y=2.34 $X2=0 $Y2=0
cc_74 N_A_M1006_g N_VPWR_c_262_n 0.00418809f $X=0.575 $Y=2.34 $X2=0 $Y2=0
cc_75 N_A_M1006_g N_VPWR_c_269_n 0.00513676f $X=0.575 $Y=2.34 $X2=0 $Y2=0
cc_76 N_A_M1006_g N_VPWR_c_261_n 0.00581878f $X=0.575 $Y=2.34 $X2=0 $Y2=0
cc_77 A N_VGND_c_345_n 0.0214717f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_78 A N_VGND_c_348_n 0.0794507f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_79 N_A_c_62_n N_VGND_c_348_n 0.0116176f $X=0.515 $Y=0.405 $X2=0 $Y2=0
cc_80 N_A_c_59_n N_VGND_c_351_n 0.00642106f $X=0.59 $Y=0.57 $X2=0 $Y2=0
cc_81 A N_VGND_c_351_n 0.0425626f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_82 N_A_c_62_n N_VGND_c_351_n 0.00862283f $X=0.515 $Y=0.405 $X2=0 $Y2=0
cc_83 N_B_M1007_g N_C_M1008_g 0.0197f $X=1.145 $Y=2.34 $X2=0 $Y2=0
cc_84 B C 0.0282664f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_85 N_B_c_92_n C 3.52745e-19 $X=1.07 $Y=1.595 $X2=0 $Y2=0
cc_86 N_B_c_92_n N_C_c_129_n 0.0316904f $X=1.07 $Y=1.595 $X2=0 $Y2=0
cc_87 B N_C_c_130_n 0.00818659f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_88 N_B_c_93_n N_C_c_130_n 0.0316904f $X=1.07 $Y=1.43 $X2=0 $Y2=0
cc_89 N_B_M1007_g N_A_41_384#_c_168_n 7.8694e-19 $X=1.145 $Y=2.34 $X2=0 $Y2=0
cc_90 B N_A_41_384#_c_168_n 0.017863f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_91 N_B_c_92_n N_A_41_384#_c_168_n 9.66961e-19 $X=1.07 $Y=1.595 $X2=0 $Y2=0
cc_92 N_B_M1007_g N_A_41_384#_c_182_n 0.0135147f $X=1.145 $Y=2.34 $X2=0 $Y2=0
cc_93 B N_A_41_384#_c_182_n 0.0214504f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_94 N_B_c_92_n N_A_41_384#_c_182_n 8.71992e-19 $X=1.07 $Y=1.595 $X2=0 $Y2=0
cc_95 B N_A_41_384#_c_169_n 0.00709791f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_96 N_B_c_93_n N_A_41_384#_c_169_n 0.0016883f $X=1.07 $Y=1.43 $X2=0 $Y2=0
cc_97 N_B_M1007_g N_A_41_384#_c_176_n 8.68654e-19 $X=1.145 $Y=2.34 $X2=0 $Y2=0
cc_98 N_B_M1007_g N_A_41_384#_c_177_n 0.0121207f $X=1.145 $Y=2.34 $X2=0 $Y2=0
cc_99 B N_A_41_384#_c_177_n 0.00709708f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_100 N_B_M1007_g N_VPWR_c_262_n 0.00623981f $X=1.145 $Y=2.34 $X2=0 $Y2=0
cc_101 N_B_M1007_g N_VPWR_c_266_n 0.00513676f $X=1.145 $Y=2.34 $X2=0 $Y2=0
cc_102 N_B_M1007_g N_VPWR_c_261_n 0.00581878f $X=1.145 $Y=2.34 $X2=0 $Y2=0
cc_103 B A_133_136# 0.00402475f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_104 B A_247_136# 0.00221309f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_105 N_B_c_93_n N_VGND_c_348_n 4.78105e-19 $X=1.07 $Y=1.43 $X2=0 $Y2=0
cc_106 N_C_c_130_n N_A_41_384#_M1000_g 0.0193095f $X=1.645 $Y=1.43 $X2=0 $Y2=0
cc_107 N_C_M1008_g N_A_41_384#_M1001_g 0.0123621f $X=1.595 $Y=2.34 $X2=0 $Y2=0
cc_108 N_C_c_129_n N_A_41_384#_M1001_g 0.00197523f $X=1.65 $Y=1.595 $X2=0 $Y2=0
cc_109 N_C_M1008_g N_A_41_384#_c_202_n 0.013956f $X=1.595 $Y=2.34 $X2=0 $Y2=0
cc_110 C N_A_41_384#_c_202_n 0.0188573f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_111 N_C_c_129_n N_A_41_384#_c_202_n 7.38901e-19 $X=1.65 $Y=1.595 $X2=0 $Y2=0
cc_112 N_C_M1008_g N_A_41_384#_c_175_n 0.00322666f $X=1.595 $Y=2.34 $X2=0 $Y2=0
cc_113 C N_A_41_384#_c_175_n 0.00689942f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_114 N_C_c_129_n N_A_41_384#_c_175_n 6.86462e-19 $X=1.65 $Y=1.595 $X2=0 $Y2=0
cc_115 N_C_M1008_g N_A_41_384#_c_177_n 0.0143622f $X=1.595 $Y=2.34 $X2=0 $Y2=0
cc_116 C N_A_41_384#_c_177_n 0.00318067f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_117 C N_A_41_384#_c_170_n 0.0157355f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_118 N_C_c_129_n N_A_41_384#_c_170_n 0.00147149f $X=1.65 $Y=1.595 $X2=0 $Y2=0
cc_119 N_C_c_130_n N_A_41_384#_c_170_n 0.00169384f $X=1.645 $Y=1.43 $X2=0 $Y2=0
cc_120 C N_A_41_384#_c_171_n 2.91011e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_121 N_C_c_129_n N_A_41_384#_c_171_n 0.0128568f $X=1.65 $Y=1.595 $X2=0 $Y2=0
cc_122 N_C_M1008_g N_VPWR_c_263_n 0.00794432f $X=1.595 $Y=2.34 $X2=0 $Y2=0
cc_123 N_C_M1008_g N_VPWR_c_266_n 0.00513676f $X=1.595 $Y=2.34 $X2=0 $Y2=0
cc_124 N_C_M1008_g N_VPWR_c_261_n 0.00581878f $X=1.595 $Y=2.34 $X2=0 $Y2=0
cc_125 N_C_M1008_g N_X_c_307_n 8.03947e-19 $X=1.595 $Y=2.34 $X2=0 $Y2=0
cc_126 C N_VGND_c_345_n 0.00794902f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_127 N_C_c_129_n N_VGND_c_345_n 9.9563e-19 $X=1.65 $Y=1.595 $X2=0 $Y2=0
cc_128 N_C_c_130_n N_VGND_c_345_n 0.0047463f $X=1.645 $Y=1.43 $X2=0 $Y2=0
cc_129 N_C_c_130_n N_VGND_c_348_n 0.0038748f $X=1.645 $Y=1.43 $X2=0 $Y2=0
cc_130 N_C_c_130_n N_VGND_c_351_n 0.00454494f $X=1.645 $Y=1.43 $X2=0 $Y2=0
cc_131 N_A_41_384#_c_182_n N_VPWR_M1006_d 0.0110071f $X=1.205 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_132 N_A_41_384#_c_202_n N_VPWR_M1008_d 0.0200575f $X=2.035 $Y=2.035 $X2=0
+ $Y2=0
cc_133 N_A_41_384#_c_175_n N_VPWR_M1008_d 0.00219679f $X=2.12 $Y=1.95 $X2=0
+ $Y2=0
cc_134 N_A_41_384#_c_182_n N_VPWR_c_262_n 0.022455f $X=1.205 $Y=2.035 $X2=0
+ $Y2=0
cc_135 N_A_41_384#_c_176_n N_VPWR_c_262_n 0.0191764f $X=0.35 $Y=2.065 $X2=0
+ $Y2=0
cc_136 N_A_41_384#_c_177_n N_VPWR_c_262_n 0.0175494f $X=1.37 $Y=2.115 $X2=0
+ $Y2=0
cc_137 N_A_41_384#_M1001_g N_VPWR_c_263_n 0.00534567f $X=2.315 $Y=2.4 $X2=0
+ $Y2=0
cc_138 N_A_41_384#_c_202_n N_VPWR_c_263_n 0.0244925f $X=2.035 $Y=2.035 $X2=0
+ $Y2=0
cc_139 N_A_41_384#_c_177_n N_VPWR_c_263_n 0.0223815f $X=1.37 $Y=2.115 $X2=0
+ $Y2=0
cc_140 N_A_41_384#_c_171_n N_VPWR_c_263_n 4.25493e-19 $X=2.765 $Y=1.505 $X2=0
+ $Y2=0
cc_141 N_A_41_384#_M1002_g N_VPWR_c_265_n 0.0284321f $X=2.765 $Y=2.4 $X2=0 $Y2=0
cc_142 N_A_41_384#_c_177_n N_VPWR_c_266_n 0.00787326f $X=1.37 $Y=2.115 $X2=0
+ $Y2=0
cc_143 N_A_41_384#_M1001_g N_VPWR_c_268_n 0.005209f $X=2.315 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A_41_384#_M1002_g N_VPWR_c_268_n 0.0049824f $X=2.765 $Y=2.4 $X2=0 $Y2=0
cc_145 N_A_41_384#_c_176_n N_VPWR_c_269_n 0.00794361f $X=0.35 $Y=2.065 $X2=0
+ $Y2=0
cc_146 N_A_41_384#_M1001_g N_VPWR_c_261_n 0.00986727f $X=2.315 $Y=2.4 $X2=0
+ $Y2=0
cc_147 N_A_41_384#_M1002_g N_VPWR_c_261_n 0.00912684f $X=2.765 $Y=2.4 $X2=0
+ $Y2=0
cc_148 N_A_41_384#_c_176_n N_VPWR_c_261_n 0.0105573f $X=0.35 $Y=2.065 $X2=0
+ $Y2=0
cc_149 N_A_41_384#_c_177_n N_VPWR_c_261_n 0.0105247f $X=1.37 $Y=2.115 $X2=0
+ $Y2=0
cc_150 N_A_41_384#_M1000_g N_X_c_304_n 0.00562723f $X=2.13 $Y=0.78 $X2=0 $Y2=0
cc_151 N_A_41_384#_M1009_g N_X_c_304_n 4.72567e-19 $X=2.6 $Y=0.78 $X2=0 $Y2=0
cc_152 N_A_41_384#_M1001_g N_X_c_307_n 0.013985f $X=2.315 $Y=2.4 $X2=0 $Y2=0
cc_153 N_A_41_384#_M1002_g N_X_c_307_n 0.0137155f $X=2.765 $Y=2.4 $X2=0 $Y2=0
cc_154 N_A_41_384#_M1001_g N_X_c_308_n 0.0026301f $X=2.315 $Y=2.4 $X2=0 $Y2=0
cc_155 N_A_41_384#_M1002_g N_X_c_308_n 0.0022984f $X=2.765 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A_41_384#_c_170_n N_X_c_308_n 7.18422e-19 $X=2.22 $Y=1.505 $X2=0 $Y2=0
cc_157 N_A_41_384#_c_171_n N_X_c_308_n 0.00204723f $X=2.765 $Y=1.505 $X2=0 $Y2=0
cc_158 N_A_41_384#_M1000_g N_X_c_305_n 9.76257e-19 $X=2.13 $Y=0.78 $X2=0 $Y2=0
cc_159 N_A_41_384#_M1001_g N_X_c_305_n 0.00132552f $X=2.315 $Y=2.4 $X2=0 $Y2=0
cc_160 N_A_41_384#_M1009_g N_X_c_305_n 0.00712292f $X=2.6 $Y=0.78 $X2=0 $Y2=0
cc_161 N_A_41_384#_M1002_g N_X_c_305_n 0.00769885f $X=2.765 $Y=2.4 $X2=0 $Y2=0
cc_162 N_A_41_384#_c_175_n N_X_c_305_n 0.0076953f $X=2.12 $Y=1.95 $X2=0 $Y2=0
cc_163 N_A_41_384#_c_170_n N_X_c_305_n 0.0236573f $X=2.22 $Y=1.505 $X2=0 $Y2=0
cc_164 N_A_41_384#_c_171_n N_X_c_305_n 0.0238914f $X=2.765 $Y=1.505 $X2=0 $Y2=0
cc_165 N_A_41_384#_M1000_g X 0.00442604f $X=2.13 $Y=0.78 $X2=0 $Y2=0
cc_166 N_A_41_384#_M1009_g X 0.0156684f $X=2.6 $Y=0.78 $X2=0 $Y2=0
cc_167 N_A_41_384#_c_170_n X 0.0162347f $X=2.22 $Y=1.505 $X2=0 $Y2=0
cc_168 N_A_41_384#_c_171_n X 0.00566308f $X=2.765 $Y=1.505 $X2=0 $Y2=0
cc_169 N_A_41_384#_M1000_g N_VGND_c_345_n 0.010364f $X=2.13 $Y=0.78 $X2=0 $Y2=0
cc_170 N_A_41_384#_M1009_g N_VGND_c_346_n 0.00878267f $X=2.6 $Y=0.78 $X2=0 $Y2=0
cc_171 N_A_41_384#_c_171_n N_VGND_c_346_n 0.00283438f $X=2.765 $Y=1.505 $X2=0
+ $Y2=0
cc_172 N_A_41_384#_M1009_g N_VGND_c_347_n 0.00565998f $X=2.6 $Y=0.78 $X2=0 $Y2=0
cc_173 N_A_41_384#_M1000_g N_VGND_c_349_n 0.00523933f $X=2.13 $Y=0.78 $X2=0
+ $Y2=0
cc_174 N_A_41_384#_M1009_g N_VGND_c_349_n 0.00548708f $X=2.6 $Y=0.78 $X2=0 $Y2=0
cc_175 N_A_41_384#_M1000_g N_VGND_c_351_n 0.00533081f $X=2.13 $Y=0.78 $X2=0
+ $Y2=0
cc_176 N_A_41_384#_M1009_g N_VGND_c_351_n 0.00533081f $X=2.6 $Y=0.78 $X2=0 $Y2=0
cc_177 N_VPWR_c_263_n N_X_c_307_n 0.0269152f $X=2.04 $Y=2.455 $X2=0 $Y2=0
cc_178 N_VPWR_c_268_n N_X_c_307_n 0.0152949f $X=2.895 $Y=3.33 $X2=0 $Y2=0
cc_179 N_VPWR_c_261_n N_X_c_307_n 0.0124766f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_180 N_VPWR_c_265_n N_X_c_305_n 0.0453496f $X=3.06 $Y=1.985 $X2=0 $Y2=0
cc_181 N_VPWR_c_265_n N_VGND_c_347_n 0.0108898f $X=3.06 $Y=1.985 $X2=0 $Y2=0
cc_182 X N_VGND_M1009_s 0.00398771f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_183 N_X_c_304_n N_VGND_c_345_n 0.0165499f $X=2.345 $Y=0.555 $X2=0 $Y2=0
cc_184 X N_VGND_c_345_n 0.0154525f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_185 N_X_c_304_n N_VGND_c_346_n 0.0016552f $X=2.345 $Y=0.555 $X2=0 $Y2=0
cc_186 X N_VGND_c_346_n 0.00191947f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_187 X N_VGND_c_347_n 0.0300887f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_188 N_X_c_304_n N_VGND_c_349_n 0.0121172f $X=2.345 $Y=0.555 $X2=0 $Y2=0
cc_189 N_X_c_304_n N_VGND_c_351_n 0.0115967f $X=2.345 $Y=0.555 $X2=0 $Y2=0
cc_190 X N_VGND_c_351_n 0.00618074f $X=2.555 $Y=0.84 $X2=0 $Y2=0

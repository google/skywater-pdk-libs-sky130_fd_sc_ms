* File: sky130_fd_sc_ms__o41a_1.spice
* Created: Fri Aug 28 18:04:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o41a_1.pex.spice"
.subckt sky130_fd_sc_ms__o41a_1  VNB VPB B1 A4 A3 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A_83_270#_M1010_g N_X_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.2109 PD=2.19 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1004 N_A_326_74#_M1004_d N_B1_M1004_g N_A_83_270#_M1004_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.112 AS=0.1824 PD=0.99 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1001_d N_A4_M1001_g N_A_326_74#_M1004_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1344 AS=0.112 PD=1.06 PS=0.99 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75000.7
+ SB=75002 A=0.096 P=1.58 MULT=1
MM1011 N_A_326_74#_M1011_d N_A3_M1011_g N_VGND_M1001_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1088 AS=0.1344 PD=0.98 PS=1.06 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75001.3
+ SB=75001.4 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g N_A_326_74#_M1011_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1792 AS=0.1088 PD=1.2 PS=0.98 NRD=20.616 NRS=11.244 M=1 R=4.26667
+ SA=75001.8 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1008 N_A_326_74#_M1008_d N_A1_M1008_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.1792 PD=1.85 PS=1.2 NRD=0 NRS=31.872 M=1 R=4.26667 SA=75002.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_A_83_270#_M1000_g N_X_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.521714 AS=0.3136 PD=2.33143 PS=2.8 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90002.7 A=0.2016 P=2.6 MULT=1
MM1002 N_A_83_270#_M1002_d N_B1_M1002_g N_VPWR_M1000_d VPB PSHORT L=0.18 W=0.84
+ AD=0.159536 AS=0.391286 PD=1.26429 PS=1.74857 NRD=18.7544 NRS=19.9167 M=1
+ R=4.66667 SA=90001.3 SB=90002.4 A=0.1512 P=2.04 MULT=1
MM1003 A_446_368# N_A4_M1003_g N_A_83_270#_M1002_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1344 AS=0.212714 PD=1.36 PS=1.68571 NRD=11.426 NRS=0 M=1 R=6.22222
+ SA=90001.4 SB=90001.9 A=0.2016 P=2.6 MULT=1
MM1007 A_530_368# N_A3_M1007_g A_446_368# VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.1344 PD=1.51 PS=1.36 NRD=24.6053 NRS=11.426 M=1 R=6.22222 SA=90001.8
+ SB=90001.4 A=0.2016 P=2.6 MULT=1
MM1005 A_644_368# N_A2_M1005_g A_530_368# VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.2184 PD=1.51 PS=1.51 NRD=24.6053 NRS=24.6053 M=1 R=6.22222 SA=90002.4
+ SB=90000.9 A=0.2016 P=2.6 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g A_644_368# VPB PSHORT L=0.18 W=1.12 AD=0.4424
+ AS=0.2184 PD=3.03 PS=1.51 NRD=0 NRS=24.6053 M=1 R=6.22222 SA=90003 SB=90000.3
+ A=0.2016 P=2.6 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__o41a_1.pxi.spice"
*
.ends
*
*

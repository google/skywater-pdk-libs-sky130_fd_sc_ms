* File: sky130_fd_sc_ms__einvp_4.pxi.spice
* Created: Fri Aug 28 17:34:16 2020
* 
x_PM_SKY130_FD_SC_MS__EINVP_4%A N_A_M1007_g N_A_M1000_g N_A_M1002_g N_A_M1009_g
+ N_A_M1003_g N_A_M1013_g N_A_c_113_n N_A_M1006_g N_A_M1016_g N_A_c_116_n A A A
+ N_A_c_117_n N_A_c_118_n PM_SKY130_FD_SC_MS__EINVP_4%A
x_PM_SKY130_FD_SC_MS__EINVP_4%A_473_323# N_A_473_323#_M1014_s
+ N_A_473_323#_M1012_s N_A_473_323#_c_210_n N_A_473_323#_M1004_g
+ N_A_473_323#_c_198_n N_A_473_323#_c_199_n N_A_473_323#_c_213_n
+ N_A_473_323#_M1005_g N_A_473_323#_c_200_n N_A_473_323#_c_215_n
+ N_A_473_323#_M1008_g N_A_473_323#_c_201_n N_A_473_323#_c_217_n
+ N_A_473_323#_M1015_g N_A_473_323#_c_202_n N_A_473_323#_c_203_n
+ N_A_473_323#_c_204_n N_A_473_323#_c_205_n N_A_473_323#_c_206_n
+ N_A_473_323#_c_207_n N_A_473_323#_c_222_n N_A_473_323#_c_208_n
+ N_A_473_323#_c_209_n PM_SKY130_FD_SC_MS__EINVP_4%A_473_323#
x_PM_SKY130_FD_SC_MS__EINVP_4%TE N_TE_c_310_n N_TE_M1001_g N_TE_c_311_n
+ N_TE_c_312_n N_TE_c_313_n N_TE_M1010_g N_TE_c_314_n N_TE_c_315_n N_TE_M1011_g
+ N_TE_c_316_n N_TE_c_317_n N_TE_M1017_g N_TE_c_318_n N_TE_M1014_g N_TE_M1012_g
+ N_TE_c_320_n N_TE_c_321_n N_TE_c_322_n TE N_TE_c_324_n N_TE_c_325_n
+ N_TE_c_326_n PM_SKY130_FD_SC_MS__EINVP_4%TE
x_PM_SKY130_FD_SC_MS__EINVP_4%A_27_368# N_A_27_368#_M1000_s N_A_27_368#_M1002_s
+ N_A_27_368#_M1006_s N_A_27_368#_M1005_s N_A_27_368#_M1015_s
+ N_A_27_368#_c_411_n N_A_27_368#_c_412_n N_A_27_368#_c_413_n
+ N_A_27_368#_c_469_p N_A_27_368#_c_414_n N_A_27_368#_c_415_n
+ N_A_27_368#_c_416_n N_A_27_368#_c_410_n N_A_27_368#_c_418_n
+ N_A_27_368#_c_419_n N_A_27_368#_c_420_n N_A_27_368#_c_421_n
+ N_A_27_368#_c_459_n PM_SKY130_FD_SC_MS__EINVP_4%A_27_368#
x_PM_SKY130_FD_SC_MS__EINVP_4%Z N_Z_M1007_s N_Z_M1013_s N_Z_M1000_d N_Z_M1003_d
+ N_Z_c_504_n N_Z_c_499_n N_Z_c_500_n N_Z_c_514_n N_Z_c_518_n N_Z_c_501_n
+ N_Z_c_526_n N_Z_c_530_n N_Z_c_502_n Z PM_SKY130_FD_SC_MS__EINVP_4%Z
x_PM_SKY130_FD_SC_MS__EINVP_4%VPWR N_VPWR_M1004_d N_VPWR_M1008_d N_VPWR_M1012_d
+ N_VPWR_c_558_n N_VPWR_c_559_n N_VPWR_c_560_n N_VPWR_c_561_n VPWR
+ N_VPWR_c_562_n N_VPWR_c_563_n N_VPWR_c_564_n N_VPWR_c_565_n N_VPWR_c_566_n
+ N_VPWR_c_557_n PM_SKY130_FD_SC_MS__EINVP_4%VPWR
x_PM_SKY130_FD_SC_MS__EINVP_4%A_27_74# N_A_27_74#_M1007_d N_A_27_74#_M1009_d
+ N_A_27_74#_M1016_d N_A_27_74#_M1010_s N_A_27_74#_M1017_s N_A_27_74#_c_619_n
+ N_A_27_74#_c_620_n N_A_27_74#_c_621_n N_A_27_74#_c_689_n N_A_27_74#_c_622_n
+ N_A_27_74#_c_623_n N_A_27_74#_c_624_n N_A_27_74#_c_625_n N_A_27_74#_c_626_n
+ N_A_27_74#_c_627_n N_A_27_74#_c_628_n N_A_27_74#_c_629_n N_A_27_74#_c_630_n
+ PM_SKY130_FD_SC_MS__EINVP_4%A_27_74#
x_PM_SKY130_FD_SC_MS__EINVP_4%VGND N_VGND_M1001_d N_VGND_M1011_d N_VGND_M1014_d
+ N_VGND_c_715_n N_VGND_c_716_n N_VGND_c_717_n N_VGND_c_718_n N_VGND_c_719_n
+ N_VGND_c_720_n VGND N_VGND_c_721_n N_VGND_c_722_n N_VGND_c_723_n
+ N_VGND_c_724_n PM_SKY130_FD_SC_MS__EINVP_4%VGND
cc_1 VNB N_A_M1007_g 0.0326264f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_M1009_g 0.0244962f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_3 VNB N_A_M1013_g 0.0240943f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=0.74
cc_4 VNB N_A_c_113_n 0.0109911f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=1.425
cc_5 VNB N_A_M1006_g 0.0114766f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_6 VNB N_A_M1016_g 0.0243622f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=0.74
cc_7 VNB N_A_c_116_n 0.00907757f $X=-0.19 $Y=-0.245 $X2=1.967 $Y2=1.425
cc_8 VNB N_A_c_117_n 0.016914f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_9 VNB N_A_c_118_n 0.0591549f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.515
cc_10 VNB N_A_473_323#_c_198_n 0.00718816f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_11 VNB N_A_473_323#_c_199_n 0.00538699f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_12 VNB N_A_473_323#_c_200_n 0.00607997f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_13 VNB N_A_473_323#_c_201_n 0.00630172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_473_323#_c_202_n 0.0174524f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=1.425
cc_15 VNB N_A_473_323#_c_203_n 0.00413151f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.5
cc_16 VNB N_A_473_323#_c_204_n 0.00413142f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_17 VNB N_A_473_323#_c_205_n 0.00413151f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_18 VNB N_A_473_323#_c_206_n 0.00909917f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=0.74
cc_19 VNB N_A_473_323#_c_207_n 0.00914505f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_20 VNB N_A_473_323#_c_208_n 2.54189e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_473_323#_c_209_n 0.00653231f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=1.515
cc_22 VNB N_TE_c_310_n 0.018325f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_23 VNB N_TE_c_311_n 0.0166678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_TE_c_312_n 0.00643851f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.68
cc_25 VNB N_TE_c_313_n 0.0180464f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_26 VNB N_TE_c_314_n 0.0105119f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.68
cc_27 VNB N_TE_c_315_n 0.0180464f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_28 VNB N_TE_c_316_n 0.0166678f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_29 VNB N_TE_c_317_n 0.0232894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_TE_c_318_n 0.0245033f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.35
cc_31 VNB N_TE_M1012_g 0.00265685f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.425
cc_32 VNB N_TE_c_320_n 0.00411221f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_33 VNB N_TE_c_321_n 0.00411221f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_34 VNB N_TE_c_322_n 0.00411221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB TE 0.0246417f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=0.74
cc_36 VNB N_TE_c_324_n 0.0497754f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_37 VNB N_TE_c_325_n 0.0768529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_TE_c_326_n 0.00245723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_368#_c_410_n 0.00443147f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_40 VNB N_Z_c_499_n 0.00388917f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=2.4
cc_41 VNB N_Z_c_500_n 0.00320239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_Z_c_501_n 0.00363957f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_43 VNB N_Z_c_502_n 9.85474e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VPWR_c_557_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_45 VNB N_A_27_74#_c_619_n 0.0302158f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=2.4
cc_46 VNB N_A_27_74#_c_620_n 0.00280532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_27_74#_c_621_n 0.00971634f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.35
cc_48 VNB N_A_27_74#_c_622_n 0.00484762f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.425
cc_49 VNB N_A_27_74#_c_623_n 0.00195492f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=1.35
cc_50 VNB N_A_27_74#_c_624_n 0.00396969f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=0.74
cc_51 VNB N_A_27_74#_c_625_n 0.00466188f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=0.74
cc_52 VNB N_A_27_74#_c_626_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_53 VNB N_A_27_74#_c_627_n 0.0078054f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_54 VNB N_A_27_74#_c_628_n 0.00962339f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_55 VNB N_A_27_74#_c_629_n 0.00244677f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.515
cc_56 VNB N_A_27_74#_c_630_n 0.00200315f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_57 VNB N_VGND_c_715_n 0.011008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_716_n 0.0114288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_717_n 0.0166826f $X=-0.19 $Y=-0.245 $X2=1.505 $Y2=2.4
cc_60 VNB N_VGND_c_718_n 0.0377021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_719_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=0.74
cc_62 VNB N_VGND_c_720_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_721_n 0.0627368f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.5
cc_64 VNB N_VGND_c_722_n 0.0334841f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_65 VNB N_VGND_c_723_n 0.00634377f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.515
cc_66 VNB N_VGND_c_724_n 0.330625f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.515
cc_67 VPB N_A_M1000_g 0.025802f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_68 VPB N_A_M1002_g 0.0207429f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_69 VPB N_A_M1003_g 0.0205822f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=2.4
cc_70 VPB N_A_M1006_g 0.0216762f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_71 VPB N_A_c_117_n 0.0144606f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_72 VPB N_A_c_118_n 0.0112617f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.515
cc_73 VPB N_A_473_323#_c_210_n 0.0166892f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_74 VPB N_A_473_323#_c_198_n 0.00755315f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_75 VPB N_A_473_323#_c_199_n 0.00356598f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_76 VPB N_A_473_323#_c_213_n 0.0166514f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_473_323#_c_200_n 0.00556401f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_78 VPB N_A_473_323#_c_215_n 0.0158745f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=1.68
cc_79 VPB N_A_473_323#_c_201_n 0.00596183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_473_323#_c_217_n 0.0199821f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=0.74
cc_81 VPB N_A_473_323#_c_202_n 0.0203617f $X=-0.19 $Y=1.66 $X2=1.865 $Y2=1.425
cc_82 VPB N_A_473_323#_c_203_n 0.00200584f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.5
cc_83 VPB N_A_473_323#_c_204_n 0.00200584f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_84 VPB N_A_473_323#_c_205_n 0.00200584f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_85 VPB N_A_473_323#_c_222_n 0.0980889f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_473_323#_c_208_n 0.0223071f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_TE_M1012_g 0.0326324f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.425
cc_88 VPB N_A_27_368#_c_411_n 0.0366851f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=2.4
cc_89 VPB N_A_27_368#_c_412_n 0.00237811f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=0.74
cc_90 VPB N_A_27_368#_c_413_n 0.00971634f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=0.74
cc_91 VPB N_A_27_368#_c_414_n 0.0045905f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_92 VPB N_A_27_368#_c_415_n 2.80234e-19 $X=-0.19 $Y=1.66 $X2=1.995 $Y2=0.74
cc_93 VPB N_A_27_368#_c_416_n 0.00474727f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_94 VPB N_A_27_368#_c_410_n 0.00149825f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_95 VPB N_A_27_368#_c_418_n 0.00226238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_27_368#_c_419_n 0.00584186f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.515
cc_97 VPB N_A_27_368#_c_420_n 0.0022364f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.515
cc_98 VPB N_A_27_368#_c_421_n 0.00181992f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_99 VPB N_Z_c_501_n 0.00151398f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_100 VPB N_VPWR_c_558_n 0.00776029f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_559_n 0.00508627f $X=-0.19 $Y=1.66 $X2=1.505 $Y2=2.4
cc_102 VPB N_VPWR_c_560_n 0.0106521f $X=-0.19 $Y=1.66 $X2=1.52 $Y2=0.74
cc_103 VPB N_VPWR_c_561_n 0.0560452f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_562_n 0.0616265f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_563_n 0.0185253f $X=-0.19 $Y=1.66 $X2=1.967 $Y2=1.425
cc_106 VPB N_VPWR_c_564_n 0.0448319f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_565_n 0.0047791f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.515
cc_108 VPB N_VPWR_c_566_n 0.00478096f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_109 VPB N_VPWR_c_557_n 0.0844912f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_110 N_A_M1006_g N_A_473_323#_c_199_n 0.014569f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_111 N_A_M1016_g N_TE_c_310_n 0.0114134f $X=1.995 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_112 N_A_c_116_n N_TE_c_312_n 0.0114134f $X=1.967 $Y=1.425 $X2=0 $Y2=0
cc_113 N_A_M1000_g N_A_27_368#_c_411_n 0.0124591f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_114 N_A_M1002_g N_A_27_368#_c_411_n 6.17159e-19 $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_115 N_A_c_117_n N_A_27_368#_c_411_n 0.0254478f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_116 N_A_M1000_g N_A_27_368#_c_412_n 0.012228f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_117 N_A_M1002_g N_A_27_368#_c_412_n 0.0144896f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A_M1000_g N_A_27_368#_c_413_n 0.00282152f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A_M1003_g N_A_27_368#_c_414_n 0.0142213f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A_M1006_g N_A_27_368#_c_414_n 0.0141884f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_121 N_A_M1006_g N_A_27_368#_c_415_n 5.21735e-19 $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_122 N_A_M1006_g N_A_27_368#_c_410_n 0.00161029f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_123 N_A_c_116_n N_A_27_368#_c_410_n 2.49919e-19 $X=1.967 $Y=1.425 $X2=0 $Y2=0
cc_124 N_A_M1009_g N_Z_c_504_n 0.00602688f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A_M1013_g N_Z_c_504_n 6.18096e-19 $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A_M1009_g N_Z_c_499_n 0.00952207f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A_M1013_g N_Z_c_499_n 0.0176893f $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A_c_117_n N_Z_c_499_n 0.0367038f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_129 N_A_c_118_n N_Z_c_499_n 0.0045887f $X=1.595 $Y=1.515 $X2=0 $Y2=0
cc_130 N_A_M1007_g N_Z_c_500_n 0.00234945f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A_M1009_g N_Z_c_500_n 0.0026663f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A_c_117_n N_Z_c_500_n 0.0276331f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_133 N_A_c_118_n N_Z_c_500_n 0.00406125f $X=1.595 $Y=1.515 $X2=0 $Y2=0
cc_134 N_A_M1002_g N_Z_c_514_n 0.0132272f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_135 N_A_M1003_g N_Z_c_514_n 0.0173197f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_136 N_A_c_117_n N_Z_c_514_n 0.0333533f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_137 N_A_c_118_n N_Z_c_514_n 7.63416e-19 $X=1.595 $Y=1.515 $X2=0 $Y2=0
cc_138 N_A_M1016_g N_Z_c_518_n 0.00395262f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A_M1013_g N_Z_c_501_n 0.00474402f $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A_c_113_n N_Z_c_501_n 0.0112863f $X=1.865 $Y=1.425 $X2=0 $Y2=0
cc_141 N_A_M1006_g N_Z_c_501_n 0.0120791f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_142 N_A_M1016_g N_Z_c_501_n 0.00156994f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A_c_116_n N_Z_c_501_n 0.00294268f $X=1.967 $Y=1.425 $X2=0 $Y2=0
cc_144 N_A_c_117_n N_Z_c_501_n 0.0326257f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_145 N_A_c_118_n N_Z_c_501_n 0.00423831f $X=1.595 $Y=1.515 $X2=0 $Y2=0
cc_146 N_A_M1002_g N_Z_c_526_n 0.0118549f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_147 N_A_M1003_g N_Z_c_526_n 5.52339e-19 $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_148 N_A_c_117_n N_Z_c_526_n 0.0244752f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_149 N_A_c_118_n N_Z_c_526_n 8.32165e-19 $X=1.595 $Y=1.515 $X2=0 $Y2=0
cc_150 N_A_M1003_g N_Z_c_530_n 0.00196977f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_151 N_A_M1006_g N_Z_c_530_n 0.00192359f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_152 N_A_M1016_g N_Z_c_502_n 0.00512787f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A_M1002_g Z 5.6976e-19 $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_154 N_A_M1003_g Z 0.011357f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_155 N_A_M1006_g Z 0.0095354f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A_M1000_g N_VPWR_c_562_n 0.00333901f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_157 N_A_M1002_g N_VPWR_c_562_n 0.00333926f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_158 N_A_M1003_g N_VPWR_c_562_n 0.00333926f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_159 N_A_M1006_g N_VPWR_c_562_n 0.00333926f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_160 N_A_M1000_g N_VPWR_c_557_n 0.00426886f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_161 N_A_M1002_g N_VPWR_c_557_n 0.00423617f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_162 N_A_M1003_g N_VPWR_c_557_n 0.00423176f $X=1.505 $Y=2.4 $X2=0 $Y2=0
cc_163 N_A_M1006_g N_VPWR_c_557_n 0.00423254f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_164 N_A_M1007_g N_A_27_74#_c_619_n 0.0114672f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A_M1009_g N_A_27_74#_c_619_n 8.28548e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A_c_117_n N_A_27_74#_c_619_n 0.023775f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_167 N_A_M1007_g N_A_27_74#_c_620_n 0.0104643f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A_M1009_g N_A_27_74#_c_620_n 0.0118001f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A_M1007_g N_A_27_74#_c_621_n 0.00282152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A_M1013_g N_A_27_74#_c_622_n 0.00938114f $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A_M1016_g N_A_27_74#_c_622_n 0.0136901f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A_M1016_g N_A_27_74#_c_623_n 0.0052852f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A_M1016_g N_A_27_74#_c_625_n 0.00392472f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A_M1013_g N_A_27_74#_c_629_n 0.00255335f $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A_M1007_g N_VGND_c_721_n 0.00278247f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A_M1009_g N_VGND_c_721_n 0.00278271f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A_M1013_g N_VGND_c_721_n 0.00278271f $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A_M1016_g N_VGND_c_721_n 0.00278271f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A_M1007_g N_VGND_c_724_n 0.00357743f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_180 N_A_M1009_g N_VGND_c_724_n 0.00354959f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_181 N_A_M1013_g N_VGND_c_724_n 0.00354734f $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A_M1016_g N_VGND_c_724_n 0.00354573f $X=1.995 $Y=0.74 $X2=0 $Y2=0
cc_183 N_A_473_323#_c_198_n N_TE_c_311_n 0.0156344f $X=2.865 $Y=1.69 $X2=0 $Y2=0
cc_184 N_A_473_323#_c_199_n N_TE_c_312_n 0.0156344f $X=2.545 $Y=1.69 $X2=0 $Y2=0
cc_185 N_A_473_323#_c_200_n N_TE_c_314_n 0.0156344f $X=3.315 $Y=1.69 $X2=0 $Y2=0
cc_186 N_A_473_323#_c_201_n N_TE_c_316_n 0.0156344f $X=3.775 $Y=1.69 $X2=0 $Y2=0
cc_187 N_A_473_323#_c_206_n N_TE_c_317_n 0.00176266f $X=4.84 $Y=0.515 $X2=0
+ $Y2=0
cc_188 N_A_473_323#_c_206_n N_TE_c_318_n 0.00812744f $X=4.84 $Y=0.515 $X2=0
+ $Y2=0
cc_189 N_A_473_323#_c_207_n N_TE_c_318_n 0.00267162f $X=4.7 $Y=1.64 $X2=0 $Y2=0
cc_190 N_A_473_323#_c_209_n N_TE_c_318_n 0.00684687f $X=4.81 $Y=1.13 $X2=0 $Y2=0
cc_191 N_A_473_323#_c_202_n N_TE_M1012_g 0.0195893f $X=4.395 $Y=1.69 $X2=0 $Y2=0
cc_192 N_A_473_323#_c_208_n N_TE_M1012_g 0.0205343f $X=5.03 $Y=2.815 $X2=0 $Y2=0
cc_193 N_A_473_323#_c_203_n N_TE_c_320_n 0.0156344f $X=2.955 $Y=1.69 $X2=0 $Y2=0
cc_194 N_A_473_323#_c_204_n N_TE_c_321_n 0.0156344f $X=3.405 $Y=1.69 $X2=0 $Y2=0
cc_195 N_A_473_323#_c_205_n N_TE_c_322_n 0.0156344f $X=3.865 $Y=1.69 $X2=0 $Y2=0
cc_196 N_A_473_323#_c_207_n TE 0.00316442f $X=4.7 $Y=1.64 $X2=0 $Y2=0
cc_197 N_A_473_323#_c_202_n N_TE_c_324_n 0.0156344f $X=4.395 $Y=1.69 $X2=0 $Y2=0
cc_198 N_A_473_323#_c_207_n N_TE_c_324_n 0.0141663f $X=4.7 $Y=1.64 $X2=0 $Y2=0
cc_199 N_A_473_323#_c_208_n N_TE_c_324_n 0.00755084f $X=5.03 $Y=2.815 $X2=0
+ $Y2=0
cc_200 N_A_473_323#_c_209_n N_TE_c_324_n 0.00468311f $X=4.81 $Y=1.13 $X2=0 $Y2=0
cc_201 N_A_473_323#_c_202_n N_TE_c_325_n 7.80231e-19 $X=4.395 $Y=1.69 $X2=0
+ $Y2=0
cc_202 N_A_473_323#_c_207_n N_TE_c_325_n 0.00166774f $X=4.7 $Y=1.64 $X2=0 $Y2=0
cc_203 N_A_473_323#_c_208_n N_TE_c_325_n 0.00487879f $X=5.03 $Y=2.815 $X2=0
+ $Y2=0
cc_204 N_A_473_323#_c_207_n N_TE_c_326_n 0.0233109f $X=4.7 $Y=1.64 $X2=0 $Y2=0
cc_205 N_A_473_323#_c_208_n N_TE_c_326_n 0.0165398f $X=5.03 $Y=2.815 $X2=0 $Y2=0
cc_206 N_A_473_323#_c_209_n N_TE_c_326_n 0.00191579f $X=4.81 $Y=1.13 $X2=0 $Y2=0
cc_207 N_A_473_323#_c_210_n N_A_27_368#_c_414_n 0.00356944f $X=2.455 $Y=1.765
+ $X2=0 $Y2=0
cc_208 N_A_473_323#_c_210_n N_A_27_368#_c_415_n 0.0147139f $X=2.455 $Y=1.765
+ $X2=0 $Y2=0
cc_209 N_A_473_323#_c_213_n N_A_27_368#_c_415_n 6.6671e-19 $X=2.955 $Y=1.765
+ $X2=0 $Y2=0
cc_210 N_A_473_323#_c_210_n N_A_27_368#_c_416_n 0.00776692f $X=2.455 $Y=1.765
+ $X2=0 $Y2=0
cc_211 N_A_473_323#_c_198_n N_A_27_368#_c_416_n 0.00740574f $X=2.865 $Y=1.69
+ $X2=0 $Y2=0
cc_212 N_A_473_323#_c_199_n N_A_27_368#_c_416_n 0.00250595f $X=2.545 $Y=1.69
+ $X2=0 $Y2=0
cc_213 N_A_473_323#_c_213_n N_A_27_368#_c_416_n 0.00776692f $X=2.955 $Y=1.765
+ $X2=0 $Y2=0
cc_214 N_A_473_323#_c_203_n N_A_27_368#_c_416_n 0.00249421f $X=2.955 $Y=1.69
+ $X2=0 $Y2=0
cc_215 N_A_473_323#_c_210_n N_A_27_368#_c_410_n 6.21913e-19 $X=2.455 $Y=1.765
+ $X2=0 $Y2=0
cc_216 N_A_473_323#_c_199_n N_A_27_368#_c_410_n 0.00193232f $X=2.545 $Y=1.69
+ $X2=0 $Y2=0
cc_217 N_A_473_323#_c_210_n N_A_27_368#_c_418_n 7.26856e-19 $X=2.455 $Y=1.765
+ $X2=0 $Y2=0
cc_218 N_A_473_323#_c_213_n N_A_27_368#_c_418_n 0.0165257f $X=2.955 $Y=1.765
+ $X2=0 $Y2=0
cc_219 N_A_473_323#_c_215_n N_A_27_368#_c_418_n 7.66408e-19 $X=3.405 $Y=1.765
+ $X2=0 $Y2=0
cc_220 N_A_473_323#_c_200_n N_A_27_368#_c_419_n 8.02435e-19 $X=3.315 $Y=1.69
+ $X2=0 $Y2=0
cc_221 N_A_473_323#_c_215_n N_A_27_368#_c_419_n 0.00880397f $X=3.405 $Y=1.765
+ $X2=0 $Y2=0
cc_222 N_A_473_323#_c_201_n N_A_27_368#_c_419_n 0.00614114f $X=3.775 $Y=1.69
+ $X2=0 $Y2=0
cc_223 N_A_473_323#_c_217_n N_A_27_368#_c_419_n 0.00836635f $X=3.865 $Y=1.765
+ $X2=0 $Y2=0
cc_224 N_A_473_323#_c_202_n N_A_27_368#_c_419_n 0.0088782f $X=4.395 $Y=1.69
+ $X2=0 $Y2=0
cc_225 N_A_473_323#_c_204_n N_A_27_368#_c_419_n 0.00301025f $X=3.405 $Y=1.69
+ $X2=0 $Y2=0
cc_226 N_A_473_323#_c_205_n N_A_27_368#_c_419_n 0.00299764f $X=3.865 $Y=1.69
+ $X2=0 $Y2=0
cc_227 N_A_473_323#_c_222_n N_A_27_368#_c_419_n 2.08714e-19 $X=4.56 $Y=1.805
+ $X2=0 $Y2=0
cc_228 N_A_473_323#_c_208_n N_A_27_368#_c_419_n 0.0113878f $X=5.03 $Y=2.815
+ $X2=0 $Y2=0
cc_229 N_A_473_323#_c_215_n N_A_27_368#_c_420_n 7.70084e-19 $X=3.405 $Y=1.765
+ $X2=0 $Y2=0
cc_230 N_A_473_323#_c_217_n N_A_27_368#_c_420_n 0.016837f $X=3.865 $Y=1.765
+ $X2=0 $Y2=0
cc_231 N_A_473_323#_c_222_n N_A_27_368#_c_420_n 0.00457539f $X=4.56 $Y=1.805
+ $X2=0 $Y2=0
cc_232 N_A_473_323#_c_208_n N_A_27_368#_c_420_n 0.0774029f $X=5.03 $Y=2.815
+ $X2=0 $Y2=0
cc_233 N_A_473_323#_c_213_n N_A_27_368#_c_459_n 6.33476e-19 $X=2.955 $Y=1.765
+ $X2=0 $Y2=0
cc_234 N_A_473_323#_c_200_n N_A_27_368#_c_459_n 0.0058398f $X=3.315 $Y=1.69
+ $X2=0 $Y2=0
cc_235 N_A_473_323#_c_203_n N_A_27_368#_c_459_n 5.03429e-19 $X=2.955 $Y=1.69
+ $X2=0 $Y2=0
cc_236 N_A_473_323#_c_199_n N_Z_c_501_n 2.98035e-19 $X=2.545 $Y=1.69 $X2=0 $Y2=0
cc_237 N_A_473_323#_c_210_n N_VPWR_c_558_n 0.00137311f $X=2.455 $Y=1.765 $X2=0
+ $Y2=0
cc_238 N_A_473_323#_c_198_n N_VPWR_c_558_n 9.95485e-19 $X=2.865 $Y=1.69 $X2=0
+ $Y2=0
cc_239 N_A_473_323#_c_213_n N_VPWR_c_558_n 0.00174963f $X=2.955 $Y=1.765 $X2=0
+ $Y2=0
cc_240 N_A_473_323#_c_213_n N_VPWR_c_559_n 6.81448e-19 $X=2.955 $Y=1.765 $X2=0
+ $Y2=0
cc_241 N_A_473_323#_c_215_n N_VPWR_c_559_n 0.0162681f $X=3.405 $Y=1.765 $X2=0
+ $Y2=0
cc_242 N_A_473_323#_c_201_n N_VPWR_c_559_n 7.11061e-19 $X=3.775 $Y=1.69 $X2=0
+ $Y2=0
cc_243 N_A_473_323#_c_217_n N_VPWR_c_559_n 0.0028988f $X=3.865 $Y=1.765 $X2=0
+ $Y2=0
cc_244 N_A_473_323#_c_208_n N_VPWR_c_559_n 2.7337e-19 $X=5.03 $Y=2.815 $X2=0
+ $Y2=0
cc_245 N_A_473_323#_c_208_n N_VPWR_c_561_n 0.0445655f $X=5.03 $Y=2.815 $X2=0
+ $Y2=0
cc_246 N_A_473_323#_c_210_n N_VPWR_c_562_n 0.00517089f $X=2.455 $Y=1.765 $X2=0
+ $Y2=0
cc_247 N_A_473_323#_c_213_n N_VPWR_c_563_n 0.005209f $X=2.955 $Y=1.765 $X2=0
+ $Y2=0
cc_248 N_A_473_323#_c_215_n N_VPWR_c_563_n 0.00460063f $X=3.405 $Y=1.765 $X2=0
+ $Y2=0
cc_249 N_A_473_323#_c_217_n N_VPWR_c_564_n 0.005209f $X=3.865 $Y=1.765 $X2=0
+ $Y2=0
cc_250 N_A_473_323#_c_222_n N_VPWR_c_564_n 0.00188351f $X=4.56 $Y=1.805 $X2=0
+ $Y2=0
cc_251 N_A_473_323#_c_208_n N_VPWR_c_564_n 0.0353308f $X=5.03 $Y=2.815 $X2=0
+ $Y2=0
cc_252 N_A_473_323#_c_210_n N_VPWR_c_557_n 0.0097786f $X=2.455 $Y=1.765 $X2=0
+ $Y2=0
cc_253 N_A_473_323#_c_213_n N_VPWR_c_557_n 0.00982754f $X=2.955 $Y=1.765 $X2=0
+ $Y2=0
cc_254 N_A_473_323#_c_215_n N_VPWR_c_557_n 0.00908554f $X=3.405 $Y=1.765 $X2=0
+ $Y2=0
cc_255 N_A_473_323#_c_217_n N_VPWR_c_557_n 0.009875f $X=3.865 $Y=1.765 $X2=0
+ $Y2=0
cc_256 N_A_473_323#_c_208_n N_VPWR_c_557_n 0.0292263f $X=5.03 $Y=2.815 $X2=0
+ $Y2=0
cc_257 N_A_473_323#_c_199_n N_A_27_74#_c_624_n 0.00426908f $X=2.545 $Y=1.69
+ $X2=0 $Y2=0
cc_258 N_A_473_323#_c_199_n N_A_27_74#_c_625_n 0.00173232f $X=2.545 $Y=1.69
+ $X2=0 $Y2=0
cc_259 N_A_473_323#_c_202_n N_A_27_74#_c_627_n 0.00700874f $X=4.395 $Y=1.69
+ $X2=0 $Y2=0
cc_260 N_A_473_323#_c_204_n N_A_27_74#_c_627_n 0.00422854f $X=3.405 $Y=1.69
+ $X2=0 $Y2=0
cc_261 N_A_473_323#_c_207_n N_A_27_74#_c_627_n 0.0137368f $X=4.7 $Y=1.64 $X2=0
+ $Y2=0
cc_262 N_A_473_323#_c_208_n N_A_27_74#_c_627_n 0.00445757f $X=5.03 $Y=2.815
+ $X2=0 $Y2=0
cc_263 N_A_473_323#_c_206_n N_A_27_74#_c_628_n 0.0785503f $X=4.84 $Y=0.515 $X2=0
+ $Y2=0
cc_264 N_A_473_323#_c_200_n N_A_27_74#_c_630_n 0.0023761f $X=3.315 $Y=1.69 $X2=0
+ $Y2=0
cc_265 N_A_473_323#_c_206_n N_VGND_c_718_n 0.026158f $X=4.84 $Y=0.515 $X2=0
+ $Y2=0
cc_266 N_A_473_323#_c_206_n N_VGND_c_722_n 0.0172412f $X=4.84 $Y=0.515 $X2=0
+ $Y2=0
cc_267 N_A_473_323#_c_206_n N_VGND_c_724_n 0.0142144f $X=4.84 $Y=0.515 $X2=0
+ $Y2=0
cc_268 N_TE_c_312_n N_A_27_368#_c_416_n 6.07857e-19 $X=2.57 $Y=1.3 $X2=0 $Y2=0
cc_269 N_TE_c_314_n N_A_27_368#_c_419_n 6.73874e-19 $X=3.42 $Y=1.3 $X2=0 $Y2=0
cc_270 N_TE_c_316_n N_A_27_368#_c_419_n 2.50455e-19 $X=3.99 $Y=1.3 $X2=0 $Y2=0
cc_271 N_TE_c_320_n N_A_27_368#_c_459_n 2.51631e-19 $X=3.065 $Y=1.3 $X2=0 $Y2=0
cc_272 N_TE_M1012_g N_VPWR_c_561_n 0.0063662f $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_273 N_TE_c_325_n N_VPWR_c_561_n 0.00595461f $X=5.485 $Y=1.465 $X2=0 $Y2=0
cc_274 N_TE_c_326_n N_VPWR_c_561_n 0.019603f $X=5.485 $Y=1.465 $X2=0 $Y2=0
cc_275 N_TE_M1012_g N_VPWR_c_564_n 0.00519767f $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_276 N_TE_M1012_g N_VPWR_c_557_n 0.00987472f $X=5.255 $Y=2.4 $X2=0 $Y2=0
cc_277 N_TE_c_310_n N_A_27_74#_c_622_n 0.00348233f $X=2.495 $Y=1.225 $X2=0 $Y2=0
cc_278 N_TE_c_310_n N_A_27_74#_c_623_n 0.011268f $X=2.495 $Y=1.225 $X2=0 $Y2=0
cc_279 N_TE_c_312_n N_A_27_74#_c_623_n 0.00315932f $X=2.57 $Y=1.3 $X2=0 $Y2=0
cc_280 N_TE_c_313_n N_A_27_74#_c_623_n 4.34235e-19 $X=3.065 $Y=1.225 $X2=0 $Y2=0
cc_281 N_TE_c_311_n N_A_27_74#_c_624_n 0.0118714f $X=2.99 $Y=1.3 $X2=0 $Y2=0
cc_282 N_TE_c_312_n N_A_27_74#_c_624_n 0.0069434f $X=2.57 $Y=1.3 $X2=0 $Y2=0
cc_283 N_TE_c_320_n N_A_27_74#_c_624_n 0.00696323f $X=3.065 $Y=1.3 $X2=0 $Y2=0
cc_284 N_TE_c_312_n N_A_27_74#_c_625_n 0.00120269f $X=2.57 $Y=1.3 $X2=0 $Y2=0
cc_285 N_TE_c_310_n N_A_27_74#_c_626_n 4.49351e-19 $X=2.495 $Y=1.225 $X2=0 $Y2=0
cc_286 N_TE_c_313_n N_A_27_74#_c_626_n 0.0125068f $X=3.065 $Y=1.225 $X2=0 $Y2=0
cc_287 N_TE_c_314_n N_A_27_74#_c_626_n 0.00434616f $X=3.42 $Y=1.3 $X2=0 $Y2=0
cc_288 N_TE_c_315_n N_A_27_74#_c_626_n 0.0125068f $X=3.495 $Y=1.225 $X2=0 $Y2=0
cc_289 N_TE_c_317_n N_A_27_74#_c_626_n 4.49351e-19 $X=4.065 $Y=1.225 $X2=0 $Y2=0
cc_290 N_TE_c_320_n N_A_27_74#_c_626_n 0.00227103f $X=3.065 $Y=1.3 $X2=0 $Y2=0
cc_291 N_TE_c_321_n N_A_27_74#_c_626_n 0.00227103f $X=3.495 $Y=1.3 $X2=0 $Y2=0
cc_292 N_TE_c_316_n N_A_27_74#_c_627_n 0.0118714f $X=3.99 $Y=1.3 $X2=0 $Y2=0
cc_293 N_TE_c_321_n N_A_27_74#_c_627_n 0.00696323f $X=3.495 $Y=1.3 $X2=0 $Y2=0
cc_294 N_TE_c_322_n N_A_27_74#_c_627_n 0.00726444f $X=4.065 $Y=1.3 $X2=0 $Y2=0
cc_295 N_TE_c_324_n N_A_27_74#_c_627_n 0.00473545f $X=4.98 $Y=1.427 $X2=0 $Y2=0
cc_296 N_TE_c_315_n N_A_27_74#_c_628_n 4.49351e-19 $X=3.495 $Y=1.225 $X2=0 $Y2=0
cc_297 N_TE_c_317_n N_A_27_74#_c_628_n 0.0140897f $X=4.065 $Y=1.225 $X2=0 $Y2=0
cc_298 N_TE_c_318_n N_A_27_74#_c_628_n 0.00123989f $X=5.055 $Y=1.225 $X2=0 $Y2=0
cc_299 N_TE_c_322_n N_A_27_74#_c_628_n 0.00227103f $X=4.065 $Y=1.3 $X2=0 $Y2=0
cc_300 N_TE_c_324_n N_A_27_74#_c_628_n 0.00830924f $X=4.98 $Y=1.427 $X2=0 $Y2=0
cc_301 N_TE_c_314_n N_A_27_74#_c_630_n 0.00334949f $X=3.42 $Y=1.3 $X2=0 $Y2=0
cc_302 N_TE_c_320_n N_A_27_74#_c_630_n 3.01213e-19 $X=3.065 $Y=1.3 $X2=0 $Y2=0
cc_303 N_TE_c_321_n N_A_27_74#_c_630_n 3.01213e-19 $X=3.495 $Y=1.3 $X2=0 $Y2=0
cc_304 N_TE_c_310_n N_VGND_c_715_n 0.00616282f $X=2.495 $Y=1.225 $X2=0 $Y2=0
cc_305 N_TE_c_311_n N_VGND_c_715_n 0.00525645f $X=2.99 $Y=1.3 $X2=0 $Y2=0
cc_306 N_TE_c_313_n N_VGND_c_715_n 0.00666821f $X=3.065 $Y=1.225 $X2=0 $Y2=0
cc_307 N_TE_c_315_n N_VGND_c_716_n 0.00666821f $X=3.495 $Y=1.225 $X2=0 $Y2=0
cc_308 N_TE_c_316_n N_VGND_c_716_n 0.00525645f $X=3.99 $Y=1.3 $X2=0 $Y2=0
cc_309 N_TE_c_317_n N_VGND_c_716_n 0.00805013f $X=4.065 $Y=1.225 $X2=0 $Y2=0
cc_310 N_TE_c_318_n N_VGND_c_718_n 0.0174858f $X=5.055 $Y=1.225 $X2=0 $Y2=0
cc_311 TE N_VGND_c_718_n 0.00881431f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_312 N_TE_c_325_n N_VGND_c_718_n 0.00679144f $X=5.485 $Y=1.465 $X2=0 $Y2=0
cc_313 N_TE_c_326_n N_VGND_c_718_n 0.0121897f $X=5.485 $Y=1.465 $X2=0 $Y2=0
cc_314 N_TE_c_313_n N_VGND_c_719_n 0.00434272f $X=3.065 $Y=1.225 $X2=0 $Y2=0
cc_315 N_TE_c_315_n N_VGND_c_719_n 0.00434272f $X=3.495 $Y=1.225 $X2=0 $Y2=0
cc_316 N_TE_c_310_n N_VGND_c_721_n 0.00430908f $X=2.495 $Y=1.225 $X2=0 $Y2=0
cc_317 N_TE_c_317_n N_VGND_c_722_n 0.00434272f $X=4.065 $Y=1.225 $X2=0 $Y2=0
cc_318 N_TE_c_318_n N_VGND_c_722_n 0.00434272f $X=5.055 $Y=1.225 $X2=0 $Y2=0
cc_319 N_TE_c_310_n N_VGND_c_724_n 0.00817403f $X=2.495 $Y=1.225 $X2=0 $Y2=0
cc_320 N_TE_c_313_n N_VGND_c_724_n 0.00821294f $X=3.065 $Y=1.225 $X2=0 $Y2=0
cc_321 N_TE_c_315_n N_VGND_c_724_n 0.00821294f $X=3.495 $Y=1.225 $X2=0 $Y2=0
cc_322 N_TE_c_317_n N_VGND_c_724_n 0.00826293f $X=4.065 $Y=1.225 $X2=0 $Y2=0
cc_323 N_TE_c_318_n N_VGND_c_724_n 0.0082925f $X=5.055 $Y=1.225 $X2=0 $Y2=0
cc_324 N_A_27_368#_c_412_n N_Z_M1000_d 0.00213667f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_325 N_A_27_368#_c_414_n N_Z_M1003_d 0.00165831f $X=2.065 $Y=2.99 $X2=0 $Y2=0
cc_326 N_A_27_368#_M1002_s N_Z_c_514_n 0.00410979f $X=1.095 $Y=1.84 $X2=0 $Y2=0
cc_327 N_A_27_368#_c_469_p N_Z_c_514_n 0.0167599f $X=1.28 $Y=2.455 $X2=0 $Y2=0
cc_328 N_A_27_368#_c_415_n N_Z_c_501_n 0.0062509f $X=2.23 $Y=1.985 $X2=0 $Y2=0
cc_329 N_A_27_368#_c_410_n N_Z_c_501_n 0.014175f $X=2.395 $Y=1.725 $X2=0 $Y2=0
cc_330 N_A_27_368#_c_412_n N_Z_c_526_n 0.0173278f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_331 N_A_27_368#_c_414_n Z 0.0159318f $X=2.065 $Y=2.99 $X2=0 $Y2=0
cc_332 N_A_27_368#_c_414_n N_VPWR_c_558_n 0.0117278f $X=2.065 $Y=2.99 $X2=0
+ $Y2=0
cc_333 N_A_27_368#_c_416_n N_VPWR_c_558_n 0.0186218f $X=3.015 $Y=1.725 $X2=0
+ $Y2=0
cc_334 N_A_27_368#_c_418_n N_VPWR_c_558_n 0.0322491f $X=3.18 $Y=1.985 $X2=0
+ $Y2=0
cc_335 N_A_27_368#_c_418_n N_VPWR_c_559_n 0.0324396f $X=3.18 $Y=1.985 $X2=0
+ $Y2=0
cc_336 N_A_27_368#_c_419_n N_VPWR_c_559_n 0.0182752f $X=3.925 $Y=1.725 $X2=0
+ $Y2=0
cc_337 N_A_27_368#_c_420_n N_VPWR_c_559_n 0.0322531f $X=4.09 $Y=1.985 $X2=0
+ $Y2=0
cc_338 N_A_27_368#_c_412_n N_VPWR_c_562_n 0.0421297f $X=1.115 $Y=2.99 $X2=0
+ $Y2=0
cc_339 N_A_27_368#_c_413_n N_VPWR_c_562_n 0.0235688f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_340 N_A_27_368#_c_414_n N_VPWR_c_562_n 0.0675378f $X=2.065 $Y=2.99 $X2=0
+ $Y2=0
cc_341 N_A_27_368#_c_421_n N_VPWR_c_562_n 0.0179217f $X=1.24 $Y=2.99 $X2=0 $Y2=0
cc_342 N_A_27_368#_c_418_n N_VPWR_c_563_n 0.0109793f $X=3.18 $Y=1.985 $X2=0
+ $Y2=0
cc_343 N_A_27_368#_c_420_n N_VPWR_c_564_n 0.0109793f $X=4.09 $Y=1.985 $X2=0
+ $Y2=0
cc_344 N_A_27_368#_c_412_n N_VPWR_c_557_n 0.0236586f $X=1.115 $Y=2.99 $X2=0
+ $Y2=0
cc_345 N_A_27_368#_c_413_n N_VPWR_c_557_n 0.0127152f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_346 N_A_27_368#_c_414_n N_VPWR_c_557_n 0.0373646f $X=2.065 $Y=2.99 $X2=0
+ $Y2=0
cc_347 N_A_27_368#_c_418_n N_VPWR_c_557_n 0.00901959f $X=3.18 $Y=1.985 $X2=0
+ $Y2=0
cc_348 N_A_27_368#_c_420_n N_VPWR_c_557_n 0.00901959f $X=4.09 $Y=1.985 $X2=0
+ $Y2=0
cc_349 N_A_27_368#_c_421_n N_VPWR_c_557_n 0.00971942f $X=1.24 $Y=2.99 $X2=0
+ $Y2=0
cc_350 N_A_27_368#_c_416_n N_A_27_74#_c_624_n 0.0406282f $X=3.015 $Y=1.725 $X2=0
+ $Y2=0
cc_351 N_A_27_368#_c_459_n N_A_27_74#_c_624_n 0.00791142f $X=3.14 $Y=1.725 $X2=0
+ $Y2=0
cc_352 N_A_27_368#_c_416_n N_A_27_74#_c_625_n 0.00399999f $X=3.015 $Y=1.725
+ $X2=0 $Y2=0
cc_353 N_A_27_368#_c_410_n N_A_27_74#_c_625_n 0.0260989f $X=2.395 $Y=1.725 $X2=0
+ $Y2=0
cc_354 N_A_27_368#_c_419_n N_A_27_74#_c_627_n 0.0546439f $X=3.925 $Y=1.725 $X2=0
+ $Y2=0
cc_355 N_A_27_368#_c_419_n N_A_27_74#_c_630_n 0.0144544f $X=3.925 $Y=1.725 $X2=0
+ $Y2=0
cc_356 N_A_27_368#_c_459_n N_A_27_74#_c_630_n 0.0133727f $X=3.14 $Y=1.725 $X2=0
+ $Y2=0
cc_357 N_Z_c_499_n N_A_27_74#_M1009_d 0.00312259f $X=1.615 $Y=1.095 $X2=0 $Y2=0
cc_358 N_Z_c_500_n N_A_27_74#_c_619_n 0.00540984f $X=0.945 $Y=1.095 $X2=0 $Y2=0
cc_359 N_Z_M1007_s N_A_27_74#_c_620_n 0.00289516f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_360 N_Z_c_504_n N_A_27_74#_c_620_n 0.0145454f $X=0.78 $Y=0.825 $X2=0 $Y2=0
cc_361 N_Z_c_499_n N_A_27_74#_c_620_n 0.00304353f $X=1.615 $Y=1.095 $X2=0 $Y2=0
cc_362 N_Z_c_499_n N_A_27_74#_c_689_n 0.0178215f $X=1.615 $Y=1.095 $X2=0 $Y2=0
cc_363 N_Z_M1013_s N_A_27_74#_c_622_n 0.00258847f $X=1.595 $Y=0.37 $X2=0 $Y2=0
cc_364 N_Z_c_499_n N_A_27_74#_c_622_n 0.00364245f $X=1.615 $Y=1.095 $X2=0 $Y2=0
cc_365 N_Z_c_518_n N_A_27_74#_c_622_n 0.0133715f $X=1.78 $Y=0.825 $X2=0 $Y2=0
cc_366 N_Z_c_501_n N_A_27_74#_c_623_n 0.00816149f $X=1.755 $Y=1.95 $X2=0 $Y2=0
cc_367 N_Z_c_502_n N_A_27_74#_c_623_n 0.0100439f $X=1.78 $Y=1.095 $X2=0 $Y2=0
cc_368 N_Z_c_501_n N_A_27_74#_c_625_n 0.0118914f $X=1.755 $Y=1.95 $X2=0 $Y2=0
cc_369 N_A_27_74#_c_622_n N_VGND_c_715_n 0.011924f $X=2.115 $Y=0.34 $X2=0 $Y2=0
cc_370 N_A_27_74#_c_623_n N_VGND_c_715_n 0.0272062f $X=2.28 $Y=0.515 $X2=0 $Y2=0
cc_371 N_A_27_74#_c_624_n N_VGND_c_715_n 0.0264638f $X=3.115 $Y=1.385 $X2=0
+ $Y2=0
cc_372 N_A_27_74#_c_626_n N_VGND_c_715_n 0.0308484f $X=3.28 $Y=0.515 $X2=0 $Y2=0
cc_373 N_A_27_74#_c_626_n N_VGND_c_716_n 0.0308485f $X=3.28 $Y=0.515 $X2=0 $Y2=0
cc_374 N_A_27_74#_c_627_n N_VGND_c_716_n 0.0264638f $X=4.115 $Y=1.385 $X2=0
+ $Y2=0
cc_375 N_A_27_74#_c_628_n N_VGND_c_716_n 0.0308485f $X=4.28 $Y=0.515 $X2=0 $Y2=0
cc_376 N_A_27_74#_c_626_n N_VGND_c_719_n 0.0144922f $X=3.28 $Y=0.515 $X2=0 $Y2=0
cc_377 N_A_27_74#_c_620_n N_VGND_c_721_n 0.0423044f $X=1.115 $Y=0.34 $X2=0 $Y2=0
cc_378 N_A_27_74#_c_621_n N_VGND_c_721_n 0.0235688f $X=0.445 $Y=0.34 $X2=0 $Y2=0
cc_379 N_A_27_74#_c_622_n N_VGND_c_721_n 0.0658004f $X=2.115 $Y=0.34 $X2=0 $Y2=0
cc_380 N_A_27_74#_c_629_n N_VGND_c_721_n 0.023268f $X=1.28 $Y=0.34 $X2=0 $Y2=0
cc_381 N_A_27_74#_c_628_n N_VGND_c_722_n 0.0145639f $X=4.28 $Y=0.515 $X2=0 $Y2=0
cc_382 N_A_27_74#_c_620_n N_VGND_c_724_n 0.0239316f $X=1.115 $Y=0.34 $X2=0 $Y2=0
cc_383 N_A_27_74#_c_621_n N_VGND_c_724_n 0.0127152f $X=0.445 $Y=0.34 $X2=0 $Y2=0
cc_384 N_A_27_74#_c_622_n N_VGND_c_724_n 0.0365331f $X=2.115 $Y=0.34 $X2=0 $Y2=0
cc_385 N_A_27_74#_c_626_n N_VGND_c_724_n 0.0118826f $X=3.28 $Y=0.515 $X2=0 $Y2=0
cc_386 N_A_27_74#_c_628_n N_VGND_c_724_n 0.0119984f $X=4.28 $Y=0.515 $X2=0 $Y2=0
cc_387 N_A_27_74#_c_629_n N_VGND_c_724_n 0.0127566f $X=1.28 $Y=0.34 $X2=0 $Y2=0

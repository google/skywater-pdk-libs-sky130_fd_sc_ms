* File: sky130_fd_sc_ms__and2_4.pex.spice
* Created: Fri Aug 28 17:10:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__AND2_4%A_83_269# 1 2 3 12 14 16 17 19 22 24 26 29 33
+ 35 37 38 47 48 49 52 54 58 60 61 63 66 68 69 80
c147 38 0 9.81068e-20 $X=1.885 $Y=1.51
c148 35 0 4.21777e-20 $X=1.935 $Y=1.345
r149 79 80 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=1.875 $Y=1.51
+ $X2=1.935 $Y2=1.51
r150 76 77 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=1.355 $Y=1.51
+ $X2=1.405 $Y2=1.51
r151 73 74 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=0.925 $Y=1.51
+ $X2=0.955 $Y2=1.51
r152 72 73 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=0.505 $Y=1.51
+ $X2=0.925 $Y2=1.51
r153 70 72 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.51
+ $X2=0.505 $Y2=1.51
r154 64 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.585 $Y=2.12
+ $X2=3.585 $Y2=2.035
r155 64 66 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.585 $Y=2.12
+ $X2=3.585 $Y2=2.19
r156 63 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.585 $Y=1.95
+ $X2=3.585 $Y2=2.035
r157 62 63 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.585 $Y=1.28
+ $X2=3.585 $Y2=1.95
r158 60 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.5 $Y=1.195
+ $X2=3.585 $Y2=1.28
r159 60 61 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.5 $Y=1.195
+ $X2=3.325 $Y2=1.195
r160 56 61 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.16 $Y=1.11
+ $X2=3.325 $Y2=1.195
r161 56 58 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=3.16 $Y=1.11
+ $X2=3.16 $Y2=0.72
r162 55 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.8 $Y=2.035
+ $X2=2.635 $Y2=2.035
r163 54 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.5 $Y=2.035
+ $X2=3.585 $Y2=2.035
r164 54 55 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.5 $Y=2.035 $X2=2.8
+ $Y2=2.035
r165 50 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.635 $Y=2.12
+ $X2=2.635 $Y2=2.035
r166 50 52 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=2.635 $Y=2.12
+ $X2=2.635 $Y2=2.19
r167 48 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.47 $Y=2.035
+ $X2=2.635 $Y2=2.035
r168 48 49 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=2.47 $Y=2.035
+ $X2=2.055 $Y2=2.035
r169 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.97 $Y=1.95
+ $X2=2.055 $Y2=2.035
r170 46 47 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.97 $Y=1.675
+ $X2=1.97 $Y2=1.95
r171 45 79 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.85 $Y=1.51
+ $X2=1.875 $Y2=1.51
r172 45 77 77.8133 $w=3.3e-07 $l=4.45e-07 $layer=POLY_cond $X=1.85 $Y=1.51
+ $X2=1.405 $Y2=1.51
r173 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.85
+ $Y=1.51 $X2=1.85 $Y2=1.51
r174 41 76 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=1.17 $Y=1.51
+ $X2=1.355 $Y2=1.51
r175 41 74 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.17 $Y=1.51
+ $X2=0.955 $Y2=1.51
r176 40 44 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.17 $Y=1.51
+ $X2=1.85 $Y2=1.51
r177 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.51 $X2=1.17 $Y2=1.51
r178 38 46 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.885 $Y=1.51
+ $X2=1.97 $Y2=1.675
r179 38 44 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=1.885 $Y=1.51
+ $X2=1.85 $Y2=1.51
r180 35 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.935 $Y=1.345
+ $X2=1.935 $Y2=1.51
r181 35 37 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.935 $Y=1.345
+ $X2=1.935 $Y2=0.865
r182 31 79 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.875 $Y=1.675
+ $X2=1.875 $Y2=1.51
r183 31 33 281.815 $w=1.8e-07 $l=7.25e-07 $layer=POLY_cond $X=1.875 $Y=1.675
+ $X2=1.875 $Y2=2.4
r184 27 77 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.675
+ $X2=1.405 $Y2=1.51
r185 27 29 281.815 $w=1.8e-07 $l=7.25e-07 $layer=POLY_cond $X=1.405 $Y=1.675
+ $X2=1.405 $Y2=2.4
r186 24 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.345
+ $X2=1.355 $Y2=1.51
r187 24 26 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.355 $Y=1.345
+ $X2=1.355 $Y2=0.865
r188 20 74 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.675
+ $X2=0.955 $Y2=1.51
r189 20 22 281.815 $w=1.8e-07 $l=7.25e-07 $layer=POLY_cond $X=0.955 $Y=1.675
+ $X2=0.955 $Y2=2.4
r190 17 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.345
+ $X2=0.925 $Y2=1.51
r191 17 19 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.925 $Y=1.345
+ $X2=0.925 $Y2=0.865
r192 14 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.345
+ $X2=0.495 $Y2=1.51
r193 14 16 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.345
+ $X2=0.495 $Y2=0.865
r194 10 72 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.675
+ $X2=0.505 $Y2=1.51
r195 10 12 281.815 $w=1.8e-07 $l=7.25e-07 $layer=POLY_cond $X=0.505 $Y=1.675
+ $X2=0.505 $Y2=2.4
r196 3 66 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.45
+ $Y=2.045 $X2=3.585 $Y2=2.19
r197 2 52 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.5
+ $Y=2.045 $X2=2.635 $Y2=2.19
r198 1 58 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=2.975
+ $Y=0.595 $X2=3.16 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_MS__AND2_4%A 3 7 11 13 15 17
c47 17 0 2.42266e-19 $X=3.12 $Y=1.665
r48 23 25 32.2928 $w=4.65e-07 $l=2.7e-07 $layer=POLY_cond $X=3.09 $Y=1.682
+ $X2=3.36 $Y2=1.682
r49 17 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.615 $X2=3.09 $Y2=1.615
r50 13 25 1.79404 $w=4.65e-07 $l=1.5e-08 $layer=POLY_cond $X=3.375 $Y=1.682
+ $X2=3.36 $Y2=1.682
r51 13 15 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=3.375 $Y=1.45
+ $X2=3.375 $Y2=0.915
r52 9 25 25.0876 $w=1.8e-07 $l=2.33e-07 $layer=POLY_cond $X=3.36 $Y=1.915
+ $X2=3.36 $Y2=1.682
r53 9 11 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=3.36 $Y=1.915 $X2=3.36
+ $Y2=2.465
r54 5 23 22.7246 $w=4.65e-07 $l=1.9e-07 $layer=POLY_cond $X=2.9 $Y=1.682
+ $X2=3.09 $Y2=1.682
r55 5 19 1.79404 $w=4.65e-07 $l=1.5e-08 $layer=POLY_cond $X=2.9 $Y=1.682
+ $X2=2.885 $Y2=1.682
r56 5 7 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.9 $Y=1.45 $X2=2.9
+ $Y2=0.915
r57 1 19 25.0876 $w=1.8e-07 $l=2.33e-07 $layer=POLY_cond $X=2.885 $Y=1.915
+ $X2=2.885 $Y2=1.682
r58 1 3 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=2.885 $Y=1.915
+ $X2=2.885 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_MS__AND2_4%B 3 8 9 10 11 13 18 20 23
c71 23 0 1.68219e-19 $X=2.42 $Y=1.51
c72 3 0 7.40463e-20 $X=2.41 $Y=2.465
r73 23 26 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.42 $Y=1.51
+ $X2=2.42 $Y2=1.675
r74 23 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.42 $Y=1.51
+ $X2=2.42 $Y2=1.345
r75 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.42
+ $Y=1.51 $X2=2.42 $Y2=1.51
r76 20 24 5.82845 $w=4.33e-07 $l=2.2e-07 $layer=LI1_cond $X=2.64 $Y=1.562
+ $X2=2.42 $Y2=1.562
r77 18 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.825 $Y=0.915
+ $X2=3.825 $Y2=1.31
r78 15 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.825 $Y=0.255
+ $X2=3.825 $Y2=0.915
r79 11 19 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.81 $Y=1.4 $X2=3.81
+ $Y2=1.31
r80 11 13 413.976 $w=1.8e-07 $l=1.065e-06 $layer=POLY_cond $X=3.81 $Y=1.4
+ $X2=3.81 $Y2=2.465
r81 9 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.75 $Y=0.18
+ $X2=3.825 $Y2=0.255
r82 9 10 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=3.75 $Y=0.18
+ $X2=2.52 $Y2=0.18
r83 8 25 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.445 $Y=0.915
+ $X2=2.445 $Y2=1.345
r84 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.445 $Y=0.255
+ $X2=2.52 $Y2=0.18
r85 5 8 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.445 $Y=0.255
+ $X2=2.445 $Y2=0.915
r86 3 26 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=2.41 $Y=2.465
+ $X2=2.41 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_MS__AND2_4%VPWR 1 2 3 4 5 16 18 24 28 32 34 36 39 40 41
+ 47 51 56 65 68 72
r73 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r74 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r75 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r76 60 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r77 60 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r78 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r79 57 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.3 $Y=3.33
+ $X2=3.135 $Y2=3.33
r80 57 59 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.3 $Y=3.33 $X2=3.6
+ $Y2=3.33
r81 56 71 4.72267 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=3.87 $Y=3.33
+ $X2=4.095 $Y2=3.33
r82 56 59 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.87 $Y=3.33 $X2=3.6
+ $Y2=3.33
r83 55 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r84 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r85 52 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=3.33
+ $X2=2.1 $Y2=3.33
r86 52 54 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.265 $Y=3.33
+ $X2=2.64 $Y2=3.33
r87 51 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.97 $Y=3.33
+ $X2=3.135 $Y2=3.33
r88 51 54 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.97 $Y=3.33
+ $X2=2.64 $Y2=3.33
r89 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r90 47 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.935 $Y=3.33
+ $X2=2.1 $Y2=3.33
r91 47 49 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.935 $Y=3.33
+ $X2=1.68 $Y2=3.33
r92 46 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r93 46 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r94 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r95 43 62 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r96 43 45 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r97 41 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r98 41 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r99 41 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r100 39 45 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r101 39 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.14 $Y2=3.33
r102 38 49 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.68 $Y2=3.33
r103 38 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.14 $Y2=3.33
r104 34 71 3.0435 $w=3.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=4.035 $Y=3.245
+ $X2=4.095 $Y2=3.33
r105 34 36 36.8433 $w=3.28e-07 $l=1.055e-06 $layer=LI1_cond $X=4.035 $Y=3.245
+ $X2=4.035 $Y2=2.19
r106 30 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=3.245
+ $X2=3.135 $Y2=3.33
r107 30 32 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.135 $Y=3.245
+ $X2=3.135 $Y2=2.415
r108 26 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.1 $Y=3.245 $X2=2.1
+ $Y2=3.33
r109 26 28 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.1 $Y=3.245
+ $X2=2.1 $Y2=2.455
r110 22 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=3.33
r111 22 24 41.2575 $w=2.48e-07 $l=8.95e-07 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=2.35
r112 18 21 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r113 16 62 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r114 16 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r115 5 36 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.9
+ $Y=2.045 $X2=4.035 $Y2=2.19
r116 4 32 300 $w=1.7e-07 $l=4.42832e-07 $layer=licon1_PDIFF $count=2 $X=2.975
+ $Y=2.045 $X2=3.135 $Y2=2.415
r117 3 28 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.965
+ $Y=1.84 $X2=2.1 $Y2=2.455
r118 2 24 300 $w=1.7e-07 $l=5.73542e-07 $layer=licon1_PDIFF $count=2 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.35
r119 1 21 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r120 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__AND2_4%X 1 2 3 4 15 21 23 25 27 29 33 36 39 42 48 50
c63 42 0 1.92991e-19 $X=0.635 $Y=1.58
r64 45 50 1.19218 $w=2.88e-07 $l=3e-08 $layer=LI1_cond $X=0.69 $Y=1.695 $X2=0.69
+ $Y2=1.665
r65 42 50 1.1127 $w=2.88e-07 $l=2.8e-08 $layer=LI1_cond $X=0.69 $Y=1.637
+ $X2=0.69 $Y2=1.665
r66 42 48 3.7084 $w=2.88e-07 $l=8.7e-08 $layer=LI1_cond $X=0.69 $Y=1.637
+ $X2=0.69 $Y2=1.55
r67 42 45 1.07296 $w=2.88e-07 $l=2.7e-08 $layer=LI1_cond $X=0.69 $Y=1.722
+ $X2=0.69 $Y2=1.695
r68 37 42 4.88795 $w=2.88e-07 $l=1.23e-07 $layer=LI1_cond $X=0.69 $Y=1.845
+ $X2=0.69 $Y2=1.722
r69 37 39 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.845 $X2=0.69
+ $Y2=1.93
r70 31 33 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=1.6 $Y=1.005
+ $X2=1.6 $Y2=0.64
r71 27 41 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=2.015
+ $X2=1.59 $Y2=1.93
r72 27 29 36.8782 $w=2.48e-07 $l=8e-07 $layer=LI1_cond $X=1.59 $Y=2.015 $X2=1.59
+ $Y2=2.815
r73 26 39 3.18746 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.835 $Y=1.93
+ $X2=0.69 $Y2=1.93
r74 25 41 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.465 $Y=1.93
+ $X2=1.59 $Y2=1.93
r75 25 26 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.465 $Y=1.93
+ $X2=0.835 $Y2=1.93
r76 24 36 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=1.09
+ $X2=0.67 $Y2=1.09
r77 23 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.475 $Y=1.09
+ $X2=1.6 $Y2=1.005
r78 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.475 $Y=1.09
+ $X2=0.795 $Y2=1.09
r79 19 39 3.351 $w=2.8e-07 $l=8.9861e-08 $layer=LI1_cond $X=0.68 $Y=2.015
+ $X2=0.69 $Y2=1.93
r80 19 21 34.1465 $w=2.68e-07 $l=8e-07 $layer=LI1_cond $X=0.68 $Y=2.015 $X2=0.68
+ $Y2=2.815
r81 17 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=1.175
+ $X2=0.67 $Y2=1.09
r82 17 48 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=0.67 $Y=1.175
+ $X2=0.67 $Y2=1.55
r83 13 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=1.005
+ $X2=0.67 $Y2=1.09
r84 13 15 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=0.67 $Y=1.005
+ $X2=0.67 $Y2=0.64
r85 4 41 400 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.84 $X2=1.63 $Y2=2.01
r86 4 29 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.84 $X2=1.63 $Y2=2.815
r87 3 39 400 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.01
r88 3 21 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.815
r89 2 33 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.43
+ $Y=0.495 $X2=1.64 $Y2=0.64
r90 1 36 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.495 $X2=0.71 $Y2=1.09
r91 1 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.495 $X2=0.71 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_MS__AND2_4%VGND 1 2 3 4 13 15 19 23 25 27 29 31 36 41 53
+ 56 60
r60 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r61 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r62 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r63 48 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r64 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r65 45 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r66 44 47 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r67 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r68 42 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.15
+ $Y2=0
r69 42 44 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.64
+ $Y2=0
r70 41 59 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=3.875 $Y=0 $X2=4.097
+ $Y2=0
r71 41 47 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.875 $Y=0 $X2=3.6
+ $Y2=0
r72 40 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r73 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r74 37 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.14
+ $Y2=0
r75 37 39 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.68
+ $Y2=0
r76 36 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.985 $Y=0 $X2=2.15
+ $Y2=0
r77 36 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=0 $X2=1.68
+ $Y2=0
r78 35 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r79 35 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r80 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r81 32 50 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r82 32 34 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.72
+ $Y2=0
r83 31 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.14
+ $Y2=0
r84 31 34 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=0.72
+ $Y2=0
r85 29 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r86 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r87 29 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r88 25 59 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.097 $Y2=0
r89 25 27 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0.74
r90 21 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=0.085
+ $X2=2.15 $Y2=0
r91 21 23 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.15 $Y=0.085
+ $X2=2.15 $Y2=0.7
r92 17 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0
r93 17 19 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0.67
r94 13 50 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r95 13 15 25.5842 $w=2.48e-07 $l=5.55e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.64
r96 4 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.9
+ $Y=0.595 $X2=4.04 $Y2=0.74
r97 3 23 91 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=2 $X=2.01
+ $Y=0.495 $X2=2.15 $Y2=0.7
r98 2 19 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.495 $X2=1.14 $Y2=0.67
r99 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.495 $X2=0.28 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_MS__AND2_4%A_504_119# 1 2 9 11 12 15
c29 12 0 4.21777e-20 $X=2.825 $Y=0.34
r30 13 15 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.59 $Y=0.425
+ $X2=3.59 $Y2=0.755
r31 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.505 $Y=0.34
+ $X2=3.59 $Y2=0.425
r32 11 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.505 $Y=0.34
+ $X2=2.825 $Y2=0.34
r33 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.66 $Y=0.425
+ $X2=2.825 $Y2=0.34
r34 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.66 $Y=0.425
+ $X2=2.66 $Y2=0.72
r35 2 15 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=3.45
+ $Y=0.595 $X2=3.59 $Y2=0.755
r36 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.52
+ $Y=0.595 $X2=2.66 $Y2=0.72
.ends


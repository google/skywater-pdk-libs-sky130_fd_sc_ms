* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fah_4 A B CI VGND VNB VPB VPWR COUT SUM
X0 VPWR a_1278_102# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 a_200_74# B a_536_114# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X2 VPWR B a_586_257# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 a_1378_125# CI VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X4 a_430_362# B a_536_114# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 SUM a_1278_102# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X6 SUM a_1278_102# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_531_362# a_586_257# a_200_74# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X8 VGND A a_200_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 VPWR a_1268_379# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X10 VPWR a_1278_102# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X11 COUT a_1268_379# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 VGND a_1268_379# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 VGND a_1268_379# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 a_1378_125# CI VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 a_200_74# B a_531_362# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X16 a_1183_102# a_531_362# a_1278_102# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X17 a_1278_102# a_536_114# a_1378_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X18 a_1183_102# a_1378_125# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X19 a_1278_102# a_536_114# a_1183_102# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X20 VGND a_27_74# a_430_362# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 VGND B a_586_257# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 COUT a_1268_379# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 VPWR A a_200_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X24 a_1268_379# a_536_114# a_1378_125# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X25 a_1183_102# a_1378_125# VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X26 VPWR a_1268_379# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X27 a_1378_125# a_531_362# a_1268_379# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X28 a_536_114# a_586_257# a_430_362# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X29 a_1378_125# a_531_362# a_1278_102# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X30 a_1268_379# a_536_114# a_586_257# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X31 VGND a_1278_102# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X32 a_586_257# a_531_362# a_1268_379# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X33 COUT a_1268_379# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X34 SUM a_1278_102# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X35 VPWR a_27_74# a_430_362# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X36 COUT a_1268_379# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X37 a_27_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X38 a_430_362# B a_531_362# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X39 a_536_114# a_586_257# a_200_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X40 a_27_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X41 VGND a_1278_102# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X42 a_531_362# a_586_257# a_430_362# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X43 SUM a_1278_102# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

* File: sky130_fd_sc_ms__sdfsbp_1.pxi.spice
* Created: Wed Sep  2 12:30:54 2020
* 
x_PM_SKY130_FD_SC_MS__SDFSBP_1%SCE N_SCE_M1010_g N_SCE_M1036_g N_SCE_c_302_n
+ N_SCE_M1011_g N_SCE_M1015_g N_SCE_c_304_n N_SCE_c_296_n N_SCE_c_297_n
+ N_SCE_c_298_n SCE N_SCE_c_299_n N_SCE_c_300_n PM_SKY130_FD_SC_MS__SDFSBP_1%SCE
x_PM_SKY130_FD_SC_MS__SDFSBP_1%A_27_74# N_A_27_74#_M1036_s N_A_27_74#_M1010_s
+ N_A_27_74#_M1039_g N_A_27_74#_M1002_g N_A_27_74#_c_372_n N_A_27_74#_c_373_n
+ N_A_27_74#_c_379_n N_A_27_74#_c_380_n N_A_27_74#_c_374_n N_A_27_74#_c_375_n
+ N_A_27_74#_c_381_n N_A_27_74#_c_382_n N_A_27_74#_c_376_n N_A_27_74#_c_383_n
+ PM_SKY130_FD_SC_MS__SDFSBP_1%A_27_74#
x_PM_SKY130_FD_SC_MS__SDFSBP_1%D N_D_M1017_g N_D_M1040_g D N_D_c_459_n
+ N_D_c_460_n PM_SKY130_FD_SC_MS__SDFSBP_1%D
x_PM_SKY130_FD_SC_MS__SDFSBP_1%SCD N_SCD_c_495_n N_SCD_M1016_g N_SCD_c_499_n
+ N_SCD_M1013_g N_SCD_c_496_n N_SCD_c_497_n SCD SCD SCD
+ PM_SKY130_FD_SC_MS__SDFSBP_1%SCD
x_PM_SKY130_FD_SC_MS__SDFSBP_1%CLK N_CLK_c_539_n N_CLK_M1023_g N_CLK_c_540_n
+ N_CLK_M1026_g CLK PM_SKY130_FD_SC_MS__SDFSBP_1%CLK
x_PM_SKY130_FD_SC_MS__SDFSBP_1%A_781_74# N_A_781_74#_M1019_d N_A_781_74#_M1030_d
+ N_A_781_74#_M1022_g N_A_781_74#_M1007_g N_A_781_74#_M1025_g
+ N_A_781_74#_M1033_g N_A_781_74#_c_574_n N_A_781_74#_c_584_n
+ N_A_781_74#_c_575_n N_A_781_74#_c_576_n N_A_781_74#_c_585_n
+ N_A_781_74#_c_586_n N_A_781_74#_c_577_n N_A_781_74#_c_587_n
+ N_A_781_74#_c_578_n N_A_781_74#_c_589_n N_A_781_74#_c_590_n
+ N_A_781_74#_c_591_n N_A_781_74#_c_592_n N_A_781_74#_c_593_n
+ N_A_781_74#_c_594_n N_A_781_74#_c_595_n N_A_781_74#_c_596_n
+ N_A_781_74#_c_597_n N_A_781_74#_c_598_n N_A_781_74#_c_579_n
+ N_A_781_74#_c_599_n N_A_781_74#_c_580_n N_A_781_74#_c_581_n
+ N_A_781_74#_c_601_n N_A_781_74#_c_602_n PM_SKY130_FD_SC_MS__SDFSBP_1%A_781_74#
x_PM_SKY130_FD_SC_MS__SDFSBP_1%A_1163_48# N_A_1163_48#_M1001_s
+ N_A_1163_48#_M1038_d N_A_1163_48#_c_779_n N_A_1163_48#_M1005_g
+ N_A_1163_48#_c_780_n N_A_1163_48#_M1021_g N_A_1163_48#_c_781_n
+ N_A_1163_48#_c_782_n N_A_1163_48#_c_786_n N_A_1163_48#_c_787_n
+ N_A_1163_48#_c_783_n PM_SKY130_FD_SC_MS__SDFSBP_1%A_1163_48#
x_PM_SKY130_FD_SC_MS__SDFSBP_1%A_995_74# N_A_995_74#_M1037_d N_A_995_74#_M1022_d
+ N_A_995_74#_c_849_n N_A_995_74#_M1038_g N_A_995_74#_M1001_g
+ N_A_995_74#_M1041_g N_A_995_74#_c_853_n N_A_995_74#_M1024_g
+ N_A_995_74#_c_854_n N_A_995_74#_c_855_n N_A_995_74#_c_856_n
+ N_A_995_74#_c_857_n N_A_995_74#_c_858_n N_A_995_74#_c_865_n
+ N_A_995_74#_c_859_n N_A_995_74#_c_860_n N_A_995_74#_c_861_n
+ PM_SKY130_FD_SC_MS__SDFSBP_1%A_995_74#
x_PM_SKY130_FD_SC_MS__SDFSBP_1%SET_B N_SET_B_M1014_g N_SET_B_M1035_g
+ N_SET_B_c_979_n N_SET_B_M1012_g N_SET_B_c_980_n N_SET_B_c_981_n
+ N_SET_B_M1032_g N_SET_B_c_982_n N_SET_B_c_995_n N_SET_B_c_983_n
+ N_SET_B_c_984_n N_SET_B_c_985_n N_SET_B_c_986_n N_SET_B_c_987_n SET_B
+ N_SET_B_c_989_n N_SET_B_c_990_n N_SET_B_c_991_n
+ PM_SKY130_FD_SC_MS__SDFSBP_1%SET_B
x_PM_SKY130_FD_SC_MS__SDFSBP_1%A_594_74# N_A_594_74#_M1023_s N_A_594_74#_M1026_s
+ N_A_594_74#_c_1124_n N_A_594_74#_M1019_g N_A_594_74#_M1030_g
+ N_A_594_74#_c_1126_n N_A_594_74#_c_1127_n N_A_594_74#_c_1128_n
+ N_A_594_74#_c_1140_n N_A_594_74#_c_1141_n N_A_594_74#_M1037_g
+ N_A_594_74#_M1020_g N_A_594_74#_c_1143_n N_A_594_74#_M1003_g
+ N_A_594_74#_c_1131_n N_A_594_74#_M1008_g N_A_594_74#_c_1132_n
+ N_A_594_74#_c_1146_n N_A_594_74#_c_1133_n N_A_594_74#_c_1134_n
+ N_A_594_74#_c_1148_n N_A_594_74#_c_1149_n N_A_594_74#_c_1135_n
+ N_A_594_74#_c_1136_n N_A_594_74#_c_1137_n N_A_594_74#_c_1151_n
+ N_A_594_74#_c_1152_n PM_SKY130_FD_SC_MS__SDFSBP_1%A_594_74#
x_PM_SKY130_FD_SC_MS__SDFSBP_1%A_1924_48# N_A_1924_48#_M1006_d
+ N_A_1924_48#_M1029_s N_A_1924_48#_M1004_g N_A_1924_48#_c_1299_n
+ N_A_1924_48#_c_1312_n N_A_1924_48#_c_1313_n N_A_1924_48#_M1028_g
+ N_A_1924_48#_c_1300_n N_A_1924_48#_c_1301_n N_A_1924_48#_c_1302_n
+ N_A_1924_48#_c_1303_n N_A_1924_48#_c_1304_n N_A_1924_48#_c_1305_n
+ N_A_1924_48#_c_1306_n N_A_1924_48#_c_1307_n N_A_1924_48#_c_1315_n
+ N_A_1924_48#_c_1316_n N_A_1924_48#_c_1317_n N_A_1924_48#_c_1308_n
+ N_A_1924_48#_c_1345_n N_A_1924_48#_c_1309_n N_A_1924_48#_c_1310_n
+ PM_SKY130_FD_SC_MS__SDFSBP_1%A_1924_48#
x_PM_SKY130_FD_SC_MS__SDFSBP_1%A_1762_74# N_A_1762_74#_M1025_d
+ N_A_1762_74#_M1033_d N_A_1762_74#_M1032_d N_A_1762_74#_c_1428_n
+ N_A_1762_74#_M1006_g N_A_1762_74#_c_1429_n N_A_1762_74#_M1029_g
+ N_A_1762_74#_M1009_g N_A_1762_74#_c_1431_n N_A_1762_74#_c_1432_n
+ N_A_1762_74#_c_1446_n N_A_1762_74#_M1000_g N_A_1762_74#_c_1433_n
+ N_A_1762_74#_M1018_g N_A_1762_74#_c_1448_n N_A_1762_74#_M1034_g
+ N_A_1762_74#_c_1435_n N_A_1762_74#_c_1436_n N_A_1762_74#_c_1437_n
+ N_A_1762_74#_c_1438_n N_A_1762_74#_c_1439_n N_A_1762_74#_c_1453_n
+ N_A_1762_74#_c_1454_n N_A_1762_74#_c_1440_n N_A_1762_74#_c_1536_n
+ N_A_1762_74#_c_1441_n N_A_1762_74#_c_1456_n N_A_1762_74#_c_1442_n
+ N_A_1762_74#_c_1458_n N_A_1762_74#_c_1459_n N_A_1762_74#_c_1460_n
+ PM_SKY130_FD_SC_MS__SDFSBP_1%A_1762_74#
x_PM_SKY130_FD_SC_MS__SDFSBP_1%A_2556_112# N_A_2556_112#_M1018_s
+ N_A_2556_112#_M1034_s N_A_2556_112#_M1031_g N_A_2556_112#_c_1616_n
+ N_A_2556_112#_M1027_g N_A_2556_112#_c_1617_n N_A_2556_112#_c_1618_n
+ N_A_2556_112#_c_1619_n N_A_2556_112#_c_1620_n N_A_2556_112#_c_1621_n
+ PM_SKY130_FD_SC_MS__SDFSBP_1%A_2556_112#
x_PM_SKY130_FD_SC_MS__SDFSBP_1%VPWR N_VPWR_M1010_d N_VPWR_M1013_d N_VPWR_M1026_d
+ N_VPWR_M1021_d N_VPWR_M1035_d N_VPWR_M1028_d N_VPWR_M1029_d N_VPWR_M1034_d
+ N_VPWR_c_1663_n N_VPWR_c_1664_n N_VPWR_c_1665_n N_VPWR_c_1666_n
+ N_VPWR_c_1667_n N_VPWR_c_1668_n N_VPWR_c_1669_n N_VPWR_c_1670_n
+ N_VPWR_c_1671_n N_VPWR_c_1672_n N_VPWR_c_1673_n N_VPWR_c_1674_n
+ N_VPWR_c_1675_n N_VPWR_c_1676_n N_VPWR_c_1677_n VPWR N_VPWR_c_1678_n
+ N_VPWR_c_1679_n N_VPWR_c_1680_n N_VPWR_c_1681_n N_VPWR_c_1682_n
+ N_VPWR_c_1662_n N_VPWR_c_1684_n N_VPWR_c_1685_n N_VPWR_c_1686_n
+ N_VPWR_c_1687_n N_VPWR_c_1688_n PM_SKY130_FD_SC_MS__SDFSBP_1%VPWR
x_PM_SKY130_FD_SC_MS__SDFSBP_1%A_293_464# N_A_293_464#_M1040_d
+ N_A_293_464#_M1037_s N_A_293_464#_M1017_d N_A_293_464#_M1022_s
+ N_A_293_464#_c_1830_n N_A_293_464#_c_1818_n N_A_293_464#_c_1819_n
+ N_A_293_464#_c_1820_n N_A_293_464#_c_1845_n N_A_293_464#_c_1821_n
+ N_A_293_464#_c_1850_n N_A_293_464#_c_1825_n N_A_293_464#_c_1826_n
+ N_A_293_464#_c_1822_n N_A_293_464#_c_1828_n N_A_293_464#_c_1851_n
+ N_A_293_464#_c_1854_n N_A_293_464#_c_1914_n N_A_293_464#_c_1823_n
+ N_A_293_464#_c_1829_n PM_SKY130_FD_SC_MS__SDFSBP_1%A_293_464#
x_PM_SKY130_FD_SC_MS__SDFSBP_1%A_1603_347# N_A_1603_347#_M1041_d
+ N_A_1603_347#_M1008_d N_A_1603_347#_c_1946_n N_A_1603_347#_c_1947_n
+ N_A_1603_347#_c_1948_n PM_SKY130_FD_SC_MS__SDFSBP_1%A_1603_347#
x_PM_SKY130_FD_SC_MS__SDFSBP_1%A_1712_374# N_A_1712_374#_M1033_s
+ N_A_1712_374#_M1028_s N_A_1712_374#_c_1980_n N_A_1712_374#_c_1981_n
+ N_A_1712_374#_c_1982_n PM_SKY130_FD_SC_MS__SDFSBP_1%A_1712_374#
x_PM_SKY130_FD_SC_MS__SDFSBP_1%Q_N N_Q_N_M1009_d N_Q_N_M1000_d N_Q_N_c_2014_n
+ N_Q_N_c_2015_n N_Q_N_c_2011_n Q_N Q_N Q_N PM_SKY130_FD_SC_MS__SDFSBP_1%Q_N
x_PM_SKY130_FD_SC_MS__SDFSBP_1%Q N_Q_M1027_d N_Q_M1031_d Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_MS__SDFSBP_1%Q
x_PM_SKY130_FD_SC_MS__SDFSBP_1%VGND N_VGND_M1036_d N_VGND_M1016_d N_VGND_M1023_d
+ N_VGND_M1005_d N_VGND_M1014_d N_VGND_M1012_d N_VGND_M1009_s N_VGND_M1018_d
+ N_VGND_c_2059_n N_VGND_c_2060_n N_VGND_c_2061_n N_VGND_c_2062_n
+ N_VGND_c_2063_n N_VGND_c_2064_n N_VGND_c_2065_n N_VGND_c_2066_n
+ N_VGND_c_2067_n N_VGND_c_2068_n VGND N_VGND_c_2069_n N_VGND_c_2070_n
+ N_VGND_c_2071_n N_VGND_c_2072_n N_VGND_c_2073_n N_VGND_c_2074_n
+ N_VGND_c_2075_n N_VGND_c_2076_n N_VGND_c_2077_n N_VGND_c_2078_n
+ N_VGND_c_2079_n N_VGND_c_2080_n N_VGND_c_2081_n N_VGND_c_2082_n
+ PM_SKY130_FD_SC_MS__SDFSBP_1%VGND
cc_1 VNB N_SCE_M1036_g 0.0641507f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_2 VNB N_SCE_M1015_g 0.035064f $X=-0.19 $Y=-0.245 $X2=1.885 $Y2=0.58
cc_3 VNB N_SCE_c_296_n 0.0234769f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.535
cc_4 VNB N_SCE_c_297_n 0.00280342f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.425
cc_5 VNB N_SCE_c_298_n 0.0318809f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.425
cc_6 VNB N_SCE_c_299_n 0.0201092f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.685
cc_7 VNB N_SCE_c_300_n 0.00254062f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.535
cc_8 VNB N_A_27_74#_M1039_g 0.0215636f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.18
cc_9 VNB N_A_27_74#_c_372_n 0.0260478f $X=-0.19 $Y=-0.245 $X2=1.885 $Y2=0.58
cc_10 VNB N_A_27_74#_c_373_n 0.0186355f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.535
cc_11 VNB N_A_27_74#_c_374_n 0.0084149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_c_375_n 0.0327363f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.685
cc_13 VNB N_A_27_74#_c_376_n 0.0182839f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.26
cc_14 VNB N_D_M1040_g 0.062081f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_15 VNB N_SCD_c_495_n 0.0176451f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.85
cc_16 VNB N_SCD_c_496_n 0.0589035f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_17 VNB N_SCD_c_497_n 0.0257799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB SCD 0.00577239f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.18
cc_19 VNB N_CLK_c_539_n 0.0191493f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.85
cc_20 VNB N_CLK_c_540_n 0.0431373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB CLK 0.00704257f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_22 VNB N_A_781_74#_M1007_g 0.0623484f $X=-0.19 $Y=-0.245 $X2=1.885 $Y2=1.26
cc_23 VNB N_A_781_74#_M1025_g 0.0315835f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.09
cc_24 VNB N_A_781_74#_c_574_n 0.00580499f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.535
cc_25 VNB N_A_781_74#_c_575_n 0.0155903f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.685
cc_26 VNB N_A_781_74#_c_576_n 0.00279267f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.685
cc_27 VNB N_A_781_74#_c_577_n 0.0011848f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.425
cc_28 VNB N_A_781_74#_c_578_n 0.0279286f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.535
cc_29 VNB N_A_781_74#_c_579_n 0.00602655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_781_74#_c_580_n 0.00206749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_781_74#_c_581_n 0.0289981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_1163_48#_c_779_n 0.0183276f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_33 VNB N_A_1163_48#_c_780_n 0.00595723f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.64
cc_34 VNB N_A_1163_48#_c_781_n 0.0254327f $X=-0.19 $Y=-0.245 $X2=1.885 $Y2=1.26
cc_35 VNB N_A_1163_48#_c_782_n 0.0220946f $X=-0.19 $Y=-0.245 $X2=1.885 $Y2=0.58
cc_36 VNB N_A_1163_48#_c_783_n 0.0607898f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.685
cc_37 VNB N_A_995_74#_c_849_n 0.0386116f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_38 VNB N_A_995_74#_M1038_g 0.00326225f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.18
cc_39 VNB N_A_995_74#_M1001_g 0.0341535f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.85
cc_40 VNB N_A_995_74#_M1041_g 0.00682949f $X=-0.19 $Y=-0.245 $X2=1.885 $Y2=0.58
cc_41 VNB N_A_995_74#_c_853_n 0.0189909f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.09
cc_42 VNB N_A_995_74#_c_854_n 0.00687291f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.425
cc_43 VNB N_A_995_74#_c_855_n 0.00207814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_995_74#_c_856_n 0.0252332f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_45 VNB N_A_995_74#_c_857_n 0.0198101f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.685
cc_46 VNB N_A_995_74#_c_858_n 0.00264222f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.685
cc_47 VNB N_A_995_74#_c_859_n 0.00350923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_995_74#_c_860_n 0.0124973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_995_74#_c_861_n 0.0577977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_SET_B_M1014_g 0.0406873f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.64
cc_51 VNB N_SET_B_M1035_g 0.00252704f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_52 VNB N_SET_B_c_979_n 0.018015f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.18
cc_53 VNB N_SET_B_c_980_n 0.0242576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_SET_B_c_981_n 0.00843777f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.85
cc_55 VNB N_SET_B_c_982_n 0.0174838f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.425
cc_56 VNB N_SET_B_c_983_n 0.00206835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_SET_B_c_984_n 0.0249121f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.535
cc_58 VNB N_SET_B_c_985_n 0.00828735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_SET_B_c_986_n 0.0184503f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.685
cc_60 VNB N_SET_B_c_987_n 0.00180662f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.685
cc_61 VNB SET_B 0.00199056f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.26
cc_62 VNB N_SET_B_c_989_n 0.0274525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_SET_B_c_990_n 0.00167402f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.665
cc_64 VNB N_SET_B_c_991_n 0.0163976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_594_74#_c_1124_n 0.0206133f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_66 VNB N_A_594_74#_M1030_g 0.00599386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_594_74#_c_1126_n 0.0266552f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.09
cc_68 VNB N_A_594_74#_c_1127_n 0.00499256f $X=-0.19 $Y=-0.245 $X2=1.885 $Y2=0.58
cc_69 VNB N_A_594_74#_c_1128_n 0.028937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_594_74#_M1037_g 0.0243464f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.425
cc_71 VNB N_A_594_74#_M1003_g 0.0562556f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.685
cc_72 VNB N_A_594_74#_c_1131_n 0.00600082f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.425
cc_73 VNB N_A_594_74#_c_1132_n 0.0256095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_594_74#_c_1133_n 0.00880724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_594_74#_c_1134_n 0.0115805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_594_74#_c_1135_n 0.00306961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_594_74#_c_1136_n 0.0201562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_594_74#_c_1137_n 0.0016464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1924_48#_c_1299_n 0.0161449f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.64
cc_80 VNB N_A_1924_48#_c_1300_n 0.0183699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1924_48#_c_1301_n 0.0165713f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.09
cc_82 VNB N_A_1924_48#_c_1302_n 0.0230002f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=1.425
cc_83 VNB N_A_1924_48#_c_1303_n 0.0243895f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.425
cc_84 VNB N_A_1924_48#_c_1304_n 0.007537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1924_48#_c_1305_n 0.00286542f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.685
cc_86 VNB N_A_1924_48#_c_1306_n 0.02238f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.685
cc_87 VNB N_A_1924_48#_c_1307_n 0.00154245f $X=-0.19 $Y=-0.245 $X2=0.67
+ $Y2=1.685
cc_88 VNB N_A_1924_48#_c_1308_n 0.00143741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1924_48#_c_1309_n 0.0181664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1924_48#_c_1310_n 0.00510964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1762_74#_c_1428_n 0.0200354f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.64
cc_92 VNB N_A_1762_74#_c_1429_n 0.0358613f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=2.09
cc_93 VNB N_A_1762_74#_M1009_g 0.0507407f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.535
cc_94 VNB N_A_1762_74#_c_1431_n 0.00282799f $X=-0.19 $Y=-0.245 $X2=1.96
+ $Y2=1.425
cc_95 VNB N_A_1762_74#_c_1432_n 0.00451186f $X=-0.19 $Y=-0.245 $X2=1.96
+ $Y2=1.425
cc_96 VNB N_A_1762_74#_c_1433_n 0.0207444f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_97 VNB N_A_1762_74#_M1018_g 0.0436388f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.685
cc_98 VNB N_A_1762_74#_c_1435_n 0.0283734f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.535
cc_99 VNB N_A_1762_74#_c_1436_n 0.00147097f $X=-0.19 $Y=-0.245 $X2=0.67
+ $Y2=1.665
cc_100 VNB N_A_1762_74#_c_1437_n 0.0100433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1762_74#_c_1438_n 0.00658164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1762_74#_c_1439_n 0.00171038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1762_74#_c_1440_n 0.00153994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1762_74#_c_1441_n 0.00938966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1762_74#_c_1442_n 0.00483919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_2556_112#_M1031_g 0.00835878f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.18
cc_107 VNB N_A_2556_112#_c_1616_n 0.023668f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.64
cc_108 VNB N_A_2556_112#_c_1617_n 0.0359811f $X=-0.19 $Y=-0.245 $X2=0.97
+ $Y2=2.09
cc_109 VNB N_A_2556_112#_c_1618_n 0.017119f $X=-0.19 $Y=-0.245 $X2=1.885
+ $Y2=1.26
cc_110 VNB N_A_2556_112#_c_1619_n 0.0138984f $X=-0.19 $Y=-0.245 $X2=1.885
+ $Y2=0.58
cc_111 VNB N_A_2556_112#_c_1620_n 0.0023636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_2556_112#_c_1621_n 0.0096015f $X=-0.19 $Y=-0.245 $X2=1.92
+ $Y2=1.425
cc_113 VNB N_VPWR_c_1662_n 0.601534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_293_464#_c_1818_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.09
cc_115 VNB N_A_293_464#_c_1819_n 0.0125835f $X=-0.19 $Y=-0.245 $X2=0.835
+ $Y2=1.535
cc_116 VNB N_A_293_464#_c_1820_n 0.0033344f $X=-0.19 $Y=-0.245 $X2=1.92
+ $Y2=1.425
cc_117 VNB N_A_293_464#_c_1821_n 0.0044818f $X=-0.19 $Y=-0.245 $X2=1.92
+ $Y2=1.535
cc_118 VNB N_A_293_464#_c_1822_n 0.00566544f $X=-0.19 $Y=-0.245 $X2=0.67
+ $Y2=1.685
cc_119 VNB N_A_293_464#_c_1823_n 0.00460204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_Q_N_c_2011_n 0.0103864f $X=-0.19 $Y=-0.245 $X2=1.885 $Y2=1.26
cc_121 VNB Q_N 0.0150197f $X=-0.19 $Y=-0.245 $X2=1.885 $Y2=0.58
cc_122 VNB Q_N 0.00781016f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_123 VNB Q 0.0547356f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_124 VNB N_VGND_c_2059_n 0.00982527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2060_n 0.0109164f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.685
cc_126 VNB N_VGND_c_2061_n 0.00600048f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.85
cc_127 VNB N_VGND_c_2062_n 0.0120969f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.535
cc_128 VNB N_VGND_c_2063_n 0.0194709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2064_n 0.0169908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2065_n 0.0411304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2066_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2067_n 0.0596655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2068_n 0.00670466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2069_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2070_n 0.0207541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2071_n 0.0583309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2072_n 0.0206359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2073_n 0.0415877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2074_n 0.0191124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2075_n 0.816858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2076_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2077_n 0.00615422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2078_n 0.0324822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2079_n 0.0266754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2080_n 0.0210309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2081_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2082_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VPB N_SCE_M1010_g 0.0431562f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_149 VPB N_SCE_c_302_n 0.00575706f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.18
cc_150 VPB N_SCE_M1011_g 0.019465f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_151 VPB N_SCE_c_304_n 0.0119787f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.09
cc_152 VPB N_SCE_c_299_n 0.0291714f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.685
cc_153 VPB N_SCE_c_300_n 0.00166152f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.535
cc_154 VPB N_A_27_74#_M1002_g 0.0228664f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.85
cc_155 VPB N_A_27_74#_c_373_n 0.0318728f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.535
cc_156 VPB N_A_27_74#_c_379_n 0.0214642f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.425
cc_157 VPB N_A_27_74#_c_380_n 0.0116291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_27_74#_c_381_n 0.00316303f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.685
cc_159 VPB N_A_27_74#_c_382_n 0.0317113f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.85
cc_160 VPB N_A_27_74#_c_383_n 0.00834358f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_D_M1017_g 0.0257642f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_162 VPB N_D_M1040_g 0.00913433f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_163 VPB N_D_c_459_n 0.0272462f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_D_c_460_n 0.00879535f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.85
cc_165 VPB N_SCD_c_499_n 0.0573101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_SCD_c_497_n 0.0258202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB SCD 0.00195322f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.18
cc_168 VPB N_CLK_c_540_n 0.0266307f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_781_74#_M1022_g 0.0281209f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.18
cc_170 VPB N_A_781_74#_M1007_g 0.00176557f $X=-0.19 $Y=1.66 $X2=1.885 $Y2=1.26
cc_171 VPB N_A_781_74#_c_584_n 0.0032477f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.685
cc_172 VPB N_A_781_74#_c_585_n 0.0226421f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.685
cc_173 VPB N_A_781_74#_c_586_n 0.00299508f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.85
cc_174 VPB N_A_781_74#_c_587_n 0.0012556f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_781_74#_c_578_n 0.0288218f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.535
cc_176 VPB N_A_781_74#_c_589_n 0.00866173f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_781_74#_c_590_n 0.00150794f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_781_74#_c_591_n 0.0232105f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_781_74#_c_592_n 0.00242474f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_781_74#_c_593_n 0.0156765f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_781_74#_c_594_n 0.00177503f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_781_74#_c_595_n 0.00330131f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_781_74#_c_596_n 0.0108876f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_781_74#_c_597_n 0.00198955f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_781_74#_c_598_n 0.00108929f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_781_74#_c_599_n 0.0367844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_781_74#_c_581_n 0.0146427f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_781_74#_c_601_n 0.0209911f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_781_74#_c_602_n 0.0178597f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_1163_48#_c_780_n 0.026024f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_191 VPB N_A_1163_48#_M1021_g 0.034101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_1163_48#_c_786_n 0.0122379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_1163_48#_c_787_n 0.00791538f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_995_74#_M1038_g 0.0502092f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.18
cc_195 VPB N_A_995_74#_M1041_g 0.0232564f $X=-0.19 $Y=1.66 $X2=1.885 $Y2=0.58
cc_196 VPB N_A_995_74#_c_855_n 0.00921227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_995_74#_c_865_n 5.32349e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_SET_B_M1035_g 0.0496257f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_199 VPB N_SET_B_M1032_g 0.0572638f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.535
cc_200 VPB N_SET_B_c_982_n 0.00938523f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.425
cc_201 VPB N_SET_B_c_995_n 0.0223199f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.425
cc_202 VPB N_SET_B_c_983_n 0.00200906f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_SET_B_c_985_n 0.00616409f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_SET_B_c_986_n 0.0153051f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.685
cc_205 VPB N_SET_B_c_987_n 0.00200016f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.685
cc_206 VPB SET_B 0.00172634f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.26
cc_207 VPB N_SET_B_c_989_n 0.00506136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_SET_B_c_990_n 0.00239196f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.665
cc_209 VPB N_A_594_74#_M1030_g 0.0221109f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_594_74#_c_1127_n 0.0728015f $X=-0.19 $Y=1.66 $X2=1.885 $Y2=0.58
cc_211 VPB N_A_594_74#_c_1140_n 0.0625467f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.535
cc_212 VPB N_A_594_74#_c_1141_n 0.0123627f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.535
cc_213 VPB N_A_594_74#_M1020_g 0.030534f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_214 VPB N_A_594_74#_c_1143_n 0.288291f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.685
cc_215 VPB N_A_594_74#_c_1131_n 0.0118122f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.425
cc_216 VPB N_A_594_74#_M1008_g 0.0197016f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.535
cc_217 VPB N_A_594_74#_c_1146_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_594_74#_c_1134_n 0.00354716f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_594_74#_c_1148_n 0.00550874f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_594_74#_c_1149_n 0.00417741f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_594_74#_c_1135_n 0.00103128f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_594_74#_c_1151_n 0.00585197f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_594_74#_c_1152_n 9.87779e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_1924_48#_c_1299_n 0.0310005f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_225 VPB N_A_1924_48#_c_1312_n 0.0317698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_1924_48#_c_1313_n 0.011056f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.85
cc_227 VPB N_A_1924_48#_M1028_g 0.0298912f $X=-0.19 $Y=1.66 $X2=1.885 $Y2=0.58
cc_228 VPB N_A_1924_48#_c_1315_n 0.0103903f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.85
cc_229 VPB N_A_1924_48#_c_1316_n 0.00493064f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.26
cc_230 VPB N_A_1924_48#_c_1317_n 0.00379531f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_1924_48#_c_1308_n 9.08496e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_1762_74#_M1029_g 0.0435597f $X=-0.19 $Y=1.66 $X2=1.885 $Y2=0.58
cc_233 VPB N_A_1762_74#_c_1431_n 0.00353145f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.425
cc_234 VPB N_A_1762_74#_c_1432_n 0.0237496f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.425
cc_235 VPB N_A_1762_74#_c_1446_n 0.0212431f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_1762_74#_c_1433_n 0.0281658f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_237 VPB N_A_1762_74#_c_1448_n 0.0177468f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.685
cc_238 VPB N_A_1762_74#_c_1436_n 0.0155417f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.665
cc_239 VPB N_A_1762_74#_c_1437_n 0.0280916f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_A_1762_74#_c_1438_n 0.00200584f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_A_1762_74#_c_1439_n 0.0334023f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_A_1762_74#_c_1453_n 0.00241768f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_1762_74#_c_1454_n 0.0173499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_A_1762_74#_c_1440_n 0.00744762f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_1762_74#_c_1456_n 0.00198749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_A_1762_74#_c_1442_n 9.77533e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_1762_74#_c_1458_n 0.00354986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_A_1762_74#_c_1459_n 0.0078305f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_A_1762_74#_c_1460_n 0.00546427f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_A_2556_112#_M1031_g 0.0305596f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.18
cc_251 VPB N_A_2556_112#_c_1620_n 0.0158606f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1663_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1664_n 0.00988271f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.685
cc_254 VPB N_VPWR_c_1665_n 0.023804f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.685
cc_255 VPB N_VPWR_c_1666_n 0.00396467f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.26
cc_256 VPB N_VPWR_c_1667_n 0.00550557f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.665
cc_257 VPB N_VPWR_c_1668_n 0.012458f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1669_n 0.00951764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1670_n 0.0070628f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1671_n 0.0115238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1672_n 0.0546335f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1673_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1674_n 0.027717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1675_n 0.00223798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1676_n 0.0685213f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1677_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1678_n 0.0180274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1679_n 0.0463631f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1680_n 0.0334651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1681_n 0.0337745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1682_n 0.0191124f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1662_n 0.130846f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1684_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1685_n 0.00507132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1686_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1687_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1688_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_A_293_464#_c_1821_n 0.00530109f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=1.535
cc_279 VPB N_A_293_464#_c_1825_n 0.0131901f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_A_293_464#_c_1826_n 0.00351062f $X=-0.19 $Y=1.66 $X2=0.505
+ $Y2=1.685
cc_281 VPB N_A_293_464#_c_1822_n 0.00402833f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.685
cc_282 VPB N_A_293_464#_c_1828_n 0.00464321f $X=-0.19 $Y=1.66 $X2=1.96 $Y2=1.26
cc_283 VPB N_A_293_464#_c_1829_n 0.00812315f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_284 VPB N_A_1603_347#_c_1946_n 0.011327f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_285 VPB N_A_1603_347#_c_1947_n 0.0114218f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.18
cc_286 VPB N_A_1603_347#_c_1948_n 0.00549831f $X=-0.19 $Y=1.66 $X2=1.885
+ $Y2=0.58
cc_287 VPB N_A_1712_374#_c_1980_n 0.0261465f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_288 VPB N_A_1712_374#_c_1981_n 0.00663462f $X=-0.19 $Y=1.66 $X2=0.955
+ $Y2=2.64
cc_289 VPB N_A_1712_374#_c_1982_n 0.0164293f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=2.09
cc_290 VPB N_Q_N_c_2014_n 0.00106684f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.18
cc_291 VPB N_Q_N_c_2015_n 0.00220173f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.64
cc_292 VPB N_Q_N_c_2011_n 5.04282e-19 $X=-0.19 $Y=1.66 $X2=1.885 $Y2=1.26
cc_293 VPB Q 0.0537246f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_294 N_SCE_M1036_g N_A_27_74#_M1039_g 0.0154087f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_295 N_SCE_M1036_g N_A_27_74#_c_372_n 0.0123507f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_296 N_SCE_M1036_g N_A_27_74#_c_373_n 0.00803467f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_297 N_SCE_c_299_n N_A_27_74#_c_373_n 0.0264823f $X=0.67 $Y=1.685 $X2=0 $Y2=0
cc_298 N_SCE_c_300_n N_A_27_74#_c_373_n 0.030623f $X=0.67 $Y=1.535 $X2=0 $Y2=0
cc_299 N_SCE_M1010_g N_A_27_74#_c_379_n 4.69176e-19 $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_300 N_SCE_M1010_g N_A_27_74#_c_380_n 0.0182123f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_301 N_SCE_M1011_g N_A_27_74#_c_380_n 0.0179896f $X=0.955 $Y=2.64 $X2=0 $Y2=0
cc_302 N_SCE_c_296_n N_A_27_74#_c_380_n 0.0125499f $X=1.795 $Y=1.535 $X2=0 $Y2=0
cc_303 N_SCE_c_299_n N_A_27_74#_c_380_n 6.8039e-19 $X=0.67 $Y=1.685 $X2=0 $Y2=0
cc_304 N_SCE_c_300_n N_A_27_74#_c_380_n 0.011957f $X=0.67 $Y=1.535 $X2=0 $Y2=0
cc_305 N_SCE_M1036_g N_A_27_74#_c_374_n 0.0168544f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_306 N_SCE_c_296_n N_A_27_74#_c_374_n 0.0229228f $X=1.795 $Y=1.535 $X2=0 $Y2=0
cc_307 N_SCE_c_297_n N_A_27_74#_c_374_n 4.79392e-19 $X=1.96 $Y=1.425 $X2=0 $Y2=0
cc_308 N_SCE_c_299_n N_A_27_74#_c_374_n 0.0014947f $X=0.67 $Y=1.685 $X2=0 $Y2=0
cc_309 N_SCE_c_300_n N_A_27_74#_c_374_n 0.0272074f $X=0.67 $Y=1.535 $X2=0 $Y2=0
cc_310 N_SCE_M1036_g N_A_27_74#_c_375_n 0.0180926f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_311 N_SCE_c_296_n N_A_27_74#_c_375_n 0.00422079f $X=1.795 $Y=1.535 $X2=0
+ $Y2=0
cc_312 N_SCE_c_299_n N_A_27_74#_c_375_n 0.00630445f $X=0.67 $Y=1.685 $X2=0 $Y2=0
cc_313 N_SCE_c_297_n N_A_27_74#_c_381_n 0.0178307f $X=1.96 $Y=1.425 $X2=0 $Y2=0
cc_314 N_SCE_c_298_n N_A_27_74#_c_381_n 2.95197e-19 $X=1.96 $Y=1.425 $X2=0 $Y2=0
cc_315 N_SCE_c_297_n N_A_27_74#_c_382_n 8.97175e-19 $X=1.96 $Y=1.425 $X2=0 $Y2=0
cc_316 N_SCE_c_298_n N_A_27_74#_c_382_n 0.019309f $X=1.96 $Y=1.425 $X2=0 $Y2=0
cc_317 N_SCE_M1036_g N_A_27_74#_c_376_n 0.00874187f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_318 N_SCE_c_299_n N_A_27_74#_c_376_n 2.24402e-19 $X=0.67 $Y=1.685 $X2=0 $Y2=0
cc_319 N_SCE_c_302_n N_D_M1017_g 0.053471f $X=0.955 $Y=2.18 $X2=0 $Y2=0
cc_320 N_SCE_M1015_g N_D_M1040_g 0.0289627f $X=1.885 $Y=0.58 $X2=0 $Y2=0
cc_321 N_SCE_c_296_n N_D_M1040_g 0.0159859f $X=1.795 $Y=1.535 $X2=0 $Y2=0
cc_322 N_SCE_c_297_n N_D_M1040_g 0.00137327f $X=1.96 $Y=1.425 $X2=0 $Y2=0
cc_323 N_SCE_c_298_n N_D_M1040_g 0.0163018f $X=1.96 $Y=1.425 $X2=0 $Y2=0
cc_324 N_SCE_c_299_n N_D_M1040_g 0.00756384f $X=0.67 $Y=1.685 $X2=0 $Y2=0
cc_325 N_SCE_c_300_n N_D_M1040_g 9.94783e-19 $X=0.67 $Y=1.535 $X2=0 $Y2=0
cc_326 N_SCE_c_296_n N_D_c_459_n 0.00440999f $X=1.795 $Y=1.535 $X2=0 $Y2=0
cc_327 N_SCE_c_299_n N_D_c_459_n 0.0196439f $X=0.67 $Y=1.685 $X2=0 $Y2=0
cc_328 N_SCE_c_296_n N_D_c_460_n 0.0377186f $X=1.795 $Y=1.535 $X2=0 $Y2=0
cc_329 N_SCE_c_299_n N_D_c_460_n 0.0083863f $X=0.67 $Y=1.685 $X2=0 $Y2=0
cc_330 N_SCE_c_300_n N_D_c_460_n 0.00363459f $X=0.67 $Y=1.535 $X2=0 $Y2=0
cc_331 N_SCE_M1015_g N_SCD_c_495_n 0.0397201f $X=1.885 $Y=0.58 $X2=-0.19
+ $Y2=-0.245
cc_332 N_SCE_M1015_g N_SCD_c_496_n 0.00623104f $X=1.885 $Y=0.58 $X2=0 $Y2=0
cc_333 N_SCE_c_297_n N_SCD_c_496_n 2.80393e-19 $X=1.96 $Y=1.425 $X2=0 $Y2=0
cc_334 N_SCE_c_298_n N_SCD_c_496_n 0.0171993f $X=1.96 $Y=1.425 $X2=0 $Y2=0
cc_335 N_SCE_M1010_g N_VPWR_c_1663_n 0.0116339f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_336 N_SCE_M1011_g N_VPWR_c_1663_n 0.0110385f $X=0.955 $Y=2.64 $X2=0 $Y2=0
cc_337 N_SCE_M1010_g N_VPWR_c_1678_n 0.00460063f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_338 N_SCE_M1011_g N_VPWR_c_1679_n 0.00460063f $X=0.955 $Y=2.64 $X2=0 $Y2=0
cc_339 N_SCE_M1010_g N_VPWR_c_1662_n 0.00912296f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_340 N_SCE_M1011_g N_VPWR_c_1662_n 0.00908371f $X=0.955 $Y=2.64 $X2=0 $Y2=0
cc_341 N_SCE_M1011_g N_A_293_464#_c_1830_n 9.27257e-19 $X=0.955 $Y=2.64 $X2=0
+ $Y2=0
cc_342 N_SCE_M1015_g N_A_293_464#_c_1818_n 0.0119647f $X=1.885 $Y=0.58 $X2=0
+ $Y2=0
cc_343 N_SCE_M1015_g N_A_293_464#_c_1819_n 0.0112369f $X=1.885 $Y=0.58 $X2=0
+ $Y2=0
cc_344 N_SCE_c_297_n N_A_293_464#_c_1819_n 0.0153887f $X=1.96 $Y=1.425 $X2=0
+ $Y2=0
cc_345 N_SCE_c_298_n N_A_293_464#_c_1819_n 0.00363502f $X=1.96 $Y=1.425 $X2=0
+ $Y2=0
cc_346 N_SCE_M1015_g N_A_293_464#_c_1820_n 0.00274486f $X=1.885 $Y=0.58 $X2=0
+ $Y2=0
cc_347 N_SCE_c_296_n N_A_293_464#_c_1820_n 0.0143345f $X=1.795 $Y=1.535 $X2=0
+ $Y2=0
cc_348 N_SCE_c_297_n N_A_293_464#_c_1820_n 0.00321217f $X=1.96 $Y=1.425 $X2=0
+ $Y2=0
cc_349 N_SCE_M1015_g N_A_293_464#_c_1821_n 0.00333921f $X=1.885 $Y=0.58 $X2=0
+ $Y2=0
cc_350 N_SCE_c_297_n N_A_293_464#_c_1821_n 0.0266104f $X=1.96 $Y=1.425 $X2=0
+ $Y2=0
cc_351 N_SCE_c_298_n N_A_293_464#_c_1821_n 0.00220024f $X=1.96 $Y=1.425 $X2=0
+ $Y2=0
cc_352 N_SCE_M1036_g N_VGND_c_2059_n 0.00586161f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_353 N_SCE_M1015_g N_VGND_c_2060_n 0.00169331f $X=1.885 $Y=0.58 $X2=0 $Y2=0
cc_354 N_SCE_M1015_g N_VGND_c_2065_n 0.00434272f $X=1.885 $Y=0.58 $X2=0 $Y2=0
cc_355 N_SCE_M1036_g N_VGND_c_2069_n 0.00434272f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_356 N_SCE_M1036_g N_VGND_c_2075_n 0.0082497f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_357 N_SCE_M1015_g N_VGND_c_2075_n 0.00821077f $X=1.885 $Y=0.58 $X2=0 $Y2=0
cc_358 N_A_27_74#_M1002_g N_D_M1017_g 0.024517f $X=2.005 $Y=2.64 $X2=0 $Y2=0
cc_359 N_A_27_74#_c_380_n N_D_M1017_g 0.0166166f $X=1.795 $Y=2.375 $X2=0 $Y2=0
cc_360 N_A_27_74#_c_381_n N_D_M1017_g 0.00281475f $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_361 N_A_27_74#_c_382_n N_D_M1017_g 0.00160977f $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_362 N_A_27_74#_M1039_g N_D_M1040_g 0.0528466f $X=1.065 $Y=0.58 $X2=0 $Y2=0
cc_363 N_A_27_74#_c_374_n N_D_M1040_g 0.0016481f $X=0.975 $Y=1.115 $X2=0 $Y2=0
cc_364 N_A_27_74#_c_380_n N_D_c_459_n 0.00361918f $X=1.795 $Y=2.375 $X2=0 $Y2=0
cc_365 N_A_27_74#_c_381_n N_D_c_459_n 3.66318e-19 $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_366 N_A_27_74#_c_382_n N_D_c_459_n 0.0182533f $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_367 N_A_27_74#_c_380_n N_D_c_460_n 0.0376063f $X=1.795 $Y=2.375 $X2=0 $Y2=0
cc_368 N_A_27_74#_c_381_n N_D_c_460_n 0.018611f $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_369 N_A_27_74#_c_382_n N_D_c_460_n 0.00100613f $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_370 N_A_27_74#_M1002_g N_SCD_c_499_n 0.0481726f $X=2.005 $Y=2.64 $X2=0 $Y2=0
cc_371 N_A_27_74#_c_382_n N_SCD_c_499_n 6.16971e-19 $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_372 N_A_27_74#_c_381_n N_SCD_c_497_n 2.71882e-19 $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_373 N_A_27_74#_c_382_n N_SCD_c_497_n 0.0166773f $X=1.96 $Y=1.995 $X2=0 $Y2=0
cc_374 N_A_27_74#_c_380_n N_VPWR_M1010_d 0.00165831f $X=1.795 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_375 N_A_27_74#_c_379_n N_VPWR_c_1663_n 0.0122069f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_376 N_A_27_74#_c_380_n N_VPWR_c_1663_n 0.0170259f $X=1.795 $Y=2.375 $X2=0
+ $Y2=0
cc_377 N_A_27_74#_c_379_n N_VPWR_c_1678_n 0.0110674f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_378 N_A_27_74#_M1002_g N_VPWR_c_1679_n 0.00373242f $X=2.005 $Y=2.64 $X2=0
+ $Y2=0
cc_379 N_A_27_74#_M1002_g N_VPWR_c_1662_n 0.0046177f $X=2.005 $Y=2.64 $X2=0
+ $Y2=0
cc_380 N_A_27_74#_c_379_n N_VPWR_c_1662_n 0.00916f $X=0.28 $Y=2.465 $X2=0 $Y2=0
cc_381 N_A_27_74#_c_380_n A_209_464# 0.0048076f $X=1.795 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_382 N_A_27_74#_c_380_n N_A_293_464#_M1017_d 0.00417746f $X=1.795 $Y=2.375
+ $X2=0 $Y2=0
cc_383 N_A_27_74#_c_380_n N_A_293_464#_c_1830_n 0.0229291f $X=1.795 $Y=2.375
+ $X2=0 $Y2=0
cc_384 N_A_27_74#_M1039_g N_A_293_464#_c_1818_n 0.00194947f $X=1.065 $Y=0.58
+ $X2=0 $Y2=0
cc_385 N_A_27_74#_c_374_n N_A_293_464#_c_1820_n 0.00633768f $X=0.975 $Y=1.115
+ $X2=0 $Y2=0
cc_386 N_A_27_74#_M1002_g N_A_293_464#_c_1845_n 0.0102664f $X=2.005 $Y=2.64
+ $X2=0 $Y2=0
cc_387 N_A_27_74#_M1002_g N_A_293_464#_c_1821_n 9.17734e-19 $X=2.005 $Y=2.64
+ $X2=0 $Y2=0
cc_388 N_A_27_74#_c_380_n N_A_293_464#_c_1821_n 0.00235954f $X=1.795 $Y=2.375
+ $X2=0 $Y2=0
cc_389 N_A_27_74#_c_381_n N_A_293_464#_c_1821_n 0.033778f $X=1.96 $Y=1.995 $X2=0
+ $Y2=0
cc_390 N_A_27_74#_c_382_n N_A_293_464#_c_1821_n 0.00219558f $X=1.96 $Y=1.995
+ $X2=0 $Y2=0
cc_391 N_A_27_74#_M1002_g N_A_293_464#_c_1850_n 0.0029949f $X=2.005 $Y=2.64
+ $X2=0 $Y2=0
cc_392 N_A_27_74#_M1002_g N_A_293_464#_c_1851_n 0.00979234f $X=2.005 $Y=2.64
+ $X2=0 $Y2=0
cc_393 N_A_27_74#_c_380_n N_A_293_464#_c_1851_n 0.0152073f $X=1.795 $Y=2.375
+ $X2=0 $Y2=0
cc_394 N_A_27_74#_c_382_n N_A_293_464#_c_1851_n 3.76263e-19 $X=1.96 $Y=1.995
+ $X2=0 $Y2=0
cc_395 N_A_27_74#_M1002_g N_A_293_464#_c_1854_n 0.00180583f $X=2.005 $Y=2.64
+ $X2=0 $Y2=0
cc_396 N_A_27_74#_c_380_n N_A_293_464#_c_1854_n 0.0122365f $X=1.795 $Y=2.375
+ $X2=0 $Y2=0
cc_397 N_A_27_74#_M1039_g N_VGND_c_2059_n 0.00597281f $X=1.065 $Y=0.58 $X2=0
+ $Y2=0
cc_398 N_A_27_74#_c_372_n N_VGND_c_2059_n 0.0169251f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_399 N_A_27_74#_c_374_n N_VGND_c_2059_n 0.0268964f $X=0.975 $Y=1.115 $X2=0
+ $Y2=0
cc_400 N_A_27_74#_c_375_n N_VGND_c_2059_n 0.0030881f $X=0.975 $Y=1.115 $X2=0
+ $Y2=0
cc_401 N_A_27_74#_M1039_g N_VGND_c_2065_n 0.00461464f $X=1.065 $Y=0.58 $X2=0
+ $Y2=0
cc_402 N_A_27_74#_c_372_n N_VGND_c_2069_n 0.0145639f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_403 N_A_27_74#_M1039_g N_VGND_c_2075_n 0.00909071f $X=1.065 $Y=0.58 $X2=0
+ $Y2=0
cc_404 N_A_27_74#_c_372_n N_VGND_c_2075_n 0.0119984f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_405 N_D_M1017_g N_VPWR_c_1663_n 0.00157859f $X=1.375 $Y=2.64 $X2=0 $Y2=0
cc_406 N_D_M1017_g N_VPWR_c_1679_n 0.00520332f $X=1.375 $Y=2.64 $X2=0 $Y2=0
cc_407 N_D_M1017_g N_VPWR_c_1662_n 0.00981564f $X=1.375 $Y=2.64 $X2=0 $Y2=0
cc_408 N_D_M1017_g N_A_293_464#_c_1830_n 0.012302f $X=1.375 $Y=2.64 $X2=0 $Y2=0
cc_409 N_D_M1040_g N_A_293_464#_c_1818_n 0.0124194f $X=1.455 $Y=0.58 $X2=0 $Y2=0
cc_410 N_D_M1040_g N_A_293_464#_c_1820_n 0.00512834f $X=1.455 $Y=0.58 $X2=0
+ $Y2=0
cc_411 N_D_M1040_g N_A_293_464#_c_1821_n 0.00342727f $X=1.455 $Y=0.58 $X2=0
+ $Y2=0
cc_412 N_D_c_460_n N_A_293_464#_c_1821_n 0.00111607f $X=1.42 $Y=1.955 $X2=0
+ $Y2=0
cc_413 N_D_M1040_g N_VGND_c_2065_n 0.00434272f $X=1.455 $Y=0.58 $X2=0 $Y2=0
cc_414 N_D_M1040_g N_VGND_c_2075_n 0.00821077f $X=1.455 $Y=0.58 $X2=0 $Y2=0
cc_415 N_SCD_c_496_n N_CLK_c_539_n 0.00165831f $X=2.597 $Y=1.372 $X2=-0.19
+ $Y2=-0.245
cc_416 N_SCD_c_496_n N_CLK_c_540_n 0.00841032f $X=2.597 $Y=1.372 $X2=0 $Y2=0
cc_417 N_SCD_c_497_n N_CLK_c_540_n 0.00596561f $X=2.597 $Y=1.918 $X2=0 $Y2=0
cc_418 N_SCD_c_495_n N_A_594_74#_c_1133_n 0.00350312f $X=2.275 $Y=0.865 $X2=0
+ $Y2=0
cc_419 N_SCD_c_496_n N_A_594_74#_c_1133_n 0.00561892f $X=2.597 $Y=1.372 $X2=0
+ $Y2=0
cc_420 N_SCD_c_496_n N_A_594_74#_c_1134_n 0.00681279f $X=2.597 $Y=1.372 $X2=0
+ $Y2=0
cc_421 SCD N_A_594_74#_c_1134_n 0.0493209f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_422 N_SCD_c_497_n N_A_594_74#_c_1148_n 0.00415065f $X=2.597 $Y=1.918 $X2=0
+ $Y2=0
cc_423 SCD N_A_594_74#_c_1148_n 0.0266661f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_424 N_SCD_c_499_n N_VPWR_c_1664_n 0.00545963f $X=2.425 $Y=2.24 $X2=0 $Y2=0
cc_425 N_SCD_c_499_n N_VPWR_c_1679_n 0.00504688f $X=2.425 $Y=2.24 $X2=0 $Y2=0
cc_426 N_SCD_c_499_n N_VPWR_c_1662_n 0.00534614f $X=2.425 $Y=2.24 $X2=0 $Y2=0
cc_427 N_SCD_c_495_n N_A_293_464#_c_1818_n 0.00199036f $X=2.275 $Y=0.865 $X2=0
+ $Y2=0
cc_428 N_SCD_c_496_n N_A_293_464#_c_1819_n 0.017869f $X=2.597 $Y=1.372 $X2=0
+ $Y2=0
cc_429 N_SCD_c_499_n N_A_293_464#_c_1845_n 0.00594919f $X=2.425 $Y=2.24 $X2=0
+ $Y2=0
cc_430 N_SCD_c_499_n N_A_293_464#_c_1821_n 0.0139631f $X=2.425 $Y=2.24 $X2=0
+ $Y2=0
cc_431 N_SCD_c_496_n N_A_293_464#_c_1821_n 0.00695808f $X=2.597 $Y=1.372 $X2=0
+ $Y2=0
cc_432 N_SCD_c_497_n N_A_293_464#_c_1821_n 0.0145162f $X=2.597 $Y=1.918 $X2=0
+ $Y2=0
cc_433 SCD N_A_293_464#_c_1821_n 0.0694511f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_434 N_SCD_c_499_n N_A_293_464#_c_1850_n 0.00668348f $X=2.425 $Y=2.24 $X2=0
+ $Y2=0
cc_435 N_SCD_c_499_n N_A_293_464#_c_1825_n 0.0189446f $X=2.425 $Y=2.24 $X2=0
+ $Y2=0
cc_436 SCD N_A_293_464#_c_1825_n 0.015765f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_437 N_SCD_c_499_n N_A_293_464#_c_1851_n 4.63834e-19 $X=2.425 $Y=2.24 $X2=0
+ $Y2=0
cc_438 N_SCD_c_499_n N_A_293_464#_c_1854_n 0.00176583f $X=2.425 $Y=2.24 $X2=0
+ $Y2=0
cc_439 N_SCD_c_495_n N_VGND_c_2060_n 0.0121542f $X=2.275 $Y=0.865 $X2=0 $Y2=0
cc_440 N_SCD_c_496_n N_VGND_c_2060_n 0.00915488f $X=2.597 $Y=1.372 $X2=0 $Y2=0
cc_441 SCD N_VGND_c_2060_n 0.00453686f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_442 N_SCD_c_495_n N_VGND_c_2065_n 0.00383152f $X=2.275 $Y=0.865 $X2=0 $Y2=0
cc_443 N_SCD_c_495_n N_VGND_c_2075_n 0.0075725f $X=2.275 $Y=0.865 $X2=0 $Y2=0
cc_444 N_CLK_c_539_n N_A_594_74#_c_1124_n 0.0188174f $X=3.33 $Y=1.22 $X2=0 $Y2=0
cc_445 CLK N_A_594_74#_c_1124_n 0.0024284f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_446 N_CLK_c_540_n N_A_594_74#_M1030_g 0.052444f $X=3.515 $Y=1.76 $X2=0 $Y2=0
cc_447 N_CLK_c_539_n N_A_594_74#_c_1133_n 6.68688e-19 $X=3.33 $Y=1.22 $X2=0
+ $Y2=0
cc_448 N_CLK_c_539_n N_A_594_74#_c_1134_n 0.00522155f $X=3.33 $Y=1.22 $X2=0
+ $Y2=0
cc_449 N_CLK_c_540_n N_A_594_74#_c_1134_n 0.00824249f $X=3.515 $Y=1.76 $X2=0
+ $Y2=0
cc_450 CLK N_A_594_74#_c_1134_n 0.028374f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_451 N_CLK_c_540_n N_A_594_74#_c_1149_n 0.00953417f $X=3.515 $Y=1.76 $X2=0
+ $Y2=0
cc_452 N_CLK_c_540_n N_A_594_74#_c_1135_n 0.00197122f $X=3.515 $Y=1.76 $X2=0
+ $Y2=0
cc_453 CLK N_A_594_74#_c_1135_n 0.0267715f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_454 N_CLK_c_540_n N_A_594_74#_c_1136_n 0.0185833f $X=3.515 $Y=1.76 $X2=0
+ $Y2=0
cc_455 CLK N_A_594_74#_c_1136_n 0.00149275f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_456 N_CLK_c_540_n N_A_594_74#_c_1151_n 0.00523766f $X=3.515 $Y=1.76 $X2=0
+ $Y2=0
cc_457 CLK N_A_594_74#_c_1151_n 0.0241043f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_458 N_CLK_c_540_n N_A_594_74#_c_1152_n 0.00585841f $X=3.515 $Y=1.76 $X2=0
+ $Y2=0
cc_459 N_CLK_c_540_n N_VPWR_c_1664_n 0.0100305f $X=3.515 $Y=1.76 $X2=0 $Y2=0
cc_460 N_CLK_c_540_n N_VPWR_c_1665_n 0.00460063f $X=3.515 $Y=1.76 $X2=0 $Y2=0
cc_461 N_CLK_c_540_n N_VPWR_c_1666_n 0.0213431f $X=3.515 $Y=1.76 $X2=0 $Y2=0
cc_462 N_CLK_c_540_n N_VPWR_c_1662_n 0.00465993f $X=3.515 $Y=1.76 $X2=0 $Y2=0
cc_463 N_CLK_c_540_n N_A_293_464#_c_1825_n 0.01471f $X=3.515 $Y=1.76 $X2=0 $Y2=0
cc_464 N_CLK_c_539_n N_VGND_c_2060_n 0.00308778f $X=3.33 $Y=1.22 $X2=0 $Y2=0
cc_465 N_CLK_c_539_n N_VGND_c_2061_n 0.0139212f $X=3.33 $Y=1.22 $X2=0 $Y2=0
cc_466 N_CLK_c_540_n N_VGND_c_2061_n 8.24718e-19 $X=3.515 $Y=1.76 $X2=0 $Y2=0
cc_467 CLK N_VGND_c_2061_n 0.0254134f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_468 N_CLK_c_539_n N_VGND_c_2070_n 0.00383152f $X=3.33 $Y=1.22 $X2=0 $Y2=0
cc_469 N_CLK_c_539_n N_VGND_c_2075_n 0.00762539f $X=3.33 $Y=1.22 $X2=0 $Y2=0
cc_470 N_A_781_74#_M1007_g N_A_1163_48#_c_779_n 0.0511043f $X=5.5 $Y=0.58 $X2=0
+ $Y2=0
cc_471 N_A_781_74#_c_589_n N_A_1163_48#_c_780_n 0.00125914f $X=5.725 $Y=2.255
+ $X2=0 $Y2=0
cc_472 N_A_781_74#_c_591_n N_A_1163_48#_c_780_n 0.00428061f $X=6.595 $Y=2.17
+ $X2=0 $Y2=0
cc_473 N_A_781_74#_c_599_n N_A_1163_48#_c_780_n 0.0197055f $X=5.645 $Y=1.855
+ $X2=0 $Y2=0
cc_474 N_A_781_74#_c_589_n N_A_1163_48#_M1021_g 0.0021815f $X=5.725 $Y=2.255
+ $X2=0 $Y2=0
cc_475 N_A_781_74#_c_590_n N_A_1163_48#_M1021_g 0.00697967f $X=5.725 $Y=2.905
+ $X2=0 $Y2=0
cc_476 N_A_781_74#_c_591_n N_A_1163_48#_M1021_g 0.0190394f $X=6.595 $Y=2.17
+ $X2=0 $Y2=0
cc_477 N_A_781_74#_c_592_n N_A_1163_48#_M1021_g 0.00358158f $X=6.68 $Y=2.905
+ $X2=0 $Y2=0
cc_478 N_A_781_74#_M1007_g N_A_1163_48#_c_781_n 0.0114125f $X=5.5 $Y=0.58 $X2=0
+ $Y2=0
cc_479 N_A_781_74#_M1007_g N_A_1163_48#_c_782_n 0.00153185f $X=5.5 $Y=0.58 $X2=0
+ $Y2=0
cc_480 N_A_781_74#_c_589_n N_A_1163_48#_c_786_n 0.0133533f $X=5.725 $Y=2.255
+ $X2=0 $Y2=0
cc_481 N_A_781_74#_c_591_n N_A_1163_48#_c_786_n 0.0541693f $X=6.595 $Y=2.17
+ $X2=0 $Y2=0
cc_482 N_A_781_74#_c_599_n N_A_1163_48#_c_786_n 2.73581e-19 $X=5.645 $Y=1.855
+ $X2=0 $Y2=0
cc_483 N_A_781_74#_c_591_n N_A_1163_48#_c_787_n 0.0135839f $X=6.595 $Y=2.17
+ $X2=0 $Y2=0
cc_484 N_A_781_74#_c_592_n N_A_1163_48#_c_787_n 0.0184532f $X=6.68 $Y=2.905
+ $X2=0 $Y2=0
cc_485 N_A_781_74#_c_593_n N_A_1163_48#_c_787_n 0.0127728f $X=7.275 $Y=2.99
+ $X2=0 $Y2=0
cc_486 N_A_781_74#_c_595_n N_A_1163_48#_c_787_n 0.0298576f $X=7.36 $Y=2.905
+ $X2=0 $Y2=0
cc_487 N_A_781_74#_c_597_n N_A_1163_48#_c_787_n 0.0143554f $X=7.445 $Y=2.035
+ $X2=0 $Y2=0
cc_488 N_A_781_74#_c_591_n N_A_995_74#_M1038_g 0.00619526f $X=6.595 $Y=2.17
+ $X2=0 $Y2=0
cc_489 N_A_781_74#_c_592_n N_A_995_74#_M1038_g 0.0162004f $X=6.68 $Y=2.905 $X2=0
+ $Y2=0
cc_490 N_A_781_74#_c_593_n N_A_995_74#_M1038_g 0.00295426f $X=7.275 $Y=2.99
+ $X2=0 $Y2=0
cc_491 N_A_781_74#_c_595_n N_A_995_74#_M1038_g 0.00120184f $X=7.36 $Y=2.905
+ $X2=0 $Y2=0
cc_492 N_A_781_74#_c_595_n N_A_995_74#_M1041_g 0.0011633f $X=7.36 $Y=2.905 $X2=0
+ $Y2=0
cc_493 N_A_781_74#_c_596_n N_A_995_74#_M1041_g 0.0204573f $X=8.66 $Y=2.035 $X2=0
+ $Y2=0
cc_494 N_A_781_74#_c_598_n N_A_995_74#_M1041_g 0.00330602f $X=8.745 $Y=1.95
+ $X2=0 $Y2=0
cc_495 N_A_781_74#_c_580_n N_A_995_74#_M1041_g 0.00181619f $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_496 N_A_781_74#_c_581_n N_A_995_74#_M1041_g 0.00661894f $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_497 N_A_781_74#_M1025_g N_A_995_74#_c_853_n 0.0322153f $X=8.735 $Y=0.69 $X2=0
+ $Y2=0
cc_498 N_A_781_74#_M1007_g N_A_995_74#_c_854_n 0.0256791f $X=5.5 $Y=0.58 $X2=0
+ $Y2=0
cc_499 N_A_781_74#_c_575_n N_A_995_74#_c_854_n 0.00381334f $X=4.86 $Y=0.34 $X2=0
+ $Y2=0
cc_500 N_A_781_74#_c_579_n N_A_995_74#_c_854_n 0.0574008f $X=4.895 $Y=1.37 $X2=0
+ $Y2=0
cc_501 N_A_781_74#_M1022_g N_A_995_74#_c_855_n 0.00646319f $X=4.985 $Y=2.525
+ $X2=0 $Y2=0
cc_502 N_A_781_74#_M1007_g N_A_995_74#_c_855_n 0.00415339f $X=5.5 $Y=0.58 $X2=0
+ $Y2=0
cc_503 N_A_781_74#_c_587_n N_A_995_74#_c_855_n 0.0378893f $X=4.925 $Y=1.535
+ $X2=0 $Y2=0
cc_504 N_A_781_74#_c_578_n N_A_995_74#_c_855_n 0.00319045f $X=4.925 $Y=1.535
+ $X2=0 $Y2=0
cc_505 N_A_781_74#_c_589_n N_A_995_74#_c_855_n 0.03794f $X=5.725 $Y=2.255 $X2=0
+ $Y2=0
cc_506 N_A_781_74#_c_590_n N_A_995_74#_c_855_n 0.00571505f $X=5.725 $Y=2.905
+ $X2=0 $Y2=0
cc_507 N_A_781_74#_c_599_n N_A_995_74#_c_855_n 0.00159541f $X=5.645 $Y=1.855
+ $X2=0 $Y2=0
cc_508 N_A_781_74#_c_601_n N_A_995_74#_c_855_n 0.0136656f $X=5.425 $Y=1.855
+ $X2=0 $Y2=0
cc_509 N_A_781_74#_M1007_g N_A_995_74#_c_856_n 0.014507f $X=5.5 $Y=0.58 $X2=0
+ $Y2=0
cc_510 N_A_781_74#_c_589_n N_A_995_74#_c_856_n 0.0210075f $X=5.725 $Y=2.255
+ $X2=0 $Y2=0
cc_511 N_A_781_74#_c_591_n N_A_995_74#_c_856_n 0.00772262f $X=6.595 $Y=2.17
+ $X2=0 $Y2=0
cc_512 N_A_781_74#_c_599_n N_A_995_74#_c_856_n 0.00165663f $X=5.645 $Y=1.855
+ $X2=0 $Y2=0
cc_513 N_A_781_74#_M1025_g N_A_995_74#_c_858_n 0.00114708f $X=8.735 $Y=0.69
+ $X2=0 $Y2=0
cc_514 N_A_781_74#_c_596_n N_A_995_74#_c_858_n 0.00418131f $X=8.66 $Y=2.035
+ $X2=0 $Y2=0
cc_515 N_A_781_74#_c_580_n N_A_995_74#_c_858_n 0.00313951f $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_516 N_A_781_74#_c_585_n N_A_995_74#_c_865_n 0.0242351f $X=5.64 $Y=2.99 $X2=0
+ $Y2=0
cc_517 N_A_781_74#_c_590_n N_A_995_74#_c_865_n 0.0120463f $X=5.725 $Y=2.905
+ $X2=0 $Y2=0
cc_518 N_A_781_74#_c_599_n N_A_995_74#_c_865_n 8.90055e-19 $X=5.645 $Y=1.855
+ $X2=0 $Y2=0
cc_519 N_A_781_74#_c_601_n N_A_995_74#_c_865_n 0.00385746f $X=5.425 $Y=1.855
+ $X2=0 $Y2=0
cc_520 N_A_781_74#_M1007_g N_A_995_74#_c_859_n 0.00354176f $X=5.5 $Y=0.58 $X2=0
+ $Y2=0
cc_521 N_A_781_74#_c_578_n N_A_995_74#_c_859_n 0.00130826f $X=4.925 $Y=1.535
+ $X2=0 $Y2=0
cc_522 N_A_781_74#_c_579_n N_A_995_74#_c_859_n 0.0140925f $X=4.895 $Y=1.37 $X2=0
+ $Y2=0
cc_523 N_A_781_74#_c_596_n N_A_995_74#_c_861_n 0.00785247f $X=8.66 $Y=2.035
+ $X2=0 $Y2=0
cc_524 N_A_781_74#_c_580_n N_A_995_74#_c_861_n 4.66986e-19 $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_525 N_A_781_74#_c_581_n N_A_995_74#_c_861_n 0.0322153f $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_526 N_A_781_74#_c_592_n N_SET_B_M1035_g 2.34711e-19 $X=6.68 $Y=2.905 $X2=0
+ $Y2=0
cc_527 N_A_781_74#_c_595_n N_SET_B_M1035_g 0.0219318f $X=7.36 $Y=2.905 $X2=0
+ $Y2=0
cc_528 N_A_781_74#_c_596_n N_SET_B_M1035_g 0.00451686f $X=8.66 $Y=2.035 $X2=0
+ $Y2=0
cc_529 N_A_781_74#_c_597_n N_SET_B_M1035_g 0.00552929f $X=7.445 $Y=2.035 $X2=0
+ $Y2=0
cc_530 N_A_781_74#_c_596_n N_SET_B_c_986_n 0.0393802f $X=8.66 $Y=2.035 $X2=0
+ $Y2=0
cc_531 N_A_781_74#_c_598_n N_SET_B_c_986_n 0.00672398f $X=8.745 $Y=1.95 $X2=0
+ $Y2=0
cc_532 N_A_781_74#_c_580_n N_SET_B_c_986_n 0.0177158f $X=8.825 $Y=1.515 $X2=0
+ $Y2=0
cc_533 N_A_781_74#_c_581_n N_SET_B_c_986_n 0.00479238f $X=8.825 $Y=1.515 $X2=0
+ $Y2=0
cc_534 N_A_781_74#_c_596_n N_SET_B_c_987_n 0.00105565f $X=8.66 $Y=2.035 $X2=0
+ $Y2=0
cc_535 N_A_781_74#_c_597_n N_SET_B_c_987_n 0.00120115f $X=7.445 $Y=2.035 $X2=0
+ $Y2=0
cc_536 N_A_781_74#_c_596_n N_SET_B_c_989_n 6.49836e-19 $X=8.66 $Y=2.035 $X2=0
+ $Y2=0
cc_537 N_A_781_74#_c_596_n N_SET_B_c_990_n 0.0120873f $X=8.66 $Y=2.035 $X2=0
+ $Y2=0
cc_538 N_A_781_74#_c_597_n N_SET_B_c_990_n 0.0100795f $X=7.445 $Y=2.035 $X2=0
+ $Y2=0
cc_539 N_A_781_74#_c_574_n N_A_594_74#_c_1124_n 0.00651805f $X=4.045 $Y=0.505
+ $X2=0 $Y2=0
cc_540 N_A_781_74#_c_576_n N_A_594_74#_c_1124_n 0.00462516f $X=4.21 $Y=0.34
+ $X2=0 $Y2=0
cc_541 N_A_781_74#_c_586_n N_A_594_74#_M1030_g 0.00112829f $X=4.355 $Y=2.99
+ $X2=0 $Y2=0
cc_542 N_A_781_74#_M1022_g N_A_594_74#_c_1127_n 0.0201046f $X=4.985 $Y=2.525
+ $X2=0 $Y2=0
cc_543 N_A_781_74#_c_584_n N_A_594_74#_c_1127_n 0.00626763f $X=4.19 $Y=2.765
+ $X2=0 $Y2=0
cc_544 N_A_781_74#_c_585_n N_A_594_74#_c_1127_n 0.0113283f $X=5.64 $Y=2.99 $X2=0
+ $Y2=0
cc_545 N_A_781_74#_c_587_n N_A_594_74#_c_1127_n 3.88824e-19 $X=4.925 $Y=1.535
+ $X2=0 $Y2=0
cc_546 N_A_781_74#_c_575_n N_A_594_74#_c_1128_n 0.00253049f $X=4.86 $Y=0.34
+ $X2=0 $Y2=0
cc_547 N_A_781_74#_c_577_n N_A_594_74#_c_1128_n 6.71829e-19 $X=4.895 $Y=1.505
+ $X2=0 $Y2=0
cc_548 N_A_781_74#_c_578_n N_A_594_74#_c_1128_n 0.0116591f $X=4.925 $Y=1.535
+ $X2=0 $Y2=0
cc_549 N_A_781_74#_c_579_n N_A_594_74#_c_1128_n 0.00664279f $X=4.895 $Y=1.37
+ $X2=0 $Y2=0
cc_550 N_A_781_74#_M1022_g N_A_594_74#_c_1140_n 0.0105864f $X=4.985 $Y=2.525
+ $X2=0 $Y2=0
cc_551 N_A_781_74#_c_585_n N_A_594_74#_c_1140_n 0.0150766f $X=5.64 $Y=2.99 $X2=0
+ $Y2=0
cc_552 N_A_781_74#_M1007_g N_A_594_74#_M1037_g 0.0160063f $X=5.5 $Y=0.58 $X2=0
+ $Y2=0
cc_553 N_A_781_74#_c_574_n N_A_594_74#_M1037_g 0.00301996f $X=4.045 $Y=0.505
+ $X2=0 $Y2=0
cc_554 N_A_781_74#_c_575_n N_A_594_74#_M1037_g 0.010044f $X=4.86 $Y=0.34 $X2=0
+ $Y2=0
cc_555 N_A_781_74#_c_579_n N_A_594_74#_M1037_g 0.0157578f $X=4.895 $Y=1.37 $X2=0
+ $Y2=0
cc_556 N_A_781_74#_M1022_g N_A_594_74#_M1020_g 0.0131318f $X=4.985 $Y=2.525
+ $X2=0 $Y2=0
cc_557 N_A_781_74#_c_585_n N_A_594_74#_M1020_g 0.0169016f $X=5.64 $Y=2.99 $X2=0
+ $Y2=0
cc_558 N_A_781_74#_c_589_n N_A_594_74#_M1020_g 7.58855e-19 $X=5.725 $Y=2.255
+ $X2=0 $Y2=0
cc_559 N_A_781_74#_c_590_n N_A_594_74#_M1020_g 0.0166185f $X=5.725 $Y=2.905
+ $X2=0 $Y2=0
cc_560 N_A_781_74#_c_599_n N_A_594_74#_M1020_g 0.0108493f $X=5.645 $Y=1.855
+ $X2=0 $Y2=0
cc_561 N_A_781_74#_c_585_n N_A_594_74#_c_1143_n 0.00206861f $X=5.64 $Y=2.99
+ $X2=0 $Y2=0
cc_562 N_A_781_74#_c_593_n N_A_594_74#_c_1143_n 0.0116627f $X=7.275 $Y=2.99
+ $X2=0 $Y2=0
cc_563 N_A_781_74#_c_594_n N_A_594_74#_c_1143_n 0.00320029f $X=6.765 $Y=2.99
+ $X2=0 $Y2=0
cc_564 N_A_781_74#_c_602_n N_A_594_74#_c_1143_n 0.00189476f $X=8.825 $Y=1.795
+ $X2=0 $Y2=0
cc_565 N_A_781_74#_M1025_g N_A_594_74#_M1003_g 0.0205499f $X=8.735 $Y=0.69 $X2=0
+ $Y2=0
cc_566 N_A_781_74#_c_580_n N_A_594_74#_M1003_g 4.68509e-19 $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_567 N_A_781_74#_c_581_n N_A_594_74#_M1003_g 0.0242476f $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_568 N_A_781_74#_c_602_n N_A_594_74#_M1008_g 0.0148225f $X=8.825 $Y=1.795
+ $X2=0 $Y2=0
cc_569 N_A_781_74#_c_574_n N_A_594_74#_c_1132_n 3.03407e-19 $X=4.045 $Y=0.505
+ $X2=0 $Y2=0
cc_570 N_A_781_74#_c_575_n N_A_594_74#_c_1132_n 5.72887e-19 $X=4.86 $Y=0.34
+ $X2=0 $Y2=0
cc_571 N_A_781_74#_c_577_n N_A_594_74#_c_1132_n 3.88824e-19 $X=4.895 $Y=1.505
+ $X2=0 $Y2=0
cc_572 N_A_781_74#_c_578_n N_A_594_74#_c_1132_n 0.0423314f $X=4.925 $Y=1.535
+ $X2=0 $Y2=0
cc_573 N_A_781_74#_c_579_n N_A_594_74#_c_1132_n 8.69379e-19 $X=4.895 $Y=1.37
+ $X2=0 $Y2=0
cc_574 N_A_781_74#_c_585_n N_A_594_74#_c_1146_n 3.42637e-19 $X=5.64 $Y=2.99
+ $X2=0 $Y2=0
cc_575 N_A_781_74#_M1030_d N_A_594_74#_c_1149_n 0.00269298f $X=4.055 $Y=1.84
+ $X2=0 $Y2=0
cc_576 N_A_781_74#_c_574_n N_A_594_74#_c_1135_n 0.0216703f $X=4.045 $Y=0.505
+ $X2=0 $Y2=0
cc_577 N_A_781_74#_c_574_n N_A_594_74#_c_1136_n 0.00163297f $X=4.045 $Y=0.505
+ $X2=0 $Y2=0
cc_578 N_A_781_74#_M1025_g N_A_1762_74#_c_1441_n 0.0185265f $X=8.735 $Y=0.69
+ $X2=0 $Y2=0
cc_579 N_A_781_74#_c_580_n N_A_1762_74#_c_1441_n 0.0100316f $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_580 N_A_781_74#_c_581_n N_A_1762_74#_c_1441_n 0.00130485f $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_581 N_A_781_74#_c_598_n N_A_1762_74#_c_1456_n 0.00345252f $X=8.745 $Y=1.95
+ $X2=0 $Y2=0
cc_582 N_A_781_74#_c_602_n N_A_1762_74#_c_1456_n 0.00187605f $X=8.825 $Y=1.795
+ $X2=0 $Y2=0
cc_583 N_A_781_74#_M1025_g N_A_1762_74#_c_1442_n 0.0041777f $X=8.735 $Y=0.69
+ $X2=0 $Y2=0
cc_584 N_A_781_74#_c_598_n N_A_1762_74#_c_1442_n 0.00405579f $X=8.745 $Y=1.95
+ $X2=0 $Y2=0
cc_585 N_A_781_74#_c_580_n N_A_1762_74#_c_1442_n 0.0195875f $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_586 N_A_781_74#_c_581_n N_A_1762_74#_c_1442_n 0.00250898f $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_587 N_A_781_74#_c_592_n N_VPWR_M1021_d 0.00437233f $X=6.68 $Y=2.905 $X2=0
+ $Y2=0
cc_588 N_A_781_74#_c_596_n N_VPWR_M1035_d 0.00533961f $X=8.66 $Y=2.035 $X2=0
+ $Y2=0
cc_589 N_A_781_74#_c_586_n N_VPWR_c_1666_n 0.0103602f $X=4.355 $Y=2.99 $X2=0
+ $Y2=0
cc_590 N_A_781_74#_c_585_n N_VPWR_c_1667_n 0.00867486f $X=5.64 $Y=2.99 $X2=0
+ $Y2=0
cc_591 N_A_781_74#_c_590_n N_VPWR_c_1667_n 0.0195575f $X=5.725 $Y=2.905 $X2=0
+ $Y2=0
cc_592 N_A_781_74#_c_591_n N_VPWR_c_1667_n 0.0177503f $X=6.595 $Y=2.17 $X2=0
+ $Y2=0
cc_593 N_A_781_74#_c_592_n N_VPWR_c_1667_n 0.0363339f $X=6.68 $Y=2.905 $X2=0
+ $Y2=0
cc_594 N_A_781_74#_c_594_n N_VPWR_c_1667_n 0.0147459f $X=6.765 $Y=2.99 $X2=0
+ $Y2=0
cc_595 N_A_781_74#_c_593_n N_VPWR_c_1668_n 0.0143583f $X=7.275 $Y=2.99 $X2=0
+ $Y2=0
cc_596 N_A_781_74#_c_595_n N_VPWR_c_1668_n 0.0431623f $X=7.36 $Y=2.905 $X2=0
+ $Y2=0
cc_597 N_A_781_74#_c_596_n N_VPWR_c_1668_n 0.0124646f $X=8.66 $Y=2.035 $X2=0
+ $Y2=0
cc_598 N_A_781_74#_c_585_n N_VPWR_c_1672_n 0.0934179f $X=5.64 $Y=2.99 $X2=0
+ $Y2=0
cc_599 N_A_781_74#_c_586_n N_VPWR_c_1672_n 0.0175791f $X=4.355 $Y=2.99 $X2=0
+ $Y2=0
cc_600 N_A_781_74#_c_593_n N_VPWR_c_1674_n 0.0443733f $X=7.275 $Y=2.99 $X2=0
+ $Y2=0
cc_601 N_A_781_74#_c_594_n N_VPWR_c_1674_n 0.0115893f $X=6.765 $Y=2.99 $X2=0
+ $Y2=0
cc_602 N_A_781_74#_c_585_n N_VPWR_c_1662_n 0.0489384f $X=5.64 $Y=2.99 $X2=0
+ $Y2=0
cc_603 N_A_781_74#_c_586_n N_VPWR_c_1662_n 0.00965514f $X=4.355 $Y=2.99 $X2=0
+ $Y2=0
cc_604 N_A_781_74#_c_593_n N_VPWR_c_1662_n 0.0229659f $X=7.275 $Y=2.99 $X2=0
+ $Y2=0
cc_605 N_A_781_74#_c_594_n N_VPWR_c_1662_n 0.00583135f $X=6.765 $Y=2.99 $X2=0
+ $Y2=0
cc_606 N_A_781_74#_c_575_n N_A_293_464#_M1037_s 0.00402708f $X=4.86 $Y=0.34
+ $X2=0 $Y2=0
cc_607 N_A_781_74#_M1030_d N_A_293_464#_c_1826_n 0.00565638f $X=4.055 $Y=1.84
+ $X2=0 $Y2=0
cc_608 N_A_781_74#_c_584_n N_A_293_464#_c_1826_n 0.0193673f $X=4.19 $Y=2.765
+ $X2=0 $Y2=0
cc_609 N_A_781_74#_c_585_n N_A_293_464#_c_1826_n 0.00206012f $X=5.64 $Y=2.99
+ $X2=0 $Y2=0
cc_610 N_A_781_74#_M1022_g N_A_293_464#_c_1822_n 0.00142806f $X=4.985 $Y=2.525
+ $X2=0 $Y2=0
cc_611 N_A_781_74#_c_574_n N_A_293_464#_c_1822_n 0.00569556f $X=4.045 $Y=0.505
+ $X2=0 $Y2=0
cc_612 N_A_781_74#_c_577_n N_A_293_464#_c_1822_n 0.0495574f $X=4.895 $Y=1.505
+ $X2=0 $Y2=0
cc_613 N_A_781_74#_c_578_n N_A_293_464#_c_1822_n 0.00362303f $X=4.925 $Y=1.535
+ $X2=0 $Y2=0
cc_614 N_A_781_74#_c_579_n N_A_293_464#_c_1822_n 0.0228629f $X=4.895 $Y=1.37
+ $X2=0 $Y2=0
cc_615 N_A_781_74#_M1022_g N_A_293_464#_c_1828_n 0.0047804f $X=4.985 $Y=2.525
+ $X2=0 $Y2=0
cc_616 N_A_781_74#_c_584_n N_A_293_464#_c_1828_n 0.0120315f $X=4.19 $Y=2.765
+ $X2=0 $Y2=0
cc_617 N_A_781_74#_c_585_n N_A_293_464#_c_1828_n 0.0230985f $X=5.64 $Y=2.99
+ $X2=0 $Y2=0
cc_618 N_A_781_74#_c_574_n N_A_293_464#_c_1823_n 0.0232909f $X=4.045 $Y=0.505
+ $X2=0 $Y2=0
cc_619 N_A_781_74#_c_575_n N_A_293_464#_c_1823_n 0.0194638f $X=4.86 $Y=0.34
+ $X2=0 $Y2=0
cc_620 N_A_781_74#_c_579_n N_A_293_464#_c_1823_n 0.0240322f $X=4.895 $Y=1.37
+ $X2=0 $Y2=0
cc_621 N_A_781_74#_M1022_g N_A_293_464#_c_1829_n 0.00432855f $X=4.985 $Y=2.525
+ $X2=0 $Y2=0
cc_622 N_A_781_74#_c_585_n N_A_293_464#_c_1829_n 0.00542945f $X=5.64 $Y=2.99
+ $X2=0 $Y2=0
cc_623 N_A_781_74#_c_587_n N_A_293_464#_c_1829_n 0.01419f $X=4.925 $Y=1.535
+ $X2=0 $Y2=0
cc_624 N_A_781_74#_c_578_n N_A_293_464#_c_1829_n 0.00102084f $X=4.925 $Y=1.535
+ $X2=0 $Y2=0
cc_625 N_A_781_74#_c_590_n A_1136_478# 0.00580115f $X=5.725 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_626 N_A_781_74#_c_596_n N_A_1603_347#_M1041_d 0.00509997f $X=8.66 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_627 N_A_781_74#_c_596_n N_A_1603_347#_c_1946_n 0.0281246f $X=8.66 $Y=2.035
+ $X2=0 $Y2=0
cc_628 N_A_781_74#_c_580_n N_A_1603_347#_c_1946_n 0.00160222f $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_629 N_A_781_74#_c_581_n N_A_1603_347#_c_1946_n 5.17038e-19 $X=8.825 $Y=1.515
+ $X2=0 $Y2=0
cc_630 N_A_781_74#_c_602_n N_A_1603_347#_c_1946_n 0.0106929f $X=8.825 $Y=1.795
+ $X2=0 $Y2=0
cc_631 N_A_781_74#_c_596_n N_A_1603_347#_c_1947_n 0.0206512f $X=8.66 $Y=2.035
+ $X2=0 $Y2=0
cc_632 N_A_781_74#_c_602_n N_A_1603_347#_c_1947_n 0.00180187f $X=8.825 $Y=1.795
+ $X2=0 $Y2=0
cc_633 N_A_781_74#_c_596_n N_A_1712_374#_M1033_s 0.00427293f $X=8.66 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_634 N_A_781_74#_c_598_n N_A_1712_374#_M1033_s 0.00137281f $X=8.745 $Y=1.95
+ $X2=-0.19 $Y2=-0.245
cc_635 N_A_781_74#_c_602_n N_A_1712_374#_c_1980_n 4.33337e-19 $X=8.825 $Y=1.795
+ $X2=0 $Y2=0
cc_636 N_A_781_74#_c_576_n N_VGND_c_2061_n 0.011924f $X=4.21 $Y=0.34 $X2=0 $Y2=0
cc_637 N_A_781_74#_M1007_g N_VGND_c_2067_n 0.00434272f $X=5.5 $Y=0.58 $X2=0
+ $Y2=0
cc_638 N_A_781_74#_c_575_n N_VGND_c_2067_n 0.0534972f $X=4.86 $Y=0.34 $X2=0
+ $Y2=0
cc_639 N_A_781_74#_c_576_n N_VGND_c_2067_n 0.0235688f $X=4.21 $Y=0.34 $X2=0
+ $Y2=0
cc_640 N_A_781_74#_M1025_g N_VGND_c_2071_n 0.00434272f $X=8.735 $Y=0.69 $X2=0
+ $Y2=0
cc_641 N_A_781_74#_M1007_g N_VGND_c_2075_n 0.00822443f $X=5.5 $Y=0.58 $X2=0
+ $Y2=0
cc_642 N_A_781_74#_M1025_g N_VGND_c_2075_n 0.00822232f $X=8.735 $Y=0.69 $X2=0
+ $Y2=0
cc_643 N_A_781_74#_c_575_n N_VGND_c_2075_n 0.0303548f $X=4.86 $Y=0.34 $X2=0
+ $Y2=0
cc_644 N_A_781_74#_c_576_n N_VGND_c_2075_n 0.0127152f $X=4.21 $Y=0.34 $X2=0
+ $Y2=0
cc_645 N_A_781_74#_M1025_g N_VGND_c_2079_n 0.00164121f $X=8.735 $Y=0.69 $X2=0
+ $Y2=0
cc_646 N_A_1163_48#_c_781_n N_A_995_74#_c_849_n 0.00856703f $X=6.125 $Y=1.635
+ $X2=0 $Y2=0
cc_647 N_A_1163_48#_c_782_n N_A_995_74#_c_849_n 9.45781e-19 $X=6.263 $Y=0.957
+ $X2=0 $Y2=0
cc_648 N_A_1163_48#_c_786_n N_A_995_74#_c_849_n 0.00129303f $X=6.935 $Y=1.802
+ $X2=0 $Y2=0
cc_649 N_A_1163_48#_c_783_n N_A_995_74#_c_849_n 0.00225195f $X=6.32 $Y=1.065
+ $X2=0 $Y2=0
cc_650 N_A_1163_48#_c_780_n N_A_995_74#_M1038_g 0.0132022f $X=6.11 $Y=1.965
+ $X2=0 $Y2=0
cc_651 N_A_1163_48#_M1021_g N_A_995_74#_M1038_g 0.015118f $X=6.11 $Y=2.525 $X2=0
+ $Y2=0
cc_652 N_A_1163_48#_c_786_n N_A_995_74#_M1038_g 0.0180333f $X=6.935 $Y=1.802
+ $X2=0 $Y2=0
cc_653 N_A_1163_48#_c_787_n N_A_995_74#_M1038_g 0.00662286f $X=7.02 $Y=2.515
+ $X2=0 $Y2=0
cc_654 N_A_1163_48#_c_782_n N_A_995_74#_M1001_g 0.0162848f $X=6.263 $Y=0.957
+ $X2=0 $Y2=0
cc_655 N_A_1163_48#_c_783_n N_A_995_74#_M1001_g 0.00719364f $X=6.32 $Y=1.065
+ $X2=0 $Y2=0
cc_656 N_A_1163_48#_c_779_n N_A_995_74#_c_854_n 0.00195661f $X=5.89 $Y=0.9 $X2=0
+ $Y2=0
cc_657 N_A_1163_48#_c_781_n N_A_995_74#_c_854_n 5.28691e-19 $X=6.125 $Y=1.635
+ $X2=0 $Y2=0
cc_658 N_A_1163_48#_c_782_n N_A_995_74#_c_854_n 0.0186822f $X=6.263 $Y=0.957
+ $X2=0 $Y2=0
cc_659 N_A_1163_48#_c_783_n N_A_995_74#_c_854_n 2.95653e-19 $X=6.32 $Y=1.065
+ $X2=0 $Y2=0
cc_660 N_A_1163_48#_M1021_g N_A_995_74#_c_855_n 6.6776e-19 $X=6.11 $Y=2.525
+ $X2=0 $Y2=0
cc_661 N_A_1163_48#_c_780_n N_A_995_74#_c_856_n 0.00190856f $X=6.11 $Y=1.965
+ $X2=0 $Y2=0
cc_662 N_A_1163_48#_c_781_n N_A_995_74#_c_856_n 0.0123773f $X=6.125 $Y=1.635
+ $X2=0 $Y2=0
cc_663 N_A_1163_48#_c_782_n N_A_995_74#_c_856_n 0.0607821f $X=6.263 $Y=0.957
+ $X2=0 $Y2=0
cc_664 N_A_1163_48#_c_786_n N_A_995_74#_c_856_n 0.0499605f $X=6.935 $Y=1.802
+ $X2=0 $Y2=0
cc_665 N_A_1163_48#_c_783_n N_A_995_74#_c_856_n 0.00984239f $X=6.32 $Y=1.065
+ $X2=0 $Y2=0
cc_666 N_A_1163_48#_c_781_n N_A_995_74#_c_860_n 6.28152e-19 $X=6.125 $Y=1.635
+ $X2=0 $Y2=0
cc_667 N_A_1163_48#_c_782_n N_A_995_74#_c_860_n 0.0172613f $X=6.263 $Y=0.957
+ $X2=0 $Y2=0
cc_668 N_A_1163_48#_c_786_n N_A_995_74#_c_860_n 0.0307973f $X=6.935 $Y=1.802
+ $X2=0 $Y2=0
cc_669 N_A_1163_48#_c_783_n N_A_995_74#_c_860_n 6.81032e-19 $X=6.32 $Y=1.065
+ $X2=0 $Y2=0
cc_670 N_A_1163_48#_c_782_n N_SET_B_M1014_g 0.00113521f $X=6.263 $Y=0.957 $X2=0
+ $Y2=0
cc_671 N_A_1163_48#_c_786_n N_SET_B_M1035_g 0.00444569f $X=6.935 $Y=1.802 $X2=0
+ $Y2=0
cc_672 N_A_1163_48#_c_787_n N_SET_B_M1035_g 0.00338211f $X=7.02 $Y=2.515 $X2=0
+ $Y2=0
cc_673 N_A_1163_48#_c_786_n N_SET_B_c_987_n 0.00248279f $X=6.935 $Y=1.802 $X2=0
+ $Y2=0
cc_674 N_A_1163_48#_c_786_n N_SET_B_c_990_n 0.00565296f $X=6.935 $Y=1.802 $X2=0
+ $Y2=0
cc_675 N_A_1163_48#_M1021_g N_A_594_74#_M1020_g 0.019239f $X=6.11 $Y=2.525 $X2=0
+ $Y2=0
cc_676 N_A_1163_48#_M1021_g N_A_594_74#_c_1143_n 0.0123939f $X=6.11 $Y=2.525
+ $X2=0 $Y2=0
cc_677 N_A_1163_48#_M1021_g N_VPWR_c_1667_n 0.00903974f $X=6.11 $Y=2.525 $X2=0
+ $Y2=0
cc_678 N_A_1163_48#_M1021_g N_VPWR_c_1662_n 9.76808e-19 $X=6.11 $Y=2.525 $X2=0
+ $Y2=0
cc_679 N_A_1163_48#_c_782_n N_VGND_M1005_d 0.0034935f $X=6.263 $Y=0.957 $X2=0
+ $Y2=0
cc_680 N_A_1163_48#_c_779_n N_VGND_c_2062_n 0.00891566f $X=5.89 $Y=0.9 $X2=0
+ $Y2=0
cc_681 N_A_1163_48#_c_782_n N_VGND_c_2062_n 0.043708f $X=6.263 $Y=0.957 $X2=0
+ $Y2=0
cc_682 N_A_1163_48#_c_783_n N_VGND_c_2062_n 0.00185009f $X=6.32 $Y=1.065 $X2=0
+ $Y2=0
cc_683 N_A_1163_48#_c_779_n N_VGND_c_2067_n 0.00336577f $X=5.89 $Y=0.9 $X2=0
+ $Y2=0
cc_684 N_A_1163_48#_c_782_n N_VGND_c_2067_n 0.00250183f $X=6.263 $Y=0.957 $X2=0
+ $Y2=0
cc_685 N_A_1163_48#_c_779_n N_VGND_c_2075_n 0.00442062f $X=5.89 $Y=0.9 $X2=0
+ $Y2=0
cc_686 N_A_1163_48#_c_782_n N_VGND_c_2075_n 0.0245359f $X=6.263 $Y=0.957 $X2=0
+ $Y2=0
cc_687 N_A_1163_48#_c_782_n N_VGND_c_2078_n 0.0178253f $X=6.263 $Y=0.957 $X2=0
+ $Y2=0
cc_688 N_A_1163_48#_c_782_n N_VGND_c_2079_n 0.00571502f $X=6.263 $Y=0.957 $X2=0
+ $Y2=0
cc_689 N_A_995_74#_M1001_g N_SET_B_M1014_g 0.0332539f $X=6.98 $Y=0.58 $X2=0
+ $Y2=0
cc_690 N_A_995_74#_c_857_n N_SET_B_M1014_g 0.0165792f $X=7.835 $Y=0.99 $X2=0
+ $Y2=0
cc_691 N_A_995_74#_c_858_n N_SET_B_M1014_g 0.00202609f $X=8 $Y=1.285 $X2=0 $Y2=0
cc_692 N_A_995_74#_c_860_n N_SET_B_M1014_g 0.00534819f $X=6.89 $Y=1.355 $X2=0
+ $Y2=0
cc_693 N_A_995_74#_c_861_n N_SET_B_M1014_g 0.0044628f $X=8.345 $Y=1.285 $X2=0
+ $Y2=0
cc_694 N_A_995_74#_M1038_g N_SET_B_M1035_g 0.0146973f $X=6.795 $Y=2.525 $X2=0
+ $Y2=0
cc_695 N_A_995_74#_M1041_g N_SET_B_M1035_g 0.035059f $X=7.925 $Y=2.235 $X2=0
+ $Y2=0
cc_696 N_A_995_74#_M1041_g N_SET_B_c_986_n 0.00689996f $X=7.925 $Y=2.235 $X2=0
+ $Y2=0
cc_697 N_A_995_74#_c_857_n N_SET_B_c_986_n 0.00699145f $X=7.835 $Y=0.99 $X2=0
+ $Y2=0
cc_698 N_A_995_74#_c_858_n N_SET_B_c_986_n 0.00966112f $X=8 $Y=1.285 $X2=0 $Y2=0
cc_699 N_A_995_74#_c_861_n N_SET_B_c_986_n 0.00683728f $X=8.345 $Y=1.285 $X2=0
+ $Y2=0
cc_700 N_A_995_74#_c_849_n N_SET_B_c_987_n 7.48901e-19 $X=6.795 $Y=1.61 $X2=0
+ $Y2=0
cc_701 N_A_995_74#_c_857_n N_SET_B_c_987_n 0.0010997f $X=7.835 $Y=0.99 $X2=0
+ $Y2=0
cc_702 N_A_995_74#_c_849_n N_SET_B_c_989_n 0.0479511f $X=6.795 $Y=1.61 $X2=0
+ $Y2=0
cc_703 N_A_995_74#_c_857_n N_SET_B_c_989_n 0.00125903f $X=7.835 $Y=0.99 $X2=0
+ $Y2=0
cc_704 N_A_995_74#_c_858_n N_SET_B_c_989_n 7.13996e-19 $X=8 $Y=1.285 $X2=0 $Y2=0
cc_705 N_A_995_74#_c_861_n N_SET_B_c_989_n 0.0211492f $X=8.345 $Y=1.285 $X2=0
+ $Y2=0
cc_706 N_A_995_74#_c_849_n N_SET_B_c_990_n 0.00180078f $X=6.795 $Y=1.61 $X2=0
+ $Y2=0
cc_707 N_A_995_74#_M1041_g N_SET_B_c_990_n 0.0038802f $X=7.925 $Y=2.235 $X2=0
+ $Y2=0
cc_708 N_A_995_74#_c_857_n N_SET_B_c_990_n 0.0242739f $X=7.835 $Y=0.99 $X2=0
+ $Y2=0
cc_709 N_A_995_74#_c_858_n N_SET_B_c_990_n 0.0129916f $X=8 $Y=1.285 $X2=0 $Y2=0
cc_710 N_A_995_74#_c_860_n N_SET_B_c_990_n 0.0213842f $X=6.89 $Y=1.355 $X2=0
+ $Y2=0
cc_711 N_A_995_74#_c_861_n N_SET_B_c_990_n 0.00163893f $X=8.345 $Y=1.285 $X2=0
+ $Y2=0
cc_712 N_A_995_74#_c_854_n N_A_594_74#_M1037_g 0.0026059f $X=5.285 $Y=0.58 $X2=0
+ $Y2=0
cc_713 N_A_995_74#_c_855_n N_A_594_74#_M1020_g 9.88425e-19 $X=5.285 $Y=2.37
+ $X2=0 $Y2=0
cc_714 N_A_995_74#_c_865_n N_A_594_74#_M1020_g 0.00237895f $X=5.285 $Y=2.55
+ $X2=0 $Y2=0
cc_715 N_A_995_74#_M1038_g N_A_594_74#_c_1143_n 0.0109545f $X=6.795 $Y=2.525
+ $X2=0 $Y2=0
cc_716 N_A_995_74#_M1041_g N_A_594_74#_c_1143_n 0.0123594f $X=7.925 $Y=2.235
+ $X2=0 $Y2=0
cc_717 N_A_995_74#_c_853_n N_A_1762_74#_c_1441_n 0.0023555f $X=8.345 $Y=1.12
+ $X2=0 $Y2=0
cc_718 N_A_995_74#_c_857_n N_A_1762_74#_c_1441_n 0.00454574f $X=7.835 $Y=0.99
+ $X2=0 $Y2=0
cc_719 N_A_995_74#_M1038_g N_VPWR_c_1667_n 0.00133128f $X=6.795 $Y=2.525 $X2=0
+ $Y2=0
cc_720 N_A_995_74#_M1041_g N_VPWR_c_1668_n 0.00322773f $X=7.925 $Y=2.235 $X2=0
+ $Y2=0
cc_721 N_A_995_74#_M1041_g N_VPWR_c_1662_n 0.00112709f $X=7.925 $Y=2.235 $X2=0
+ $Y2=0
cc_722 N_A_995_74#_c_855_n N_A_293_464#_c_1822_n 0.0051899f $X=5.285 $Y=2.37
+ $X2=0 $Y2=0
cc_723 N_A_995_74#_c_855_n N_A_293_464#_c_1829_n 0.00879291f $X=5.285 $Y=2.37
+ $X2=0 $Y2=0
cc_724 N_A_995_74#_M1041_g N_A_1603_347#_c_1947_n 0.00794322f $X=7.925 $Y=2.235
+ $X2=0 $Y2=0
cc_725 N_A_995_74#_M1041_g N_A_1712_374#_c_1982_n 0.00309824f $X=7.925 $Y=2.235
+ $X2=0 $Y2=0
cc_726 N_A_995_74#_c_857_n N_VGND_M1014_d 0.00962076f $X=7.835 $Y=0.99 $X2=0
+ $Y2=0
cc_727 N_A_995_74#_M1001_g N_VGND_c_2062_n 0.00317476f $X=6.98 $Y=0.58 $X2=0
+ $Y2=0
cc_728 N_A_995_74#_c_854_n N_VGND_c_2062_n 0.00319235f $X=5.285 $Y=0.58 $X2=0
+ $Y2=0
cc_729 N_A_995_74#_c_854_n N_VGND_c_2067_n 0.0109942f $X=5.285 $Y=0.58 $X2=0
+ $Y2=0
cc_730 N_A_995_74#_c_853_n N_VGND_c_2071_n 0.00383152f $X=8.345 $Y=1.12 $X2=0
+ $Y2=0
cc_731 N_A_995_74#_M1001_g N_VGND_c_2075_n 0.0082231f $X=6.98 $Y=0.58 $X2=0
+ $Y2=0
cc_732 N_A_995_74#_c_853_n N_VGND_c_2075_n 0.00752635f $X=8.345 $Y=1.12 $X2=0
+ $Y2=0
cc_733 N_A_995_74#_c_854_n N_VGND_c_2075_n 0.00904371f $X=5.285 $Y=0.58 $X2=0
+ $Y2=0
cc_734 N_A_995_74#_M1001_g N_VGND_c_2078_n 0.00433139f $X=6.98 $Y=0.58 $X2=0
+ $Y2=0
cc_735 N_A_995_74#_c_853_n N_VGND_c_2079_n 0.0135277f $X=8.345 $Y=1.12 $X2=0
+ $Y2=0
cc_736 N_A_995_74#_c_857_n N_VGND_c_2079_n 0.0561832f $X=7.835 $Y=0.99 $X2=0
+ $Y2=0
cc_737 N_A_995_74#_c_861_n N_VGND_c_2079_n 0.00421324f $X=8.345 $Y=1.285 $X2=0
+ $Y2=0
cc_738 N_SET_B_M1035_g N_A_594_74#_c_1143_n 0.0118199f $X=7.385 $Y=2.525 $X2=0
+ $Y2=0
cc_739 N_SET_B_c_985_n N_A_594_74#_M1003_g 5.49097e-19 $X=10.585 $Y=1.665 $X2=0
+ $Y2=0
cc_740 N_SET_B_c_986_n N_A_594_74#_M1003_g 4.75412e-19 $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_741 SET_B N_A_594_74#_M1003_g 6.71157e-19 $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_742 N_SET_B_c_985_n N_A_594_74#_c_1131_n 9.87584e-19 $X=10.585 $Y=1.665 $X2=0
+ $Y2=0
cc_743 N_SET_B_c_986_n N_A_594_74#_c_1131_n 0.00361779f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_744 SET_B N_A_594_74#_c_1131_n 7.37013e-19 $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_745 N_SET_B_c_982_n N_A_1924_48#_c_1299_n 0.00789413f $X=10.765 $Y=1.775
+ $X2=0 $Y2=0
cc_746 N_SET_B_c_983_n N_A_1924_48#_c_1299_n 8.51789e-19 $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_747 N_SET_B_c_985_n N_A_1924_48#_c_1299_n 0.0133161f $X=10.585 $Y=1.665 $X2=0
+ $Y2=0
cc_748 SET_B N_A_1924_48#_c_1299_n 0.0020819f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_749 N_SET_B_M1032_g N_A_1924_48#_c_1312_n 0.0247122f $X=10.89 $Y=2.75 $X2=0
+ $Y2=0
cc_750 N_SET_B_c_985_n N_A_1924_48#_c_1312_n 0.00262055f $X=10.585 $Y=1.665
+ $X2=0 $Y2=0
cc_751 N_SET_B_c_981_n N_A_1924_48#_c_1300_n 0.0101943f $X=10.31 $Y=0.94 $X2=0
+ $Y2=0
cc_752 N_SET_B_c_991_n N_A_1924_48#_c_1300_n 0.00487711f $X=10.75 $Y=1.255 $X2=0
+ $Y2=0
cc_753 N_SET_B_c_979_n N_A_1924_48#_c_1301_n 0.0212296f $X=10.235 $Y=0.865 $X2=0
+ $Y2=0
cc_754 N_SET_B_c_983_n N_A_1924_48#_c_1302_n 0.00158234f $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_755 N_SET_B_c_984_n N_A_1924_48#_c_1302_n 0.00789413f $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_756 N_SET_B_c_985_n N_A_1924_48#_c_1302_n 0.00419833f $X=10.585 $Y=1.665
+ $X2=0 $Y2=0
cc_757 N_SET_B_c_986_n N_A_1924_48#_c_1302_n 0.00205438f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_758 SET_B N_A_1924_48#_c_1302_n 0.00539133f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_759 N_SET_B_c_980_n N_A_1924_48#_c_1303_n 0.0117431f $X=10.55 $Y=0.94 $X2=0
+ $Y2=0
cc_760 N_SET_B_c_981_n N_A_1924_48#_c_1303_n 0.0106933f $X=10.31 $Y=0.94 $X2=0
+ $Y2=0
cc_761 N_SET_B_c_983_n N_A_1924_48#_c_1303_n 0.02412f $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_762 N_SET_B_c_984_n N_A_1924_48#_c_1303_n 0.00273565f $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_763 N_SET_B_c_985_n N_A_1924_48#_c_1303_n 0.0227767f $X=10.585 $Y=1.665 $X2=0
+ $Y2=0
cc_764 SET_B N_A_1924_48#_c_1303_n 6.64033e-19 $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_765 N_SET_B_c_991_n N_A_1924_48#_c_1303_n 0.00520213f $X=10.75 $Y=1.255 $X2=0
+ $Y2=0
cc_766 N_SET_B_c_983_n N_A_1924_48#_c_1305_n 0.00196616f $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_767 N_SET_B_c_991_n N_A_1924_48#_c_1305_n 9.74678e-19 $X=10.75 $Y=1.255 $X2=0
+ $Y2=0
cc_768 N_SET_B_c_983_n N_A_1924_48#_c_1307_n 0.00835006f $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_769 N_SET_B_c_984_n N_A_1924_48#_c_1307_n 6.8943e-19 $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_770 N_SET_B_M1032_g N_A_1924_48#_c_1315_n 8.9375e-19 $X=10.89 $Y=2.75 $X2=0
+ $Y2=0
cc_771 N_SET_B_c_985_n N_A_1924_48#_c_1345_n 0.00742107f $X=10.585 $Y=1.665
+ $X2=0 $Y2=0
cc_772 N_SET_B_c_986_n N_A_1924_48#_c_1345_n 0.00267727f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_773 SET_B N_A_1924_48#_c_1345_n 0.00653525f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_774 N_SET_B_c_991_n N_A_1924_48#_c_1345_n 8.32131e-19 $X=10.75 $Y=1.255 $X2=0
+ $Y2=0
cc_775 N_SET_B_c_979_n N_A_1762_74#_c_1428_n 0.00514966f $X=10.235 $Y=0.865
+ $X2=0 $Y2=0
cc_776 N_SET_B_c_983_n N_A_1762_74#_c_1429_n 0.00136743f $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_777 N_SET_B_c_984_n N_A_1762_74#_c_1429_n 0.01211f $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_778 N_SET_B_c_991_n N_A_1762_74#_c_1429_n 0.00524052f $X=10.75 $Y=1.255 $X2=0
+ $Y2=0
cc_779 N_SET_B_c_980_n N_A_1762_74#_c_1435_n 0.00859503f $X=10.55 $Y=0.94 $X2=0
+ $Y2=0
cc_780 N_SET_B_c_984_n N_A_1762_74#_c_1435_n 5.62189e-19 $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_781 N_SET_B_c_982_n N_A_1762_74#_c_1436_n 0.01211f $X=10.765 $Y=1.775 $X2=0
+ $Y2=0
cc_782 N_SET_B_c_995_n N_A_1762_74#_c_1436_n 0.0100137f $X=10.765 $Y=1.925 $X2=0
+ $Y2=0
cc_783 N_SET_B_c_983_n N_A_1762_74#_c_1436_n 2.72084e-19 $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_784 N_SET_B_c_985_n N_A_1762_74#_c_1453_n 0.0175055f $X=10.585 $Y=1.665 $X2=0
+ $Y2=0
cc_785 N_SET_B_c_986_n N_A_1762_74#_c_1453_n 0.0125497f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_786 SET_B N_A_1762_74#_c_1453_n 0.008126f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_787 N_SET_B_M1032_g N_A_1762_74#_c_1454_n 0.0199132f $X=10.89 $Y=2.75 $X2=0
+ $Y2=0
cc_788 N_SET_B_c_995_n N_A_1762_74#_c_1454_n 0.00251056f $X=10.765 $Y=1.925
+ $X2=0 $Y2=0
cc_789 N_SET_B_c_983_n N_A_1762_74#_c_1454_n 0.0257549f $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_790 N_SET_B_c_985_n N_A_1762_74#_c_1454_n 0.0207168f $X=10.585 $Y=1.665 $X2=0
+ $Y2=0
cc_791 N_SET_B_M1032_g N_A_1762_74#_c_1440_n 0.0102771f $X=10.89 $Y=2.75 $X2=0
+ $Y2=0
cc_792 N_SET_B_c_982_n N_A_1762_74#_c_1440_n 9.04429e-19 $X=10.765 $Y=1.775
+ $X2=0 $Y2=0
cc_793 N_SET_B_c_995_n N_A_1762_74#_c_1440_n 0.00657737f $X=10.765 $Y=1.925
+ $X2=0 $Y2=0
cc_794 N_SET_B_c_983_n N_A_1762_74#_c_1440_n 0.0192851f $X=10.75 $Y=1.42 $X2=0
+ $Y2=0
cc_795 N_SET_B_c_986_n N_A_1762_74#_c_1441_n 0.00926935f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_796 N_SET_B_c_986_n N_A_1762_74#_c_1456_n 0.00844651f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_797 N_SET_B_c_985_n N_A_1762_74#_c_1442_n 0.00721247f $X=10.585 $Y=1.665
+ $X2=0 $Y2=0
cc_798 N_SET_B_c_986_n N_A_1762_74#_c_1442_n 0.0193428f $X=9.695 $Y=1.665 $X2=0
+ $Y2=0
cc_799 SET_B N_A_1762_74#_c_1442_n 0.00234368f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_800 N_SET_B_M1032_g N_A_1762_74#_c_1458_n 0.00332493f $X=10.89 $Y=2.75 $X2=0
+ $Y2=0
cc_801 N_SET_B_c_985_n N_A_1762_74#_c_1458_n 0.0133991f $X=10.585 $Y=1.665 $X2=0
+ $Y2=0
cc_802 N_SET_B_M1032_g N_A_1762_74#_c_1459_n 0.0076098f $X=10.89 $Y=2.75 $X2=0
+ $Y2=0
cc_803 N_SET_B_c_986_n N_VPWR_M1035_d 0.00175187f $X=9.695 $Y=1.665 $X2=0 $Y2=0
cc_804 N_SET_B_c_990_n N_VPWR_M1035_d 0.00101131f $X=7.46 $Y=1.41 $X2=0 $Y2=0
cc_805 N_SET_B_M1035_g N_VPWR_c_1668_n 0.00395223f $X=7.385 $Y=2.525 $X2=0 $Y2=0
cc_806 N_SET_B_M1032_g N_VPWR_c_1669_n 0.0030528f $X=10.89 $Y=2.75 $X2=0 $Y2=0
cc_807 N_SET_B_M1032_g N_VPWR_c_1680_n 0.005209f $X=10.89 $Y=2.75 $X2=0 $Y2=0
cc_808 N_SET_B_M1032_g N_VPWR_c_1662_n 0.00987509f $X=10.89 $Y=2.75 $X2=0 $Y2=0
cc_809 N_SET_B_c_986_n N_A_1603_347#_M1041_d 0.00228324f $X=9.695 $Y=1.665
+ $X2=-0.19 $Y2=-0.245
cc_810 N_SET_B_c_986_n N_A_1603_347#_c_1946_n 0.00581237f $X=9.695 $Y=1.665
+ $X2=0 $Y2=0
cc_811 N_SET_B_c_979_n N_VGND_c_2071_n 0.00384553f $X=10.235 $Y=0.865 $X2=0
+ $Y2=0
cc_812 N_SET_B_M1014_g N_VGND_c_2075_n 0.00913019f $X=7.37 $Y=0.58 $X2=0 $Y2=0
cc_813 N_SET_B_c_979_n N_VGND_c_2075_n 0.00758569f $X=10.235 $Y=0.865 $X2=0
+ $Y2=0
cc_814 N_SET_B_M1014_g N_VGND_c_2078_n 0.00461464f $X=7.37 $Y=0.58 $X2=0 $Y2=0
cc_815 N_SET_B_M1014_g N_VGND_c_2079_n 0.00576207f $X=7.37 $Y=0.58 $X2=0 $Y2=0
cc_816 N_SET_B_c_979_n N_VGND_c_2080_n 0.0127134f $X=10.235 $Y=0.865 $X2=0 $Y2=0
cc_817 N_SET_B_c_980_n N_VGND_c_2080_n 0.00878086f $X=10.55 $Y=0.94 $X2=0 $Y2=0
cc_818 N_A_594_74#_M1003_g N_A_1924_48#_c_1299_n 0.00544029f $X=9.305 $Y=0.58
+ $X2=0 $Y2=0
cc_819 N_A_594_74#_c_1131_n N_A_1924_48#_c_1299_n 0.0120712f $X=9.44 $Y=1.795
+ $X2=0 $Y2=0
cc_820 N_A_594_74#_M1008_g N_A_1924_48#_c_1313_n 0.0120712f $X=9.44 $Y=2.37
+ $X2=0 $Y2=0
cc_821 N_A_594_74#_M1003_g N_A_1924_48#_c_1301_n 0.06105f $X=9.305 $Y=0.58 $X2=0
+ $Y2=0
cc_822 N_A_594_74#_M1003_g N_A_1924_48#_c_1345_n 0.00104919f $X=9.305 $Y=0.58
+ $X2=0 $Y2=0
cc_823 N_A_594_74#_M1008_g N_A_1762_74#_c_1453_n 0.00985565f $X=9.44 $Y=2.37
+ $X2=0 $Y2=0
cc_824 N_A_594_74#_M1003_g N_A_1762_74#_c_1441_n 0.0256745f $X=9.305 $Y=0.58
+ $X2=0 $Y2=0
cc_825 N_A_594_74#_M1008_g N_A_1762_74#_c_1456_n 0.00487272f $X=9.44 $Y=2.37
+ $X2=0 $Y2=0
cc_826 N_A_594_74#_M1003_g N_A_1762_74#_c_1442_n 0.0174369f $X=9.305 $Y=0.58
+ $X2=0 $Y2=0
cc_827 N_A_594_74#_c_1131_n N_A_1762_74#_c_1442_n 0.0065831f $X=9.44 $Y=1.795
+ $X2=0 $Y2=0
cc_828 N_A_594_74#_M1008_g N_A_1762_74#_c_1442_n 0.00178445f $X=9.44 $Y=2.37
+ $X2=0 $Y2=0
cc_829 N_A_594_74#_M1008_g N_A_1762_74#_c_1458_n 6.92524e-19 $X=9.44 $Y=2.37
+ $X2=0 $Y2=0
cc_830 N_A_594_74#_c_1149_n N_VPWR_M1026_d 0.00184478f $X=3.885 $Y=1.905 $X2=0
+ $Y2=0
cc_831 N_A_594_74#_M1030_g N_VPWR_c_1666_n 0.00786105f $X=3.965 $Y=2.4 $X2=0
+ $Y2=0
cc_832 N_A_594_74#_c_1141_n N_VPWR_c_1666_n 0.00246093f $X=4.55 $Y=3.15 $X2=0
+ $Y2=0
cc_833 N_A_594_74#_M1020_g N_VPWR_c_1667_n 0.00144272f $X=5.59 $Y=2.6 $X2=0
+ $Y2=0
cc_834 N_A_594_74#_c_1143_n N_VPWR_c_1667_n 0.0211465f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_835 N_A_594_74#_c_1143_n N_VPWR_c_1668_n 0.0170937f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_836 N_A_594_74#_M1030_g N_VPWR_c_1672_n 0.00460063f $X=3.965 $Y=2.4 $X2=0
+ $Y2=0
cc_837 N_A_594_74#_c_1141_n N_VPWR_c_1672_n 0.0434218f $X=4.55 $Y=3.15 $X2=0
+ $Y2=0
cc_838 N_A_594_74#_c_1143_n N_VPWR_c_1674_n 0.0290731f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_839 N_A_594_74#_c_1143_n N_VPWR_c_1676_n 0.0437144f $X=9.35 $Y=3.15 $X2=0
+ $Y2=0
cc_840 N_A_594_74#_M1030_g N_VPWR_c_1662_n 0.0090927f $X=3.965 $Y=2.4 $X2=0
+ $Y2=0
cc_841 N_A_594_74#_c_1140_n N_VPWR_c_1662_n 0.0223434f $X=5.5 $Y=3.15 $X2=0
+ $Y2=0
cc_842 N_A_594_74#_c_1141_n N_VPWR_c_1662_n 0.00599845f $X=4.55 $Y=3.15 $X2=0
+ $Y2=0
cc_843 N_A_594_74#_c_1143_n N_VPWR_c_1662_n 0.10486f $X=9.35 $Y=3.15 $X2=0 $Y2=0
cc_844 N_A_594_74#_c_1146_n N_VPWR_c_1662_n 0.00445012f $X=5.59 $Y=3.15 $X2=0
+ $Y2=0
cc_845 N_A_594_74#_c_1137_n N_A_293_464#_c_1819_n 0.00564313f $X=3.067 $Y=1.01
+ $X2=0 $Y2=0
cc_846 N_A_594_74#_c_1134_n N_A_293_464#_c_1821_n 0.00146536f $X=3.02 $Y=1.82
+ $X2=0 $Y2=0
cc_847 N_A_594_74#_M1026_s N_A_293_464#_c_1825_n 0.00758929f $X=3.15 $Y=1.84
+ $X2=0 $Y2=0
cc_848 N_A_594_74#_c_1148_n N_A_293_464#_c_1825_n 0.014265f $X=3.105 $Y=1.985
+ $X2=0 $Y2=0
cc_849 N_A_594_74#_c_1149_n N_A_293_464#_c_1825_n 0.00595683f $X=3.885 $Y=1.905
+ $X2=0 $Y2=0
cc_850 N_A_594_74#_c_1151_n N_A_293_464#_c_1825_n 0.0222509f $X=3.29 $Y=1.985
+ $X2=0 $Y2=0
cc_851 N_A_594_74#_M1030_g N_A_293_464#_c_1826_n 0.0161063f $X=3.965 $Y=2.4
+ $X2=0 $Y2=0
cc_852 N_A_594_74#_c_1126_n N_A_293_464#_c_1826_n 0.00236726f $X=4.4 $Y=1.385
+ $X2=0 $Y2=0
cc_853 N_A_594_74#_c_1127_n N_A_293_464#_c_1826_n 0.00393837f $X=4.475 $Y=3.075
+ $X2=0 $Y2=0
cc_854 N_A_594_74#_c_1149_n N_A_293_464#_c_1826_n 0.0193151f $X=3.885 $Y=1.905
+ $X2=0 $Y2=0
cc_855 N_A_594_74#_c_1124_n N_A_293_464#_c_1822_n 0.00100658f $X=3.83 $Y=1.22
+ $X2=0 $Y2=0
cc_856 N_A_594_74#_M1030_g N_A_293_464#_c_1822_n 0.00173466f $X=3.965 $Y=2.4
+ $X2=0 $Y2=0
cc_857 N_A_594_74#_c_1127_n N_A_293_464#_c_1822_n 0.0157324f $X=4.475 $Y=3.075
+ $X2=0 $Y2=0
cc_858 N_A_594_74#_c_1128_n N_A_293_464#_c_1822_n 0.00466065f $X=4.825 $Y=1.055
+ $X2=0 $Y2=0
cc_859 N_A_594_74#_M1037_g N_A_293_464#_c_1822_n 0.00101293f $X=4.9 $Y=0.58
+ $X2=0 $Y2=0
cc_860 N_A_594_74#_c_1132_n N_A_293_464#_c_1822_n 0.0200212f $X=4.475 $Y=1.055
+ $X2=0 $Y2=0
cc_861 N_A_594_74#_c_1149_n N_A_293_464#_c_1822_n 0.011652f $X=3.885 $Y=1.905
+ $X2=0 $Y2=0
cc_862 N_A_594_74#_c_1135_n N_A_293_464#_c_1822_n 0.0379515f $X=4.05 $Y=1.385
+ $X2=0 $Y2=0
cc_863 N_A_594_74#_c_1127_n N_A_293_464#_c_1828_n 0.00662564f $X=4.475 $Y=3.075
+ $X2=0 $Y2=0
cc_864 N_A_594_74#_M1030_g N_A_293_464#_c_1914_n 0.00283204f $X=3.965 $Y=2.4
+ $X2=0 $Y2=0
cc_865 N_A_594_74#_c_1149_n N_A_293_464#_c_1914_n 0.00826352f $X=3.885 $Y=1.905
+ $X2=0 $Y2=0
cc_866 N_A_594_74#_c_1128_n N_A_293_464#_c_1823_n 0.00424734f $X=4.825 $Y=1.055
+ $X2=0 $Y2=0
cc_867 N_A_594_74#_M1037_g N_A_293_464#_c_1823_n 0.00662014f $X=4.9 $Y=0.58
+ $X2=0 $Y2=0
cc_868 N_A_594_74#_c_1132_n N_A_293_464#_c_1823_n 0.00145165f $X=4.475 $Y=1.055
+ $X2=0 $Y2=0
cc_869 N_A_594_74#_c_1127_n N_A_293_464#_c_1829_n 0.00791487f $X=4.475 $Y=3.075
+ $X2=0 $Y2=0
cc_870 N_A_594_74#_c_1143_n N_A_1603_347#_c_1946_n 0.00686321f $X=9.35 $Y=3.15
+ $X2=0 $Y2=0
cc_871 N_A_594_74#_c_1131_n N_A_1603_347#_c_1946_n 3.12245e-19 $X=9.44 $Y=1.795
+ $X2=0 $Y2=0
cc_872 N_A_594_74#_M1008_g N_A_1603_347#_c_1946_n 0.0127656f $X=9.44 $Y=2.37
+ $X2=0 $Y2=0
cc_873 N_A_594_74#_c_1143_n N_A_1603_347#_c_1947_n 0.00598911f $X=9.35 $Y=3.15
+ $X2=0 $Y2=0
cc_874 N_A_594_74#_c_1143_n N_A_1712_374#_c_1980_n 0.00796669f $X=9.35 $Y=3.15
+ $X2=0 $Y2=0
cc_875 N_A_594_74#_M1008_g N_A_1712_374#_c_1980_n 0.0160595f $X=9.44 $Y=2.37
+ $X2=0 $Y2=0
cc_876 N_A_594_74#_M1008_g N_A_1712_374#_c_1981_n 0.00481013f $X=9.44 $Y=2.37
+ $X2=0 $Y2=0
cc_877 N_A_594_74#_c_1143_n N_A_1712_374#_c_1982_n 0.00738175f $X=9.35 $Y=3.15
+ $X2=0 $Y2=0
cc_878 N_A_594_74#_M1008_g N_A_1712_374#_c_1982_n 0.00623466f $X=9.44 $Y=2.37
+ $X2=0 $Y2=0
cc_879 N_A_594_74#_c_1133_n N_VGND_c_2060_n 0.0237473f $X=3.115 $Y=0.505 $X2=0
+ $Y2=0
cc_880 N_A_594_74#_c_1124_n N_VGND_c_2061_n 0.00470925f $X=3.83 $Y=1.22 $X2=0
+ $Y2=0
cc_881 N_A_594_74#_c_1133_n N_VGND_c_2061_n 0.0251347f $X=3.115 $Y=0.505 $X2=0
+ $Y2=0
cc_882 N_A_594_74#_c_1124_n N_VGND_c_2067_n 0.00430908f $X=3.83 $Y=1.22 $X2=0
+ $Y2=0
cc_883 N_A_594_74#_M1037_g N_VGND_c_2067_n 0.00278159f $X=4.9 $Y=0.58 $X2=0
+ $Y2=0
cc_884 N_A_594_74#_c_1133_n N_VGND_c_2070_n 0.0122205f $X=3.115 $Y=0.505 $X2=0
+ $Y2=0
cc_885 N_A_594_74#_M1003_g N_VGND_c_2071_n 0.00292646f $X=9.305 $Y=0.58 $X2=0
+ $Y2=0
cc_886 N_A_594_74#_c_1124_n N_VGND_c_2075_n 0.00821169f $X=3.83 $Y=1.22 $X2=0
+ $Y2=0
cc_887 N_A_594_74#_M1037_g N_VGND_c_2075_n 0.00359882f $X=4.9 $Y=0.58 $X2=0
+ $Y2=0
cc_888 N_A_594_74#_M1003_g N_VGND_c_2075_n 0.00359032f $X=9.305 $Y=0.58 $X2=0
+ $Y2=0
cc_889 N_A_594_74#_c_1133_n N_VGND_c_2075_n 0.00976972f $X=3.115 $Y=0.505 $X2=0
+ $Y2=0
cc_890 N_A_1924_48#_c_1304_n N_A_1762_74#_c_1428_n 0.0142415f $X=11.23 $Y=0.58
+ $X2=0 $Y2=0
cc_891 N_A_1924_48#_c_1305_n N_A_1762_74#_c_1429_n 0.00858132f $X=11.31 $Y=1.3
+ $X2=0 $Y2=0
cc_892 N_A_1924_48#_c_1307_n N_A_1762_74#_c_1429_n 0.0084379f $X=11.395 $Y=1.385
+ $X2=0 $Y2=0
cc_893 N_A_1924_48#_c_1308_n N_A_1762_74#_c_1429_n 6.40251e-19 $X=12.15 $Y=2.18
+ $X2=0 $Y2=0
cc_894 N_A_1924_48#_c_1310_n N_A_1762_74#_c_1429_n 0.00224676f $X=11.23 $Y=0.985
+ $X2=0 $Y2=0
cc_895 N_A_1924_48#_c_1315_n N_A_1762_74#_M1029_g 0.00860477f $X=11.665 $Y=2.75
+ $X2=0 $Y2=0
cc_896 N_A_1924_48#_c_1316_n N_A_1762_74#_M1029_g 0.0201094f $X=12.065 $Y=2.265
+ $X2=0 $Y2=0
cc_897 N_A_1924_48#_c_1305_n N_A_1762_74#_M1009_g 0.00247796f $X=11.31 $Y=1.3
+ $X2=0 $Y2=0
cc_898 N_A_1924_48#_c_1306_n N_A_1762_74#_M1009_g 0.0175404f $X=12.065 $Y=1.385
+ $X2=0 $Y2=0
cc_899 N_A_1924_48#_c_1308_n N_A_1762_74#_M1009_g 0.00604112f $X=12.15 $Y=2.18
+ $X2=0 $Y2=0
cc_900 N_A_1924_48#_c_1308_n N_A_1762_74#_c_1431_n 0.00497859f $X=12.15 $Y=2.18
+ $X2=0 $Y2=0
cc_901 N_A_1924_48#_c_1306_n N_A_1762_74#_c_1432_n 8.5035e-19 $X=12.065 $Y=1.385
+ $X2=0 $Y2=0
cc_902 N_A_1924_48#_c_1316_n N_A_1762_74#_c_1432_n 7.87495e-19 $X=12.065
+ $Y=2.265 $X2=0 $Y2=0
cc_903 N_A_1924_48#_c_1308_n N_A_1762_74#_c_1432_n 0.0127667f $X=12.15 $Y=2.18
+ $X2=0 $Y2=0
cc_904 N_A_1924_48#_c_1316_n N_A_1762_74#_c_1446_n 0.00161327f $X=12.065
+ $Y=2.265 $X2=0 $Y2=0
cc_905 N_A_1924_48#_c_1308_n N_A_1762_74#_c_1446_n 0.00347689f $X=12.15 $Y=2.18
+ $X2=0 $Y2=0
cc_906 N_A_1924_48#_c_1303_n N_A_1762_74#_c_1435_n 0.00958405f $X=11.065
+ $Y=0.985 $X2=0 $Y2=0
cc_907 N_A_1924_48#_c_1304_n N_A_1762_74#_c_1435_n 0.00829222f $X=11.23 $Y=0.58
+ $X2=0 $Y2=0
cc_908 N_A_1924_48#_c_1310_n N_A_1762_74#_c_1435_n 0.00686615f $X=11.23 $Y=0.985
+ $X2=0 $Y2=0
cc_909 N_A_1924_48#_c_1306_n N_A_1762_74#_c_1437_n 0.0110481f $X=12.065 $Y=1.385
+ $X2=0 $Y2=0
cc_910 N_A_1924_48#_c_1316_n N_A_1762_74#_c_1437_n 0.00108592f $X=12.065
+ $Y=2.265 $X2=0 $Y2=0
cc_911 N_A_1924_48#_c_1317_n N_A_1762_74#_c_1437_n 0.00578596f $X=11.75 $Y=2.265
+ $X2=0 $Y2=0
cc_912 N_A_1924_48#_c_1299_n N_A_1762_74#_c_1453_n 0.0110264f $X=9.955 $Y=2.165
+ $X2=0 $Y2=0
cc_913 N_A_1924_48#_c_1302_n N_A_1762_74#_c_1453_n 0.00311771f $X=9.825 $Y=1.405
+ $X2=0 $Y2=0
cc_914 N_A_1924_48#_c_1299_n N_A_1762_74#_c_1454_n 3.79939e-19 $X=9.955 $Y=2.165
+ $X2=0 $Y2=0
cc_915 N_A_1924_48#_c_1312_n N_A_1762_74#_c_1454_n 0.0193659f $X=10.35 $Y=2.24
+ $X2=0 $Y2=0
cc_916 N_A_1924_48#_c_1307_n N_A_1762_74#_c_1440_n 0.00457115f $X=11.395
+ $Y=1.385 $X2=0 $Y2=0
cc_917 N_A_1924_48#_c_1317_n N_A_1762_74#_c_1440_n 0.0119447f $X=11.75 $Y=2.265
+ $X2=0 $Y2=0
cc_918 N_A_1924_48#_c_1310_n N_A_1762_74#_c_1440_n 0.00460453f $X=11.23 $Y=0.985
+ $X2=0 $Y2=0
cc_919 N_A_1924_48#_c_1306_n N_A_1762_74#_c_1536_n 0.0375032f $X=12.065 $Y=1.385
+ $X2=0 $Y2=0
cc_920 N_A_1924_48#_c_1307_n N_A_1762_74#_c_1536_n 0.00923271f $X=11.395
+ $Y=1.385 $X2=0 $Y2=0
cc_921 N_A_1924_48#_c_1316_n N_A_1762_74#_c_1536_n 0.0088719f $X=12.065 $Y=2.265
+ $X2=0 $Y2=0
cc_922 N_A_1924_48#_c_1317_n N_A_1762_74#_c_1536_n 0.0179959f $X=11.75 $Y=2.265
+ $X2=0 $Y2=0
cc_923 N_A_1924_48#_c_1308_n N_A_1762_74#_c_1536_n 0.0253686f $X=12.15 $Y=2.18
+ $X2=0 $Y2=0
cc_924 N_A_1924_48#_c_1301_n N_A_1762_74#_c_1441_n 0.00300533f $X=9.785 $Y=0.865
+ $X2=0 $Y2=0
cc_925 N_A_1924_48#_c_1345_n N_A_1762_74#_c_1441_n 0.0189516f $X=9.785 $Y=0.985
+ $X2=0 $Y2=0
cc_926 N_A_1924_48#_c_1299_n N_A_1762_74#_c_1456_n 2.64746e-19 $X=9.955 $Y=2.165
+ $X2=0 $Y2=0
cc_927 N_A_1924_48#_c_1299_n N_A_1762_74#_c_1442_n 0.00183767f $X=9.955 $Y=2.165
+ $X2=0 $Y2=0
cc_928 N_A_1924_48#_c_1309_n N_A_1762_74#_c_1442_n 0.00300533f $X=9.785 $Y=1.065
+ $X2=0 $Y2=0
cc_929 N_A_1924_48#_c_1299_n N_A_1762_74#_c_1458_n 0.00593027f $X=9.955 $Y=2.165
+ $X2=0 $Y2=0
cc_930 N_A_1924_48#_c_1312_n N_A_1762_74#_c_1458_n 0.00552372f $X=10.35 $Y=2.24
+ $X2=0 $Y2=0
cc_931 N_A_1924_48#_c_1313_n N_A_1762_74#_c_1458_n 0.00237768f $X=10.03 $Y=2.24
+ $X2=0 $Y2=0
cc_932 N_A_1924_48#_c_1315_n N_A_1762_74#_c_1460_n 0.0422692f $X=11.665 $Y=2.75
+ $X2=0 $Y2=0
cc_933 N_A_1924_48#_c_1316_n N_VPWR_M1029_d 0.00437093f $X=12.065 $Y=2.265 $X2=0
+ $Y2=0
cc_934 N_A_1924_48#_c_1308_n N_VPWR_M1029_d 0.00764262f $X=12.15 $Y=2.18 $X2=0
+ $Y2=0
cc_935 N_A_1924_48#_M1028_g N_VPWR_c_1669_n 0.0014827f $X=10.44 $Y=2.75 $X2=0
+ $Y2=0
cc_936 N_A_1924_48#_c_1315_n N_VPWR_c_1670_n 0.0165069f $X=11.665 $Y=2.75 $X2=0
+ $Y2=0
cc_937 N_A_1924_48#_c_1316_n N_VPWR_c_1670_n 0.0245581f $X=12.065 $Y=2.265 $X2=0
+ $Y2=0
cc_938 N_A_1924_48#_M1028_g N_VPWR_c_1676_n 0.00517089f $X=10.44 $Y=2.75 $X2=0
+ $Y2=0
cc_939 N_A_1924_48#_c_1315_n N_VPWR_c_1680_n 0.011066f $X=11.665 $Y=2.75 $X2=0
+ $Y2=0
cc_940 N_A_1924_48#_M1028_g N_VPWR_c_1662_n 0.00982721f $X=10.44 $Y=2.75 $X2=0
+ $Y2=0
cc_941 N_A_1924_48#_c_1315_n N_VPWR_c_1662_n 0.00915947f $X=11.665 $Y=2.75 $X2=0
+ $Y2=0
cc_942 N_A_1924_48#_c_1313_n N_A_1603_347#_c_1948_n 7.20281e-19 $X=10.03 $Y=2.24
+ $X2=0 $Y2=0
cc_943 N_A_1924_48#_M1028_g N_A_1603_347#_c_1948_n 0.00560766f $X=10.44 $Y=2.75
+ $X2=0 $Y2=0
cc_944 N_A_1924_48#_c_1313_n N_A_1712_374#_c_1980_n 0.00406826f $X=10.03 $Y=2.24
+ $X2=0 $Y2=0
cc_945 N_A_1924_48#_M1028_g N_A_1712_374#_c_1980_n 0.00532912f $X=10.44 $Y=2.75
+ $X2=0 $Y2=0
cc_946 N_A_1924_48#_c_1312_n N_A_1712_374#_c_1981_n 0.00603289f $X=10.35 $Y=2.24
+ $X2=0 $Y2=0
cc_947 N_A_1924_48#_M1028_g N_A_1712_374#_c_1981_n 0.00578543f $X=10.44 $Y=2.75
+ $X2=0 $Y2=0
cc_948 N_A_1924_48#_c_1316_n N_Q_N_c_2015_n 0.0115069f $X=12.065 $Y=2.265 $X2=0
+ $Y2=0
cc_949 N_A_1924_48#_c_1306_n N_Q_N_c_2011_n 0.0121685f $X=12.065 $Y=1.385 $X2=0
+ $Y2=0
cc_950 N_A_1924_48#_c_1308_n N_Q_N_c_2011_n 0.0426161f $X=12.15 $Y=2.18 $X2=0
+ $Y2=0
cc_951 N_A_1924_48#_c_1306_n Q_N 0.00999592f $X=12.065 $Y=1.385 $X2=0 $Y2=0
cc_952 N_A_1924_48#_c_1304_n N_VGND_c_2063_n 0.0370462f $X=11.23 $Y=0.58 $X2=0
+ $Y2=0
cc_953 N_A_1924_48#_c_1305_n N_VGND_c_2063_n 0.00382008f $X=11.31 $Y=1.3 $X2=0
+ $Y2=0
cc_954 N_A_1924_48#_c_1306_n N_VGND_c_2063_n 0.0277028f $X=12.065 $Y=1.385 $X2=0
+ $Y2=0
cc_955 N_A_1924_48#_c_1310_n N_VGND_c_2063_n 0.0121589f $X=11.23 $Y=0.985 $X2=0
+ $Y2=0
cc_956 N_A_1924_48#_c_1301_n N_VGND_c_2071_n 0.00461464f $X=9.785 $Y=0.865 $X2=0
+ $Y2=0
cc_957 N_A_1924_48#_c_1304_n N_VGND_c_2072_n 0.0145931f $X=11.23 $Y=0.58 $X2=0
+ $Y2=0
cc_958 N_A_1924_48#_c_1300_n N_VGND_c_2075_n 0.00441445f $X=9.785 $Y=1.03 $X2=0
+ $Y2=0
cc_959 N_A_1924_48#_c_1301_n N_VGND_c_2075_n 0.00910057f $X=9.785 $Y=0.865 $X2=0
+ $Y2=0
cc_960 N_A_1924_48#_c_1304_n N_VGND_c_2075_n 0.0120099f $X=11.23 $Y=0.58 $X2=0
+ $Y2=0
cc_961 N_A_1924_48#_c_1301_n N_VGND_c_2080_n 0.00203578f $X=9.785 $Y=0.865 $X2=0
+ $Y2=0
cc_962 N_A_1924_48#_c_1303_n N_VGND_c_2080_n 0.0374282f $X=11.065 $Y=0.985 $X2=0
+ $Y2=0
cc_963 N_A_1924_48#_c_1304_n N_VGND_c_2080_n 0.0132497f $X=11.23 $Y=0.58 $X2=0
+ $Y2=0
cc_964 N_A_1762_74#_M1018_g N_A_2556_112#_M1031_g 0.00350851f $X=13.14 $Y=0.835
+ $X2=0 $Y2=0
cc_965 N_A_1762_74#_c_1439_n N_A_2556_112#_M1031_g 0.0163785f $X=13.14 $Y=1.79
+ $X2=0 $Y2=0
cc_966 N_A_1762_74#_M1018_g N_A_2556_112#_c_1616_n 0.0093401f $X=13.14 $Y=0.835
+ $X2=0 $Y2=0
cc_967 N_A_1762_74#_M1018_g N_A_2556_112#_c_1617_n 0.0181387f $X=13.14 $Y=0.835
+ $X2=0 $Y2=0
cc_968 N_A_1762_74#_c_1439_n N_A_2556_112#_c_1617_n 0.00172362f $X=13.14 $Y=1.79
+ $X2=0 $Y2=0
cc_969 N_A_1762_74#_M1009_g N_A_2556_112#_c_1619_n 9.40127e-19 $X=12.075 $Y=0.74
+ $X2=0 $Y2=0
cc_970 N_A_1762_74#_c_1433_n N_A_2556_112#_c_1619_n 0.00388219f $X=13.065
+ $Y=1.69 $X2=0 $Y2=0
cc_971 N_A_1762_74#_M1018_g N_A_2556_112#_c_1619_n 0.0367305f $X=13.14 $Y=0.835
+ $X2=0 $Y2=0
cc_972 N_A_1762_74#_c_1446_n N_A_2556_112#_c_1620_n 0.00255732f $X=12.395
+ $Y=1.765 $X2=0 $Y2=0
cc_973 N_A_1762_74#_c_1433_n N_A_2556_112#_c_1620_n 0.00554698f $X=13.065
+ $Y=1.69 $X2=0 $Y2=0
cc_974 N_A_1762_74#_M1018_g N_A_2556_112#_c_1620_n 0.00246233f $X=13.14 $Y=0.835
+ $X2=0 $Y2=0
cc_975 N_A_1762_74#_c_1448_n N_A_2556_112#_c_1620_n 0.00642329f $X=13.395
+ $Y=1.94 $X2=0 $Y2=0
cc_976 N_A_1762_74#_c_1439_n N_A_2556_112#_c_1620_n 0.0170146f $X=13.14 $Y=1.79
+ $X2=0 $Y2=0
cc_977 N_A_1762_74#_c_1439_n N_A_2556_112#_c_1621_n 0.00801933f $X=13.14 $Y=1.79
+ $X2=0 $Y2=0
cc_978 N_A_1762_74#_c_1454_n N_VPWR_c_1669_n 0.0106837f $X=11.11 $Y=2.18 $X2=0
+ $Y2=0
cc_979 N_A_1762_74#_c_1459_n N_VPWR_c_1669_n 0.01643f $X=11.115 $Y=2.75 $X2=0
+ $Y2=0
cc_980 N_A_1762_74#_M1029_g N_VPWR_c_1670_n 0.01359f $X=11.89 $Y=2.75 $X2=0
+ $Y2=0
cc_981 N_A_1762_74#_c_1446_n N_VPWR_c_1670_n 0.00359954f $X=12.395 $Y=1.765
+ $X2=0 $Y2=0
cc_982 N_A_1762_74#_c_1448_n N_VPWR_c_1671_n 0.0204993f $X=13.395 $Y=1.94 $X2=0
+ $Y2=0
cc_983 N_A_1762_74#_M1029_g N_VPWR_c_1680_n 0.00460063f $X=11.89 $Y=2.75 $X2=0
+ $Y2=0
cc_984 N_A_1762_74#_c_1459_n N_VPWR_c_1680_n 0.0143566f $X=11.115 $Y=2.75 $X2=0
+ $Y2=0
cc_985 N_A_1762_74#_c_1446_n N_VPWR_c_1681_n 0.00515235f $X=12.395 $Y=1.765
+ $X2=0 $Y2=0
cc_986 N_A_1762_74#_c_1448_n N_VPWR_c_1681_n 0.00502645f $X=13.395 $Y=1.94 $X2=0
+ $Y2=0
cc_987 N_A_1762_74#_M1029_g N_VPWR_c_1662_n 0.00913687f $X=11.89 $Y=2.75 $X2=0
+ $Y2=0
cc_988 N_A_1762_74#_c_1446_n N_VPWR_c_1662_n 0.0096903f $X=12.395 $Y=1.765 $X2=0
+ $Y2=0
cc_989 N_A_1762_74#_c_1448_n N_VPWR_c_1662_n 0.00516335f $X=13.395 $Y=1.94 $X2=0
+ $Y2=0
cc_990 N_A_1762_74#_c_1459_n N_VPWR_c_1662_n 0.011899f $X=11.115 $Y=2.75 $X2=0
+ $Y2=0
cc_991 N_A_1762_74#_c_1453_n N_A_1603_347#_M1008_d 0.00405263f $X=10 $Y=2.035
+ $X2=0 $Y2=0
cc_992 N_A_1762_74#_M1033_d N_A_1603_347#_c_1946_n 0.00460527f $X=8.99 $Y=1.87
+ $X2=0 $Y2=0
cc_993 N_A_1762_74#_c_1453_n N_A_1603_347#_c_1946_n 0.00755336f $X=10 $Y=2.035
+ $X2=0 $Y2=0
cc_994 N_A_1762_74#_c_1456_n N_A_1603_347#_c_1946_n 0.0210899f $X=9.21 $Y=2.015
+ $X2=0 $Y2=0
cc_995 N_A_1762_74#_c_1453_n N_A_1603_347#_c_1948_n 0.0184544f $X=10 $Y=2.035
+ $X2=0 $Y2=0
cc_996 N_A_1762_74#_c_1458_n N_A_1712_374#_c_1980_n 0.00131213f $X=10.085
+ $Y=2.035 $X2=0 $Y2=0
cc_997 N_A_1762_74#_c_1454_n N_A_1712_374#_c_1981_n 0.0120968f $X=11.11 $Y=2.18
+ $X2=0 $Y2=0
cc_998 N_A_1762_74#_c_1458_n N_A_1712_374#_c_1981_n 0.00723033f $X=10.085
+ $Y=2.035 $X2=0 $Y2=0
cc_999 N_A_1762_74#_c_1446_n N_Q_N_c_2014_n 0.00188854f $X=12.395 $Y=1.765 $X2=0
+ $Y2=0
cc_1000 N_A_1762_74#_c_1433_n N_Q_N_c_2014_n 0.00391459f $X=13.065 $Y=1.69 $X2=0
+ $Y2=0
cc_1001 N_A_1762_74#_c_1448_n N_Q_N_c_2014_n 0.00421522f $X=13.395 $Y=1.94 $X2=0
+ $Y2=0
cc_1002 N_A_1762_74#_c_1439_n N_Q_N_c_2014_n 4.52148e-19 $X=13.14 $Y=1.79 $X2=0
+ $Y2=0
cc_1003 N_A_1762_74#_M1029_g N_Q_N_c_2015_n 0.00112542f $X=11.89 $Y=2.75 $X2=0
+ $Y2=0
cc_1004 N_A_1762_74#_c_1446_n N_Q_N_c_2015_n 0.0154106f $X=12.395 $Y=1.765 $X2=0
+ $Y2=0
cc_1005 N_A_1762_74#_M1009_g N_Q_N_c_2011_n 0.00681469f $X=12.075 $Y=0.74 $X2=0
+ $Y2=0
cc_1006 N_A_1762_74#_c_1446_n N_Q_N_c_2011_n 0.00133028f $X=12.395 $Y=1.765
+ $X2=0 $Y2=0
cc_1007 N_A_1762_74#_c_1433_n N_Q_N_c_2011_n 0.0115f $X=13.065 $Y=1.69 $X2=0
+ $Y2=0
cc_1008 N_A_1762_74#_c_1438_n N_Q_N_c_2011_n 0.00365808f $X=12.395 $Y=1.69 $X2=0
+ $Y2=0
cc_1009 N_A_1762_74#_M1009_g Q_N 0.00766778f $X=12.075 $Y=0.74 $X2=0 $Y2=0
cc_1010 N_A_1762_74#_M1018_g Q_N 0.00756882f $X=13.14 $Y=0.835 $X2=0 $Y2=0
cc_1011 N_A_1762_74#_M1009_g Q_N 0.0034024f $X=12.075 $Y=0.74 $X2=0 $Y2=0
cc_1012 N_A_1762_74#_c_1431_n Q_N 0.00728143f $X=12.305 $Y=1.69 $X2=0 $Y2=0
cc_1013 N_A_1762_74#_c_1448_n Q 3.68595e-19 $X=13.395 $Y=1.94 $X2=0 $Y2=0
cc_1014 N_A_1762_74#_c_1439_n Q 0.00103644f $X=13.14 $Y=1.79 $X2=0 $Y2=0
cc_1015 N_A_1762_74#_c_1428_n N_VGND_c_2063_n 0.00389959f $X=11.015 $Y=0.865
+ $X2=0 $Y2=0
cc_1016 N_A_1762_74#_M1009_g N_VGND_c_2063_n 0.0169409f $X=12.075 $Y=0.74 $X2=0
+ $Y2=0
cc_1017 N_A_1762_74#_c_1435_n N_VGND_c_2063_n 0.00114561f $X=11.3 $Y=0.94 $X2=0
+ $Y2=0
cc_1018 N_A_1762_74#_M1018_g N_VGND_c_2064_n 0.0047492f $X=13.14 $Y=0.835 $X2=0
+ $Y2=0
cc_1019 N_A_1762_74#_c_1441_n N_VGND_c_2071_n 0.025983f $X=9.09 $Y=0.515 $X2=0
+ $Y2=0
cc_1020 N_A_1762_74#_c_1428_n N_VGND_c_2072_n 0.00434272f $X=11.015 $Y=0.865
+ $X2=0 $Y2=0
cc_1021 N_A_1762_74#_M1009_g N_VGND_c_2073_n 0.00434272f $X=12.075 $Y=0.74 $X2=0
+ $Y2=0
cc_1022 N_A_1762_74#_M1018_g N_VGND_c_2073_n 0.00340575f $X=13.14 $Y=0.835 $X2=0
+ $Y2=0
cc_1023 N_A_1762_74#_c_1428_n N_VGND_c_2075_n 0.00827575f $X=11.015 $Y=0.865
+ $X2=0 $Y2=0
cc_1024 N_A_1762_74#_M1009_g N_VGND_c_2075_n 0.00830058f $X=12.075 $Y=0.74 $X2=0
+ $Y2=0
cc_1025 N_A_1762_74#_M1018_g N_VGND_c_2075_n 0.00487769f $X=13.14 $Y=0.835 $X2=0
+ $Y2=0
cc_1026 N_A_1762_74#_c_1441_n N_VGND_c_2075_n 0.0210826f $X=9.09 $Y=0.515 $X2=0
+ $Y2=0
cc_1027 N_A_1762_74#_c_1441_n N_VGND_c_2079_n 0.0134766f $X=9.09 $Y=0.515 $X2=0
+ $Y2=0
cc_1028 N_A_1762_74#_c_1428_n N_VGND_c_2080_n 0.00405065f $X=11.015 $Y=0.865
+ $X2=0 $Y2=0
cc_1029 N_A_2556_112#_M1031_g N_VPWR_c_1671_n 0.00607507f $X=13.9 $Y=2.4 $X2=0
+ $Y2=0
cc_1030 N_A_2556_112#_c_1617_n N_VPWR_c_1671_n 0.00578125f $X=13.81 $Y=1.385
+ $X2=0 $Y2=0
cc_1031 N_A_2556_112#_c_1620_n N_VPWR_c_1671_n 0.030344f $X=13.17 $Y=2.16 $X2=0
+ $Y2=0
cc_1032 N_A_2556_112#_c_1621_n N_VPWR_c_1671_n 0.0122557f $X=13.62 $Y=1.385
+ $X2=0 $Y2=0
cc_1033 N_A_2556_112#_c_1620_n N_VPWR_c_1681_n 0.00775887f $X=13.17 $Y=2.16
+ $X2=0 $Y2=0
cc_1034 N_A_2556_112#_M1031_g N_VPWR_c_1682_n 0.00515235f $X=13.9 $Y=2.4 $X2=0
+ $Y2=0
cc_1035 N_A_2556_112#_M1031_g N_VPWR_c_1662_n 0.0097222f $X=13.9 $Y=2.4 $X2=0
+ $Y2=0
cc_1036 N_A_2556_112#_c_1620_n N_VPWR_c_1662_n 0.00855956f $X=13.17 $Y=2.16
+ $X2=0 $Y2=0
cc_1037 N_A_2556_112#_c_1620_n N_Q_N_c_2014_n 0.0552251f $X=13.17 $Y=2.16 $X2=0
+ $Y2=0
cc_1038 N_A_2556_112#_c_1619_n N_Q_N_c_2011_n 0.0197595f $X=13.13 $Y=1.55 $X2=0
+ $Y2=0
cc_1039 N_A_2556_112#_c_1620_n N_Q_N_c_2011_n 0.0106741f $X=13.17 $Y=2.16 $X2=0
+ $Y2=0
cc_1040 N_A_2556_112#_c_1619_n Q_N 0.0422235f $X=13.13 $Y=1.55 $X2=0 $Y2=0
cc_1041 N_A_2556_112#_M1031_g Q 0.0338237f $X=13.9 $Y=2.4 $X2=0 $Y2=0
cc_1042 N_A_2556_112#_c_1616_n Q 0.0188373f $X=13.905 $Y=1.22 $X2=0 $Y2=0
cc_1043 N_A_2556_112#_c_1618_n Q 0.0125549f $X=13.9 $Y=1.385 $X2=0 $Y2=0
cc_1044 N_A_2556_112#_c_1621_n Q 0.026211f $X=13.62 $Y=1.385 $X2=0 $Y2=0
cc_1045 N_A_2556_112#_c_1616_n N_VGND_c_2064_n 0.0113395f $X=13.905 $Y=1.22
+ $X2=0 $Y2=0
cc_1046 N_A_2556_112#_c_1617_n N_VGND_c_2064_n 0.00760746f $X=13.81 $Y=1.385
+ $X2=0 $Y2=0
cc_1047 N_A_2556_112#_c_1619_n N_VGND_c_2064_n 0.0189646f $X=13.13 $Y=1.55 $X2=0
+ $Y2=0
cc_1048 N_A_2556_112#_c_1621_n N_VGND_c_2064_n 0.0265928f $X=13.62 $Y=1.385
+ $X2=0 $Y2=0
cc_1049 N_A_2556_112#_c_1619_n N_VGND_c_2073_n 0.0099752f $X=13.13 $Y=1.55 $X2=0
+ $Y2=0
cc_1050 N_A_2556_112#_c_1616_n N_VGND_c_2074_n 0.00434272f $X=13.905 $Y=1.22
+ $X2=0 $Y2=0
cc_1051 N_A_2556_112#_c_1616_n N_VGND_c_2075_n 0.00828717f $X=13.905 $Y=1.22
+ $X2=0 $Y2=0
cc_1052 N_A_2556_112#_c_1619_n N_VGND_c_2075_n 0.0132953f $X=13.13 $Y=1.55 $X2=0
+ $Y2=0
cc_1053 N_VPWR_c_1663_n N_A_293_464#_c_1830_n 0.0100033f $X=0.73 $Y=2.805 $X2=0
+ $Y2=0
cc_1054 N_VPWR_c_1679_n N_A_293_464#_c_1830_n 0.0173809f $X=2.555 $Y=3.33 $X2=0
+ $Y2=0
cc_1055 N_VPWR_c_1662_n N_A_293_464#_c_1830_n 0.0178497f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1056 N_VPWR_c_1679_n N_A_293_464#_c_1845_n 0.00875362f $X=2.555 $Y=3.33 $X2=0
+ $Y2=0
cc_1057 N_VPWR_c_1662_n N_A_293_464#_c_1845_n 0.0129168f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1058 N_VPWR_M1013_d N_A_293_464#_c_1825_n 0.00616563f $X=2.515 $Y=2.32 $X2=0
+ $Y2=0
cc_1059 N_VPWR_c_1664_n N_A_293_464#_c_1825_n 0.0196553f $X=2.655 $Y=2.825 $X2=0
+ $Y2=0
cc_1060 N_VPWR_c_1666_n N_A_293_464#_c_1825_n 0.0021187f $X=3.74 $Y=2.78 $X2=0
+ $Y2=0
cc_1061 N_VPWR_c_1662_n N_A_293_464#_c_1825_n 0.0310339f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1062 N_VPWR_M1026_d N_A_293_464#_c_1826_n 9.89723e-19 $X=3.605 $Y=1.84 $X2=0
+ $Y2=0
cc_1063 N_VPWR_c_1666_n N_A_293_464#_c_1826_n 0.00274559f $X=3.74 $Y=2.78 $X2=0
+ $Y2=0
cc_1064 N_VPWR_M1026_d N_A_293_464#_c_1914_n 0.00462404f $X=3.605 $Y=1.84 $X2=0
+ $Y2=0
cc_1065 N_VPWR_c_1666_n N_A_293_464#_c_1914_n 0.0109162f $X=3.74 $Y=2.78 $X2=0
+ $Y2=0
cc_1066 N_VPWR_c_1662_n N_A_293_464#_c_1914_n 5.62582e-19 $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1067 N_VPWR_c_1662_n N_A_1603_347#_c_1946_n 0.0094792f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1068 N_VPWR_c_1668_n N_A_1603_347#_c_1947_n 0.0157924f $X=7.7 $Y=2.525 $X2=0
+ $Y2=0
cc_1069 N_VPWR_c_1676_n N_A_1603_347#_c_1947_n 0.00727677f $X=10.58 $Y=3.33
+ $X2=0 $Y2=0
cc_1070 N_VPWR_c_1662_n N_A_1603_347#_c_1947_n 0.00889546f $X=14.16 $Y=3.33
+ $X2=0 $Y2=0
cc_1071 N_VPWR_c_1669_n N_A_1712_374#_c_1980_n 0.0101219f $X=10.665 $Y=2.75
+ $X2=0 $Y2=0
cc_1072 N_VPWR_c_1676_n N_A_1712_374#_c_1980_n 0.0992665f $X=10.58 $Y=3.33 $X2=0
+ $Y2=0
cc_1073 N_VPWR_c_1662_n N_A_1712_374#_c_1980_n 0.054558f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1074 N_VPWR_c_1669_n N_A_1712_374#_c_1981_n 0.0132886f $X=10.665 $Y=2.75
+ $X2=0 $Y2=0
cc_1075 N_VPWR_c_1676_n N_A_1712_374#_c_1982_n 0.0214714f $X=10.58 $Y=3.33 $X2=0
+ $Y2=0
cc_1076 N_VPWR_c_1662_n N_A_1712_374#_c_1982_n 0.0110721f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1077 N_VPWR_c_1670_n N_Q_N_c_2015_n 0.0173821f $X=12.115 $Y=2.75 $X2=0 $Y2=0
cc_1078 N_VPWR_c_1681_n N_Q_N_c_2015_n 0.0111875f $X=13.455 $Y=3.33 $X2=0 $Y2=0
cc_1079 N_VPWR_c_1662_n N_Q_N_c_2015_n 0.00918014f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1080 N_VPWR_c_1671_n Q 0.0378352f $X=13.62 $Y=2.16 $X2=0 $Y2=0
cc_1081 N_VPWR_c_1682_n Q 0.0147571f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1082 N_VPWR_c_1662_n Q 0.0121348f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1083 N_A_293_464#_c_1845_n A_419_464# 0.00431352f $X=2.215 $Y=2.715 $X2=-0.19
+ $Y2=-0.245
cc_1084 N_A_293_464#_c_1850_n A_419_464# 0.00155419f $X=2.3 $Y=2.63 $X2=-0.19
+ $Y2=-0.245
cc_1085 N_A_293_464#_c_1854_n A_419_464# 0.00159805f $X=2.3 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_1086 N_A_293_464#_c_1818_n N_VGND_c_2059_n 0.00639088f $X=1.67 $Y=0.58 $X2=0
+ $Y2=0
cc_1087 N_A_293_464#_c_1818_n N_VGND_c_2060_n 0.0126723f $X=1.67 $Y=0.58 $X2=0
+ $Y2=0
cc_1088 N_A_293_464#_c_1819_n N_VGND_c_2060_n 0.00351301f $X=2.215 $Y=1.005
+ $X2=0 $Y2=0
cc_1089 N_A_293_464#_c_1818_n N_VGND_c_2065_n 0.0144922f $X=1.67 $Y=0.58 $X2=0
+ $Y2=0
cc_1090 N_A_293_464#_c_1818_n N_VGND_c_2075_n 0.0118826f $X=1.67 $Y=0.58 $X2=0
+ $Y2=0
cc_1091 N_A_1603_347#_c_1946_n N_A_1712_374#_M1033_s 0.00379272f $X=9.58
+ $Y=2.435 $X2=-0.19 $Y2=1.66
cc_1092 N_A_1603_347#_c_1946_n N_A_1712_374#_c_1980_n 0.0234493f $X=9.58
+ $Y=2.435 $X2=0 $Y2=0
cc_1093 N_A_1603_347#_c_1948_n N_A_1712_374#_c_1980_n 0.0184181f $X=9.665
+ $Y=2.51 $X2=0 $Y2=0
cc_1094 N_A_1603_347#_c_1948_n N_A_1712_374#_c_1981_n 0.0146403f $X=9.665
+ $Y=2.51 $X2=0 $Y2=0
cc_1095 N_A_1603_347#_c_1946_n N_A_1712_374#_c_1982_n 0.0253437f $X=9.58
+ $Y=2.435 $X2=0 $Y2=0
cc_1096 N_A_1603_347#_c_1947_n N_A_1712_374#_c_1982_n 0.00459189f $X=8.15
+ $Y=2.435 $X2=0 $Y2=0
cc_1097 Q_N N_VGND_c_2063_n 0.0326809f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1098 Q_N N_VGND_c_2073_n 0.0219264f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1099 Q_N N_VGND_c_2075_n 0.0180924f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_1100 Q N_VGND_c_2064_n 0.0271167f $X=14.075 $Y=0.47 $X2=0 $Y2=0
cc_1101 Q N_VGND_c_2074_n 0.014787f $X=14.075 $Y=0.47 $X2=0 $Y2=0
cc_1102 Q N_VGND_c_2075_n 0.012183f $X=14.075 $Y=0.47 $X2=0 $Y2=0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and4b_4 A_N B C D VGND VNB VPB VPWR X
X0 VPWR B a_199_294# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X1 VPWR D a_199_294# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X2 a_199_294# a_27_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X3 a_751_125# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 VPWR C a_199_294# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X5 a_199_294# D VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X6 a_199_294# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X7 VGND a_199_294# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 VGND a_199_294# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_664_125# C a_751_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X10 VPWR a_199_294# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X11 X a_199_294# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X12 a_1136_125# a_27_368# a_199_294# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 a_199_294# a_27_368# a_1136_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X14 a_1136_125# B a_664_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 a_27_368# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X16 a_27_368# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X17 X a_199_294# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 VPWR a_27_368# a_199_294# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X19 a_199_294# C VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X20 a_664_125# B a_1136_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X21 a_751_125# C a_664_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X22 VGND D a_751_125# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X23 VPWR a_199_294# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X24 X a_199_294# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 X a_199_294# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
.ends

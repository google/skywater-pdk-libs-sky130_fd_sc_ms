* File: sky130_fd_sc_ms__xnor3_4.spice
* Created: Fri Aug 28 18:18:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__xnor3_4.pex.spice"
.subckt sky130_fd_sc_ms__xnor3_4  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1016 N_VGND_M1016_d N_A_75_227#_M1016_g N_A_27_373#_M1016_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.112 AS=0.1824 PD=0.99 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1003 N_A_75_227#_M1003_d N_A_M1003_g N_VGND_M1016_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1072 AS=0.112 PD=0.975 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.7
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1024 N_A_321_77#_M1024_d N_B_M1024_g N_A_75_227#_M1003_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.115623 AS=0.1072 PD=1.16528 PS=0.975 NRD=8.436 NRS=10.308 M=1
+ R=4.26667 SA=75001.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1006 N_A_27_373#_M1006_d N_A_386_23#_M1006_g N_A_321_77#_M1024_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.111379 AS=0.0758774 PD=0.87566 PS=0.764717 NRD=60.048 NRS=0
+ M=1 R=2.8 SA=75001.7 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1005 N_A_327_373#_M1005_d N_B_M1005_g N_A_27_373#_M1006_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.096 AS=0.169721 PD=0.94 PS=1.33434 NRD=1.872 NRS=19.68 M=1
+ R=4.26667 SA=75001.6 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1009 N_A_75_227#_M1009_d N_A_386_23#_M1009_g N_A_327_373#_M1005_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.3467 AS=0.096 PD=2.79 PS=0.94 NRD=91.248 NRS=1.872 M=1
+ R=4.26667 SA=75002.1 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1022 N_VGND_M1022_d N_B_M1022_g N_A_386_23#_M1022_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.3368 AS=0.2109 PD=2.67 PS=2.05 NRD=64.884 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1027 N_A_1057_74#_M1027_d N_A_1024_300#_M1027_g N_A_321_77#_M1027_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1296 AS=0.1824 PD=1.045 PS=1.85 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1010 N_A_327_373#_M1010_d N_C_M1010_g N_A_1057_74#_M1027_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.192 AS=0.1296 PD=1.88 PS=1.045 NRD=2.808 NRS=10.308 M=1 R=4.26667
+ SA=75000.8 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1017 N_VGND_M1017_d N_C_M1017_g N_A_1024_300#_M1017_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.497211 AS=0.1197 PD=1.75603 PS=1.41 NRD=312.852 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_1057_74#_M1001_g N_VGND_M1017_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.876039 PD=1.02 PS=3.09397 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1004 N_X_M1001_d N_A_1057_74#_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1011 N_X_M1011_d N_A_1057_74#_M1011_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.4
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1013 N_X_M1011_d N_A_1057_74#_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1020 N_VPWR_M1020_d N_A_75_227#_M1020_g N_A_27_373#_M1020_s VPB PSHORT L=0.18
+ W=1 AD=0.16 AS=0.28 PD=1.32 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90002.3 A=0.18 P=2.36 MULT=1
MM1018 N_A_75_227#_M1018_d N_A_M1018_g N_VPWR_M1020_d VPB PSHORT L=0.18 W=1
+ AD=0.188696 AS=0.16 PD=1.47826 PS=1.32 NRD=0 NRS=8.8453 M=1 R=5.55556
+ SA=90000.7 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1025 N_A_327_373#_M1025_d N_B_M1025_g N_A_75_227#_M1018_d VPB PSHORT L=0.18
+ W=0.84 AD=0.217265 AS=0.158504 PD=1.54378 PS=1.24174 NRD=57.4452 NRS=20.3107
+ M=1 R=4.66667 SA=90001.2 SB=90001.5 A=0.1512 P=2.04 MULT=1
MM1014 N_A_27_373#_M1014_d N_A_386_23#_M1014_g N_A_327_373#_M1025_d VPB PSHORT
+ L=0.18 W=0.64 AD=0.0864 AS=0.165535 PD=0.91 PS=1.17622 NRD=0 NRS=0 M=1
+ R=3.55556 SA=90001.9 SB=90001.2 A=0.1152 P=1.64 MULT=1
MM1015 N_A_321_77#_M1015_d N_B_M1015_g N_A_27_373#_M1014_d VPB PSHORT L=0.18
+ W=0.64 AD=0.112951 AS=0.0864 PD=1.01189 PS=0.91 NRD=16.9223 NRS=0 M=1
+ R=3.55556 SA=90002.4 SB=90000.8 A=0.1152 P=1.64 MULT=1
MM1000 N_A_75_227#_M1000_d N_A_386_23#_M1000_g N_A_321_77#_M1015_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.37475 AS=0.148249 PD=2.88 PS=1.32811 NRD=91.7232 NRS=0 M=1
+ R=4.66667 SA=90002.2 SB=90000.3 A=0.1512 P=2.04 MULT=1
MM1007 N_VPWR_M1007_d N_B_M1007_g N_A_386_23#_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.3136 PD=2.8 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1021 N_A_1057_74#_M1021_d N_A_1024_300#_M1021_g N_A_327_373#_M1021_s VPB
+ PSHORT L=0.18 W=0.84 AD=0.21525 AS=0.2352 PD=1.49 PS=2.24 NRD=47.1815 NRS=0
+ M=1 R=4.66667 SA=90000.2 SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1019 N_A_321_77#_M1019_d N_C_M1019_g N_A_1057_74#_M1021_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.21525 PD=2.24 PS=1.49 NRD=0 NRS=47.1815 M=1 R=4.66667
+ SA=90000.8 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1012 N_VPWR_M1012_d N_C_M1012_g N_A_1024_300#_M1012_s VPB PSHORT L=0.18 W=0.64
+ AD=0.377018 AS=0.1792 PD=1.55636 PS=1.84 NRD=160.062 NRS=0 M=1 R=3.55556
+ SA=90000.2 SB=90002.7 A=0.1152 P=1.64 MULT=1
MM1002 N_X_M1002_d N_A_1057_74#_M1002_g N_VPWR_M1012_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.659782 PD=1.39 PS=2.72364 NRD=0 NRS=18.8923 M=1 R=6.22222
+ SA=90001.1 SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1008 N_X_M1002_d N_A_1057_74#_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1023 N_X_M1023_d N_A_1057_74#_M1023_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1026 N_X_M1023_d N_A_1057_74#_M1026_g N_VPWR_M1026_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.4
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX28_noxref VNB VPB NWDIODE A=19.4556 P=24.64
c_98 VNB 0 1.89638e-19 $X=0 $Y=0
c_186 VPB 0 1.87651e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__xnor3_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__or2b_4.pex.spice
* Created: Fri Aug 28 18:07:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__OR2B_4%A_81_296# 1 2 3 12 16 22 26 30 34 38 42 44 45
+ 53 57 59 63 67 69 73 74 77 84
c139 42 0 1.88904e-19 $X=1.88 $Y=0.74
r140 83 84 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=1.845 $Y=1.465
+ $X2=1.88 $Y2=1.465
r141 80 81 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=1.395 $Y=1.465
+ $X2=1.425 $Y2=1.465
r142 76 78 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=0.925 $Y=1.465
+ $X2=0.945 $Y2=1.465
r143 76 77 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.925 $Y=1.465
+ $X2=0.85 $Y2=1.465
r144 74 75 18.9664 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.63 $Y=1.28 $X2=4
+ $Y2=1.28
r145 65 75 0.414291 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=4 $Y=1.45 $X2=4
+ $Y2=1.28
r146 65 67 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=4 $Y=1.45 $X2=4
+ $Y2=2.08
r147 61 74 0.414291 $w=2.5e-07 $l=1.7e-07 $layer=LI1_cond $X=3.63 $Y=1.11
+ $X2=3.63 $Y2=1.28
r148 61 63 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=3.63 $Y=1.11
+ $X2=3.63 $Y2=0.515
r149 60 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=1.195
+ $X2=2.64 $Y2=1.195
r150 59 74 7.42157 $w=2.38e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.505 $Y=1.195
+ $X2=3.63 $Y2=1.28
r151 59 60 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.505 $Y=1.195
+ $X2=2.805 $Y2=1.195
r152 55 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=1.11
+ $X2=2.64 $Y2=1.195
r153 55 57 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=2.64 $Y=1.11
+ $X2=2.64 $Y2=0.515
r154 54 69 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=1.195
+ $X2=2.06 $Y2=1.195
r155 53 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=1.195
+ $X2=2.64 $Y2=1.195
r156 53 54 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.475 $Y=1.195
+ $X2=2.145 $Y2=1.195
r157 52 83 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=1.79 $Y=1.465
+ $X2=1.845 $Y2=1.465
r158 52 81 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=1.79 $Y=1.465
+ $X2=1.425 $Y2=1.465
r159 51 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.79
+ $Y=1.465 $X2=1.79 $Y2=1.465
r160 48 80 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=1.11 $Y=1.465
+ $X2=1.395 $Y2=1.465
r161 48 78 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.11 $Y=1.465
+ $X2=0.945 $Y2=1.465
r162 47 51 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.11 $Y=1.465
+ $X2=1.79 $Y2=1.465
r163 47 48 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.11
+ $Y=1.465 $X2=1.11 $Y2=1.465
r164 45 69 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.06 $Y=1.465
+ $X2=2.06 $Y2=1.195
r165 45 51 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.975 $Y=1.465
+ $X2=1.79 $Y2=1.465
r166 40 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.88 $Y=1.3
+ $X2=1.88 $Y2=1.465
r167 40 42 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.88 $Y=1.3
+ $X2=1.88 $Y2=0.74
r168 36 83 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.63
+ $X2=1.845 $Y2=1.465
r169 36 38 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.845 $Y=1.63
+ $X2=1.845 $Y2=2.4
r170 32 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.3
+ $X2=1.425 $Y2=1.465
r171 32 34 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.425 $Y=1.3
+ $X2=1.425 $Y2=0.74
r172 28 80 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.395 $Y=1.63
+ $X2=1.395 $Y2=1.465
r173 28 30 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.395 $Y=1.63
+ $X2=1.395 $Y2=2.4
r174 24 78 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=1.63
+ $X2=0.945 $Y2=1.465
r175 24 26 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.945 $Y=1.63
+ $X2=0.945 $Y2=2.4
r176 20 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.3
+ $X2=0.925 $Y2=1.465
r177 20 22 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.925 $Y=1.3
+ $X2=0.925 $Y2=0.74
r178 19 44 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.585 $Y=1.555
+ $X2=0.495 $Y2=1.555
r179 19 77 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.585 $Y=1.555
+ $X2=0.85 $Y2=1.555
r180 14 44 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=1.48
+ $X2=0.495 $Y2=1.555
r181 14 16 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.495 $Y=1.48
+ $X2=0.495 $Y2=0.74
r182 10 44 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=1.63
+ $X2=0.495 $Y2=1.555
r183 10 12 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.495 $Y=1.63
+ $X2=0.495 $Y2=2.4
r184 3 67 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.905
+ $Y=1.935 $X2=4.04 $Y2=2.08
r185 2 63 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.53
+ $Y=0.37 $X2=3.67 $Y2=0.515
r186 1 57 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=2.43
+ $Y=0.37 $X2=2.64 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR2B_4%A 3 7 9 13 17 19 20 21 24
r59 27 29 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.615
+ $X2=2.865 $Y2=1.78
r60 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.865
+ $Y=1.615 $X2=2.865 $Y2=1.615
r61 24 27 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=2.865 $Y=1.515
+ $X2=2.865 $Y2=1.615
r62 24 25 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.865 $Y=1.515
+ $X2=2.865 $Y2=1.44
r63 21 28 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=3.12 $Y=1.615
+ $X2=2.865 $Y2=1.615
r64 20 28 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=2.64 $Y=1.615
+ $X2=2.865 $Y2=1.615
r65 17 25 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=2.955 $Y=0.69
+ $X2=2.955 $Y2=1.44
r66 13 29 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=2.82 $Y=2.46
+ $X2=2.82 $Y2=1.78
r67 10 19 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.46 $Y=1.515 $X2=2.37
+ $Y2=1.515
r68 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=1.515
+ $X2=2.865 $Y2=1.515
r69 9 10 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.7 $Y=1.515 $X2=2.46
+ $Y2=1.515
r70 5 19 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=2.37 $Y=1.59
+ $X2=2.37 $Y2=1.515
r71 5 7 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=2.37 $Y=1.59 $X2=2.37
+ $Y2=2.46
r72 1 19 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=2.355 $Y=1.44
+ $X2=2.37 $Y2=1.515
r73 1 3 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=2.355 $Y=1.44
+ $X2=2.355 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__OR2B_4%A_676_48# 1 2 9 11 12 15 19 25 27 28 30 36 41
+ 42 43 48
c87 25 0 7.62661e-20 $X=4.265 $Y=2.435
r88 47 48 33.0969 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.265 $Y=1.61
+ $X2=4.175 $Y2=1.61
r89 42 47 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=4.46 $Y=1.61
+ $X2=4.265 $Y2=1.61
r90 41 43 7.81899 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.46 $Y=1.61
+ $X2=4.46 $Y2=1.445
r91 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.46
+ $Y=1.61 $X2=4.46 $Y2=1.61
r92 36 38 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=5.53 $Y=2.105
+ $X2=5.53 $Y2=2.815
r93 34 36 53.2429 $w=2.48e-07 $l=1.155e-06 $layer=LI1_cond $X=5.53 $Y=0.95
+ $X2=5.53 $Y2=2.105
r94 31 46 2.29372 $w=6e-07 $l=9.5e-08 $layer=LI1_cond $X=4.625 $Y=0.65 $X2=4.53
+ $Y2=0.65
r95 31 33 13.3562 $w=5.98e-07 $l=6.7e-07 $layer=LI1_cond $X=4.625 $Y=0.65
+ $X2=5.295 $Y2=0.65
r96 30 34 8.44061 $w=6e-07 $l=3.57071e-07 $layer=LI1_cond $X=5.405 $Y=0.65
+ $X2=5.53 $Y2=0.95
r97 30 33 2.19281 $w=5.98e-07 $l=1.1e-07 $layer=LI1_cond $X=5.405 $Y=0.65
+ $X2=5.295 $Y2=0.65
r98 28 46 7.24332 $w=1.9e-07 $l=3e-07 $layer=LI1_cond $X=4.53 $Y=0.95 $X2=4.53
+ $Y2=0.65
r99 28 43 28.8947 $w=1.88e-07 $l=4.95e-07 $layer=LI1_cond $X=4.53 $Y=0.95
+ $X2=4.53 $Y2=1.445
r100 23 47 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=1.775
+ $X2=4.265 $Y2=1.61
r101 23 25 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=4.265 $Y=1.775
+ $X2=4.265 $Y2=2.435
r102 22 27 13.2179 $w=1.5e-07 $l=1.18e-07 $layer=POLY_cond $X=3.96 $Y=1.52
+ $X2=3.842 $Y2=1.52
r103 22 48 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=3.96 $Y=1.52
+ $X2=4.175 $Y2=1.52
r104 17 27 10.9219 $w=1.5e-07 $l=9.40744e-08 $layer=POLY_cond $X=3.885 $Y=1.445
+ $X2=3.842 $Y2=1.52
r105 17 19 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=3.885 $Y=1.445
+ $X2=3.885 $Y2=0.69
r106 13 27 10.9219 $w=1.8e-07 $l=8.74643e-08 $layer=POLY_cond $X=3.815 $Y=1.595
+ $X2=3.842 $Y2=1.52
r107 13 15 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=3.815 $Y=1.595
+ $X2=3.815 $Y2=2.435
r108 11 27 13.2179 $w=1.5e-07 $l=1.17e-07 $layer=POLY_cond $X=3.725 $Y=1.52
+ $X2=3.842 $Y2=1.52
r109 11 12 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=3.725 $Y=1.52
+ $X2=3.53 $Y2=1.52
r110 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.455 $Y=1.445
+ $X2=3.53 $Y2=1.52
r111 7 9 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=3.455 $Y=1.445
+ $X2=3.455 $Y2=0.69
r112 2 38 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.355
+ $Y=1.96 $X2=5.49 $Y2=2.815
r113 2 36 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.355
+ $Y=1.96 $X2=5.49 $Y2=2.105
r114 1 46 60.6667 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=3 $X=4.46
+ $Y=0.37 $X2=4.6 $Y2=0.515
r115 1 33 60.6667 $w=1.7e-07 $l=9.04599e-07 $layer=licon1_NDIFF $count=3 $X=4.46
+ $Y=0.37 $X2=5.295 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR2B_4%B_N 1 3 4 5 6 8 10 11 12 16
c36 11 0 7.62661e-20 $X=5.04 $Y=1.295
r37 11 12 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=5.07 $Y=1.285
+ $X2=5.07 $Y2=1.665
r38 11 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.07
+ $Y=1.285 $X2=5.07 $Y2=1.285
r39 10 16 39.0632 $w=4.2e-07 $l=2.95e-07 $layer=POLY_cond $X=5.115 $Y=1.58
+ $X2=5.115 $Y2=1.285
r40 9 16 6.62088 $w=4.2e-07 $l=5e-08 $layer=POLY_cond $X=5.115 $Y=1.235
+ $X2=5.115 $Y2=1.285
r41 6 10 41.5517 $w=3.48e-07 $l=3.67423e-07 $layer=POLY_cond $X=5.265 $Y=1.88
+ $X2=5.115 $Y2=1.58
r42 6 8 155.311 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=5.265 $Y=1.88
+ $X2=5.265 $Y2=2.46
r43 4 9 35.6662 $w=1.5e-07 $l=2.44643e-07 $layer=POLY_cond $X=4.905 $Y=1.16
+ $X2=5.115 $Y2=1.235
r44 4 5 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.905 $Y=1.16
+ $X2=4.46 $Y2=1.16
r45 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.385 $Y=1.085
+ $X2=4.46 $Y2=1.16
r46 1 3 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.385 $Y=1.085
+ $X2=4.385 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__OR2B_4%VPWR 1 2 3 4 5 16 18 24 28 34 38 43 44 46 47
+ 48 57 61 71 72 78 81
r78 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r79 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r80 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r81 72 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r82 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r83 69 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.205 $Y=3.33
+ $X2=5.04 $Y2=3.33
r84 69 71 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.205 $Y=3.33
+ $X2=5.52 $Y2=3.33
r85 68 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r86 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r87 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r88 65 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r89 64 67 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r90 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r91 62 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.21 $Y=3.33
+ $X2=3.085 $Y2=3.33
r92 62 64 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.21 $Y=3.33 $X2=3.6
+ $Y2=3.33
r93 61 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.875 $Y=3.33
+ $X2=5.04 $Y2=3.33
r94 61 67 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.875 $Y=3.33
+ $X2=4.56 $Y2=3.33
r95 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r96 57 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.96 $Y=3.33
+ $X2=3.085 $Y2=3.33
r97 57 59 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.96 $Y=3.33 $X2=2.64
+ $Y2=3.33
r98 56 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r99 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r100 53 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r101 53 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r102 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r103 50 75 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.217 $Y2=3.33
r104 50 52 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.72 $Y2=3.33
r105 48 79 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r106 48 60 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r107 46 55 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=1.68 $Y2=3.33
r108 46 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=2.11 $Y2=3.33
r109 45 59 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.235 $Y=3.33
+ $X2=2.64 $Y2=3.33
r110 45 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.235 $Y=3.33
+ $X2=2.11 $Y2=3.33
r111 43 52 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.72 $Y2=3.33
r112 43 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.13 $Y2=3.33
r113 42 55 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.255 $Y=3.33
+ $X2=1.68 $Y2=3.33
r114 42 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.255 $Y=3.33
+ $X2=1.13 $Y2=3.33
r115 38 41 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=5.04 $Y=2.125
+ $X2=5.04 $Y2=2.815
r116 36 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.04 $Y=3.245
+ $X2=5.04 $Y2=3.33
r117 36 41 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.04 $Y=3.245
+ $X2=5.04 $Y2=2.815
r118 32 78 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=3.245
+ $X2=3.085 $Y2=3.33
r119 32 34 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=3.085 $Y=3.245
+ $X2=3.085 $Y2=2.455
r120 28 31 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=2.11 $Y=2.105
+ $X2=2.11 $Y2=2.815
r121 26 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=3.245
+ $X2=2.11 $Y2=3.33
r122 26 31 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.11 $Y=3.245
+ $X2=2.11 $Y2=2.815
r123 22 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=3.245
+ $X2=1.13 $Y2=3.33
r124 22 24 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=1.13 $Y=3.245
+ $X2=1.13 $Y2=2.305
r125 18 21 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.27 $Y=1.985
+ $X2=0.27 $Y2=2.815
r126 16 75 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.217 $Y2=3.33
r127 16 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.27 $Y2=2.815
r128 5 41 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=4.9
+ $Y=1.96 $X2=5.04 $Y2=2.815
r129 5 38 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=4.9
+ $Y=1.96 $X2=5.04 $Y2=2.125
r130 4 34 300 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=2 $X=2.91
+ $Y=1.96 $X2=3.045 $Y2=2.455
r131 3 31 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=1.84 $X2=2.07 $Y2=2.815
r132 3 28 400 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=1.84 $X2=2.07 $Y2=2.105
r133 2 24 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=1.035
+ $Y=1.84 $X2=1.17 $Y2=2.305
r134 1 21 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.815
r135 1 18 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__OR2B_4%X 1 2 3 4 15 17 18 21 25 27 31 37 41 42 43
c69 25 0 1.88904e-19 $X=1.475 $Y=1.045
r70 41 43 15.2824 $w=2.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=1.295
+ $X2=0.24 $Y2=1.295
r71 40 41 0.898652 $w=2.3e-07 $l=1.25e-07 $layer=LI1_cond $X=0.67 $Y=1.295
+ $X2=0.545 $Y2=1.295
r72 39 40 12.8692 $w=2.37e-07 $l=2.5e-07 $layer=LI1_cond $X=0.67 $Y=1.045
+ $X2=0.67 $Y2=1.295
r73 35 37 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=1.64 $Y=0.96
+ $X2=1.64 $Y2=0.515
r74 31 33 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.62 $Y=1.985
+ $X2=1.62 $Y2=2.815
r75 29 31 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.62 $Y=1.97
+ $X2=1.62 $Y2=1.985
r76 28 42 1.64875 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.805 $Y=1.885
+ $X2=0.705 $Y2=1.885
r77 27 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.455 $Y=1.885
+ $X2=1.62 $Y2=1.97
r78 27 28 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.455 $Y=1.885
+ $X2=0.805 $Y2=1.885
r79 26 39 2.684 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=1.045
+ $X2=0.67 $Y2=1.045
r80 25 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.475 $Y=1.045
+ $X2=1.64 $Y2=0.96
r81 25 26 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.475 $Y=1.045
+ $X2=0.795 $Y2=1.045
r82 21 23 46.0273 $w=1.98e-07 $l=8.3e-07 $layer=LI1_cond $X=0.705 $Y=1.985
+ $X2=0.705 $Y2=2.815
r83 19 42 4.81226 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=1.97
+ $X2=0.705 $Y2=1.885
r84 19 21 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=0.705 $Y=1.97
+ $X2=0.705 $Y2=1.985
r85 18 42 4.81226 $w=1.85e-07 $l=9.21954e-08 $layer=LI1_cond $X=0.69 $Y=1.8
+ $X2=0.705 $Y2=1.885
r86 17 40 6.91381 $w=2.37e-07 $l=1.24599e-07 $layer=LI1_cond $X=0.69 $Y=1.41
+ $X2=0.67 $Y2=1.295
r87 17 18 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.69 $Y=1.41
+ $X2=0.69 $Y2=1.8
r88 13 39 4.19367 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.96 $X2=0.67
+ $Y2=1.045
r89 13 15 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.67 $Y=0.96
+ $X2=0.67 $Y2=0.515
r90 4 33 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.84 $X2=1.62 $Y2=2.815
r91 4 31 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.84 $X2=1.62 $Y2=1.985
r92 3 23 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.72 $Y2=2.815
r93 3 21 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.72 $Y2=1.985
r94 2 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.5
+ $Y=0.37 $X2=1.64 $Y2=0.515
r95 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR2B_4%A_492_392# 1 2 3 10 12 14 16 19 20 21 24
r54 24 27 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.49 $Y=2.11
+ $X2=4.49 $Y2=2.79
r55 22 27 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=4.49 $Y=2.905
+ $X2=4.49 $Y2=2.79
r56 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.325 $Y=2.99
+ $X2=4.49 $Y2=2.905
r57 20 21 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.325 $Y=2.99
+ $X2=3.675 $Y2=2.99
r58 17 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.55 $Y=2.905
+ $X2=3.675 $Y2=2.99
r59 17 19 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=3.55 $Y=2.905
+ $X2=3.55 $Y2=2.79
r60 16 31 2.99084 $w=2.5e-07 $l=1.03e-07 $layer=LI1_cond $X=3.55 $Y=2.12
+ $X2=3.55 $Y2=2.017
r61 16 19 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=3.55 $Y=2.12
+ $X2=3.55 $Y2=2.79
r62 15 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.76 $Y=2.035
+ $X2=2.595 $Y2=2.035
r63 14 31 4.15233 $w=1.7e-07 $l=1.33697e-07 $layer=LI1_cond $X=3.425 $Y=2.035
+ $X2=3.55 $Y2=2.017
r64 14 15 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.425 $Y=2.035
+ $X2=2.76 $Y2=2.035
r65 10 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=2.12
+ $X2=2.595 $Y2=2.035
r66 10 12 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.595 $Y=2.12
+ $X2=2.595 $Y2=2.815
r67 3 27 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.355
+ $Y=1.935 $X2=4.49 $Y2=2.79
r68 3 24 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=4.355
+ $Y=1.935 $X2=4.49 $Y2=2.11
r69 2 31 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.45
+ $Y=1.935 $X2=3.59 $Y2=2.08
r70 2 19 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.45
+ $Y=1.935 $X2=3.59 $Y2=2.79
r71 1 29 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=2.46
+ $Y=1.96 $X2=2.595 $Y2=2.115
r72 1 12 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.46
+ $Y=1.96 $X2=2.595 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__OR2B_4%VGND 1 2 3 4 5 16 18 22 26 30 34 36 38 43 48
+ 53 63 64 70 73 76 79
r78 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r79 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r80 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r81 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r82 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r83 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r84 61 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r85 61 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r86 60 63 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r87 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r88 58 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.265 $Y=0 $X2=4.1
+ $Y2=0
r89 58 60 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.265 $Y=0 $X2=4.56
+ $Y2=0
r90 57 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r91 57 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r92 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r93 54 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.335 $Y=0 $X2=3.17
+ $Y2=0
r94 54 56 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.335 $Y=0 $X2=3.6
+ $Y2=0
r95 53 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.935 $Y=0 $X2=4.1
+ $Y2=0
r96 53 56 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.935 $Y=0 $X2=3.6
+ $Y2=0
r97 52 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r98 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r99 49 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.14
+ $Y2=0
r100 49 51 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.305 $Y=0
+ $X2=2.64 $Y2=0
r101 48 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.005 $Y=0 $X2=3.17
+ $Y2=0
r102 48 51 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.005 $Y=0
+ $X2=2.64 $Y2=0
r103 47 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r104 47 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r105 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r106 44 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.14
+ $Y2=0
r107 44 46 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.305 $Y=0
+ $X2=1.68 $Y2=0
r108 43 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=2.14
+ $Y2=0
r109 43 46 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=1.68
+ $Y2=0
r110 42 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r111 42 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r112 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r113 39 67 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r114 39 41 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.72 $Y2=0
r115 38 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.14
+ $Y2=0
r116 38 41 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0
+ $X2=0.72 $Y2=0
r117 36 77 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=3.12 $Y2=0
r118 36 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=2.64 $Y2=0
r119 32 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.1 $Y=0.085 $X2=4.1
+ $Y2=0
r120 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.1 $Y=0.085
+ $X2=4.1 $Y2=0.515
r121 28 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.17 $Y=0.085
+ $X2=3.17 $Y2=0
r122 28 30 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.17 $Y=0.085
+ $X2=3.17 $Y2=0.515
r123 24 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0
r124 24 26 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0.515
r125 20 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0
r126 20 22 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0.6
r127 16 67 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r128 16 18 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.505
r129 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.96
+ $Y=0.37 $X2=4.1 $Y2=0.515
r130 4 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.03
+ $Y=0.37 $X2=3.17 $Y2=0.515
r131 3 26 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=1.955
+ $Y=0.37 $X2=2.14 $Y2=0.515
r132 2 22 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.37 $X2=1.14 $Y2=0.6
r133 1 18 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.505
.ends


* File: sky130_fd_sc_ms__einvp_1.pxi.spice
* Created: Wed Sep  2 12:08:39 2020
* 
x_PM_SKY130_FD_SC_MS__EINVP_1%A_44_549# N_A_44_549#_M1003_s N_A_44_549#_M1005_s
+ N_A_44_549#_c_48_n N_A_44_549#_c_49_n N_A_44_549#_M1000_g N_A_44_549#_c_45_n
+ N_A_44_549#_c_46_n N_A_44_549#_c_47_n N_A_44_549#_c_51_n N_A_44_549#_c_52_n
+ N_A_44_549#_c_53_n PM_SKY130_FD_SC_MS__EINVP_1%A_44_549#
x_PM_SKY130_FD_SC_MS__EINVP_1%TE N_TE_M1005_g N_TE_M1003_g N_TE_c_90_n
+ N_TE_M1001_g TE TE N_TE_c_93_n N_TE_c_94_n PM_SKY130_FD_SC_MS__EINVP_1%TE
x_PM_SKY130_FD_SC_MS__EINVP_1%A N_A_c_139_n N_A_M1004_g N_A_M1002_g N_A_c_136_n
+ A N_A_c_137_n N_A_c_138_n PM_SKY130_FD_SC_MS__EINVP_1%A
x_PM_SKY130_FD_SC_MS__EINVP_1%VPWR N_VPWR_M1005_d N_VPWR_c_163_n VPWR
+ N_VPWR_c_164_n N_VPWR_c_165_n N_VPWR_c_162_n N_VPWR_c_167_n
+ PM_SKY130_FD_SC_MS__EINVP_1%VPWR
x_PM_SKY130_FD_SC_MS__EINVP_1%Z N_Z_M1002_d N_Z_M1004_d N_Z_c_191_n N_Z_c_192_n
+ N_Z_c_204_n N_Z_c_193_n N_Z_c_195_n Z Z PM_SKY130_FD_SC_MS__EINVP_1%Z
x_PM_SKY130_FD_SC_MS__EINVP_1%VGND N_VGND_M1003_d N_VGND_c_226_n VGND
+ N_VGND_c_227_n N_VGND_c_228_n N_VGND_c_229_n N_VGND_c_230_n
+ PM_SKY130_FD_SC_MS__EINVP_1%VGND
cc_1 VNB N_A_44_549#_c_45_n 0.0311176f $X=-0.19 $Y=-0.245 $X2=0.19 $Y2=2.01
cc_2 VNB N_A_44_549#_c_46_n 0.0321729f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=0.735
cc_3 VNB N_A_44_549#_c_47_n 0.0209133f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.575
cc_4 VNB N_TE_M1003_g 0.0564205f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_5 VNB N_TE_c_90_n 0.0265752f $X=-0.19 $Y=-0.245 $X2=1.385 $Y2=3.11
cc_6 VNB N_TE_M1001_g 0.0293931f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.46
cc_7 VNB TE 0.00267865f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=0.735
cc_8 VNB N_TE_c_93_n 0.027005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_TE_c_94_n 0.0111472f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.965
cc_10 VNB N_A_M1002_g 0.0297146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_c_136_n 0.00216621f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=3.11
cc_12 VNB N_A_c_137_n 0.0560277f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.735
cc_13 VNB N_A_c_138_n 0.00385705f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.575
cc_14 VNB N_VPWR_c_162_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.497 $Y2=2.175
cc_15 VNB N_Z_c_191_n 0.0103948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_Z_c_192_n 0.0111859f $X=-0.19 $Y=-0.245 $X2=1.385 $Y2=3.11
cc_17 VNB N_Z_c_193_n 0.02581f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.46
cc_18 VNB N_VGND_c_226_n 0.0166561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_227_n 0.032472f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=2.46
cc_20 VNB N_VGND_c_228_n 0.0307665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_229_n 0.171006f $X=-0.19 $Y=-0.245 $X2=0.497 $Y2=2.175
cc_22 VNB N_VGND_c_230_n 0.00548191f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.91
cc_23 VPB N_A_44_549#_c_48_n 0.0459397f $X=-0.19 $Y=1.66 $X2=1.385 $Y2=3.11
cc_24 VPB N_A_44_549#_c_49_n 0.0150919f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=3.035
cc_25 VPB N_A_44_549#_c_45_n 0.0171975f $X=-0.19 $Y=1.66 $X2=0.19 $Y2=2.01
cc_26 VPB N_A_44_549#_c_51_n 0.0540047f $X=-0.19 $Y=1.66 $X2=0.715 $Y2=2.175
cc_27 VPB N_A_44_549#_c_52_n 0.0624106f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=2.91
cc_28 VPB N_A_44_549#_c_53_n 0.0291717f $X=-0.19 $Y=1.66 $X2=0.89 $Y2=2.965
cc_29 VPB N_TE_M1005_g 0.0286367f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_30 VPB TE 0.0108738f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=0.735
cc_31 VPB N_TE_c_93_n 0.019406f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB N_TE_c_94_n 0.00815262f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=2.965
cc_33 VPB N_A_c_139_n 0.0285966f $X=-0.19 $Y=1.66 $X2=0.33 $Y2=0.37
cc_34 VPB N_A_c_136_n 0.013048f $X=-0.19 $Y=1.66 $X2=0.89 $Y2=3.11
cc_35 VPB N_A_c_138_n 0.00716996f $X=-0.19 $Y=1.66 $X2=0.81 $Y2=0.575
cc_36 VPB N_VPWR_c_163_n 0.00683642f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_164_n 0.02821f $X=-0.19 $Y=1.66 $X2=1.475 $Y2=2.46
cc_38 VPB N_VPWR_c_165_n 0.0301422f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_162_n 0.0575286f $X=-0.19 $Y=1.66 $X2=0.497 $Y2=2.175
cc_40 VPB N_VPWR_c_167_n 0.00485691f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=2.91
cc_41 VPB N_Z_c_191_n 0.0063016f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_Z_c_195_n 0.0175065f $X=-0.19 $Y=1.66 $X2=0.81 $Y2=0.575
cc_43 VPB Z 0.0294608f $X=-0.19 $Y=1.66 $X2=0.715 $Y2=2.175
cc_44 N_A_44_549#_c_48_n N_TE_M1005_g 0.00141874f $X=1.385 $Y=3.11 $X2=0 $Y2=0
cc_45 N_A_44_549#_c_49_n N_TE_M1005_g 0.0120776f $X=1.475 $Y=3.035 $X2=0 $Y2=0
cc_46 N_A_44_549#_c_45_n N_TE_M1005_g 0.00496506f $X=0.19 $Y=2.01 $X2=0 $Y2=0
cc_47 N_A_44_549#_c_51_n N_TE_M1005_g 0.0104766f $X=0.715 $Y=2.175 $X2=0 $Y2=0
cc_48 N_A_44_549#_c_53_n N_TE_M1005_g 0.00228475f $X=0.89 $Y=2.965 $X2=0 $Y2=0
cc_49 N_A_44_549#_c_45_n N_TE_M1003_g 0.00771354f $X=0.19 $Y=2.01 $X2=0 $Y2=0
cc_50 N_A_44_549#_c_47_n N_TE_M1003_g 0.00711567f $X=0.81 $Y=0.575 $X2=0 $Y2=0
cc_51 N_A_44_549#_c_49_n N_TE_c_90_n 0.0130357f $X=1.475 $Y=3.035 $X2=0 $Y2=0
cc_52 N_A_44_549#_c_45_n TE 0.0270525f $X=0.19 $Y=2.01 $X2=0 $Y2=0
cc_53 N_A_44_549#_c_47_n TE 0.0228364f $X=0.81 $Y=0.575 $X2=0 $Y2=0
cc_54 N_A_44_549#_c_51_n TE 0.028084f $X=0.715 $Y=2.175 $X2=0 $Y2=0
cc_55 N_A_44_549#_c_45_n N_TE_c_93_n 0.00228985f $X=0.19 $Y=2.01 $X2=0 $Y2=0
cc_56 N_A_44_549#_c_47_n N_TE_c_93_n 0.0103428f $X=0.81 $Y=0.575 $X2=0 $Y2=0
cc_57 N_A_44_549#_c_51_n N_TE_c_93_n 0.00281856f $X=0.715 $Y=2.175 $X2=0 $Y2=0
cc_58 N_A_44_549#_c_49_n N_A_c_139_n 0.0633571f $X=1.475 $Y=3.035 $X2=-0.19
+ $Y2=-0.245
cc_59 N_A_44_549#_c_48_n N_VPWR_c_163_n 0.022096f $X=1.385 $Y=3.11 $X2=0 $Y2=0
cc_60 N_A_44_549#_c_49_n N_VPWR_c_163_n 0.0185739f $X=1.475 $Y=3.035 $X2=0 $Y2=0
cc_61 N_A_44_549#_c_51_n N_VPWR_c_163_n 0.0654877f $X=0.715 $Y=2.175 $X2=0 $Y2=0
cc_62 N_A_44_549#_c_53_n N_VPWR_c_163_n 0.00120066f $X=0.89 $Y=2.965 $X2=0 $Y2=0
cc_63 N_A_44_549#_c_51_n N_VPWR_c_164_n 0.0538165f $X=0.715 $Y=2.175 $X2=0 $Y2=0
cc_64 N_A_44_549#_c_52_n N_VPWR_c_164_n 0.0207159f $X=0.725 $Y=2.91 $X2=0 $Y2=0
cc_65 N_A_44_549#_c_48_n N_VPWR_c_165_n 0.00543892f $X=1.385 $Y=3.11 $X2=0 $Y2=0
cc_66 N_A_44_549#_c_48_n N_VPWR_c_162_n 0.0186893f $X=1.385 $Y=3.11 $X2=0 $Y2=0
cc_67 N_A_44_549#_c_51_n N_VPWR_c_162_n 0.0274069f $X=0.715 $Y=2.175 $X2=0 $Y2=0
cc_68 N_A_44_549#_c_52_n N_VPWR_c_162_n 0.011903f $X=0.725 $Y=2.91 $X2=0 $Y2=0
cc_69 N_A_44_549#_c_53_n N_VPWR_c_162_n 0.00526618f $X=0.89 $Y=2.965 $X2=0 $Y2=0
cc_70 N_A_44_549#_c_49_n N_Z_c_191_n 0.00287181f $X=1.475 $Y=3.035 $X2=0 $Y2=0
cc_71 N_A_44_549#_c_49_n N_Z_c_195_n 0.0014979f $X=1.475 $Y=3.035 $X2=0 $Y2=0
cc_72 N_A_44_549#_c_49_n Z 0.00199884f $X=1.475 $Y=3.035 $X2=0 $Y2=0
cc_73 N_A_44_549#_c_49_n N_VGND_c_226_n 5.3302e-19 $X=1.475 $Y=3.035 $X2=0 $Y2=0
cc_74 N_A_44_549#_c_47_n N_VGND_c_226_n 0.0212724f $X=0.81 $Y=0.575 $X2=0 $Y2=0
cc_75 N_A_44_549#_c_46_n N_VGND_c_227_n 0.00610681f $X=0.275 $Y=0.735 $X2=0
+ $Y2=0
cc_76 N_A_44_549#_c_47_n N_VGND_c_227_n 0.0222861f $X=0.81 $Y=0.575 $X2=0 $Y2=0
cc_77 N_A_44_549#_c_46_n N_VGND_c_229_n 0.00604639f $X=0.275 $Y=0.735 $X2=0
+ $Y2=0
cc_78 N_A_44_549#_c_47_n N_VGND_c_229_n 0.0235867f $X=0.81 $Y=0.575 $X2=0 $Y2=0
cc_79 N_TE_M1001_g N_A_M1002_g 0.0329902f $X=1.515 $Y=0.74 $X2=0 $Y2=0
cc_80 N_TE_c_90_n N_A_c_137_n 0.0329902f $X=1.44 $Y=1.515 $X2=0 $Y2=0
cc_81 N_TE_c_94_n N_A_c_137_n 0.00156384f $X=0.95 $Y=1.605 $X2=0 $Y2=0
cc_82 N_TE_M1005_g N_VPWR_c_163_n 0.00313349f $X=0.94 $Y=2.17 $X2=0 $Y2=0
cc_83 N_TE_c_90_n N_VPWR_c_163_n 0.002513f $X=1.44 $Y=1.515 $X2=0 $Y2=0
cc_84 TE N_VPWR_c_163_n 0.0154758f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_85 N_TE_c_94_n N_VPWR_c_163_n 2.09729e-19 $X=0.95 $Y=1.605 $X2=0 $Y2=0
cc_86 N_TE_M1005_g N_VPWR_c_162_n 0.00177544f $X=0.94 $Y=2.17 $X2=0 $Y2=0
cc_87 N_TE_M1005_g N_Z_c_191_n 0.00145277f $X=0.94 $Y=2.17 $X2=0 $Y2=0
cc_88 N_TE_M1001_g N_Z_c_191_n 0.0091827f $X=1.515 $Y=0.74 $X2=0 $Y2=0
cc_89 TE N_Z_c_191_n 0.0189581f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_90 N_TE_c_94_n N_Z_c_191_n 4.99808e-19 $X=0.95 $Y=1.605 $X2=0 $Y2=0
cc_91 N_TE_M1001_g N_Z_c_204_n 7.6545e-19 $X=1.515 $Y=0.74 $X2=0 $Y2=0
cc_92 N_TE_M1001_g N_Z_c_193_n 0.00176373f $X=1.515 $Y=0.74 $X2=0 $Y2=0
cc_93 N_TE_M1003_g N_VGND_c_226_n 0.0101098f $X=1.025 $Y=0.58 $X2=0 $Y2=0
cc_94 N_TE_c_90_n N_VGND_c_226_n 0.00356442f $X=1.44 $Y=1.515 $X2=0 $Y2=0
cc_95 N_TE_M1001_g N_VGND_c_226_n 0.00387195f $X=1.515 $Y=0.74 $X2=0 $Y2=0
cc_96 TE N_VGND_c_226_n 0.00967694f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_97 N_TE_M1003_g N_VGND_c_227_n 0.00461464f $X=1.025 $Y=0.58 $X2=0 $Y2=0
cc_98 N_TE_M1001_g N_VGND_c_228_n 0.00461464f $X=1.515 $Y=0.74 $X2=0 $Y2=0
cc_99 N_TE_M1003_g N_VGND_c_229_n 0.00913453f $X=1.025 $Y=0.58 $X2=0 $Y2=0
cc_100 N_TE_M1001_g N_VGND_c_229_n 0.00907828f $X=1.515 $Y=0.74 $X2=0 $Y2=0
cc_101 N_A_c_139_n N_VPWR_c_163_n 0.0027306f $X=1.895 $Y=1.92 $X2=0 $Y2=0
cc_102 N_A_c_139_n N_VPWR_c_165_n 0.005209f $X=1.895 $Y=1.92 $X2=0 $Y2=0
cc_103 N_A_c_139_n N_VPWR_c_162_n 0.00986922f $X=1.895 $Y=1.92 $X2=0 $Y2=0
cc_104 N_A_c_139_n N_Z_c_191_n 0.00290451f $X=1.895 $Y=1.92 $X2=0 $Y2=0
cc_105 N_A_M1002_g N_Z_c_191_n 0.0104807f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_106 N_A_c_138_n N_Z_c_191_n 0.0360328f $X=2.11 $Y=1.465 $X2=0 $Y2=0
cc_107 N_A_M1002_g N_Z_c_192_n 0.0151759f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_108 N_A_c_137_n N_Z_c_192_n 0.00232646f $X=2.11 $Y=1.465 $X2=0 $Y2=0
cc_109 N_A_c_138_n N_Z_c_192_n 0.0282627f $X=2.11 $Y=1.465 $X2=0 $Y2=0
cc_110 N_A_M1002_g N_Z_c_193_n 0.0123878f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_111 N_A_c_139_n N_Z_c_195_n 0.0224443f $X=1.895 $Y=1.92 $X2=0 $Y2=0
cc_112 N_A_c_137_n N_Z_c_195_n 0.00148544f $X=2.11 $Y=1.465 $X2=0 $Y2=0
cc_113 N_A_c_138_n N_Z_c_195_n 0.027873f $X=2.11 $Y=1.465 $X2=0 $Y2=0
cc_114 N_A_c_139_n Z 0.0138139f $X=1.895 $Y=1.92 $X2=0 $Y2=0
cc_115 N_A_M1002_g N_VGND_c_228_n 0.00434272f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A_M1002_g N_VGND_c_229_n 0.00824638f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_117 N_VPWR_c_163_n Z 0.0205004f $X=1.25 $Y=2.105 $X2=0 $Y2=0
cc_118 N_VPWR_c_165_n Z 0.0145873f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_119 N_VPWR_c_162_n Z 0.0119893f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_120 A_313_392# N_Z_c_195_n 0.00525124f $X=1.565 $Y=1.96 $X2=2.12 $Y2=2.115
cc_121 N_Z_c_204_n N_VGND_c_226_n 0.00156525f $X=1.775 $Y=1.045 $X2=0 $Y2=0
cc_122 N_Z_c_193_n N_VGND_c_226_n 0.00927251f $X=2.12 $Y=0.515 $X2=0 $Y2=0
cc_123 N_Z_c_193_n N_VGND_c_228_n 0.0145639f $X=2.12 $Y=0.515 $X2=0 $Y2=0
cc_124 N_Z_c_193_n N_VGND_c_229_n 0.0119984f $X=2.12 $Y=0.515 $X2=0 $Y2=0
cc_125 N_Z_c_204_n A_318_74# 0.00570883f $X=1.775 $Y=1.045 $X2=-0.19 $Y2=-0.245

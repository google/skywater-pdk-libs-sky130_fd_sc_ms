* File: sky130_fd_sc_ms__conb_1.spice
* Created: Wed Sep  2 12:02:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__conb_1.pex.spice"
.subckt sky130_fd_sc_ms__conb_1  VNB VPB HI VPWR VGND LO
* 
* LO	LO
* VGND	VGND
* VPWR	VPWR
* HI	HI
* VPB	VPB
* VNB	VNB
DX0_noxref VNB VPB NWDIODE A=3.3852 P=7.36
R0 N_HI_R0_pos N_VPWR_R0_neg SHORT 0.01 M=1
R1 N_VGND_R1_pos N_LO_R1_neg SHORT 0.01 M=1
*
.include "sky130_fd_sc_ms__conb_1.pxi.spice"
*
.ends
*
*

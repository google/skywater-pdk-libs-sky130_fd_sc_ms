* File: sky130_fd_sc_ms__dfrtp_1.pxi.spice
* Created: Wed Sep  2 12:03:03 2020
* 
x_PM_SKY130_FD_SC_MS__DFRTP_1%D N_D_c_232_n N_D_M1018_g N_D_M1026_g D D D
+ N_D_c_234_n N_D_c_235_n N_D_c_239_n PM_SKY130_FD_SC_MS__DFRTP_1%D
x_PM_SKY130_FD_SC_MS__DFRTP_1%CLK N_CLK_M1021_g N_CLK_M1023_g CLK N_CLK_c_265_n
+ N_CLK_c_266_n PM_SKY130_FD_SC_MS__DFRTP_1%CLK
x_PM_SKY130_FD_SC_MS__DFRTP_1%A_493_387# N_A_493_387#_M1001_d
+ N_A_493_387#_M1025_d N_A_493_387#_M1014_g N_A_493_387#_c_309_n
+ N_A_493_387#_c_310_n N_A_493_387#_M1002_g N_A_493_387#_c_312_n
+ N_A_493_387#_M1027_g N_A_493_387#_c_313_n N_A_493_387#_c_314_n
+ N_A_493_387#_M1010_g N_A_493_387#_c_315_n N_A_493_387#_c_316_n
+ N_A_493_387#_c_317_n N_A_493_387#_c_318_n N_A_493_387#_c_319_n
+ N_A_493_387#_c_338_p N_A_493_387#_c_320_n N_A_493_387#_c_321_n
+ N_A_493_387#_c_322_n N_A_493_387#_c_323_n N_A_493_387#_c_324_n
+ N_A_493_387#_c_325_n N_A_493_387#_c_326_n N_A_493_387#_c_327_n
+ N_A_493_387#_c_328_n N_A_493_387#_c_336_n
+ PM_SKY130_FD_SC_MS__DFRTP_1%A_493_387#
x_PM_SKY130_FD_SC_MS__DFRTP_1%A_833_400# N_A_833_400#_M1031_d
+ N_A_833_400#_M1029_d N_A_833_400#_c_506_n N_A_833_400#_M1008_g
+ N_A_833_400#_M1012_g N_A_833_400#_c_503_n N_A_833_400#_c_524_n
+ N_A_833_400#_c_527_n N_A_833_400#_c_510_n N_A_833_400#_c_504_n
+ N_A_833_400#_c_505_n PM_SKY130_FD_SC_MS__DFRTP_1%A_833_400#
x_PM_SKY130_FD_SC_MS__DFRTP_1%RESET_B N_RESET_B_M1009_g N_RESET_B_c_591_n
+ N_RESET_B_M1019_g N_RESET_B_c_592_n N_RESET_B_c_593_n N_RESET_B_M1006_g
+ N_RESET_B_c_602_n N_RESET_B_M1030_g N_RESET_B_c_595_n N_RESET_B_M1000_g
+ N_RESET_B_M1020_g N_RESET_B_c_597_n N_RESET_B_c_606_n N_RESET_B_c_607_n
+ N_RESET_B_c_608_n N_RESET_B_c_609_n N_RESET_B_c_610_n N_RESET_B_c_611_n
+ RESET_B N_RESET_B_c_598_n N_RESET_B_c_599_n N_RESET_B_c_613_n
+ N_RESET_B_c_614_n N_RESET_B_c_615_n PM_SKY130_FD_SC_MS__DFRTP_1%RESET_B
x_PM_SKY130_FD_SC_MS__DFRTP_1%A_701_463# N_A_701_463#_M1007_d
+ N_A_701_463#_M1014_d N_A_701_463#_M1030_d N_A_701_463#_M1031_g
+ N_A_701_463#_M1029_g N_A_701_463#_c_814_n N_A_701_463#_c_839_n
+ N_A_701_463#_c_805_n N_A_701_463#_c_806_n N_A_701_463#_c_807_n
+ N_A_701_463#_c_808_n N_A_701_463#_c_809_n N_A_701_463#_c_810_n
+ N_A_701_463#_c_817_n N_A_701_463#_c_811_n N_A_701_463#_c_819_n
+ N_A_701_463#_c_812_n PM_SKY130_FD_SC_MS__DFRTP_1%A_701_463#
x_PM_SKY130_FD_SC_MS__DFRTP_1%A_299_387# N_A_299_387#_M1023_s
+ N_A_299_387#_M1021_s N_A_299_387#_M1025_g N_A_299_387#_c_934_n
+ N_A_299_387#_M1001_g N_A_299_387#_c_946_n N_A_299_387#_c_947_n
+ N_A_299_387#_c_948_n N_A_299_387#_c_935_n N_A_299_387#_c_936_n
+ N_A_299_387#_M1007_g N_A_299_387#_M1022_g N_A_299_387#_c_951_n
+ N_A_299_387#_M1004_g N_A_299_387#_c_938_n N_A_299_387#_c_939_n
+ N_A_299_387#_M1016_g N_A_299_387#_c_955_n N_A_299_387#_c_941_n
+ N_A_299_387#_c_942_n N_A_299_387#_c_971_n N_A_299_387#_c_943_n
+ N_A_299_387#_c_944_n N_A_299_387#_c_958_n
+ PM_SKY130_FD_SC_MS__DFRTP_1%A_299_387#
x_PM_SKY130_FD_SC_MS__DFRTP_1%A_1518_203# N_A_1518_203#_M1017_d
+ N_A_1518_203#_M1020_d N_A_1518_203#_c_1119_n N_A_1518_203#_M1015_g
+ N_A_1518_203#_M1013_g N_A_1518_203#_c_1112_n N_A_1518_203#_c_1113_n
+ N_A_1518_203#_c_1114_n N_A_1518_203#_c_1122_n N_A_1518_203#_c_1123_n
+ N_A_1518_203#_c_1115_n N_A_1518_203#_c_1116_n N_A_1518_203#_c_1117_n
+ N_A_1518_203#_c_1125_n N_A_1518_203#_c_1126_n N_A_1518_203#_c_1118_n
+ PM_SKY130_FD_SC_MS__DFRTP_1%A_1518_203#
x_PM_SKY130_FD_SC_MS__DFRTP_1%A_1266_74# N_A_1266_74#_M1027_d
+ N_A_1266_74#_M1004_d N_A_1266_74#_M1017_g N_A_1266_74#_M1024_g
+ N_A_1266_74#_c_1226_n N_A_1266_74#_c_1227_n N_A_1266_74#_c_1228_n
+ N_A_1266_74#_M1011_g N_A_1266_74#_c_1229_n N_A_1266_74#_c_1230_n
+ N_A_1266_74#_c_1231_n N_A_1266_74#_M1028_g N_A_1266_74#_c_1232_n
+ N_A_1266_74#_c_1250_n N_A_1266_74#_c_1233_n N_A_1266_74#_c_1244_n
+ N_A_1266_74#_c_1234_n N_A_1266_74#_c_1267_n N_A_1266_74#_c_1363_p
+ N_A_1266_74#_c_1245_n N_A_1266_74#_c_1235_n N_A_1266_74#_c_1236_n
+ N_A_1266_74#_c_1237_n N_A_1266_74#_c_1238_n
+ PM_SKY130_FD_SC_MS__DFRTP_1%A_1266_74#
x_PM_SKY130_FD_SC_MS__DFRTP_1%A_1867_409# N_A_1867_409#_M1028_d
+ N_A_1867_409#_M1011_d N_A_1867_409#_c_1385_n N_A_1867_409#_M1005_g
+ N_A_1867_409#_M1003_g N_A_1867_409#_c_1381_n N_A_1867_409#_c_1382_n
+ N_A_1867_409#_c_1388_n N_A_1867_409#_c_1383_n N_A_1867_409#_c_1384_n
+ PM_SKY130_FD_SC_MS__DFRTP_1%A_1867_409#
x_PM_SKY130_FD_SC_MS__DFRTP_1%VPWR N_VPWR_M1018_s N_VPWR_M1019_d N_VPWR_M1021_d
+ N_VPWR_M1008_d N_VPWR_M1029_s N_VPWR_M1015_d N_VPWR_M1024_d N_VPWR_M1005_d
+ N_VPWR_c_1432_n N_VPWR_c_1433_n N_VPWR_c_1434_n N_VPWR_c_1435_n
+ N_VPWR_c_1436_n N_VPWR_c_1437_n N_VPWR_c_1438_n N_VPWR_c_1439_n
+ N_VPWR_c_1440_n N_VPWR_c_1441_n N_VPWR_c_1442_n N_VPWR_c_1443_n VPWR
+ N_VPWR_c_1444_n N_VPWR_c_1445_n N_VPWR_c_1446_n N_VPWR_c_1447_n
+ N_VPWR_c_1448_n N_VPWR_c_1449_n N_VPWR_c_1450_n N_VPWR_c_1451_n
+ N_VPWR_c_1452_n N_VPWR_c_1453_n N_VPWR_c_1454_n N_VPWR_c_1431_n
+ PM_SKY130_FD_SC_MS__DFRTP_1%VPWR
x_PM_SKY130_FD_SC_MS__DFRTP_1%A_30_78# N_A_30_78#_M1026_s N_A_30_78#_M1007_s
+ N_A_30_78#_M1018_d N_A_30_78#_M1014_s N_A_30_78#_c_1568_n N_A_30_78#_c_1574_n
+ N_A_30_78#_c_1569_n N_A_30_78#_c_1576_n N_A_30_78#_c_1570_n
+ N_A_30_78#_c_1577_n N_A_30_78#_c_1571_n N_A_30_78#_c_1572_n
+ N_A_30_78#_c_1579_n N_A_30_78#_c_1580_n N_A_30_78#_c_1573_n
+ PM_SKY130_FD_SC_MS__DFRTP_1%A_30_78#
x_PM_SKY130_FD_SC_MS__DFRTP_1%Q N_Q_M1003_s N_Q_M1005_s N_Q_c_1683_n
+ N_Q_c_1684_n Q Q Q N_Q_c_1685_n PM_SKY130_FD_SC_MS__DFRTP_1%Q
x_PM_SKY130_FD_SC_MS__DFRTP_1%VGND N_VGND_M1009_d N_VGND_M1023_d N_VGND_M1006_d
+ N_VGND_M1013_d N_VGND_M1028_s N_VGND_M1003_d N_VGND_c_1712_n N_VGND_c_1713_n
+ N_VGND_c_1714_n N_VGND_c_1715_n N_VGND_c_1716_n N_VGND_c_1717_n
+ N_VGND_c_1718_n N_VGND_c_1719_n VGND N_VGND_c_1720_n N_VGND_c_1721_n
+ N_VGND_c_1722_n N_VGND_c_1723_n N_VGND_c_1724_n N_VGND_c_1725_n
+ N_VGND_c_1726_n N_VGND_c_1727_n N_VGND_c_1728_n
+ PM_SKY130_FD_SC_MS__DFRTP_1%VGND
cc_1 VNB N_D_c_232_n 0.0406028f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.828
cc_2 VNB N_D_M1026_g 0.0286471f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_3 VNB N_D_c_234_n 0.0216279f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_4 VNB N_D_c_235_n 0.0281582f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_5 VNB CLK 0.00356247f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_6 VNB N_CLK_c_265_n 0.0265092f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB N_CLK_c_266_n 0.0166711f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_8 VNB N_A_493_387#_c_309_n 0.0102637f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_9 VNB N_A_493_387#_c_310_n 0.0246981f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_10 VNB N_A_493_387#_M1002_g 0.0243281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_493_387#_c_312_n 0.0192767f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.165
cc_12 VNB N_A_493_387#_c_313_n 0.0205614f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1
cc_13 VNB N_A_493_387#_c_314_n 0.0110769f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.845
cc_14 VNB N_A_493_387#_c_315_n 0.0081907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_493_387#_c_316_n 0.0369929f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.665
cc_16 VNB N_A_493_387#_c_317_n 0.0059887f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=2.035
cc_17 VNB N_A_493_387#_c_318_n 0.00293095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_493_387#_c_319_n 9.76188e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_493_387#_c_320_n 0.0169659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_493_387#_c_321_n 9.76919e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_493_387#_c_322_n 0.00385029f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_493_387#_c_323_n 0.0019226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_493_387#_c_324_n 0.00390484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_493_387#_c_325_n 0.0176845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_493_387#_c_326_n 0.0313598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_493_387#_c_327_n 0.00797767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_493_387#_c_328_n 0.00714349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_833_400#_M1012_g 0.0374366f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_29 VNB N_A_833_400#_c_503_n 0.00393175f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=1.165
cc_30 VNB N_A_833_400#_c_504_n 0.00275035f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.665
cc_31 VNB N_A_833_400#_c_505_n 0.00959482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_RESET_B_M1009_g 0.0204705f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.825
cc_33 VNB N_RESET_B_c_591_n 0.029225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_RESET_B_c_592_n 0.282729f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_35 VNB N_RESET_B_c_593_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_36 VNB N_RESET_B_M1006_g 0.0304415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_RESET_B_c_595_n 0.0270062f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.845
cc_38 VNB N_RESET_B_M1000_g 0.0510668f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=2.01
cc_39 VNB N_RESET_B_c_597_n 0.0144541f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=2.035
cc_40 VNB N_RESET_B_c_598_n 0.0349041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_RESET_B_c_599_n 0.00330649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_701_463#_M1031_g 0.0231233f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_43 VNB N_A_701_463#_c_805_n 0.00267896f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.295
cc_44 VNB N_A_701_463#_c_806_n 0.0027521f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.665
cc_45 VNB N_A_701_463#_c_807_n 0.00375429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_701_463#_c_808_n 0.0015235f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=2.035
cc_47 VNB N_A_701_463#_c_809_n 0.0418231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_701_463#_c_810_n 0.00322075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_701_463#_c_811_n 0.00336472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_701_463#_c_812_n 0.00442778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_299_387#_c_934_n 0.0140606f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_52 VNB N_A_299_387#_c_935_n 0.0365647f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_53 VNB N_A_299_387#_c_936_n 0.0619838f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.165
cc_54 VNB N_A_299_387#_M1007_g 0.0247999f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.845
cc_55 VNB N_A_299_387#_c_938_n 0.0226279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_299_387#_c_939_n 0.00146492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_299_387#_M1016_g 0.0517191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_299_387#_c_941_n 0.00905459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_299_387#_c_942_n 0.00910913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_299_387#_c_943_n 4.56385e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_299_387#_c_944_n 0.00289971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1518_203#_M1013_g 0.0207732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1518_203#_c_1112_n 0.0156636f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=1.165
cc_64 VNB N_A_1518_203#_c_1113_n 0.0155514f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_65 VNB N_A_1518_203#_c_1114_n 0.0105463f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=2.01
cc_66 VNB N_A_1518_203#_c_1115_n 0.0023345f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=1.665
cc_67 VNB N_A_1518_203#_c_1116_n 0.00392193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1518_203#_c_1117_n 0.0310153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1518_203#_c_1118_n 0.0124417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1266_74#_M1017_g 0.04091f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_71 VNB N_A_1266_74#_c_1226_n 0.0182931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1266_74#_c_1227_n 0.016718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1266_74#_c_1228_n 0.0126324f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.165
cc_74 VNB N_A_1266_74#_c_1229_n 0.0232568f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.845
cc_75 VNB N_A_1266_74#_c_1230_n 0.0100399f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=2.01
cc_76 VNB N_A_1266_74#_c_1231_n 0.0210614f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.165
cc_77 VNB N_A_1266_74#_c_1232_n 0.0123873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1266_74#_c_1233_n 0.00445288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1266_74#_c_1234_n 0.00403288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1266_74#_c_1235_n 0.00637997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1266_74#_c_1236_n 0.00599516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1266_74#_c_1237_n 0.00266453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1266_74#_c_1238_n 0.00109446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1867_409#_M1003_g 0.0383367f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_85 VNB N_A_1867_409#_c_1381_n 0.0564146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1867_409#_c_1382_n 0.0212821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1867_409#_c_1383_n 0.014962f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.845
cc_88 VNB N_A_1867_409#_c_1384_n 0.00445066f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=1.295
cc_89 VNB N_VPWR_c_1431_n 0.462217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_30_78#_c_1568_n 0.003401f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_91 VNB N_A_30_78#_c_1569_n 0.00542054f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1
cc_92 VNB N_A_30_78#_c_1570_n 0.00390068f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.165
cc_93 VNB N_A_30_78#_c_1571_n 0.00425886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_30_78#_c_1572_n 0.0223919f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=2.035
cc_95 VNB N_A_30_78#_c_1573_n 0.00551376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_Q_c_1683_n 0.00811762f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.6
cc_97 VNB N_Q_c_1684_n 0.00208381f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_98 VNB N_Q_c_1685_n 0.00535471f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.665
cc_99 VNB N_VGND_c_1712_n 0.0156373f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.845
cc_100 VNB N_VGND_c_1713_n 0.0140007f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.165
cc_101 VNB N_VGND_c_1714_n 0.0111809f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.665
cc_102 VNB N_VGND_c_1715_n 0.0145996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1716_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1717_n 0.0505973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1718_n 0.0297253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1719_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1720_n 0.0201695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1721_n 0.0744823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1722_n 0.0580863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1723_n 0.0325483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1724_n 0.0345892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1725_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1726_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1727_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1728_n 0.588959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VPB N_D_c_232_n 0.0142152f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.828
cc_117 VPB N_D_M1018_g 0.0623425f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.825
cc_118 VPB N_D_c_235_n 0.0248233f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_119 VPB N_D_c_239_n 0.0207718f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.845
cc_120 VPB N_CLK_M1021_g 0.0244552f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.01
cc_121 VPB CLK 0.00401162f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_122 VPB N_CLK_c_265_n 0.00555141f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_123 VPB N_A_493_387#_M1014_g 0.0280354f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_124 VPB N_A_493_387#_c_309_n 0.0113258f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_125 VPB N_A_493_387#_c_310_n 0.00567462f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_126 VPB N_A_493_387#_M1010_g 0.0245724f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=2.01
cc_127 VPB N_A_493_387#_c_322_n 0.00558147f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_493_387#_c_324_n 0.0070351f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_493_387#_c_328_n 0.0214675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_493_387#_c_336_n 0.0372848f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_833_400#_c_506_n 0.0402397f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1
cc_132 VPB N_A_833_400#_M1008_g 0.0225347f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_133 VPB N_A_833_400#_M1012_g 0.00203513f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_134 VPB N_A_833_400#_c_503_n 0.00130319f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.165
cc_135 VPB N_A_833_400#_c_510_n 0.00183167f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_833_400#_c_505_n 0.00377517f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_RESET_B_c_591_n 0.016789f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_RESET_B_M1019_g 0.0476635f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_139 VPB N_RESET_B_c_602_n 0.0722175f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.165
cc_140 VPB N_RESET_B_c_595_n 0.00254578f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.845
cc_141 VPB N_RESET_B_M1000_g 0.0151047f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=2.01
cc_142 VPB N_RESET_B_M1020_g 0.0252514f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_RESET_B_c_606_n 0.020403f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_RESET_B_c_607_n 0.00405114f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_RESET_B_c_608_n 0.0198788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_RESET_B_c_609_n 0.00168948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_RESET_B_c_610_n 0.00493802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_RESET_B_c_611_n 0.00335799f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_RESET_B_c_599_n 0.00152246f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_RESET_B_c_613_n 0.0303933f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_RESET_B_c_614_n 0.0318865f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_RESET_B_c_615_n 0.00620787f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_701_463#_M1029_g 0.0257157f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_701_463#_c_814_n 0.00250947f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_155 VPB N_A_701_463#_c_805_n 0.00374508f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.295
cc_156 VPB N_A_701_463#_c_809_n 0.0158423f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_701_463#_c_817_n 0.0020626f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_701_463#_c_811_n 0.00518095f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_701_463#_c_819_n 0.00350781f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_299_387#_M1025_g 0.0214025f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_161 VPB N_A_299_387#_c_946_n 0.0735552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_299_387#_c_947_n 0.0550828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_299_387#_c_948_n 0.0106469f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.165
cc_164 VPB N_A_299_387#_c_936_n 0.00654266f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.165
cc_165 VPB N_A_299_387#_M1022_g 0.0366772f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_299_387#_c_951_n 0.184481f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_299_387#_M1004_g 0.0249381f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_299_387#_c_938_n 0.0299618f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_299_387#_c_939_n 0.00685394f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_299_387#_c_955_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_299_387#_c_942_n 0.00389213f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_299_387#_c_943_n 9.98016e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_299_387#_c_958_n 0.00304845f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_1518_203#_c_1119_n 0.0069195f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.6
cc_175 VPB N_A_1518_203#_M1015_g 0.0455905f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_176 VPB N_A_1518_203#_c_1112_n 0.0041544f $X=-0.19 $Y=1.66 $X2=0.402
+ $Y2=1.165
cc_177 VPB N_A_1518_203#_c_1122_n 0.00691219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_1518_203#_c_1123_n 0.00198797f $X=-0.19 $Y=1.66 $X2=0.32
+ $Y2=1.295
cc_179 VPB N_A_1518_203#_c_1115_n 0.00168296f $X=-0.19 $Y=1.66 $X2=0.32
+ $Y2=1.665
cc_180 VPB N_A_1518_203#_c_1125_n 0.00902162f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_1518_203#_c_1126_n 0.00311963f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_1266_74#_M1024_g 0.0537663f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.95
cc_183 VPB N_A_1266_74#_c_1226_n 0.00533618f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_1266_74#_c_1227_n 0.003846f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_1266_74#_M1011_g 0.0339505f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.845
cc_186 VPB N_A_1266_74#_c_1232_n 9.60226e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_1266_74#_c_1244_n 0.00279595f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=2.035
cc_188 VPB N_A_1266_74#_c_1245_n 0.00553317f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_1266_74#_c_1235_n 0.00921317f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_1266_74#_c_1237_n 2.00274e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_1266_74#_c_1238_n 9.16426e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_1867_409#_c_1385_n 0.0283402f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1
cc_193 VPB N_A_1867_409#_c_1381_n 0.0304841f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_1867_409#_c_1382_n 0.00409062f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_1867_409#_c_1388_n 0.00987001f $X=-0.19 $Y=1.66 $X2=0.385
+ $Y2=1.165
cc_196 VPB N_A_1867_409#_c_1384_n 0.00279207f $X=-0.19 $Y=1.66 $X2=0.32
+ $Y2=1.295
cc_197 VPB N_VPWR_c_1432_n 0.0103331f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.165
cc_198 VPB N_VPWR_c_1433_n 0.0226189f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.295
cc_199 VPB N_VPWR_c_1434_n 0.00667138f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.845
cc_200 VPB N_VPWR_c_1435_n 0.00129922f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1436_n 0.0142067f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1437_n 0.0207312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1438_n 0.0233415f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1439_n 0.0190165f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1440_n 0.0204007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1441_n 0.0142652f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1442_n 0.0120013f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1443_n 0.0657363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1444_n 0.0166261f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1445_n 0.0173826f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1446_n 0.0563378f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1447_n 0.0543442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1448_n 0.0380491f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1449_n 0.00554228f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1450_n 0.00485433f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1451_n 0.00436844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1452_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1453_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1454_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1431_n 0.106488f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_30_78#_c_1574_n 0.00121614f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.165
cc_222 VPB N_A_30_78#_c_1569_n 0.00823629f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1
cc_223 VPB N_A_30_78#_c_1576_n 0.0162192f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.845
cc_224 VPB N_A_30_78#_c_1577_n 0.00148503f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.295
cc_225 VPB N_A_30_78#_c_1571_n 0.00480328f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_30_78#_c_1579_n 0.00475722f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_30_78#_c_1580_n 0.00637881f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB Q 0.0106512f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB Q 0.0224653f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_Q_c_1685_n 0.00312989f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.665
cc_231 N_D_M1026_g N_RESET_B_M1009_g 0.0245154f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_232 N_D_c_235_n N_RESET_B_M1009_g 9.92331e-19 $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_233 N_D_c_232_n N_RESET_B_c_591_n 0.0245154f $X=0.402 $Y=1.828 $X2=0 $Y2=0
cc_234 N_D_M1018_g N_RESET_B_M1019_g 0.0270074f $X=0.495 $Y=2.825 $X2=0 $Y2=0
cc_235 N_D_c_234_n N_RESET_B_c_598_n 0.0245154f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_236 N_D_c_239_n N_RESET_B_c_613_n 0.0245154f $X=0.385 $Y=1.845 $X2=0 $Y2=0
cc_237 N_D_M1018_g N_VPWR_c_1433_n 0.00385528f $X=0.495 $Y=2.825 $X2=0 $Y2=0
cc_238 N_D_c_235_n N_VPWR_c_1433_n 0.00974499f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_239 N_D_c_239_n N_VPWR_c_1433_n 6.71306e-19 $X=0.385 $Y=1.845 $X2=0 $Y2=0
cc_240 N_D_M1018_g N_VPWR_c_1434_n 5.02639e-19 $X=0.495 $Y=2.825 $X2=0 $Y2=0
cc_241 N_D_M1018_g N_VPWR_c_1444_n 0.00553346f $X=0.495 $Y=2.825 $X2=0 $Y2=0
cc_242 N_D_M1018_g N_VPWR_c_1431_n 0.0104464f $X=0.495 $Y=2.825 $X2=0 $Y2=0
cc_243 N_D_M1026_g N_A_30_78#_c_1568_n 0.0108589f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_244 N_D_c_235_n N_A_30_78#_c_1568_n 0.00411346f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_245 N_D_M1018_g N_A_30_78#_c_1574_n 0.00599391f $X=0.495 $Y=2.825 $X2=0 $Y2=0
cc_246 N_D_M1026_g N_A_30_78#_c_1569_n 0.0175726f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_247 N_D_c_235_n N_A_30_78#_c_1569_n 0.0884076f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_248 N_D_M1026_g N_A_30_78#_c_1572_n 0.00806237f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_249 N_D_c_234_n N_A_30_78#_c_1572_n 0.00161806f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_250 N_D_c_235_n N_A_30_78#_c_1572_n 0.0286676f $X=0.385 $Y=1.165 $X2=0 $Y2=0
cc_251 N_D_M1018_g N_A_30_78#_c_1579_n 0.0128371f $X=0.495 $Y=2.825 $X2=0 $Y2=0
cc_252 N_D_M1026_g N_VGND_c_1712_n 0.00190636f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_253 N_D_M1026_g N_VGND_c_1718_n 0.00429844f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_254 N_D_M1026_g N_VGND_c_1728_n 0.00539454f $X=0.51 $Y=0.6 $X2=0 $Y2=0
cc_255 N_CLK_M1021_g N_RESET_B_c_591_n 0.00732518f $X=1.925 $Y=2.495 $X2=0 $Y2=0
cc_256 N_CLK_c_265_n N_RESET_B_c_591_n 0.00731614f $X=1.91 $Y=1.61 $X2=0 $Y2=0
cc_257 N_CLK_c_266_n N_RESET_B_c_592_n 0.0104164f $X=1.91 $Y=1.445 $X2=0 $Y2=0
cc_258 N_CLK_M1021_g N_RESET_B_c_606_n 0.00664186f $X=1.925 $Y=2.495 $X2=0 $Y2=0
cc_259 CLK N_RESET_B_c_606_n 0.0148408f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_260 N_CLK_c_265_n N_RESET_B_c_606_n 2.28173e-19 $X=1.91 $Y=1.61 $X2=0 $Y2=0
cc_261 N_CLK_c_266_n N_RESET_B_c_598_n 0.0037388f $X=1.91 $Y=1.445 $X2=0 $Y2=0
cc_262 CLK N_A_299_387#_M1023_s 5.48149e-19 $X=2.075 $Y=1.58 $X2=-0.19
+ $Y2=-0.245
cc_263 N_CLK_M1021_g N_A_299_387#_M1025_g 0.0511553f $X=1.925 $Y=2.495 $X2=0
+ $Y2=0
cc_264 CLK N_A_299_387#_c_934_n 7.66037e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_265 N_CLK_c_266_n N_A_299_387#_c_934_n 0.0187918f $X=1.91 $Y=1.445 $X2=0
+ $Y2=0
cc_266 CLK N_A_299_387#_c_936_n 0.00368307f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_267 N_CLK_c_265_n N_A_299_387#_c_936_n 0.0214802f $X=1.91 $Y=1.61 $X2=0 $Y2=0
cc_268 N_CLK_c_266_n N_A_299_387#_c_936_n 0.00174202f $X=1.91 $Y=1.445 $X2=0
+ $Y2=0
cc_269 N_CLK_c_266_n N_A_299_387#_c_941_n 0.00108005f $X=1.91 $Y=1.445 $X2=0
+ $Y2=0
cc_270 N_CLK_M1021_g N_A_299_387#_c_942_n 0.00368352f $X=1.925 $Y=2.495 $X2=0
+ $Y2=0
cc_271 CLK N_A_299_387#_c_942_n 0.0368639f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_272 N_CLK_c_265_n N_A_299_387#_c_942_n 0.00288465f $X=1.91 $Y=1.61 $X2=0
+ $Y2=0
cc_273 N_CLK_c_266_n N_A_299_387#_c_942_n 0.00340676f $X=1.91 $Y=1.445 $X2=0
+ $Y2=0
cc_274 CLK N_A_299_387#_c_971_n 0.0258828f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_275 N_CLK_c_266_n N_A_299_387#_c_971_n 0.0129975f $X=1.91 $Y=1.445 $X2=0
+ $Y2=0
cc_276 CLK N_A_299_387#_c_943_n 0.0328411f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_277 N_CLK_c_265_n N_A_299_387#_c_943_n 2.23279e-19 $X=1.91 $Y=1.61 $X2=0
+ $Y2=0
cc_278 N_CLK_c_266_n N_A_299_387#_c_943_n 0.00102506f $X=1.91 $Y=1.445 $X2=0
+ $Y2=0
cc_279 CLK N_A_299_387#_c_944_n 0.00242903f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_280 N_CLK_c_265_n N_A_299_387#_c_944_n 0.0021895f $X=1.91 $Y=1.61 $X2=0 $Y2=0
cc_281 N_CLK_M1021_g N_A_299_387#_c_958_n 0.00525582f $X=1.925 $Y=2.495 $X2=0
+ $Y2=0
cc_282 N_CLK_c_265_n N_A_299_387#_c_958_n 0.00147562f $X=1.91 $Y=1.61 $X2=0
+ $Y2=0
cc_283 N_CLK_M1021_g N_VPWR_c_1434_n 0.00615221f $X=1.925 $Y=2.495 $X2=0 $Y2=0
cc_284 N_CLK_M1021_g N_VPWR_c_1435_n 0.0109019f $X=1.925 $Y=2.495 $X2=0 $Y2=0
cc_285 N_CLK_M1021_g N_VPWR_c_1445_n 0.0040249f $X=1.925 $Y=2.495 $X2=0 $Y2=0
cc_286 N_CLK_M1021_g N_VPWR_c_1431_n 0.0059177f $X=1.925 $Y=2.495 $X2=0 $Y2=0
cc_287 N_CLK_M1021_g N_A_30_78#_c_1576_n 0.0177613f $X=1.925 $Y=2.495 $X2=0
+ $Y2=0
cc_288 CLK N_A_30_78#_c_1576_n 0.0041586f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_289 N_CLK_c_265_n N_A_30_78#_c_1576_n 2.11571e-19 $X=1.91 $Y=1.61 $X2=0 $Y2=0
cc_290 CLK N_VGND_M1023_d 0.00227476f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_291 N_CLK_c_266_n N_VGND_c_1712_n 0.00226704f $X=1.91 $Y=1.445 $X2=0 $Y2=0
cc_292 N_CLK_c_266_n N_VGND_c_1713_n 0.00293245f $X=1.91 $Y=1.445 $X2=0 $Y2=0
cc_293 N_CLK_c_266_n N_VGND_c_1728_n 9.39239e-19 $X=1.91 $Y=1.445 $X2=0 $Y2=0
cc_294 N_A_493_387#_c_318_n N_A_833_400#_M1031_d 0.00330812f $X=5.48 $Y=0.65
+ $X2=-0.19 $Y2=-0.245
cc_295 N_A_493_387#_c_338_p N_A_833_400#_M1031_d 0.00218198f $X=5.565 $Y=0.565
+ $X2=-0.19 $Y2=-0.245
cc_296 N_A_493_387#_c_320_n N_A_833_400#_M1031_d 0.00764003f $X=7.25 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_297 N_A_493_387#_c_310_n N_A_833_400#_c_506_n 0.00241246f $X=4.03 $Y=1.435
+ $X2=0 $Y2=0
cc_298 N_A_493_387#_c_328_n N_A_833_400#_c_506_n 0.00302769f $X=3.337 $Y=1.76
+ $X2=0 $Y2=0
cc_299 N_A_493_387#_M1014_g N_A_833_400#_M1008_g 0.00125103f $X=3.415 $Y=2.525
+ $X2=0 $Y2=0
cc_300 N_A_493_387#_c_310_n N_A_833_400#_M1012_g 0.00734359f $X=4.03 $Y=1.435
+ $X2=0 $Y2=0
cc_301 N_A_493_387#_M1002_g N_A_833_400#_M1012_g 0.0603967f $X=4.03 $Y=0.9 $X2=0
+ $Y2=0
cc_302 N_A_493_387#_c_317_n N_A_833_400#_M1012_g 0.00198166f $X=4.395 $Y=0.565
+ $X2=0 $Y2=0
cc_303 N_A_493_387#_c_319_n N_A_833_400#_M1012_g 0.00653413f $X=4.48 $Y=0.65
+ $X2=0 $Y2=0
cc_304 N_A_493_387#_c_310_n N_A_833_400#_c_503_n 5.4926e-19 $X=4.03 $Y=1.435
+ $X2=0 $Y2=0
cc_305 N_A_493_387#_M1002_g N_A_833_400#_c_503_n 0.00243635f $X=4.03 $Y=0.9
+ $X2=0 $Y2=0
cc_306 N_A_493_387#_c_318_n N_A_833_400#_c_524_n 0.0642391f $X=5.48 $Y=0.65
+ $X2=0 $Y2=0
cc_307 N_A_493_387#_c_319_n N_A_833_400#_c_524_n 0.00181597f $X=4.48 $Y=0.65
+ $X2=0 $Y2=0
cc_308 N_A_493_387#_c_320_n N_A_833_400#_c_524_n 0.00571426f $X=7.25 $Y=0.34
+ $X2=0 $Y2=0
cc_309 N_A_493_387#_c_319_n N_A_833_400#_c_527_n 0.0103082f $X=4.48 $Y=0.65
+ $X2=0 $Y2=0
cc_310 N_A_493_387#_c_314_n N_A_833_400#_c_510_n 0.00391868f $X=6.33 $Y=1.27
+ $X2=0 $Y2=0
cc_311 N_A_493_387#_c_312_n N_A_833_400#_c_504_n 0.00184952f $X=6.255 $Y=1.195
+ $X2=0 $Y2=0
cc_312 N_A_493_387#_c_318_n N_A_833_400#_c_504_n 0.00596144f $X=5.48 $Y=0.65
+ $X2=0 $Y2=0
cc_313 N_A_493_387#_c_320_n N_A_833_400#_c_504_n 0.0168368f $X=7.25 $Y=0.34
+ $X2=0 $Y2=0
cc_314 N_A_493_387#_c_314_n N_A_833_400#_c_505_n 0.00184952f $X=6.33 $Y=1.27
+ $X2=0 $Y2=0
cc_315 N_A_493_387#_M1002_g N_RESET_B_c_592_n 0.00530602f $X=4.03 $Y=0.9 $X2=0
+ $Y2=0
cc_316 N_A_493_387#_c_316_n N_RESET_B_c_592_n 0.0272042f $X=4.31 $Y=0.34 $X2=0
+ $Y2=0
cc_317 N_A_493_387#_c_318_n N_RESET_B_c_592_n 0.00262578f $X=5.48 $Y=0.65 $X2=0
+ $Y2=0
cc_318 N_A_493_387#_c_325_n N_RESET_B_c_592_n 0.0118629f $X=2.792 $Y=0.34 $X2=0
+ $Y2=0
cc_319 N_A_493_387#_c_316_n N_RESET_B_M1006_g 0.00423981f $X=4.31 $Y=0.34 $X2=0
+ $Y2=0
cc_320 N_A_493_387#_c_317_n N_RESET_B_M1006_g 0.00439495f $X=4.395 $Y=0.565
+ $X2=0 $Y2=0
cc_321 N_A_493_387#_c_318_n N_RESET_B_M1006_g 0.0122094f $X=5.48 $Y=0.65 $X2=0
+ $Y2=0
cc_322 N_A_493_387#_c_338_p N_RESET_B_M1006_g 6.19914e-19 $X=5.565 $Y=0.565
+ $X2=0 $Y2=0
cc_323 N_A_493_387#_M1025_d N_RESET_B_c_606_n 9.76131e-19 $X=2.465 $Y=1.935
+ $X2=0 $Y2=0
cc_324 N_A_493_387#_M1014_g N_RESET_B_c_606_n 0.00320728f $X=3.415 $Y=2.525
+ $X2=0 $Y2=0
cc_325 N_A_493_387#_c_309_n N_RESET_B_c_606_n 0.00446894f $X=3.83 $Y=1.76 $X2=0
+ $Y2=0
cc_326 N_A_493_387#_c_324_n N_RESET_B_c_606_n 0.0514449f $X=2.945 $Y=1.925 $X2=0
+ $Y2=0
cc_327 N_A_493_387#_c_328_n N_RESET_B_c_606_n 0.00311319f $X=3.337 $Y=1.76 $X2=0
+ $Y2=0
cc_328 N_A_493_387#_c_322_n N_RESET_B_c_608_n 0.0220527f $X=7.13 $Y=2.14 $X2=0
+ $Y2=0
cc_329 N_A_493_387#_c_336_n N_RESET_B_c_608_n 0.00268118f $X=7.265 $Y=2.14 $X2=0
+ $Y2=0
cc_330 N_A_493_387#_c_312_n N_A_701_463#_M1031_g 0.00895705f $X=6.255 $Y=1.195
+ $X2=0 $Y2=0
cc_331 N_A_493_387#_c_318_n N_A_701_463#_M1031_g 0.0118282f $X=5.48 $Y=0.65
+ $X2=0 $Y2=0
cc_332 N_A_493_387#_c_338_p N_A_701_463#_M1031_g 0.0047339f $X=5.565 $Y=0.565
+ $X2=0 $Y2=0
cc_333 N_A_493_387#_c_321_n N_A_701_463#_M1031_g 0.00591041f $X=5.65 $Y=0.34
+ $X2=0 $Y2=0
cc_334 N_A_493_387#_M1014_g N_A_701_463#_c_814_n 0.00358967f $X=3.415 $Y=2.525
+ $X2=0 $Y2=0
cc_335 N_A_493_387#_c_309_n N_A_701_463#_c_814_n 0.00101726f $X=3.83 $Y=1.76
+ $X2=0 $Y2=0
cc_336 N_A_493_387#_c_314_n N_A_701_463#_c_809_n 0.00168855f $X=6.33 $Y=1.27
+ $X2=0 $Y2=0
cc_337 N_A_493_387#_c_309_n N_A_701_463#_c_810_n 0.00151485f $X=3.83 $Y=1.76
+ $X2=0 $Y2=0
cc_338 N_A_493_387#_c_310_n N_A_701_463#_c_810_n 0.00288816f $X=4.03 $Y=1.435
+ $X2=0 $Y2=0
cc_339 N_A_493_387#_M1002_g N_A_701_463#_c_810_n 0.00929992f $X=4.03 $Y=0.9
+ $X2=0 $Y2=0
cc_340 N_A_493_387#_c_316_n N_A_701_463#_c_810_n 0.0328447f $X=4.31 $Y=0.34
+ $X2=0 $Y2=0
cc_341 N_A_493_387#_c_319_n N_A_701_463#_c_810_n 0.00854511f $X=4.48 $Y=0.65
+ $X2=0 $Y2=0
cc_342 N_A_493_387#_M1014_g N_A_701_463#_c_811_n 3.85628e-19 $X=3.415 $Y=2.525
+ $X2=0 $Y2=0
cc_343 N_A_493_387#_c_310_n N_A_701_463#_c_811_n 0.014385f $X=4.03 $Y=1.435
+ $X2=0 $Y2=0
cc_344 N_A_493_387#_M1002_g N_A_701_463#_c_811_n 0.0100691f $X=4.03 $Y=0.9 $X2=0
+ $Y2=0
cc_345 N_A_493_387#_c_324_n N_A_299_387#_M1025_g 0.00166699f $X=2.945 $Y=1.925
+ $X2=0 $Y2=0
cc_346 N_A_493_387#_c_315_n N_A_299_387#_c_934_n 0.00537196f $X=2.945 $Y=1.575
+ $X2=0 $Y2=0
cc_347 N_A_493_387#_c_325_n N_A_299_387#_c_934_n 0.00313928f $X=2.792 $Y=0.34
+ $X2=0 $Y2=0
cc_348 N_A_493_387#_M1014_g N_A_299_387#_c_946_n 0.0202399f $X=3.415 $Y=2.525
+ $X2=0 $Y2=0
cc_349 N_A_493_387#_c_324_n N_A_299_387#_c_946_n 0.020856f $X=2.945 $Y=1.925
+ $X2=0 $Y2=0
cc_350 N_A_493_387#_M1014_g N_A_299_387#_c_947_n 0.0123549f $X=3.415 $Y=2.525
+ $X2=0 $Y2=0
cc_351 N_A_493_387#_c_310_n N_A_299_387#_c_935_n 0.00244951f $X=4.03 $Y=1.435
+ $X2=0 $Y2=0
cc_352 N_A_493_387#_c_324_n N_A_299_387#_c_935_n 0.00778364f $X=2.945 $Y=1.925
+ $X2=0 $Y2=0
cc_353 N_A_493_387#_c_328_n N_A_299_387#_c_935_n 0.0284449f $X=3.337 $Y=1.76
+ $X2=0 $Y2=0
cc_354 N_A_493_387#_c_315_n N_A_299_387#_c_936_n 0.0168867f $X=2.945 $Y=1.575
+ $X2=0 $Y2=0
cc_355 N_A_493_387#_c_324_n N_A_299_387#_c_936_n 0.0112143f $X=2.945 $Y=1.925
+ $X2=0 $Y2=0
cc_356 N_A_493_387#_c_325_n N_A_299_387#_c_936_n 0.00537248f $X=2.792 $Y=0.34
+ $X2=0 $Y2=0
cc_357 N_A_493_387#_c_328_n N_A_299_387#_c_936_n 0.0213791f $X=3.337 $Y=1.76
+ $X2=0 $Y2=0
cc_358 N_A_493_387#_M1002_g N_A_299_387#_M1007_g 0.0175066f $X=4.03 $Y=0.9 $X2=0
+ $Y2=0
cc_359 N_A_493_387#_c_315_n N_A_299_387#_M1007_g 4.88505e-19 $X=2.945 $Y=1.575
+ $X2=0 $Y2=0
cc_360 N_A_493_387#_c_316_n N_A_299_387#_M1007_g 0.00315349f $X=4.31 $Y=0.34
+ $X2=0 $Y2=0
cc_361 N_A_493_387#_c_325_n N_A_299_387#_M1007_g 0.00248325f $X=2.792 $Y=0.34
+ $X2=0 $Y2=0
cc_362 N_A_493_387#_M1014_g N_A_299_387#_M1022_g 0.0167726f $X=3.415 $Y=2.525
+ $X2=0 $Y2=0
cc_363 N_A_493_387#_c_309_n N_A_299_387#_M1022_g 0.00727013f $X=3.83 $Y=1.76
+ $X2=0 $Y2=0
cc_364 N_A_493_387#_M1010_g N_A_299_387#_M1004_g 0.00551007f $X=7.265 $Y=2.675
+ $X2=0 $Y2=0
cc_365 N_A_493_387#_c_336_n N_A_299_387#_M1004_g 0.00690574f $X=7.265 $Y=2.14
+ $X2=0 $Y2=0
cc_366 N_A_493_387#_c_313_n N_A_299_387#_c_938_n 0.0196707f $X=6.69 $Y=1.27
+ $X2=0 $Y2=0
cc_367 N_A_493_387#_c_322_n N_A_299_387#_c_938_n 0.0164562f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_368 N_A_493_387#_c_327_n N_A_299_387#_c_938_n 0.00266664f $X=7.335 $Y=1.18
+ $X2=0 $Y2=0
cc_369 N_A_493_387#_c_336_n N_A_299_387#_c_938_n 0.0220885f $X=7.265 $Y=2.14
+ $X2=0 $Y2=0
cc_370 N_A_493_387#_c_314_n N_A_299_387#_c_939_n 0.0196707f $X=6.33 $Y=1.27
+ $X2=0 $Y2=0
cc_371 N_A_493_387#_c_320_n N_A_299_387#_M1016_g 0.0088085f $X=7.25 $Y=0.34
+ $X2=0 $Y2=0
cc_372 N_A_493_387#_c_322_n N_A_299_387#_M1016_g 0.00923892f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_373 N_A_493_387#_c_323_n N_A_299_387#_M1016_g 0.0233298f $X=7.335 $Y=1.015
+ $X2=0 $Y2=0
cc_374 N_A_493_387#_c_326_n N_A_299_387#_M1016_g 0.0213806f $X=6.855 $Y=1.18
+ $X2=0 $Y2=0
cc_375 N_A_493_387#_c_327_n N_A_299_387#_M1016_g 0.011895f $X=7.335 $Y=1.18
+ $X2=0 $Y2=0
cc_376 N_A_493_387#_M1001_d N_A_299_387#_c_971_n 0.00269359f $X=2.55 $Y=0.595
+ $X2=0 $Y2=0
cc_377 N_A_493_387#_c_315_n N_A_299_387#_c_971_n 0.0137394f $X=2.945 $Y=1.575
+ $X2=0 $Y2=0
cc_378 N_A_493_387#_c_325_n N_A_299_387#_c_971_n 0.00692369f $X=2.792 $Y=0.34
+ $X2=0 $Y2=0
cc_379 N_A_493_387#_M1001_d N_A_299_387#_c_943_n 0.00205608f $X=2.55 $Y=0.595
+ $X2=0 $Y2=0
cc_380 N_A_493_387#_c_315_n N_A_299_387#_c_943_n 0.0320469f $X=2.945 $Y=1.575
+ $X2=0 $Y2=0
cc_381 N_A_493_387#_c_324_n N_A_299_387#_c_943_n 0.0276081f $X=2.945 $Y=1.925
+ $X2=0 $Y2=0
cc_382 N_A_493_387#_c_322_n N_A_1518_203#_M1015_g 3.63622e-19 $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_383 N_A_493_387#_c_336_n N_A_1518_203#_M1015_g 0.0562924f $X=7.265 $Y=2.14
+ $X2=0 $Y2=0
cc_384 N_A_493_387#_c_320_n N_A_1518_203#_M1013_g 0.00107872f $X=7.25 $Y=0.34
+ $X2=0 $Y2=0
cc_385 N_A_493_387#_c_323_n N_A_1518_203#_M1013_g 0.0045389f $X=7.335 $Y=1.015
+ $X2=0 $Y2=0
cc_386 N_A_493_387#_c_322_n N_A_1518_203#_c_1112_n 0.00240511f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_387 N_A_493_387#_c_327_n N_A_1518_203#_c_1116_n 0.0276613f $X=7.335 $Y=1.18
+ $X2=0 $Y2=0
cc_388 N_A_493_387#_c_327_n N_A_1518_203#_c_1117_n 0.00201148f $X=7.335 $Y=1.18
+ $X2=0 $Y2=0
cc_389 N_A_493_387#_c_320_n N_A_1266_74#_M1027_d 0.00949775f $X=7.25 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_390 N_A_493_387#_c_312_n N_A_1266_74#_c_1250_n 0.0033591f $X=6.255 $Y=1.195
+ $X2=0 $Y2=0
cc_391 N_A_493_387#_c_318_n N_A_1266_74#_c_1250_n 0.00205017f $X=5.48 $Y=0.65
+ $X2=0 $Y2=0
cc_392 N_A_493_387#_c_320_n N_A_1266_74#_c_1250_n 0.00851496f $X=7.25 $Y=0.34
+ $X2=0 $Y2=0
cc_393 N_A_493_387#_c_312_n N_A_1266_74#_c_1233_n 0.00750067f $X=6.255 $Y=1.195
+ $X2=0 $Y2=0
cc_394 N_A_493_387#_c_313_n N_A_1266_74#_c_1233_n 0.00921579f $X=6.69 $Y=1.27
+ $X2=0 $Y2=0
cc_395 N_A_493_387#_c_314_n N_A_1266_74#_c_1233_n 0.00149681f $X=6.33 $Y=1.27
+ $X2=0 $Y2=0
cc_396 N_A_493_387#_c_322_n N_A_1266_74#_c_1233_n 0.00662434f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_397 N_A_493_387#_c_326_n N_A_1266_74#_c_1233_n 6.18001e-19 $X=6.855 $Y=1.18
+ $X2=0 $Y2=0
cc_398 N_A_493_387#_c_327_n N_A_1266_74#_c_1233_n 0.0224751f $X=7.335 $Y=1.18
+ $X2=0 $Y2=0
cc_399 N_A_493_387#_M1010_g N_A_1266_74#_c_1244_n 0.00266968f $X=7.265 $Y=2.675
+ $X2=0 $Y2=0
cc_400 N_A_493_387#_c_322_n N_A_1266_74#_c_1244_n 0.0279378f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_401 N_A_493_387#_c_336_n N_A_1266_74#_c_1244_n 0.00232018f $X=7.265 $Y=2.14
+ $X2=0 $Y2=0
cc_402 N_A_493_387#_c_313_n N_A_1266_74#_c_1234_n 0.00430336f $X=6.69 $Y=1.27
+ $X2=0 $Y2=0
cc_403 N_A_493_387#_c_320_n N_A_1266_74#_c_1234_n 0.0414158f $X=7.25 $Y=0.34
+ $X2=0 $Y2=0
cc_404 N_A_493_387#_c_323_n N_A_1266_74#_c_1234_n 0.0196081f $X=7.335 $Y=1.015
+ $X2=0 $Y2=0
cc_405 N_A_493_387#_c_326_n N_A_1266_74#_c_1234_n 0.00746605f $X=6.855 $Y=1.18
+ $X2=0 $Y2=0
cc_406 N_A_493_387#_c_327_n N_A_1266_74#_c_1234_n 0.030444f $X=7.335 $Y=1.18
+ $X2=0 $Y2=0
cc_407 N_A_493_387#_M1010_g N_A_1266_74#_c_1267_n 0.0146227f $X=7.265 $Y=2.675
+ $X2=0 $Y2=0
cc_408 N_A_493_387#_c_322_n N_A_1266_74#_c_1267_n 0.0232328f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_409 N_A_493_387#_c_336_n N_A_1266_74#_c_1267_n 0.00140365f $X=7.265 $Y=2.14
+ $X2=0 $Y2=0
cc_410 N_A_493_387#_c_322_n N_A_1266_74#_c_1245_n 0.0462528f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_411 N_A_493_387#_c_336_n N_A_1266_74#_c_1245_n 0.00567651f $X=7.265 $Y=2.14
+ $X2=0 $Y2=0
cc_412 N_A_493_387#_c_322_n N_A_1266_74#_c_1236_n 0.0142973f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_413 N_A_493_387#_c_313_n N_A_1266_74#_c_1237_n 0.0016242f $X=6.69 $Y=1.27
+ $X2=0 $Y2=0
cc_414 N_A_493_387#_c_322_n N_A_1266_74#_c_1237_n 0.00830682f $X=7.13 $Y=2.14
+ $X2=0 $Y2=0
cc_415 N_A_493_387#_M1010_g N_VPWR_c_1447_n 0.00469675f $X=7.265 $Y=2.675 $X2=0
+ $Y2=0
cc_416 N_A_493_387#_M1014_g N_VPWR_c_1431_n 0.00112709f $X=3.415 $Y=2.525 $X2=0
+ $Y2=0
cc_417 N_A_493_387#_M1010_g N_VPWR_c_1431_n 0.00626544f $X=7.265 $Y=2.675 $X2=0
+ $Y2=0
cc_418 N_A_493_387#_M1025_d N_A_30_78#_c_1576_n 0.0060793f $X=2.465 $Y=1.935
+ $X2=0 $Y2=0
cc_419 N_A_493_387#_c_324_n N_A_30_78#_c_1576_n 0.0332008f $X=2.945 $Y=1.925
+ $X2=0 $Y2=0
cc_420 N_A_493_387#_M1002_g N_A_30_78#_c_1570_n 3.15604e-19 $X=4.03 $Y=0.9 $X2=0
+ $Y2=0
cc_421 N_A_493_387#_c_316_n N_A_30_78#_c_1570_n 0.0224516f $X=4.31 $Y=0.34 $X2=0
+ $Y2=0
cc_422 N_A_493_387#_c_325_n N_A_30_78#_c_1570_n 0.0483059f $X=2.792 $Y=0.34
+ $X2=0 $Y2=0
cc_423 N_A_493_387#_M1014_g N_A_30_78#_c_1577_n 0.0150772f $X=3.415 $Y=2.525
+ $X2=0 $Y2=0
cc_424 N_A_493_387#_c_309_n N_A_30_78#_c_1577_n 0.00251615f $X=3.83 $Y=1.76
+ $X2=0 $Y2=0
cc_425 N_A_493_387#_c_324_n N_A_30_78#_c_1577_n 0.00718765f $X=2.945 $Y=1.925
+ $X2=0 $Y2=0
cc_426 N_A_493_387#_c_309_n N_A_30_78#_c_1571_n 0.0132826f $X=3.83 $Y=1.76 $X2=0
+ $Y2=0
cc_427 N_A_493_387#_c_310_n N_A_30_78#_c_1571_n 0.005114f $X=4.03 $Y=1.435 $X2=0
+ $Y2=0
cc_428 N_A_493_387#_M1002_g N_A_30_78#_c_1571_n 2.04804e-19 $X=4.03 $Y=0.9 $X2=0
+ $Y2=0
cc_429 N_A_493_387#_c_315_n N_A_30_78#_c_1571_n 0.00580219f $X=2.945 $Y=1.575
+ $X2=0 $Y2=0
cc_430 N_A_493_387#_c_324_n N_A_30_78#_c_1571_n 0.0380096f $X=2.945 $Y=1.925
+ $X2=0 $Y2=0
cc_431 N_A_493_387#_c_328_n N_A_30_78#_c_1571_n 0.00455231f $X=3.337 $Y=1.76
+ $X2=0 $Y2=0
cc_432 N_A_493_387#_M1014_g N_A_30_78#_c_1580_n 2.18709e-19 $X=3.415 $Y=2.525
+ $X2=0 $Y2=0
cc_433 N_A_493_387#_c_324_n N_A_30_78#_c_1580_n 0.0217947f $X=2.945 $Y=1.925
+ $X2=0 $Y2=0
cc_434 N_A_493_387#_c_328_n N_A_30_78#_c_1580_n 0.00104726f $X=3.337 $Y=1.76
+ $X2=0 $Y2=0
cc_435 N_A_493_387#_c_309_n N_A_30_78#_c_1573_n 4.93811e-19 $X=3.83 $Y=1.76
+ $X2=0 $Y2=0
cc_436 N_A_493_387#_M1002_g N_A_30_78#_c_1573_n 6.43133e-19 $X=4.03 $Y=0.9 $X2=0
+ $Y2=0
cc_437 N_A_493_387#_c_315_n N_A_30_78#_c_1573_n 0.0136584f $X=2.945 $Y=1.575
+ $X2=0 $Y2=0
cc_438 N_A_493_387#_c_324_n N_A_30_78#_c_1573_n 0.014334f $X=2.945 $Y=1.925
+ $X2=0 $Y2=0
cc_439 N_A_493_387#_c_328_n N_A_30_78#_c_1573_n 0.00115865f $X=3.337 $Y=1.76
+ $X2=0 $Y2=0
cc_440 N_A_493_387#_c_318_n N_VGND_M1006_d 0.00922416f $X=5.48 $Y=0.65 $X2=0
+ $Y2=0
cc_441 N_A_493_387#_c_325_n N_VGND_c_1713_n 0.0381058f $X=2.792 $Y=0.34 $X2=0
+ $Y2=0
cc_442 N_A_493_387#_c_320_n N_VGND_c_1714_n 0.00831292f $X=7.25 $Y=0.34 $X2=0
+ $Y2=0
cc_443 N_A_493_387#_c_323_n N_VGND_c_1714_n 0.00983536f $X=7.335 $Y=1.015 $X2=0
+ $Y2=0
cc_444 N_A_493_387#_c_316_n N_VGND_c_1721_n 0.0998821f $X=4.31 $Y=0.34 $X2=0
+ $Y2=0
cc_445 N_A_493_387#_c_318_n N_VGND_c_1721_n 0.0381943f $X=5.48 $Y=0.65 $X2=0
+ $Y2=0
cc_446 N_A_493_387#_c_321_n N_VGND_c_1721_n 0.0107916f $X=5.65 $Y=0.34 $X2=0
+ $Y2=0
cc_447 N_A_493_387#_c_325_n N_VGND_c_1721_n 0.0326115f $X=2.792 $Y=0.34 $X2=0
+ $Y2=0
cc_448 N_A_493_387#_c_312_n N_VGND_c_1722_n 0.00278271f $X=6.255 $Y=1.195 $X2=0
+ $Y2=0
cc_449 N_A_493_387#_c_318_n N_VGND_c_1722_n 0.00286598f $X=5.48 $Y=0.65 $X2=0
+ $Y2=0
cc_450 N_A_493_387#_c_320_n N_VGND_c_1722_n 0.114761f $X=7.25 $Y=0.34 $X2=0
+ $Y2=0
cc_451 N_A_493_387#_c_321_n N_VGND_c_1722_n 0.0117553f $X=5.65 $Y=0.34 $X2=0
+ $Y2=0
cc_452 N_A_493_387#_c_312_n N_VGND_c_1728_n 0.00361111f $X=6.255 $Y=1.195 $X2=0
+ $Y2=0
cc_453 N_A_493_387#_c_316_n N_VGND_c_1728_n 0.0486258f $X=4.31 $Y=0.34 $X2=0
+ $Y2=0
cc_454 N_A_493_387#_c_318_n N_VGND_c_1728_n 0.0180862f $X=5.48 $Y=0.65 $X2=0
+ $Y2=0
cc_455 N_A_493_387#_c_320_n N_VGND_c_1728_n 0.0660751f $X=7.25 $Y=0.34 $X2=0
+ $Y2=0
cc_456 N_A_493_387#_c_321_n N_VGND_c_1728_n 0.00639038f $X=5.65 $Y=0.34 $X2=0
+ $Y2=0
cc_457 N_A_493_387#_c_325_n N_VGND_c_1728_n 0.0165036f $X=2.792 $Y=0.34 $X2=0
+ $Y2=0
cc_458 N_A_493_387#_c_318_n A_894_138# 0.00134267f $X=5.48 $Y=0.65 $X2=-0.19
+ $Y2=-0.245
cc_459 N_A_833_400#_M1012_g N_RESET_B_c_592_n 0.00610028f $X=4.395 $Y=0.9 $X2=0
+ $Y2=0
cc_460 N_A_833_400#_M1012_g N_RESET_B_M1006_g 0.0421141f $X=4.395 $Y=0.9 $X2=0
+ $Y2=0
cc_461 N_A_833_400#_c_503_n N_RESET_B_M1006_g 0.00164083f $X=4.36 $Y=1.96 $X2=0
+ $Y2=0
cc_462 N_A_833_400#_c_524_n N_RESET_B_M1006_g 0.011669f $X=5.82 $Y=0.99 $X2=0
+ $Y2=0
cc_463 N_A_833_400#_c_506_n N_RESET_B_c_602_n 0.0171884f $X=4.255 $Y=2.125 $X2=0
+ $Y2=0
cc_464 N_A_833_400#_M1008_g N_RESET_B_c_602_n 0.0177981f $X=4.255 $Y=2.525 $X2=0
+ $Y2=0
cc_465 N_A_833_400#_c_503_n N_RESET_B_c_602_n 3.33923e-19 $X=4.36 $Y=1.96 $X2=0
+ $Y2=0
cc_466 N_A_833_400#_M1012_g N_RESET_B_c_595_n 0.0141928f $X=4.395 $Y=0.9 $X2=0
+ $Y2=0
cc_467 N_A_833_400#_c_503_n N_RESET_B_c_595_n 6.38323e-19 $X=4.36 $Y=1.96 $X2=0
+ $Y2=0
cc_468 N_A_833_400#_c_524_n N_RESET_B_c_597_n 0.00246935f $X=5.82 $Y=0.99 $X2=0
+ $Y2=0
cc_469 N_A_833_400#_c_506_n N_RESET_B_c_606_n 0.0104284f $X=4.255 $Y=2.125 $X2=0
+ $Y2=0
cc_470 N_A_833_400#_c_503_n N_RESET_B_c_606_n 0.0161444f $X=4.36 $Y=1.96 $X2=0
+ $Y2=0
cc_471 N_A_833_400#_M1029_d N_RESET_B_c_608_n 6.08559e-19 $X=5.97 $Y=1.735 $X2=0
+ $Y2=0
cc_472 N_A_833_400#_c_510_n N_RESET_B_c_608_n 0.0388437f $X=6.145 $Y=2.03 $X2=0
+ $Y2=0
cc_473 N_A_833_400#_c_524_n N_A_701_463#_M1031_g 0.0124811f $X=5.82 $Y=0.99
+ $X2=0 $Y2=0
cc_474 N_A_833_400#_c_504_n N_A_701_463#_M1031_g 0.00563857f $X=5.985 $Y=0.855
+ $X2=0 $Y2=0
cc_475 N_A_833_400#_c_505_n N_A_701_463#_M1031_g 0.0019205f $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_476 N_A_833_400#_c_510_n N_A_701_463#_M1029_g 0.00560705f $X=6.145 $Y=2.03
+ $X2=0 $Y2=0
cc_477 N_A_833_400#_c_506_n N_A_701_463#_c_839_n 0.00348386f $X=4.255 $Y=2.125
+ $X2=0 $Y2=0
cc_478 N_A_833_400#_M1008_g N_A_701_463#_c_839_n 0.00943891f $X=4.255 $Y=2.525
+ $X2=0 $Y2=0
cc_479 N_A_833_400#_c_503_n N_A_701_463#_c_839_n 0.00775184f $X=4.36 $Y=1.96
+ $X2=0 $Y2=0
cc_480 N_A_833_400#_c_506_n N_A_701_463#_c_805_n 0.00206044f $X=4.255 $Y=2.125
+ $X2=0 $Y2=0
cc_481 N_A_833_400#_M1008_g N_A_701_463#_c_805_n 0.0017364f $X=4.255 $Y=2.525
+ $X2=0 $Y2=0
cc_482 N_A_833_400#_M1012_g N_A_701_463#_c_805_n 0.00139327f $X=4.395 $Y=0.9
+ $X2=0 $Y2=0
cc_483 N_A_833_400#_c_503_n N_A_701_463#_c_805_n 0.0385458f $X=4.36 $Y=1.96
+ $X2=0 $Y2=0
cc_484 N_A_833_400#_M1012_g N_A_701_463#_c_806_n 0.00123542f $X=4.395 $Y=0.9
+ $X2=0 $Y2=0
cc_485 N_A_833_400#_c_503_n N_A_701_463#_c_806_n 0.0137157f $X=4.36 $Y=1.96
+ $X2=0 $Y2=0
cc_486 N_A_833_400#_c_524_n N_A_701_463#_c_806_n 0.00734087f $X=5.82 $Y=0.99
+ $X2=0 $Y2=0
cc_487 N_A_833_400#_c_524_n N_A_701_463#_c_807_n 0.0251784f $X=5.82 $Y=0.99
+ $X2=0 $Y2=0
cc_488 N_A_833_400#_c_505_n N_A_701_463#_c_808_n 0.013796f $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_489 N_A_833_400#_c_524_n N_A_701_463#_c_809_n 0.00647112f $X=5.82 $Y=0.99
+ $X2=0 $Y2=0
cc_490 N_A_833_400#_c_504_n N_A_701_463#_c_809_n 0.00600822f $X=5.985 $Y=0.855
+ $X2=0 $Y2=0
cc_491 N_A_833_400#_c_505_n N_A_701_463#_c_809_n 0.00713814f $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_492 N_A_833_400#_M1012_g N_A_701_463#_c_810_n 0.00144193f $X=4.395 $Y=0.9
+ $X2=0 $Y2=0
cc_493 N_A_833_400#_M1008_g N_A_701_463#_c_817_n 0.0108411f $X=4.255 $Y=2.525
+ $X2=0 $Y2=0
cc_494 N_A_833_400#_c_506_n N_A_701_463#_c_811_n 0.00631548f $X=4.255 $Y=2.125
+ $X2=0 $Y2=0
cc_495 N_A_833_400#_M1012_g N_A_701_463#_c_811_n 0.0012738f $X=4.395 $Y=0.9
+ $X2=0 $Y2=0
cc_496 N_A_833_400#_c_503_n N_A_701_463#_c_811_n 0.0739669f $X=4.36 $Y=1.96
+ $X2=0 $Y2=0
cc_497 N_A_833_400#_M1008_g N_A_701_463#_c_819_n 4.25665e-19 $X=4.255 $Y=2.525
+ $X2=0 $Y2=0
cc_498 N_A_833_400#_c_524_n N_A_701_463#_c_812_n 0.0165891f $X=5.82 $Y=0.99
+ $X2=0 $Y2=0
cc_499 N_A_833_400#_M1008_g N_A_299_387#_M1022_g 0.0428347f $X=4.255 $Y=2.525
+ $X2=0 $Y2=0
cc_500 N_A_833_400#_M1008_g N_A_299_387#_c_951_n 0.0118761f $X=4.255 $Y=2.525
+ $X2=0 $Y2=0
cc_501 N_A_833_400#_c_510_n N_A_299_387#_c_951_n 0.00455019f $X=6.145 $Y=2.03
+ $X2=0 $Y2=0
cc_502 N_A_833_400#_c_510_n N_A_299_387#_M1004_g 0.0117311f $X=6.145 $Y=2.03
+ $X2=0 $Y2=0
cc_503 N_A_833_400#_c_505_n N_A_299_387#_c_939_n 0.00239037f $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_504 N_A_833_400#_c_504_n N_A_1266_74#_c_1233_n 0.03852f $X=5.985 $Y=0.855
+ $X2=0 $Y2=0
cc_505 N_A_833_400#_c_510_n N_A_1266_74#_c_1244_n 0.0253543f $X=6.145 $Y=2.03
+ $X2=0 $Y2=0
cc_506 N_A_833_400#_c_505_n N_A_1266_74#_c_1244_n 0.00813908f $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_507 N_A_833_400#_c_505_n N_A_1266_74#_c_1237_n 0.0129729f $X=6.145 $Y=1.865
+ $X2=0 $Y2=0
cc_508 N_A_833_400#_M1008_g N_VPWR_c_1436_n 0.00339674f $X=4.255 $Y=2.525 $X2=0
+ $Y2=0
cc_509 N_A_833_400#_c_524_n N_VPWR_c_1438_n 0.00359959f $X=5.82 $Y=0.99 $X2=0
+ $Y2=0
cc_510 N_A_833_400#_c_510_n N_VPWR_c_1438_n 0.0405057f $X=6.145 $Y=2.03 $X2=0
+ $Y2=0
cc_511 N_A_833_400#_c_510_n N_VPWR_c_1447_n 0.00666645f $X=6.145 $Y=2.03 $X2=0
+ $Y2=0
cc_512 N_A_833_400#_M1008_g N_VPWR_c_1431_n 0.00112709f $X=4.255 $Y=2.525 $X2=0
+ $Y2=0
cc_513 N_A_833_400#_c_510_n N_VPWR_c_1431_n 0.00905011f $X=6.145 $Y=2.03 $X2=0
+ $Y2=0
cc_514 N_A_833_400#_c_524_n N_VGND_M1006_d 0.0107327f $X=5.82 $Y=0.99 $X2=0
+ $Y2=0
cc_515 N_A_833_400#_c_524_n A_894_138# 0.00517725f $X=5.82 $Y=0.99 $X2=-0.19
+ $Y2=-0.245
cc_516 N_RESET_B_c_592_n N_A_701_463#_M1031_g 0.0212385f $X=4.71 $Y=0.18 $X2=0
+ $Y2=0
cc_517 N_RESET_B_c_597_n N_A_701_463#_M1031_g 0.00219471f $X=4.875 $Y=1.26 $X2=0
+ $Y2=0
cc_518 N_RESET_B_c_608_n N_A_701_463#_M1029_g 0.0125673f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_519 N_RESET_B_c_606_n N_A_701_463#_c_814_n 0.00665963f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_520 N_RESET_B_c_606_n N_A_701_463#_c_839_n 0.0102468f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_521 N_RESET_B_c_602_n N_A_701_463#_c_805_n 0.0153662f $X=4.86 $Y=2.275 $X2=0
+ $Y2=0
cc_522 N_RESET_B_c_595_n N_A_701_463#_c_805_n 0.0056545f $X=4.875 $Y=1.795 $X2=0
+ $Y2=0
cc_523 N_RESET_B_c_606_n N_A_701_463#_c_805_n 0.0206062f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_524 N_RESET_B_c_609_n N_A_701_463#_c_805_n 0.00237384f $X=5.185 $Y=2.035
+ $X2=0 $Y2=0
cc_525 N_RESET_B_c_610_n N_A_701_463#_c_805_n 0.0234789f $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_526 N_RESET_B_c_597_n N_A_701_463#_c_806_n 0.00235031f $X=4.875 $Y=1.26 $X2=0
+ $Y2=0
cc_527 N_RESET_B_c_597_n N_A_701_463#_c_807_n 0.00287348f $X=4.875 $Y=1.26 $X2=0
+ $Y2=0
cc_528 N_RESET_B_c_608_n N_A_701_463#_c_807_n 0.00696682f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_529 N_RESET_B_c_608_n N_A_701_463#_c_808_n 7.66226e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_530 N_RESET_B_c_597_n N_A_701_463#_c_809_n 0.0104866f $X=4.875 $Y=1.26 $X2=0
+ $Y2=0
cc_531 N_RESET_B_c_608_n N_A_701_463#_c_809_n 0.00379376f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_532 N_RESET_B_c_602_n N_A_701_463#_c_817_n 9.30965e-19 $X=4.86 $Y=2.275 $X2=0
+ $Y2=0
cc_533 N_RESET_B_c_606_n N_A_701_463#_c_817_n 0.00460206f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_534 N_RESET_B_c_606_n N_A_701_463#_c_811_n 0.0184579f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_535 N_RESET_B_c_602_n N_A_701_463#_c_819_n 0.0139724f $X=4.86 $Y=2.275 $X2=0
+ $Y2=0
cc_536 N_RESET_B_c_606_n N_A_701_463#_c_819_n 0.00411593f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_537 N_RESET_B_c_608_n N_A_701_463#_c_819_n 4.71937e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_538 N_RESET_B_c_609_n N_A_701_463#_c_819_n 0.00893678f $X=5.185 $Y=2.035
+ $X2=0 $Y2=0
cc_539 N_RESET_B_c_610_n N_A_701_463#_c_819_n 0.019232f $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_540 N_RESET_B_c_602_n N_A_701_463#_c_812_n 0.00769376f $X=4.86 $Y=2.275 $X2=0
+ $Y2=0
cc_541 N_RESET_B_c_595_n N_A_701_463#_c_812_n 0.0118026f $X=4.875 $Y=1.795 $X2=0
+ $Y2=0
cc_542 N_RESET_B_c_597_n N_A_701_463#_c_812_n 2.01544e-19 $X=4.875 $Y=1.26 $X2=0
+ $Y2=0
cc_543 N_RESET_B_c_606_n N_A_701_463#_c_812_n 0.0032742f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_544 N_RESET_B_c_608_n N_A_701_463#_c_812_n 5.46313e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_545 N_RESET_B_c_609_n N_A_701_463#_c_812_n 0.00327889f $X=5.185 $Y=2.035
+ $X2=0 $Y2=0
cc_546 N_RESET_B_c_610_n N_A_701_463#_c_812_n 0.0188004f $X=5.04 $Y=2.035 $X2=0
+ $Y2=0
cc_547 N_RESET_B_c_606_n N_A_299_387#_M1021_s 9.41382e-19 $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_548 N_RESET_B_c_606_n N_A_299_387#_M1025_g 0.0100292f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_549 N_RESET_B_c_592_n N_A_299_387#_c_934_n 0.0104164f $X=4.71 $Y=0.18 $X2=0
+ $Y2=0
cc_550 N_RESET_B_c_606_n N_A_299_387#_c_935_n 3.18309e-19 $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_551 N_RESET_B_c_592_n N_A_299_387#_M1007_g 0.00530602f $X=4.71 $Y=0.18 $X2=0
+ $Y2=0
cc_552 N_RESET_B_c_606_n N_A_299_387#_M1022_g 0.00254899f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_553 N_RESET_B_c_602_n N_A_299_387#_c_951_n 0.0119613f $X=4.86 $Y=2.275 $X2=0
+ $Y2=0
cc_554 N_RESET_B_c_608_n N_A_299_387#_M1004_g 0.00983659f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_555 N_RESET_B_c_608_n N_A_299_387#_c_938_n 0.00802201f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_556 N_RESET_B_M1009_g N_A_299_387#_c_941_n 0.00279512f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_557 N_RESET_B_c_592_n N_A_299_387#_c_941_n 0.00848569f $X=4.71 $Y=0.18 $X2=0
+ $Y2=0
cc_558 N_RESET_B_c_606_n N_A_299_387#_c_942_n 0.00308596f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_559 N_RESET_B_c_607_n N_A_299_387#_c_942_n 7.65024e-19 $X=1.345 $Y=2.035
+ $X2=0 $Y2=0
cc_560 N_RESET_B_c_598_n N_A_299_387#_c_942_n 0.00796133f $X=1.155 $Y=1.295
+ $X2=0 $Y2=0
cc_561 N_RESET_B_c_599_n N_A_299_387#_c_942_n 0.0590176f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_562 N_RESET_B_c_606_n N_A_299_387#_c_943_n 0.00375674f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_563 N_RESET_B_M1009_g N_A_299_387#_c_944_n 0.00122712f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_564 N_RESET_B_c_599_n N_A_299_387#_c_944_n 8.29766e-19 $X=1.155 $Y=1.295
+ $X2=0 $Y2=0
cc_565 N_RESET_B_M1019_g N_A_299_387#_c_958_n 0.00245957f $X=0.945 $Y=2.825
+ $X2=0 $Y2=0
cc_566 N_RESET_B_c_606_n N_A_299_387#_c_958_n 0.0235216f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_567 N_RESET_B_c_607_n N_A_299_387#_c_958_n 0.00206236f $X=1.345 $Y=2.035
+ $X2=0 $Y2=0
cc_568 N_RESET_B_c_599_n N_A_299_387#_c_958_n 0.0132215f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_569 N_RESET_B_c_613_n N_A_299_387#_c_958_n 0.00153975f $X=1.155 $Y=1.975
+ $X2=0 $Y2=0
cc_570 N_RESET_B_M1000_g N_A_1518_203#_c_1119_n 0.00652196f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_571 N_RESET_B_M1020_g N_A_1518_203#_M1015_g 0.0143049f $X=8.26 $Y=2.675 $X2=0
+ $Y2=0
cc_572 N_RESET_B_c_608_n N_A_1518_203#_M1015_g 0.00713109f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_573 N_RESET_B_c_611_n N_A_1518_203#_M1015_g 0.00231702f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_574 N_RESET_B_c_614_n N_A_1518_203#_M1015_g 0.0181717f $X=8.18 $Y=2.09 $X2=0
+ $Y2=0
cc_575 N_RESET_B_c_615_n N_A_1518_203#_M1015_g 0.00228452f $X=8.18 $Y=2.09 $X2=0
+ $Y2=0
cc_576 N_RESET_B_M1000_g N_A_1518_203#_M1013_g 0.0166359f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_577 N_RESET_B_M1000_g N_A_1518_203#_c_1112_n 0.0133984f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_578 N_RESET_B_M1000_g N_A_1518_203#_c_1113_n 0.0149634f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_579 N_RESET_B_M1000_g N_A_1518_203#_c_1114_n 0.00216035f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_580 N_RESET_B_M1000_g N_A_1518_203#_c_1123_n 0.00169886f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_581 N_RESET_B_c_611_n N_A_1518_203#_c_1123_n 4.76192e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_582 N_RESET_B_c_614_n N_A_1518_203#_c_1123_n 6.9451e-19 $X=8.18 $Y=2.09 $X2=0
+ $Y2=0
cc_583 N_RESET_B_c_615_n N_A_1518_203#_c_1123_n 0.00873148f $X=8.18 $Y=2.09
+ $X2=0 $Y2=0
cc_584 N_RESET_B_M1000_g N_A_1518_203#_c_1116_n 0.00118187f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_585 N_RESET_B_c_608_n N_A_1518_203#_c_1116_n 3.17521e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_586 N_RESET_B_M1000_g N_A_1518_203#_c_1117_n 0.021263f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_587 N_RESET_B_M1020_g N_A_1518_203#_c_1125_n 0.00713508f $X=8.26 $Y=2.675
+ $X2=0 $Y2=0
cc_588 N_RESET_B_c_615_n N_A_1518_203#_c_1125_n 0.0017001f $X=8.18 $Y=2.09 $X2=0
+ $Y2=0
cc_589 N_RESET_B_c_611_n N_A_1518_203#_c_1126_n 5.01506e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_590 N_RESET_B_c_614_n N_A_1518_203#_c_1126_n 0.00535994f $X=8.18 $Y=2.09
+ $X2=0 $Y2=0
cc_591 N_RESET_B_c_615_n N_A_1518_203#_c_1126_n 0.0175397f $X=8.18 $Y=2.09 $X2=0
+ $Y2=0
cc_592 N_RESET_B_c_608_n N_A_1266_74#_M1004_d 0.00197859f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_593 N_RESET_B_M1000_g N_A_1266_74#_M1017_g 0.0757442f $X=8.205 $Y=0.615 $X2=0
+ $Y2=0
cc_594 N_RESET_B_M1000_g N_A_1266_74#_M1024_g 0.00953304f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_595 N_RESET_B_c_614_n N_A_1266_74#_M1024_g 0.0313246f $X=8.18 $Y=2.09 $X2=0
+ $Y2=0
cc_596 N_RESET_B_c_615_n N_A_1266_74#_M1024_g 3.48207e-19 $X=8.18 $Y=2.09 $X2=0
+ $Y2=0
cc_597 N_RESET_B_M1000_g N_A_1266_74#_c_1227_n 0.00996674f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_598 N_RESET_B_c_608_n N_A_1266_74#_c_1244_n 0.0174694f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_599 N_RESET_B_c_608_n N_A_1266_74#_c_1267_n 0.0206114f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_600 N_RESET_B_M1000_g N_A_1266_74#_c_1245_n 0.00109662f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_601 N_RESET_B_M1020_g N_A_1266_74#_c_1245_n 8.85939e-19 $X=8.26 $Y=2.675
+ $X2=0 $Y2=0
cc_602 N_RESET_B_c_608_n N_A_1266_74#_c_1245_n 0.0211228f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_603 N_RESET_B_c_611_n N_A_1266_74#_c_1245_n 0.00228452f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_604 N_RESET_B_c_614_n N_A_1266_74#_c_1245_n 2.85076e-19 $X=8.18 $Y=2.09 $X2=0
+ $Y2=0
cc_605 N_RESET_B_c_615_n N_A_1266_74#_c_1245_n 0.0236542f $X=8.18 $Y=2.09 $X2=0
+ $Y2=0
cc_606 N_RESET_B_M1000_g N_A_1266_74#_c_1235_n 0.011972f $X=8.205 $Y=0.615 $X2=0
+ $Y2=0
cc_607 N_RESET_B_c_608_n N_A_1266_74#_c_1235_n 0.00476106f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_608 N_RESET_B_c_611_n N_A_1266_74#_c_1235_n 0.00823149f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_609 N_RESET_B_c_614_n N_A_1266_74#_c_1235_n 0.00136037f $X=8.18 $Y=2.09 $X2=0
+ $Y2=0
cc_610 N_RESET_B_c_615_n N_A_1266_74#_c_1235_n 0.02904f $X=8.18 $Y=2.09 $X2=0
+ $Y2=0
cc_611 N_RESET_B_c_608_n N_A_1266_74#_c_1237_n 0.00594354f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_612 N_RESET_B_M1000_g N_A_1266_74#_c_1238_n 0.00110907f $X=8.205 $Y=0.615
+ $X2=0 $Y2=0
cc_613 N_RESET_B_c_606_n N_VPWR_M1021_d 0.00508462f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_614 N_RESET_B_M1019_g N_VPWR_c_1434_n 0.0086413f $X=0.945 $Y=2.825 $X2=0
+ $Y2=0
cc_615 N_RESET_B_c_602_n N_VPWR_c_1436_n 0.00366918f $X=4.86 $Y=2.275 $X2=0
+ $Y2=0
cc_616 N_RESET_B_c_602_n N_VPWR_c_1438_n 0.0104488f $X=4.86 $Y=2.275 $X2=0 $Y2=0
cc_617 N_RESET_B_c_595_n N_VPWR_c_1438_n 0.00126145f $X=4.875 $Y=1.795 $X2=0
+ $Y2=0
cc_618 N_RESET_B_c_608_n N_VPWR_c_1438_n 0.0322565f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_619 N_RESET_B_c_609_n N_VPWR_c_1438_n 5.51604e-19 $X=5.185 $Y=2.035 $X2=0
+ $Y2=0
cc_620 N_RESET_B_c_610_n N_VPWR_c_1438_n 0.023147f $X=5.04 $Y=2.035 $X2=0 $Y2=0
cc_621 N_RESET_B_M1020_g N_VPWR_c_1439_n 0.00621399f $X=8.26 $Y=2.675 $X2=0
+ $Y2=0
cc_622 N_RESET_B_c_611_n N_VPWR_c_1439_n 0.00171912f $X=7.92 $Y=2.035 $X2=0
+ $Y2=0
cc_623 N_RESET_B_c_614_n N_VPWR_c_1439_n 0.00275991f $X=8.18 $Y=2.09 $X2=0 $Y2=0
cc_624 N_RESET_B_c_615_n N_VPWR_c_1439_n 0.0244512f $X=8.18 $Y=2.09 $X2=0 $Y2=0
cc_625 N_RESET_B_M1020_g N_VPWR_c_1440_n 0.00601158f $X=8.26 $Y=2.675 $X2=0
+ $Y2=0
cc_626 N_RESET_B_M1019_g N_VPWR_c_1444_n 0.00386446f $X=0.945 $Y=2.825 $X2=0
+ $Y2=0
cc_627 N_RESET_B_M1019_g N_VPWR_c_1431_n 0.00480274f $X=0.945 $Y=2.825 $X2=0
+ $Y2=0
cc_628 N_RESET_B_c_602_n N_VPWR_c_1431_n 0.00112687f $X=4.86 $Y=2.275 $X2=0
+ $Y2=0
cc_629 N_RESET_B_M1020_g N_VPWR_c_1431_n 0.00626544f $X=8.26 $Y=2.675 $X2=0
+ $Y2=0
cc_630 N_RESET_B_M1009_g N_A_30_78#_c_1568_n 0.00433444f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_631 N_RESET_B_M1009_g N_A_30_78#_c_1569_n 0.0089809f $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_632 N_RESET_B_c_591_n N_A_30_78#_c_1569_n 0.0116119f $X=1.072 $Y=1.893 $X2=0
+ $Y2=0
cc_633 N_RESET_B_M1019_g N_A_30_78#_c_1569_n 0.00621241f $X=0.945 $Y=2.825 $X2=0
+ $Y2=0
cc_634 N_RESET_B_c_607_n N_A_30_78#_c_1569_n 0.00172785f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_635 N_RESET_B_c_598_n N_A_30_78#_c_1569_n 0.00558005f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_636 N_RESET_B_c_599_n N_A_30_78#_c_1569_n 0.069302f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_637 N_RESET_B_c_613_n N_A_30_78#_c_1569_n 0.00614539f $X=1.155 $Y=1.975 $X2=0
+ $Y2=0
cc_638 N_RESET_B_M1019_g N_A_30_78#_c_1576_n 0.0161123f $X=0.945 $Y=2.825 $X2=0
+ $Y2=0
cc_639 N_RESET_B_c_606_n N_A_30_78#_c_1576_n 0.0292189f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_640 N_RESET_B_c_607_n N_A_30_78#_c_1576_n 0.00844426f $X=1.345 $Y=2.035 $X2=0
+ $Y2=0
cc_641 N_RESET_B_c_599_n N_A_30_78#_c_1576_n 0.00915778f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_642 N_RESET_B_c_613_n N_A_30_78#_c_1576_n 0.00253837f $X=1.155 $Y=1.975 $X2=0
+ $Y2=0
cc_643 N_RESET_B_c_606_n N_A_30_78#_c_1577_n 0.0107558f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_644 N_RESET_B_c_606_n N_A_30_78#_c_1571_n 0.0129345f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_645 N_RESET_B_M1009_g N_A_30_78#_c_1572_n 9.29579e-19 $X=0.9 $Y=0.6 $X2=0
+ $Y2=0
cc_646 N_RESET_B_M1019_g N_A_30_78#_c_1579_n 0.0058061f $X=0.945 $Y=2.825 $X2=0
+ $Y2=0
cc_647 N_RESET_B_c_606_n N_A_30_78#_c_1580_n 0.00767864f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_648 N_RESET_B_c_606_n N_A_30_78#_c_1573_n 0.005403f $X=4.895 $Y=2.035 $X2=0
+ $Y2=0
cc_649 N_RESET_B_M1009_g N_VGND_c_1712_n 0.00257803f $X=0.9 $Y=0.6 $X2=0 $Y2=0
cc_650 N_RESET_B_c_592_n N_VGND_c_1712_n 0.0200565f $X=4.71 $Y=0.18 $X2=0 $Y2=0
cc_651 N_RESET_B_c_598_n N_VGND_c_1712_n 0.00181416f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_652 N_RESET_B_c_599_n N_VGND_c_1712_n 0.0144384f $X=1.155 $Y=1.295 $X2=0
+ $Y2=0
cc_653 N_RESET_B_c_592_n N_VGND_c_1713_n 0.0257653f $X=4.71 $Y=0.18 $X2=0 $Y2=0
cc_654 N_RESET_B_M1000_g N_VGND_c_1714_n 0.0058325f $X=8.205 $Y=0.615 $X2=0
+ $Y2=0
cc_655 N_RESET_B_c_593_n N_VGND_c_1718_n 0.00764766f $X=0.975 $Y=0.18 $X2=0
+ $Y2=0
cc_656 N_RESET_B_c_592_n N_VGND_c_1720_n 0.0223671f $X=4.71 $Y=0.18 $X2=0 $Y2=0
cc_657 N_RESET_B_c_592_n N_VGND_c_1721_n 0.0625127f $X=4.71 $Y=0.18 $X2=0 $Y2=0
cc_658 N_RESET_B_M1000_g N_VGND_c_1723_n 0.00552345f $X=8.205 $Y=0.615 $X2=0
+ $Y2=0
cc_659 N_RESET_B_c_592_n N_VGND_c_1728_n 0.0926626f $X=4.71 $Y=0.18 $X2=0 $Y2=0
cc_660 N_RESET_B_c_593_n N_VGND_c_1728_n 0.0105042f $X=0.975 $Y=0.18 $X2=0 $Y2=0
cc_661 N_RESET_B_M1000_g N_VGND_c_1728_n 0.00534666f $X=8.205 $Y=0.615 $X2=0
+ $Y2=0
cc_662 N_A_701_463#_c_814_n N_A_299_387#_c_947_n 0.00349469f $X=3.935 $Y=2.64
+ $X2=0 $Y2=0
cc_663 N_A_701_463#_c_810_n N_A_299_387#_M1007_g 8.00721e-19 $X=4.02 $Y=0.812
+ $X2=0 $Y2=0
cc_664 N_A_701_463#_c_811_n N_A_299_387#_M1007_g 0.0011886f $X=4.075 $Y=2.36
+ $X2=0 $Y2=0
cc_665 N_A_701_463#_c_814_n N_A_299_387#_M1022_g 0.00916834f $X=3.935 $Y=2.64
+ $X2=0 $Y2=0
cc_666 N_A_701_463#_c_817_n N_A_299_387#_M1022_g 0.00822981f $X=4.075 $Y=2.46
+ $X2=0 $Y2=0
cc_667 N_A_701_463#_c_811_n N_A_299_387#_M1022_g 0.00303502f $X=4.075 $Y=2.36
+ $X2=0 $Y2=0
cc_668 N_A_701_463#_M1029_g N_A_299_387#_c_951_n 0.0124167f $X=5.88 $Y=2.235
+ $X2=0 $Y2=0
cc_669 N_A_701_463#_c_839_n N_A_299_387#_c_951_n 0.00124604f $X=4.615 $Y=2.46
+ $X2=0 $Y2=0
cc_670 N_A_701_463#_c_817_n N_A_299_387#_c_951_n 0.00253247f $X=4.075 $Y=2.46
+ $X2=0 $Y2=0
cc_671 N_A_701_463#_c_819_n N_A_299_387#_c_951_n 0.00625565f $X=4.7 $Y=2.5 $X2=0
+ $Y2=0
cc_672 N_A_701_463#_M1029_g N_A_299_387#_c_939_n 0.0182076f $X=5.88 $Y=2.235
+ $X2=0 $Y2=0
cc_673 N_A_701_463#_c_839_n N_VPWR_M1008_d 0.00477669f $X=4.615 $Y=2.46 $X2=0
+ $Y2=0
cc_674 N_A_701_463#_c_819_n N_VPWR_M1008_d 0.0014715f $X=4.7 $Y=2.5 $X2=0 $Y2=0
cc_675 N_A_701_463#_c_839_n N_VPWR_c_1436_n 0.0167043f $X=4.615 $Y=2.46 $X2=0
+ $Y2=0
cc_676 N_A_701_463#_c_817_n N_VPWR_c_1436_n 0.00114764f $X=4.075 $Y=2.46 $X2=0
+ $Y2=0
cc_677 N_A_701_463#_c_819_n N_VPWR_c_1436_n 0.00841104f $X=4.7 $Y=2.5 $X2=0
+ $Y2=0
cc_678 N_A_701_463#_c_819_n N_VPWR_c_1437_n 0.00488601f $X=4.7 $Y=2.5 $X2=0
+ $Y2=0
cc_679 N_A_701_463#_M1029_g N_VPWR_c_1438_n 0.0156464f $X=5.88 $Y=2.235 $X2=0
+ $Y2=0
cc_680 N_A_701_463#_c_808_n N_VPWR_c_1438_n 0.0132253f $X=5.485 $Y=1.41 $X2=0
+ $Y2=0
cc_681 N_A_701_463#_c_809_n N_VPWR_c_1438_n 0.00726322f $X=5.485 $Y=1.41 $X2=0
+ $Y2=0
cc_682 N_A_701_463#_c_819_n N_VPWR_c_1438_n 0.0252145f $X=4.7 $Y=2.5 $X2=0 $Y2=0
cc_683 N_A_701_463#_c_814_n N_VPWR_c_1446_n 0.0093859f $X=3.935 $Y=2.64 $X2=0
+ $Y2=0
cc_684 N_A_701_463#_c_817_n N_VPWR_c_1446_n 0.00615345f $X=4.075 $Y=2.46 $X2=0
+ $Y2=0
cc_685 N_A_701_463#_M1029_g N_VPWR_c_1431_n 0.00100812f $X=5.88 $Y=2.235 $X2=0
+ $Y2=0
cc_686 N_A_701_463#_c_814_n N_VPWR_c_1431_n 0.0118816f $X=3.935 $Y=2.64 $X2=0
+ $Y2=0
cc_687 N_A_701_463#_c_839_n N_VPWR_c_1431_n 0.00626132f $X=4.615 $Y=2.46 $X2=0
+ $Y2=0
cc_688 N_A_701_463#_c_817_n N_VPWR_c_1431_n 0.0075359f $X=4.075 $Y=2.46 $X2=0
+ $Y2=0
cc_689 N_A_701_463#_c_819_n N_VPWR_c_1431_n 0.015479f $X=4.7 $Y=2.5 $X2=0 $Y2=0
cc_690 N_A_701_463#_c_810_n N_A_30_78#_c_1570_n 0.0200654f $X=4.02 $Y=0.812
+ $X2=0 $Y2=0
cc_691 N_A_701_463#_c_811_n N_A_30_78#_c_1570_n 0.00462959f $X=4.075 $Y=2.36
+ $X2=0 $Y2=0
cc_692 N_A_701_463#_M1014_d N_A_30_78#_c_1577_n 0.00176212f $X=3.505 $Y=2.315
+ $X2=0 $Y2=0
cc_693 N_A_701_463#_c_814_n N_A_30_78#_c_1577_n 0.014029f $X=3.935 $Y=2.64 $X2=0
+ $Y2=0
cc_694 N_A_701_463#_c_811_n N_A_30_78#_c_1577_n 0.0117396f $X=4.075 $Y=2.36
+ $X2=0 $Y2=0
cc_695 N_A_701_463#_c_811_n N_A_30_78#_c_1571_n 0.05859f $X=4.075 $Y=2.36 $X2=0
+ $Y2=0
cc_696 N_A_701_463#_c_814_n N_A_30_78#_c_1580_n 0.00983037f $X=3.935 $Y=2.64
+ $X2=0 $Y2=0
cc_697 N_A_701_463#_c_811_n N_A_30_78#_c_1580_n 0.002121f $X=4.075 $Y=2.36 $X2=0
+ $Y2=0
cc_698 N_A_701_463#_c_810_n N_A_30_78#_c_1573_n 0.00744272f $X=4.02 $Y=0.812
+ $X2=0 $Y2=0
cc_699 N_A_701_463#_c_811_n N_A_30_78#_c_1573_n 0.0139602f $X=4.075 $Y=2.36
+ $X2=0 $Y2=0
cc_700 N_A_701_463#_c_811_n A_791_463# 5.2133e-19 $X=4.075 $Y=2.36 $X2=-0.19
+ $Y2=-0.245
cc_701 N_A_701_463#_M1031_g N_VGND_c_1721_n 0.00178007f $X=5.44 $Y=0.74 $X2=0
+ $Y2=0
cc_702 N_A_701_463#_M1031_g N_VGND_c_1722_n 0.00309023f $X=5.44 $Y=0.74 $X2=0
+ $Y2=0
cc_703 N_A_701_463#_M1031_g N_VGND_c_1728_n 0.00390562f $X=5.44 $Y=0.74 $X2=0
+ $Y2=0
cc_704 N_A_299_387#_M1016_g N_A_1518_203#_M1013_g 0.0368892f $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_705 N_A_299_387#_M1016_g N_A_1518_203#_c_1112_n 0.0235039f $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_706 N_A_299_387#_M1016_g N_A_1518_203#_c_1116_n 3.81559e-19 $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_707 N_A_299_387#_M1016_g N_A_1518_203#_c_1117_n 0.0205557f $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_708 N_A_299_387#_c_939_n N_A_1266_74#_c_1233_n 2.47725e-19 $X=6.475 $Y=1.66
+ $X2=0 $Y2=0
cc_709 N_A_299_387#_M1004_g N_A_1266_74#_c_1244_n 0.00984585f $X=6.385 $Y=2.385
+ $X2=0 $Y2=0
cc_710 N_A_299_387#_c_938_n N_A_1266_74#_c_1244_n 0.00695316f $X=7.23 $Y=1.66
+ $X2=0 $Y2=0
cc_711 N_A_299_387#_M1016_g N_A_1266_74#_c_1234_n 0.00507341f $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_712 N_A_299_387#_c_938_n N_A_1266_74#_c_1245_n 3.51038e-19 $X=7.23 $Y=1.66
+ $X2=0 $Y2=0
cc_713 N_A_299_387#_M1016_g N_A_1266_74#_c_1236_n 0.00127921f $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_714 N_A_299_387#_c_938_n N_A_1266_74#_c_1237_n 0.00490084f $X=7.23 $Y=1.66
+ $X2=0 $Y2=0
cc_715 N_A_299_387#_c_939_n N_A_1266_74#_c_1237_n 0.00531722f $X=6.475 $Y=1.66
+ $X2=0 $Y2=0
cc_716 N_A_299_387#_M1016_g N_A_1266_74#_c_1237_n 2.86702e-19 $X=7.305 $Y=0.615
+ $X2=0 $Y2=0
cc_717 N_A_299_387#_M1025_g N_VPWR_c_1435_n 0.0107256f $X=2.375 $Y=2.495 $X2=0
+ $Y2=0
cc_718 N_A_299_387#_c_946_n N_VPWR_c_1435_n 0.00207208f $X=2.885 $Y=3.075 $X2=0
+ $Y2=0
cc_719 N_A_299_387#_c_948_n N_VPWR_c_1435_n 7.02368e-19 $X=2.96 $Y=3.15 $X2=0
+ $Y2=0
cc_720 N_A_299_387#_M1022_g N_VPWR_c_1436_n 0.00617059f $X=3.865 $Y=2.525 $X2=0
+ $Y2=0
cc_721 N_A_299_387#_c_951_n N_VPWR_c_1436_n 0.0250293f $X=6.295 $Y=3.15 $X2=0
+ $Y2=0
cc_722 N_A_299_387#_c_951_n N_VPWR_c_1437_n 0.0236268f $X=6.295 $Y=3.15 $X2=0
+ $Y2=0
cc_723 N_A_299_387#_c_951_n N_VPWR_c_1438_n 0.0257967f $X=6.295 $Y=3.15 $X2=0
+ $Y2=0
cc_724 N_A_299_387#_M1004_g N_VPWR_c_1438_n 0.00637792f $X=6.385 $Y=2.385 $X2=0
+ $Y2=0
cc_725 N_A_299_387#_M1025_g N_VPWR_c_1446_n 0.0040249f $X=2.375 $Y=2.495 $X2=0
+ $Y2=0
cc_726 N_A_299_387#_c_948_n N_VPWR_c_1446_n 0.0442898f $X=2.96 $Y=3.15 $X2=0
+ $Y2=0
cc_727 N_A_299_387#_c_951_n N_VPWR_c_1447_n 0.0207332f $X=6.295 $Y=3.15 $X2=0
+ $Y2=0
cc_728 N_A_299_387#_M1025_g N_VPWR_c_1431_n 0.00503418f $X=2.375 $Y=2.495 $X2=0
+ $Y2=0
cc_729 N_A_299_387#_c_947_n N_VPWR_c_1431_n 0.0231327f $X=3.775 $Y=3.15 $X2=0
+ $Y2=0
cc_730 N_A_299_387#_c_948_n N_VPWR_c_1431_n 0.0059101f $X=2.96 $Y=3.15 $X2=0
+ $Y2=0
cc_731 N_A_299_387#_c_951_n N_VPWR_c_1431_n 0.0651362f $X=6.295 $Y=3.15 $X2=0
+ $Y2=0
cc_732 N_A_299_387#_c_955_n N_VPWR_c_1431_n 0.00499121f $X=3.865 $Y=3.15 $X2=0
+ $Y2=0
cc_733 N_A_299_387#_c_941_n N_A_30_78#_c_1569_n 0.00414764f $X=1.695 $Y=0.715
+ $X2=0 $Y2=0
cc_734 N_A_299_387#_c_944_n N_A_30_78#_c_1569_n 0.00499576f $X=1.695 $Y=1.055
+ $X2=0 $Y2=0
cc_735 N_A_299_387#_c_958_n N_A_30_78#_c_1569_n 0.00418053f $X=1.62 $Y=2.1 $X2=0
+ $Y2=0
cc_736 N_A_299_387#_M1021_s N_A_30_78#_c_1576_n 0.00624686f $X=1.495 $Y=1.935
+ $X2=0 $Y2=0
cc_737 N_A_299_387#_M1025_g N_A_30_78#_c_1576_n 0.0146133f $X=2.375 $Y=2.495
+ $X2=0 $Y2=0
cc_738 N_A_299_387#_c_946_n N_A_30_78#_c_1576_n 0.0128192f $X=2.885 $Y=3.075
+ $X2=0 $Y2=0
cc_739 N_A_299_387#_c_958_n N_A_30_78#_c_1576_n 0.0234284f $X=1.62 $Y=2.1 $X2=0
+ $Y2=0
cc_740 N_A_299_387#_c_935_n N_A_30_78#_c_1570_n 0.00156397f $X=3.47 $Y=1.4 $X2=0
+ $Y2=0
cc_741 N_A_299_387#_M1007_g N_A_30_78#_c_1570_n 0.0116369f $X=3.545 $Y=0.9 $X2=0
+ $Y2=0
cc_742 N_A_299_387#_M1022_g N_A_30_78#_c_1577_n 0.00132842f $X=3.865 $Y=2.525
+ $X2=0 $Y2=0
cc_743 N_A_299_387#_c_935_n N_A_30_78#_c_1571_n 0.00406894f $X=3.47 $Y=1.4 $X2=0
+ $Y2=0
cc_744 N_A_299_387#_c_936_n N_A_30_78#_c_1571_n 0.00150989f $X=3.04 $Y=1.4 $X2=0
+ $Y2=0
cc_745 N_A_299_387#_c_946_n N_A_30_78#_c_1580_n 0.00884165f $X=2.885 $Y=3.075
+ $X2=0 $Y2=0
cc_746 N_A_299_387#_c_947_n N_A_30_78#_c_1580_n 0.0050544f $X=3.775 $Y=3.15
+ $X2=0 $Y2=0
cc_747 N_A_299_387#_c_935_n N_A_30_78#_c_1573_n 0.0102217f $X=3.47 $Y=1.4 $X2=0
+ $Y2=0
cc_748 N_A_299_387#_M1007_g N_A_30_78#_c_1573_n 0.010712f $X=3.545 $Y=0.9 $X2=0
+ $Y2=0
cc_749 N_A_299_387#_c_971_n N_VGND_M1023_d 0.00592101f $X=2.445 $Y=1.055 $X2=0
+ $Y2=0
cc_750 N_A_299_387#_c_941_n N_VGND_c_1712_n 0.0227757f $X=1.695 $Y=0.715 $X2=0
+ $Y2=0
cc_751 N_A_299_387#_c_934_n N_VGND_c_1713_n 0.00119784f $X=2.475 $Y=1.41 $X2=0
+ $Y2=0
cc_752 N_A_299_387#_c_941_n N_VGND_c_1713_n 0.00357823f $X=1.695 $Y=0.715 $X2=0
+ $Y2=0
cc_753 N_A_299_387#_c_971_n N_VGND_c_1713_n 0.0208278f $X=2.445 $Y=1.055 $X2=0
+ $Y2=0
cc_754 N_A_299_387#_M1016_g N_VGND_c_1714_n 5.78056e-19 $X=7.305 $Y=0.615 $X2=0
+ $Y2=0
cc_755 N_A_299_387#_c_941_n N_VGND_c_1720_n 0.0100123f $X=1.695 $Y=0.715 $X2=0
+ $Y2=0
cc_756 N_A_299_387#_M1016_g N_VGND_c_1722_n 9.33926e-19 $X=7.305 $Y=0.615 $X2=0
+ $Y2=0
cc_757 N_A_299_387#_c_934_n N_VGND_c_1728_n 9.39239e-19 $X=2.475 $Y=1.41 $X2=0
+ $Y2=0
cc_758 N_A_299_387#_c_941_n N_VGND_c_1728_n 0.0116439f $X=1.695 $Y=0.715 $X2=0
+ $Y2=0
cc_759 N_A_1518_203#_c_1113_n N_A_1266_74#_M1017_g 0.0107164f $X=8.615 $Y=1.1
+ $X2=0 $Y2=0
cc_760 N_A_1518_203#_c_1114_n N_A_1266_74#_M1017_g 0.0159617f $X=8.78 $Y=0.615
+ $X2=0 $Y2=0
cc_761 N_A_1518_203#_c_1115_n N_A_1266_74#_M1017_g 0.00301146f $X=9.105 $Y=1.855
+ $X2=0 $Y2=0
cc_762 N_A_1518_203#_c_1118_n N_A_1266_74#_M1017_g 0.00389282f $X=9.105 $Y=1.1
+ $X2=0 $Y2=0
cc_763 N_A_1518_203#_c_1122_n N_A_1266_74#_M1024_g 0.0108266f $X=9.02 $Y=1.94
+ $X2=0 $Y2=0
cc_764 N_A_1518_203#_c_1123_n N_A_1266_74#_M1024_g 0.00310966f $X=8.685 $Y=1.94
+ $X2=0 $Y2=0
cc_765 N_A_1518_203#_c_1115_n N_A_1266_74#_M1024_g 0.00343619f $X=9.105 $Y=1.855
+ $X2=0 $Y2=0
cc_766 N_A_1518_203#_c_1125_n N_A_1266_74#_M1024_g 0.00786363f $X=8.485 $Y=2.675
+ $X2=0 $Y2=0
cc_767 N_A_1518_203#_c_1126_n N_A_1266_74#_M1024_g 0.00961954f $X=8.502 $Y=2.445
+ $X2=0 $Y2=0
cc_768 N_A_1518_203#_c_1122_n N_A_1266_74#_c_1226_n 0.00354772f $X=9.02 $Y=1.94
+ $X2=0 $Y2=0
cc_769 N_A_1518_203#_c_1115_n N_A_1266_74#_c_1226_n 0.0103302f $X=9.105 $Y=1.855
+ $X2=0 $Y2=0
cc_770 N_A_1518_203#_c_1118_n N_A_1266_74#_c_1226_n 0.00508985f $X=9.105 $Y=1.1
+ $X2=0 $Y2=0
cc_771 N_A_1518_203#_c_1123_n N_A_1266_74#_c_1227_n 7.74206e-19 $X=8.685 $Y=1.94
+ $X2=0 $Y2=0
cc_772 N_A_1518_203#_c_1118_n N_A_1266_74#_c_1227_n 8.2291e-19 $X=9.105 $Y=1.1
+ $X2=0 $Y2=0
cc_773 N_A_1518_203#_c_1115_n N_A_1266_74#_c_1228_n 0.00511666f $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_774 N_A_1518_203#_c_1118_n N_A_1266_74#_c_1228_n 0.00147647f $X=9.105 $Y=1.1
+ $X2=0 $Y2=0
cc_775 N_A_1518_203#_c_1122_n N_A_1266_74#_M1011_g 0.00526703f $X=9.02 $Y=1.94
+ $X2=0 $Y2=0
cc_776 N_A_1518_203#_c_1115_n N_A_1266_74#_M1011_g 0.00358035f $X=9.105 $Y=1.855
+ $X2=0 $Y2=0
cc_777 N_A_1518_203#_c_1126_n N_A_1266_74#_M1011_g 9.41942e-19 $X=8.502 $Y=2.445
+ $X2=0 $Y2=0
cc_778 N_A_1518_203#_c_1114_n N_A_1266_74#_c_1230_n 2.88416e-19 $X=8.78 $Y=0.615
+ $X2=0 $Y2=0
cc_779 N_A_1518_203#_c_1118_n N_A_1266_74#_c_1230_n 0.00670166f $X=9.105 $Y=1.1
+ $X2=0 $Y2=0
cc_780 N_A_1518_203#_c_1114_n N_A_1266_74#_c_1231_n 0.00317724f $X=8.78 $Y=0.615
+ $X2=0 $Y2=0
cc_781 N_A_1518_203#_c_1115_n N_A_1266_74#_c_1232_n 0.00419613f $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_782 N_A_1518_203#_M1015_g N_A_1266_74#_c_1267_n 0.00803155f $X=7.685 $Y=2.675
+ $X2=0 $Y2=0
cc_783 N_A_1518_203#_c_1119_n N_A_1266_74#_c_1245_n 0.00331106f $X=7.685
+ $Y=1.835 $X2=0 $Y2=0
cc_784 N_A_1518_203#_M1015_g N_A_1266_74#_c_1245_n 0.01469f $X=7.685 $Y=2.675
+ $X2=0 $Y2=0
cc_785 N_A_1518_203#_c_1112_n N_A_1266_74#_c_1245_n 0.0015543f $X=7.685 $Y=1.745
+ $X2=0 $Y2=0
cc_786 N_A_1518_203#_c_1119_n N_A_1266_74#_c_1235_n 8.29273e-19 $X=7.685
+ $Y=1.835 $X2=0 $Y2=0
cc_787 N_A_1518_203#_c_1112_n N_A_1266_74#_c_1235_n 0.00762694f $X=7.685
+ $Y=1.745 $X2=0 $Y2=0
cc_788 N_A_1518_203#_c_1113_n N_A_1266_74#_c_1235_n 0.0272699f $X=8.615 $Y=1.1
+ $X2=0 $Y2=0
cc_789 N_A_1518_203#_c_1123_n N_A_1266_74#_c_1235_n 4.22281e-19 $X=8.685 $Y=1.94
+ $X2=0 $Y2=0
cc_790 N_A_1518_203#_c_1116_n N_A_1266_74#_c_1235_n 0.0204811f $X=7.755 $Y=1.1
+ $X2=0 $Y2=0
cc_791 N_A_1518_203#_c_1117_n N_A_1266_74#_c_1235_n 0.00111936f $X=7.755 $Y=1.18
+ $X2=0 $Y2=0
cc_792 N_A_1518_203#_c_1112_n N_A_1266_74#_c_1236_n 0.00211774f $X=7.685
+ $Y=1.745 $X2=0 $Y2=0
cc_793 N_A_1518_203#_c_1116_n N_A_1266_74#_c_1236_n 0.0034757f $X=7.755 $Y=1.1
+ $X2=0 $Y2=0
cc_794 N_A_1518_203#_c_1113_n N_A_1266_74#_c_1238_n 0.0242574f $X=8.615 $Y=1.1
+ $X2=0 $Y2=0
cc_795 N_A_1518_203#_c_1122_n N_A_1266_74#_c_1238_n 0.0118853f $X=9.02 $Y=1.94
+ $X2=0 $Y2=0
cc_796 N_A_1518_203#_c_1123_n N_A_1266_74#_c_1238_n 0.0136054f $X=8.685 $Y=1.94
+ $X2=0 $Y2=0
cc_797 N_A_1518_203#_c_1115_n N_A_1266_74#_c_1238_n 0.0235661f $X=9.105 $Y=1.855
+ $X2=0 $Y2=0
cc_798 N_A_1518_203#_c_1115_n N_A_1867_409#_c_1381_n 2.38456e-19 $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_799 N_A_1518_203#_c_1122_n N_A_1867_409#_c_1388_n 0.0122325f $X=9.02 $Y=1.94
+ $X2=0 $Y2=0
cc_800 N_A_1518_203#_c_1115_n N_A_1867_409#_c_1388_n 0.00900265f $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_801 N_A_1518_203#_c_1114_n N_A_1867_409#_c_1383_n 0.00478045f $X=8.78
+ $Y=0.615 $X2=0 $Y2=0
cc_802 N_A_1518_203#_c_1115_n N_A_1867_409#_c_1383_n 0.0077671f $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_803 N_A_1518_203#_c_1118_n N_A_1867_409#_c_1383_n 0.00665068f $X=9.105 $Y=1.1
+ $X2=0 $Y2=0
cc_804 N_A_1518_203#_c_1115_n N_A_1867_409#_c_1384_n 0.0234089f $X=9.105
+ $Y=1.855 $X2=0 $Y2=0
cc_805 N_A_1518_203#_M1015_g N_VPWR_c_1439_n 0.004218f $X=7.685 $Y=2.675 $X2=0
+ $Y2=0
cc_806 N_A_1518_203#_c_1125_n N_VPWR_c_1439_n 0.0178695f $X=8.485 $Y=2.675 $X2=0
+ $Y2=0
cc_807 N_A_1518_203#_c_1125_n N_VPWR_c_1440_n 0.0119999f $X=8.485 $Y=2.675 $X2=0
+ $Y2=0
cc_808 N_A_1518_203#_c_1122_n N_VPWR_c_1441_n 0.0258104f $X=9.02 $Y=1.94 $X2=0
+ $Y2=0
cc_809 N_A_1518_203#_c_1126_n N_VPWR_c_1441_n 0.0379498f $X=8.502 $Y=2.445 $X2=0
+ $Y2=0
cc_810 N_A_1518_203#_M1015_g N_VPWR_c_1447_n 0.00593406f $X=7.685 $Y=2.675 $X2=0
+ $Y2=0
cc_811 N_A_1518_203#_M1015_g N_VPWR_c_1431_n 0.00626544f $X=7.685 $Y=2.675 $X2=0
+ $Y2=0
cc_812 N_A_1518_203#_c_1125_n N_VPWR_c_1431_n 0.0125964f $X=8.485 $Y=2.675 $X2=0
+ $Y2=0
cc_813 N_A_1518_203#_M1013_g N_VGND_c_1714_n 0.0107187f $X=7.695 $Y=0.615 $X2=0
+ $Y2=0
cc_814 N_A_1518_203#_c_1113_n N_VGND_c_1714_n 0.0130069f $X=8.615 $Y=1.1 $X2=0
+ $Y2=0
cc_815 N_A_1518_203#_c_1114_n N_VGND_c_1714_n 0.00738736f $X=8.78 $Y=0.615 $X2=0
+ $Y2=0
cc_816 N_A_1518_203#_c_1116_n N_VGND_c_1714_n 0.0145528f $X=7.755 $Y=1.1 $X2=0
+ $Y2=0
cc_817 N_A_1518_203#_c_1117_n N_VGND_c_1714_n 0.0011793f $X=7.755 $Y=1.18 $X2=0
+ $Y2=0
cc_818 N_A_1518_203#_c_1114_n N_VGND_c_1715_n 0.0303742f $X=8.78 $Y=0.615 $X2=0
+ $Y2=0
cc_819 N_A_1518_203#_c_1118_n N_VGND_c_1715_n 0.00112954f $X=9.105 $Y=1.1 $X2=0
+ $Y2=0
cc_820 N_A_1518_203#_M1013_g N_VGND_c_1722_n 0.0045897f $X=7.695 $Y=0.615 $X2=0
+ $Y2=0
cc_821 N_A_1518_203#_c_1114_n N_VGND_c_1723_n 0.0126905f $X=8.78 $Y=0.615 $X2=0
+ $Y2=0
cc_822 N_A_1518_203#_M1013_g N_VGND_c_1728_n 0.0044912f $X=7.695 $Y=0.615 $X2=0
+ $Y2=0
cc_823 N_A_1518_203#_c_1114_n N_VGND_c_1728_n 0.0118012f $X=8.78 $Y=0.615 $X2=0
+ $Y2=0
cc_824 N_A_1266_74#_c_1229_n N_A_1867_409#_c_1381_n 0.00139534f $X=9.48 $Y=1.07
+ $X2=0 $Y2=0
cc_825 N_A_1266_74#_c_1232_n N_A_1867_409#_c_1381_n 0.0154815f $X=9.245 $Y=1.52
+ $X2=0 $Y2=0
cc_826 N_A_1266_74#_M1011_g N_A_1867_409#_c_1388_n 0.0116614f $X=9.245 $Y=2.465
+ $X2=0 $Y2=0
cc_827 N_A_1266_74#_c_1228_n N_A_1867_409#_c_1383_n 0.00400367f $X=9.23 $Y=1.355
+ $X2=0 $Y2=0
cc_828 N_A_1266_74#_c_1229_n N_A_1867_409#_c_1383_n 0.00708838f $X=9.48 $Y=1.07
+ $X2=0 $Y2=0
cc_829 N_A_1266_74#_c_1231_n N_A_1867_409#_c_1383_n 0.0140899f $X=9.555 $Y=0.995
+ $X2=0 $Y2=0
cc_830 N_A_1266_74#_c_1232_n N_A_1867_409#_c_1383_n 7.91947e-19 $X=9.245 $Y=1.52
+ $X2=0 $Y2=0
cc_831 N_A_1266_74#_c_1229_n N_A_1867_409#_c_1384_n 0.0079216f $X=9.48 $Y=1.07
+ $X2=0 $Y2=0
cc_832 N_A_1266_74#_c_1232_n N_A_1867_409#_c_1384_n 0.00324958f $X=9.245 $Y=1.52
+ $X2=0 $Y2=0
cc_833 N_A_1266_74#_c_1245_n N_VPWR_c_1439_n 0.0017733f $X=7.55 $Y=2.475 $X2=0
+ $Y2=0
cc_834 N_A_1266_74#_M1024_g N_VPWR_c_1440_n 0.00567808f $X=8.71 $Y=2.675 $X2=0
+ $Y2=0
cc_835 N_A_1266_74#_M1024_g N_VPWR_c_1441_n 0.00787004f $X=8.71 $Y=2.675 $X2=0
+ $Y2=0
cc_836 N_A_1266_74#_c_1226_n N_VPWR_c_1441_n 3.97376e-19 $X=9.155 $Y=1.52 $X2=0
+ $Y2=0
cc_837 N_A_1266_74#_M1011_g N_VPWR_c_1441_n 0.0145837f $X=9.245 $Y=2.465 $X2=0
+ $Y2=0
cc_838 N_A_1266_74#_c_1267_n N_VPWR_c_1447_n 0.0213217f $X=7.465 $Y=2.64 $X2=0
+ $Y2=0
cc_839 N_A_1266_74#_c_1363_p N_VPWR_c_1447_n 0.00361811f $X=6.65 $Y=2.64 $X2=0
+ $Y2=0
cc_840 N_A_1266_74#_M1011_g N_VPWR_c_1448_n 0.00522765f $X=9.245 $Y=2.465 $X2=0
+ $Y2=0
cc_841 N_A_1266_74#_M1024_g N_VPWR_c_1431_n 0.00626544f $X=8.71 $Y=2.675 $X2=0
+ $Y2=0
cc_842 N_A_1266_74#_M1011_g N_VPWR_c_1431_n 0.005256f $X=9.245 $Y=2.465 $X2=0
+ $Y2=0
cc_843 N_A_1266_74#_c_1267_n N_VPWR_c_1431_n 0.0312985f $X=7.465 $Y=2.64 $X2=0
+ $Y2=0
cc_844 N_A_1266_74#_c_1363_p N_VPWR_c_1431_n 0.00557315f $X=6.65 $Y=2.64 $X2=0
+ $Y2=0
cc_845 N_A_1266_74#_c_1267_n A_1471_493# 0.00285115f $X=7.465 $Y=2.64 $X2=-0.19
+ $Y2=-0.245
cc_846 N_A_1266_74#_c_1231_n N_Q_c_1683_n 0.00112501f $X=9.555 $Y=0.995 $X2=0
+ $Y2=0
cc_847 N_A_1266_74#_c_1229_n N_Q_c_1684_n 0.00112501f $X=9.48 $Y=1.07 $X2=0
+ $Y2=0
cc_848 N_A_1266_74#_M1011_g Q 0.00350879f $X=9.245 $Y=2.465 $X2=0 $Y2=0
cc_849 N_A_1266_74#_M1017_g N_VGND_c_1715_n 0.00359522f $X=8.565 $Y=0.615 $X2=0
+ $Y2=0
cc_850 N_A_1266_74#_c_1230_n N_VGND_c_1715_n 0.0104251f $X=9.305 $Y=1.07 $X2=0
+ $Y2=0
cc_851 N_A_1266_74#_c_1231_n N_VGND_c_1715_n 0.0065091f $X=9.555 $Y=0.995 $X2=0
+ $Y2=0
cc_852 N_A_1266_74#_M1017_g N_VGND_c_1723_n 0.00527282f $X=8.565 $Y=0.615 $X2=0
+ $Y2=0
cc_853 N_A_1266_74#_c_1231_n N_VGND_c_1724_n 0.00434272f $X=9.555 $Y=0.995 $X2=0
+ $Y2=0
cc_854 N_A_1266_74#_M1017_g N_VGND_c_1728_n 0.00534666f $X=8.565 $Y=0.615 $X2=0
+ $Y2=0
cc_855 N_A_1266_74#_c_1231_n N_VGND_c_1728_n 0.00830282f $X=9.555 $Y=0.995 $X2=0
+ $Y2=0
cc_856 N_A_1867_409#_c_1388_n N_VPWR_c_1441_n 0.0240288f $X=9.47 $Y=2.19 $X2=0
+ $Y2=0
cc_857 N_A_1867_409#_c_1385_n N_VPWR_c_1443_n 0.023669f $X=10.53 $Y=1.715 $X2=0
+ $Y2=0
cc_858 N_A_1867_409#_c_1385_n N_VPWR_c_1448_n 0.00475445f $X=10.53 $Y=1.715
+ $X2=0 $Y2=0
cc_859 N_A_1867_409#_c_1388_n N_VPWR_c_1448_n 0.00575213f $X=9.47 $Y=2.19 $X2=0
+ $Y2=0
cc_860 N_A_1867_409#_c_1385_n N_VPWR_c_1431_n 0.00943794f $X=10.53 $Y=1.715
+ $X2=0 $Y2=0
cc_861 N_A_1867_409#_c_1388_n N_VPWR_c_1431_n 0.00591657f $X=9.47 $Y=2.19 $X2=0
+ $Y2=0
cc_862 N_A_1867_409#_M1003_g N_Q_c_1683_n 0.00853833f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_863 N_A_1867_409#_c_1383_n N_Q_c_1683_n 0.0694074f $X=9.77 $Y=0.645 $X2=0
+ $Y2=0
cc_864 N_A_1867_409#_M1003_g N_Q_c_1684_n 0.00343176f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_865 N_A_1867_409#_c_1381_n N_Q_c_1684_n 0.00191508f $X=10.44 $Y=1.55 $X2=0
+ $Y2=0
cc_866 N_A_1867_409#_c_1381_n Q 0.0150903f $X=10.44 $Y=1.55 $X2=0 $Y2=0
cc_867 N_A_1867_409#_c_1388_n Q 0.0848079f $X=9.47 $Y=2.19 $X2=0 $Y2=0
cc_868 N_A_1867_409#_c_1384_n Q 0.017588f $X=9.77 $Y=1.55 $X2=0 $Y2=0
cc_869 N_A_1867_409#_c_1385_n N_Q_c_1685_n 0.00584027f $X=10.53 $Y=1.715 $X2=0
+ $Y2=0
cc_870 N_A_1867_409#_M1003_g N_Q_c_1685_n 0.0104864f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_871 N_A_1867_409#_c_1381_n N_Q_c_1685_n 0.0395686f $X=10.44 $Y=1.55 $X2=0
+ $Y2=0
cc_872 N_A_1867_409#_c_1388_n N_Q_c_1685_n 0.00535008f $X=9.47 $Y=2.19 $X2=0
+ $Y2=0
cc_873 N_A_1867_409#_c_1384_n N_Q_c_1685_n 0.0198451f $X=9.77 $Y=1.55 $X2=0
+ $Y2=0
cc_874 N_A_1867_409#_c_1383_n N_VGND_c_1715_n 0.0184694f $X=9.77 $Y=0.645 $X2=0
+ $Y2=0
cc_875 N_A_1867_409#_c_1384_n N_VGND_c_1715_n 0.00144181f $X=9.77 $Y=1.55 $X2=0
+ $Y2=0
cc_876 N_A_1867_409#_M1003_g N_VGND_c_1717_n 0.00647412f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_877 N_A_1867_409#_M1003_g N_VGND_c_1724_n 0.00434272f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_878 N_A_1867_409#_c_1383_n N_VGND_c_1724_n 0.0145639f $X=9.77 $Y=0.645 $X2=0
+ $Y2=0
cc_879 N_A_1867_409#_M1003_g N_VGND_c_1728_n 0.00828941f $X=10.545 $Y=0.74 $X2=0
+ $Y2=0
cc_880 N_A_1867_409#_c_1383_n N_VGND_c_1728_n 0.0119984f $X=9.77 $Y=0.645 $X2=0
+ $Y2=0
cc_881 N_VPWR_c_1444_n N_A_30_78#_c_1574_n 0.0144625f $X=1.005 $Y=3.33 $X2=0
+ $Y2=0
cc_882 N_VPWR_c_1431_n N_A_30_78#_c_1574_n 0.011411f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_883 N_VPWR_M1021_d N_A_30_78#_c_1576_n 0.00445472f $X=2.015 $Y=1.935 $X2=0
+ $Y2=0
cc_884 N_VPWR_c_1434_n N_A_30_78#_c_1576_n 0.0232756f $X=1.17 $Y=2.89 $X2=0
+ $Y2=0
cc_885 N_VPWR_c_1435_n N_A_30_78#_c_1576_n 0.0163245f $X=2.15 $Y=2.87 $X2=0
+ $Y2=0
cc_886 N_VPWR_c_1444_n N_A_30_78#_c_1576_n 0.00162466f $X=1.005 $Y=3.33 $X2=0
+ $Y2=0
cc_887 N_VPWR_c_1445_n N_A_30_78#_c_1576_n 0.00920625f $X=1.985 $Y=3.33 $X2=0
+ $Y2=0
cc_888 N_VPWR_c_1446_n N_A_30_78#_c_1576_n 0.00984423f $X=4.39 $Y=3.33 $X2=0
+ $Y2=0
cc_889 N_VPWR_c_1431_n N_A_30_78#_c_1576_n 0.0392722f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_890 N_VPWR_c_1444_n N_A_30_78#_c_1579_n 5.98759e-19 $X=1.005 $Y=3.33 $X2=0
+ $Y2=0
cc_891 N_VPWR_c_1431_n N_A_30_78#_c_1579_n 0.00124618f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_892 N_VPWR_c_1446_n N_A_30_78#_c_1580_n 0.00627421f $X=4.39 $Y=3.33 $X2=0
+ $Y2=0
cc_893 N_VPWR_c_1431_n N_A_30_78#_c_1580_n 0.00762703f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_894 N_VPWR_c_1441_n Q 0.00265691f $X=9.02 $Y=2.36 $X2=0 $Y2=0
cc_895 N_VPWR_c_1448_n Q 0.0311454f $X=10.595 $Y=3.33 $X2=0 $Y2=0
cc_896 N_VPWR_c_1431_n Q 0.0257795f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_897 N_VPWR_c_1443_n N_Q_c_1685_n 0.0451739f $X=10.76 $Y=1.985 $X2=0 $Y2=0
cc_898 N_A_30_78#_c_1568_n A_117_78# 0.00231141f $X=0.685 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_899 N_A_30_78#_c_1568_n N_VGND_c_1712_n 0.00719261f $X=0.685 $Y=0.745 $X2=0
+ $Y2=0
cc_900 N_A_30_78#_c_1572_n N_VGND_c_1712_n 0.00436551f $X=0.295 $Y=0.6 $X2=0
+ $Y2=0
cc_901 N_A_30_78#_c_1568_n N_VGND_c_1718_n 0.00570266f $X=0.685 $Y=0.745 $X2=0
+ $Y2=0
cc_902 N_A_30_78#_c_1572_n N_VGND_c_1718_n 0.0131067f $X=0.295 $Y=0.6 $X2=0
+ $Y2=0
cc_903 N_A_30_78#_c_1568_n N_VGND_c_1728_n 0.0110739f $X=0.685 $Y=0.745 $X2=0
+ $Y2=0
cc_904 N_A_30_78#_c_1572_n N_VGND_c_1728_n 0.0117869f $X=0.295 $Y=0.6 $X2=0
+ $Y2=0
cc_905 N_Q_c_1683_n N_VGND_c_1717_n 0.0293763f $X=10.33 $Y=0.515 $X2=0 $Y2=0
cc_906 N_Q_c_1683_n N_VGND_c_1724_n 0.0145639f $X=10.33 $Y=0.515 $X2=0 $Y2=0
cc_907 N_Q_c_1683_n N_VGND_c_1728_n 0.0119984f $X=10.33 $Y=0.515 $X2=0 $Y2=0

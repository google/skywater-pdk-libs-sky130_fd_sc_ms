* File: sky130_fd_sc_ms__dfsbp_1.spice
* Created: Wed Sep  2 12:03:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dfsbp_1.pex.spice"
.subckt sky130_fd_sc_ms__dfsbp_1  VNB VPB D CLK SET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* D	D
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_D_M1003_g N_A_27_80#_M1003_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1032 N_VGND_M1032_d N_CLK_M1032_g N_A_225_74#_M1032_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1013 N_A_398_74#_M1013_d N_A_225_74#_M1013_g N_VGND_M1032_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_A_596_81#_M1004_d N_A_225_74#_M1004_g N_A_27_80#_M1004_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1281 AS=0.1197 PD=1.03 PS=1.41 NRD=94.284 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1022 A_748_81# N_A_398_74#_M1022_g N_A_596_81#_M1004_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.1281 PD=0.66 PS=1.03 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_779_380#_M1006_g A_748_81# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 A_1061_74# N_A_596_81#_M1015_g N_A_779_380#_M1015_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.1113 PD=0.66 PS=1.37 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.9 A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_SET_B_M1026_g A_1061_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.102226 AS=0.0504 PD=0.87566 PS=0.66 NRD=53.568 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1000 A_1262_74# N_A_596_81#_M1000_g N_VGND_M1026_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1088 AS=0.155774 PD=0.98 PS=1.33434 NRD=21.552 NRS=0 M=1 R=4.26667
+ SA=75000.9 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1018 N_A_1358_377#_M1018_d N_A_398_74#_M1018_g A_1262_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.129147 AS=0.1088 PD=1.20755 PS=0.98 NRD=0 NRS=21.552 M=1 R=4.26667
+ SA=75001.3 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1031 A_1462_74# N_A_225_74#_M1031_g N_A_1358_377#_M1018_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0847528 PD=0.66 PS=0.792453 NRD=18.564 NRS=24.276 M=1
+ R=2.8 SA=75002.2 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1028 A_1540_74# N_A_1510_48#_M1028_g A_1462_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75002.6
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_SET_B_M1024_g A_1540_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1491 AS=0.0504 PD=1.13 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75003
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1011 N_A_1510_48#_M1011_d N_A_1358_377#_M1011_g N_VGND_M1024_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1197 AS=0.1491 PD=1.41 PS=1.13 NRD=0 NRS=19.992 M=1 R=2.8
+ SA=75003.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_Q_N_M1008_d N_A_1358_377#_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.2627 PD=2.05 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1025 N_VGND_M1025_d N_A_1358_377#_M1025_g N_A_2113_74#_M1025_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.129591 AS=0.15675 PD=0.997674 PS=1.67 NRD=17.988 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1021 N_Q_M1021_d N_A_2113_74#_M1021_g N_VGND_M1025_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1023 N_VPWR_M1023_d N_D_M1023_g N_A_27_80#_M1023_s VPB PSHORT L=0.18 W=0.42
+ AD=0.1176 AS=0.1176 PD=1.4 PS=1.4 NRD=0 NRS=0 M=1 R=2.33333 SA=90000.2
+ SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1012 N_VPWR_M1012_d N_CLK_M1012_g N_A_225_74#_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1019 N_A_398_74#_M1019_d N_A_225_74#_M1019_g N_VPWR_M1012_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1009 N_A_596_81#_M1009_d N_A_398_74#_M1009_g N_A_27_80#_M1009_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0672 AS=0.1176 PD=0.74 PS=1.4 NRD=21.0987 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90004.4 A=0.0756 P=1.2 MULT=1
MM1007 A_731_463# N_A_225_74#_M1007_g N_A_596_81#_M1009_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0672 PD=0.66 PS=0.74 NRD=30.4759 NRS=0 M=1 R=2.33333
+ SA=90000.7 SB=90003.9 A=0.0756 P=1.2 MULT=1
MM1020 N_VPWR_M1020_d N_A_779_380#_M1020_g A_731_463# VPB PSHORT L=0.18 W=0.42
+ AD=0.15225 AS=0.0504 PD=1.145 PS=0.66 NRD=11.7215 NRS=30.4759 M=1 R=2.33333
+ SA=90001.1 SB=90003.5 A=0.0756 P=1.2 MULT=1
MM1029 N_A_779_380#_M1029_d N_A_596_81#_M1029_g N_VPWR_M1020_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0693 AS=0.15225 PD=0.75 PS=1.145 NRD=0 NRS=197 M=1 R=2.33333
+ SA=90002 SB=90002.6 A=0.0756 P=1.2 MULT=1
MM1016 N_VPWR_M1016_d N_SET_B_M1016_g N_A_779_380#_M1029_d VPB PSHORT L=0.18
+ W=0.42 AD=0.125335 AS=0.0693 PD=0.996761 PS=0.75 NRD=98.4803 NRS=25.7873 M=1
+ R=2.33333 SA=90002.5 SB=90002.1 A=0.0756 P=1.2 MULT=1
MM1001 A_1257_341# N_A_596_81#_M1001_g N_VPWR_M1016_d VPB PSHORT L=0.18 W=1
+ AD=0.17825 AS=0.298415 PD=1.505 PS=2.37324 NRD=24.2704 NRS=25.5903 M=1
+ R=5.55556 SA=90001.4 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1002 N_A_1358_377#_M1002_d N_A_225_74#_M1002_g A_1257_341# VPB PSHORT L=0.18
+ W=1 AD=0.295423 AS=0.17825 PD=2.40141 PS=1.505 NRD=0 NRS=24.2704 M=1 R=5.55556
+ SA=90001.8 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1005 A_1520_508# N_A_398_74#_M1005_g N_A_1358_377#_M1002_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.124077 PD=0.66 PS=1.00859 NRD=30.4759 NRS=0 M=1
+ R=2.33333 SA=90002.3 SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1010_d N_A_1510_48#_M1010_g A_1520_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.0567 AS=0.0504 PD=0.69 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.33333 SA=90002.7
+ SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1014 N_A_1358_377#_M1014_d N_SET_B_M1014_g N_VPWR_M1010_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1176 AS=0.0567 PD=1.4 PS=0.69 NRD=0 NRS=0 M=1 R=2.33333 SA=90003.1
+ SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1017 N_VPWR_M1017_d N_A_1358_377#_M1017_g N_A_1510_48#_M1017_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0849545 AS=0.1533 PD=0.788182 PS=1.57 NRD=14.0658
+ NRS=37.5088 M=1 R=2.33333 SA=90000.3 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1030 N_Q_N_M1030_d N_A_1358_377#_M1030_g N_VPWR_M1017_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.226545 PD=2.8 PS=2.10182 NRD=0 NRS=2.6201 M=1 R=6.22222
+ SA=90000.4 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1033 N_VPWR_M1033_d N_A_1358_377#_M1033_g N_A_2113_74#_M1033_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.147 AS=0.2352 PD=1.23857 PS=2.24 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1027 N_Q_M1027_d N_A_2113_74#_M1027_g N_VPWR_M1033_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.196 PD=2.8 PS=1.65143 NRD=0 NRS=8.7862 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX34_noxref VNB VPB NWDIODE A=23.4027 P=28.75
*
.include "sky130_fd_sc_ms__dfsbp_1.pxi.spice"
*
.ends
*
*

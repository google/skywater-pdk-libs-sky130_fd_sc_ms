* File: sky130_fd_sc_ms__dlrtn_2.spice
* Created: Fri Aug 28 17:27:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dlrtn_2.pex.spice"
.subckt sky130_fd_sc_ms__dlrtn_2  VNB VPB D GATE_N RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_D_M1017_g N_A_27_136#_M1017_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.171076 AS=0.15675 PD=1.27054 PS=1.67 NRD=55.86 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1001 N_A_232_98#_M1001_d N_GATE_N_M1001_g N_VGND_M1017_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2257 AS=0.230174 PD=2.09 PS=1.70946 NRD=0 NRS=41.52 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_232_98#_M1007_g N_A_373_82#_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.4514 AS=0.2294 PD=2.12348 PS=2.1 NRD=89.988 NRS=2.424 M=1
+ R=4.93333 SA=75000.2 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1016 A_697_74# N_A_27_136#_M1016_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.3904 PD=0.88 PS=1.83652 NRD=12.18 NRS=15.936 M=1 R=4.26667
+ SA=75001.4 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1014 N_A_673_392#_M1014_d N_A_232_98#_M1014_g A_697_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.115623 AS=0.0768 PD=1.16528 PS=0.88 NRD=8.436 NRS=12.18 M=1
+ R=4.26667 SA=75001.8 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1020 A_870_74# N_A_373_82#_M1020_g N_A_673_392#_M1014_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.05775 AS=0.0758774 PD=0.695 PS=0.764717 NRD=23.568 NRS=0 M=1 R=2.8
+ SA=75002.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1018_d N_A_913_406#_M1018_g A_870_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.05775 PD=1.41 PS=0.695 NRD=0 NRS=23.568 M=1 R=2.8 SA=75002.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_1153_74# N_A_673_392#_M1002_g N_A_913_406#_M1002_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.2 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_RESET_B_M1000_g A_1153_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.34225 AS=0.0888 PD=1.665 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333
+ SA=75000.6 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1004 N_Q_M1004_d N_A_913_406#_M1004_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.34225 PD=1.02 PS=1.665 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.7
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1013 N_Q_M1004_d N_A_913_406#_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.1
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1015 N_VPWR_M1015_d N_D_M1015_g N_A_27_136#_M1015_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1554 AS=0.2352 PD=1.21 PS=2.24 NRD=10.5395 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1011 N_A_232_98#_M1011_d N_GATE_N_M1011_g N_VPWR_M1015_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.1554 PD=2.24 PS=1.21 NRD=0 NRS=10.5395 M=1 R=4.66667
+ SA=90000.7 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1021 N_VPWR_M1021_d N_A_232_98#_M1021_g N_A_373_82#_M1021_s VPB PSHORT L=0.18
+ W=0.84 AD=0.223193 AS=0.2352 PD=1.50652 PS=2.24 NRD=49.4076 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90002.7 A=0.1512 P=2.04 MULT=1
MM1003 A_589_392# N_A_27_136#_M1003_g N_VPWR_M1021_d VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.265707 PD=1.24 PS=1.79348 NRD=12.7853 NRS=16.7253 M=1 R=5.55556
+ SA=90000.7 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1010 N_A_673_392#_M1010_d N_A_373_82#_M1010_g A_589_392# VPB PSHORT L=0.18 W=1
+ AD=0.222394 AS=0.12 PD=1.91549 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556
+ SA=90001.1 SB=90002 A=0.18 P=2.36 MULT=1
MM1012 A_781_504# N_A_232_98#_M1012_g N_A_673_392#_M1010_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1386 AS=0.0934056 PD=1.08 PS=0.804507 NRD=128.976 NRS=78.5045 M=1
+ R=2.33333 SA=90001.6 SB=90004 A=0.0756 P=1.2 MULT=1
MM1005 N_VPWR_M1005_d N_A_913_406#_M1005_g A_781_504# VPB PSHORT L=0.18 W=0.42
+ AD=0.140509 AS=0.1386 PD=1.05273 PS=1.08 NRD=0 NRS=128.976 M=1 R=2.33333
+ SA=90002.4 SB=90003.2 A=0.0756 P=1.2 MULT=1
MM1008 N_A_913_406#_M1008_d N_A_673_392#_M1008_g N_VPWR_M1005_d VPB PSHORT
+ L=0.18 W=1.12 AD=0.1568 AS=0.374691 PD=1.4 PS=2.80727 NRD=0.8668 NRS=6.1464
+ M=1 R=6.22222 SA=90001.4 SB=90002.2 A=0.2016 P=2.6 MULT=1
MM1019 N_VPWR_M1019_d N_RESET_B_M1019_g N_A_913_406#_M1008_d VPB PSHORT L=0.18
+ W=1.12 AD=0.4816 AS=0.1568 PD=1.98 PS=1.4 NRD=26.3783 NRS=0 M=1 R=6.22222
+ SA=90001.8 SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1006 N_Q_M1006_d N_A_913_406#_M1006_g N_VPWR_M1019_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.4816 PD=1.39 PS=1.98 NRD=0 NRS=75.6283 M=1 R=6.22222 SA=90002.9
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1009 N_Q_M1006_d N_A_913_406#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3808 PD=1.39 PS=2.92 NRD=0 NRS=8.7862 M=1 R=6.22222 SA=90003.3
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX22_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_ms__dlrtn_2.pxi.spice"
*
.ends
*
*

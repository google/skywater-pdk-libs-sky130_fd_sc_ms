* File: sky130_fd_sc_ms__mux2_2.spice
* Created: Wed Sep  2 12:11:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__mux2_2.pex.spice"
.subckt sky130_fd_sc_ms__mux2_2  VNB VPB A0 A1 S VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* S	S
* A1	A1
* A0	A0
* VPB	VPB
* VNB	VNB
MM1002 N_A_119_368#_M1002_d N_A0_M1002_g N_A_38_74#_M1002_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.21275 AS=0.2109 PD=1.315 PS=2.05 NRD=25.128 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002 A=0.111 P=1.78 MULT=1
MM1006 A_270_74# N_A1_M1006_g N_A_119_368#_M1002_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.0888 AS=0.21275 PD=0.98 PS=1.315 NRD=10.536 NRS=22.692 M=1 R=4.93333
+ SA=75000.9 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_S_M1009_g A_270_74# VNB NLOWVT L=0.15 W=0.74 AD=0.20535
+ AS=0.0888 PD=1.295 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75001.3
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1004 N_A_38_74#_M1004_d N_A_459_48#_M1004_g N_VGND_M1009_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2183 AS=0.20535 PD=2.07 PS=1.295 NRD=0 NRS=44.592 M=1 R=4.93333
+ SA=75002 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_S_M1012_g N_A_459_48#_M1012_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.117568 AS=0.15675 PD=0.984884 PS=1.67 NRD=21.816 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75001.3 A=0.0825 P=1.4 MULT=1
MM1003 N_X_M1003_d N_A_119_368#_M1003_g N_VGND_M1012_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.158182 PD=1.02 PS=1.32512 NRD=0 NRS=5.664 M=1 R=4.93333
+ SA=75000.6 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1013 N_X_M1003_d N_A_119_368#_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1000 N_A_119_368#_M1000_d N_A0_M1000_g N_A_27_368#_M1000_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1001 N_A_209_368#_M1001_d N_A1_M1001_g N_A_119_368#_M1000_d VPB PSHORT L=0.18
+ W=1 AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_S_M1007_g N_A_27_368#_M1007_s VPB PSHORT L=0.18 W=1
+ AD=0.185 AS=0.28 PD=1.37 PS=2.56 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1005 N_A_209_368#_M1005_d N_A_459_48#_M1005_g N_VPWR_M1007_d VPB PSHORT L=0.18
+ W=1 AD=0.28 AS=0.185 PD=2.56 PS=1.37 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90000.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_S_M1008_g N_A_459_48#_M1008_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1662 AS=0.2352 PD=1.27286 PS=2.24 NRD=33.49 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90001.2 A=0.1512 P=2.04 MULT=1
MM1010 N_X_M1010_d N_A_119_368#_M1010_g N_VPWR_M1008_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2216 PD=1.39 PS=1.69714 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1011 N_X_M1010_d N_A_119_368#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3752 PD=1.39 PS=2.91 NRD=0 NRS=3.5066 M=1 R=6.22222 SA=90001.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX14_noxref VNB VPB NWDIODE A=10.5276 P=15.04
c_591 A_270_74# 0 1.6439e-20 $X=1.35 $Y=0.37
*
.include "sky130_fd_sc_ms__mux2_2.pxi.spice"
*
.ends
*
*

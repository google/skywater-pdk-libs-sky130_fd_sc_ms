* File: sky130_fd_sc_ms__and2b_4.pxi.spice
* Created: Fri Aug 28 17:11:47 2020
* 
x_PM_SKY130_FD_SC_MS__AND2B_4%A_N N_A_N_M1008_g N_A_N_M1010_g A_N N_A_N_c_113_n
+ PM_SKY130_FD_SC_MS__AND2B_4%A_N
x_PM_SKY130_FD_SC_MS__AND2B_4%B N_B_M1009_g N_B_c_153_n N_B_M1000_g N_B_c_154_n
+ N_B_c_155_n N_B_c_147_n N_B_c_157_n N_B_M1017_g N_B_M1015_g N_B_c_158_n
+ N_B_c_149_n N_B_c_160_n N_B_c_150_n B B N_B_c_152_n
+ PM_SKY130_FD_SC_MS__AND2B_4%B
x_PM_SKY130_FD_SC_MS__AND2B_4%A_27_392# N_A_27_392#_M1010_s N_A_27_392#_M1008_s
+ N_A_27_392#_c_259_n N_A_27_392#_M1014_g N_A_27_392#_c_260_n
+ N_A_27_392#_c_261_n N_A_27_392#_c_262_n N_A_27_392#_M1016_g
+ N_A_27_392#_c_250_n N_A_27_392#_M1007_g N_A_27_392#_c_251_n
+ N_A_27_392#_c_252_n N_A_27_392#_M1013_g N_A_27_392#_c_264_n
+ N_A_27_392#_c_253_n N_A_27_392#_c_265_n N_A_27_392#_c_266_n
+ N_A_27_392#_c_254_n N_A_27_392#_c_255_n N_A_27_392#_c_256_n
+ N_A_27_392#_c_257_n N_A_27_392#_c_258_n PM_SKY130_FD_SC_MS__AND2B_4%A_27_392#
x_PM_SKY130_FD_SC_MS__AND2B_4%A_221_424# N_A_221_424#_M1007_d
+ N_A_221_424#_M1014_d N_A_221_424#_M1000_s N_A_221_424#_M1002_g
+ N_A_221_424#_M1001_g N_A_221_424#_M1003_g N_A_221_424#_M1006_g
+ N_A_221_424#_M1004_g N_A_221_424#_c_350_n N_A_221_424#_M1011_g
+ N_A_221_424#_c_351_n N_A_221_424#_c_352_n N_A_221_424#_c_353_n
+ N_A_221_424#_M1012_g N_A_221_424#_M1005_g N_A_221_424#_c_355_n
+ N_A_221_424#_c_362_n N_A_221_424#_c_363_n N_A_221_424#_c_368_n
+ N_A_221_424#_c_383_n N_A_221_424#_c_364_n N_A_221_424#_c_365_n
+ N_A_221_424#_c_356_n N_A_221_424#_c_366_n N_A_221_424#_c_457_p
+ N_A_221_424#_c_398_n N_A_221_424#_c_357_n
+ PM_SKY130_FD_SC_MS__AND2B_4%A_221_424#
x_PM_SKY130_FD_SC_MS__AND2B_4%VPWR N_VPWR_M1008_d N_VPWR_M1016_s N_VPWR_M1017_d
+ N_VPWR_M1003_s N_VPWR_M1005_s N_VPWR_c_515_n N_VPWR_c_516_n N_VPWR_c_517_n
+ N_VPWR_c_518_n N_VPWR_c_519_n N_VPWR_c_520_n N_VPWR_c_521_n N_VPWR_c_522_n
+ VPWR N_VPWR_c_523_n N_VPWR_c_524_n N_VPWR_c_525_n N_VPWR_c_526_n
+ N_VPWR_c_527_n N_VPWR_c_528_n N_VPWR_c_529_n N_VPWR_c_514_n
+ PM_SKY130_FD_SC_MS__AND2B_4%VPWR
x_PM_SKY130_FD_SC_MS__AND2B_4%X N_X_M1001_s N_X_M1011_s N_X_M1002_d N_X_M1004_d
+ N_X_c_594_n N_X_c_603_n N_X_c_604_n N_X_c_595_n N_X_c_596_n N_X_c_605_n
+ N_X_c_597_n N_X_c_606_n N_X_c_607_n N_X_c_598_n N_X_c_599_n N_X_c_600_n
+ N_X_c_601_n N_X_c_658_n X PM_SKY130_FD_SC_MS__AND2B_4%X
x_PM_SKY130_FD_SC_MS__AND2B_4%VGND N_VGND_M1010_d N_VGND_M1015_s N_VGND_M1006_d
+ N_VGND_M1012_d N_VGND_c_671_n N_VGND_c_672_n N_VGND_c_673_n N_VGND_c_674_n
+ N_VGND_c_675_n VGND N_VGND_c_676_n N_VGND_c_677_n N_VGND_c_678_n
+ N_VGND_c_679_n N_VGND_c_680_n N_VGND_c_681_n N_VGND_c_682_n
+ PM_SKY130_FD_SC_MS__AND2B_4%VGND
x_PM_SKY130_FD_SC_MS__AND2B_4%A_233_74# N_A_233_74#_M1009_d N_A_233_74#_M1013_s
+ N_A_233_74#_c_744_n N_A_233_74#_c_740_n N_A_233_74#_c_741_n
+ PM_SKY130_FD_SC_MS__AND2B_4%A_233_74#
cc_1 VNB N_A_N_M1010_g 0.0425761f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.69
cc_2 VNB A_N 0.00184438f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_3 VNB N_A_N_c_113_n 0.0197932f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.615
cc_4 VNB N_B_M1009_g 0.030296f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.46
cc_5 VNB N_B_c_147_n 0.00618265f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.615
cc_6 VNB N_B_M1015_g 0.0236056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_B_c_149_n 0.00619883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B_c_150_n 0.0253169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB B 0.00880776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B_c_152_n 0.0329693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_392#_c_250_n 0.0176057f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.78
cc_12 VNB N_A_27_392#_c_251_n 0.0123802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_392#_c_252_n 0.0173846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_392#_c_253_n 0.0368859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_392#_c_254_n 0.0179929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_392#_c_255_n 0.0154055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_392#_c_256_n 0.0189908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_392#_c_257_n 0.00357485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_392#_c_258_n 0.0432998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_221_424#_M1002_g 4.86301e-19 $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.615
cc_21 VNB N_A_221_424#_M1001_g 0.0212213f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.615
cc_22 VNB N_A_221_424#_M1003_g 4.77886e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_221_424#_M1006_g 0.0218136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_221_424#_M1004_g 4.76207e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_221_424#_c_350_n 0.0151946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_221_424#_c_351_n 0.0084015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_221_424#_c_352_n 0.0629841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_221_424#_c_353_n 0.0170341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_221_424#_M1005_g 0.0141907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_221_424#_c_355_n 0.0120724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_221_424#_c_356_n 0.00151958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_221_424#_c_357_n 0.00204131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_514_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_X_c_594_n 0.00179817f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.78
cc_35 VNB N_X_c_595_n 0.00296071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_X_c_596_n 0.00151717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_X_c_597_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_X_c_598_n 0.00879366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_X_c_599_n 0.0127874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_X_c_600_n 0.00248839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_601_n 0.00212146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB X 0.0161443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_671_n 0.00641543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_672_n 0.00568769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_673_n 0.00420532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_674_n 0.0125057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_675_n 0.0262963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_676_n 0.0383162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_677_n 0.0155668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_678_n 0.0183662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_679_n 0.027356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_680_n 0.00613614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_681_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_682_n 0.275826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_233_74#_c_740_n 0.00250269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_233_74#_c_741_n 0.00513172f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.615
cc_57 VPB N_A_N_M1008_g 0.0301726f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.46
cc_58 VPB A_N 0.0017388f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_59 VPB N_A_N_c_113_n 0.0146325f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.615
cc_60 VPB N_B_c_153_n 0.0168764f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.45
cc_61 VPB N_B_c_154_n 0.011729f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_B_c_155_n 0.0102749f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_63 VPB N_B_c_147_n 0.0145753f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.615
cc_64 VPB N_B_c_157_n 0.0168764f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.615
cc_65 VPB N_B_c_158_n 0.00761042f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_B_c_149_n 0.00562027f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_B_c_160_n 0.00327454f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_B_c_150_n 0.00489863f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB B 0.0039893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_27_392#_c_259_n 0.0173287f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=0.69
cc_71 VPB N_A_27_392#_c_260_n 0.0118759f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_27_392#_c_261_n 0.0102027f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=1.615
cc_73 VPB N_A_27_392#_c_262_n 0.016877f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.615
cc_74 VPB N_A_27_392#_c_251_n 0.0180254f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_27_392#_c_264_n 0.0134257f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_27_392#_c_265_n 0.00931663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_27_392#_c_266_n 0.0367061f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_27_392#_c_256_n 0.013946f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_221_424#_M1002_g 0.0223074f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.615
cc_80 VPB N_A_221_424#_M1003_g 0.0215928f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_221_424#_M1004_g 0.021563f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_221_424#_M1005_g 0.0289586f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_221_424#_c_362_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_221_424#_c_363_n 0.00167726f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_221_424#_c_364_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_221_424#_c_365_n 7.68838e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_221_424#_c_366_n 0.00136909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_515_n 0.00794822f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_89 VPB N_VPWR_c_516_n 0.0202859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_517_n 0.00891431f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_518_n 0.0199421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_519_n 0.00575094f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_520_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_521_n 0.0116777f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_522_n 0.0564386f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_523_n 0.0175529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_524_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_525_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_526_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_527_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_528_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_529_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_514_n 0.06954f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_X_c_603_n 0.00142836f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_X_c_604_n 0.00179594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_X_c_605_n 0.00338871f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_X_c_606_n 0.0028845f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_X_c_607_n 0.00179594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 N_A_N_M1010_g N_B_M1009_g 0.0251047f $X=0.59 $Y=0.69 $X2=0 $Y2=0
cc_110 N_A_N_M1008_g N_B_c_160_n 2.8555e-19 $X=0.495 $Y=2.46 $X2=0 $Y2=0
cc_111 A_N N_B_c_160_n 0.0267667f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_112 N_A_N_c_113_n N_B_c_160_n 8.54572e-19 $X=0.58 $Y=1.615 $X2=0 $Y2=0
cc_113 N_A_N_M1010_g N_B_c_150_n 0.00456823f $X=0.59 $Y=0.69 $X2=0 $Y2=0
cc_114 A_N N_B_c_150_n 0.00140103f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_115 N_A_N_c_113_n N_B_c_150_n 0.0130918f $X=0.58 $Y=1.615 $X2=0 $Y2=0
cc_116 N_A_N_M1008_g N_A_27_392#_c_261_n 0.0259267f $X=0.495 $Y=2.46 $X2=0 $Y2=0
cc_117 N_A_N_M1010_g N_A_27_392#_c_253_n 0.0117205f $X=0.59 $Y=0.69 $X2=0 $Y2=0
cc_118 N_A_N_M1008_g N_A_27_392#_c_265_n 8.69055e-19 $X=0.495 $Y=2.46 $X2=0
+ $Y2=0
cc_119 N_A_N_M1010_g N_A_27_392#_c_254_n 0.0115584f $X=0.59 $Y=0.69 $X2=0 $Y2=0
cc_120 A_N N_A_27_392#_c_254_n 0.0184339f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_121 N_A_N_c_113_n N_A_27_392#_c_254_n 0.00177632f $X=0.58 $Y=1.615 $X2=0
+ $Y2=0
cc_122 N_A_N_M1010_g N_A_27_392#_c_255_n 0.00449058f $X=0.59 $Y=0.69 $X2=0 $Y2=0
cc_123 A_N N_A_27_392#_c_255_n 0.00898631f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_124 N_A_N_c_113_n N_A_27_392#_c_255_n 0.00338244f $X=0.58 $Y=1.615 $X2=0
+ $Y2=0
cc_125 N_A_N_M1010_g N_A_27_392#_c_256_n 0.00572006f $X=0.59 $Y=0.69 $X2=0 $Y2=0
cc_126 A_N N_A_27_392#_c_256_n 0.0250408f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_127 N_A_N_c_113_n N_A_27_392#_c_256_n 0.0136844f $X=0.58 $Y=1.615 $X2=0 $Y2=0
cc_128 N_A_N_M1008_g N_A_221_424#_c_362_n 2.92115e-19 $X=0.495 $Y=2.46 $X2=0
+ $Y2=0
cc_129 N_A_N_M1008_g N_A_221_424#_c_368_n 5.72362e-19 $X=0.495 $Y=2.46 $X2=0
+ $Y2=0
cc_130 N_A_N_M1008_g N_VPWR_c_515_n 0.0203479f $X=0.495 $Y=2.46 $X2=0 $Y2=0
cc_131 A_N N_VPWR_c_515_n 0.0111957f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_132 N_A_N_c_113_n N_VPWR_c_515_n 0.00344958f $X=0.58 $Y=1.615 $X2=0 $Y2=0
cc_133 N_A_N_M1008_g N_VPWR_c_523_n 0.00460063f $X=0.495 $Y=2.46 $X2=0 $Y2=0
cc_134 N_A_N_M1008_g N_VPWR_c_514_n 0.00912261f $X=0.495 $Y=2.46 $X2=0 $Y2=0
cc_135 N_A_N_M1010_g N_VGND_c_671_n 0.00615346f $X=0.59 $Y=0.69 $X2=0 $Y2=0
cc_136 N_A_N_M1010_g N_VGND_c_679_n 0.00434272f $X=0.59 $Y=0.69 $X2=0 $Y2=0
cc_137 N_A_N_M1010_g N_VGND_c_682_n 0.00824713f $X=0.59 $Y=0.69 $X2=0 $Y2=0
cc_138 N_B_c_149_n N_A_27_392#_c_260_n 0.00594459f $X=2.045 $Y=1.705 $X2=0 $Y2=0
cc_139 N_B_c_160_n N_A_27_392#_c_261_n 0.00412153f $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_140 N_B_c_150_n N_A_27_392#_c_261_n 0.0210707f $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_141 N_B_c_153_n N_A_27_392#_c_262_n 0.0206104f $X=1.985 $Y=2.045 $X2=0 $Y2=0
cc_142 N_B_M1009_g N_A_27_392#_c_250_n 0.0251644f $X=1.09 $Y=0.69 $X2=0 $Y2=0
cc_143 N_B_c_149_n N_A_27_392#_c_251_n 0.0118894f $X=2.045 $Y=1.705 $X2=0 $Y2=0
cc_144 N_B_c_160_n N_A_27_392#_c_251_n 4.97671e-19 $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_145 B N_A_27_392#_c_251_n 0.0040484f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_146 N_B_c_152_n N_A_27_392#_c_251_n 0.00646392f $X=2.47 $Y=1.385 $X2=0 $Y2=0
cc_147 N_B_M1015_g N_A_27_392#_c_252_n 0.0283032f $X=2.47 $Y=0.69 $X2=0 $Y2=0
cc_148 N_B_c_155_n N_A_27_392#_c_264_n 0.00993433f $X=2.075 $Y=1.97 $X2=0 $Y2=0
cc_149 N_B_M1009_g N_A_27_392#_c_253_n 7.4234e-19 $X=1.09 $Y=0.69 $X2=0 $Y2=0
cc_150 N_B_M1009_g N_A_27_392#_c_254_n 0.0149394f $X=1.09 $Y=0.69 $X2=0 $Y2=0
cc_151 N_B_c_149_n N_A_27_392#_c_254_n 0.00950432f $X=2.045 $Y=1.705 $X2=0 $Y2=0
cc_152 N_B_c_160_n N_A_27_392#_c_254_n 0.0243488f $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_153 N_B_c_150_n N_A_27_392#_c_254_n 0.00446668f $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_154 N_B_M1009_g N_A_27_392#_c_257_n 6.47392e-19 $X=1.09 $Y=0.69 $X2=0 $Y2=0
cc_155 N_B_M1015_g N_A_27_392#_c_257_n 2.55667e-19 $X=2.47 $Y=0.69 $X2=0 $Y2=0
cc_156 N_B_c_149_n N_A_27_392#_c_257_n 0.0243539f $X=2.045 $Y=1.705 $X2=0 $Y2=0
cc_157 N_B_c_160_n N_A_27_392#_c_257_n 9.50602e-19 $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_158 N_B_c_150_n N_A_27_392#_c_257_n 6.23084e-19 $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_159 B N_A_27_392#_c_257_n 0.0192912f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_160 N_B_c_155_n N_A_27_392#_c_258_n 0.00272f $X=2.075 $Y=1.97 $X2=0 $Y2=0
cc_161 N_B_c_149_n N_A_27_392#_c_258_n 0.00607751f $X=2.045 $Y=1.705 $X2=0 $Y2=0
cc_162 N_B_c_160_n N_A_27_392#_c_258_n 0.00118989f $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_163 N_B_c_150_n N_A_27_392#_c_258_n 0.0214109f $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_164 B N_A_27_392#_c_258_n 0.00619253f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_165 N_B_c_152_n N_A_27_392#_c_258_n 0.00703692f $X=2.47 $Y=1.385 $X2=0 $Y2=0
cc_166 N_B_c_158_n N_A_221_424#_M1002_g 0.0264877f $X=2.415 $Y=1.97 $X2=0 $Y2=0
cc_167 N_B_M1015_g N_A_221_424#_M1001_g 0.0220476f $X=2.47 $Y=0.69 $X2=0 $Y2=0
cc_168 B N_A_221_424#_M1001_g 3.49507e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_169 N_B_c_152_n N_A_221_424#_M1001_g 0.0127101f $X=2.47 $Y=1.385 $X2=0 $Y2=0
cc_170 N_B_c_147_n N_A_221_424#_c_352_n 0.00894968f $X=2.38 $Y=1.895 $X2=0 $Y2=0
cc_171 B N_A_221_424#_c_352_n 8.4263e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_172 N_B_c_152_n N_A_221_424#_c_352_n 0.00443805f $X=2.47 $Y=1.385 $X2=0 $Y2=0
cc_173 N_B_c_153_n N_A_221_424#_c_362_n 6.99406e-19 $X=1.985 $Y=2.045 $X2=0
+ $Y2=0
cc_174 N_B_c_153_n N_A_221_424#_c_363_n 0.00888896f $X=1.985 $Y=2.045 $X2=0
+ $Y2=0
cc_175 N_B_c_155_n N_A_221_424#_c_363_n 0.00301435f $X=2.075 $Y=1.97 $X2=0 $Y2=0
cc_176 N_B_c_149_n N_A_221_424#_c_363_n 0.0460131f $X=2.045 $Y=1.705 $X2=0 $Y2=0
cc_177 N_B_c_149_n N_A_221_424#_c_368_n 0.00794883f $X=2.045 $Y=1.705 $X2=0
+ $Y2=0
cc_178 N_B_c_160_n N_A_221_424#_c_368_n 0.019374f $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_179 N_B_c_150_n N_A_221_424#_c_368_n 2.06523e-19 $X=1.14 $Y=1.52 $X2=0 $Y2=0
cc_180 N_B_M1015_g N_A_221_424#_c_383_n 0.0129721f $X=2.47 $Y=0.69 $X2=0 $Y2=0
cc_181 B N_A_221_424#_c_383_n 0.0275877f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_182 N_B_c_152_n N_A_221_424#_c_383_n 0.00178839f $X=2.47 $Y=1.385 $X2=0 $Y2=0
cc_183 N_B_c_153_n N_A_221_424#_c_364_n 0.0138613f $X=1.985 $Y=2.045 $X2=0 $Y2=0
cc_184 N_B_c_157_n N_A_221_424#_c_364_n 0.0137813f $X=2.435 $Y=2.045 $X2=0 $Y2=0
cc_185 N_B_c_157_n N_A_221_424#_c_365_n 0.00888896f $X=2.435 $Y=2.045 $X2=0
+ $Y2=0
cc_186 N_B_c_158_n N_A_221_424#_c_365_n 0.00387425f $X=2.415 $Y=1.97 $X2=0 $Y2=0
cc_187 B N_A_221_424#_c_365_n 0.0165376f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_188 N_B_c_152_n N_A_221_424#_c_365_n 0.00178207f $X=2.47 $Y=1.385 $X2=0 $Y2=0
cc_189 N_B_M1015_g N_A_221_424#_c_356_n 0.0052622f $X=2.47 $Y=0.69 $X2=0 $Y2=0
cc_190 B N_A_221_424#_c_356_n 0.0110703f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_191 N_B_c_152_n N_A_221_424#_c_356_n 6.31866e-19 $X=2.47 $Y=1.385 $X2=0 $Y2=0
cc_192 N_B_c_147_n N_A_221_424#_c_366_n 0.0023229f $X=2.38 $Y=1.895 $X2=0 $Y2=0
cc_193 N_B_c_158_n N_A_221_424#_c_366_n 0.00135928f $X=2.415 $Y=1.97 $X2=0 $Y2=0
cc_194 B N_A_221_424#_c_366_n 0.0115106f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_195 N_B_c_153_n N_A_221_424#_c_398_n 0.00108113f $X=1.985 $Y=2.045 $X2=0
+ $Y2=0
cc_196 N_B_c_154_n N_A_221_424#_c_398_n 0.00553073f $X=2.305 $Y=1.97 $X2=0 $Y2=0
cc_197 N_B_c_155_n N_A_221_424#_c_398_n 4.31578e-19 $X=2.075 $Y=1.97 $X2=0 $Y2=0
cc_198 N_B_c_157_n N_A_221_424#_c_398_n 0.00108113f $X=2.435 $Y=2.045 $X2=0
+ $Y2=0
cc_199 N_B_c_158_n N_A_221_424#_c_398_n 0.00157192f $X=2.415 $Y=1.97 $X2=0 $Y2=0
cc_200 B N_A_221_424#_c_398_n 0.0286849f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_201 N_B_c_147_n N_A_221_424#_c_357_n 3.22534e-19 $X=2.38 $Y=1.895 $X2=0 $Y2=0
cc_202 B N_A_221_424#_c_357_n 0.029241f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_203 N_B_c_152_n N_A_221_424#_c_357_n 0.00166039f $X=2.47 $Y=1.385 $X2=0 $Y2=0
cc_204 N_B_c_153_n N_VPWR_c_517_n 0.00667684f $X=1.985 $Y=2.045 $X2=0 $Y2=0
cc_205 N_B_c_153_n N_VPWR_c_518_n 0.005209f $X=1.985 $Y=2.045 $X2=0 $Y2=0
cc_206 N_B_c_157_n N_VPWR_c_518_n 0.005209f $X=2.435 $Y=2.045 $X2=0 $Y2=0
cc_207 N_B_c_157_n N_VPWR_c_519_n 0.00683535f $X=2.435 $Y=2.045 $X2=0 $Y2=0
cc_208 N_B_c_153_n N_VPWR_c_514_n 0.00982779f $X=1.985 $Y=2.045 $X2=0 $Y2=0
cc_209 N_B_c_157_n N_VPWR_c_514_n 0.00982779f $X=2.435 $Y=2.045 $X2=0 $Y2=0
cc_210 N_B_M1009_g N_VGND_c_671_n 0.0102293f $X=1.09 $Y=0.69 $X2=0 $Y2=0
cc_211 N_B_M1015_g N_VGND_c_672_n 0.00303986f $X=2.47 $Y=0.69 $X2=0 $Y2=0
cc_212 N_B_M1009_g N_VGND_c_676_n 0.00383152f $X=1.09 $Y=0.69 $X2=0 $Y2=0
cc_213 N_B_M1015_g N_VGND_c_676_n 0.00336923f $X=2.47 $Y=0.69 $X2=0 $Y2=0
cc_214 N_B_M1009_g N_VGND_c_682_n 0.00758251f $X=1.09 $Y=0.69 $X2=0 $Y2=0
cc_215 N_B_M1015_g N_VGND_c_682_n 0.00439691f $X=2.47 $Y=0.69 $X2=0 $Y2=0
cc_216 N_B_M1009_g N_A_233_74#_c_740_n 7.34787e-19 $X=1.09 $Y=0.69 $X2=0 $Y2=0
cc_217 N_B_M1015_g N_A_233_74#_c_741_n 0.0026545f $X=2.47 $Y=0.69 $X2=0 $Y2=0
cc_218 N_A_27_392#_c_259_n N_A_221_424#_c_362_n 0.0123686f $X=1.015 $Y=2.045
+ $X2=0 $Y2=0
cc_219 N_A_27_392#_c_262_n N_A_221_424#_c_362_n 0.0140218f $X=1.465 $Y=2.045
+ $X2=0 $Y2=0
cc_220 N_A_27_392#_c_262_n N_A_221_424#_c_363_n 0.00888896f $X=1.465 $Y=2.045
+ $X2=0 $Y2=0
cc_221 N_A_27_392#_c_264_n N_A_221_424#_c_363_n 0.00742071f $X=1.52 $Y=1.97
+ $X2=0 $Y2=0
cc_222 N_A_27_392#_c_259_n N_A_221_424#_c_368_n 0.00238091f $X=1.015 $Y=2.045
+ $X2=0 $Y2=0
cc_223 N_A_27_392#_c_260_n N_A_221_424#_c_368_n 0.0059939f $X=1.375 $Y=1.97
+ $X2=0 $Y2=0
cc_224 N_A_27_392#_c_261_n N_A_221_424#_c_368_n 0.0020407f $X=1.105 $Y=1.97
+ $X2=0 $Y2=0
cc_225 N_A_27_392#_c_262_n N_A_221_424#_c_368_n 0.00108113f $X=1.465 $Y=2.045
+ $X2=0 $Y2=0
cc_226 N_A_27_392#_c_264_n N_A_221_424#_c_368_n 4.43608e-19 $X=1.52 $Y=1.97
+ $X2=0 $Y2=0
cc_227 N_A_27_392#_c_250_n N_A_221_424#_c_383_n 0.00237855f $X=1.59 $Y=1.12
+ $X2=0 $Y2=0
cc_228 N_A_27_392#_c_252_n N_A_221_424#_c_383_n 0.0113406f $X=2.02 $Y=1.12 $X2=0
+ $Y2=0
cc_229 N_A_27_392#_c_257_n N_A_221_424#_c_383_n 0.0137945f $X=1.68 $Y=1.18 $X2=0
+ $Y2=0
cc_230 N_A_27_392#_c_258_n N_A_221_424#_c_383_n 9.53947e-19 $X=1.68 $Y=1.285
+ $X2=0 $Y2=0
cc_231 N_A_27_392#_c_262_n N_A_221_424#_c_364_n 6.21402e-19 $X=1.465 $Y=2.045
+ $X2=0 $Y2=0
cc_232 N_A_27_392#_c_259_n N_VPWR_c_515_n 0.00797656f $X=1.015 $Y=2.045 $X2=0
+ $Y2=0
cc_233 N_A_27_392#_c_266_n N_VPWR_c_515_n 0.0296759f $X=0.27 $Y=2.115 $X2=0
+ $Y2=0
cc_234 N_A_27_392#_c_259_n N_VPWR_c_516_n 0.005209f $X=1.015 $Y=2.045 $X2=0
+ $Y2=0
cc_235 N_A_27_392#_c_262_n N_VPWR_c_516_n 0.005209f $X=1.465 $Y=2.045 $X2=0
+ $Y2=0
cc_236 N_A_27_392#_c_262_n N_VPWR_c_517_n 0.00310234f $X=1.465 $Y=2.045 $X2=0
+ $Y2=0
cc_237 N_A_27_392#_c_264_n N_VPWR_c_517_n 3.56539e-19 $X=1.52 $Y=1.97 $X2=0
+ $Y2=0
cc_238 N_A_27_392#_c_266_n N_VPWR_c_523_n 0.0119584f $X=0.27 $Y=2.115 $X2=0
+ $Y2=0
cc_239 N_A_27_392#_c_259_n N_VPWR_c_514_n 0.00982779f $X=1.015 $Y=2.045 $X2=0
+ $Y2=0
cc_240 N_A_27_392#_c_262_n N_VPWR_c_514_n 0.00983003f $X=1.465 $Y=2.045 $X2=0
+ $Y2=0
cc_241 N_A_27_392#_c_266_n N_VPWR_c_514_n 0.00989813f $X=0.27 $Y=2.115 $X2=0
+ $Y2=0
cc_242 N_A_27_392#_c_250_n N_VGND_c_671_n 5.74073e-19 $X=1.59 $Y=1.12 $X2=0
+ $Y2=0
cc_243 N_A_27_392#_c_253_n N_VGND_c_671_n 0.0234524f $X=0.375 $Y=0.515 $X2=0
+ $Y2=0
cc_244 N_A_27_392#_c_254_n N_VGND_c_671_n 0.0238718f $X=1.515 $Y=1.18 $X2=0
+ $Y2=0
cc_245 N_A_27_392#_c_250_n N_VGND_c_676_n 0.00289603f $X=1.59 $Y=1.12 $X2=0
+ $Y2=0
cc_246 N_A_27_392#_c_252_n N_VGND_c_676_n 0.00289603f $X=2.02 $Y=1.12 $X2=0
+ $Y2=0
cc_247 N_A_27_392#_c_253_n N_VGND_c_679_n 0.0201415f $X=0.375 $Y=0.515 $X2=0
+ $Y2=0
cc_248 N_A_27_392#_c_250_n N_VGND_c_682_n 0.0035835f $X=1.59 $Y=1.12 $X2=0 $Y2=0
cc_249 N_A_27_392#_c_252_n N_VGND_c_682_n 0.00357919f $X=2.02 $Y=1.12 $X2=0
+ $Y2=0
cc_250 N_A_27_392#_c_253_n N_VGND_c_682_n 0.016615f $X=0.375 $Y=0.515 $X2=0
+ $Y2=0
cc_251 N_A_27_392#_c_254_n N_A_233_74#_c_744_n 0.0201258f $X=1.515 $Y=1.18 $X2=0
+ $Y2=0
cc_252 N_A_27_392#_c_250_n N_A_233_74#_c_741_n 0.0127013f $X=1.59 $Y=1.12 $X2=0
+ $Y2=0
cc_253 N_A_27_392#_c_252_n N_A_233_74#_c_741_n 0.0103014f $X=2.02 $Y=1.12 $X2=0
+ $Y2=0
cc_254 N_A_27_392#_c_257_n N_A_233_74#_c_741_n 0.00374521f $X=1.68 $Y=1.18 $X2=0
+ $Y2=0
cc_255 N_A_221_424#_c_363_n N_VPWR_M1016_s 0.00240242f $X=2.045 $Y=2.045 $X2=0
+ $Y2=0
cc_256 N_A_221_424#_c_365_n N_VPWR_M1017_d 0.00722852f $X=2.755 $Y=2.045 $X2=0
+ $Y2=0
cc_257 N_A_221_424#_c_366_n N_VPWR_M1017_d 0.00148303f $X=2.84 $Y=1.96 $X2=0
+ $Y2=0
cc_258 N_A_221_424#_c_362_n N_VPWR_c_515_n 0.0298716f $X=1.24 $Y=2.265 $X2=0
+ $Y2=0
cc_259 N_A_221_424#_c_368_n N_VPWR_c_515_n 0.00188897f $X=1.405 $Y=2.045 $X2=0
+ $Y2=0
cc_260 N_A_221_424#_c_362_n N_VPWR_c_516_n 0.0144623f $X=1.24 $Y=2.265 $X2=0
+ $Y2=0
cc_261 N_A_221_424#_c_362_n N_VPWR_c_517_n 0.0230789f $X=1.24 $Y=2.265 $X2=0
+ $Y2=0
cc_262 N_A_221_424#_c_363_n N_VPWR_c_517_n 0.018387f $X=2.045 $Y=2.045 $X2=0
+ $Y2=0
cc_263 N_A_221_424#_c_364_n N_VPWR_c_517_n 0.0240408f $X=2.21 $Y=2.265 $X2=0
+ $Y2=0
cc_264 N_A_221_424#_c_364_n N_VPWR_c_518_n 0.0144623f $X=2.21 $Y=2.265 $X2=0
+ $Y2=0
cc_265 N_A_221_424#_M1002_g N_VPWR_c_519_n 0.0126824f $X=2.955 $Y=2.4 $X2=0
+ $Y2=0
cc_266 N_A_221_424#_M1003_g N_VPWR_c_519_n 5.38044e-19 $X=3.405 $Y=2.4 $X2=0
+ $Y2=0
cc_267 N_A_221_424#_c_364_n N_VPWR_c_519_n 0.0240709f $X=2.21 $Y=2.265 $X2=0
+ $Y2=0
cc_268 N_A_221_424#_c_365_n N_VPWR_c_519_n 0.0211846f $X=2.755 $Y=2.045 $X2=0
+ $Y2=0
cc_269 N_A_221_424#_M1002_g N_VPWR_c_520_n 5.82312e-19 $X=2.955 $Y=2.4 $X2=0
+ $Y2=0
cc_270 N_A_221_424#_M1003_g N_VPWR_c_520_n 0.0154938f $X=3.405 $Y=2.4 $X2=0
+ $Y2=0
cc_271 N_A_221_424#_M1004_g N_VPWR_c_520_n 0.0154938f $X=3.855 $Y=2.4 $X2=0
+ $Y2=0
cc_272 N_A_221_424#_M1005_g N_VPWR_c_520_n 5.82312e-19 $X=4.305 $Y=2.4 $X2=0
+ $Y2=0
cc_273 N_A_221_424#_M1004_g N_VPWR_c_522_n 6.97239e-19 $X=3.855 $Y=2.4 $X2=0
+ $Y2=0
cc_274 N_A_221_424#_M1005_g N_VPWR_c_522_n 0.0208524f $X=4.305 $Y=2.4 $X2=0
+ $Y2=0
cc_275 N_A_221_424#_M1002_g N_VPWR_c_524_n 0.00460063f $X=2.955 $Y=2.4 $X2=0
+ $Y2=0
cc_276 N_A_221_424#_M1003_g N_VPWR_c_524_n 0.00460063f $X=3.405 $Y=2.4 $X2=0
+ $Y2=0
cc_277 N_A_221_424#_M1004_g N_VPWR_c_525_n 0.00460063f $X=3.855 $Y=2.4 $X2=0
+ $Y2=0
cc_278 N_A_221_424#_M1005_g N_VPWR_c_525_n 0.00460063f $X=4.305 $Y=2.4 $X2=0
+ $Y2=0
cc_279 N_A_221_424#_M1002_g N_VPWR_c_514_n 0.00908554f $X=2.955 $Y=2.4 $X2=0
+ $Y2=0
cc_280 N_A_221_424#_M1003_g N_VPWR_c_514_n 0.00908554f $X=3.405 $Y=2.4 $X2=0
+ $Y2=0
cc_281 N_A_221_424#_M1004_g N_VPWR_c_514_n 0.00908554f $X=3.855 $Y=2.4 $X2=0
+ $Y2=0
cc_282 N_A_221_424#_M1005_g N_VPWR_c_514_n 0.00908554f $X=4.305 $Y=2.4 $X2=0
+ $Y2=0
cc_283 N_A_221_424#_c_362_n N_VPWR_c_514_n 0.0118344f $X=1.24 $Y=2.265 $X2=0
+ $Y2=0
cc_284 N_A_221_424#_c_364_n N_VPWR_c_514_n 0.0118344f $X=2.21 $Y=2.265 $X2=0
+ $Y2=0
cc_285 N_A_221_424#_M1001_g N_X_c_594_n 0.00497662f $X=2.955 $Y=0.74 $X2=0 $Y2=0
cc_286 N_A_221_424#_M1006_g N_X_c_594_n 4.02861e-19 $X=3.395 $Y=0.74 $X2=0 $Y2=0
cc_287 N_A_221_424#_c_383_n N_X_c_594_n 0.0133617f $X=2.755 $Y=0.84 $X2=0 $Y2=0
cc_288 N_A_221_424#_c_356_n N_X_c_594_n 0.00379102f $X=2.84 $Y=1.32 $X2=0 $Y2=0
cc_289 N_A_221_424#_c_352_n N_X_c_603_n 0.00209661f $X=3.945 $Y=1.26 $X2=0 $Y2=0
cc_290 N_A_221_424#_c_366_n N_X_c_603_n 0.00561888f $X=2.84 $Y=1.96 $X2=0 $Y2=0
cc_291 N_A_221_424#_c_457_p N_X_c_603_n 0.0143383f $X=3.725 $Y=1.485 $X2=0 $Y2=0
cc_292 N_A_221_424#_M1002_g N_X_c_604_n 3.62369e-19 $X=2.955 $Y=2.4 $X2=0 $Y2=0
cc_293 N_A_221_424#_M1003_g N_X_c_604_n 3.62369e-19 $X=3.405 $Y=2.4 $X2=0 $Y2=0
cc_294 N_A_221_424#_M1006_g N_X_c_595_n 0.0128363f $X=3.395 $Y=0.74 $X2=0 $Y2=0
cc_295 N_A_221_424#_c_350_n N_X_c_595_n 0.01254f $X=3.86 $Y=1.185 $X2=0 $Y2=0
cc_296 N_A_221_424#_c_352_n N_X_c_595_n 0.00320407f $X=3.945 $Y=1.26 $X2=0 $Y2=0
cc_297 N_A_221_424#_c_457_p N_X_c_595_n 0.0413425f $X=3.725 $Y=1.485 $X2=0 $Y2=0
cc_298 N_A_221_424#_M1001_g N_X_c_596_n 8.1288e-19 $X=2.955 $Y=0.74 $X2=0 $Y2=0
cc_299 N_A_221_424#_c_352_n N_X_c_596_n 0.00264141f $X=3.945 $Y=1.26 $X2=0 $Y2=0
cc_300 N_A_221_424#_c_356_n N_X_c_596_n 0.0134877f $X=2.84 $Y=1.32 $X2=0 $Y2=0
cc_301 N_A_221_424#_c_457_p N_X_c_596_n 0.0143379f $X=3.725 $Y=1.485 $X2=0 $Y2=0
cc_302 N_A_221_424#_M1003_g N_X_c_605_n 0.0143902f $X=3.405 $Y=2.4 $X2=0 $Y2=0
cc_303 N_A_221_424#_M1004_g N_X_c_605_n 0.0161584f $X=3.855 $Y=2.4 $X2=0 $Y2=0
cc_304 N_A_221_424#_c_352_n N_X_c_605_n 0.00201785f $X=3.945 $Y=1.26 $X2=0 $Y2=0
cc_305 N_A_221_424#_c_457_p N_X_c_605_n 0.0411552f $X=3.725 $Y=1.485 $X2=0 $Y2=0
cc_306 N_A_221_424#_M1006_g N_X_c_597_n 6.54757e-19 $X=3.395 $Y=0.74 $X2=0 $Y2=0
cc_307 N_A_221_424#_c_350_n N_X_c_597_n 0.00939704f $X=3.86 $Y=1.185 $X2=0 $Y2=0
cc_308 N_A_221_424#_c_353_n N_X_c_597_n 3.97481e-19 $X=4.29 $Y=1.185 $X2=0 $Y2=0
cc_309 N_A_221_424#_M1004_g N_X_c_606_n 0.00404608f $X=3.855 $Y=2.4 $X2=0 $Y2=0
cc_310 N_A_221_424#_M1005_g N_X_c_606_n 0.00405038f $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_311 N_A_221_424#_M1004_g N_X_c_607_n 3.62369e-19 $X=3.855 $Y=2.4 $X2=0 $Y2=0
cc_312 N_A_221_424#_M1005_g N_X_c_607_n 3.62369e-19 $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_313 N_A_221_424#_c_353_n N_X_c_598_n 0.0148317f $X=4.29 $Y=1.185 $X2=0 $Y2=0
cc_314 N_A_221_424#_c_355_n N_X_c_598_n 8.29489e-19 $X=4.215 $Y=1.185 $X2=0
+ $Y2=0
cc_315 N_A_221_424#_M1005_g N_X_c_599_n 0.017865f $X=4.305 $Y=2.4 $X2=0 $Y2=0
cc_316 N_A_221_424#_c_351_n N_X_c_600_n 0.00208718f $X=4.215 $Y=1.26 $X2=0 $Y2=0
cc_317 N_A_221_424#_c_352_n N_X_c_600_n 0.00167782f $X=3.945 $Y=1.26 $X2=0 $Y2=0
cc_318 N_A_221_424#_c_457_p N_X_c_600_n 0.015065f $X=3.725 $Y=1.485 $X2=0 $Y2=0
cc_319 N_A_221_424#_c_350_n N_X_c_601_n 0.00156393f $X=3.86 $Y=1.185 $X2=0 $Y2=0
cc_320 N_A_221_424#_c_351_n N_X_c_601_n 0.00276997f $X=4.215 $Y=1.26 $X2=0 $Y2=0
cc_321 N_A_221_424#_c_353_n X 0.00806324f $X=4.29 $Y=1.185 $X2=0 $Y2=0
cc_322 N_A_221_424#_c_355_n X 0.00418807f $X=4.215 $Y=1.185 $X2=0 $Y2=0
cc_323 N_A_221_424#_c_457_p X 0.00476845f $X=3.725 $Y=1.485 $X2=0 $Y2=0
cc_324 N_A_221_424#_c_383_n N_VGND_M1015_s 0.00728075f $X=2.755 $Y=0.84 $X2=0
+ $Y2=0
cc_325 N_A_221_424#_c_356_n N_VGND_M1015_s 0.00219581f $X=2.84 $Y=1.32 $X2=0
+ $Y2=0
cc_326 N_A_221_424#_M1001_g N_VGND_c_672_n 0.00650608f $X=2.955 $Y=0.74 $X2=0
+ $Y2=0
cc_327 N_A_221_424#_M1006_g N_VGND_c_672_n 3.97853e-19 $X=3.395 $Y=0.74 $X2=0
+ $Y2=0
cc_328 N_A_221_424#_c_383_n N_VGND_c_672_n 0.0194555f $X=2.755 $Y=0.84 $X2=0
+ $Y2=0
cc_329 N_A_221_424#_M1001_g N_VGND_c_673_n 4.63452e-19 $X=2.955 $Y=0.74 $X2=0
+ $Y2=0
cc_330 N_A_221_424#_M1006_g N_VGND_c_673_n 0.00960479f $X=3.395 $Y=0.74 $X2=0
+ $Y2=0
cc_331 N_A_221_424#_c_350_n N_VGND_c_673_n 0.00347183f $X=3.86 $Y=1.185 $X2=0
+ $Y2=0
cc_332 N_A_221_424#_c_350_n N_VGND_c_675_n 5.14978e-19 $X=3.86 $Y=1.185 $X2=0
+ $Y2=0
cc_333 N_A_221_424#_c_353_n N_VGND_c_675_n 0.011928f $X=4.29 $Y=1.185 $X2=0
+ $Y2=0
cc_334 N_A_221_424#_c_383_n N_VGND_c_676_n 0.00199065f $X=2.755 $Y=0.84 $X2=0
+ $Y2=0
cc_335 N_A_221_424#_M1001_g N_VGND_c_677_n 0.00378853f $X=2.955 $Y=0.74 $X2=0
+ $Y2=0
cc_336 N_A_221_424#_M1006_g N_VGND_c_677_n 0.00383152f $X=3.395 $Y=0.74 $X2=0
+ $Y2=0
cc_337 N_A_221_424#_c_383_n N_VGND_c_677_n 3.38697e-19 $X=2.755 $Y=0.84 $X2=0
+ $Y2=0
cc_338 N_A_221_424#_c_350_n N_VGND_c_678_n 0.00434272f $X=3.86 $Y=1.185 $X2=0
+ $Y2=0
cc_339 N_A_221_424#_c_353_n N_VGND_c_678_n 0.00383152f $X=4.29 $Y=1.185 $X2=0
+ $Y2=0
cc_340 N_A_221_424#_M1001_g N_VGND_c_682_n 0.00706821f $X=2.955 $Y=0.74 $X2=0
+ $Y2=0
cc_341 N_A_221_424#_M1006_g N_VGND_c_682_n 0.0075764f $X=3.395 $Y=0.74 $X2=0
+ $Y2=0
cc_342 N_A_221_424#_c_350_n N_VGND_c_682_n 0.00821408f $X=3.86 $Y=1.185 $X2=0
+ $Y2=0
cc_343 N_A_221_424#_c_353_n N_VGND_c_682_n 0.0075754f $X=4.29 $Y=1.185 $X2=0
+ $Y2=0
cc_344 N_A_221_424#_c_383_n N_VGND_c_682_n 0.00675954f $X=2.755 $Y=0.84 $X2=0
+ $Y2=0
cc_345 N_A_221_424#_c_383_n N_A_233_74#_M1013_s 0.00423148f $X=2.755 $Y=0.84
+ $X2=0 $Y2=0
cc_346 N_A_221_424#_M1007_d N_A_233_74#_c_741_n 0.00168037f $X=1.665 $Y=0.37
+ $X2=0 $Y2=0
cc_347 N_A_221_424#_c_383_n N_A_233_74#_c_741_n 0.037476f $X=2.755 $Y=0.84 $X2=0
+ $Y2=0
cc_348 N_VPWR_c_519_n N_X_c_604_n 0.0230404f $X=2.73 $Y=2.465 $X2=0 $Y2=0
cc_349 N_VPWR_c_520_n N_X_c_604_n 0.0276528f $X=3.63 $Y=2.325 $X2=0 $Y2=0
cc_350 N_VPWR_c_524_n N_X_c_604_n 0.00749631f $X=3.465 $Y=3.33 $X2=0 $Y2=0
cc_351 N_VPWR_c_514_n N_X_c_604_n 0.0062048f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_352 N_VPWR_M1003_s N_X_c_605_n 0.00165831f $X=3.495 $Y=1.84 $X2=0 $Y2=0
cc_353 N_VPWR_c_520_n N_X_c_605_n 0.0170259f $X=3.63 $Y=2.325 $X2=0 $Y2=0
cc_354 N_VPWR_c_520_n N_X_c_607_n 0.0276528f $X=3.63 $Y=2.325 $X2=0 $Y2=0
cc_355 N_VPWR_c_522_n N_X_c_607_n 0.0332535f $X=4.53 $Y=1.985 $X2=0 $Y2=0
cc_356 N_VPWR_c_525_n N_X_c_607_n 0.00749631f $X=4.365 $Y=3.33 $X2=0 $Y2=0
cc_357 N_VPWR_c_514_n N_X_c_607_n 0.0062048f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_358 N_VPWR_c_522_n N_X_c_599_n 0.0279208f $X=4.53 $Y=1.985 $X2=0 $Y2=0
cc_359 N_VPWR_c_522_n N_X_c_658_n 0.00641267f $X=4.53 $Y=1.985 $X2=0 $Y2=0
cc_360 N_X_c_595_n N_VGND_M1006_d 0.00307253f $X=3.91 $Y=1.065 $X2=0 $Y2=0
cc_361 N_X_c_598_n N_VGND_M1012_d 0.00325695f $X=4.445 $Y=1.065 $X2=0 $Y2=0
cc_362 N_X_c_594_n N_VGND_c_672_n 0.0156353f $X=3.18 $Y=0.515 $X2=0 $Y2=0
cc_363 N_X_c_594_n N_VGND_c_673_n 0.0164868f $X=3.18 $Y=0.515 $X2=0 $Y2=0
cc_364 N_X_c_595_n N_VGND_c_673_n 0.015373f $X=3.91 $Y=1.065 $X2=0 $Y2=0
cc_365 N_X_c_597_n N_VGND_c_673_n 0.0286138f $X=4.075 $Y=0.515 $X2=0 $Y2=0
cc_366 N_X_c_597_n N_VGND_c_675_n 0.017215f $X=4.075 $Y=0.515 $X2=0 $Y2=0
cc_367 N_X_c_598_n N_VGND_c_675_n 0.023862f $X=4.445 $Y=1.065 $X2=0 $Y2=0
cc_368 N_X_c_594_n N_VGND_c_677_n 0.00749631f $X=3.18 $Y=0.515 $X2=0 $Y2=0
cc_369 N_X_c_597_n N_VGND_c_678_n 0.0109942f $X=4.075 $Y=0.515 $X2=0 $Y2=0
cc_370 N_X_c_594_n N_VGND_c_682_n 0.0062048f $X=3.18 $Y=0.515 $X2=0 $Y2=0
cc_371 N_X_c_597_n N_VGND_c_682_n 0.00904371f $X=4.075 $Y=0.515 $X2=0 $Y2=0
cc_372 N_VGND_c_671_n N_A_233_74#_c_740_n 0.0110102f $X=0.875 $Y=0.495 $X2=0
+ $Y2=0
cc_373 N_VGND_c_676_n N_A_233_74#_c_740_n 0.0122168f $X=2.57 $Y=0 $X2=0 $Y2=0
cc_374 N_VGND_c_682_n N_A_233_74#_c_740_n 0.00964373f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_375 N_VGND_c_672_n N_A_233_74#_c_741_n 0.0118255f $X=2.735 $Y=0.5 $X2=0 $Y2=0
cc_376 N_VGND_c_676_n N_A_233_74#_c_741_n 0.0401098f $X=2.57 $Y=0 $X2=0 $Y2=0
cc_377 N_VGND_c_682_n N_A_233_74#_c_741_n 0.0321234f $X=4.56 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__or4b_1.spice
* Created: Fri Aug 28 18:09:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__or4b_1.pex.spice"
.subckt sky130_fd_sc_ms__or4b_1  VNB VPB D_N C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_D_N_M1008_g N_A_27_74#_M1008_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.1155 AS=0.15675 PD=0.97 PS=1.67 NRD=15.264 NRS=0 M=1 R=3.66667 SA=75000.2
+ SB=75003.5 A=0.0825 P=1.4 MULT=1
MM1010 N_A_228_74#_M1010_d N_A_27_74#_M1010_g N_VGND_M1008_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.254375 AS=0.1155 PD=1.475 PS=0.97 NRD=0 NRS=15.264 M=1 R=3.66667
+ SA=75000.8 SB=75002.9 A=0.0825 P=1.4 MULT=1
MM1000 N_VGND_M1000_d N_C_M1000_g N_A_228_74#_M1010_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.1155 AS=0.254375 PD=0.97 PS=1.475 NRD=15.264 NRS=0 M=1 R=3.66667
+ SA=75001.9 SB=75001.9 A=0.0825 P=1.4 MULT=1
MM1006 N_A_228_74#_M1006_d N_B_M1006_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.077 AS=0.1155 PD=0.83 PS=0.97 NRD=0 NRS=15.264 M=1 R=3.66667 SA=75002.4
+ SB=75001.3 A=0.0825 P=1.4 MULT=1
MM1011 N_VGND_M1011_d N_A_M1011_g N_A_228_74#_M1006_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.136328 AS=0.077 PD=1.0531 PS=0.83 NRD=22.908 NRS=0 M=1 R=3.66667
+ SA=75002.9 SB=75000.9 A=0.0825 P=1.4 MULT=1
MM1002 N_X_M1002_d N_A_228_74#_M1002_g N_VGND_M1011_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.183422 PD=2.05 PS=1.4169 NRD=0 NRS=17.832 M=1 R=4.93333
+ SA=75002.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VPWR_M1001_d N_D_N_M1001_g N_A_27_74#_M1001_s VPB PSHORT L=0.18 W=0.84
+ AD=0.2772 AS=0.2352 PD=2.34 PS=2.24 NRD=10.5395 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1007 A_359_368# N_A_27_74#_M1007_g N_A_228_74#_M1007_s VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.28 PD=1.24 PS=2.56 NRD=12.7853 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90002.3 A=0.18 P=2.36 MULT=1
MM1009 A_443_368# N_C_M1009_g A_359_368# VPB PSHORT L=0.18 W=1 AD=0.12 AS=0.12
+ PD=1.24 PS=1.24 NRD=12.7853 NRS=12.7853 M=1 R=5.55556 SA=90000.6 SB=90001.8
+ A=0.18 P=2.36 MULT=1
MM1003 A_527_368# N_B_M1003_g A_443_368# VPB PSHORT L=0.18 W=1 AD=0.18 AS=0.12
+ PD=1.36 PS=1.24 NRD=24.6053 NRS=12.7853 M=1 R=5.55556 SA=90001 SB=90001.4
+ A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g A_527_368# VPB PSHORT L=0.18 W=1 AD=0.259245
+ AS=0.18 PD=1.53774 PS=1.36 NRD=36.9375 NRS=24.6053 M=1 R=5.55556 SA=90001.6
+ SB=90000.9 A=0.18 P=2.36 MULT=1
MM1005 N_X_M1005_d N_A_228_74#_M1005_g N_VPWR_M1004_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.290355 PD=2.8 PS=1.72226 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90002 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__or4b_1.pxi.spice"
*
.ends
*
*

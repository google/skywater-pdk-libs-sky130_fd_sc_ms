* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sedfxtp_4 CLK D DE SCD SCE VGND VNB VPB VPWR Q
X0 a_37_464# D a_129_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X1 a_1902_508# a_1943_53# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X2 a_1858_79# a_1943_53# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 VPWR CLK a_1313_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X4 a_1756_97# a_1313_74# a_1902_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X5 VGND a_2403_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VGND SCD a_1044_125# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X7 Q a_2403_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_631_87# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X9 a_2403_74# a_1510_74# a_2589_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X10 a_129_464# a_177_290# VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X11 a_37_464# D a_135_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X12 VPWR a_2403_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X13 a_37_464# SCE a_661_113# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X14 a_2589_508# a_545_87# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X15 a_497_113# a_545_87# a_37_464# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X16 VGND a_2403_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 a_177_290# DE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X18 VPWR a_2403_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X19 VGND a_2403_74# a_545_87# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X20 VPWR DE a_575_463# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X21 a_661_113# a_1510_74# a_1756_97# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X22 Q a_2403_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 VPWR SCD a_1074_455# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X24 a_1756_97# a_1510_74# a_1858_79# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X25 VPWR a_1313_74# a_1510_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X26 a_37_464# a_631_87# a_661_113# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X27 VPWR a_2403_74# a_545_87# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X28 a_1044_125# SCE a_661_113# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X29 VGND a_1943_53# a_2331_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X30 VPWR a_1756_97# a_1943_53# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X31 VGND a_1756_97# a_1943_53# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X32 VGND a_1313_74# a_1510_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X33 a_2295_392# a_1313_74# a_2403_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X34 a_2331_74# a_1510_74# a_2403_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X35 Q a_2403_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X36 a_575_463# a_545_87# a_37_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X37 a_661_113# a_1313_74# a_1756_97# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X38 a_2498_74# a_545_87# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X39 a_1074_455# a_631_87# a_661_113# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X40 VGND a_177_290# a_497_113# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X41 VGND CLK a_1313_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X42 VPWR a_1943_53# a_2295_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X43 Q a_2403_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X44 a_177_290# DE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X45 a_2403_74# a_1313_74# a_2498_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X46 a_631_87# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X47 a_135_74# DE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
.ends

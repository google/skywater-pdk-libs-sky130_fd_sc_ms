* NGSPICE file created from sky130_fd_sc_ms__mux2_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__mux2_2 A0 A1 S VGND VNB VPB VPWR X
M1000 a_119_368# A0 a_27_368# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=5.6e+11p ps=5.12e+06u
M1001 a_209_368# A1 a_119_368# VPB pshort w=1e+06u l=180000u
+  ad=5.6e+11p pd=5.12e+06u as=0p ps=0u
M1002 a_119_368# A0 a_38_74# VNB nlowvt w=740000u l=150000u
+  ad=4.255e+11p pd=2.63e+06u as=4.292e+11p ps=4.12e+06u
M1003 X a_119_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=9.4915e+11p ps=7.09e+06u
M1004 a_38_74# a_459_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_209_368# a_459_48# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=1.133e+12p ps=8.62e+06u
M1006 a_270_74# A1 a_119_368# VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=0p ps=0u
M1007 VPWR S a_27_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR S a_459_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1009 VGND S a_270_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_119_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1011 VPWR a_119_368# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND S a_459_48# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1013 VGND a_119_368# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


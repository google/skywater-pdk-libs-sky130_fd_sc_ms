* File: sky130_fd_sc_ms__or3_4.spice
* Created: Wed Sep  2 12:28:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__or3_4.pex.spice"
.subckt sky130_fd_sc_ms__or3_4  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_C_M1008_g N_A_305_388#_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1332 AS=0.2109 PD=1.1 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1015 N_A_305_388#_M1015_d N_B_M1015_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1258 AS=0.1332 PD=1.08 PS=1.1 NRD=9.72 NRS=1.62 M=1 R=4.93333 SA=75000.7
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A_M1001_g N_A_305_388#_M1015_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1258 PD=1.09 PS=1.08 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1000 N_X_M1000_d N_A_305_388#_M1000_g N_VGND_M1001_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.10545 AS=0.1295 PD=1.025 PS=1.09 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75001.7
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1002 N_X_M1000_d N_A_305_388#_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10545 AS=0.1258 PD=1.025 PS=1.08 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1010 N_X_M1010_d N_A_305_388#_M1010_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1258 PD=1.02 PS=1.08 NRD=0 NRS=9.72 M=1 R=4.93333 SA=75002.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1016 N_X_M1010_d N_A_305_388#_M1016_g N_VGND_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_A_119_388#_M1006_s VPB PSHORT L=0.18 W=1
+ AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90004.5 A=0.18 P=2.36 MULT=1
MM1009 N_A_119_388#_M1006_s N_B_M1009_g N_A_209_388#_M1009_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.15 PD=1.27 PS=1.3 NRD=0 NRS=1.9503 M=1 R=5.55556 SA=90000.6
+ SB=90004 A=0.18 P=2.36 MULT=1
MM1003 N_A_305_388#_M1003_d N_C_M1003_g N_A_209_388#_M1009_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.15 PD=1.27 PS=1.3 NRD=0 NRS=1.9503 M=1 R=5.55556 SA=90001.1
+ SB=90003.5 A=0.18 P=2.36 MULT=1
MM1005 N_A_305_388#_M1003_d N_C_M1005_g N_A_209_388#_M1005_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.1625 PD=1.27 PS=1.325 NRD=0 NRS=3.9203 M=1 R=5.55556
+ SA=90001.6 SB=90003.1 A=0.18 P=2.36 MULT=1
MM1014 N_A_119_388#_M1014_d N_B_M1014_g N_A_209_388#_M1005_s VPB PSHORT L=0.18
+ W=1 AD=0.16 AS=0.1625 PD=1.32 PS=1.325 NRD=8.8453 NRS=4.9053 M=1 R=5.55556
+ SA=90002.1 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1013_d N_A_M1013_g N_A_119_388#_M1014_d VPB PSHORT L=0.18 W=1
+ AD=0.181887 AS=0.16 PD=1.39151 PS=1.32 NRD=15.7403 NRS=0 M=1 R=5.55556
+ SA=90002.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1004 N_X_M1004_d N_A_305_388#_M1004_g N_VPWR_M1013_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.203713 PD=1.39 PS=1.55849 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.8
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1007 N_X_M1004_d N_A_305_388#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.2
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1011 N_X_M1011_d N_A_305_388#_M1011_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.7
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1012 N_X_M1011_d N_A_305_388#_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX17_noxref VNB VPB NWDIODE A=10.5276 P=15.04
*
.include "sky130_fd_sc_ms__or3_4.pxi.spice"
*
.ends
*
*

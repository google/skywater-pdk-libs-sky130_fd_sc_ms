* File: sky130_fd_sc_ms__o311ai_2.spice
* Created: Fri Aug 28 18:01:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o311ai_2.pex.spice"
.subckt sky130_fd_sc_ms__o311ai_2  VNB VPB A1 A2 A3 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1003 N_A_27_74#_M1003_d N_A1_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1258 PD=2.05 PS=1.08 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.6 A=0.111 P=1.78 MULT=1
MM1018 N_A_27_74#_M1018_d N_A1_M1018_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1258 AS=0.1258 PD=1.08 PS=1.08 NRD=0 NRS=9.72 M=1 R=4.93333 SA=75000.7
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_A2_M1012_g N_A_27_74#_M1018_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1073 AS=0.1258 PD=1.03 PS=1.08 NRD=1.62 NRS=9.72 M=1 R=4.93333 SA=75001.2
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1012_d N_A2_M1013_g N_A_27_74#_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1073 AS=0.1184 PD=1.03 PS=1.06 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A3_M1009_g N_A_27_74#_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1147 AS=0.1184 PD=1.05 PS=1.06 NRD=4.86 NRS=6.48 M=1 R=4.93333 SA=75002.1
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1009_d N_A3_M1016_g N_A_27_74#_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1147 AS=0.1036 PD=1.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.6
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1008 N_A_670_74#_M1008_d N_B1_M1008_g N_A_27_74#_M1016_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75003 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1015 N_A_670_74#_M1008_d N_B1_M1015_g N_A_27_74#_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1554 AS=0.2109 PD=1.16 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75003.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_A_670_74#_M1004_d N_C1_M1004_g N_Y_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1011 N_A_670_74#_M1004_d N_C1_M1011_g N_Y_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g N_A_28_368#_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1568 AS=0.3136 PD=1.4 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1014 N_VPWR_M1005_d N_A1_M1014_g N_A_28_368#_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1568 AS=0.1736 PD=1.4 PS=1.43 NRD=0.8668 NRS=6.1464 M=1 R=6.22222
+ SA=90000.6 SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1001 N_A_310_368#_M1001_d N_A2_M1001_g N_A_28_368#_M1014_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1904 AS=0.1736 PD=1.46 PS=1.43 NRD=11.426 NRS=0 M=1 R=6.22222
+ SA=90001.1 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1002 N_A_310_368#_M1001_d N_A2_M1002_g N_A_28_368#_M1002_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1904 AS=0.3136 PD=1.46 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.7
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1017 N_A_310_368#_M1017_d N_A3_M1017_g N_Y_M1017_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1019 N_A_310_368#_M1017_d N_A3_M1019_g N_Y_M1019_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90002 A=0.2016 P=2.6 MULT=1
MM1000 N_VPWR_M1000_d N_B1_M1000_g N_Y_M1019_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1006 N_VPWR_M1000_d N_B1_M1006_g N_Y_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1007 N_VPWR_M1007_d N_C1_M1007_g N_Y_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1010 N_VPWR_M1007_d N_C1_M1010_g N_Y_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.4
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ms__o311ai_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__o221a_4.pxi.spice
* Created: Fri Aug 28 17:57:13 2020
* 
x_PM_SKY130_FD_SC_MS__O221A_4%C1 N_C1_M1015_g N_C1_M1012_g N_C1_M1014_g
+ N_C1_M1016_g C1 C1 N_C1_c_144_n PM_SKY130_FD_SC_MS__O221A_4%C1
x_PM_SKY130_FD_SC_MS__O221A_4%B2 N_B2_M1004_g N_B2_M1019_g N_B2_M1021_g
+ N_B2_M1025_g B2 B2 N_B2_c_189_n PM_SKY130_FD_SC_MS__O221A_4%B2
x_PM_SKY130_FD_SC_MS__O221A_4%B1 N_B1_c_233_n N_B1_M1008_g N_B1_M1001_g
+ N_B1_c_236_n N_B1_c_237_n N_B1_M1011_g N_B1_M1023_g N_B1_c_240_n N_B1_c_241_n
+ B1 B1 B1 N_B1_c_243_n N_B1_c_244_n PM_SKY130_FD_SC_MS__O221A_4%B1
x_PM_SKY130_FD_SC_MS__O221A_4%A2 N_A2_M1007_g N_A2_M1009_g N_A2_M1010_g
+ N_A2_M1017_g A2 N_A2_c_321_n PM_SKY130_FD_SC_MS__O221A_4%A2
x_PM_SKY130_FD_SC_MS__O221A_4%A1 N_A1_M1013_g N_A1_M1006_g N_A1_c_368_n
+ N_A1_c_369_n N_A1_M1018_g N_A1_M1024_g N_A1_c_371_n A1 N_A1_c_372_n
+ N_A1_c_373_n PM_SKY130_FD_SC_MS__O221A_4%A1
x_PM_SKY130_FD_SC_MS__O221A_4%A_114_125# N_A_114_125#_M1012_s
+ N_A_114_125#_M1015_d N_A_114_125#_M1019_d N_A_114_125#_M1007_d
+ N_A_114_125#_c_441_n N_A_114_125#_M1002_g N_A_114_125#_M1000_g
+ N_A_114_125#_c_442_n N_A_114_125#_M1005_g N_A_114_125#_M1003_g
+ N_A_114_125#_M1020_g N_A_114_125#_c_443_n N_A_114_125#_M1022_g
+ N_A_114_125#_c_444_n N_A_114_125#_c_445_n N_A_114_125#_M1027_g
+ N_A_114_125#_M1026_g N_A_114_125#_c_447_n N_A_114_125#_c_448_n
+ N_A_114_125#_c_458_n N_A_114_125#_c_449_n N_A_114_125#_c_450_n
+ N_A_114_125#_c_451_n N_A_114_125#_c_478_n N_A_114_125#_c_474_n
+ N_A_114_125#_c_479_n N_A_114_125#_c_493_n N_A_114_125#_c_460_n
+ N_A_114_125#_c_452_n N_A_114_125#_c_556_p N_A_114_125#_c_481_n
+ N_A_114_125#_c_495_n N_A_114_125#_c_453_n
+ PM_SKY130_FD_SC_MS__O221A_4%A_114_125#
x_PM_SKY130_FD_SC_MS__O221A_4%VPWR N_VPWR_M1015_s N_VPWR_M1016_s N_VPWR_M1023_s
+ N_VPWR_M1024_s N_VPWR_M1003_s N_VPWR_M1026_s N_VPWR_c_618_n N_VPWR_c_619_n
+ N_VPWR_c_620_n N_VPWR_c_621_n N_VPWR_c_622_n N_VPWR_c_623_n N_VPWR_c_624_n
+ N_VPWR_c_625_n VPWR N_VPWR_c_626_n N_VPWR_c_627_n N_VPWR_c_628_n
+ N_VPWR_c_629_n N_VPWR_c_630_n N_VPWR_c_631_n N_VPWR_c_632_n N_VPWR_c_633_n
+ N_VPWR_c_634_n N_VPWR_c_617_n PM_SKY130_FD_SC_MS__O221A_4%VPWR
x_PM_SKY130_FD_SC_MS__O221A_4%A_300_387# N_A_300_387#_M1008_d
+ N_A_300_387#_M1021_s N_A_300_387#_c_714_n N_A_300_387#_c_712_n
+ N_A_300_387#_c_713_n N_A_300_387#_c_719_n
+ PM_SKY130_FD_SC_MS__O221A_4%A_300_387#
x_PM_SKY130_FD_SC_MS__O221A_4%A_766_387# N_A_766_387#_M1013_d
+ N_A_766_387#_M1017_s N_A_766_387#_c_738_n N_A_766_387#_c_736_n
+ N_A_766_387#_c_737_n N_A_766_387#_c_746_n
+ PM_SKY130_FD_SC_MS__O221A_4%A_766_387#
x_PM_SKY130_FD_SC_MS__O221A_4%X N_X_M1002_s N_X_M1022_s N_X_M1000_d N_X_M1020_d
+ N_X_c_760_n N_X_c_770_n N_X_c_765_n N_X_c_776_n N_X_c_780_n N_X_c_783_n
+ N_X_c_761_n N_X_c_766_n N_X_c_792_n N_X_c_762_n N_X_c_763_n X
+ PM_SKY130_FD_SC_MS__O221A_4%X
x_PM_SKY130_FD_SC_MS__O221A_4%A_27_125# N_A_27_125#_M1012_d N_A_27_125#_M1014_d
+ N_A_27_125#_M1004_s N_A_27_125#_M1011_d N_A_27_125#_c_828_n
+ N_A_27_125#_c_829_n N_A_27_125#_c_830_n N_A_27_125#_c_831_n
+ N_A_27_125#_c_832_n N_A_27_125#_c_833_n N_A_27_125#_c_834_n
+ N_A_27_125#_c_835_n N_A_27_125#_c_836_n N_A_27_125#_c_837_n
+ PM_SKY130_FD_SC_MS__O221A_4%A_27_125#
x_PM_SKY130_FD_SC_MS__O221A_4%A_300_125# N_A_300_125#_M1001_s
+ N_A_300_125#_M1025_d N_A_300_125#_M1006_s N_A_300_125#_M1010_s
+ N_A_300_125#_c_896_n N_A_300_125#_c_897_n N_A_300_125#_c_898_n
+ N_A_300_125#_c_948_n N_A_300_125#_c_899_n N_A_300_125#_c_900_n
+ N_A_300_125#_c_920_n N_A_300_125#_c_932_n N_A_300_125#_c_901_n
+ N_A_300_125#_c_902_n N_A_300_125#_c_903_n
+ PM_SKY130_FD_SC_MS__O221A_4%A_300_125#
x_PM_SKY130_FD_SC_MS__O221A_4%VGND N_VGND_M1006_d N_VGND_M1009_d N_VGND_M1018_d
+ N_VGND_M1005_d N_VGND_M1027_d N_VGND_c_965_n N_VGND_c_966_n N_VGND_c_967_n
+ N_VGND_c_968_n N_VGND_c_969_n N_VGND_c_970_n N_VGND_c_971_n N_VGND_c_972_n
+ N_VGND_c_973_n N_VGND_c_974_n VGND N_VGND_c_975_n N_VGND_c_976_n
+ N_VGND_c_977_n N_VGND_c_978_n N_VGND_c_979_n N_VGND_c_980_n
+ PM_SKY130_FD_SC_MS__O221A_4%VGND
cc_1 VNB N_C1_M1012_g 0.0248304f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.945
cc_2 VNB N_C1_M1014_g 0.0197165f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.945
cc_3 VNB C1 0.00959695f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_C1_c_144_n 0.0391224f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.61
cc_5 VNB N_B2_M1004_g 0.0195673f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.435
cc_6 VNB N_B2_M1025_g 0.0185522f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.435
cc_7 VNB B2 0.00250521f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_8 VNB N_B2_c_189_n 0.0254617f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.61
cc_9 VNB N_B1_c_233_n 0.00706085f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.775
cc_10 VNB N_B1_M1008_g 0.0133785f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.435
cc_11 VNB N_B1_M1001_g 0.0287863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B1_c_236_n 0.126455f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.445
cc_13 VNB N_B1_c_237_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.945
cc_14 VNB N_B1_M1011_g 0.0211117f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.775
cc_15 VNB N_B1_M1023_g 0.00296389f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_16 VNB N_B1_c_240_n 0.0634657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B1_c_241_n 0.00478553f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.61
cc_18 VNB B1 0.00468429f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.61
cc_19 VNB N_B1_c_243_n 0.0124943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B1_c_244_n 0.0125846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A2_M1009_g 0.0196145f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.945
cc_22 VNB N_A2_M1010_g 0.0194573f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.945
cc_23 VNB A2 0.0010959f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_24 VNB N_A2_c_321_n 0.0262754f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.61
cc_25 VNB N_A1_M1013_g 0.00865647f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.435
cc_26 VNB N_A1_M1006_g 0.0226908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A1_c_368_n 0.0923141f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.445
cc_28 VNB N_A1_c_369_n 0.00976419f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.945
cc_29 VNB N_A1_M1018_g 0.0277553f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.435
cc_30 VNB N_A1_c_371_n 0.0129769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A1_c_372_n 0.0255242f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.61
cc_32 VNB N_A1_c_373_n 0.00635152f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.61
cc_33 VNB N_A_114_125#_c_441_n 0.0181187f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.775
cc_34 VNB N_A_114_125#_c_442_n 0.0173169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_114_125#_c_443_n 0.0176839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_114_125#_c_444_n 0.0151179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_114_125#_c_445_n 0.0193836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_114_125#_M1026_g 0.00213502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_114_125#_c_447_n 0.0230631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_114_125#_c_448_n 0.00200866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_114_125#_c_449_n 0.00119414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_114_125#_c_450_n 0.00177795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_114_125#_c_451_n 0.00781354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_114_125#_c_452_n 0.00426668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_114_125#_c_453_n 0.0515424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VPWR_c_617_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_X_c_760_n 0.00256408f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.435
cc_48 VNB N_X_c_761_n 0.0029512f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.61
cc_49 VNB N_X_c_762_n 2.03777e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_X_c_763_n 0.00109461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB X 0.00795563f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_27_125#_c_828_n 0.0362546f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.435
cc_53 VNB N_A_27_125#_c_829_n 0.0145686f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_54 VNB N_A_27_125#_c_830_n 0.0103479f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_55 VNB N_A_27_125#_c_831_n 0.0024541f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.61
cc_56 VNB N_A_27_125#_c_832_n 0.0104965f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.61
cc_57 VNB N_A_27_125#_c_833_n 0.00275908f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.61
cc_58 VNB N_A_27_125#_c_834_n 0.013376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_27_125#_c_835_n 0.00433773f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.612
cc_60 VNB N_A_27_125#_c_836_n 0.00279016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_27_125#_c_837_n 0.00380446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_300_125#_c_896_n 0.00535119f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=1.775
cc_63 VNB N_A_300_125#_c_897_n 0.0022314f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.435
cc_64 VNB N_A_300_125#_c_898_n 0.00361466f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_65 VNB N_A_300_125#_c_899_n 0.0111664f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.61
cc_66 VNB N_A_300_125#_c_900_n 0.00174318f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.61
cc_67 VNB N_A_300_125#_c_901_n 0.00223616f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.612
cc_68 VNB N_A_300_125#_c_902_n 0.00222589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_300_125#_c_903_n 0.00204476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_965_n 0.00996043f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_71 VNB N_VGND_c_966_n 0.0043165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_967_n 0.0133036f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.61
cc_73 VNB N_VGND_c_968_n 0.0110731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_969_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_970_n 0.0537609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_971_n 0.014017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_972_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_973_n 0.0170938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_974_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_975_n 0.0834355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_976_n 0.0175142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_977_n 0.0192529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_978_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_979_n 0.0076939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_980_n 0.405249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VPB N_C1_M1015_g 0.0253237f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.435
cc_87 VPB N_C1_M1016_g 0.0204461f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.435
cc_88 VPB C1 0.0114774f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_89 VPB N_C1_c_144_n 0.0237392f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.61
cc_90 VPB N_B2_M1019_g 0.0201486f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.945
cc_91 VPB N_B2_M1021_g 0.019544f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.945
cc_92 VPB B2 0.00455134f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_93 VPB N_B2_c_189_n 0.0141956f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.61
cc_94 VPB N_B1_M1008_g 0.0276273f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.435
cc_95 VPB N_B1_M1023_g 0.0305681f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_96 VPB B1 0.00954549f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.61
cc_97 VPB N_B1_c_244_n 0.0158044f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A2_M1007_g 0.0201024f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.435
cc_99 VPB N_A2_M1017_g 0.0203783f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.435
cc_100 VPB A2 0.00216666f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_101 VPB N_A2_c_321_n 0.0152296f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.61
cc_102 VPB N_A1_M1013_g 0.0305262f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.435
cc_103 VPB N_A1_M1024_g 0.026112f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_104 VPB N_A1_c_372_n 0.00555062f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.61
cc_105 VPB N_A1_c_373_n 0.00342849f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.61
cc_106 VPB N_A_114_125#_M1000_g 0.0218995f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_107 VPB N_A_114_125#_M1003_g 0.0221559f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.61
cc_108 VPB N_A_114_125#_M1020_g 0.0212859f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_114_125#_M1026_g 0.0263227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_114_125#_c_458_n 0.00241627f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_114_125#_c_451_n 0.00526214f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_114_125#_c_460_n 0.00119912f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_114_125#_c_453_n 0.00943905f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_618_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_619_n 0.050625f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.61
cc_116 VPB N_VPWR_c_620_n 0.00692241f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.61
cc_117 VPB N_VPWR_c_621_n 0.0145886f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_622_n 0.00649384f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_623_n 0.00554449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_624_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_625_n 0.0498587f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_626_n 0.0207267f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_627_n 0.0383359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_628_n 0.0405655f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_629_n 0.0204461f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_630_n 0.0196506f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_631_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_632_n 0.013727f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_633_n 0.00613202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_634_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_617_n 0.104024f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_300_387#_c_712_n 0.00654042f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.945
cc_133 VPB N_A_300_387#_c_713_n 0.0038297f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_766_387#_c_736_n 0.00723084f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.945
cc_135 VPB N_A_766_387#_c_737_n 0.0024962f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_X_c_765_n 0.00276927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_X_c_766_n 0.00276145f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.612
cc_138 VPB N_X_c_762_n 0.00166836f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB X 0.00910174f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 N_C1_M1014_g N_B1_c_233_n 0.00304803f $X=0.925 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_141 N_C1_c_144_n N_B1_M1008_g 0.0400131f $X=0.955 $Y=1.61 $X2=0 $Y2=0
cc_142 N_C1_M1014_g N_B1_M1001_g 0.019296f $X=0.925 $Y=0.945 $X2=0 $Y2=0
cc_143 N_C1_M1012_g N_A_114_125#_c_448_n 0.00580887f $X=0.495 $Y=0.945 $X2=0
+ $Y2=0
cc_144 N_C1_M1015_g N_A_114_125#_c_458_n 0.0110696f $X=0.505 $Y=2.435 $X2=0
+ $Y2=0
cc_145 N_C1_M1016_g N_A_114_125#_c_458_n 0.0117191f $X=0.955 $Y=2.435 $X2=0
+ $Y2=0
cc_146 N_C1_M1014_g N_A_114_125#_c_449_n 0.011584f $X=0.925 $Y=0.945 $X2=0 $Y2=0
cc_147 C1 N_A_114_125#_c_449_n 0.00696157f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_148 N_C1_c_144_n N_A_114_125#_c_449_n 0.00140962f $X=0.955 $Y=1.61 $X2=0
+ $Y2=0
cc_149 N_C1_M1012_g N_A_114_125#_c_450_n 0.00231577f $X=0.495 $Y=0.945 $X2=0
+ $Y2=0
cc_150 C1 N_A_114_125#_c_450_n 0.0209693f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_151 N_C1_c_144_n N_A_114_125#_c_450_n 0.00242321f $X=0.955 $Y=1.61 $X2=0
+ $Y2=0
cc_152 N_C1_M1014_g N_A_114_125#_c_451_n 0.00411919f $X=0.925 $Y=0.945 $X2=0
+ $Y2=0
cc_153 C1 N_A_114_125#_c_451_n 0.026566f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_154 N_C1_c_144_n N_A_114_125#_c_451_n 0.00715063f $X=0.955 $Y=1.61 $X2=0
+ $Y2=0
cc_155 N_C1_M1015_g N_A_114_125#_c_474_n 0.00259641f $X=0.505 $Y=2.435 $X2=0
+ $Y2=0
cc_156 N_C1_M1016_g N_A_114_125#_c_474_n 0.0161623f $X=0.955 $Y=2.435 $X2=0
+ $Y2=0
cc_157 C1 N_A_114_125#_c_474_n 0.020797f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_158 N_C1_c_144_n N_A_114_125#_c_474_n 6.24812e-19 $X=0.955 $Y=1.61 $X2=0
+ $Y2=0
cc_159 N_C1_M1015_g N_VPWR_c_619_n 0.00505401f $X=0.505 $Y=2.435 $X2=0 $Y2=0
cc_160 C1 N_VPWR_c_619_n 0.02049f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_161 N_C1_c_144_n N_VPWR_c_619_n 0.00110779f $X=0.955 $Y=1.61 $X2=0 $Y2=0
cc_162 N_C1_M1016_g N_VPWR_c_620_n 0.003011f $X=0.955 $Y=2.435 $X2=0 $Y2=0
cc_163 N_C1_M1015_g N_VPWR_c_626_n 0.00640648f $X=0.505 $Y=2.435 $X2=0 $Y2=0
cc_164 N_C1_M1016_g N_VPWR_c_626_n 0.00640648f $X=0.955 $Y=2.435 $X2=0 $Y2=0
cc_165 N_C1_M1015_g N_VPWR_c_617_n 0.00645424f $X=0.505 $Y=2.435 $X2=0 $Y2=0
cc_166 N_C1_M1016_g N_VPWR_c_617_n 0.00645424f $X=0.955 $Y=2.435 $X2=0 $Y2=0
cc_167 N_C1_M1012_g N_A_27_125#_c_828_n 0.00376028f $X=0.495 $Y=0.945 $X2=0
+ $Y2=0
cc_168 C1 N_A_27_125#_c_828_n 0.0205694f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_169 N_C1_c_144_n N_A_27_125#_c_828_n 0.00335457f $X=0.955 $Y=1.61 $X2=0 $Y2=0
cc_170 N_C1_M1012_g N_A_27_125#_c_829_n 0.00661564f $X=0.495 $Y=0.945 $X2=0
+ $Y2=0
cc_171 N_C1_M1014_g N_A_27_125#_c_829_n 0.00448896f $X=0.925 $Y=0.945 $X2=0
+ $Y2=0
cc_172 N_C1_M1012_g N_A_27_125#_c_831_n 4.41984e-19 $X=0.495 $Y=0.945 $X2=0
+ $Y2=0
cc_173 N_C1_M1014_g N_A_27_125#_c_831_n 0.00781575f $X=0.925 $Y=0.945 $X2=0
+ $Y2=0
cc_174 N_C1_M1014_g N_A_300_125#_c_896_n 5.16104e-19 $X=0.925 $Y=0.945 $X2=0
+ $Y2=0
cc_175 N_C1_M1014_g N_A_300_125#_c_897_n 4.39727e-19 $X=0.925 $Y=0.945 $X2=0
+ $Y2=0
cc_176 N_C1_M1014_g N_VGND_c_975_n 2.28708e-19 $X=0.925 $Y=0.945 $X2=0 $Y2=0
cc_177 N_B2_c_189_n N_B1_c_233_n 0.0162786f $X=2.355 $Y=1.61 $X2=-0.19
+ $Y2=-0.245
cc_178 N_B2_M1019_g N_B1_M1008_g 0.0162786f $X=1.905 $Y=2.435 $X2=0 $Y2=0
cc_179 B2 N_B1_M1008_g 0.00133285f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_180 N_B2_M1004_g N_B1_M1001_g 0.0162786f $X=1.89 $Y=0.945 $X2=0 $Y2=0
cc_181 N_B2_M1004_g N_B1_c_236_n 0.00737233f $X=1.89 $Y=0.945 $X2=0 $Y2=0
cc_182 N_B2_M1025_g N_B1_c_236_n 0.00737481f $X=2.355 $Y=0.945 $X2=0 $Y2=0
cc_183 N_B2_M1025_g N_B1_M1011_g 0.0140397f $X=2.355 $Y=0.945 $X2=0 $Y2=0
cc_184 N_B2_M1021_g N_B1_M1023_g 0.0221343f $X=2.355 $Y=2.435 $X2=0 $Y2=0
cc_185 B2 N_B1_M1023_g 0.00505672f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_186 B2 N_B1_c_241_n 0.00550809f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_187 N_B2_c_189_n N_B1_c_241_n 0.0221343f $X=2.355 $Y=1.61 $X2=0 $Y2=0
cc_188 B2 B1 0.0215428f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_189 N_B2_M1019_g N_A_114_125#_c_478_n 0.017215f $X=1.905 $Y=2.435 $X2=0 $Y2=0
cc_190 N_B2_M1021_g N_A_114_125#_c_479_n 0.0142175f $X=2.355 $Y=2.435 $X2=0
+ $Y2=0
cc_191 B2 N_A_114_125#_c_479_n 0.0347148f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_192 B2 N_A_114_125#_c_481_n 0.0141251f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_193 N_B2_c_189_n N_A_114_125#_c_481_n 7.03681e-19 $X=2.355 $Y=1.61 $X2=0
+ $Y2=0
cc_194 N_B2_M1019_g N_VPWR_c_620_n 2.41446e-19 $X=1.905 $Y=2.435 $X2=0 $Y2=0
cc_195 N_B2_M1019_g N_VPWR_c_627_n 0.00115241f $X=1.905 $Y=2.435 $X2=0 $Y2=0
cc_196 N_B2_M1021_g N_VPWR_c_627_n 0.00115241f $X=2.355 $Y=2.435 $X2=0 $Y2=0
cc_197 N_B2_M1019_g N_A_300_387#_c_714_n 0.00892729f $X=1.905 $Y=2.435 $X2=0
+ $Y2=0
cc_198 N_B2_M1021_g N_A_300_387#_c_714_n 5.73047e-19 $X=2.355 $Y=2.435 $X2=0
+ $Y2=0
cc_199 N_B2_M1019_g N_A_300_387#_c_712_n 0.0127415f $X=1.905 $Y=2.435 $X2=0
+ $Y2=0
cc_200 N_B2_M1021_g N_A_300_387#_c_712_n 0.0150734f $X=2.355 $Y=2.435 $X2=0
+ $Y2=0
cc_201 N_B2_M1019_g N_A_300_387#_c_713_n 0.00231365f $X=1.905 $Y=2.435 $X2=0
+ $Y2=0
cc_202 N_B2_M1019_g N_A_300_387#_c_719_n 5.73047e-19 $X=1.905 $Y=2.435 $X2=0
+ $Y2=0
cc_203 N_B2_M1021_g N_A_300_387#_c_719_n 0.00892729f $X=2.355 $Y=2.435 $X2=0
+ $Y2=0
cc_204 N_B2_M1004_g N_A_27_125#_c_832_n 0.00197096f $X=1.89 $Y=0.945 $X2=0 $Y2=0
cc_205 N_B2_M1004_g N_A_27_125#_c_833_n 0.00196596f $X=1.89 $Y=0.945 $X2=0 $Y2=0
cc_206 N_B2_M1025_g N_A_27_125#_c_833_n 0.00667575f $X=2.355 $Y=0.945 $X2=0
+ $Y2=0
cc_207 N_B2_M1025_g N_A_27_125#_c_834_n 0.00167488f $X=2.355 $Y=0.945 $X2=0
+ $Y2=0
cc_208 N_B2_M1025_g N_A_27_125#_c_835_n 4.53441e-19 $X=2.355 $Y=0.945 $X2=0
+ $Y2=0
cc_209 N_B2_M1004_g N_A_300_125#_c_896_n 2.9258e-19 $X=1.89 $Y=0.945 $X2=0 $Y2=0
cc_210 N_B2_M1004_g N_A_300_125#_c_898_n 0.0149567f $X=1.89 $Y=0.945 $X2=0 $Y2=0
cc_211 N_B2_M1025_g N_A_300_125#_c_898_n 0.0122769f $X=2.355 $Y=0.945 $X2=0
+ $Y2=0
cc_212 B2 N_A_300_125#_c_898_n 0.0328248f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_213 N_B2_c_189_n N_A_300_125#_c_898_n 0.00363005f $X=2.355 $Y=1.61 $X2=0
+ $Y2=0
cc_214 B2 N_A_300_125#_c_899_n 0.0010386f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_215 B2 N_A_300_125#_c_902_n 0.0227277f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_216 B1 N_A2_M1007_g 9.30501e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_217 B1 A2 0.0265558f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_218 B1 N_A2_c_321_n 0.0117853f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_219 B1 N_A1_M1013_g 0.0146519f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_220 N_B1_c_240_n N_A1_M1006_g 0.0160145f $X=3.3 $Y=1.445 $X2=0 $Y2=0
cc_221 N_B1_c_236_n N_A1_c_369_n 0.0160145f $X=3.225 $Y=0.18 $X2=0 $Y2=0
cc_222 N_B1_c_240_n N_A1_c_371_n 0.00776698f $X=3.3 $Y=1.445 $X2=0 $Y2=0
cc_223 B1 N_A1_c_371_n 0.00456294f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_224 N_B1_c_244_n N_A1_c_371_n 0.0207512f $X=3.3 $Y=1.61 $X2=0 $Y2=0
cc_225 N_B1_M1008_g N_A_114_125#_c_458_n 9.59636e-19 $X=1.41 $Y=2.435 $X2=0
+ $Y2=0
cc_226 N_B1_M1001_g N_A_114_125#_c_449_n 0.00155158f $X=1.425 $Y=0.945 $X2=0
+ $Y2=0
cc_227 N_B1_c_233_n N_A_114_125#_c_451_n 0.0140456f $X=1.41 $Y=1.43 $X2=0 $Y2=0
cc_228 N_B1_M1001_g N_A_114_125#_c_451_n 0.00132407f $X=1.425 $Y=0.945 $X2=0
+ $Y2=0
cc_229 N_B1_M1008_g N_A_114_125#_c_478_n 0.0216983f $X=1.41 $Y=2.435 $X2=0 $Y2=0
cc_230 N_B1_M1023_g N_A_114_125#_c_479_n 0.0205002f $X=2.805 $Y=2.435 $X2=0
+ $Y2=0
cc_231 B1 N_A_114_125#_c_479_n 0.0850278f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_232 N_B1_c_243_n N_A_114_125#_c_479_n 0.00259684f $X=3.105 $Y=1.61 $X2=0
+ $Y2=0
cc_233 N_B1_c_244_n N_A_114_125#_c_479_n 0.00227385f $X=3.3 $Y=1.61 $X2=0 $Y2=0
cc_234 N_B1_M1008_g N_VPWR_c_620_n 0.0104513f $X=1.41 $Y=2.435 $X2=0 $Y2=0
cc_235 N_B1_M1023_g N_VPWR_c_621_n 0.00323248f $X=2.805 $Y=2.435 $X2=0 $Y2=0
cc_236 N_B1_M1008_g N_VPWR_c_627_n 0.00577018f $X=1.41 $Y=2.435 $X2=0 $Y2=0
cc_237 N_B1_M1023_g N_VPWR_c_627_n 0.00578564f $X=2.805 $Y=2.435 $X2=0 $Y2=0
cc_238 N_B1_M1008_g N_VPWR_c_617_n 0.00559367f $X=1.41 $Y=2.435 $X2=0 $Y2=0
cc_239 N_B1_M1023_g N_VPWR_c_617_n 0.00537853f $X=2.805 $Y=2.435 $X2=0 $Y2=0
cc_240 N_B1_M1023_g N_A_300_387#_c_712_n 0.00378099f $X=2.805 $Y=2.435 $X2=0
+ $Y2=0
cc_241 N_B1_M1008_g N_A_300_387#_c_713_n 0.00123098f $X=1.41 $Y=2.435 $X2=0
+ $Y2=0
cc_242 N_B1_M1023_g N_A_300_387#_c_719_n 0.00761611f $X=2.805 $Y=2.435 $X2=0
+ $Y2=0
cc_243 N_B1_M1001_g N_A_27_125#_c_831_n 0.00528809f $X=1.425 $Y=0.945 $X2=0
+ $Y2=0
cc_244 N_B1_M1001_g N_A_27_125#_c_832_n 0.0177276f $X=1.425 $Y=0.945 $X2=0 $Y2=0
cc_245 N_B1_c_236_n N_A_27_125#_c_832_n 0.00657408f $X=3.225 $Y=0.18 $X2=0 $Y2=0
cc_246 N_B1_M1001_g N_A_27_125#_c_833_n 9.16073e-19 $X=1.425 $Y=0.945 $X2=0
+ $Y2=0
cc_247 N_B1_M1011_g N_A_27_125#_c_833_n 4.53441e-19 $X=2.79 $Y=0.945 $X2=0 $Y2=0
cc_248 N_B1_c_236_n N_A_27_125#_c_834_n 0.0151295f $X=3.225 $Y=0.18 $X2=0 $Y2=0
cc_249 N_B1_M1011_g N_A_27_125#_c_834_n 0.00175679f $X=2.79 $Y=0.945 $X2=0 $Y2=0
cc_250 N_B1_c_240_n N_A_27_125#_c_834_n 0.00273287f $X=3.3 $Y=1.445 $X2=0 $Y2=0
cc_251 N_B1_M1011_g N_A_27_125#_c_835_n 0.00686346f $X=2.79 $Y=0.945 $X2=0 $Y2=0
cc_252 N_B1_c_240_n N_A_27_125#_c_835_n 0.00454226f $X=3.3 $Y=1.445 $X2=0 $Y2=0
cc_253 N_B1_M1001_g N_A_27_125#_c_837_n 3.62868e-19 $X=1.425 $Y=0.945 $X2=0
+ $Y2=0
cc_254 N_B1_c_236_n N_A_27_125#_c_837_n 0.00766105f $X=3.225 $Y=0.18 $X2=0 $Y2=0
cc_255 N_B1_M1001_g N_A_300_125#_c_896_n 0.00477879f $X=1.425 $Y=0.945 $X2=0
+ $Y2=0
cc_256 N_B1_M1001_g N_A_300_125#_c_897_n 0.00564861f $X=1.425 $Y=0.945 $X2=0
+ $Y2=0
cc_257 N_B1_M1011_g N_A_300_125#_c_899_n 0.0108083f $X=2.79 $Y=0.945 $X2=0 $Y2=0
cc_258 N_B1_c_240_n N_A_300_125#_c_899_n 0.0158987f $X=3.3 $Y=1.445 $X2=0 $Y2=0
cc_259 B1 N_A_300_125#_c_899_n 0.0702714f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_260 N_B1_c_243_n N_A_300_125#_c_899_n 0.00376758f $X=3.105 $Y=1.61 $X2=0
+ $Y2=0
cc_261 N_B1_c_244_n N_A_300_125#_c_899_n 0.00134523f $X=3.3 $Y=1.61 $X2=0 $Y2=0
cc_262 B1 N_A_300_125#_c_920_n 0.00272347f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_263 N_B1_M1011_g N_A_300_125#_c_902_n 0.00310616f $X=2.79 $Y=0.945 $X2=0
+ $Y2=0
cc_264 N_B1_c_240_n N_A_300_125#_c_902_n 3.73248e-19 $X=3.3 $Y=1.445 $X2=0 $Y2=0
cc_265 B1 N_A_300_125#_c_903_n 0.0155152f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_266 N_B1_c_236_n N_VGND_c_965_n 0.01258f $X=3.225 $Y=0.18 $X2=0 $Y2=0
cc_267 N_B1_c_237_n N_VGND_c_975_n 0.0461037f $X=1.5 $Y=0.18 $X2=0 $Y2=0
cc_268 N_B1_c_236_n N_VGND_c_980_n 0.0526956f $X=3.225 $Y=0.18 $X2=0 $Y2=0
cc_269 N_B1_c_237_n N_VGND_c_980_n 0.00604685f $X=1.5 $Y=0.18 $X2=0 $Y2=0
cc_270 N_A2_c_321_n N_A1_M1013_g 0.0391913f $X=4.675 $Y=1.61 $X2=0 $Y2=0
cc_271 N_A2_M1009_g N_A1_M1006_g 0.0153432f $X=4.245 $Y=0.915 $X2=0 $Y2=0
cc_272 N_A2_M1009_g N_A1_c_368_n 0.0103107f $X=4.245 $Y=0.915 $X2=0 $Y2=0
cc_273 N_A2_M1010_g N_A1_c_368_n 0.0103107f $X=4.675 $Y=0.915 $X2=0 $Y2=0
cc_274 N_A2_M1010_g N_A1_M1018_g 0.0111633f $X=4.675 $Y=0.915 $X2=0 $Y2=0
cc_275 N_A2_c_321_n N_A1_M1024_g 0.0270732f $X=4.675 $Y=1.61 $X2=0 $Y2=0
cc_276 N_A2_c_321_n N_A1_c_371_n 8.38744e-19 $X=4.675 $Y=1.61 $X2=0 $Y2=0
cc_277 N_A2_M1010_g N_A1_c_372_n 0.0130117f $X=4.675 $Y=0.915 $X2=0 $Y2=0
cc_278 A2 N_A1_c_372_n 2.40741e-19 $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_279 N_A2_c_321_n N_A1_c_372_n 0.00557182f $X=4.675 $Y=1.61 $X2=0 $Y2=0
cc_280 N_A2_M1010_g N_A1_c_373_n 0.0033787f $X=4.675 $Y=0.915 $X2=0 $Y2=0
cc_281 A2 N_A1_c_373_n 0.0214356f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_282 N_A2_c_321_n N_A1_c_373_n 0.00154554f $X=4.675 $Y=1.61 $X2=0 $Y2=0
cc_283 N_A2_M1007_g N_A_114_125#_c_479_n 0.0178828f $X=4.215 $Y=2.435 $X2=0
+ $Y2=0
cc_284 N_A2_M1017_g N_A_114_125#_c_493_n 0.0156925f $X=4.69 $Y=2.435 $X2=0 $Y2=0
cc_285 A2 N_A_114_125#_c_493_n 0.00456582f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_286 N_A2_M1007_g N_A_114_125#_c_495_n 0.0106162f $X=4.215 $Y=2.435 $X2=0
+ $Y2=0
cc_287 N_A2_M1017_g N_A_114_125#_c_495_n 0.011221f $X=4.69 $Y=2.435 $X2=0 $Y2=0
cc_288 A2 N_A_114_125#_c_495_n 0.0202023f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_289 N_A2_c_321_n N_A_114_125#_c_495_n 8.95858e-19 $X=4.675 $Y=1.61 $X2=0
+ $Y2=0
cc_290 N_A2_M1007_g N_VPWR_c_628_n 0.00115264f $X=4.215 $Y=2.435 $X2=0 $Y2=0
cc_291 N_A2_M1017_g N_VPWR_c_628_n 0.00113339f $X=4.69 $Y=2.435 $X2=0 $Y2=0
cc_292 N_A2_M1007_g N_A_766_387#_c_738_n 0.00928566f $X=4.215 $Y=2.435 $X2=0
+ $Y2=0
cc_293 N_A2_M1017_g N_A_766_387#_c_738_n 4.61476e-19 $X=4.69 $Y=2.435 $X2=0
+ $Y2=0
cc_294 N_A2_M1007_g N_A_766_387#_c_736_n 0.0145385f $X=4.215 $Y=2.435 $X2=0
+ $Y2=0
cc_295 N_A2_M1017_g N_A_766_387#_c_736_n 0.0159033f $X=4.69 $Y=2.435 $X2=0 $Y2=0
cc_296 N_A2_M1007_g N_A_766_387#_c_737_n 0.00171894f $X=4.215 $Y=2.435 $X2=0
+ $Y2=0
cc_297 N_A2_M1009_g N_A_300_125#_c_920_n 0.0158989f $X=4.245 $Y=0.915 $X2=0
+ $Y2=0
cc_298 N_A2_M1010_g N_A_300_125#_c_920_n 0.0139892f $X=4.675 $Y=0.915 $X2=0
+ $Y2=0
cc_299 A2 N_A_300_125#_c_920_n 0.015287f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_300 N_A2_c_321_n N_A_300_125#_c_920_n 6.42129e-19 $X=4.675 $Y=1.61 $X2=0
+ $Y2=0
cc_301 N_A2_M1009_g N_A_300_125#_c_903_n 0.00124096f $X=4.245 $Y=0.915 $X2=0
+ $Y2=0
cc_302 N_A2_M1009_g N_VGND_c_965_n 4.57735e-19 $X=4.245 $Y=0.915 $X2=0 $Y2=0
cc_303 N_A2_M1009_g N_VGND_c_966_n 0.00680324f $X=4.245 $Y=0.915 $X2=0 $Y2=0
cc_304 N_A2_M1010_g N_VGND_c_966_n 0.00702747f $X=4.675 $Y=0.915 $X2=0 $Y2=0
cc_305 N_A2_M1009_g N_VGND_c_980_n 7.88961e-19 $X=4.245 $Y=0.915 $X2=0 $Y2=0
cc_306 N_A2_M1010_g N_VGND_c_980_n 7.88961e-19 $X=4.675 $Y=0.915 $X2=0 $Y2=0
cc_307 N_A1_M1018_g N_A_114_125#_c_441_n 0.0210564f $X=5.105 $Y=0.915 $X2=0
+ $Y2=0
cc_308 N_A1_M1024_g N_A_114_125#_M1000_g 0.0236947f $X=5.19 $Y=2.435 $X2=0 $Y2=0
cc_309 N_A1_c_373_n N_A_114_125#_M1000_g 2.85661e-19 $X=5.155 $Y=1.515 $X2=0
+ $Y2=0
cc_310 N_A1_M1013_g N_A_114_125#_c_479_n 0.0185061f $X=3.74 $Y=2.435 $X2=0 $Y2=0
cc_311 N_A1_M1024_g N_A_114_125#_c_493_n 0.0167879f $X=5.19 $Y=2.435 $X2=0 $Y2=0
cc_312 N_A1_c_372_n N_A_114_125#_c_493_n 4.91416e-19 $X=5.155 $Y=1.515 $X2=0
+ $Y2=0
cc_313 N_A1_c_373_n N_A_114_125#_c_493_n 0.0267438f $X=5.155 $Y=1.515 $X2=0
+ $Y2=0
cc_314 N_A1_M1024_g N_A_114_125#_c_460_n 0.00372702f $X=5.19 $Y=2.435 $X2=0
+ $Y2=0
cc_315 N_A1_c_373_n N_A_114_125#_c_460_n 0.00800366f $X=5.155 $Y=1.515 $X2=0
+ $Y2=0
cc_316 N_A1_c_372_n N_A_114_125#_c_452_n 0.00234848f $X=5.155 $Y=1.515 $X2=0
+ $Y2=0
cc_317 N_A1_c_373_n N_A_114_125#_c_452_n 0.028177f $X=5.155 $Y=1.515 $X2=0 $Y2=0
cc_318 N_A1_M1013_g N_A_114_125#_c_495_n 6.17306e-19 $X=3.74 $Y=2.435 $X2=0
+ $Y2=0
cc_319 N_A1_M1024_g N_A_114_125#_c_495_n 6.3351e-19 $X=5.19 $Y=2.435 $X2=0 $Y2=0
cc_320 N_A1_c_372_n N_A_114_125#_c_453_n 0.0139319f $X=5.155 $Y=1.515 $X2=0
+ $Y2=0
cc_321 N_A1_c_373_n N_A_114_125#_c_453_n 3.39156e-19 $X=5.155 $Y=1.515 $X2=0
+ $Y2=0
cc_322 N_A1_M1013_g N_VPWR_c_621_n 0.00323248f $X=3.74 $Y=2.435 $X2=0 $Y2=0
cc_323 N_A1_M1024_g N_VPWR_c_622_n 0.00114594f $X=5.19 $Y=2.435 $X2=0 $Y2=0
cc_324 N_A1_M1013_g N_VPWR_c_628_n 0.00578564f $X=3.74 $Y=2.435 $X2=0 $Y2=0
cc_325 N_A1_M1024_g N_VPWR_c_628_n 0.00578564f $X=5.19 $Y=2.435 $X2=0 $Y2=0
cc_326 N_A1_M1013_g N_VPWR_c_617_n 0.00537853f $X=3.74 $Y=2.435 $X2=0 $Y2=0
cc_327 N_A1_M1024_g N_VPWR_c_617_n 0.00537853f $X=5.19 $Y=2.435 $X2=0 $Y2=0
cc_328 N_A1_M1013_g N_A_766_387#_c_738_n 0.00761611f $X=3.74 $Y=2.435 $X2=0
+ $Y2=0
cc_329 N_A1_M1024_g N_A_766_387#_c_736_n 0.00392636f $X=5.19 $Y=2.435 $X2=0
+ $Y2=0
cc_330 N_A1_M1013_g N_A_766_387#_c_737_n 0.00389438f $X=3.74 $Y=2.435 $X2=0
+ $Y2=0
cc_331 N_A1_M1024_g N_A_766_387#_c_746_n 0.00732993f $X=5.19 $Y=2.435 $X2=0
+ $Y2=0
cc_332 N_A1_M1006_g N_A_300_125#_c_899_n 0.0130111f $X=3.81 $Y=0.915 $X2=0 $Y2=0
cc_333 N_A1_c_371_n N_A_300_125#_c_899_n 0.00262703f $X=3.767 $Y=1.46 $X2=0
+ $Y2=0
cc_334 N_A1_c_368_n N_A_300_125#_c_900_n 0.0027941f $X=5.03 $Y=0.18 $X2=0 $Y2=0
cc_335 N_A1_M1018_g N_A_300_125#_c_932_n 0.00213302f $X=5.105 $Y=0.915 $X2=0
+ $Y2=0
cc_336 N_A1_c_373_n N_A_300_125#_c_932_n 0.00843415f $X=5.155 $Y=1.515 $X2=0
+ $Y2=0
cc_337 N_A1_c_368_n N_A_300_125#_c_901_n 0.0026558f $X=5.03 $Y=0.18 $X2=0 $Y2=0
cc_338 N_A1_M1018_g N_A_300_125#_c_901_n 0.00494004f $X=5.105 $Y=0.915 $X2=0
+ $Y2=0
cc_339 N_A1_M1006_g N_VGND_c_965_n 0.0143118f $X=3.81 $Y=0.915 $X2=0 $Y2=0
cc_340 N_A1_c_369_n N_VGND_c_965_n 0.00541156f $X=3.885 $Y=0.18 $X2=0 $Y2=0
cc_341 N_A1_M1006_g N_VGND_c_966_n 0.00412296f $X=3.81 $Y=0.915 $X2=0 $Y2=0
cc_342 N_A1_c_368_n N_VGND_c_966_n 0.0232758f $X=5.03 $Y=0.18 $X2=0 $Y2=0
cc_343 N_A1_M1018_g N_VGND_c_966_n 0.00428233f $X=5.105 $Y=0.915 $X2=0 $Y2=0
cc_344 N_A1_c_368_n N_VGND_c_967_n 0.0144414f $X=5.03 $Y=0.18 $X2=0 $Y2=0
cc_345 N_A1_c_372_n N_VGND_c_967_n 6.49736e-19 $X=5.155 $Y=1.515 $X2=0 $Y2=0
cc_346 N_A1_c_373_n N_VGND_c_967_n 0.00697284f $X=5.155 $Y=1.515 $X2=0 $Y2=0
cc_347 N_A1_c_369_n N_VGND_c_971_n 0.0176917f $X=3.885 $Y=0.18 $X2=0 $Y2=0
cc_348 N_A1_c_368_n N_VGND_c_973_n 0.0176813f $X=5.03 $Y=0.18 $X2=0 $Y2=0
cc_349 N_A1_c_368_n N_VGND_c_980_n 0.0384141f $X=5.03 $Y=0.18 $X2=0 $Y2=0
cc_350 N_A1_c_369_n N_VGND_c_980_n 0.00749832f $X=3.885 $Y=0.18 $X2=0 $Y2=0
cc_351 N_A_114_125#_c_451_n N_VPWR_M1016_s 5.42186e-19 $X=1.145 $Y=1.95 $X2=0
+ $Y2=0
cc_352 N_A_114_125#_c_478_n N_VPWR_M1016_s 0.00156114f $X=2.045 $Y=2.035 $X2=0
+ $Y2=0
cc_353 N_A_114_125#_c_474_n N_VPWR_M1016_s 0.00172556f $X=1.23 $Y=2.035 $X2=0
+ $Y2=0
cc_354 N_A_114_125#_c_479_n N_VPWR_M1023_s 0.0166081f $X=4.3 $Y=2.035 $X2=0
+ $Y2=0
cc_355 N_A_114_125#_c_493_n N_VPWR_M1024_s 0.00804621f $X=5.49 $Y=2.035 $X2=0
+ $Y2=0
cc_356 N_A_114_125#_c_460_n N_VPWR_M1024_s 0.00130078f $X=5.575 $Y=1.95 $X2=0
+ $Y2=0
cc_357 N_A_114_125#_c_458_n N_VPWR_c_619_n 0.0281854f $X=0.73 $Y=2.79 $X2=0
+ $Y2=0
cc_358 N_A_114_125#_c_458_n N_VPWR_c_620_n 0.0225847f $X=0.73 $Y=2.79 $X2=0
+ $Y2=0
cc_359 N_A_114_125#_c_474_n N_VPWR_c_620_n 0.0148119f $X=1.23 $Y=2.035 $X2=0
+ $Y2=0
cc_360 N_A_114_125#_c_479_n N_VPWR_c_621_n 0.0521508f $X=4.3 $Y=2.035 $X2=0
+ $Y2=0
cc_361 N_A_114_125#_M1000_g N_VPWR_c_622_n 0.0127792f $X=5.695 $Y=2.4 $X2=0
+ $Y2=0
cc_362 N_A_114_125#_M1003_g N_VPWR_c_622_n 7.06477e-19 $X=6.22 $Y=2.4 $X2=0
+ $Y2=0
cc_363 N_A_114_125#_c_493_n N_VPWR_c_622_n 0.019585f $X=5.49 $Y=2.035 $X2=0
+ $Y2=0
cc_364 N_A_114_125#_M1003_g N_VPWR_c_623_n 0.00327951f $X=6.22 $Y=2.4 $X2=0
+ $Y2=0
cc_365 N_A_114_125#_M1020_g N_VPWR_c_623_n 0.0138991f $X=6.67 $Y=2.4 $X2=0 $Y2=0
cc_366 N_A_114_125#_M1026_g N_VPWR_c_623_n 7.44604e-19 $X=7.175 $Y=2.4 $X2=0
+ $Y2=0
cc_367 N_A_114_125#_M1026_g N_VPWR_c_625_n 0.00501904f $X=7.175 $Y=2.4 $X2=0
+ $Y2=0
cc_368 N_A_114_125#_c_458_n N_VPWR_c_626_n 0.013132f $X=0.73 $Y=2.79 $X2=0 $Y2=0
cc_369 N_A_114_125#_M1000_g N_VPWR_c_629_n 0.00475445f $X=5.695 $Y=2.4 $X2=0
+ $Y2=0
cc_370 N_A_114_125#_M1003_g N_VPWR_c_629_n 0.005209f $X=6.22 $Y=2.4 $X2=0 $Y2=0
cc_371 N_A_114_125#_M1020_g N_VPWR_c_630_n 0.00460063f $X=6.67 $Y=2.4 $X2=0
+ $Y2=0
cc_372 N_A_114_125#_M1026_g N_VPWR_c_630_n 0.005209f $X=7.175 $Y=2.4 $X2=0 $Y2=0
cc_373 N_A_114_125#_M1000_g N_VPWR_c_617_n 0.00939376f $X=5.695 $Y=2.4 $X2=0
+ $Y2=0
cc_374 N_A_114_125#_M1003_g N_VPWR_c_617_n 0.00982981f $X=6.22 $Y=2.4 $X2=0
+ $Y2=0
cc_375 N_A_114_125#_M1020_g N_VPWR_c_617_n 0.00909089f $X=6.67 $Y=2.4 $X2=0
+ $Y2=0
cc_376 N_A_114_125#_M1026_g N_VPWR_c_617_n 0.00986542f $X=7.175 $Y=2.4 $X2=0
+ $Y2=0
cc_377 N_A_114_125#_c_458_n N_VPWR_c_617_n 0.0118799f $X=0.73 $Y=2.79 $X2=0
+ $Y2=0
cc_378 N_A_114_125#_c_478_n N_A_300_387#_M1008_d 0.00635864f $X=2.045 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_379 N_A_114_125#_c_479_n N_A_300_387#_M1021_s 0.00332066f $X=4.3 $Y=2.035
+ $X2=0 $Y2=0
cc_380 N_A_114_125#_c_478_n N_A_300_387#_c_714_n 0.01852f $X=2.045 $Y=2.035
+ $X2=0 $Y2=0
cc_381 N_A_114_125#_M1019_d N_A_300_387#_c_712_n 0.00165831f $X=1.995 $Y=1.935
+ $X2=0 $Y2=0
cc_382 N_A_114_125#_c_481_n N_A_300_387#_c_712_n 0.0118736f $X=2.13 $Y=2.115
+ $X2=0 $Y2=0
cc_383 N_A_114_125#_c_479_n N_A_300_387#_c_719_n 0.0170259f $X=4.3 $Y=2.035
+ $X2=0 $Y2=0
cc_384 N_A_114_125#_c_479_n N_A_766_387#_M1013_d 0.00385282f $X=4.3 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_385 N_A_114_125#_c_493_n N_A_766_387#_M1017_s 0.00672557f $X=5.49 $Y=2.035
+ $X2=0 $Y2=0
cc_386 N_A_114_125#_c_479_n N_A_766_387#_c_738_n 0.0171554f $X=4.3 $Y=2.035
+ $X2=0 $Y2=0
cc_387 N_A_114_125#_c_495_n N_A_766_387#_c_738_n 0.0333949f $X=4.465 $Y=2.115
+ $X2=0 $Y2=0
cc_388 N_A_114_125#_M1007_d N_A_766_387#_c_736_n 0.00192406f $X=4.305 $Y=1.935
+ $X2=0 $Y2=0
cc_389 N_A_114_125#_c_495_n N_A_766_387#_c_736_n 0.0160534f $X=4.465 $Y=2.115
+ $X2=0 $Y2=0
cc_390 N_A_114_125#_c_493_n N_A_766_387#_c_746_n 0.0189268f $X=5.49 $Y=2.035
+ $X2=0 $Y2=0
cc_391 N_A_114_125#_c_441_n N_X_c_760_n 0.00575016f $X=5.68 $Y=1.35 $X2=0 $Y2=0
cc_392 N_A_114_125#_M1003_g N_X_c_770_n 8.84614e-19 $X=6.22 $Y=2.4 $X2=0 $Y2=0
cc_393 N_A_114_125#_c_556_p N_X_c_770_n 0.0240302f $X=6.45 $Y=1.515 $X2=0 $Y2=0
cc_394 N_A_114_125#_c_453_n N_X_c_770_n 0.00419876f $X=6.76 $Y=1.515 $X2=0 $Y2=0
cc_395 N_A_114_125#_M1000_g N_X_c_765_n 0.00522625f $X=5.695 $Y=2.4 $X2=0 $Y2=0
cc_396 N_A_114_125#_M1003_g N_X_c_765_n 0.0135076f $X=6.22 $Y=2.4 $X2=0 $Y2=0
cc_397 N_A_114_125#_M1020_g N_X_c_765_n 7.3056e-19 $X=6.67 $Y=2.4 $X2=0 $Y2=0
cc_398 N_A_114_125#_c_442_n N_X_c_776_n 0.0128266f $X=6.115 $Y=1.35 $X2=0 $Y2=0
cc_399 N_A_114_125#_c_443_n N_X_c_776_n 0.013439f $X=6.685 $Y=1.35 $X2=0 $Y2=0
cc_400 N_A_114_125#_c_556_p N_X_c_776_n 0.0399707f $X=6.45 $Y=1.515 $X2=0 $Y2=0
cc_401 N_A_114_125#_c_453_n N_X_c_776_n 0.00597192f $X=6.76 $Y=1.515 $X2=0 $Y2=0
cc_402 N_A_114_125#_c_441_n N_X_c_780_n 0.00196505f $X=5.68 $Y=1.35 $X2=0 $Y2=0
cc_403 N_A_114_125#_c_556_p N_X_c_780_n 0.0179455f $X=6.45 $Y=1.515 $X2=0 $Y2=0
cc_404 N_A_114_125#_c_453_n N_X_c_780_n 0.00256284f $X=6.76 $Y=1.515 $X2=0 $Y2=0
cc_405 N_A_114_125#_M1003_g N_X_c_783_n 0.0128923f $X=6.22 $Y=2.4 $X2=0 $Y2=0
cc_406 N_A_114_125#_M1020_g N_X_c_783_n 0.0163784f $X=6.67 $Y=2.4 $X2=0 $Y2=0
cc_407 N_A_114_125#_c_556_p N_X_c_783_n 0.0289737f $X=6.45 $Y=1.515 $X2=0 $Y2=0
cc_408 N_A_114_125#_c_453_n N_X_c_783_n 0.00201785f $X=6.76 $Y=1.515 $X2=0 $Y2=0
cc_409 N_A_114_125#_c_442_n N_X_c_761_n 9.34645e-19 $X=6.115 $Y=1.35 $X2=0 $Y2=0
cc_410 N_A_114_125#_c_443_n N_X_c_761_n 0.00809381f $X=6.685 $Y=1.35 $X2=0 $Y2=0
cc_411 N_A_114_125#_c_445_n N_X_c_761_n 0.00622602f $X=7.115 $Y=1.35 $X2=0 $Y2=0
cc_412 N_A_114_125#_M1020_g N_X_c_766_n 4.39447e-19 $X=6.67 $Y=2.4 $X2=0 $Y2=0
cc_413 N_A_114_125#_M1026_g N_X_c_766_n 0.0130882f $X=7.175 $Y=2.4 $X2=0 $Y2=0
cc_414 N_A_114_125#_c_443_n N_X_c_792_n 0.00103753f $X=6.685 $Y=1.35 $X2=0 $Y2=0
cc_415 N_A_114_125#_c_445_n N_X_c_792_n 0.00181823f $X=7.115 $Y=1.35 $X2=0 $Y2=0
cc_416 N_A_114_125#_c_444_n N_X_c_762_n 0.00642043f $X=7.04 $Y=1.487 $X2=0 $Y2=0
cc_417 N_A_114_125#_M1026_g N_X_c_762_n 0.0117574f $X=7.175 $Y=2.4 $X2=0 $Y2=0
cc_418 N_A_114_125#_c_447_n N_X_c_762_n 0.00329975f $X=7.152 $Y=1.487 $X2=0
+ $Y2=0
cc_419 N_A_114_125#_c_453_n N_X_c_762_n 0.00521865f $X=6.76 $Y=1.515 $X2=0 $Y2=0
cc_420 N_A_114_125#_c_443_n N_X_c_763_n 0.00322108f $X=6.685 $Y=1.35 $X2=0 $Y2=0
cc_421 N_A_114_125#_c_444_n N_X_c_763_n 0.00995134f $X=7.04 $Y=1.487 $X2=0 $Y2=0
cc_422 N_A_114_125#_c_445_n N_X_c_763_n 0.00613906f $X=7.115 $Y=1.35 $X2=0 $Y2=0
cc_423 N_A_114_125#_c_447_n N_X_c_763_n 0.00867018f $X=7.152 $Y=1.487 $X2=0
+ $Y2=0
cc_424 N_A_114_125#_c_556_p N_X_c_763_n 0.0261795f $X=6.45 $Y=1.515 $X2=0 $Y2=0
cc_425 N_A_114_125#_M1026_g X 0.0128155f $X=7.175 $Y=2.4 $X2=0 $Y2=0
cc_426 N_A_114_125#_c_447_n X 0.00843911f $X=7.152 $Y=1.487 $X2=0 $Y2=0
cc_427 N_A_114_125#_c_449_n N_A_27_125#_M1014_d 0.00391046f $X=1.06 $Y=1.19
+ $X2=0 $Y2=0
cc_428 N_A_114_125#_c_448_n N_A_27_125#_c_828_n 0.0178678f $X=0.71 $Y=0.77 $X2=0
+ $Y2=0
cc_429 N_A_114_125#_c_450_n N_A_27_125#_c_828_n 0.00719222f $X=0.795 $Y=1.19
+ $X2=0 $Y2=0
cc_430 N_A_114_125#_c_448_n N_A_27_125#_c_829_n 0.0195166f $X=0.71 $Y=0.77 $X2=0
+ $Y2=0
cc_431 N_A_114_125#_c_449_n N_A_27_125#_c_829_n 0.00388263f $X=1.06 $Y=1.19
+ $X2=0 $Y2=0
cc_432 N_A_114_125#_c_448_n N_A_27_125#_c_831_n 0.0125556f $X=0.71 $Y=0.77 $X2=0
+ $Y2=0
cc_433 N_A_114_125#_c_449_n N_A_27_125#_c_831_n 0.0172289f $X=1.06 $Y=1.19 $X2=0
+ $Y2=0
cc_434 N_A_114_125#_c_449_n N_A_300_125#_c_896_n 0.0112178f $X=1.06 $Y=1.19
+ $X2=0 $Y2=0
cc_435 N_A_114_125#_c_451_n N_A_300_125#_c_896_n 5.44422e-19 $X=1.145 $Y=1.95
+ $X2=0 $Y2=0
cc_436 N_A_114_125#_c_478_n N_A_300_125#_c_896_n 0.00869791f $X=2.045 $Y=2.035
+ $X2=0 $Y2=0
cc_437 N_A_114_125#_c_478_n N_A_300_125#_c_898_n 0.0049714f $X=2.045 $Y=2.035
+ $X2=0 $Y2=0
cc_438 N_A_114_125#_c_479_n N_A_300_125#_c_899_n 0.00535038f $X=4.3 $Y=2.035
+ $X2=0 $Y2=0
cc_439 N_A_114_125#_c_441_n N_VGND_c_967_n 0.00618447f $X=5.68 $Y=1.35 $X2=0
+ $Y2=0
cc_440 N_A_114_125#_c_452_n N_VGND_c_967_n 0.0060815f $X=5.66 $Y=1.515 $X2=0
+ $Y2=0
cc_441 N_A_114_125#_c_441_n N_VGND_c_968_n 4.38995e-19 $X=5.68 $Y=1.35 $X2=0
+ $Y2=0
cc_442 N_A_114_125#_c_442_n N_VGND_c_968_n 0.00821436f $X=6.115 $Y=1.35 $X2=0
+ $Y2=0
cc_443 N_A_114_125#_c_443_n N_VGND_c_968_n 0.00394182f $X=6.685 $Y=1.35 $X2=0
+ $Y2=0
cc_444 N_A_114_125#_c_445_n N_VGND_c_970_n 0.0185143f $X=7.115 $Y=1.35 $X2=0
+ $Y2=0
cc_445 N_A_114_125#_c_447_n N_VGND_c_970_n 9.30454e-19 $X=7.152 $Y=1.487 $X2=0
+ $Y2=0
cc_446 N_A_114_125#_c_441_n N_VGND_c_976_n 0.00474666f $X=5.68 $Y=1.35 $X2=0
+ $Y2=0
cc_447 N_A_114_125#_c_442_n N_VGND_c_976_n 0.00407914f $X=6.115 $Y=1.35 $X2=0
+ $Y2=0
cc_448 N_A_114_125#_c_443_n N_VGND_c_977_n 0.00470409f $X=6.685 $Y=1.35 $X2=0
+ $Y2=0
cc_449 N_A_114_125#_c_445_n N_VGND_c_977_n 0.00470409f $X=7.115 $Y=1.35 $X2=0
+ $Y2=0
cc_450 N_A_114_125#_c_441_n N_VGND_c_980_n 0.00506877f $X=5.68 $Y=1.35 $X2=0
+ $Y2=0
cc_451 N_A_114_125#_c_442_n N_VGND_c_980_n 0.00425776f $X=6.115 $Y=1.35 $X2=0
+ $Y2=0
cc_452 N_A_114_125#_c_443_n N_VGND_c_980_n 0.00506877f $X=6.685 $Y=1.35 $X2=0
+ $Y2=0
cc_453 N_A_114_125#_c_445_n N_VGND_c_980_n 0.00506877f $X=7.115 $Y=1.35 $X2=0
+ $Y2=0
cc_454 N_VPWR_c_621_n N_A_300_387#_c_712_n 0.0137331f $X=3.515 $Y=2.455 $X2=0
+ $Y2=0
cc_455 N_VPWR_c_627_n N_A_300_387#_c_712_n 0.0603168f $X=2.915 $Y=3.33 $X2=0
+ $Y2=0
cc_456 N_VPWR_c_617_n N_A_300_387#_c_712_n 0.0342523f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_457 N_VPWR_c_620_n N_A_300_387#_c_713_n 0.012662f $X=1.18 $Y=2.455 $X2=0
+ $Y2=0
cc_458 N_VPWR_c_627_n N_A_300_387#_c_713_n 0.0236566f $X=2.915 $Y=3.33 $X2=0
+ $Y2=0
cc_459 N_VPWR_c_617_n N_A_300_387#_c_713_n 0.0128296f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_460 N_VPWR_c_622_n N_A_766_387#_c_736_n 0.0130139f $X=5.465 $Y=2.415 $X2=0
+ $Y2=0
cc_461 N_VPWR_c_628_n N_A_766_387#_c_736_n 0.0667586f $X=5.3 $Y=3.33 $X2=0 $Y2=0
cc_462 N_VPWR_c_617_n N_A_766_387#_c_736_n 0.0380121f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_463 N_VPWR_c_621_n N_A_766_387#_c_737_n 0.0137331f $X=3.515 $Y=2.455 $X2=0
+ $Y2=0
cc_464 N_VPWR_c_628_n N_A_766_387#_c_737_n 0.0236566f $X=5.3 $Y=3.33 $X2=0 $Y2=0
cc_465 N_VPWR_c_617_n N_A_766_387#_c_737_n 0.0128296f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_466 N_VPWR_c_622_n N_X_c_765_n 0.0234373f $X=5.465 $Y=2.415 $X2=0 $Y2=0
cc_467 N_VPWR_c_623_n N_X_c_765_n 0.0267028f $X=6.445 $Y=2.355 $X2=0 $Y2=0
cc_468 N_VPWR_c_629_n N_X_c_765_n 0.014549f $X=6.36 $Y=3.33 $X2=0 $Y2=0
cc_469 N_VPWR_c_617_n N_X_c_765_n 0.0119743f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_470 N_VPWR_M1003_s N_X_c_783_n 0.00311483f $X=6.31 $Y=1.84 $X2=0 $Y2=0
cc_471 N_VPWR_c_623_n N_X_c_783_n 0.0148589f $X=6.445 $Y=2.355 $X2=0 $Y2=0
cc_472 N_VPWR_c_623_n N_X_c_766_n 0.0285293f $X=6.445 $Y=2.355 $X2=0 $Y2=0
cc_473 N_VPWR_c_630_n N_X_c_766_n 0.014549f $X=7.315 $Y=3.33 $X2=0 $Y2=0
cc_474 N_VPWR_c_617_n N_X_c_766_n 0.0119743f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_475 N_VPWR_c_625_n N_X_c_762_n 0.0345768f $X=7.4 $Y=2.115 $X2=0 $Y2=0
cc_476 N_VPWR_c_625_n X 0.0199358f $X=7.4 $Y=2.115 $X2=0 $Y2=0
cc_477 N_VPWR_c_619_n N_A_27_125#_c_828_n 3.19761e-19 $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_478 N_X_c_776_n N_VGND_M1005_d 0.00676949f $X=6.735 $Y=1.095 $X2=0 $Y2=0
cc_479 N_X_c_760_n N_VGND_c_967_n 0.0199928f $X=5.9 $Y=0.64 $X2=0 $Y2=0
cc_480 N_X_c_760_n N_VGND_c_968_n 0.0129089f $X=5.9 $Y=0.64 $X2=0 $Y2=0
cc_481 N_X_c_776_n N_VGND_c_968_n 0.0231921f $X=6.735 $Y=1.095 $X2=0 $Y2=0
cc_482 N_X_c_761_n N_VGND_c_968_n 0.0131962f $X=6.9 $Y=0.64 $X2=0 $Y2=0
cc_483 N_X_c_761_n N_VGND_c_970_n 0.0208274f $X=6.9 $Y=0.64 $X2=0 $Y2=0
cc_484 N_X_c_763_n N_VGND_c_970_n 0.00349814f $X=6.95 $Y=1.55 $X2=0 $Y2=0
cc_485 X N_VGND_c_970_n 0.0186157f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_486 N_X_c_760_n N_VGND_c_976_n 0.0073038f $X=5.9 $Y=0.64 $X2=0 $Y2=0
cc_487 N_X_c_761_n N_VGND_c_977_n 0.00957956f $X=6.9 $Y=0.64 $X2=0 $Y2=0
cc_488 N_X_c_760_n N_VGND_c_980_n 0.00843588f $X=5.9 $Y=0.64 $X2=0 $Y2=0
cc_489 N_X_c_761_n N_VGND_c_980_n 0.0111194f $X=6.9 $Y=0.64 $X2=0 $Y2=0
cc_490 N_A_27_125#_c_831_n N_A_300_125#_c_897_n 0.0131729f $X=1.14 $Y=0.77 $X2=0
+ $Y2=0
cc_491 N_A_27_125#_c_832_n N_A_300_125#_c_897_n 0.0257832f $X=1.975 $Y=0.35
+ $X2=0 $Y2=0
cc_492 N_A_27_125#_c_833_n N_A_300_125#_c_897_n 0.00158095f $X=2.14 $Y=0.77
+ $X2=0 $Y2=0
cc_493 N_A_27_125#_M1004_s N_A_300_125#_c_898_n 0.00216221f $X=1.965 $Y=0.625
+ $X2=0 $Y2=0
cc_494 N_A_27_125#_c_832_n N_A_300_125#_c_898_n 0.00456055f $X=1.975 $Y=0.35
+ $X2=0 $Y2=0
cc_495 N_A_27_125#_c_833_n N_A_300_125#_c_898_n 0.0184164f $X=2.14 $Y=0.77 $X2=0
+ $Y2=0
cc_496 N_A_27_125#_c_834_n N_A_300_125#_c_898_n 0.00436498f $X=2.84 $Y=0.37
+ $X2=0 $Y2=0
cc_497 N_A_27_125#_c_834_n N_A_300_125#_c_948_n 0.0134462f $X=2.84 $Y=0.37 $X2=0
+ $Y2=0
cc_498 N_A_27_125#_M1011_d N_A_300_125#_c_899_n 0.00288015f $X=2.865 $Y=0.625
+ $X2=0 $Y2=0
cc_499 N_A_27_125#_c_834_n N_A_300_125#_c_899_n 0.00253018f $X=2.84 $Y=0.37
+ $X2=0 $Y2=0
cc_500 N_A_27_125#_c_835_n N_A_300_125#_c_899_n 0.0162401f $X=3.005 $Y=0.77
+ $X2=0 $Y2=0
cc_501 N_A_27_125#_c_834_n N_A_300_125#_c_902_n 0.00145328f $X=2.84 $Y=0.37
+ $X2=0 $Y2=0
cc_502 N_A_27_125#_c_834_n N_VGND_c_965_n 0.0111551f $X=2.84 $Y=0.37 $X2=0 $Y2=0
cc_503 N_A_27_125#_c_835_n N_VGND_c_965_n 0.0247045f $X=3.005 $Y=0.77 $X2=0
+ $Y2=0
cc_504 N_A_27_125#_c_829_n N_VGND_c_975_n 0.0369325f $X=0.975 $Y=0.35 $X2=0
+ $Y2=0
cc_505 N_A_27_125#_c_830_n N_VGND_c_975_n 0.0168561f $X=0.365 $Y=0.35 $X2=0
+ $Y2=0
cc_506 N_A_27_125#_c_832_n N_VGND_c_975_n 0.0401321f $X=1.975 $Y=0.35 $X2=0
+ $Y2=0
cc_507 N_A_27_125#_c_834_n N_VGND_c_975_n 0.0485706f $X=2.84 $Y=0.37 $X2=0 $Y2=0
cc_508 N_A_27_125#_c_836_n N_VGND_c_975_n 0.0222253f $X=1.14 $Y=0.35 $X2=0 $Y2=0
cc_509 N_A_27_125#_c_837_n N_VGND_c_975_n 0.022006f $X=2.14 $Y=0.36 $X2=0 $Y2=0
cc_510 N_A_27_125#_c_829_n N_VGND_c_980_n 0.0227893f $X=0.975 $Y=0.35 $X2=0
+ $Y2=0
cc_511 N_A_27_125#_c_830_n N_VGND_c_980_n 0.00967329f $X=0.365 $Y=0.35 $X2=0
+ $Y2=0
cc_512 N_A_27_125#_c_832_n N_VGND_c_980_n 0.022421f $X=1.975 $Y=0.35 $X2=0 $Y2=0
cc_513 N_A_27_125#_c_834_n N_VGND_c_980_n 0.0288613f $X=2.84 $Y=0.37 $X2=0 $Y2=0
cc_514 N_A_27_125#_c_836_n N_VGND_c_980_n 0.0127636f $X=1.14 $Y=0.35 $X2=0 $Y2=0
cc_515 N_A_27_125#_c_837_n N_VGND_c_980_n 0.0114038f $X=2.14 $Y=0.36 $X2=0 $Y2=0
cc_516 N_A_300_125#_c_899_n N_VGND_M1006_d 0.00242368f $X=3.94 $Y=1.19 $X2=-0.19
+ $Y2=-0.245
cc_517 N_A_300_125#_c_920_n N_VGND_M1009_d 0.00365842f $X=4.805 $Y=1.095 $X2=0
+ $Y2=0
cc_518 N_A_300_125#_c_899_n N_VGND_c_965_n 0.0219406f $X=3.94 $Y=1.19 $X2=0
+ $Y2=0
cc_519 N_A_300_125#_c_900_n N_VGND_c_965_n 0.0128711f $X=4.025 $Y=0.75 $X2=0
+ $Y2=0
cc_520 N_A_300_125#_c_900_n N_VGND_c_966_n 0.00946619f $X=4.025 $Y=0.75 $X2=0
+ $Y2=0
cc_521 N_A_300_125#_c_920_n N_VGND_c_966_n 0.0170777f $X=4.805 $Y=1.095 $X2=0
+ $Y2=0
cc_522 N_A_300_125#_c_901_n N_VGND_c_966_n 0.00911358f $X=4.89 $Y=0.755 $X2=0
+ $Y2=0
cc_523 N_A_300_125#_c_901_n N_VGND_c_967_n 0.0145518f $X=4.89 $Y=0.755 $X2=0
+ $Y2=0
cc_524 N_A_300_125#_c_900_n N_VGND_c_971_n 0.00389986f $X=4.025 $Y=0.75 $X2=0
+ $Y2=0
cc_525 N_A_300_125#_c_901_n N_VGND_c_973_n 0.0054105f $X=4.89 $Y=0.755 $X2=0
+ $Y2=0
cc_526 N_A_300_125#_c_900_n N_VGND_c_980_n 0.00476452f $X=4.025 $Y=0.75 $X2=0
+ $Y2=0
cc_527 N_A_300_125#_c_901_n N_VGND_c_980_n 0.00669947f $X=4.89 $Y=0.755 $X2=0
+ $Y2=0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or4b_4 A B C D_N VGND VNB VPB VPWR X
M1000 VGND a_27_74# X VNB nlowvt w=740000u l=150000u
+  ad=1.3615e+12p pd=1.11e+07u as=5.069e+11p ps=4.33e+06u
M1001 a_119_392# B a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=8.8e+11p ps=7.76e+06u
M1002 VPWR A a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=1.269e+12p pd=1.106e+07u as=0p ps=0u
M1003 a_499_392# C a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=0p ps=0u
M1004 a_27_74# a_563_48# a_499_392# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1005 a_27_392# B a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_119_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_499_392# a_563_48# a_27_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_392# C a_499_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND D_N a_563_48# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=3.2135e+11p ps=2.98e+06u
M1012 VGND a_27_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND C a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.2395e+12p ps=7.79e+06u
M1014 X a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1015 VPWR a_27_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_74# a_563_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND B a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR D_N a_563_48# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1020 VPWR a_27_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_27_74# A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

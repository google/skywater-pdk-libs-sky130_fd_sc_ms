* File: sky130_fd_sc_ms__o21a_2.pxi.spice
* Created: Wed Sep  2 12:21:37 2020
* 
x_PM_SKY130_FD_SC_MS__O21A_2%A1 N_A1_c_63_n N_A1_M1006_g N_A1_M1008_g
+ N_A1_c_65_n N_A1_c_66_n A1 A1 PM_SKY130_FD_SC_MS__O21A_2%A1
x_PM_SKY130_FD_SC_MS__O21A_2%A2 N_A2_M1001_g N_A2_M1005_g A2 N_A2_c_90_n
+ N_A2_c_91_n PM_SKY130_FD_SC_MS__O21A_2%A2
x_PM_SKY130_FD_SC_MS__O21A_2%B1 N_B1_M1000_g N_B1_M1009_g B1 N_B1_c_120_n
+ N_B1_c_121_n N_B1_c_122_n PM_SKY130_FD_SC_MS__O21A_2%B1
x_PM_SKY130_FD_SC_MS__O21A_2%A_247_368# N_A_247_368#_M1009_d
+ N_A_247_368#_M1001_d N_A_247_368#_M1002_g N_A_247_368#_M1004_g
+ N_A_247_368#_c_160_n N_A_247_368#_M1003_g N_A_247_368#_c_161_n
+ N_A_247_368#_c_162_n N_A_247_368#_c_163_n N_A_247_368#_M1007_g
+ N_A_247_368#_c_171_n N_A_247_368#_c_172_n N_A_247_368#_c_173_n
+ N_A_247_368#_c_164_n N_A_247_368#_c_165_n N_A_247_368#_c_166_n
+ N_A_247_368#_c_167_n N_A_247_368#_c_168_n
+ PM_SKY130_FD_SC_MS__O21A_2%A_247_368#
x_PM_SKY130_FD_SC_MS__O21A_2%VPWR N_VPWR_M1008_s N_VPWR_M1000_d N_VPWR_M1004_s
+ N_VPWR_c_237_n N_VPWR_c_238_n N_VPWR_c_239_n N_VPWR_c_240_n N_VPWR_c_241_n
+ VPWR N_VPWR_c_242_n N_VPWR_c_243_n N_VPWR_c_244_n N_VPWR_c_236_n
+ N_VPWR_c_246_n N_VPWR_c_247_n PM_SKY130_FD_SC_MS__O21A_2%VPWR
x_PM_SKY130_FD_SC_MS__O21A_2%X N_X_M1003_d N_X_M1002_d N_X_c_279_n X X X X
+ N_X_c_281_n X PM_SKY130_FD_SC_MS__O21A_2%X
x_PM_SKY130_FD_SC_MS__O21A_2%A_54_74# N_A_54_74#_M1006_s N_A_54_74#_M1005_d
+ N_A_54_74#_c_309_n N_A_54_74#_c_310_n N_A_54_74#_c_315_n N_A_54_74#_c_321_n
+ N_A_54_74#_c_311_n PM_SKY130_FD_SC_MS__O21A_2%A_54_74#
x_PM_SKY130_FD_SC_MS__O21A_2%VGND N_VGND_M1006_d N_VGND_M1003_s N_VGND_M1007_s
+ N_VGND_c_335_n N_VGND_c_336_n N_VGND_c_337_n N_VGND_c_338_n VGND
+ N_VGND_c_339_n N_VGND_c_340_n N_VGND_c_341_n N_VGND_c_342_n N_VGND_c_343_n
+ N_VGND_c_344_n PM_SKY130_FD_SC_MS__O21A_2%VGND
cc_1 VNB N_A1_c_63_n 0.0234618f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.22
cc_2 VNB N_A1_M1008_g 0.00923934f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.34
cc_3 VNB N_A1_c_65_n 0.0616222f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.385
cc_4 VNB N_A1_c_66_n 0.0114302f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.22
cc_5 VNB A1 0.0278098f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_6 VNB N_A2_M1001_g 0.00654075f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.74
cc_7 VNB A2 0.00587703f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.385
cc_8 VNB N_A2_c_90_n 0.0328928f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_9 VNB N_A2_c_91_n 0.0194558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B1_M1000_g 0.00748692f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.74
cc_11 VNB N_B1_c_120_n 0.0295946f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_12 VNB N_B1_c_121_n 0.00895346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B1_c_122_n 0.0199025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_247_368#_M1002_g 0.00674104f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.22
cc_15 VNB N_A_247_368#_M1004_g 0.00282595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_247_368#_c_160_n 0.0184836f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_17 VNB N_A_247_368#_c_161_n 0.0335612f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_18 VNB N_A_247_368#_c_162_n 0.0591743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_247_368#_c_163_n 0.0199304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_247_368#_c_164_n 0.00868066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_247_368#_c_165_n 0.0039379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_247_368#_c_166_n 0.00271468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_247_368#_c_167_n 0.00201793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_247_368#_c_168_n 0.00452572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_236_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB X 0.0162439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_54_74#_c_309_n 0.0071683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_54_74#_c_310_n 0.0222165f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.22
cc_29 VNB N_A_54_74#_c_311_n 0.00286839f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_30 VNB N_VGND_c_335_n 0.00811421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_336_n 0.0160569f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_32 VNB N_VGND_c_337_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_33 VNB N_VGND_c_338_n 0.0505973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_339_n 0.0232388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_340_n 0.0333734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_341_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_342_n 0.00911377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_343_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_344_n 0.238533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VPB N_A1_M1008_g 0.0283435f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=2.34
cc_41 VPB N_A2_M1001_g 0.0235529f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=0.74
cc_42 VPB N_B1_M1000_g 0.0246488f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=0.74
cc_43 VPB N_A_247_368#_M1002_g 0.02421f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.22
cc_44 VPB N_A_247_368#_M1004_g 0.0241923f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A_247_368#_c_171_n 0.00340823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_247_368#_c_172_n 0.0086276f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_247_368#_c_173_n 0.0100705f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_247_368#_c_166_n 0.00119878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_237_n 0.0610756f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_238_n 0.0123089f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.365
cc_51 VPB N_VPWR_c_239_n 0.0469031f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_240_n 0.0128037f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_241_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_242_n 0.0392809f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_243_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_244_n 0.0194863f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_236_n 0.107567f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_246_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_247_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_X_c_279_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.22
cc_61 VPB X 0.00412425f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_X_c_281_n 0.0116776f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.365
cc_63 N_A1_M1008_g N_A2_M1001_g 0.041709f $X=0.725 $Y=2.34 $X2=0 $Y2=0
cc_64 N_A1_c_66_n A2 3.8796e-19 $X=0.625 $Y=1.22 $X2=0 $Y2=0
cc_65 A1 A2 0.0257541f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_66 N_A1_c_66_n N_A2_c_90_n 0.0495672f $X=0.625 $Y=1.22 $X2=0 $Y2=0
cc_67 A1 N_A2_c_90_n 0.00227871f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_68 N_A1_c_63_n N_A2_c_91_n 0.0226983f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_69 N_A1_M1008_g N_VPWR_c_237_n 0.0273006f $X=0.725 $Y=2.34 $X2=0 $Y2=0
cc_70 N_A1_c_65_n N_VPWR_c_237_n 0.00660418f $X=0.625 $Y=1.385 $X2=0 $Y2=0
cc_71 A1 N_VPWR_c_237_n 0.0195859f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_72 N_A1_M1008_g N_VPWR_c_242_n 0.00492916f $X=0.725 $Y=2.34 $X2=0 $Y2=0
cc_73 N_A1_M1008_g N_VPWR_c_236_n 0.00511769f $X=0.725 $Y=2.34 $X2=0 $Y2=0
cc_74 N_A1_c_65_n N_A_54_74#_c_309_n 0.00229997f $X=0.625 $Y=1.385 $X2=0 $Y2=0
cc_75 A1 N_A_54_74#_c_309_n 0.0283136f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_76 N_A1_c_63_n N_A_54_74#_c_310_n 0.00977947f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_77 N_A1_c_63_n N_A_54_74#_c_315_n 0.0140987f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_78 A1 N_A_54_74#_c_315_n 0.0153682f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_79 N_A1_c_63_n N_VGND_c_335_n 0.0138709f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_80 N_A1_c_63_n N_VGND_c_339_n 0.00383152f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_81 N_A1_c_63_n N_VGND_c_344_n 0.00388149f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_82 N_A2_M1001_g N_B1_M1000_g 0.0254135f $X=1.145 $Y=2.34 $X2=0 $Y2=0
cc_83 A2 N_B1_c_120_n 3.71725e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_84 N_A2_c_90_n N_B1_c_120_n 0.0174273f $X=1.22 $Y=1.385 $X2=0 $Y2=0
cc_85 A2 N_B1_c_121_n 0.0283697f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_86 N_A2_c_91_n N_B1_c_121_n 0.00227475f $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_87 N_A2_c_91_n N_B1_c_122_n 0.0103208f $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_88 N_A2_M1001_g N_A_247_368#_c_171_n 0.0144897f $X=1.145 $Y=2.34 $X2=0 $Y2=0
cc_89 N_A2_M1001_g N_A_247_368#_c_173_n 0.00436267f $X=1.145 $Y=2.34 $X2=0 $Y2=0
cc_90 A2 N_A_247_368#_c_173_n 0.00503923f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_91 N_A2_c_90_n N_A_247_368#_c_173_n 4.61395e-19 $X=1.22 $Y=1.385 $X2=0 $Y2=0
cc_92 N_A2_M1001_g N_VPWR_c_237_n 0.00363017f $X=1.145 $Y=2.34 $X2=0 $Y2=0
cc_93 N_A2_M1001_g N_VPWR_c_242_n 0.0059286f $X=1.145 $Y=2.34 $X2=0 $Y2=0
cc_94 N_A2_M1001_g N_VPWR_c_236_n 0.00610055f $X=1.145 $Y=2.34 $X2=0 $Y2=0
cc_95 A2 N_A_54_74#_c_315_n 0.0228656f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_96 N_A2_c_90_n N_A_54_74#_c_315_n 9.98643e-19 $X=1.22 $Y=1.385 $X2=0 $Y2=0
cc_97 N_A2_c_91_n N_A_54_74#_c_315_n 0.0106434f $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_98 N_A2_c_91_n N_A_54_74#_c_311_n 4.10343e-19 $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_99 N_A2_c_91_n N_VGND_c_335_n 0.00532072f $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_100 N_A2_c_91_n N_VGND_c_340_n 0.00460063f $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_101 N_A2_c_91_n N_VGND_c_344_n 0.00464404f $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_102 N_B1_M1000_g N_A_247_368#_M1002_g 0.0146212f $X=1.715 $Y=2.34 $X2=0 $Y2=0
cc_103 N_B1_c_120_n N_A_247_368#_c_162_n 0.0107914f $X=1.79 $Y=1.385 $X2=0 $Y2=0
cc_104 N_B1_c_121_n N_A_247_368#_c_162_n 3.0788e-19 $X=1.79 $Y=1.385 $X2=0 $Y2=0
cc_105 N_B1_M1000_g N_A_247_368#_c_171_n 0.0163699f $X=1.715 $Y=2.34 $X2=0 $Y2=0
cc_106 N_B1_M1000_g N_A_247_368#_c_172_n 0.013848f $X=1.715 $Y=2.34 $X2=0 $Y2=0
cc_107 N_B1_c_120_n N_A_247_368#_c_172_n 0.00357978f $X=1.79 $Y=1.385 $X2=0
+ $Y2=0
cc_108 N_B1_c_121_n N_A_247_368#_c_172_n 0.0221503f $X=1.79 $Y=1.385 $X2=0 $Y2=0
cc_109 N_B1_M1000_g N_A_247_368#_c_173_n 0.00242377f $X=1.715 $Y=2.34 $X2=0
+ $Y2=0
cc_110 N_B1_c_121_n N_A_247_368#_c_173_n 0.00776619f $X=1.79 $Y=1.385 $X2=0
+ $Y2=0
cc_111 N_B1_c_122_n N_A_247_368#_c_164_n 6.80643e-19 $X=1.79 $Y=1.22 $X2=0 $Y2=0
cc_112 N_B1_c_121_n N_A_247_368#_c_165_n 0.00314775f $X=1.79 $Y=1.385 $X2=0
+ $Y2=0
cc_113 N_B1_c_122_n N_A_247_368#_c_165_n 0.00502808f $X=1.79 $Y=1.22 $X2=0 $Y2=0
cc_114 N_B1_M1000_g N_A_247_368#_c_166_n 0.00324601f $X=1.715 $Y=2.34 $X2=0
+ $Y2=0
cc_115 N_B1_c_120_n N_A_247_368#_c_167_n 3.15972e-19 $X=1.79 $Y=1.385 $X2=0
+ $Y2=0
cc_116 N_B1_c_121_n N_A_247_368#_c_167_n 0.00378611f $X=1.79 $Y=1.385 $X2=0
+ $Y2=0
cc_117 N_B1_c_120_n N_A_247_368#_c_168_n 0.00131824f $X=1.79 $Y=1.385 $X2=0
+ $Y2=0
cc_118 N_B1_c_121_n N_A_247_368#_c_168_n 0.0275093f $X=1.79 $Y=1.385 $X2=0 $Y2=0
cc_119 N_B1_M1000_g N_VPWR_c_238_n 0.0112281f $X=1.715 $Y=2.34 $X2=0 $Y2=0
cc_120 N_B1_M1000_g N_VPWR_c_242_n 0.00567889f $X=1.715 $Y=2.34 $X2=0 $Y2=0
cc_121 N_B1_M1000_g N_VPWR_c_236_n 0.00610055f $X=1.715 $Y=2.34 $X2=0 $Y2=0
cc_122 N_B1_M1000_g N_X_c_279_n 8.67015e-19 $X=1.715 $Y=2.34 $X2=0 $Y2=0
cc_123 N_B1_c_120_n N_A_54_74#_c_321_n 4.36016e-19 $X=1.79 $Y=1.385 $X2=0 $Y2=0
cc_124 N_B1_c_121_n N_A_54_74#_c_321_n 0.012077f $X=1.79 $Y=1.385 $X2=0 $Y2=0
cc_125 N_B1_c_122_n N_A_54_74#_c_321_n 0.00215143f $X=1.79 $Y=1.22 $X2=0 $Y2=0
cc_126 N_B1_c_122_n N_A_54_74#_c_311_n 0.00622341f $X=1.79 $Y=1.22 $X2=0 $Y2=0
cc_127 N_B1_c_122_n N_VGND_c_336_n 0.00313679f $X=1.79 $Y=1.22 $X2=0 $Y2=0
cc_128 N_B1_c_122_n N_VGND_c_340_n 0.00434054f $X=1.79 $Y=1.22 $X2=0 $Y2=0
cc_129 N_B1_c_122_n N_VGND_c_344_n 0.0082661f $X=1.79 $Y=1.22 $X2=0 $Y2=0
cc_130 N_A_247_368#_c_172_n N_VPWR_M1000_d 0.007823f $X=2.125 $Y=1.805 $X2=0
+ $Y2=0
cc_131 N_A_247_368#_c_171_n N_VPWR_c_237_n 0.0255922f $X=1.49 $Y=1.985 $X2=0
+ $Y2=0
cc_132 N_A_247_368#_c_173_n N_VPWR_c_237_n 0.00199752f $X=1.655 $Y=1.805 $X2=0
+ $Y2=0
cc_133 N_A_247_368#_M1002_g N_VPWR_c_238_n 0.00381877f $X=2.405 $Y=2.4 $X2=0
+ $Y2=0
cc_134 N_A_247_368#_c_171_n N_VPWR_c_238_n 0.0391818f $X=1.49 $Y=1.985 $X2=0
+ $Y2=0
cc_135 N_A_247_368#_c_172_n N_VPWR_c_238_n 0.0243097f $X=2.125 $Y=1.805 $X2=0
+ $Y2=0
cc_136 N_A_247_368#_M1004_g N_VPWR_c_239_n 0.00809945f $X=2.855 $Y=2.4 $X2=0
+ $Y2=0
cc_137 N_A_247_368#_c_171_n N_VPWR_c_242_n 0.00975961f $X=1.49 $Y=1.985 $X2=0
+ $Y2=0
cc_138 N_A_247_368#_M1002_g N_VPWR_c_243_n 0.005209f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A_247_368#_M1004_g N_VPWR_c_243_n 0.005209f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A_247_368#_M1002_g N_VPWR_c_236_n 0.00986727f $X=2.405 $Y=2.4 $X2=0
+ $Y2=0
cc_141 N_A_247_368#_M1004_g N_VPWR_c_236_n 0.00986727f $X=2.855 $Y=2.4 $X2=0
+ $Y2=0
cc_142 N_A_247_368#_c_171_n N_VPWR_c_236_n 0.0111753f $X=1.49 $Y=1.985 $X2=0
+ $Y2=0
cc_143 N_A_247_368#_M1002_g N_X_c_279_n 0.0157148f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A_247_368#_M1004_g N_X_c_279_n 0.0195696f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_145 N_A_247_368#_M1004_g X 0.00347091f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_146 N_A_247_368#_c_160_n X 0.0137211f $X=2.915 $Y=1.22 $X2=0 $Y2=0
cc_147 N_A_247_368#_c_161_n X 0.0191488f $X=3.27 $Y=1.295 $X2=0 $Y2=0
cc_148 N_A_247_368#_c_162_n X 0.012068f $X=2.99 $Y=1.295 $X2=0 $Y2=0
cc_149 N_A_247_368#_c_163_n X 0.0148558f $X=3.345 $Y=1.22 $X2=0 $Y2=0
cc_150 N_A_247_368#_c_165_n X 0.00446539f $X=2.21 $Y=1.22 $X2=0 $Y2=0
cc_151 N_A_247_368#_c_166_n X 0.00504242f $X=2.21 $Y=1.72 $X2=0 $Y2=0
cc_152 N_A_247_368#_c_168_n X 0.0161585f $X=2.48 $Y=1.385 $X2=0 $Y2=0
cc_153 N_A_247_368#_M1002_g N_X_c_281_n 0.0037987f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_154 N_A_247_368#_M1004_g N_X_c_281_n 0.0217953f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_155 N_A_247_368#_c_162_n N_X_c_281_n 0.00403718f $X=2.99 $Y=1.295 $X2=0 $Y2=0
cc_156 N_A_247_368#_c_172_n N_X_c_281_n 0.0126349f $X=2.125 $Y=1.805 $X2=0 $Y2=0
cc_157 N_A_247_368#_c_168_n N_X_c_281_n 0.0134173f $X=2.48 $Y=1.385 $X2=0 $Y2=0
cc_158 N_A_247_368#_c_164_n N_A_54_74#_c_311_n 0.0199611f $X=2 $Y=0.505 $X2=0
+ $Y2=0
cc_159 N_A_247_368#_c_160_n N_VGND_c_336_n 0.0182605f $X=2.915 $Y=1.22 $X2=0
+ $Y2=0
cc_160 N_A_247_368#_c_162_n N_VGND_c_336_n 0.0094957f $X=2.99 $Y=1.295 $X2=0
+ $Y2=0
cc_161 N_A_247_368#_c_164_n N_VGND_c_336_n 0.0595951f $X=2 $Y=0.505 $X2=0 $Y2=0
cc_162 N_A_247_368#_c_168_n N_VGND_c_336_n 0.0148152f $X=2.48 $Y=1.385 $X2=0
+ $Y2=0
cc_163 N_A_247_368#_c_163_n N_VGND_c_338_n 0.00647412f $X=3.345 $Y=1.22 $X2=0
+ $Y2=0
cc_164 N_A_247_368#_c_164_n N_VGND_c_340_n 0.0180247f $X=2 $Y=0.505 $X2=0 $Y2=0
cc_165 N_A_247_368#_c_160_n N_VGND_c_341_n 0.00434272f $X=2.915 $Y=1.22 $X2=0
+ $Y2=0
cc_166 N_A_247_368#_c_163_n N_VGND_c_341_n 0.00434272f $X=3.345 $Y=1.22 $X2=0
+ $Y2=0
cc_167 N_A_247_368#_c_160_n N_VGND_c_344_n 0.00825059f $X=2.915 $Y=1.22 $X2=0
+ $Y2=0
cc_168 N_A_247_368#_c_163_n N_VGND_c_344_n 0.00823942f $X=3.345 $Y=1.22 $X2=0
+ $Y2=0
cc_169 N_A_247_368#_c_164_n N_VGND_c_344_n 0.0144116f $X=2 $Y=0.505 $X2=0 $Y2=0
cc_170 N_VPWR_c_238_n N_X_c_279_n 0.0353111f $X=2.13 $Y=2.145 $X2=0 $Y2=0
cc_171 N_VPWR_c_239_n N_X_c_279_n 0.0353111f $X=3.13 $Y=2.225 $X2=0 $Y2=0
cc_172 N_VPWR_c_243_n N_X_c_279_n 0.0144623f $X=2.965 $Y=3.33 $X2=0 $Y2=0
cc_173 N_VPWR_c_236_n N_X_c_279_n 0.0118344f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_174 N_VPWR_M1004_s N_X_c_281_n 0.00330887f $X=2.945 $Y=1.84 $X2=0 $Y2=0
cc_175 N_VPWR_c_239_n N_X_c_281_n 0.0238156f $X=3.13 $Y=2.225 $X2=0 $Y2=0
cc_176 X N_VGND_c_336_n 0.0270562f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_177 N_X_c_281_n N_VGND_c_336_n 0.00421771f $X=3.13 $Y=1.72 $X2=0 $Y2=0
cc_178 X N_VGND_c_338_n 0.0294122f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_179 X N_VGND_c_341_n 0.0144922f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_180 X N_VGND_c_344_n 0.0118826f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_181 N_A_54_74#_c_315_n N_VGND_M1006_d 0.0146092f $X=1.405 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_182 N_A_54_74#_c_310_n N_VGND_c_335_n 0.0115542f $X=0.415 $Y=0.505 $X2=0
+ $Y2=0
cc_183 N_A_54_74#_c_315_n N_VGND_c_335_n 0.0219781f $X=1.405 $Y=0.925 $X2=0
+ $Y2=0
cc_184 N_A_54_74#_c_311_n N_VGND_c_335_n 0.00248533f $X=1.57 $Y=0.505 $X2=0
+ $Y2=0
cc_185 N_A_54_74#_c_310_n N_VGND_c_339_n 0.0152302f $X=0.415 $Y=0.505 $X2=0
+ $Y2=0
cc_186 N_A_54_74#_c_311_n N_VGND_c_340_n 0.0151574f $X=1.57 $Y=0.505 $X2=0 $Y2=0
cc_187 N_A_54_74#_c_310_n N_VGND_c_344_n 0.0121804f $X=0.415 $Y=0.505 $X2=0
+ $Y2=0
cc_188 N_A_54_74#_c_315_n N_VGND_c_344_n 0.0115606f $X=1.405 $Y=0.925 $X2=0
+ $Y2=0
cc_189 N_A_54_74#_c_311_n N_VGND_c_344_n 0.0120652f $X=1.57 $Y=0.505 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__nor2_8.spice
* Created: Wed Sep  2 12:15:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nor2_8.pex.spice"
.subckt sky130_fd_sc_ms__nor2_8  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_M1002_g N_Y_M1002_s VNB NLOWVT L=0.15 W=0.74 AD=0.7881
+ AS=0.1295 PD=3.61 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75001 SB=75004.8
+ A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_A_M1005_g N_Y_M1002_s VNB NLOWVT L=0.15 W=0.74 AD=0.2775
+ AS=0.1295 PD=1.49 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.5 SB=75004.3
+ A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1005_d N_A_M1014_g N_Y_M1014_s VNB NLOWVT L=0.15 W=0.74 AD=0.2775
+ AS=0.1295 PD=1.49 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.4 SB=75003.4
+ A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1016_d N_A_M1016_g N_Y_M1014_s VNB NLOWVT L=0.15 W=0.74 AD=0.1295
+ AS=0.1295 PD=1.09 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.9 SB=75002.9
+ A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1016_d N_B_M1000_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74 AD=0.1295
+ AS=0.35705 PD=1.09 PS=1.705 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75003.4
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_B_M1008_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.35705 PD=1.16 PS=1.705 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75004.5
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1008_d N_B_M1009_g N_Y_M1009_s VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75005.1 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1023 N_VGND_M1023_d N_B_M1023_g N_Y_M1009_s VNB NLOWVT L=0.15 W=0.74 AD=0.2627
+ AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75005.5 SB=75000.3
+ A=0.111 P=1.78 MULT=1
MM1001 N_A_27_368#_M1001_d N_A_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1792 PD=2.8 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.2
+ SB=90007.3 A=0.2016 P=2.6 MULT=1
MM1003 N_A_27_368#_M1003_d N_A_M1003_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.7
+ SB=90006.8 A=0.2016 P=2.6 MULT=1
MM1004 N_A_27_368#_M1003_d N_A_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90006.4 A=0.2016 P=2.6 MULT=1
MM1006 N_A_27_368#_M1006_d N_A_M1006_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.6
+ SB=90005.9 A=0.2016 P=2.6 MULT=1
MM1007 N_A_27_368#_M1006_d N_A_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002
+ SB=90005.5 A=0.2016 P=2.6 MULT=1
MM1010 N_A_27_368#_M1010_d N_A_M1010_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.5
+ SB=90005 A=0.2016 P=2.6 MULT=1
MM1011 N_A_27_368#_M1010_d N_A_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003
+ SB=90004.5 A=0.2016 P=2.6 MULT=1
MM1015 N_A_27_368#_M1015_d N_A_M1015_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003.5
+ SB=90004 A=0.2016 P=2.6 MULT=1
MM1012 N_Y_M1012_d N_B_M1012_g N_A_27_368#_M1015_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90004
+ SB=90003.5 A=0.2016 P=2.6 MULT=1
MM1013 N_Y_M1012_d N_B_M1013_g N_A_27_368#_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90004.5
+ SB=90003 A=0.2016 P=2.6 MULT=1
MM1017 N_Y_M1017_d N_B_M1017_g N_A_27_368#_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90005
+ SB=90002.5 A=0.2016 P=2.6 MULT=1
MM1018 N_Y_M1017_d N_B_M1018_g N_A_27_368#_M1018_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90005.4
+ SB=90002.1 A=0.2016 P=2.6 MULT=1
MM1019 N_Y_M1019_d N_B_M1019_g N_A_27_368#_M1018_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90005.9
+ SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1020 N_Y_M1019_d N_B_M1020_g N_A_27_368#_M1020_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90006.3
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1021 N_Y_M1021_d N_B_M1021_g N_A_27_368#_M1020_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90006.8
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1022 N_Y_M1021_d N_B_M1022_g N_A_27_368#_M1022_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90007.3
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX24_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_ms__nor2_8.pxi.spice"
*
.ends
*
*

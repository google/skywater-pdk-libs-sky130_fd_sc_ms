* File: sky130_fd_sc_ms__dfsbp_2.pxi.spice
* Created: Fri Aug 28 17:23:40 2020
* 
x_PM_SKY130_FD_SC_MS__DFSBP_2%D N_D_c_278_n N_D_M1029_g N_D_M1033_g D D
+ N_D_c_280_n N_D_c_281_n N_D_c_285_n PM_SKY130_FD_SC_MS__DFSBP_2%D
x_PM_SKY130_FD_SC_MS__DFSBP_2%CLK N_CLK_M1035_g N_CLK_M1018_g CLK N_CLK_c_314_n
+ N_CLK_c_315_n PM_SKY130_FD_SC_MS__DFSBP_2%CLK
x_PM_SKY130_FD_SC_MS__DFSBP_2%A_398_74# N_A_398_74#_M1019_d N_A_398_74#_M1021_d
+ N_A_398_74#_c_351_n N_A_398_74#_c_370_n N_A_398_74#_M1001_g
+ N_A_398_74#_c_352_n N_A_398_74#_M1036_g N_A_398_74#_M1022_g
+ N_A_398_74#_M1010_g N_A_398_74#_c_374_n N_A_398_74#_c_354_n
+ N_A_398_74#_c_478_p N_A_398_74#_c_355_n N_A_398_74#_c_356_n
+ N_A_398_74#_c_375_n N_A_398_74#_c_376_n N_A_398_74#_c_357_n
+ N_A_398_74#_c_358_n N_A_398_74#_c_359_n N_A_398_74#_c_380_n
+ N_A_398_74#_c_393_p N_A_398_74#_c_381_n N_A_398_74#_c_382_n
+ N_A_398_74#_c_383_n N_A_398_74#_c_384_n N_A_398_74#_c_385_n
+ N_A_398_74#_c_386_n N_A_398_74#_c_360_n N_A_398_74#_c_361_n
+ N_A_398_74#_c_362_n N_A_398_74#_c_363_n N_A_398_74#_c_364_n
+ N_A_398_74#_c_395_p N_A_398_74#_c_365_n N_A_398_74#_c_366_n
+ N_A_398_74#_c_388_n N_A_398_74#_c_367_n N_A_398_74#_c_368_n
+ N_A_398_74#_c_390_n PM_SKY130_FD_SC_MS__DFSBP_2%A_398_74#
x_PM_SKY130_FD_SC_MS__DFSBP_2%A_757_401# N_A_757_401#_M1032_s
+ N_A_757_401#_M1020_d N_A_757_401#_M1009_g N_A_757_401#_c_621_n
+ N_A_757_401#_M1025_g N_A_757_401#_c_627_n N_A_757_401#_c_628_n
+ N_A_757_401#_c_622_n N_A_757_401#_c_623_n N_A_757_401#_c_629_n
+ N_A_757_401#_c_630_n N_A_757_401#_c_631_n N_A_757_401#_c_624_n
+ N_A_757_401#_c_632_n N_A_757_401#_c_625_n
+ PM_SKY130_FD_SC_MS__DFSBP_2%A_757_401#
x_PM_SKY130_FD_SC_MS__DFSBP_2%A_595_97# N_A_595_97#_M1017_d N_A_595_97#_M1001_d
+ N_A_595_97#_M1020_g N_A_595_97#_M1032_g N_A_595_97#_c_710_n
+ N_A_595_97#_M1006_g N_A_595_97#_c_712_n N_A_595_97#_M1012_g
+ N_A_595_97#_c_713_n N_A_595_97#_c_714_n N_A_595_97#_c_715_n
+ N_A_595_97#_c_716_n N_A_595_97#_c_717_n N_A_595_97#_c_718_n
+ N_A_595_97#_c_719_n N_A_595_97#_c_720_n N_A_595_97#_c_732_n
+ N_A_595_97#_c_773_n N_A_595_97#_c_721_n N_A_595_97#_c_722_n
+ N_A_595_97#_c_723_n N_A_595_97#_c_724_n N_A_595_97#_c_725_n
+ N_A_595_97#_c_726_n PM_SKY130_FD_SC_MS__DFSBP_2%A_595_97#
x_PM_SKY130_FD_SC_MS__DFSBP_2%SET_B N_SET_B_M1028_g N_SET_B_M1000_g
+ N_SET_B_c_872_n N_SET_B_M1002_g N_SET_B_c_873_n N_SET_B_c_874_n
+ N_SET_B_M1034_g N_SET_B_c_876_n N_SET_B_c_877_n N_SET_B_c_878_n
+ N_SET_B_c_879_n N_SET_B_c_880_n SET_B N_SET_B_c_891_n N_SET_B_c_882_n
+ N_SET_B_c_883_n N_SET_B_c_884_n PM_SKY130_FD_SC_MS__DFSBP_2%SET_B
x_PM_SKY130_FD_SC_MS__DFSBP_2%A_225_74# N_A_225_74#_M1035_s N_A_225_74#_M1018_s
+ N_A_225_74#_M1019_g N_A_225_74#_M1021_g N_A_225_74#_c_1006_n
+ N_A_225_74#_c_994_n N_A_225_74#_c_1007_n N_A_225_74#_c_1008_n
+ N_A_225_74#_M1017_g N_A_225_74#_M1005_g N_A_225_74#_c_1010_n
+ N_A_225_74#_M1027_g N_A_225_74#_c_996_n N_A_225_74#_c_997_n
+ N_A_225_74#_M1037_g N_A_225_74#_c_999_n N_A_225_74#_c_1000_n
+ N_A_225_74#_c_1001_n N_A_225_74#_c_1017_n N_A_225_74#_c_1002_n
+ N_A_225_74#_c_1019_n N_A_225_74#_c_1020_n N_A_225_74#_c_1021_n
+ N_A_225_74#_c_1003_n N_A_225_74#_c_1004_n N_A_225_74#_c_1023_n
+ PM_SKY130_FD_SC_MS__DFSBP_2%A_225_74#
x_PM_SKY130_FD_SC_MS__DFSBP_2%A_1501_92# N_A_1501_92#_M1003_d
+ N_A_1501_92#_M1026_s N_A_1501_92#_M1023_g N_A_1501_92#_M1031_g
+ N_A_1501_92#_c_1175_n N_A_1501_92#_c_1176_n N_A_1501_92#_c_1209_n
+ N_A_1501_92#_c_1193_n N_A_1501_92#_c_1183_n N_A_1501_92#_c_1177_n
+ N_A_1501_92#_c_1178_n N_A_1501_92#_c_1185_n N_A_1501_92#_c_1179_n
+ PM_SKY130_FD_SC_MS__DFSBP_2%A_1501_92#
x_PM_SKY130_FD_SC_MS__DFSBP_2%A_1339_74# N_A_1339_74#_M1022_d
+ N_A_1339_74#_M1027_d N_A_1339_74#_M1034_d N_A_1339_74#_M1003_g
+ N_A_1339_74#_c_1274_n N_A_1339_74#_c_1275_n N_A_1339_74#_M1026_g
+ N_A_1339_74#_c_1276_n N_A_1339_74#_M1008_g N_A_1339_74#_M1013_g
+ N_A_1339_74#_M1030_g N_A_1339_74#_M1024_g N_A_1339_74#_c_1281_n
+ N_A_1339_74#_c_1282_n N_A_1339_74#_M1015_g N_A_1339_74#_M1007_g
+ N_A_1339_74#_c_1285_n N_A_1339_74#_c_1305_n N_A_1339_74#_c_1295_n
+ N_A_1339_74#_c_1286_n N_A_1339_74#_c_1296_n N_A_1339_74#_c_1287_n
+ N_A_1339_74#_c_1298_n N_A_1339_74#_c_1299_n N_A_1339_74#_c_1300_n
+ N_A_1339_74#_c_1301_n N_A_1339_74#_c_1302_n N_A_1339_74#_c_1288_n
+ PM_SKY130_FD_SC_MS__DFSBP_2%A_1339_74#
x_PM_SKY130_FD_SC_MS__DFSBP_2%A_2221_74# N_A_2221_74#_M1007_s
+ N_A_2221_74#_M1015_s N_A_2221_74#_M1011_g N_A_2221_74#_M1004_g
+ N_A_2221_74#_M1014_g N_A_2221_74#_M1016_g N_A_2221_74#_c_1462_n
+ N_A_2221_74#_c_1463_n N_A_2221_74#_c_1464_n N_A_2221_74#_c_1465_n
+ N_A_2221_74#_c_1466_n PM_SKY130_FD_SC_MS__DFSBP_2%A_2221_74#
x_PM_SKY130_FD_SC_MS__DFSBP_2%A_27_74# N_A_27_74#_M1033_s N_A_27_74#_M1017_s
+ N_A_27_74#_M1029_s N_A_27_74#_M1001_s N_A_27_74#_c_1529_n N_A_27_74#_c_1530_n
+ N_A_27_74#_c_1535_n N_A_27_74#_c_1536_n N_A_27_74#_c_1537_n
+ N_A_27_74#_c_1531_n N_A_27_74#_c_1532_n N_A_27_74#_c_1539_n
+ N_A_27_74#_c_1581_n N_A_27_74#_c_1533_n PM_SKY130_FD_SC_MS__DFSBP_2%A_27_74#
x_PM_SKY130_FD_SC_MS__DFSBP_2%VPWR N_VPWR_M1029_d N_VPWR_M1018_d N_VPWR_M1009_d
+ N_VPWR_M1000_d N_VPWR_M1031_d N_VPWR_M1026_d N_VPWR_M1030_s N_VPWR_M1015_d
+ N_VPWR_M1014_s N_VPWR_c_1599_n N_VPWR_c_1600_n N_VPWR_c_1601_n N_VPWR_c_1602_n
+ N_VPWR_c_1603_n N_VPWR_c_1604_n N_VPWR_c_1605_n N_VPWR_c_1606_n
+ N_VPWR_c_1607_n N_VPWR_c_1608_n N_VPWR_c_1609_n N_VPWR_c_1610_n
+ N_VPWR_c_1611_n N_VPWR_c_1612_n VPWR N_VPWR_c_1613_n N_VPWR_c_1614_n
+ N_VPWR_c_1615_n N_VPWR_c_1616_n N_VPWR_c_1617_n N_VPWR_c_1618_n
+ N_VPWR_c_1619_n N_VPWR_c_1620_n N_VPWR_c_1621_n N_VPWR_c_1622_n
+ N_VPWR_c_1623_n N_VPWR_c_1624_n N_VPWR_c_1625_n N_VPWR_c_1598_n
+ PM_SKY130_FD_SC_MS__DFSBP_2%VPWR
x_PM_SKY130_FD_SC_MS__DFSBP_2%Q_N N_Q_N_M1013_d N_Q_N_M1008_d Q_N Q_N Q_N Q_N
+ Q_N Q_N PM_SKY130_FD_SC_MS__DFSBP_2%Q_N
x_PM_SKY130_FD_SC_MS__DFSBP_2%Q N_Q_M1004_s N_Q_M1011_d N_Q_c_1779_n
+ N_Q_c_1780_n N_Q_c_1776_n Q Q Q PM_SKY130_FD_SC_MS__DFSBP_2%Q
x_PM_SKY130_FD_SC_MS__DFSBP_2%VGND N_VGND_M1033_d N_VGND_M1035_d N_VGND_M1025_d
+ N_VGND_M1028_d N_VGND_M1002_d N_VGND_M1013_s N_VGND_M1024_s N_VGND_M1007_d
+ N_VGND_M1016_d N_VGND_c_1809_n N_VGND_c_1810_n N_VGND_c_1811_n N_VGND_c_1812_n
+ N_VGND_c_1813_n N_VGND_c_1814_n N_VGND_c_1815_n N_VGND_c_1816_n
+ N_VGND_c_1817_n N_VGND_c_1818_n N_VGND_c_1819_n VGND N_VGND_c_1820_n
+ N_VGND_c_1821_n N_VGND_c_1822_n N_VGND_c_1823_n N_VGND_c_1824_n
+ N_VGND_c_1825_n N_VGND_c_1826_n N_VGND_c_1827_n N_VGND_c_1828_n
+ N_VGND_c_1829_n N_VGND_c_1830_n N_VGND_c_1831_n N_VGND_c_1832_n
+ N_VGND_c_1833_n N_VGND_c_1834_n PM_SKY130_FD_SC_MS__DFSBP_2%VGND
cc_1 VNB N_D_c_278_n 0.0447809f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.795
cc_2 VNB N_D_M1033_g 0.0283644f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_3 VNB N_D_c_280_n 0.025337f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_4 VNB N_D_c_281_n 0.00250659f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_5 VNB N_CLK_M1018_g 0.00385449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB CLK 0.00845272f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_7 VNB N_CLK_c_314_n 0.0322132f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_8 VNB N_CLK_c_315_n 0.0199636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_398_74#_c_351_n 0.0152453f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.98
cc_10 VNB N_A_398_74#_c_352_n 0.0218688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_398_74#_M1036_g 0.0428034f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_12 VNB N_A_398_74#_c_354_n 0.00150841f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_13 VNB N_A_398_74#_c_355_n 0.0225218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_398_74#_c_356_n 0.00264685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_398_74#_c_357_n 0.00184302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_398_74#_c_358_n 0.0017748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_398_74#_c_359_n 0.0180595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_398_74#_c_360_n 0.00252917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_398_74#_c_361_n 0.00213435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_398_74#_c_362_n 0.0185305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_398_74#_c_363_n 0.00189911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_398_74#_c_364_n 0.00652496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_398_74#_c_365_n 0.00733674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_398_74#_c_366_n 0.0309266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_398_74#_c_367_n 0.00534817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_398_74#_c_368_n 0.0194713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_757_401#_c_621_n 0.0184264f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_28 VNB N_A_757_401#_c_622_n 0.0584491f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_29 VNB N_A_757_401#_c_623_n 0.00815564f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_30 VNB N_A_757_401#_c_624_n 0.018262f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_31 VNB N_A_757_401#_c_625_n 0.0154979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_595_97#_M1032_g 0.0511561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_595_97#_c_710_n 0.0160274f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_34 VNB N_A_595_97#_M1006_g 0.0157366f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.825
cc_35 VNB N_A_595_97#_c_712_n 0.021832f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_36 VNB N_A_595_97#_c_713_n 0.00651763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_595_97#_c_714_n 0.00248621f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.665
cc_38 VNB N_A_595_97#_c_715_n 0.0013452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_595_97#_c_716_n 0.00289252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_595_97#_c_717_n 0.0134003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_595_97#_c_718_n 0.00439152f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_595_97#_c_719_n 0.00427182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_595_97#_c_720_n 8.90541e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_595_97#_c_721_n 0.00213571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_595_97#_c_722_n 0.00547595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_595_97#_c_723_n 0.00856211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_595_97#_c_724_n 0.00247208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_595_97#_c_725_n 0.0185631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_595_97#_c_726_n 0.0380798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_SET_B_c_872_n 0.016029f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_SET_B_c_873_n 0.0185076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_SET_B_c_874_n 0.00564647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_SET_B_M1034_g 0.00734157f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_54 VNB N_SET_B_c_876_n 0.0186942f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.825
cc_55 VNB N_SET_B_c_877_n 0.012641f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_56 VNB N_SET_B_c_878_n 0.0137927f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_57 VNB N_SET_B_c_879_n 0.00275558f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.99
cc_58 VNB N_SET_B_c_880_n 0.00127012f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.295
cc_59 VNB SET_B 6.91838e-19 $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.665
cc_60 VNB N_SET_B_c_882_n 0.0341432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_SET_B_c_883_n 0.0405859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_SET_B_c_884_n 0.00406556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_225_74#_M1019_g 0.0224523f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_64 VNB N_A_225_74#_c_994_n 0.0289831f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_65 VNB N_A_225_74#_M1017_g 0.0210047f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_66 VNB N_A_225_74#_c_996_n 0.00841887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_225_74#_c_997_n 8.10579e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_225_74#_M1037_g 0.0446676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_225_74#_c_999_n 0.0123708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_225_74#_c_1000_n 0.0254751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_225_74#_c_1001_n 0.0195044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_225_74#_c_1002_n 0.0104758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_225_74#_c_1003_n 0.00365457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_225_74#_c_1004_n 0.0130637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1501_92#_M1023_g 0.0323321f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_76 VNB N_A_1501_92#_c_1175_n 0.00698987f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.145
cc_77 VNB N_A_1501_92#_c_1176_n 0.0327285f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.98
cc_78 VNB N_A_1501_92#_c_1177_n 0.0133421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1501_92#_c_1178_n 0.00405333f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.665
cc_80 VNB N_A_1501_92#_c_1179_n 0.0100146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1339_74#_M1003_g 0.0361264f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_82 VNB N_A_1339_74#_c_1274_n 0.0185463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1339_74#_c_1275_n 0.00960128f $X=-0.19 $Y=-0.245 $X2=0.61
+ $Y2=1.145
cc_84 VNB N_A_1339_74#_c_1276_n 0.0238846f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_85 VNB N_A_1339_74#_M1008_g 0.00161699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1339_74#_M1013_g 0.0259325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1339_74#_M1030_g 0.00177582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1339_74#_M1024_g 0.0258655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1339_74#_c_1281_n 0.0698362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1339_74#_c_1282_n 0.0241532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1339_74#_M1015_g 0.00201707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1339_74#_M1007_g 0.0364692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1339_74#_c_1285_n 0.00889457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1339_74#_c_1286_n 0.00581877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1339_74#_c_1287_n 0.00629293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1339_74#_c_1288_n 0.011619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_2221_74#_M1011_g 0.00167302f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_98 VNB N_A_2221_74#_M1004_g 0.0230317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_2221_74#_M1014_g 0.00231818f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_100 VNB N_A_2221_74#_M1016_g 0.0260184f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_101 VNB N_A_2221_74#_c_1462_n 0.0123246f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.295
cc_102 VNB N_A_2221_74#_c_1463_n 3.56488e-19 $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.825
cc_103 VNB N_A_2221_74#_c_1464_n 0.0072339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_2221_74#_c_1465_n 6.27903e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_2221_74#_c_1466_n 0.0645911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_27_74#_c_1529_n 0.0146704f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_107 VNB N_A_27_74#_c_1530_n 0.040185f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.98
cc_108 VNB N_A_27_74#_c_1531_n 0.00621313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_27_74#_c_1532_n 0.00791533f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_110 VNB N_A_27_74#_c_1533_n 0.00628546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VPWR_c_1598_n 0.541827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB Q_N 0.00397681f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.98
cc_113 VNB N_Q_c_1776_n 0.00141953f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.145
cc_114 VNB Q 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_115 VNB Q 0.00429087f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_116 VNB N_VGND_c_1809_n 0.0077412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1810_n 0.0221343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1811_n 0.00564229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1812_n 0.0119517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1813_n 0.0176142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1814_n 0.0194608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1815_n 0.0112908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1816_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1817_n 0.0505285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1818_n 0.0171743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1819_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1820_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1821_n 0.0558487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1822_n 0.0245702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1823_n 0.0206041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1824_n 0.0189349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1825_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1826_n 0.00481148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1827_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1828_n 0.0311101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1829_n 0.0239278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1830_n 0.0493081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1831_n 0.0419048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_1832_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_1833_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_1834_n 0.720699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VPB N_D_c_278_n 0.0126737f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.795
cc_143 VPB N_D_M1029_g 0.0635978f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.75
cc_144 VPB N_D_c_281_n 0.00207792f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_145 VPB N_D_c_285_n 0.0244074f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_146 VPB N_CLK_M1018_g 0.0238474f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_398_74#_c_351_n 0.00815295f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.98
cc_148 VPB N_A_398_74#_c_370_n 0.0132143f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_149 VPB N_A_398_74#_M1001_g 0.0239798f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_150 VPB N_A_398_74#_c_352_n 0.0167993f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_398_74#_M1010_g 0.0262284f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_398_74#_c_374_n 0.017404f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_398_74#_c_375_n 0.0225094f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_398_74#_c_376_n 0.00313547f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_398_74#_c_357_n 0.00298749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_398_74#_c_358_n 0.00604873f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_398_74#_c_359_n 0.021928f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_398_74#_c_380_n 0.00195993f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_398_74#_c_381_n 0.00400201f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_398_74#_c_382_n 0.0152159f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_398_74#_c_383_n 0.00260501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_398_74#_c_384_n 0.00197523f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_398_74#_c_385_n 0.00567462f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_398_74#_c_386_n 6.92221e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_398_74#_c_361_n 0.00428605f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_398_74#_c_388_n 0.00176185f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_398_74#_c_367_n 0.00576515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_398_74#_c_390_n 0.0408875f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_757_401#_M1009_g 0.0205265f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_170 VPB N_A_757_401#_c_627_n 0.012156f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_757_401#_c_628_n 0.0116824f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.145
cc_172 VPB N_A_757_401#_c_629_n 0.00575682f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_173 VPB N_A_757_401#_c_630_n 0.00369936f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_174 VPB N_A_757_401#_c_631_n 0.0358692f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_757_401#_c_632_n 0.0110022f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_757_401#_c_625_n 0.0114856f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_595_97#_M1020_g 0.0373067f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_178 VPB N_A_595_97#_M1006_g 0.0264745f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.825
cc_179 VPB N_A_595_97#_c_716_n 0.00764653f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_595_97#_c_719_n 0.00348451f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_595_97#_c_720_n 0.00251531f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_595_97#_c_732_n 0.00283654f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_595_97#_c_722_n 0.00116107f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_595_97#_c_723_n 0.0227484f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_SET_B_M1000_g 0.0314086f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_186 VPB N_SET_B_M1034_g 0.0712589f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_187 VPB N_SET_B_c_878_n 0.0194185f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_188 VPB N_SET_B_c_879_n 0.00103021f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.99
cc_189 VPB N_SET_B_c_880_n 0.00772355f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.295
cc_190 VPB SET_B 0.00113364f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_191 VPB N_SET_B_c_891_n 0.0343035f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_SET_B_c_882_n 0.00480279f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_SET_B_c_884_n 0.00291878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_225_74#_M1021_g 0.0197043f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_225_74#_c_1006_n 0.0734122f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_196 VPB N_A_225_74#_c_1007_n 0.0522732f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.825
cc_197 VPB N_A_225_74#_c_1008_n 0.0125859f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_198 VPB N_A_225_74#_M1005_g 0.0339302f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_199 VPB N_A_225_74#_c_1010_n 0.243267f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_200 VPB N_A_225_74#_M1027_g 0.0189716f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_225_74#_c_996_n 0.0321991f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_225_74#_c_997_n 0.00757347f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_225_74#_c_999_n 0.00170265f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_225_74#_c_1000_n 5.35904e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_225_74#_c_1001_n 0.00577555f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_225_74#_c_1017_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_225_74#_c_1002_n 0.00240536f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_225_74#_c_1019_n 0.0058961f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_225_74#_c_1020_n 0.00539283f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_225_74#_c_1021_n 0.00446037f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_225_74#_c_1003_n 5.33031e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_225_74#_c_1023_n 7.70291e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_1501_92#_M1031_g 0.0512647f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_1501_92#_c_1175_n 0.00214188f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_215 VPB N_A_1501_92#_c_1176_n 0.0128253f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_216 VPB N_A_1501_92#_c_1183_n 0.0134314f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.99
cc_217 VPB N_A_1501_92#_c_1178_n 0.00243604f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_218 VPB N_A_1501_92#_c_1185_n 0.0108998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_1339_74#_c_1274_n 0.010501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_1339_74#_c_1275_n 0.00495563f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.145
cc_221 VPB N_A_1339_74#_M1026_g 0.0243319f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_222 VPB N_A_1339_74#_M1008_g 0.0243291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_1339_74#_M1030_g 0.0244465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_1339_74#_M1015_g 0.0265411f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_1339_74#_c_1295_n 0.00170136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_1339_74#_c_1296_n 0.00684463f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_1339_74#_c_1287_n 0.0317634f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_1339_74#_c_1298_n 0.013245f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_1339_74#_c_1299_n 0.00363179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_1339_74#_c_1300_n 0.00904383f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_1339_74#_c_1301_n 0.00443161f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_1339_74#_c_1302_n 0.0048782f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_1339_74#_c_1288_n 7.82331e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_2221_74#_M1011_g 0.0238629f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_235 VPB N_A_2221_74#_M1014_g 0.0274022f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_236 VPB N_A_2221_74#_c_1463_n 0.014381f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_237 VPB N_A_27_74#_c_1530_n 0.0250181f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.98
cc_238 VPB N_A_27_74#_c_1535_n 0.0274742f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_239 VPB N_A_27_74#_c_1536_n 0.0257471f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_240 VPB N_A_27_74#_c_1537_n 0.0154585f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.295
cc_241 VPB N_A_27_74#_c_1531_n 0.00269752f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_A_27_74#_c_1539_n 0.0109364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1599_n 0.0169911f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1600_n 0.00646119f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1601_n 0.00578178f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1602_n 0.00906458f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1603_n 0.00808814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1604_n 0.0220673f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1605_n 0.0265971f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1606_n 0.0157534f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1607_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1608_n 0.0644823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1609_n 0.0559624f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1610_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1611_n 0.0179825f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1612_n 0.00487897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1613_n 0.0180274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1614_n 0.0215753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1615_n 0.049432f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1616_n 0.0312072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1617_n 0.0400196f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1618_n 0.0219379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1619_n 0.0203698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1620_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1621_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1622_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1623_n 0.00490136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1624_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1625_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1598_n 0.14639f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB Q_N 0.00107351f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.98
cc_272 VPB Q_N 0.00196166f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_273 VPB Q_N 0.00224648f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_Q_c_1779_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_275 VPB N_Q_c_1780_n 0.00447264f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_Q_c_1776_n 0.0010488f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.145
cc_277 N_D_c_278_n N_CLK_M1018_g 0.00408937f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_278 N_D_c_278_n N_CLK_c_314_n 0.00572583f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_279 N_D_c_280_n N_CLK_c_315_n 0.00232413f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_280 N_D_c_278_n N_A_225_74#_c_1002_n 0.003576f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_281 N_D_c_278_n N_A_225_74#_c_1020_n 0.00298111f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_282 N_D_M1029_g N_A_225_74#_c_1020_n 9.40485e-19 $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_283 N_D_c_281_n N_A_225_74#_c_1020_n 0.0224944f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_284 N_D_M1033_g N_A_225_74#_c_1004_n 0.00616966f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_285 N_D_c_280_n N_A_225_74#_c_1004_n 0.003576f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_286 N_D_c_281_n N_A_225_74#_c_1004_n 0.0556869f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_287 N_D_M1033_g N_A_27_74#_c_1529_n 0.00146243f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_288 N_D_M1033_g N_A_27_74#_c_1530_n 0.00600966f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_289 N_D_c_280_n N_A_27_74#_c_1530_n 0.0320429f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_290 N_D_c_281_n N_A_27_74#_c_1530_n 0.0697394f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_291 N_D_M1029_g N_A_27_74#_c_1535_n 0.0083684f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_292 N_D_M1029_g N_A_27_74#_c_1536_n 0.0218367f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_293 N_D_c_281_n N_A_27_74#_c_1536_n 0.0227191f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_294 N_D_c_285_n N_A_27_74#_c_1536_n 0.00140505f $X=0.64 $Y=1.825 $X2=0 $Y2=0
cc_295 N_D_M1029_g N_VPWR_c_1599_n 0.0148304f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_296 N_D_M1029_g N_VPWR_c_1613_n 0.00460063f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_297 N_D_M1029_g N_VPWR_c_1598_n 0.00912296f $X=0.505 $Y=2.75 $X2=0 $Y2=0
cc_298 N_D_M1033_g N_VGND_c_1809_n 0.0137856f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_299 N_D_c_280_n N_VGND_c_1809_n 0.00175174f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_300 N_D_c_281_n N_VGND_c_1809_n 0.0220022f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_301 N_D_M1033_g N_VGND_c_1820_n 0.00383152f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_302 N_D_M1033_g N_VGND_c_1834_n 0.00761198f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_303 CLK N_A_225_74#_M1019_g 0.00369616f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_304 N_CLK_c_314_n N_A_225_74#_M1019_g 0.0210236f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_305 N_CLK_c_315_n N_A_225_74#_M1019_g 0.0131368f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_306 N_CLK_M1018_g N_A_225_74#_M1021_g 0.0488038f $X=1.515 $Y=2.35 $X2=0 $Y2=0
cc_307 N_CLK_M1018_g N_A_225_74#_c_999_n 0.00479904f $X=1.515 $Y=2.35 $X2=0
+ $Y2=0
cc_308 N_CLK_M1018_g N_A_225_74#_c_1002_n 0.00354737f $X=1.515 $Y=2.35 $X2=0
+ $Y2=0
cc_309 CLK N_A_225_74#_c_1002_n 0.0286813f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_310 N_CLK_c_314_n N_A_225_74#_c_1002_n 0.00297156f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_311 N_CLK_c_315_n N_A_225_74#_c_1002_n 0.00330079f $X=1.465 $Y=1.22 $X2=0
+ $Y2=0
cc_312 N_CLK_c_314_n N_A_225_74#_c_1019_n 0.00313913f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_313 N_CLK_M1018_g N_A_225_74#_c_1021_n 0.009076f $X=1.515 $Y=2.35 $X2=0 $Y2=0
cc_314 N_CLK_c_314_n N_A_225_74#_c_1021_n 5.60514e-19 $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_315 N_CLK_M1018_g N_A_225_74#_c_1003_n 9.11681e-19 $X=1.515 $Y=2.35 $X2=0
+ $Y2=0
cc_316 CLK N_A_225_74#_c_1003_n 0.0203335f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_317 N_CLK_c_314_n N_A_225_74#_c_1003_n 2.00661e-19 $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_318 CLK N_A_225_74#_c_1004_n 0.00762435f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_319 N_CLK_c_314_n N_A_225_74#_c_1004_n 0.00114511f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_320 N_CLK_c_315_n N_A_225_74#_c_1004_n 0.00765617f $X=1.465 $Y=1.22 $X2=0
+ $Y2=0
cc_321 N_CLK_M1018_g N_A_225_74#_c_1023_n 0.00508679f $X=1.515 $Y=2.35 $X2=0
+ $Y2=0
cc_322 CLK N_A_225_74#_c_1023_n 0.0352423f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_323 N_CLK_M1018_g N_A_27_74#_c_1536_n 0.0177479f $X=1.515 $Y=2.35 $X2=0 $Y2=0
cc_324 CLK N_A_27_74#_c_1531_n 0.00324184f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_325 N_CLK_M1018_g N_VPWR_c_1599_n 0.0132363f $X=1.515 $Y=2.35 $X2=0 $Y2=0
cc_326 N_CLK_M1018_g N_VPWR_c_1600_n 0.025074f $X=1.515 $Y=2.35 $X2=0 $Y2=0
cc_327 N_CLK_M1018_g N_VPWR_c_1614_n 0.00540231f $X=1.515 $Y=2.35 $X2=0 $Y2=0
cc_328 N_CLK_M1018_g N_VPWR_c_1598_n 0.00533457f $X=1.515 $Y=2.35 $X2=0 $Y2=0
cc_329 N_CLK_c_315_n N_VGND_c_1809_n 0.00299692f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_330 N_CLK_c_315_n N_VGND_c_1810_n 0.00434272f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_331 CLK N_VGND_c_1811_n 0.0142803f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_332 N_CLK_c_315_n N_VGND_c_1811_n 0.00300619f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_333 N_CLK_c_315_n N_VGND_c_1834_n 0.00825157f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_334 N_A_398_74#_c_358_n N_A_757_401#_M1009_g 0.0105331f $X=3.735 $Y=1.6 $X2=0
+ $Y2=0
cc_335 N_A_398_74#_c_380_n N_A_757_401#_M1009_g 0.00869165f $X=3.735 $Y=2.905
+ $X2=0 $Y2=0
cc_336 N_A_398_74#_c_393_p N_A_757_401#_M1009_g 0.0106925f $X=4.52 $Y=2.48 $X2=0
+ $Y2=0
cc_337 N_A_398_74#_c_381_n N_A_757_401#_M1009_g 0.00277482f $X=4.605 $Y=2.905
+ $X2=0 $Y2=0
cc_338 N_A_398_74#_c_395_p N_A_757_401#_M1009_g 0.00209717f $X=3.735 $Y=2.48
+ $X2=0 $Y2=0
cc_339 N_A_398_74#_M1036_g N_A_757_401#_c_621_n 0.0485648f $X=3.58 $Y=0.695
+ $X2=0 $Y2=0
cc_340 N_A_398_74#_c_393_p N_A_757_401#_c_627_n 0.00464419f $X=4.52 $Y=2.48
+ $X2=0 $Y2=0
cc_341 N_A_398_74#_M1001_g N_A_757_401#_c_628_n 7.56368e-19 $X=3.005 $Y=2.525
+ $X2=0 $Y2=0
cc_342 N_A_398_74#_c_374_n N_A_757_401#_c_628_n 0.00105872f $X=2.95 $Y=2.105
+ $X2=0 $Y2=0
cc_343 N_A_398_74#_c_358_n N_A_757_401#_c_628_n 0.00634699f $X=3.735 $Y=1.6
+ $X2=0 $Y2=0
cc_344 N_A_398_74#_c_359_n N_A_757_401#_c_628_n 0.00700889f $X=3.735 $Y=1.6
+ $X2=0 $Y2=0
cc_345 N_A_398_74#_M1036_g N_A_757_401#_c_622_n 0.00296636f $X=3.58 $Y=0.695
+ $X2=0 $Y2=0
cc_346 N_A_398_74#_c_359_n N_A_757_401#_c_623_n 0.00158807f $X=3.735 $Y=1.6
+ $X2=0 $Y2=0
cc_347 N_A_398_74#_c_393_p N_A_757_401#_c_629_n 0.0160587f $X=4.52 $Y=2.48 $X2=0
+ $Y2=0
cc_348 N_A_398_74#_c_358_n N_A_757_401#_c_630_n 0.018204f $X=3.735 $Y=1.6 $X2=0
+ $Y2=0
cc_349 N_A_398_74#_c_393_p N_A_757_401#_c_630_n 0.0259281f $X=4.52 $Y=2.48 $X2=0
+ $Y2=0
cc_350 N_A_398_74#_c_358_n N_A_757_401#_c_631_n 0.00412226f $X=3.735 $Y=1.6
+ $X2=0 $Y2=0
cc_351 N_A_398_74#_c_393_p N_A_757_401#_c_631_n 0.00190513f $X=4.52 $Y=2.48
+ $X2=0 $Y2=0
cc_352 N_A_398_74#_M1036_g N_A_757_401#_c_624_n 3.1275e-19 $X=3.58 $Y=0.695
+ $X2=0 $Y2=0
cc_353 N_A_398_74#_c_382_n N_A_757_401#_c_632_n 0.0220094f $X=5.36 $Y=2.99 $X2=0
+ $Y2=0
cc_354 N_A_398_74#_c_386_n N_A_757_401#_c_632_n 0.00882225f $X=5.53 $Y=2.275
+ $X2=0 $Y2=0
cc_355 N_A_398_74#_c_358_n N_A_757_401#_c_625_n 0.00214471f $X=3.735 $Y=1.6
+ $X2=0 $Y2=0
cc_356 N_A_398_74#_c_359_n N_A_757_401#_c_625_n 0.00953288f $X=3.735 $Y=1.6
+ $X2=0 $Y2=0
cc_357 N_A_398_74#_c_364_n N_A_595_97#_M1017_d 0.00383506f $X=2.95 $Y=1.435
+ $X2=-0.19 $Y2=-0.245
cc_358 N_A_398_74#_c_381_n N_A_595_97#_M1020_g 0.00744321f $X=4.605 $Y=2.905
+ $X2=0 $Y2=0
cc_359 N_A_398_74#_c_382_n N_A_595_97#_M1020_g 0.00394744f $X=5.36 $Y=2.99 $X2=0
+ $Y2=0
cc_360 N_A_398_74#_c_384_n N_A_595_97#_M1020_g 5.16056e-19 $X=5.445 $Y=2.905
+ $X2=0 $Y2=0
cc_361 N_A_398_74#_c_384_n N_A_595_97#_M1006_g 0.00282974f $X=5.445 $Y=2.905
+ $X2=0 $Y2=0
cc_362 N_A_398_74#_c_385_n N_A_595_97#_M1006_g 0.019251f $X=6.33 $Y=2.275 $X2=0
+ $Y2=0
cc_363 N_A_398_74#_c_361_n N_A_595_97#_M1006_g 0.012049f $X=6.415 $Y=2.19 $X2=0
+ $Y2=0
cc_364 N_A_398_74#_c_360_n N_A_595_97#_c_712_n 0.00482959f $X=6.415 $Y=1.12
+ $X2=0 $Y2=0
cc_365 N_A_398_74#_c_363_n N_A_595_97#_c_712_n 0.00103022f $X=6.5 $Y=0.365 $X2=0
+ $Y2=0
cc_366 N_A_398_74#_c_368_n N_A_595_97#_c_712_n 0.0283274f $X=6.71 $Y=1.12 $X2=0
+ $Y2=0
cc_367 N_A_398_74#_c_365_n N_A_595_97#_c_713_n 0.00505169f $X=6.71 $Y=1.285
+ $X2=0 $Y2=0
cc_368 N_A_398_74#_c_366_n N_A_595_97#_c_713_n 0.0283274f $X=6.71 $Y=1.285 $X2=0
+ $Y2=0
cc_369 N_A_398_74#_M1036_g N_A_595_97#_c_714_n 0.00609952f $X=3.58 $Y=0.695
+ $X2=0 $Y2=0
cc_370 N_A_398_74#_c_364_n N_A_595_97#_c_714_n 0.0344769f $X=2.95 $Y=1.435 $X2=0
+ $Y2=0
cc_371 N_A_398_74#_M1036_g N_A_595_97#_c_715_n 0.00510302f $X=3.58 $Y=0.695
+ $X2=0 $Y2=0
cc_372 N_A_398_74#_c_364_n N_A_595_97#_c_715_n 0.0128205f $X=2.95 $Y=1.435 $X2=0
+ $Y2=0
cc_373 N_A_398_74#_c_370_n N_A_595_97#_c_716_n 0.00638833f $X=2.95 $Y=1.94 $X2=0
+ $Y2=0
cc_374 N_A_398_74#_M1001_g N_A_595_97#_c_716_n 0.00222137f $X=3.005 $Y=2.525
+ $X2=0 $Y2=0
cc_375 N_A_398_74#_c_352_n N_A_595_97#_c_716_n 0.0216127f $X=3.505 $Y=1.6 $X2=0
+ $Y2=0
cc_376 N_A_398_74#_M1036_g N_A_595_97#_c_716_n 0.00457084f $X=3.58 $Y=0.695
+ $X2=0 $Y2=0
cc_377 N_A_398_74#_c_357_n N_A_595_97#_c_716_n 0.0490068f $X=2.95 $Y=1.6 $X2=0
+ $Y2=0
cc_378 N_A_398_74#_c_358_n N_A_595_97#_c_716_n 0.0631091f $X=3.735 $Y=1.6 $X2=0
+ $Y2=0
cc_379 N_A_398_74#_c_364_n N_A_595_97#_c_716_n 0.0124678f $X=2.95 $Y=1.435 $X2=0
+ $Y2=0
cc_380 N_A_398_74#_M1036_g N_A_595_97#_c_717_n 0.0143046f $X=3.58 $Y=0.695 $X2=0
+ $Y2=0
cc_381 N_A_398_74#_c_358_n N_A_595_97#_c_717_n 0.0173132f $X=3.735 $Y=1.6 $X2=0
+ $Y2=0
cc_382 N_A_398_74#_c_359_n N_A_595_97#_c_717_n 0.00286357f $X=3.735 $Y=1.6 $X2=0
+ $Y2=0
cc_383 N_A_398_74#_M1036_g N_A_595_97#_c_718_n 0.0015524f $X=3.58 $Y=0.695 $X2=0
+ $Y2=0
cc_384 N_A_398_74#_c_358_n N_A_595_97#_c_718_n 0.00579354f $X=3.735 $Y=1.6 $X2=0
+ $Y2=0
cc_385 N_A_398_74#_c_359_n N_A_595_97#_c_718_n 7.68037e-19 $X=3.735 $Y=1.6 $X2=0
+ $Y2=0
cc_386 N_A_398_74#_c_358_n N_A_595_97#_c_720_n 0.0139492f $X=3.735 $Y=1.6 $X2=0
+ $Y2=0
cc_387 N_A_398_74#_c_359_n N_A_595_97#_c_720_n 0.00180184f $X=3.735 $Y=1.6 $X2=0
+ $Y2=0
cc_388 N_A_398_74#_M1001_g N_A_595_97#_c_732_n 0.00651612f $X=3.005 $Y=2.525
+ $X2=0 $Y2=0
cc_389 N_A_398_74#_c_352_n N_A_595_97#_c_732_n 0.0051059f $X=3.505 $Y=1.6 $X2=0
+ $Y2=0
cc_390 N_A_398_74#_c_375_n N_A_595_97#_c_732_n 0.0242202f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_391 N_A_398_74#_c_357_n N_A_595_97#_c_732_n 0.00373424f $X=2.95 $Y=1.6 $X2=0
+ $Y2=0
cc_392 N_A_398_74#_c_358_n N_A_595_97#_c_732_n 0.00757352f $X=3.735 $Y=1.6 $X2=0
+ $Y2=0
cc_393 N_A_398_74#_c_380_n N_A_595_97#_c_732_n 0.0129105f $X=3.735 $Y=2.905
+ $X2=0 $Y2=0
cc_394 N_A_398_74#_c_395_p N_A_595_97#_c_732_n 0.0142748f $X=3.735 $Y=2.48 $X2=0
+ $Y2=0
cc_395 N_A_398_74#_M1036_g N_A_595_97#_c_773_n 0.00254046f $X=3.58 $Y=0.695
+ $X2=0 $Y2=0
cc_396 N_A_398_74#_c_352_n N_A_595_97#_c_721_n 0.00220182f $X=3.505 $Y=1.6 $X2=0
+ $Y2=0
cc_397 N_A_398_74#_M1036_g N_A_595_97#_c_721_n 0.00428676f $X=3.58 $Y=0.695
+ $X2=0 $Y2=0
cc_398 N_A_398_74#_c_364_n N_A_595_97#_c_721_n 0.0140647f $X=2.95 $Y=1.435 $X2=0
+ $Y2=0
cc_399 N_A_398_74#_c_365_n N_A_595_97#_c_724_n 0.0126088f $X=6.71 $Y=1.285 $X2=0
+ $Y2=0
cc_400 N_A_398_74#_c_382_n N_SET_B_M1000_g 0.00332604f $X=5.36 $Y=2.99 $X2=0
+ $Y2=0
cc_401 N_A_398_74#_c_384_n N_SET_B_M1000_g 0.014868f $X=5.445 $Y=2.905 $X2=0
+ $Y2=0
cc_402 N_A_398_74#_c_386_n N_SET_B_M1000_g 0.00670868f $X=5.53 $Y=2.275 $X2=0
+ $Y2=0
cc_403 N_A_398_74#_c_367_n N_SET_B_c_872_n 0.00186884f $X=7.415 $Y=2.02 $X2=0
+ $Y2=0
cc_404 N_A_398_74#_c_385_n N_SET_B_c_878_n 0.0216423f $X=6.33 $Y=2.275 $X2=0
+ $Y2=0
cc_405 N_A_398_74#_c_361_n N_SET_B_c_878_n 0.0209674f $X=6.415 $Y=2.19 $X2=0
+ $Y2=0
cc_406 N_A_398_74#_c_365_n N_SET_B_c_878_n 0.0165581f $X=6.71 $Y=1.285 $X2=0
+ $Y2=0
cc_407 N_A_398_74#_c_366_n N_SET_B_c_878_n 0.00557641f $X=6.71 $Y=1.285 $X2=0
+ $Y2=0
cc_408 N_A_398_74#_c_388_n N_SET_B_c_878_n 0.00611943f $X=7.415 $Y=2.185 $X2=0
+ $Y2=0
cc_409 N_A_398_74#_c_367_n N_SET_B_c_878_n 0.0189131f $X=7.415 $Y=2.02 $X2=0
+ $Y2=0
cc_410 N_A_398_74#_c_390_n N_SET_B_c_878_n 5.97324e-19 $X=7.53 $Y=2.185 $X2=0
+ $Y2=0
cc_411 N_A_398_74#_c_385_n N_SET_B_c_879_n 0.00163184f $X=6.33 $Y=2.275 $X2=0
+ $Y2=0
cc_412 N_A_398_74#_c_386_n N_SET_B_c_879_n 7.6844e-19 $X=5.53 $Y=2.275 $X2=0
+ $Y2=0
cc_413 N_A_398_74#_c_385_n N_SET_B_c_880_n 0.00795886f $X=6.33 $Y=2.275 $X2=0
+ $Y2=0
cc_414 N_A_398_74#_c_386_n N_SET_B_c_880_n 0.0138178f $X=5.53 $Y=2.275 $X2=0
+ $Y2=0
cc_415 N_A_398_74#_c_386_n N_SET_B_c_891_n 9.89342e-19 $X=5.53 $Y=2.275 $X2=0
+ $Y2=0
cc_416 N_A_398_74#_c_354_n N_A_225_74#_M1019_g 0.00164183f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_417 N_A_398_74#_c_356_n N_A_225_74#_M1019_g 0.00266901f $X=2.215 $Y=0.34
+ $X2=0 $Y2=0
cc_418 N_A_398_74#_c_376_n N_A_225_74#_M1021_g 0.00132039f $X=2.275 $Y=2.99
+ $X2=0 $Y2=0
cc_419 N_A_398_74#_c_370_n N_A_225_74#_c_1006_n 0.019666f $X=2.95 $Y=1.94 $X2=0
+ $Y2=0
cc_420 N_A_398_74#_M1001_g N_A_225_74#_c_1006_n 0.0185309f $X=3.005 $Y=2.525
+ $X2=0 $Y2=0
cc_421 N_A_398_74#_c_478_p N_A_225_74#_c_1006_n 0.00605299f $X=2.19 $Y=2.665
+ $X2=0 $Y2=0
cc_422 N_A_398_74#_c_375_n N_A_225_74#_c_1006_n 0.0104492f $X=3.625 $Y=2.99
+ $X2=0 $Y2=0
cc_423 N_A_398_74#_c_357_n N_A_225_74#_c_1006_n 3.80029e-19 $X=2.95 $Y=1.6 $X2=0
+ $Y2=0
cc_424 N_A_398_74#_c_351_n N_A_225_74#_c_994_n 0.0105031f $X=2.95 $Y=1.765 $X2=0
+ $Y2=0
cc_425 N_A_398_74#_c_355_n N_A_225_74#_c_994_n 0.00132303f $X=2.94 $Y=0.34 $X2=0
+ $Y2=0
cc_426 N_A_398_74#_c_357_n N_A_225_74#_c_994_n 0.00111273f $X=2.95 $Y=1.6 $X2=0
+ $Y2=0
cc_427 N_A_398_74#_c_364_n N_A_225_74#_c_994_n 0.00549547f $X=2.95 $Y=1.435
+ $X2=0 $Y2=0
cc_428 N_A_398_74#_M1001_g N_A_225_74#_c_1007_n 0.0105864f $X=3.005 $Y=2.525
+ $X2=0 $Y2=0
cc_429 N_A_398_74#_c_375_n N_A_225_74#_c_1007_n 0.0116715f $X=3.625 $Y=2.99
+ $X2=0 $Y2=0
cc_430 N_A_398_74#_M1036_g N_A_225_74#_M1017_g 0.0110915f $X=3.58 $Y=0.695 $X2=0
+ $Y2=0
cc_431 N_A_398_74#_c_354_n N_A_225_74#_M1017_g 0.00397637f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_432 N_A_398_74#_c_355_n N_A_225_74#_M1017_g 0.0109068f $X=2.94 $Y=0.34 $X2=0
+ $Y2=0
cc_433 N_A_398_74#_c_364_n N_A_225_74#_M1017_g 0.0197485f $X=2.95 $Y=1.435 $X2=0
+ $Y2=0
cc_434 N_A_398_74#_M1001_g N_A_225_74#_M1005_g 0.0136242f $X=3.005 $Y=2.525
+ $X2=0 $Y2=0
cc_435 N_A_398_74#_c_352_n N_A_225_74#_M1005_g 0.00622413f $X=3.505 $Y=1.6 $X2=0
+ $Y2=0
cc_436 N_A_398_74#_c_375_n N_A_225_74#_M1005_g 0.017045f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_437 N_A_398_74#_c_358_n N_A_225_74#_M1005_g 0.00136341f $X=3.735 $Y=1.6 $X2=0
+ $Y2=0
cc_438 N_A_398_74#_c_380_n N_A_225_74#_M1005_g 0.00578433f $X=3.735 $Y=2.905
+ $X2=0 $Y2=0
cc_439 N_A_398_74#_c_395_p N_A_225_74#_M1005_g 0.00123784f $X=3.735 $Y=2.48
+ $X2=0 $Y2=0
cc_440 N_A_398_74#_c_375_n N_A_225_74#_c_1010_n 0.00603546f $X=3.625 $Y=2.99
+ $X2=0 $Y2=0
cc_441 N_A_398_74#_c_393_p N_A_225_74#_c_1010_n 0.00565527f $X=4.52 $Y=2.48
+ $X2=0 $Y2=0
cc_442 N_A_398_74#_c_382_n N_A_225_74#_c_1010_n 0.0139188f $X=5.36 $Y=2.99 $X2=0
+ $Y2=0
cc_443 N_A_398_74#_c_383_n N_A_225_74#_c_1010_n 0.00419347f $X=4.69 $Y=2.99
+ $X2=0 $Y2=0
cc_444 N_A_398_74#_M1010_g N_A_225_74#_M1027_g 0.0046362f $X=7.53 $Y=2.75 $X2=0
+ $Y2=0
cc_445 N_A_398_74#_c_385_n N_A_225_74#_M1027_g 0.0016151f $X=6.33 $Y=2.275 $X2=0
+ $Y2=0
cc_446 N_A_398_74#_c_367_n N_A_225_74#_M1027_g 6.92741e-19 $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_447 N_A_398_74#_c_390_n N_A_225_74#_c_996_n 0.00100919f $X=7.53 $Y=2.185
+ $X2=0 $Y2=0
cc_448 N_A_398_74#_c_361_n N_A_225_74#_c_997_n 0.0043502f $X=6.415 $Y=2.19 $X2=0
+ $Y2=0
cc_449 N_A_398_74#_c_365_n N_A_225_74#_c_997_n 0.00122906f $X=6.71 $Y=1.285
+ $X2=0 $Y2=0
cc_450 N_A_398_74#_c_366_n N_A_225_74#_c_997_n 0.0172932f $X=6.71 $Y=1.285 $X2=0
+ $Y2=0
cc_451 N_A_398_74#_c_361_n N_A_225_74#_M1037_g 9.168e-19 $X=6.415 $Y=2.19 $X2=0
+ $Y2=0
cc_452 N_A_398_74#_c_362_n N_A_225_74#_M1037_g 0.00565608f $X=7.385 $Y=0.365
+ $X2=0 $Y2=0
cc_453 N_A_398_74#_c_365_n N_A_225_74#_M1037_g 3.65769e-19 $X=6.71 $Y=1.285
+ $X2=0 $Y2=0
cc_454 N_A_398_74#_c_366_n N_A_225_74#_M1037_g 0.0180888f $X=6.71 $Y=1.285 $X2=0
+ $Y2=0
cc_455 N_A_398_74#_c_367_n N_A_225_74#_M1037_g 0.0107513f $X=7.415 $Y=2.02 $X2=0
+ $Y2=0
cc_456 N_A_398_74#_c_368_n N_A_225_74#_M1037_g 0.016767f $X=6.71 $Y=1.12 $X2=0
+ $Y2=0
cc_457 N_A_398_74#_c_351_n N_A_225_74#_c_1000_n 0.019666f $X=2.95 $Y=1.765 $X2=0
+ $Y2=0
cc_458 N_A_398_74#_c_354_n N_A_225_74#_c_1000_n 7.55533e-19 $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_459 N_A_398_74#_c_355_n N_A_225_74#_c_1000_n 9.27593e-19 $X=2.94 $Y=0.34
+ $X2=0 $Y2=0
cc_460 N_A_398_74#_c_357_n N_A_225_74#_c_1000_n 3.80029e-19 $X=2.95 $Y=1.6 $X2=0
+ $Y2=0
cc_461 N_A_398_74#_c_364_n N_A_225_74#_c_1000_n 8.1877e-19 $X=2.95 $Y=1.435
+ $X2=0 $Y2=0
cc_462 N_A_398_74#_c_354_n N_A_225_74#_c_1001_n 0.00105443f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_463 N_A_398_74#_M1021_d N_A_225_74#_c_1021_n 0.00277287f $X=2.055 $Y=1.79
+ $X2=0 $Y2=0
cc_464 N_A_398_74#_c_354_n N_A_225_74#_c_1003_n 0.0147852f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_465 N_A_398_74#_c_367_n N_A_1501_92#_M1023_g 0.0209879f $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_466 N_A_398_74#_c_388_n N_A_1501_92#_M1031_g 2.82185e-19 $X=7.415 $Y=2.185
+ $X2=0 $Y2=0
cc_467 N_A_398_74#_c_367_n N_A_1501_92#_M1031_g 0.00523185f $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_468 N_A_398_74#_c_390_n N_A_1501_92#_M1031_g 0.0561902f $X=7.53 $Y=2.185
+ $X2=0 $Y2=0
cc_469 N_A_398_74#_c_367_n N_A_1501_92#_c_1175_n 0.0563716f $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_470 N_A_398_74#_c_367_n N_A_1501_92#_c_1176_n 0.00557226f $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_471 N_A_398_74#_c_390_n N_A_1501_92#_c_1176_n 0.00343339f $X=7.53 $Y=2.185
+ $X2=0 $Y2=0
cc_472 N_A_398_74#_c_367_n N_A_1501_92#_c_1193_n 0.013418f $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_473 N_A_398_74#_c_362_n N_A_1339_74#_M1022_d 0.00226519f $X=7.385 $Y=0.365
+ $X2=-0.19 $Y2=-0.245
cc_474 N_A_398_74#_c_362_n N_A_1339_74#_c_1305_n 0.0335956f $X=7.385 $Y=0.365
+ $X2=0 $Y2=0
cc_475 N_A_398_74#_c_365_n N_A_1339_74#_c_1305_n 0.0135629f $X=6.71 $Y=1.285
+ $X2=0 $Y2=0
cc_476 N_A_398_74#_c_366_n N_A_1339_74#_c_1305_n 0.00395514f $X=6.71 $Y=1.285
+ $X2=0 $Y2=0
cc_477 N_A_398_74#_c_367_n N_A_1339_74#_c_1305_n 0.02548f $X=7.415 $Y=2.02 $X2=0
+ $Y2=0
cc_478 N_A_398_74#_c_368_n N_A_1339_74#_c_1305_n 0.00921999f $X=6.71 $Y=1.12
+ $X2=0 $Y2=0
cc_479 N_A_398_74#_M1010_g N_A_1339_74#_c_1295_n 0.00249406f $X=7.53 $Y=2.75
+ $X2=0 $Y2=0
cc_480 N_A_398_74#_c_385_n N_A_1339_74#_c_1295_n 0.00938849f $X=6.33 $Y=2.275
+ $X2=0 $Y2=0
cc_481 N_A_398_74#_c_361_n N_A_1339_74#_c_1295_n 0.0167305f $X=6.415 $Y=2.19
+ $X2=0 $Y2=0
cc_482 N_A_398_74#_c_388_n N_A_1339_74#_c_1295_n 0.0180759f $X=7.415 $Y=2.185
+ $X2=0 $Y2=0
cc_483 N_A_398_74#_c_367_n N_A_1339_74#_c_1295_n 0.00780712f $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_484 N_A_398_74#_c_390_n N_A_1339_74#_c_1295_n 0.00334148f $X=7.53 $Y=2.185
+ $X2=0 $Y2=0
cc_485 N_A_398_74#_c_360_n N_A_1339_74#_c_1286_n 0.00454611f $X=6.415 $Y=1.12
+ $X2=0 $Y2=0
cc_486 N_A_398_74#_c_361_n N_A_1339_74#_c_1286_n 0.0064862f $X=6.415 $Y=2.19
+ $X2=0 $Y2=0
cc_487 N_A_398_74#_c_365_n N_A_1339_74#_c_1286_n 0.0257548f $X=6.71 $Y=1.285
+ $X2=0 $Y2=0
cc_488 N_A_398_74#_c_366_n N_A_1339_74#_c_1286_n 9.90303e-19 $X=6.71 $Y=1.285
+ $X2=0 $Y2=0
cc_489 N_A_398_74#_c_367_n N_A_1339_74#_c_1286_n 0.0517761f $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_490 N_A_398_74#_c_368_n N_A_1339_74#_c_1286_n 0.00131891f $X=6.71 $Y=1.12
+ $X2=0 $Y2=0
cc_491 N_A_398_74#_c_361_n N_A_1339_74#_c_1299_n 0.00799661f $X=6.415 $Y=2.19
+ $X2=0 $Y2=0
cc_492 N_A_398_74#_c_365_n N_A_1339_74#_c_1299_n 0.00416021f $X=6.71 $Y=1.285
+ $X2=0 $Y2=0
cc_493 N_A_398_74#_c_366_n N_A_1339_74#_c_1299_n 3.84168e-19 $X=6.71 $Y=1.285
+ $X2=0 $Y2=0
cc_494 N_A_398_74#_c_367_n N_A_1339_74#_c_1299_n 0.012655f $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_495 N_A_398_74#_M1010_g N_A_1339_74#_c_1300_n 0.0108199f $X=7.53 $Y=2.75
+ $X2=0 $Y2=0
cc_496 N_A_398_74#_c_388_n N_A_1339_74#_c_1300_n 0.0262994f $X=7.415 $Y=2.185
+ $X2=0 $Y2=0
cc_497 N_A_398_74#_c_390_n N_A_1339_74#_c_1300_n 0.00460932f $X=7.53 $Y=2.185
+ $X2=0 $Y2=0
cc_498 N_A_398_74#_M1010_g N_A_1339_74#_c_1301_n 0.0106687f $X=7.53 $Y=2.75
+ $X2=0 $Y2=0
cc_499 N_A_398_74#_c_388_n N_A_1339_74#_c_1302_n 0.0244552f $X=7.415 $Y=2.185
+ $X2=0 $Y2=0
cc_500 N_A_398_74#_c_367_n N_A_1339_74#_c_1302_n 0.00525436f $X=7.415 $Y=2.02
+ $X2=0 $Y2=0
cc_501 N_A_398_74#_c_390_n N_A_1339_74#_c_1302_n 0.00695557f $X=7.53 $Y=2.185
+ $X2=0 $Y2=0
cc_502 N_A_398_74#_M1021_d N_A_27_74#_c_1537_n 0.00575804f $X=2.055 $Y=1.79
+ $X2=0 $Y2=0
cc_503 N_A_398_74#_M1001_g N_A_27_74#_c_1537_n 0.00235893f $X=3.005 $Y=2.525
+ $X2=0 $Y2=0
cc_504 N_A_398_74#_c_374_n N_A_27_74#_c_1537_n 8.6797e-19 $X=2.95 $Y=2.105 $X2=0
+ $Y2=0
cc_505 N_A_398_74#_c_478_p N_A_27_74#_c_1537_n 0.0385051f $X=2.19 $Y=2.665 $X2=0
+ $Y2=0
cc_506 N_A_398_74#_c_375_n N_A_27_74#_c_1537_n 0.0354334f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_507 N_A_398_74#_c_357_n N_A_27_74#_c_1537_n 0.0100447f $X=2.95 $Y=1.6 $X2=0
+ $Y2=0
cc_508 N_A_398_74#_c_351_n N_A_27_74#_c_1531_n 0.00362357f $X=2.95 $Y=1.765
+ $X2=0 $Y2=0
cc_509 N_A_398_74#_c_354_n N_A_27_74#_c_1531_n 0.0119039f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_510 N_A_398_74#_c_357_n N_A_27_74#_c_1531_n 0.0468227f $X=2.95 $Y=1.6 $X2=0
+ $Y2=0
cc_511 N_A_398_74#_c_364_n N_A_27_74#_c_1531_n 0.0228448f $X=2.95 $Y=1.435 $X2=0
+ $Y2=0
cc_512 N_A_398_74#_c_354_n N_A_27_74#_c_1533_n 0.0206338f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_513 N_A_398_74#_c_355_n N_A_27_74#_c_1533_n 0.0237903f $X=2.94 $Y=0.34 $X2=0
+ $Y2=0
cc_514 N_A_398_74#_c_364_n N_A_27_74#_c_1533_n 0.0119198f $X=2.95 $Y=1.435 $X2=0
+ $Y2=0
cc_515 N_A_398_74#_c_393_p N_VPWR_M1009_d 0.0152684f $X=4.52 $Y=2.48 $X2=0 $Y2=0
cc_516 N_A_398_74#_c_381_n N_VPWR_M1009_d 0.00408793f $X=4.605 $Y=2.905 $X2=0
+ $Y2=0
cc_517 N_A_398_74#_c_384_n N_VPWR_M1000_d 0.00481679f $X=5.445 $Y=2.905 $X2=0
+ $Y2=0
cc_518 N_A_398_74#_c_385_n N_VPWR_M1000_d 0.0151494f $X=6.33 $Y=2.275 $X2=0
+ $Y2=0
cc_519 N_A_398_74#_c_376_n N_VPWR_c_1600_n 0.0125862f $X=2.275 $Y=2.99 $X2=0
+ $Y2=0
cc_520 N_A_398_74#_c_375_n N_VPWR_c_1601_n 0.0147319f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_521 N_A_398_74#_c_380_n N_VPWR_c_1601_n 0.0129053f $X=3.735 $Y=2.905 $X2=0
+ $Y2=0
cc_522 N_A_398_74#_c_393_p N_VPWR_c_1601_n 0.0258766f $X=4.52 $Y=2.48 $X2=0
+ $Y2=0
cc_523 N_A_398_74#_c_381_n N_VPWR_c_1601_n 0.0134404f $X=4.605 $Y=2.905 $X2=0
+ $Y2=0
cc_524 N_A_398_74#_c_383_n N_VPWR_c_1601_n 0.0150385f $X=4.69 $Y=2.99 $X2=0
+ $Y2=0
cc_525 N_A_398_74#_c_382_n N_VPWR_c_1602_n 0.0151625f $X=5.36 $Y=2.99 $X2=0
+ $Y2=0
cc_526 N_A_398_74#_c_384_n N_VPWR_c_1602_n 0.0293714f $X=5.445 $Y=2.905 $X2=0
+ $Y2=0
cc_527 N_A_398_74#_c_385_n N_VPWR_c_1602_n 0.0298586f $X=6.33 $Y=2.275 $X2=0
+ $Y2=0
cc_528 N_A_398_74#_M1010_g N_VPWR_c_1609_n 0.00389302f $X=7.53 $Y=2.75 $X2=0
+ $Y2=0
cc_529 N_A_398_74#_c_375_n N_VPWR_c_1615_n 0.10093f $X=3.625 $Y=2.99 $X2=0 $Y2=0
cc_530 N_A_398_74#_c_376_n N_VPWR_c_1615_n 0.01218f $X=2.275 $Y=2.99 $X2=0 $Y2=0
cc_531 N_A_398_74#_c_382_n N_VPWR_c_1616_n 0.0546768f $X=5.36 $Y=2.99 $X2=0
+ $Y2=0
cc_532 N_A_398_74#_c_383_n N_VPWR_c_1616_n 0.0115893f $X=4.69 $Y=2.99 $X2=0
+ $Y2=0
cc_533 N_A_398_74#_M1010_g N_VPWR_c_1598_n 0.00497526f $X=7.53 $Y=2.75 $X2=0
+ $Y2=0
cc_534 N_A_398_74#_c_375_n N_VPWR_c_1598_n 0.0531785f $X=3.625 $Y=2.99 $X2=0
+ $Y2=0
cc_535 N_A_398_74#_c_376_n N_VPWR_c_1598_n 0.00660793f $X=2.275 $Y=2.99 $X2=0
+ $Y2=0
cc_536 N_A_398_74#_c_393_p N_VPWR_c_1598_n 0.0122156f $X=4.52 $Y=2.48 $X2=0
+ $Y2=0
cc_537 N_A_398_74#_c_382_n N_VPWR_c_1598_n 0.028344f $X=5.36 $Y=2.99 $X2=0 $Y2=0
cc_538 N_A_398_74#_c_383_n N_VPWR_c_1598_n 0.00583135f $X=4.69 $Y=2.99 $X2=0
+ $Y2=0
cc_539 N_A_398_74#_c_358_n A_709_463# 6.49096e-19 $X=3.735 $Y=1.6 $X2=-0.19
+ $Y2=-0.245
cc_540 N_A_398_74#_c_380_n A_709_463# 0.00138036f $X=3.735 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_541 N_A_398_74#_c_395_p A_709_463# 0.00144266f $X=3.735 $Y=2.48 $X2=-0.19
+ $Y2=-0.245
cc_542 N_A_398_74#_c_385_n A_1261_341# 0.00811299f $X=6.33 $Y=2.275 $X2=-0.19
+ $Y2=-0.245
cc_543 N_A_398_74#_c_361_n A_1261_341# 0.00725647f $X=6.415 $Y=2.19 $X2=-0.19
+ $Y2=-0.245
cc_544 N_A_398_74#_c_356_n N_VGND_c_1811_n 0.0110038f $X=2.215 $Y=0.34 $X2=0
+ $Y2=0
cc_545 N_A_398_74#_M1036_g N_VGND_c_1812_n 0.00159069f $X=3.58 $Y=0.695 $X2=0
+ $Y2=0
cc_546 N_A_398_74#_M1036_g N_VGND_c_1821_n 0.00476381f $X=3.58 $Y=0.695 $X2=0
+ $Y2=0
cc_547 N_A_398_74#_c_355_n N_VGND_c_1821_n 0.0588317f $X=2.94 $Y=0.34 $X2=0
+ $Y2=0
cc_548 N_A_398_74#_c_356_n N_VGND_c_1821_n 0.0121867f $X=2.215 $Y=0.34 $X2=0
+ $Y2=0
cc_549 N_A_398_74#_c_363_n N_VGND_c_1829_n 0.0113619f $X=6.5 $Y=0.365 $X2=0
+ $Y2=0
cc_550 N_A_398_74#_c_368_n N_VGND_c_1829_n 3.97182e-19 $X=6.71 $Y=1.12 $X2=0
+ $Y2=0
cc_551 N_A_398_74#_c_362_n N_VGND_c_1830_n 0.0593621f $X=7.385 $Y=0.365 $X2=0
+ $Y2=0
cc_552 N_A_398_74#_c_363_n N_VGND_c_1830_n 0.0105206f $X=6.5 $Y=0.365 $X2=0
+ $Y2=0
cc_553 N_A_398_74#_c_368_n N_VGND_c_1830_n 0.00281891f $X=6.71 $Y=1.12 $X2=0
+ $Y2=0
cc_554 N_A_398_74#_c_362_n N_VGND_c_1831_n 0.0070631f $X=7.385 $Y=0.365 $X2=0
+ $Y2=0
cc_555 N_A_398_74#_c_367_n N_VGND_c_1831_n 0.00572644f $X=7.415 $Y=2.02 $X2=0
+ $Y2=0
cc_556 N_A_398_74#_M1036_g N_VGND_c_1834_n 0.00509887f $X=3.58 $Y=0.695 $X2=0
+ $Y2=0
cc_557 N_A_398_74#_c_355_n N_VGND_c_1834_n 0.0338596f $X=2.94 $Y=0.34 $X2=0
+ $Y2=0
cc_558 N_A_398_74#_c_356_n N_VGND_c_1834_n 0.00660921f $X=2.215 $Y=0.34 $X2=0
+ $Y2=0
cc_559 N_A_398_74#_c_362_n N_VGND_c_1834_n 0.0385992f $X=7.385 $Y=0.365 $X2=0
+ $Y2=0
cc_560 N_A_398_74#_c_363_n N_VGND_c_1834_n 0.00652894f $X=6.5 $Y=0.365 $X2=0
+ $Y2=0
cc_561 N_A_398_74#_c_368_n N_VGND_c_1834_n 0.00358754f $X=6.71 $Y=1.12 $X2=0
+ $Y2=0
cc_562 N_A_398_74#_c_360_n A_1261_74# 0.00221695f $X=6.415 $Y=1.12 $X2=-0.19
+ $Y2=-0.245
cc_563 N_A_398_74#_c_367_n A_1453_118# 0.00353049f $X=7.415 $Y=2.02 $X2=-0.19
+ $Y2=-0.245
cc_564 N_A_757_401#_c_629_n N_A_595_97#_M1020_g 0.0133637f $X=4.86 $Y=2.14 $X2=0
+ $Y2=0
cc_565 N_A_757_401#_c_630_n N_A_595_97#_M1020_g 0.00146526f $X=4.305 $Y=1.99
+ $X2=0 $Y2=0
cc_566 N_A_757_401#_c_631_n N_A_595_97#_M1020_g 0.0152862f $X=4.305 $Y=1.99
+ $X2=0 $Y2=0
cc_567 N_A_757_401#_c_632_n N_A_595_97#_M1020_g 0.0150626f $X=5.025 $Y=2.14
+ $X2=0 $Y2=0
cc_568 N_A_757_401#_c_622_n N_A_595_97#_M1032_g 0.0201634f $X=4.295 $Y=1.09
+ $X2=0 $Y2=0
cc_569 N_A_757_401#_c_624_n N_A_595_97#_M1032_g 0.0194663f $X=4.715 $Y=0.58
+ $X2=0 $Y2=0
cc_570 N_A_757_401#_c_625_n N_A_595_97#_M1032_g 0.00519936f $X=4.305 $Y=1.825
+ $X2=0 $Y2=0
cc_571 N_A_757_401#_c_621_n N_A_595_97#_c_714_n 0.00117593f $X=3.94 $Y=1.015
+ $X2=0 $Y2=0
cc_572 N_A_757_401#_c_628_n N_A_595_97#_c_716_n 4.97762e-19 $X=3.965 $Y=2.08
+ $X2=0 $Y2=0
cc_573 N_A_757_401#_c_622_n N_A_595_97#_c_717_n 0.00856275f $X=4.295 $Y=1.09
+ $X2=0 $Y2=0
cc_574 N_A_757_401#_c_623_n N_A_595_97#_c_717_n 0.00961364f $X=4.015 $Y=1.09
+ $X2=0 $Y2=0
cc_575 N_A_757_401#_c_624_n N_A_595_97#_c_717_n 0.0137257f $X=4.715 $Y=0.58
+ $X2=0 $Y2=0
cc_576 N_A_757_401#_c_622_n N_A_595_97#_c_718_n 0.00316276f $X=4.295 $Y=1.09
+ $X2=0 $Y2=0
cc_577 N_A_757_401#_c_624_n N_A_595_97#_c_718_n 0.005833f $X=4.715 $Y=0.58 $X2=0
+ $Y2=0
cc_578 N_A_757_401#_c_622_n N_A_595_97#_c_719_n 0.00378094f $X=4.295 $Y=1.09
+ $X2=0 $Y2=0
cc_579 N_A_757_401#_c_629_n N_A_595_97#_c_719_n 0.0119117f $X=4.86 $Y=2.14 $X2=0
+ $Y2=0
cc_580 N_A_757_401#_c_630_n N_A_595_97#_c_719_n 0.0210386f $X=4.305 $Y=1.99
+ $X2=0 $Y2=0
cc_581 N_A_757_401#_c_631_n N_A_595_97#_c_719_n 0.00144642f $X=4.305 $Y=1.99
+ $X2=0 $Y2=0
cc_582 N_A_757_401#_c_624_n N_A_595_97#_c_719_n 0.0239403f $X=4.715 $Y=0.58
+ $X2=0 $Y2=0
cc_583 N_A_757_401#_c_625_n N_A_595_97#_c_719_n 0.0120775f $X=4.305 $Y=1.825
+ $X2=0 $Y2=0
cc_584 N_A_757_401#_c_627_n N_A_595_97#_c_720_n 0.00424988f $X=4.14 $Y=2.08
+ $X2=0 $Y2=0
cc_585 N_A_757_401#_c_630_n N_A_595_97#_c_720_n 0.0037144f $X=4.305 $Y=1.99
+ $X2=0 $Y2=0
cc_586 N_A_757_401#_c_631_n N_A_595_97#_c_720_n 5.49386e-19 $X=4.305 $Y=1.99
+ $X2=0 $Y2=0
cc_587 N_A_757_401#_M1009_g N_A_595_97#_c_732_n 3.68447e-19 $X=3.875 $Y=2.525
+ $X2=0 $Y2=0
cc_588 N_A_757_401#_c_623_n N_A_595_97#_c_773_n 0.00117593f $X=4.015 $Y=1.09
+ $X2=0 $Y2=0
cc_589 N_A_757_401#_c_622_n N_A_595_97#_c_722_n 6.62687e-19 $X=4.295 $Y=1.09
+ $X2=0 $Y2=0
cc_590 N_A_757_401#_c_629_n N_A_595_97#_c_722_n 0.00823228f $X=4.86 $Y=2.14
+ $X2=0 $Y2=0
cc_591 N_A_757_401#_c_630_n N_A_595_97#_c_722_n 0.00148595f $X=4.305 $Y=1.99
+ $X2=0 $Y2=0
cc_592 N_A_757_401#_c_631_n N_A_595_97#_c_722_n 2.79593e-19 $X=4.305 $Y=1.99
+ $X2=0 $Y2=0
cc_593 N_A_757_401#_c_624_n N_A_595_97#_c_722_n 0.017608f $X=4.715 $Y=0.58 $X2=0
+ $Y2=0
cc_594 N_A_757_401#_c_632_n N_A_595_97#_c_722_n 0.0135425f $X=5.025 $Y=2.14
+ $X2=0 $Y2=0
cc_595 N_A_757_401#_c_625_n N_A_595_97#_c_722_n 0.00244526f $X=4.305 $Y=1.825
+ $X2=0 $Y2=0
cc_596 N_A_757_401#_c_629_n N_A_595_97#_c_723_n 6.15625e-19 $X=4.86 $Y=2.14
+ $X2=0 $Y2=0
cc_597 N_A_757_401#_c_631_n N_A_595_97#_c_723_n 0.00379936f $X=4.305 $Y=1.99
+ $X2=0 $Y2=0
cc_598 N_A_757_401#_c_624_n N_A_595_97#_c_723_n 8.22799e-19 $X=4.715 $Y=0.58
+ $X2=0 $Y2=0
cc_599 N_A_757_401#_c_632_n N_A_595_97#_c_723_n 9.65695e-19 $X=5.025 $Y=2.14
+ $X2=0 $Y2=0
cc_600 N_A_757_401#_c_625_n N_A_595_97#_c_723_n 0.0150128f $X=4.305 $Y=1.825
+ $X2=0 $Y2=0
cc_601 N_A_757_401#_c_632_n N_A_595_97#_c_725_n 4.98461e-19 $X=5.025 $Y=2.14
+ $X2=0 $Y2=0
cc_602 N_A_757_401#_c_632_n N_SET_B_M1000_g 0.00679845f $X=5.025 $Y=2.14 $X2=0
+ $Y2=0
cc_603 N_A_757_401#_c_624_n N_SET_B_c_876_n 0.00257545f $X=4.715 $Y=0.58 $X2=0
+ $Y2=0
cc_604 N_A_757_401#_M1009_g N_A_225_74#_M1005_g 0.0338123f $X=3.875 $Y=2.525
+ $X2=0 $Y2=0
cc_605 N_A_757_401#_M1009_g N_A_225_74#_c_1010_n 0.0118682f $X=3.875 $Y=2.525
+ $X2=0 $Y2=0
cc_606 N_A_757_401#_M1009_g N_VPWR_c_1601_n 0.00302798f $X=3.875 $Y=2.525 $X2=0
+ $Y2=0
cc_607 N_A_757_401#_M1009_g N_VPWR_c_1598_n 7.53851e-19 $X=3.875 $Y=2.525 $X2=0
+ $Y2=0
cc_608 N_A_757_401#_c_621_n N_VGND_c_1812_n 0.0112772f $X=3.94 $Y=1.015 $X2=0
+ $Y2=0
cc_609 N_A_757_401#_c_622_n N_VGND_c_1812_n 0.00479662f $X=4.295 $Y=1.09 $X2=0
+ $Y2=0
cc_610 N_A_757_401#_c_624_n N_VGND_c_1812_n 0.0411686f $X=4.715 $Y=0.58 $X2=0
+ $Y2=0
cc_611 N_A_757_401#_c_621_n N_VGND_c_1821_n 0.00413255f $X=3.94 $Y=1.015 $X2=0
+ $Y2=0
cc_612 N_A_757_401#_c_624_n N_VGND_c_1828_n 0.0208755f $X=4.715 $Y=0.58 $X2=0
+ $Y2=0
cc_613 N_A_757_401#_c_624_n N_VGND_c_1829_n 0.0120077f $X=4.715 $Y=0.58 $X2=0
+ $Y2=0
cc_614 N_A_757_401#_c_621_n N_VGND_c_1834_n 0.00428305f $X=3.94 $Y=1.015 $X2=0
+ $Y2=0
cc_615 N_A_757_401#_c_624_n N_VGND_c_1834_n 0.0172297f $X=4.715 $Y=0.58 $X2=0
+ $Y2=0
cc_616 N_A_595_97#_M1006_g N_SET_B_M1000_g 0.0095631f $X=6.215 $Y=2.205 $X2=0
+ $Y2=0
cc_617 N_A_595_97#_M1032_g N_SET_B_c_876_n 0.0460006f $X=4.93 $Y=0.58 $X2=0
+ $Y2=0
cc_618 N_A_595_97#_c_725_n N_SET_B_c_877_n 3.91223e-19 $X=5.585 $Y=1.265 $X2=0
+ $Y2=0
cc_619 N_A_595_97#_c_710_n N_SET_B_c_878_n 0.0040413f $X=6.125 $Y=1.195 $X2=0
+ $Y2=0
cc_620 N_A_595_97#_M1006_g N_SET_B_c_878_n 0.0138145f $X=6.215 $Y=2.205 $X2=0
+ $Y2=0
cc_621 N_A_595_97#_c_724_n N_SET_B_c_878_n 0.010821f $X=5.75 $Y=1.285 $X2=0
+ $Y2=0
cc_622 N_A_595_97#_c_726_n N_SET_B_c_878_n 0.00611328f $X=5.75 $Y=1.195 $X2=0
+ $Y2=0
cc_623 N_A_595_97#_M1006_g N_SET_B_c_879_n 0.00155289f $X=6.215 $Y=2.205 $X2=0
+ $Y2=0
cc_624 N_A_595_97#_c_722_n N_SET_B_c_879_n 0.00204547f $X=4.882 $Y=1.325 $X2=0
+ $Y2=0
cc_625 N_A_595_97#_c_725_n N_SET_B_c_879_n 0.00882985f $X=5.585 $Y=1.265 $X2=0
+ $Y2=0
cc_626 N_A_595_97#_c_726_n N_SET_B_c_879_n 0.00215733f $X=5.75 $Y=1.195 $X2=0
+ $Y2=0
cc_627 N_A_595_97#_M1020_g N_SET_B_c_880_n 8.23032e-19 $X=4.8 $Y=2.525 $X2=0
+ $Y2=0
cc_628 N_A_595_97#_M1006_g N_SET_B_c_880_n 0.00744603f $X=6.215 $Y=2.205 $X2=0
+ $Y2=0
cc_629 N_A_595_97#_c_722_n N_SET_B_c_880_n 0.0182485f $X=4.882 $Y=1.325 $X2=0
+ $Y2=0
cc_630 N_A_595_97#_c_723_n N_SET_B_c_880_n 0.0010606f $X=4.85 $Y=1.72 $X2=0
+ $Y2=0
cc_631 N_A_595_97#_c_725_n N_SET_B_c_880_n 0.0282062f $X=5.585 $Y=1.265 $X2=0
+ $Y2=0
cc_632 N_A_595_97#_c_726_n N_SET_B_c_880_n 0.00114191f $X=5.75 $Y=1.195 $X2=0
+ $Y2=0
cc_633 N_A_595_97#_M1020_g N_SET_B_c_891_n 0.0261038f $X=4.8 $Y=2.525 $X2=0
+ $Y2=0
cc_634 N_A_595_97#_M1006_g N_SET_B_c_891_n 0.00521148f $X=6.215 $Y=2.205 $X2=0
+ $Y2=0
cc_635 N_A_595_97#_c_725_n N_SET_B_c_891_n 9.55679e-19 $X=5.585 $Y=1.265 $X2=0
+ $Y2=0
cc_636 N_A_595_97#_M1032_g N_SET_B_c_882_n 0.0317616f $X=4.93 $Y=0.58 $X2=0
+ $Y2=0
cc_637 N_A_595_97#_c_722_n N_SET_B_c_882_n 0.00434007f $X=4.882 $Y=1.325 $X2=0
+ $Y2=0
cc_638 N_A_595_97#_c_723_n N_SET_B_c_882_n 0.0197563f $X=4.85 $Y=1.72 $X2=0
+ $Y2=0
cc_639 N_A_595_97#_c_724_n N_SET_B_c_882_n 7.95332e-19 $X=5.75 $Y=1.285 $X2=0
+ $Y2=0
cc_640 N_A_595_97#_c_725_n N_SET_B_c_882_n 0.0131004f $X=5.585 $Y=1.265 $X2=0
+ $Y2=0
cc_641 N_A_595_97#_c_726_n N_SET_B_c_882_n 0.0208717f $X=5.75 $Y=1.195 $X2=0
+ $Y2=0
cc_642 N_A_595_97#_c_732_n N_A_225_74#_c_1006_n 3.02281e-19 $X=3.37 $Y=2.515
+ $X2=0 $Y2=0
cc_643 N_A_595_97#_c_721_n N_A_225_74#_c_994_n 3.39751e-19 $X=3.407 $Y=1.18
+ $X2=0 $Y2=0
cc_644 N_A_595_97#_c_714_n N_A_225_74#_M1017_g 0.001333f $X=3.365 $Y=0.695 $X2=0
+ $Y2=0
cc_645 N_A_595_97#_c_715_n N_A_225_74#_M1017_g 4.88269e-19 $X=3.407 $Y=1.095
+ $X2=0 $Y2=0
cc_646 N_A_595_97#_c_716_n N_A_225_74#_M1005_g 0.00398609f $X=3.37 $Y=2.295
+ $X2=0 $Y2=0
cc_647 N_A_595_97#_c_732_n N_A_225_74#_M1005_g 0.00875861f $X=3.37 $Y=2.515
+ $X2=0 $Y2=0
cc_648 N_A_595_97#_M1020_g N_A_225_74#_c_1010_n 0.0105864f $X=4.8 $Y=2.525 $X2=0
+ $Y2=0
cc_649 N_A_595_97#_M1006_g N_A_225_74#_c_1010_n 0.0108881f $X=6.215 $Y=2.205
+ $X2=0 $Y2=0
cc_650 N_A_595_97#_M1006_g N_A_225_74#_c_997_n 0.0402996f $X=6.215 $Y=2.205
+ $X2=0 $Y2=0
cc_651 N_A_595_97#_M1006_g N_A_1339_74#_c_1295_n 8.31258e-19 $X=6.215 $Y=2.205
+ $X2=0 $Y2=0
cc_652 N_A_595_97#_M1006_g N_A_1339_74#_c_1300_n 0.00163913f $X=6.215 $Y=2.205
+ $X2=0 $Y2=0
cc_653 N_A_595_97#_c_716_n N_A_27_74#_c_1537_n 0.00584669f $X=3.37 $Y=2.295
+ $X2=0 $Y2=0
cc_654 N_A_595_97#_c_732_n N_A_27_74#_c_1537_n 0.0156328f $X=3.37 $Y=2.515 $X2=0
+ $Y2=0
cc_655 N_A_595_97#_M1006_g N_VPWR_c_1602_n 0.0059048f $X=6.215 $Y=2.205 $X2=0
+ $Y2=0
cc_656 N_A_595_97#_M1006_g N_VPWR_c_1598_n 0.00113998f $X=6.215 $Y=2.205 $X2=0
+ $Y2=0
cc_657 N_A_595_97#_M1032_g N_VGND_c_1812_n 0.00316744f $X=4.93 $Y=0.58 $X2=0
+ $Y2=0
cc_658 N_A_595_97#_c_714_n N_VGND_c_1812_n 0.0121682f $X=3.365 $Y=0.695 $X2=0
+ $Y2=0
cc_659 N_A_595_97#_c_717_n N_VGND_c_1812_n 0.0102353f $X=4.015 $Y=1.18 $X2=0
+ $Y2=0
cc_660 N_A_595_97#_c_719_n N_VGND_c_1812_n 0.00161263f $X=4.75 $Y=1.6 $X2=0
+ $Y2=0
cc_661 N_A_595_97#_c_714_n N_VGND_c_1821_n 0.00747853f $X=3.365 $Y=0.695 $X2=0
+ $Y2=0
cc_662 N_A_595_97#_M1032_g N_VGND_c_1828_n 0.00433139f $X=4.93 $Y=0.58 $X2=0
+ $Y2=0
cc_663 N_A_595_97#_M1032_g N_VGND_c_1829_n 0.00145723f $X=4.93 $Y=0.58 $X2=0
+ $Y2=0
cc_664 N_A_595_97#_c_712_n N_VGND_c_1829_n 0.00739087f $X=6.23 $Y=1.12 $X2=0
+ $Y2=0
cc_665 N_A_595_97#_c_724_n N_VGND_c_1829_n 0.0129342f $X=5.75 $Y=1.285 $X2=0
+ $Y2=0
cc_666 N_A_595_97#_c_725_n N_VGND_c_1829_n 0.0072628f $X=5.585 $Y=1.265 $X2=0
+ $Y2=0
cc_667 N_A_595_97#_c_726_n N_VGND_c_1829_n 0.0129788f $X=5.75 $Y=1.195 $X2=0
+ $Y2=0
cc_668 N_A_595_97#_c_712_n N_VGND_c_1830_n 0.00292261f $X=6.23 $Y=1.12 $X2=0
+ $Y2=0
cc_669 N_A_595_97#_M1032_g N_VGND_c_1834_n 0.00822f $X=4.93 $Y=0.58 $X2=0 $Y2=0
cc_670 N_A_595_97#_c_712_n N_VGND_c_1834_n 0.00872613f $X=6.23 $Y=1.12 $X2=0
+ $Y2=0
cc_671 N_A_595_97#_c_714_n N_VGND_c_1834_n 0.00847688f $X=3.365 $Y=0.695 $X2=0
+ $Y2=0
cc_672 N_SET_B_M1000_g N_A_225_74#_c_1010_n 0.0108634f $X=5.315 $Y=2.525 $X2=0
+ $Y2=0
cc_673 N_SET_B_c_878_n N_A_225_74#_c_996_n 0.00362468f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_674 N_SET_B_c_878_n N_A_225_74#_c_997_n 0.00687396f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_675 N_SET_B_c_878_n N_A_225_74#_M1037_g 0.00266496f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_676 N_SET_B_c_872_n N_A_1501_92#_M1023_g 0.0389792f $X=7.97 $Y=1.09 $X2=0
+ $Y2=0
cc_677 N_SET_B_c_883_n N_A_1501_92#_M1023_g 0.00214118f $X=8.475 $Y=1.165 $X2=0
+ $Y2=0
cc_678 N_SET_B_M1034_g N_A_1501_92#_M1031_g 0.0452756f $X=8.4 $Y=2.75 $X2=0
+ $Y2=0
cc_679 N_SET_B_c_872_n N_A_1501_92#_c_1175_n 0.00272879f $X=7.97 $Y=1.09 $X2=0
+ $Y2=0
cc_680 N_SET_B_c_873_n N_A_1501_92#_c_1175_n 0.00543494f $X=8.31 $Y=1.165 $X2=0
+ $Y2=0
cc_681 N_SET_B_c_874_n N_A_1501_92#_c_1175_n 0.00453006f $X=8.045 $Y=1.165 $X2=0
+ $Y2=0
cc_682 N_SET_B_c_878_n N_A_1501_92#_c_1175_n 0.0259693f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_683 SET_B N_A_1501_92#_c_1175_n 0.00256053f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_684 N_SET_B_c_883_n N_A_1501_92#_c_1175_n 0.00140589f $X=8.475 $Y=1.165 $X2=0
+ $Y2=0
cc_685 N_SET_B_c_884_n N_A_1501_92#_c_1175_n 0.0354924f $X=8.475 $Y=1.345 $X2=0
+ $Y2=0
cc_686 N_SET_B_c_874_n N_A_1501_92#_c_1176_n 0.0104285f $X=8.045 $Y=1.165 $X2=0
+ $Y2=0
cc_687 N_SET_B_c_878_n N_A_1501_92#_c_1176_n 0.01006f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_688 SET_B N_A_1501_92#_c_1176_n 0.00139253f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_689 N_SET_B_c_883_n N_A_1501_92#_c_1176_n 0.0171448f $X=8.475 $Y=1.165 $X2=0
+ $Y2=0
cc_690 N_SET_B_c_884_n N_A_1501_92#_c_1176_n 0.00179807f $X=8.475 $Y=1.345 $X2=0
+ $Y2=0
cc_691 N_SET_B_c_873_n N_A_1501_92#_c_1209_n 0.0175303f $X=8.31 $Y=1.165 $X2=0
+ $Y2=0
cc_692 N_SET_B_c_878_n N_A_1501_92#_c_1209_n 0.00610939f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_693 SET_B N_A_1501_92#_c_1209_n 0.00196951f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_694 N_SET_B_c_884_n N_A_1501_92#_c_1209_n 0.0268551f $X=8.475 $Y=1.345 $X2=0
+ $Y2=0
cc_695 N_SET_B_c_872_n N_A_1501_92#_c_1193_n 0.0115671f $X=7.97 $Y=1.09 $X2=0
+ $Y2=0
cc_696 N_SET_B_M1034_g N_A_1501_92#_c_1185_n 0.00116659f $X=8.4 $Y=2.75 $X2=0
+ $Y2=0
cc_697 N_SET_B_c_883_n N_A_1339_74#_M1003_g 0.0217685f $X=8.475 $Y=1.165 $X2=0
+ $Y2=0
cc_698 N_SET_B_c_884_n N_A_1339_74#_M1003_g 0.00107899f $X=8.475 $Y=1.345 $X2=0
+ $Y2=0
cc_699 N_SET_B_M1034_g N_A_1339_74#_c_1275_n 0.00455626f $X=8.4 $Y=2.75 $X2=0
+ $Y2=0
cc_700 N_SET_B_c_884_n N_A_1339_74#_c_1275_n 9.08428e-19 $X=8.475 $Y=1.345 $X2=0
+ $Y2=0
cc_701 N_SET_B_c_878_n N_A_1339_74#_c_1295_n 0.00158223f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_702 N_SET_B_c_878_n N_A_1339_74#_c_1286_n 0.0132819f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_703 N_SET_B_M1034_g N_A_1339_74#_c_1296_n 0.0193931f $X=8.4 $Y=2.75 $X2=0
+ $Y2=0
cc_704 N_SET_B_c_878_n N_A_1339_74#_c_1296_n 0.00979116f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_705 SET_B N_A_1339_74#_c_1296_n 0.0030363f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_706 N_SET_B_c_884_n N_A_1339_74#_c_1296_n 0.0116201f $X=8.475 $Y=1.345 $X2=0
+ $Y2=0
cc_707 N_SET_B_M1034_g N_A_1339_74#_c_1287_n 0.0194714f $X=8.4 $Y=2.75 $X2=0
+ $Y2=0
cc_708 SET_B N_A_1339_74#_c_1287_n 0.00218127f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_709 N_SET_B_c_883_n N_A_1339_74#_c_1287_n 0.00125511f $X=8.475 $Y=1.165 $X2=0
+ $Y2=0
cc_710 N_SET_B_c_884_n N_A_1339_74#_c_1287_n 0.0392467f $X=8.475 $Y=1.345 $X2=0
+ $Y2=0
cc_711 N_SET_B_M1034_g N_A_1339_74#_c_1298_n 0.00814108f $X=8.4 $Y=2.75 $X2=0
+ $Y2=0
cc_712 N_SET_B_c_878_n N_A_1339_74#_c_1299_n 0.0177625f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_713 N_SET_B_M1034_g N_A_1339_74#_c_1302_n 4.5108e-19 $X=8.4 $Y=2.75 $X2=0
+ $Y2=0
cc_714 N_SET_B_c_878_n N_A_1339_74#_c_1302_n 0.00223482f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_715 N_SET_B_c_878_n N_VPWR_M1000_d 0.00286361f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_716 N_SET_B_M1000_g N_VPWR_c_1602_n 0.00121603f $X=5.315 $Y=2.525 $X2=0 $Y2=0
cc_717 N_SET_B_M1034_g N_VPWR_c_1603_n 0.00308998f $X=8.4 $Y=2.75 $X2=0 $Y2=0
cc_718 N_SET_B_M1034_g N_VPWR_c_1617_n 0.00522561f $X=8.4 $Y=2.75 $X2=0 $Y2=0
cc_719 N_SET_B_M1034_g N_VPWR_c_1598_n 0.00542307f $X=8.4 $Y=2.75 $X2=0 $Y2=0
cc_720 N_SET_B_c_878_n A_1261_341# 0.00239809f $X=8.255 $Y=1.665 $X2=-0.19
+ $Y2=-0.245
cc_721 N_SET_B_c_876_n N_VGND_c_1828_n 0.00383152f $X=5.295 $Y=0.865 $X2=0 $Y2=0
cc_722 N_SET_B_c_876_n N_VGND_c_1829_n 0.0116257f $X=5.295 $Y=0.865 $X2=0 $Y2=0
cc_723 N_SET_B_c_872_n N_VGND_c_1830_n 0.00434252f $X=7.97 $Y=1.09 $X2=0 $Y2=0
cc_724 N_SET_B_c_872_n N_VGND_c_1831_n 0.00536598f $X=7.97 $Y=1.09 $X2=0 $Y2=0
cc_725 N_SET_B_c_872_n N_VGND_c_1834_n 0.00479212f $X=7.97 $Y=1.09 $X2=0 $Y2=0
cc_726 N_SET_B_c_876_n N_VGND_c_1834_n 0.00752325f $X=5.295 $Y=0.865 $X2=0 $Y2=0
cc_727 N_A_225_74#_M1037_g N_A_1501_92#_M1023_g 0.0562485f $X=7.19 $Y=0.8 $X2=0
+ $Y2=0
cc_728 N_A_225_74#_c_996_n N_A_1501_92#_M1031_g 3.89004e-19 $X=7.115 $Y=1.735
+ $X2=0 $Y2=0
cc_729 N_A_225_74#_M1037_g N_A_1501_92#_c_1176_n 0.00477807f $X=7.19 $Y=0.8
+ $X2=0 $Y2=0
cc_730 N_A_225_74#_M1037_g N_A_1339_74#_c_1305_n 0.0111291f $X=7.19 $Y=0.8 $X2=0
+ $Y2=0
cc_731 N_A_225_74#_M1027_g N_A_1339_74#_c_1295_n 0.0116581f $X=6.72 $Y=2.46
+ $X2=0 $Y2=0
cc_732 N_A_225_74#_c_996_n N_A_1339_74#_c_1295_n 0.00229379f $X=7.115 $Y=1.735
+ $X2=0 $Y2=0
cc_733 N_A_225_74#_c_996_n N_A_1339_74#_c_1286_n 0.00233299f $X=7.115 $Y=1.735
+ $X2=0 $Y2=0
cc_734 N_A_225_74#_M1037_g N_A_1339_74#_c_1286_n 0.0164602f $X=7.19 $Y=0.8 $X2=0
+ $Y2=0
cc_735 N_A_225_74#_M1027_g N_A_1339_74#_c_1299_n 0.00144122f $X=6.72 $Y=2.46
+ $X2=0 $Y2=0
cc_736 N_A_225_74#_c_996_n N_A_1339_74#_c_1299_n 0.0144662f $X=7.115 $Y=1.735
+ $X2=0 $Y2=0
cc_737 N_A_225_74#_c_997_n N_A_1339_74#_c_1299_n 0.00165844f $X=6.81 $Y=1.735
+ $X2=0 $Y2=0
cc_738 N_A_225_74#_M1027_g N_A_1339_74#_c_1300_n 0.0153547f $X=6.72 $Y=2.46
+ $X2=0 $Y2=0
cc_739 N_A_225_74#_c_996_n N_A_1339_74#_c_1300_n 0.00199244f $X=7.115 $Y=1.735
+ $X2=0 $Y2=0
cc_740 N_A_225_74#_M1018_s N_A_27_74#_c_1536_n 0.0117593f $X=1.145 $Y=1.79 $X2=0
+ $Y2=0
cc_741 N_A_225_74#_c_1019_n N_A_27_74#_c_1536_n 0.0189258f $X=1.305 $Y=1.87
+ $X2=0 $Y2=0
cc_742 N_A_225_74#_c_1020_n N_A_27_74#_c_1536_n 0.0142272f $X=1.145 $Y=1.87
+ $X2=0 $Y2=0
cc_743 N_A_225_74#_c_1021_n N_A_27_74#_c_1536_n 0.00643406f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_744 N_A_225_74#_M1021_g N_A_27_74#_c_1537_n 0.0165916f $X=1.965 $Y=2.35 $X2=0
+ $Y2=0
cc_745 N_A_225_74#_c_1006_n N_A_27_74#_c_1537_n 0.0254037f $X=2.485 $Y=3.075
+ $X2=0 $Y2=0
cc_746 N_A_225_74#_c_1001_n N_A_27_74#_c_1537_n 0.00180813f $X=2.41 $Y=1.465
+ $X2=0 $Y2=0
cc_747 N_A_225_74#_c_1021_n N_A_27_74#_c_1537_n 0.0277303f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_748 N_A_225_74#_M1019_g N_A_27_74#_c_1531_n 7.39226e-19 $X=1.915 $Y=0.74
+ $X2=0 $Y2=0
cc_749 N_A_225_74#_M1021_g N_A_27_74#_c_1531_n 0.00119828f $X=1.965 $Y=2.35
+ $X2=0 $Y2=0
cc_750 N_A_225_74#_c_1006_n N_A_27_74#_c_1531_n 0.00985083f $X=2.485 $Y=3.075
+ $X2=0 $Y2=0
cc_751 N_A_225_74#_c_994_n N_A_27_74#_c_1531_n 0.00583176f $X=2.825 $Y=1.12
+ $X2=0 $Y2=0
cc_752 N_A_225_74#_M1017_g N_A_27_74#_c_1531_n 0.00236295f $X=2.9 $Y=0.695 $X2=0
+ $Y2=0
cc_753 N_A_225_74#_c_1000_n N_A_27_74#_c_1531_n 0.0188485f $X=2.485 $Y=1.12
+ $X2=0 $Y2=0
cc_754 N_A_225_74#_c_1021_n N_A_27_74#_c_1531_n 0.0135406f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_755 N_A_225_74#_c_1003_n N_A_27_74#_c_1531_n 0.0302859f $X=2.11 $Y=1.465
+ $X2=0 $Y2=0
cc_756 N_A_225_74#_M1021_g N_A_27_74#_c_1581_n 0.00187706f $X=1.965 $Y=2.35
+ $X2=0 $Y2=0
cc_757 N_A_225_74#_c_1021_n N_A_27_74#_c_1581_n 0.0100622f $X=1.945 $Y=1.805
+ $X2=0 $Y2=0
cc_758 N_A_225_74#_c_994_n N_A_27_74#_c_1533_n 0.00610954f $X=2.825 $Y=1.12
+ $X2=0 $Y2=0
cc_759 N_A_225_74#_M1017_g N_A_27_74#_c_1533_n 4.22296e-19 $X=2.9 $Y=0.695 $X2=0
+ $Y2=0
cc_760 N_A_225_74#_c_1000_n N_A_27_74#_c_1533_n 9.83875e-19 $X=2.485 $Y=1.12
+ $X2=0 $Y2=0
cc_761 N_A_225_74#_c_1021_n N_VPWR_M1018_d 0.00164828f $X=1.945 $Y=1.805 $X2=0
+ $Y2=0
cc_762 N_A_225_74#_M1021_g N_VPWR_c_1600_n 0.00884461f $X=1.965 $Y=2.35 $X2=0
+ $Y2=0
cc_763 N_A_225_74#_c_1006_n N_VPWR_c_1600_n 3.19321e-19 $X=2.485 $Y=3.075 $X2=0
+ $Y2=0
cc_764 N_A_225_74#_c_1008_n N_VPWR_c_1600_n 0.00272925f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_765 N_A_225_74#_M1005_g N_VPWR_c_1601_n 7.29299e-19 $X=3.455 $Y=2.525 $X2=0
+ $Y2=0
cc_766 N_A_225_74#_c_1010_n N_VPWR_c_1601_n 0.0250524f $X=6.63 $Y=3.15 $X2=0
+ $Y2=0
cc_767 N_A_225_74#_c_1010_n N_VPWR_c_1602_n 0.027981f $X=6.63 $Y=3.15 $X2=0
+ $Y2=0
cc_768 N_A_225_74#_M1027_g N_VPWR_c_1602_n 0.00672258f $X=6.72 $Y=2.46 $X2=0
+ $Y2=0
cc_769 N_A_225_74#_c_1010_n N_VPWR_c_1609_n 0.0266714f $X=6.63 $Y=3.15 $X2=0
+ $Y2=0
cc_770 N_A_225_74#_M1021_g N_VPWR_c_1615_n 0.00540231f $X=1.965 $Y=2.35 $X2=0
+ $Y2=0
cc_771 N_A_225_74#_c_1008_n N_VPWR_c_1615_n 0.0372177f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_772 N_A_225_74#_c_1010_n N_VPWR_c_1616_n 0.0322942f $X=6.63 $Y=3.15 $X2=0
+ $Y2=0
cc_773 N_A_225_74#_M1021_g N_VPWR_c_1598_n 0.00533457f $X=1.965 $Y=2.35 $X2=0
+ $Y2=0
cc_774 N_A_225_74#_c_1007_n N_VPWR_c_1598_n 0.0189646f $X=3.365 $Y=3.15 $X2=0
+ $Y2=0
cc_775 N_A_225_74#_c_1008_n N_VPWR_c_1598_n 0.00604517f $X=2.56 $Y=3.15 $X2=0
+ $Y2=0
cc_776 N_A_225_74#_c_1010_n N_VPWR_c_1598_n 0.0883164f $X=6.63 $Y=3.15 $X2=0
+ $Y2=0
cc_777 N_A_225_74#_c_1017_n N_VPWR_c_1598_n 0.00445015f $X=3.455 $Y=3.15 $X2=0
+ $Y2=0
cc_778 N_A_225_74#_c_1004_n N_VGND_c_1809_n 0.0363632f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_779 N_A_225_74#_c_1004_n N_VGND_c_1810_n 0.0203368f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_780 N_A_225_74#_M1019_g N_VGND_c_1811_n 0.0115939f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_781 N_A_225_74#_c_1004_n N_VGND_c_1811_n 0.0268179f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_782 N_A_225_74#_M1019_g N_VGND_c_1821_n 0.00383152f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_783 N_A_225_74#_M1017_g N_VGND_c_1821_n 7.53287e-19 $X=2.9 $Y=0.695 $X2=0
+ $Y2=0
cc_784 N_A_225_74#_M1019_g N_VGND_c_1834_n 0.00762539f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_785 N_A_225_74#_c_1004_n N_VGND_c_1834_n 0.0167889f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_786 N_A_1501_92#_c_1209_n N_A_1339_74#_M1003_g 0.0152859f $X=9.105 $Y=0.925
+ $X2=0 $Y2=0
cc_787 N_A_1501_92#_c_1178_n N_A_1339_74#_M1003_g 0.00338973f $X=9.825 $Y=2.29
+ $X2=0 $Y2=0
cc_788 N_A_1501_92#_c_1179_n N_A_1339_74#_M1003_g 0.00714524f $X=9.27 $Y=0.8
+ $X2=0 $Y2=0
cc_789 N_A_1501_92#_c_1179_n N_A_1339_74#_c_1274_n 0.00226353f $X=9.27 $Y=0.8
+ $X2=0 $Y2=0
cc_790 N_A_1501_92#_c_1185_n N_A_1339_74#_c_1275_n 9.92746e-19 $X=9.18 $Y=2.375
+ $X2=0 $Y2=0
cc_791 N_A_1501_92#_c_1183_n N_A_1339_74#_M1026_g 0.00980989f $X=9.74 $Y=2.375
+ $X2=0 $Y2=0
cc_792 N_A_1501_92#_c_1185_n N_A_1339_74#_M1026_g 9.23576e-19 $X=9.18 $Y=2.375
+ $X2=0 $Y2=0
cc_793 N_A_1501_92#_c_1183_n N_A_1339_74#_c_1276_n 0.00165546f $X=9.74 $Y=2.375
+ $X2=0 $Y2=0
cc_794 N_A_1501_92#_c_1178_n N_A_1339_74#_c_1276_n 0.0184193f $X=9.825 $Y=2.29
+ $X2=0 $Y2=0
cc_795 N_A_1501_92#_c_1178_n N_A_1339_74#_M1008_g 0.00473493f $X=9.825 $Y=2.29
+ $X2=0 $Y2=0
cc_796 N_A_1501_92#_c_1185_n N_A_1339_74#_M1008_g 0.0038423f $X=9.18 $Y=2.375
+ $X2=0 $Y2=0
cc_797 N_A_1501_92#_c_1177_n N_A_1339_74#_M1013_g 0.00412514f $X=9.74 $Y=1.095
+ $X2=0 $Y2=0
cc_798 N_A_1501_92#_c_1178_n N_A_1339_74#_M1013_g 0.00391208f $X=9.825 $Y=2.29
+ $X2=0 $Y2=0
cc_799 N_A_1501_92#_c_1179_n N_A_1339_74#_M1013_g 0.00398937f $X=9.27 $Y=0.8
+ $X2=0 $Y2=0
cc_800 N_A_1501_92#_M1023_g N_A_1339_74#_c_1305_n 3.11108e-19 $X=7.58 $Y=0.8
+ $X2=0 $Y2=0
cc_801 N_A_1501_92#_M1023_g N_A_1339_74#_c_1286_n 6.18383e-19 $X=7.58 $Y=0.8
+ $X2=0 $Y2=0
cc_802 N_A_1501_92#_M1031_g N_A_1339_74#_c_1296_n 0.0167055f $X=7.95 $Y=2.75
+ $X2=0 $Y2=0
cc_803 N_A_1501_92#_M1026_s N_A_1339_74#_c_1287_n 0.00594347f $X=9.035 $Y=1.84
+ $X2=0 $Y2=0
cc_804 N_A_1501_92#_c_1209_n N_A_1339_74#_c_1287_n 0.00784261f $X=9.105 $Y=0.925
+ $X2=0 $Y2=0
cc_805 N_A_1501_92#_c_1183_n N_A_1339_74#_c_1287_n 0.0152211f $X=9.74 $Y=2.375
+ $X2=0 $Y2=0
cc_806 N_A_1501_92#_c_1177_n N_A_1339_74#_c_1287_n 0.0107886f $X=9.74 $Y=1.095
+ $X2=0 $Y2=0
cc_807 N_A_1501_92#_c_1178_n N_A_1339_74#_c_1287_n 0.0600201f $X=9.825 $Y=2.29
+ $X2=0 $Y2=0
cc_808 N_A_1501_92#_c_1185_n N_A_1339_74#_c_1287_n 0.0417001f $X=9.18 $Y=2.375
+ $X2=0 $Y2=0
cc_809 N_A_1501_92#_c_1179_n N_A_1339_74#_c_1287_n 0.0286983f $X=9.27 $Y=0.8
+ $X2=0 $Y2=0
cc_810 N_A_1501_92#_M1031_g N_A_1339_74#_c_1298_n 5.1186e-19 $X=7.95 $Y=2.75
+ $X2=0 $Y2=0
cc_811 N_A_1501_92#_c_1185_n N_A_1339_74#_c_1298_n 0.00954913f $X=9.18 $Y=2.375
+ $X2=0 $Y2=0
cc_812 N_A_1501_92#_M1031_g N_A_1339_74#_c_1300_n 9.61445e-19 $X=7.95 $Y=2.75
+ $X2=0 $Y2=0
cc_813 N_A_1501_92#_M1031_g N_A_1339_74#_c_1302_n 0.0140867f $X=7.95 $Y=2.75
+ $X2=0 $Y2=0
cc_814 N_A_1501_92#_c_1175_n N_A_1339_74#_c_1302_n 0.0237116f $X=7.89 $Y=1.615
+ $X2=0 $Y2=0
cc_815 N_A_1501_92#_c_1176_n N_A_1339_74#_c_1302_n 8.67582e-19 $X=7.89 $Y=1.615
+ $X2=0 $Y2=0
cc_816 N_A_1501_92#_c_1177_n N_A_1339_74#_c_1288_n 0.00760222f $X=9.74 $Y=1.095
+ $X2=0 $Y2=0
cc_817 N_A_1501_92#_c_1178_n N_A_1339_74#_c_1288_n 0.00695766f $X=9.825 $Y=2.29
+ $X2=0 $Y2=0
cc_818 N_A_1501_92#_c_1183_n N_VPWR_M1026_d 0.00532511f $X=9.74 $Y=2.375 $X2=0
+ $Y2=0
cc_819 N_A_1501_92#_c_1178_n N_VPWR_M1026_d 0.00729559f $X=9.825 $Y=2.29 $X2=0
+ $Y2=0
cc_820 N_A_1501_92#_M1031_g N_VPWR_c_1603_n 0.00288539f $X=7.95 $Y=2.75 $X2=0
+ $Y2=0
cc_821 N_A_1501_92#_c_1183_n N_VPWR_c_1604_n 0.020837f $X=9.74 $Y=2.375 $X2=0
+ $Y2=0
cc_822 N_A_1501_92#_M1031_g N_VPWR_c_1609_n 0.0050156f $X=7.95 $Y=2.75 $X2=0
+ $Y2=0
cc_823 N_A_1501_92#_c_1185_n N_VPWR_c_1617_n 0.00541079f $X=9.18 $Y=2.375 $X2=0
+ $Y2=0
cc_824 N_A_1501_92#_M1031_g N_VPWR_c_1598_n 0.00540938f $X=7.95 $Y=2.75 $X2=0
+ $Y2=0
cc_825 N_A_1501_92#_c_1185_n N_VPWR_c_1598_n 0.00910369f $X=9.18 $Y=2.375 $X2=0
+ $Y2=0
cc_826 N_A_1501_92#_c_1177_n Q_N 0.00736666f $X=9.74 $Y=1.095 $X2=0 $Y2=0
cc_827 N_A_1501_92#_c_1178_n Q_N 0.0342329f $X=9.825 $Y=2.29 $X2=0 $Y2=0
cc_828 N_A_1501_92#_c_1178_n Q_N 0.00124832f $X=9.825 $Y=2.29 $X2=0 $Y2=0
cc_829 N_A_1501_92#_c_1209_n N_VGND_M1002_d 0.0237418f $X=9.105 $Y=0.925 $X2=0
+ $Y2=0
cc_830 N_A_1501_92#_c_1177_n N_VGND_M1013_s 0.00461825f $X=9.74 $Y=1.095 $X2=0
+ $Y2=0
cc_831 N_A_1501_92#_c_1177_n N_VGND_c_1813_n 0.0213705f $X=9.74 $Y=1.095 $X2=0
+ $Y2=0
cc_832 N_A_1501_92#_c_1179_n N_VGND_c_1813_n 0.0138209f $X=9.27 $Y=0.8 $X2=0
+ $Y2=0
cc_833 N_A_1501_92#_c_1179_n N_VGND_c_1822_n 0.00623106f $X=9.27 $Y=0.8 $X2=0
+ $Y2=0
cc_834 N_A_1501_92#_M1023_g N_VGND_c_1830_n 0.00311027f $X=7.58 $Y=0.8 $X2=0
+ $Y2=0
cc_835 N_A_1501_92#_c_1209_n N_VGND_c_1831_n 0.0586839f $X=9.105 $Y=0.925 $X2=0
+ $Y2=0
cc_836 N_A_1501_92#_M1023_g N_VGND_c_1834_n 0.00321167f $X=7.58 $Y=0.8 $X2=0
+ $Y2=0
cc_837 N_A_1501_92#_c_1209_n N_VGND_c_1834_n 0.0123962f $X=9.105 $Y=0.925 $X2=0
+ $Y2=0
cc_838 N_A_1501_92#_c_1193_n N_VGND_c_1834_n 0.0124246f $X=8.055 $Y=0.925 $X2=0
+ $Y2=0
cc_839 N_A_1501_92#_c_1179_n N_VGND_c_1834_n 0.00984494f $X=9.27 $Y=0.8 $X2=0
+ $Y2=0
cc_840 N_A_1501_92#_c_1193_n A_1531_118# 0.00412701f $X=8.055 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_841 N_A_1339_74#_M1015_g N_A_2221_74#_M1011_g 0.0227319f $X=11.475 $Y=2.34
+ $X2=0 $Y2=0
cc_842 N_A_1339_74#_M1007_g N_A_2221_74#_M1004_g 0.0226536f $X=11.465 $Y=0.69
+ $X2=0 $Y2=0
cc_843 N_A_1339_74#_M1024_g N_A_2221_74#_c_1462_n 0.00404932f $X=10.475 $Y=0.74
+ $X2=0 $Y2=0
cc_844 N_A_1339_74#_M1007_g N_A_2221_74#_c_1462_n 0.0189532f $X=11.465 $Y=0.69
+ $X2=0 $Y2=0
cc_845 N_A_1339_74#_M1030_g N_A_2221_74#_c_1463_n 0.00492925f $X=10.47 $Y=2.4
+ $X2=0 $Y2=0
cc_846 N_A_1339_74#_M1015_g N_A_2221_74#_c_1463_n 0.0212962f $X=11.475 $Y=2.34
+ $X2=0 $Y2=0
cc_847 N_A_1339_74#_M1007_g N_A_2221_74#_c_1464_n 0.00696112f $X=11.465 $Y=0.69
+ $X2=0 $Y2=0
cc_848 N_A_1339_74#_c_1285_n N_A_2221_74#_c_1464_n 0.0139657f $X=11.475 $Y=1.49
+ $X2=0 $Y2=0
cc_849 N_A_1339_74#_M1024_g N_A_2221_74#_c_1465_n 8.258e-19 $X=10.475 $Y=0.74
+ $X2=0 $Y2=0
cc_850 N_A_1339_74#_c_1281_n N_A_2221_74#_c_1465_n 0.0267893f $X=11.385 $Y=1.49
+ $X2=0 $Y2=0
cc_851 N_A_1339_74#_M1007_g N_A_2221_74#_c_1465_n 0.00110532f $X=11.465 $Y=0.69
+ $X2=0 $Y2=0
cc_852 N_A_1339_74#_c_1285_n N_A_2221_74#_c_1465_n 7.90981e-19 $X=11.475 $Y=1.49
+ $X2=0 $Y2=0
cc_853 N_A_1339_74#_M1007_g N_A_2221_74#_c_1466_n 0.00280567f $X=11.465 $Y=0.69
+ $X2=0 $Y2=0
cc_854 N_A_1339_74#_c_1285_n N_A_2221_74#_c_1466_n 0.0183328f $X=11.475 $Y=1.49
+ $X2=0 $Y2=0
cc_855 N_A_1339_74#_c_1296_n N_VPWR_c_1603_n 0.0141918f $X=8.46 $Y=2.215 $X2=0
+ $Y2=0
cc_856 N_A_1339_74#_c_1300_n N_VPWR_c_1603_n 0.00499852f $X=7.47 $Y=2.73 $X2=0
+ $Y2=0
cc_857 N_A_1339_74#_M1008_g N_VPWR_c_1604_n 0.0108651f $X=10.02 $Y=2.4 $X2=0
+ $Y2=0
cc_858 N_A_1339_74#_M1030_g N_VPWR_c_1604_n 4.59615e-19 $X=10.47 $Y=2.4 $X2=0
+ $Y2=0
cc_859 N_A_1339_74#_M1030_g N_VPWR_c_1605_n 0.0050513f $X=10.47 $Y=2.4 $X2=0
+ $Y2=0
cc_860 N_A_1339_74#_c_1281_n N_VPWR_c_1605_n 0.0089376f $X=11.385 $Y=1.49 $X2=0
+ $Y2=0
cc_861 N_A_1339_74#_M1015_g N_VPWR_c_1605_n 0.00456525f $X=11.475 $Y=2.34 $X2=0
+ $Y2=0
cc_862 N_A_1339_74#_M1015_g N_VPWR_c_1606_n 0.00869729f $X=11.475 $Y=2.34 $X2=0
+ $Y2=0
cc_863 N_A_1339_74#_c_1300_n N_VPWR_c_1609_n 0.0298117f $X=7.47 $Y=2.73 $X2=0
+ $Y2=0
cc_864 N_A_1339_74#_c_1301_n N_VPWR_c_1609_n 0.00624867f $X=7.75 $Y=2.3 $X2=0
+ $Y2=0
cc_865 N_A_1339_74#_M1008_g N_VPWR_c_1611_n 0.00460063f $X=10.02 $Y=2.4 $X2=0
+ $Y2=0
cc_866 N_A_1339_74#_M1030_g N_VPWR_c_1611_n 0.00493061f $X=10.47 $Y=2.4 $X2=0
+ $Y2=0
cc_867 N_A_1339_74#_c_1298_n N_VPWR_c_1617_n 0.0102883f $X=8.625 $Y=2.75 $X2=0
+ $Y2=0
cc_868 N_A_1339_74#_M1015_g N_VPWR_c_1618_n 0.00567889f $X=11.475 $Y=2.34 $X2=0
+ $Y2=0
cc_869 N_A_1339_74#_M1008_g N_VPWR_c_1598_n 0.00908554f $X=10.02 $Y=2.4 $X2=0
+ $Y2=0
cc_870 N_A_1339_74#_M1030_g N_VPWR_c_1598_n 0.00895963f $X=10.47 $Y=2.4 $X2=0
+ $Y2=0
cc_871 N_A_1339_74#_M1015_g N_VPWR_c_1598_n 0.00610055f $X=11.475 $Y=2.34 $X2=0
+ $Y2=0
cc_872 N_A_1339_74#_c_1296_n N_VPWR_c_1598_n 0.0126768f $X=8.46 $Y=2.215 $X2=0
+ $Y2=0
cc_873 N_A_1339_74#_c_1298_n N_VPWR_c_1598_n 0.0114715f $X=8.625 $Y=2.75 $X2=0
+ $Y2=0
cc_874 N_A_1339_74#_c_1300_n N_VPWR_c_1598_n 0.0249157f $X=7.47 $Y=2.73 $X2=0
+ $Y2=0
cc_875 N_A_1339_74#_c_1301_n N_VPWR_c_1598_n 0.0116485f $X=7.75 $Y=2.3 $X2=0
+ $Y2=0
cc_876 N_A_1339_74#_c_1301_n A_1524_508# 0.00131813f $X=7.75 $Y=2.3 $X2=-0.19
+ $Y2=-0.245
cc_877 N_A_1339_74#_c_1302_n A_1524_508# 0.00101982f $X=7.92 $Y=2.3 $X2=-0.19
+ $Y2=-0.245
cc_878 N_A_1339_74#_M1008_g Q_N 0.00163201f $X=10.02 $Y=2.4 $X2=0 $Y2=0
cc_879 N_A_1339_74#_M1013_g Q_N 0.00249434f $X=10.045 $Y=0.74 $X2=0 $Y2=0
cc_880 N_A_1339_74#_M1030_g Q_N 0.00625782f $X=10.47 $Y=2.4 $X2=0 $Y2=0
cc_881 N_A_1339_74#_M1024_g Q_N 0.0170389f $X=10.475 $Y=0.74 $X2=0 $Y2=0
cc_882 N_A_1339_74#_c_1282_n Q_N 0.0245493f $X=10.56 $Y=1.49 $X2=0 $Y2=0
cc_883 N_A_1339_74#_M1008_g Q_N 4.33031e-19 $X=10.02 $Y=2.4 $X2=0 $Y2=0
cc_884 N_A_1339_74#_M1030_g Q_N 0.002227f $X=10.47 $Y=2.4 $X2=0 $Y2=0
cc_885 N_A_1339_74#_M1030_g Q_N 0.0144554f $X=10.47 $Y=2.4 $X2=0 $Y2=0
cc_886 N_A_1339_74#_M1007_g Q 4.4789e-19 $X=11.465 $Y=0.69 $X2=0 $Y2=0
cc_887 N_A_1339_74#_M1003_g N_VGND_c_1813_n 0.00440494f $X=8.975 $Y=0.8 $X2=0
+ $Y2=0
cc_888 N_A_1339_74#_c_1276_n N_VGND_c_1813_n 6.71793e-19 $X=9.93 $Y=1.49 $X2=0
+ $Y2=0
cc_889 N_A_1339_74#_M1013_g N_VGND_c_1813_n 0.0136519f $X=10.045 $Y=0.74 $X2=0
+ $Y2=0
cc_890 N_A_1339_74#_M1024_g N_VGND_c_1813_n 5.19194e-19 $X=10.475 $Y=0.74 $X2=0
+ $Y2=0
cc_891 N_A_1339_74#_M1024_g N_VGND_c_1814_n 0.00510543f $X=10.475 $Y=0.74 $X2=0
+ $Y2=0
cc_892 N_A_1339_74#_c_1281_n N_VGND_c_1814_n 0.00890562f $X=11.385 $Y=1.49 $X2=0
+ $Y2=0
cc_893 N_A_1339_74#_M1007_g N_VGND_c_1814_n 0.00422013f $X=11.465 $Y=0.69 $X2=0
+ $Y2=0
cc_894 N_A_1339_74#_M1007_g N_VGND_c_1815_n 0.00744279f $X=11.465 $Y=0.69 $X2=0
+ $Y2=0
cc_895 N_A_1339_74#_M1013_g N_VGND_c_1818_n 0.00383152f $X=10.045 $Y=0.74 $X2=0
+ $Y2=0
cc_896 N_A_1339_74#_M1024_g N_VGND_c_1818_n 0.00422942f $X=10.475 $Y=0.74 $X2=0
+ $Y2=0
cc_897 N_A_1339_74#_M1003_g N_VGND_c_1822_n 0.00434252f $X=8.975 $Y=0.8 $X2=0
+ $Y2=0
cc_898 N_A_1339_74#_M1007_g N_VGND_c_1823_n 0.00434272f $X=11.465 $Y=0.69 $X2=0
+ $Y2=0
cc_899 N_A_1339_74#_M1003_g N_VGND_c_1831_n 0.00754579f $X=8.975 $Y=0.8 $X2=0
+ $Y2=0
cc_900 N_A_1339_74#_M1003_g N_VGND_c_1834_n 0.00479212f $X=8.975 $Y=0.8 $X2=0
+ $Y2=0
cc_901 N_A_1339_74#_M1013_g N_VGND_c_1834_n 0.0075754f $X=10.045 $Y=0.74 $X2=0
+ $Y2=0
cc_902 N_A_1339_74#_M1024_g N_VGND_c_1834_n 0.00788596f $X=10.475 $Y=0.74 $X2=0
+ $Y2=0
cc_903 N_A_1339_74#_M1007_g N_VGND_c_1834_n 0.00826311f $X=11.465 $Y=0.69 $X2=0
+ $Y2=0
cc_904 N_A_2221_74#_c_1463_n N_VPWR_c_1605_n 0.0698268f $X=11.25 $Y=1.985 $X2=0
+ $Y2=0
cc_905 N_A_2221_74#_M1011_g N_VPWR_c_1606_n 0.00542375f $X=12.005 $Y=2.4 $X2=0
+ $Y2=0
cc_906 N_A_2221_74#_c_1463_n N_VPWR_c_1606_n 0.0356152f $X=11.25 $Y=1.985 $X2=0
+ $Y2=0
cc_907 N_A_2221_74#_c_1464_n N_VPWR_c_1606_n 0.0199046f $X=11.94 $Y=1.465 $X2=0
+ $Y2=0
cc_908 N_A_2221_74#_c_1466_n N_VPWR_c_1606_n 0.00205259f $X=12.465 $Y=1.465
+ $X2=0 $Y2=0
cc_909 N_A_2221_74#_M1014_g N_VPWR_c_1608_n 0.00647357f $X=12.455 $Y=2.4 $X2=0
+ $Y2=0
cc_910 N_A_2221_74#_c_1463_n N_VPWR_c_1618_n 0.00975961f $X=11.25 $Y=1.985 $X2=0
+ $Y2=0
cc_911 N_A_2221_74#_M1011_g N_VPWR_c_1619_n 0.005209f $X=12.005 $Y=2.4 $X2=0
+ $Y2=0
cc_912 N_A_2221_74#_M1014_g N_VPWR_c_1619_n 0.0048691f $X=12.455 $Y=2.4 $X2=0
+ $Y2=0
cc_913 N_A_2221_74#_M1011_g N_VPWR_c_1598_n 0.00987399f $X=12.005 $Y=2.4 $X2=0
+ $Y2=0
cc_914 N_A_2221_74#_M1014_g N_VPWR_c_1598_n 0.00875947f $X=12.455 $Y=2.4 $X2=0
+ $Y2=0
cc_915 N_A_2221_74#_c_1463_n N_VPWR_c_1598_n 0.0111753f $X=11.25 $Y=1.985 $X2=0
+ $Y2=0
cc_916 N_A_2221_74#_c_1462_n Q_N 0.00476669f $X=11.25 $Y=0.515 $X2=0 $Y2=0
cc_917 N_A_2221_74#_c_1463_n Q_N 0.00530528f $X=11.25 $Y=1.985 $X2=0 $Y2=0
cc_918 N_A_2221_74#_c_1465_n Q_N 0.00865359f $X=11.25 $Y=1.465 $X2=0 $Y2=0
cc_919 N_A_2221_74#_M1011_g N_Q_c_1779_n 0.0128686f $X=12.005 $Y=2.4 $X2=0 $Y2=0
cc_920 N_A_2221_74#_M1014_g N_Q_c_1779_n 0.0149161f $X=12.455 $Y=2.4 $X2=0 $Y2=0
cc_921 N_A_2221_74#_M1011_g N_Q_c_1780_n 0.00319737f $X=12.005 $Y=2.4 $X2=0
+ $Y2=0
cc_922 N_A_2221_74#_M1014_g N_Q_c_1780_n 0.00270934f $X=12.455 $Y=2.4 $X2=0
+ $Y2=0
cc_923 N_A_2221_74#_c_1464_n N_Q_c_1780_n 0.00138666f $X=11.94 $Y=1.465 $X2=0
+ $Y2=0
cc_924 N_A_2221_74#_c_1466_n N_Q_c_1780_n 0.00310238f $X=12.465 $Y=1.465 $X2=0
+ $Y2=0
cc_925 N_A_2221_74#_M1011_g N_Q_c_1776_n 0.00293165f $X=12.005 $Y=2.4 $X2=0
+ $Y2=0
cc_926 N_A_2221_74#_M1004_g N_Q_c_1776_n 0.0025553f $X=12.035 $Y=0.74 $X2=0
+ $Y2=0
cc_927 N_A_2221_74#_M1014_g N_Q_c_1776_n 0.00994275f $X=12.455 $Y=2.4 $X2=0
+ $Y2=0
cc_928 N_A_2221_74#_M1016_g N_Q_c_1776_n 0.00866774f $X=12.465 $Y=0.74 $X2=0
+ $Y2=0
cc_929 N_A_2221_74#_c_1464_n N_Q_c_1776_n 0.0249855f $X=11.94 $Y=1.465 $X2=0
+ $Y2=0
cc_930 N_A_2221_74#_c_1466_n N_Q_c_1776_n 0.0237264f $X=12.465 $Y=1.465 $X2=0
+ $Y2=0
cc_931 N_A_2221_74#_M1004_g Q 0.00746865f $X=12.035 $Y=0.74 $X2=0 $Y2=0
cc_932 N_A_2221_74#_M1016_g Q 0.0081896f $X=12.465 $Y=0.74 $X2=0 $Y2=0
cc_933 N_A_2221_74#_M1004_g Q 0.00423302f $X=12.035 $Y=0.74 $X2=0 $Y2=0
cc_934 N_A_2221_74#_M1016_g Q 0.00215589f $X=12.465 $Y=0.74 $X2=0 $Y2=0
cc_935 N_A_2221_74#_c_1462_n Q 0.00238899f $X=11.25 $Y=0.515 $X2=0 $Y2=0
cc_936 N_A_2221_74#_c_1466_n Q 0.00244427f $X=12.465 $Y=1.465 $X2=0 $Y2=0
cc_937 N_A_2221_74#_c_1462_n N_VGND_c_1814_n 0.051504f $X=11.25 $Y=0.515 $X2=0
+ $Y2=0
cc_938 N_A_2221_74#_M1004_g N_VGND_c_1815_n 0.00737997f $X=12.035 $Y=0.74 $X2=0
+ $Y2=0
cc_939 N_A_2221_74#_c_1462_n N_VGND_c_1815_n 0.0270962f $X=11.25 $Y=0.515 $X2=0
+ $Y2=0
cc_940 N_A_2221_74#_c_1464_n N_VGND_c_1815_n 0.019673f $X=11.94 $Y=1.465 $X2=0
+ $Y2=0
cc_941 N_A_2221_74#_c_1466_n N_VGND_c_1815_n 0.00301993f $X=12.465 $Y=1.465
+ $X2=0 $Y2=0
cc_942 N_A_2221_74#_M1016_g N_VGND_c_1817_n 0.00646793f $X=12.465 $Y=0.74 $X2=0
+ $Y2=0
cc_943 N_A_2221_74#_c_1462_n N_VGND_c_1823_n 0.0145639f $X=11.25 $Y=0.515 $X2=0
+ $Y2=0
cc_944 N_A_2221_74#_M1004_g N_VGND_c_1824_n 0.00434272f $X=12.035 $Y=0.74 $X2=0
+ $Y2=0
cc_945 N_A_2221_74#_M1016_g N_VGND_c_1824_n 0.00422942f $X=12.465 $Y=0.74 $X2=0
+ $Y2=0
cc_946 N_A_2221_74#_M1004_g N_VGND_c_1834_n 0.00821312f $X=12.035 $Y=0.74 $X2=0
+ $Y2=0
cc_947 N_A_2221_74#_M1016_g N_VGND_c_1834_n 0.00787255f $X=12.465 $Y=0.74 $X2=0
+ $Y2=0
cc_948 N_A_2221_74#_c_1462_n N_VGND_c_1834_n 0.0119984f $X=11.25 $Y=0.515 $X2=0
+ $Y2=0
cc_949 N_A_27_74#_c_1537_n N_VPWR_M1018_d 9.71305e-19 $X=2.445 $Y=2.145 $X2=0
+ $Y2=0
cc_950 N_A_27_74#_c_1581_n N_VPWR_M1018_d 0.00499461f $X=1.71 $Y=2.145 $X2=0
+ $Y2=0
cc_951 N_A_27_74#_c_1535_n N_VPWR_c_1599_n 0.0158217f $X=0.28 $Y=2.75 $X2=0
+ $Y2=0
cc_952 N_A_27_74#_c_1536_n N_VPWR_c_1599_n 0.0274627f $X=1.625 $Y=2.275 $X2=0
+ $Y2=0
cc_953 N_A_27_74#_c_1536_n N_VPWR_c_1600_n 0.00220908f $X=1.625 $Y=2.275 $X2=0
+ $Y2=0
cc_954 N_A_27_74#_c_1537_n N_VPWR_c_1600_n 0.00262985f $X=2.445 $Y=2.145 $X2=0
+ $Y2=0
cc_955 N_A_27_74#_c_1581_n N_VPWR_c_1600_n 0.0112212f $X=1.71 $Y=2.145 $X2=0
+ $Y2=0
cc_956 N_A_27_74#_c_1535_n N_VPWR_c_1613_n 0.011066f $X=0.28 $Y=2.75 $X2=0 $Y2=0
cc_957 N_A_27_74#_c_1535_n N_VPWR_c_1598_n 0.00915947f $X=0.28 $Y=2.75 $X2=0
+ $Y2=0
cc_958 N_A_27_74#_c_1529_n N_VGND_c_1809_n 0.0172562f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_959 N_A_27_74#_c_1529_n N_VGND_c_1820_n 0.0109681f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_960 N_A_27_74#_c_1529_n N_VGND_c_1834_n 0.00912188f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_961 N_VPWR_c_1605_n Q_N 0.0437165f $X=10.695 $Y=1.985 $X2=0 $Y2=0
cc_962 N_VPWR_c_1604_n Q_N 0.0131276f $X=9.795 $Y=2.805 $X2=0 $Y2=0
cc_963 N_VPWR_c_1611_n Q_N 0.0128394f $X=10.605 $Y=3.33 $X2=0 $Y2=0
cc_964 N_VPWR_c_1598_n Q_N 0.0108616f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_965 N_VPWR_c_1619_n N_Q_c_1779_n 0.0157112f $X=12.595 $Y=3.33 $X2=0 $Y2=0
cc_966 N_VPWR_c_1598_n N_Q_c_1779_n 0.0127977f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_967 N_VPWR_c_1606_n N_Q_c_1780_n 0.0400476f $X=11.78 $Y=1.985 $X2=0 $Y2=0
cc_968 N_VPWR_c_1608_n N_Q_c_1780_n 0.0455874f $X=12.68 $Y=1.985 $X2=0 $Y2=0
cc_969 Q_N N_VGND_c_1813_n 0.0182946f $X=10.235 $Y=0.47 $X2=0 $Y2=0
cc_970 Q_N N_VGND_c_1814_n 0.0297335f $X=10.235 $Y=0.47 $X2=0 $Y2=0
cc_971 Q_N N_VGND_c_1818_n 0.0114106f $X=10.235 $Y=0.47 $X2=0 $Y2=0
cc_972 Q_N N_VGND_c_1834_n 0.00936481f $X=10.235 $Y=0.47 $X2=0 $Y2=0
cc_973 Q N_VGND_c_1815_n 0.0263849f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_974 Q N_VGND_c_1817_n 0.0308798f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_975 Q N_VGND_c_1824_n 0.0149085f $X=12.155 $Y=0.47 $X2=0 $Y2=0
cc_976 Q N_VGND_c_1834_n 0.0122037f $X=12.155 $Y=0.47 $X2=0 $Y2=0

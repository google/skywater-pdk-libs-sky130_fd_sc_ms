* File: sky130_fd_sc_ms__xnor3_1.pxi.spice
* Created: Fri Aug 28 18:18:00 2020
* 
x_PM_SKY130_FD_SC_MS__XNOR3_1%A_81_268# N_A_81_268#_M1008_d N_A_81_268#_M1000_d
+ N_A_81_268#_M1016_g N_A_81_268#_M1003_g N_A_81_268#_c_177_n
+ N_A_81_268#_c_168_n N_A_81_268#_c_254_p N_A_81_268#_c_186_p
+ N_A_81_268#_c_225_p N_A_81_268#_c_178_n N_A_81_268#_c_179_n
+ N_A_81_268#_c_180_n N_A_81_268#_c_169_n N_A_81_268#_c_170_n
+ N_A_81_268#_c_171_n N_A_81_268#_c_208_p N_A_81_268#_c_172_n
+ N_A_81_268#_c_173_n N_A_81_268#_c_174_n N_A_81_268#_c_183_n
+ N_A_81_268#_c_175_n PM_SKY130_FD_SC_MS__XNOR3_1%A_81_268#
x_PM_SKY130_FD_SC_MS__XNOR3_1%C N_C_M1013_g N_C_M1018_g N_C_c_270_n N_C_c_271_n
+ N_C_M1000_g N_C_c_273_n N_C_M1008_g C N_C_c_274_n N_C_c_275_n N_C_c_276_n
+ PM_SKY130_FD_SC_MS__XNOR3_1%C
x_PM_SKY130_FD_SC_MS__XNOR3_1%A_232_162# N_A_232_162#_M1013_d
+ N_A_232_162#_M1018_d N_A_232_162#_M1006_g N_A_232_162#_M1019_g
+ N_A_232_162#_c_352_n N_A_232_162#_c_359_n N_A_232_162#_c_353_n
+ N_A_232_162#_c_360_n N_A_232_162#_c_354_n N_A_232_162#_c_355_n
+ N_A_232_162#_c_356_n N_A_232_162#_c_357_n
+ PM_SKY130_FD_SC_MS__XNOR3_1%A_232_162#
x_PM_SKY130_FD_SC_MS__XNOR3_1%A_786_100# N_A_786_100#_M1001_d
+ N_A_786_100#_M1002_d N_A_786_100#_M1009_g N_A_786_100#_M1007_g
+ N_A_786_100#_c_441_n N_A_786_100#_c_442_n N_A_786_100#_M1012_g
+ N_A_786_100#_M1021_g N_A_786_100#_c_445_n N_A_786_100#_c_446_n
+ N_A_786_100#_c_452_n N_A_786_100#_c_447_n N_A_786_100#_c_453_n
+ N_A_786_100#_c_448_n N_A_786_100#_c_449_n
+ PM_SKY130_FD_SC_MS__XNOR3_1%A_786_100#
x_PM_SKY130_FD_SC_MS__XNOR3_1%B N_B_M1002_g N_B_c_561_n N_B_M1001_g N_B_c_568_n
+ N_B_c_569_n N_B_c_570_n N_B_M1010_g N_B_M1004_g N_B_c_573_n N_B_c_574_n
+ N_B_M1015_g N_B_M1014_g N_B_c_564_n N_B_c_565_n N_B_c_579_n N_B_c_580_n B
+ N_B_c_566_n PM_SKY130_FD_SC_MS__XNOR3_1%B
x_PM_SKY130_FD_SC_MS__XNOR3_1%A N_A_M1017_g N_A_M1020_g A N_A_c_691_n
+ PM_SKY130_FD_SC_MS__XNOR3_1%A
x_PM_SKY130_FD_SC_MS__XNOR3_1%A_897_54# N_A_897_54#_M1007_s N_A_897_54#_M1014_d
+ N_A_897_54#_M1009_s N_A_897_54#_M1015_d N_A_897_54#_M1011_g
+ N_A_897_54#_M1005_g N_A_897_54#_c_742_n N_A_897_54#_c_734_n
+ N_A_897_54#_c_735_n N_A_897_54#_c_767_n N_A_897_54#_c_743_n
+ N_A_897_54#_c_736_n N_A_897_54#_c_737_n N_A_897_54#_c_788_n
+ N_A_897_54#_c_744_n N_A_897_54#_c_738_n N_A_897_54#_c_745_n
+ N_A_897_54#_c_791_n N_A_897_54#_c_739_n N_A_897_54#_c_740_n
+ PM_SKY130_FD_SC_MS__XNOR3_1%A_897_54#
x_PM_SKY130_FD_SC_MS__XNOR3_1%X N_X_M1003_s N_X_M1016_s N_X_c_861_n N_X_c_862_n
+ N_X_c_858_n X X X PM_SKY130_FD_SC_MS__XNOR3_1%X
x_PM_SKY130_FD_SC_MS__XNOR3_1%VPWR N_VPWR_M1016_d N_VPWR_M1002_s N_VPWR_M1020_d
+ N_VPWR_c_880_n N_VPWR_c_881_n N_VPWR_c_882_n VPWR N_VPWR_c_883_n
+ N_VPWR_c_884_n N_VPWR_c_885_n N_VPWR_c_886_n N_VPWR_c_879_n N_VPWR_c_888_n
+ N_VPWR_c_889_n N_VPWR_c_890_n PM_SKY130_FD_SC_MS__XNOR3_1%VPWR
x_PM_SKY130_FD_SC_MS__XNOR3_1%A_363_394# N_A_363_394#_M1006_d
+ N_A_363_394#_M1021_d N_A_363_394#_M1000_s N_A_363_394#_M1009_d
+ N_A_363_394#_c_961_n N_A_363_394#_c_962_n N_A_363_394#_c_970_n
+ N_A_363_394#_c_955_n N_A_363_394#_c_956_n N_A_363_394#_c_964_n
+ N_A_363_394#_c_965_n N_A_363_394#_c_957_n N_A_363_394#_c_958_n
+ N_A_363_394#_c_966_n N_A_363_394#_c_959_n N_A_363_394#_c_960_n
+ PM_SKY130_FD_SC_MS__XNOR3_1%A_363_394#
x_PM_SKY130_FD_SC_MS__XNOR3_1%A_371_74# N_A_371_74#_M1008_s N_A_371_74#_M1007_d
+ N_A_371_74#_M1019_d N_A_371_74#_M1012_d N_A_371_74#_c_1086_n
+ N_A_371_74#_c_1087_n N_A_371_74#_c_1088_n N_A_371_74#_c_1134_n
+ N_A_371_74#_c_1089_n N_A_371_74#_c_1090_n N_A_371_74#_c_1097_n
+ N_A_371_74#_c_1148_n N_A_371_74#_c_1166_n N_A_371_74#_c_1098_n
+ N_A_371_74#_c_1091_n N_A_371_74#_c_1092_n N_A_371_74#_c_1093_n
+ N_A_371_74#_c_1094_n PM_SKY130_FD_SC_MS__XNOR3_1%A_371_74#
x_PM_SKY130_FD_SC_MS__XNOR3_1%A_1116_383# N_A_1116_383#_M1004_d
+ N_A_1116_383#_M1005_d N_A_1116_383#_M1010_d N_A_1116_383#_M1011_d
+ N_A_1116_383#_c_1227_n N_A_1116_383#_c_1221_n N_A_1116_383#_c_1222_n
+ N_A_1116_383#_c_1212_n N_A_1116_383#_c_1213_n N_A_1116_383#_c_1214_n
+ N_A_1116_383#_c_1224_n N_A_1116_383#_c_1225_n N_A_1116_383#_c_1215_n
+ N_A_1116_383#_c_1216_n N_A_1116_383#_c_1217_n N_A_1116_383#_c_1237_n
+ N_A_1116_383#_c_1218_n N_A_1116_383#_c_1219_n N_A_1116_383#_c_1220_n
+ PM_SKY130_FD_SC_MS__XNOR3_1%A_1116_383#
x_PM_SKY130_FD_SC_MS__XNOR3_1%VGND N_VGND_M1003_d N_VGND_M1001_s N_VGND_M1017_d
+ N_VGND_c_1327_n N_VGND_c_1328_n N_VGND_c_1329_n VGND N_VGND_c_1330_n
+ N_VGND_c_1331_n N_VGND_c_1332_n N_VGND_c_1333_n N_VGND_c_1334_n
+ N_VGND_c_1335_n N_VGND_c_1336_n N_VGND_c_1337_n
+ PM_SKY130_FD_SC_MS__XNOR3_1%VGND
cc_1 VNB N_A_81_268#_c_168_n 0.0113669f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=0.745
cc_2 VNB N_A_81_268#_c_169_n 0.0104919f $X=-0.19 $Y=-0.245 $X2=1.58 $Y2=0.66
cc_3 VNB N_A_81_268#_c_170_n 0.0135346f $X=-0.19 $Y=-0.245 $X2=2.335 $Y2=0.34
cc_4 VNB N_A_81_268#_c_171_n 0.00494049f $X=-0.19 $Y=-0.245 $X2=1.665 $Y2=0.34
cc_5 VNB N_A_81_268#_c_172_n 0.00384286f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.505
cc_6 VNB N_A_81_268#_c_173_n 0.0289515f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.505
cc_7 VNB N_A_81_268#_c_174_n 0.00189669f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.34
cc_8 VNB N_A_81_268#_c_175_n 0.0209671f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.34
cc_9 VNB N_C_c_270_n 0.0526962f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_10 VNB N_C_c_271_n 0.0309647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_C_M1000_g 0.00409515f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.86
cc_12 VNB N_C_c_273_n 0.0180813f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.83
cc_13 VNB N_C_c_274_n 0.0228235f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.035
cc_14 VNB N_C_c_275_n 0.0201289f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=2.035
cc_15 VNB N_C_c_276_n 9.1398e-19 $X=-0.19 $Y=-0.245 $X2=2.325 $Y2=2.99
cc_16 VNB N_A_232_162#_M1006_g 0.0429487f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_17 VNB N_A_232_162#_c_352_n 0.00323147f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.34
cc_18 VNB N_A_232_162#_c_353_n 0.00384589f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=2.905
cc_19 VNB N_A_232_162#_c_354_n 4.91183e-19 $X=-0.19 $Y=-0.245 $X2=1.665 $Y2=0.34
cc_20 VNB N_A_232_162#_c_355_n 0.00109233f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=0.545
cc_21 VNB N_A_232_162#_c_356_n 0.0187643f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=0.545
cc_22 VNB N_A_232_162#_c_357_n 0.00523187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_786_100#_M1007_g 0.0337529f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.83
cc_24 VNB N_A_786_100#_c_441_n 0.0811869f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.34
cc_25 VNB N_A_786_100#_c_442_n 0.0127779f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.67
cc_26 VNB N_A_786_100#_M1012_g 0.0103348f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=0.745
cc_27 VNB N_A_786_100#_M1021_g 0.0393244f $X=-0.19 $Y=-0.245 $X2=2.325 $Y2=2.99
cc_28 VNB N_A_786_100#_c_445_n 0.0183891f $X=-0.19 $Y=-0.245 $X2=1.58 $Y2=0.66
cc_29 VNB N_A_786_100#_c_446_n 0.00541476f $X=-0.19 $Y=-0.245 $X2=1.665 $Y2=0.34
cc_30 VNB N_A_786_100#_c_447_n 0.00232667f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.67
cc_31 VNB N_A_786_100#_c_448_n 0.00450057f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.505
cc_32 VNB N_A_786_100#_c_449_n 0.026185f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.34
cc_33 VNB N_B_c_561_n 0.0219042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_B_M1004_g 0.031515f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=0.745
cc_35 VNB N_B_M1014_g 0.0326237f $X=-0.19 $Y=-0.245 $X2=2.335 $Y2=0.34
cc_36 VNB N_B_c_564_n 0.0190224f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=0.545
cc_37 VNB N_B_c_565_n 0.0366081f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=0.545
cc_38 VNB N_B_c_566_n 0.00210104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_M1017_g 0.0213947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB A 0.00339401f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_41 VNB N_A_c_691_n 0.0174305f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.86
cc_42 VNB N_A_897_54#_M1005_g 0.025997f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=0.745
cc_43 VNB N_A_897_54#_c_734_n 0.0261652f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=2.905
cc_44 VNB N_A_897_54#_c_735_n 0.00314505f $X=-0.19 $Y=-0.245 $X2=2.335 $Y2=0.34
cc_45 VNB N_A_897_54#_c_736_n 0.00282973f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=0.545
cc_46 VNB N_A_897_54#_c_737_n 0.00245736f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=0.545
cc_47 VNB N_A_897_54#_c_738_n 0.0106808f $X=-0.19 $Y=-0.245 $X2=2.49 $Y2=2.99
cc_48 VNB N_A_897_54#_c_739_n 0.0227391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_897_54#_c_740_n 0.00201658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_X_c_858_n 0.0221881f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.34
cc_51 VNB X 0.0251976f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.67
cc_52 VNB X 0.00710642f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.95
cc_53 VNB N_VPWR_c_879_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_363_394#_c_955_n 0.0119754f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.035
cc_55 VNB N_A_363_394#_c_956_n 0.0161108f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=2.12
cc_56 VNB N_A_363_394#_c_957_n 0.00931374f $X=-0.19 $Y=-0.245 $X2=1.665 $Y2=0.34
cc_57 VNB N_A_363_394#_c_958_n 5.75182e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_363_394#_c_959_n 0.00700879f $X=-0.19 $Y=-0.245 $X2=2.49 $Y2=2.795
cc_59 VNB N_A_363_394#_c_960_n 9.95883e-19 $X=-0.19 $Y=-0.245 $X2=2.49 $Y2=2.795
cc_60 VNB N_A_371_74#_c_1086_n 0.00659688f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.34
cc_61 VNB N_A_371_74#_c_1087_n 0.0154078f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.95
cc_62 VNB N_A_371_74#_c_1088_n 0.00727053f $X=-0.19 $Y=-0.245 $X2=0.975
+ $Y2=2.035
cc_63 VNB N_A_371_74#_c_1089_n 0.00440829f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=2.99
cc_64 VNB N_A_371_74#_c_1090_n 0.00226213f $X=-0.19 $Y=-0.245 $X2=1.58 $Y2=0.425
cc_65 VNB N_A_371_74#_c_1091_n 0.0288161f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.34
cc_66 VNB N_A_371_74#_c_1092_n 0.00112558f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.67
cc_67 VNB N_A_371_74#_c_1093_n 0.00254106f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.505
cc_68 VNB N_A_371_74#_c_1094_n 0.00313006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1116_383#_c_1212_n 0.0102941f $X=-0.19 $Y=-0.245 $X2=0.785
+ $Y2=0.745
cc_70 VNB N_A_1116_383#_c_1213_n 0.00220528f $X=-0.19 $Y=-0.245 $X2=0.975
+ $Y2=2.035
cc_71 VNB N_A_1116_383#_c_1214_n 7.41744e-19 $X=-0.19 $Y=-0.245 $X2=1.06
+ $Y2=2.12
cc_72 VNB N_A_1116_383#_c_1215_n 0.0240083f $X=-0.19 $Y=-0.245 $X2=1.665
+ $Y2=0.34
cc_73 VNB N_A_1116_383#_c_1216_n 0.00596711f $X=-0.19 $Y=-0.245 $X2=0.59
+ $Y2=1.505
cc_74 VNB N_A_1116_383#_c_1217_n 0.0117474f $X=-0.19 $Y=-0.245 $X2=0.59
+ $Y2=1.505
cc_75 VNB N_A_1116_383#_c_1218_n 0.00259632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1116_383#_c_1219_n 0.0200335f $X=-0.19 $Y=-0.245 $X2=0.58
+ $Y2=1.505
cc_77 VNB N_A_1116_383#_c_1220_n 8.74794e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1327_n 0.015181f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.86
cc_79 VNB N_VGND_c_1328_n 0.0147615f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.67
cc_80 VNB N_VGND_c_1329_n 0.0214927f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.035
cc_81 VNB N_VGND_c_1330_n 0.0196503f $X=-0.19 $Y=-0.245 $X2=2.325 $Y2=2.99
cc_82 VNB N_VGND_c_1331_n 0.0605039f $X=-0.19 $Y=-0.245 $X2=1.665 $Y2=0.34
cc_83 VNB N_VGND_c_1332_n 0.0829908f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.34
cc_84 VNB N_VGND_c_1333_n 0.0181195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1334_n 0.445941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1335_n 0.00631593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1336_n 0.00631651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1337_n 0.00788625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VPB N_A_81_268#_M1016_g 0.0290559f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_90 VPB N_A_81_268#_c_177_n 0.00263861f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.95
cc_91 VPB N_A_81_268#_c_178_n 0.0136763f $X=-0.19 $Y=1.66 $X2=1.06 $Y2=2.905
cc_92 VPB N_A_81_268#_c_179_n 0.0310815f $X=-0.19 $Y=1.66 $X2=2.325 $Y2=2.99
cc_93 VPB N_A_81_268#_c_180_n 0.00348146f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=2.99
cc_94 VPB N_A_81_268#_c_172_n 5.57459e-19 $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.505
cc_95 VPB N_A_81_268#_c_173_n 0.00555941f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.505
cc_96 VPB N_A_81_268#_c_183_n 0.0111754f $X=-0.19 $Y=1.66 $X2=2.49 $Y2=2.795
cc_97 VPB N_C_M1018_g 0.0248718f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_C_M1000_g 0.0365283f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.86
cc_99 VPB N_C_c_274_n 0.00582698f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=2.035
cc_100 VPB N_C_c_276_n 0.00453434f $X=-0.19 $Y=1.66 $X2=2.325 $Y2=2.99
cc_101 VPB N_A_232_162#_M1019_g 0.0249402f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.86
cc_102 VPB N_A_232_162#_c_359_n 0.0111292f $X=-0.19 $Y=1.66 $X2=0.785 $Y2=0.745
cc_103 VPB N_A_232_162#_c_360_n 0.00417031f $X=-0.19 $Y=1.66 $X2=2.335 $Y2=0.34
cc_104 VPB N_A_232_162#_c_354_n 9.82239e-19 $X=-0.19 $Y=1.66 $X2=1.665 $Y2=0.34
cc_105 VPB N_A_232_162#_c_355_n 6.47771e-19 $X=-0.19 $Y=1.66 $X2=2.5 $Y2=0.545
cc_106 VPB N_A_232_162#_c_356_n 0.0171909f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=0.545
cc_107 VPB N_A_232_162#_c_357_n 0.013886f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_786_100#_M1009_g 0.023037f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_109 VPB N_A_786_100#_M1012_g 0.023759f $X=-0.19 $Y=1.66 $X2=0.785 $Y2=0.745
cc_110 VPB N_A_786_100#_c_452_n 0.00338753f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_786_100#_c_453_n 0.00345271f $X=-0.19 $Y=1.66 $X2=2.49 $Y2=2.795
cc_112 VPB N_A_786_100#_c_448_n 8.48419e-19 $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.505
cc_113 VPB N_A_786_100#_c_449_n 0.00678153f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.34
cc_114 VPB N_B_M1002_g 0.0240607f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_B_c_568_n 0.0778069f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_116 VPB N_B_c_569_n 0.0652201f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_B_c_570_n 0.012363f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.34
cc_118 VPB N_B_M1010_g 0.0430692f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.34
cc_119 VPB N_B_M1004_g 0.00149491f $X=-0.19 $Y=1.66 $X2=1.495 $Y2=0.745
cc_120 VPB N_B_c_573_n 0.0745877f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=2.035
cc_121 VPB N_B_c_574_n 0.00587777f $X=-0.19 $Y=1.66 $X2=1.06 $Y2=2.12
cc_122 VPB N_B_M1015_g 0.0325588f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=2.99
cc_123 VPB N_B_M1014_g 0.00150828f $X=-0.19 $Y=1.66 $X2=2.335 $Y2=0.34
cc_124 VPB N_B_c_564_n 0.00287621f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=0.545
cc_125 VPB N_B_c_565_n 0.00615023f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=0.545
cc_126 VPB N_B_c_579_n 0.0112504f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.505
cc_127 VPB N_B_c_580_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.505
cc_128 VPB N_B_c_566_n 0.00520205f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_M1020_g 0.0220202f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.67
cc_130 VPB A 0.0032939f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_131 VPB N_A_c_691_n 0.00954793f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.86
cc_132 VPB N_A_897_54#_M1011_g 0.0242992f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.34
cc_133 VPB N_A_897_54#_c_742_n 0.0370795f $X=-0.19 $Y=1.66 $X2=0.785 $Y2=2.035
cc_134 VPB N_A_897_54#_c_743_n 0.00148809f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=0.425
cc_135 VPB N_A_897_54#_c_744_n 0.00152579f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.67
cc_136 VPB N_A_897_54#_c_745_n 0.00892558f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.505
cc_137 VPB N_A_897_54#_c_739_n 0.0114884f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_X_c_861_n 0.00656497f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_139 VPB N_X_c_862_n 0.0409054f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.34
cc_140 VPB N_X_c_858_n 0.00857113f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.34
cc_141 VPB N_VPWR_c_880_n 0.00585142f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.86
cc_142 VPB N_VPWR_c_881_n 0.0173465f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.67
cc_143 VPB N_VPWR_c_882_n 0.0082002f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=2.035
cc_144 VPB N_VPWR_c_883_n 0.0175529f $X=-0.19 $Y=1.66 $X2=2.325 $Y2=2.99
cc_145 VPB N_VPWR_c_884_n 0.0665747f $X=-0.19 $Y=1.66 $X2=1.665 $Y2=0.34
cc_146 VPB N_VPWR_c_885_n 0.0876859f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.34
cc_147 VPB N_VPWR_c_886_n 0.0182776f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_879_n 0.0987141f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_888_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_889_n 0.00632279f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_890_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_363_394#_c_961_n 0.00179965f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.34
cc_153 VPB N_A_363_394#_c_962_n 0.0105867f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.95
cc_154 VPB N_A_363_394#_c_955_n 0.00977296f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=2.035
cc_155 VPB N_A_363_394#_c_964_n 0.00362121f $X=-0.19 $Y=1.66 $X2=1.06 $Y2=2.905
cc_156 VPB N_A_363_394#_c_965_n 0.00337867f $X=-0.19 $Y=1.66 $X2=1.58 $Y2=0.66
cc_157 VPB N_A_363_394#_c_966_n 0.00147614f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.67
cc_158 VPB N_A_371_74#_c_1088_n 0.00696615f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=2.035
cc_159 VPB N_A_371_74#_c_1090_n 2.87575e-19 $X=-0.19 $Y=1.66 $X2=1.58 $Y2=0.425
cc_160 VPB N_A_371_74#_c_1097_n 0.00782132f $X=-0.19 $Y=1.66 $X2=1.58 $Y2=0.66
cc_161 VPB N_A_371_74#_c_1098_n 0.00179963f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.505
cc_162 VPB N_A_1116_383#_c_1221_n 0.00375705f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.95
cc_163 VPB N_A_1116_383#_c_1222_n 0.00198282f $X=-0.19 $Y=1.66 $X2=1.495
+ $Y2=0.745
cc_164 VPB N_A_1116_383#_c_1214_n 0.002223f $X=-0.19 $Y=1.66 $X2=1.06 $Y2=2.12
cc_165 VPB N_A_1116_383#_c_1224_n 0.00545527f $X=-0.19 $Y=1.66 $X2=1.06
+ $Y2=2.905
cc_166 VPB N_A_1116_383#_c_1225_n 0.0257916f $X=-0.19 $Y=1.66 $X2=1.145 $Y2=2.99
cc_167 VPB N_A_1116_383#_c_1219_n 0.0231953f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.505
cc_168 N_A_81_268#_M1016_g N_C_M1018_g 0.0132293f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_169 N_A_81_268#_c_177_n N_C_M1018_g 0.00362599f $X=0.7 $Y=1.95 $X2=0 $Y2=0
cc_170 N_A_81_268#_c_186_p N_C_M1018_g 0.00607771f $X=0.975 $Y=2.035 $X2=0 $Y2=0
cc_171 N_A_81_268#_c_178_n N_C_M1018_g 0.0165132f $X=1.06 $Y=2.905 $X2=0 $Y2=0
cc_172 N_A_81_268#_c_179_n N_C_M1018_g 0.00434263f $X=2.325 $Y=2.99 $X2=0 $Y2=0
cc_173 N_A_81_268#_c_168_n N_C_c_270_n 6.31839e-19 $X=1.495 $Y=0.745 $X2=0 $Y2=0
cc_174 N_A_81_268#_c_179_n N_C_M1000_g 0.00824549f $X=2.325 $Y=2.99 $X2=0 $Y2=0
cc_175 N_A_81_268#_c_183_n N_C_M1000_g 0.00352829f $X=2.49 $Y=2.795 $X2=0 $Y2=0
cc_176 N_A_81_268#_c_169_n N_C_c_273_n 0.00292421f $X=1.58 $Y=0.66 $X2=0 $Y2=0
cc_177 N_A_81_268#_c_170_n N_C_c_273_n 0.0153137f $X=2.335 $Y=0.34 $X2=0 $Y2=0
cc_178 N_A_81_268#_M1016_g N_C_c_274_n 2.09353e-19 $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_179 N_A_81_268#_c_186_p N_C_c_274_n 3.99897e-19 $X=0.975 $Y=2.035 $X2=0 $Y2=0
cc_180 N_A_81_268#_c_172_n N_C_c_274_n 0.00213403f $X=0.59 $Y=1.505 $X2=0 $Y2=0
cc_181 N_A_81_268#_c_173_n N_C_c_274_n 0.0174684f $X=0.59 $Y=1.505 $X2=0 $Y2=0
cc_182 N_A_81_268#_c_168_n N_C_c_275_n 0.0133267f $X=1.495 $Y=0.745 $X2=0 $Y2=0
cc_183 N_A_81_268#_c_173_n N_C_c_275_n 4.44706e-19 $X=0.59 $Y=1.505 $X2=0 $Y2=0
cc_184 N_A_81_268#_c_174_n N_C_c_275_n 0.00868243f $X=0.605 $Y=1.34 $X2=0 $Y2=0
cc_185 N_A_81_268#_c_175_n N_C_c_275_n 0.012441f $X=0.58 $Y=1.34 $X2=0 $Y2=0
cc_186 N_A_81_268#_c_168_n N_C_c_276_n 0.00388368f $X=1.495 $Y=0.745 $X2=0 $Y2=0
cc_187 N_A_81_268#_c_186_p N_C_c_276_n 0.0102424f $X=0.975 $Y=2.035 $X2=0 $Y2=0
cc_188 N_A_81_268#_c_172_n N_C_c_276_n 0.0292202f $X=0.59 $Y=1.505 $X2=0 $Y2=0
cc_189 N_A_81_268#_c_173_n N_C_c_276_n 3.86162e-19 $X=0.59 $Y=1.505 $X2=0 $Y2=0
cc_190 N_A_81_268#_c_168_n N_A_232_162#_M1013_d 0.00326701f $X=1.495 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_191 N_A_81_268#_c_170_n N_A_232_162#_M1006_g 0.00698889f $X=2.335 $Y=0.34
+ $X2=0 $Y2=0
cc_192 N_A_81_268#_c_208_p N_A_232_162#_M1006_g 0.00610641f $X=2.5 $Y=0.545
+ $X2=0 $Y2=0
cc_193 N_A_81_268#_c_183_n N_A_232_162#_M1019_g 0.00445699f $X=2.49 $Y=2.795
+ $X2=0 $Y2=0
cc_194 N_A_81_268#_c_168_n N_A_232_162#_c_352_n 0.0373712f $X=1.495 $Y=0.745
+ $X2=0 $Y2=0
cc_195 N_A_81_268#_c_174_n N_A_232_162#_c_352_n 0.00740263f $X=0.605 $Y=1.34
+ $X2=0 $Y2=0
cc_196 N_A_81_268#_c_178_n N_A_232_162#_c_359_n 0.0136419f $X=1.06 $Y=2.905
+ $X2=0 $Y2=0
cc_197 N_A_81_268#_c_179_n N_A_232_162#_c_359_n 0.0134564f $X=2.325 $Y=2.99
+ $X2=0 $Y2=0
cc_198 N_A_81_268#_M1016_g N_X_c_862_n 0.00107274f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_199 N_A_81_268#_c_177_n N_X_c_858_n 0.00752377f $X=0.7 $Y=1.95 $X2=0 $Y2=0
cc_200 N_A_81_268#_c_172_n N_X_c_858_n 0.024967f $X=0.59 $Y=1.505 $X2=0 $Y2=0
cc_201 N_A_81_268#_c_173_n N_X_c_858_n 0.0114633f $X=0.59 $Y=1.505 $X2=0 $Y2=0
cc_202 N_A_81_268#_c_174_n N_X_c_858_n 0.00610084f $X=0.605 $Y=1.34 $X2=0 $Y2=0
cc_203 N_A_81_268#_c_175_n N_X_c_858_n 0.0030945f $X=0.58 $Y=1.34 $X2=0 $Y2=0
cc_204 N_A_81_268#_c_175_n X 0.012666f $X=0.58 $Y=1.34 $X2=0 $Y2=0
cc_205 N_A_81_268#_c_172_n X 0.00144434f $X=0.59 $Y=1.505 $X2=0 $Y2=0
cc_206 N_A_81_268#_c_175_n X 0.00238049f $X=0.58 $Y=1.34 $X2=0 $Y2=0
cc_207 N_A_81_268#_c_177_n N_VPWR_M1016_d 0.00217984f $X=0.7 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_208 N_A_81_268#_c_186_p N_VPWR_M1016_d 0.0161937f $X=0.975 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_209 N_A_81_268#_c_225_p N_VPWR_M1016_d 0.00284944f $X=0.785 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_210 N_A_81_268#_c_178_n N_VPWR_M1016_d 0.00442522f $X=1.06 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_211 N_A_81_268#_M1016_g N_VPWR_c_880_n 0.0170998f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_212 N_A_81_268#_c_186_p N_VPWR_c_880_n 0.00150934f $X=0.975 $Y=2.035 $X2=0
+ $Y2=0
cc_213 N_A_81_268#_c_225_p N_VPWR_c_880_n 0.0128481f $X=0.785 $Y=2.035 $X2=0
+ $Y2=0
cc_214 N_A_81_268#_c_178_n N_VPWR_c_880_n 0.0465257f $X=1.06 $Y=2.905 $X2=0
+ $Y2=0
cc_215 N_A_81_268#_c_180_n N_VPWR_c_880_n 0.0146661f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_216 N_A_81_268#_c_172_n N_VPWR_c_880_n 0.0011623f $X=0.59 $Y=1.505 $X2=0
+ $Y2=0
cc_217 N_A_81_268#_c_173_n N_VPWR_c_880_n 4.1218e-19 $X=0.59 $Y=1.505 $X2=0
+ $Y2=0
cc_218 N_A_81_268#_M1016_g N_VPWR_c_883_n 0.00460063f $X=0.495 $Y=2.4 $X2=0
+ $Y2=0
cc_219 N_A_81_268#_c_179_n N_VPWR_c_884_n 0.0759845f $X=2.325 $Y=2.99 $X2=0
+ $Y2=0
cc_220 N_A_81_268#_c_180_n N_VPWR_c_884_n 0.0121867f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_221 N_A_81_268#_c_183_n N_VPWR_c_884_n 0.0224527f $X=2.49 $Y=2.795 $X2=0
+ $Y2=0
cc_222 N_A_81_268#_M1016_g N_VPWR_c_879_n 0.00912261f $X=0.495 $Y=2.4 $X2=0
+ $Y2=0
cc_223 N_A_81_268#_c_179_n N_VPWR_c_879_n 0.0443614f $X=2.325 $Y=2.99 $X2=0
+ $Y2=0
cc_224 N_A_81_268#_c_180_n N_VPWR_c_879_n 0.00660921f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_225 N_A_81_268#_c_183_n N_VPWR_c_879_n 0.0125544f $X=2.49 $Y=2.795 $X2=0
+ $Y2=0
cc_226 N_A_81_268#_M1000_d N_A_363_394#_c_962_n 0.00965907f $X=2.275 $Y=1.97
+ $X2=0 $Y2=0
cc_227 N_A_81_268#_c_179_n N_A_363_394#_c_962_n 0.00586468f $X=2.325 $Y=2.99
+ $X2=0 $Y2=0
cc_228 N_A_81_268#_c_183_n N_A_363_394#_c_962_n 0.0234024f $X=2.49 $Y=2.795
+ $X2=0 $Y2=0
cc_229 N_A_81_268#_c_179_n N_A_363_394#_c_970_n 0.0168392f $X=2.325 $Y=2.99
+ $X2=0 $Y2=0
cc_230 N_A_81_268#_c_170_n N_A_363_394#_c_956_n 0.00397229f $X=2.335 $Y=0.34
+ $X2=0 $Y2=0
cc_231 N_A_81_268#_c_170_n N_A_371_74#_M1008_s 0.00273752f $X=2.335 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_232 N_A_81_268#_c_168_n N_A_371_74#_c_1086_n 0.0150383f $X=1.495 $Y=0.745
+ $X2=0 $Y2=0
cc_233 N_A_81_268#_c_169_n N_A_371_74#_c_1086_n 0.00511585f $X=1.58 $Y=0.66
+ $X2=0 $Y2=0
cc_234 N_A_81_268#_c_170_n N_A_371_74#_c_1086_n 0.020565f $X=2.335 $Y=0.34 $X2=0
+ $Y2=0
cc_235 N_A_81_268#_c_208_p N_A_371_74#_c_1087_n 0.0221626f $X=2.5 $Y=0.545 $X2=0
+ $Y2=0
cc_236 N_A_81_268#_c_208_p N_A_371_74#_c_1091_n 0.00229444f $X=2.5 $Y=0.545
+ $X2=0 $Y2=0
cc_237 N_A_81_268#_c_168_n N_VGND_M1003_d 0.00831043f $X=1.495 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_238 N_A_81_268#_c_254_p N_VGND_M1003_d 0.00317478f $X=0.785 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_239 N_A_81_268#_c_174_n N_VGND_M1003_d 0.00758042f $X=0.605 $Y=1.34 $X2=-0.19
+ $Y2=-0.245
cc_240 N_A_81_268#_c_168_n N_VGND_c_1327_n 0.0130057f $X=1.495 $Y=0.745 $X2=0
+ $Y2=0
cc_241 N_A_81_268#_c_254_p N_VGND_c_1327_n 0.0134514f $X=0.785 $Y=0.745 $X2=0
+ $Y2=0
cc_242 N_A_81_268#_c_169_n N_VGND_c_1327_n 0.00229662f $X=1.58 $Y=0.66 $X2=0
+ $Y2=0
cc_243 N_A_81_268#_c_171_n N_VGND_c_1327_n 0.00673184f $X=1.665 $Y=0.34 $X2=0
+ $Y2=0
cc_244 N_A_81_268#_c_175_n N_VGND_c_1327_n 0.00449249f $X=0.58 $Y=1.34 $X2=0
+ $Y2=0
cc_245 N_A_81_268#_c_175_n N_VGND_c_1330_n 0.00472938f $X=0.58 $Y=1.34 $X2=0
+ $Y2=0
cc_246 N_A_81_268#_c_168_n N_VGND_c_1331_n 0.00932679f $X=1.495 $Y=0.745 $X2=0
+ $Y2=0
cc_247 N_A_81_268#_c_170_n N_VGND_c_1331_n 0.0663235f $X=2.335 $Y=0.34 $X2=0
+ $Y2=0
cc_248 N_A_81_268#_c_171_n N_VGND_c_1331_n 0.0120335f $X=1.665 $Y=0.34 $X2=0
+ $Y2=0
cc_249 N_A_81_268#_c_168_n N_VGND_c_1334_n 0.0158896f $X=1.495 $Y=0.745 $X2=0
+ $Y2=0
cc_250 N_A_81_268#_c_254_p N_VGND_c_1334_n 0.00111722f $X=0.785 $Y=0.745 $X2=0
+ $Y2=0
cc_251 N_A_81_268#_c_170_n N_VGND_c_1334_n 0.0372321f $X=2.335 $Y=0.34 $X2=0
+ $Y2=0
cc_252 N_A_81_268#_c_171_n N_VGND_c_1334_n 0.00658039f $X=1.665 $Y=0.34 $X2=0
+ $Y2=0
cc_253 N_A_81_268#_c_175_n N_VGND_c_1334_n 0.00508379f $X=0.58 $Y=1.34 $X2=0
+ $Y2=0
cc_254 N_C_c_271_n N_A_232_162#_M1006_g 0.00796043f $X=2.185 $Y=1.59 $X2=0 $Y2=0
cc_255 N_C_c_273_n N_A_232_162#_M1006_g 0.0210141f $X=2.215 $Y=1.085 $X2=0 $Y2=0
cc_256 N_C_M1000_g N_A_232_162#_M1019_g 0.0311125f $X=2.185 $Y=2.39 $X2=0 $Y2=0
cc_257 N_C_c_271_n N_A_232_162#_c_352_n 3.82753e-19 $X=2.185 $Y=1.59 $X2=0 $Y2=0
cc_258 N_C_c_273_n N_A_232_162#_c_352_n 3.29455e-19 $X=2.215 $Y=1.085 $X2=0
+ $Y2=0
cc_259 N_C_c_274_n N_A_232_162#_c_352_n 0.00627487f $X=1.16 $Y=1.425 $X2=0 $Y2=0
cc_260 N_C_c_275_n N_A_232_162#_c_352_n 0.00311959f $X=1.16 $Y=1.35 $X2=0 $Y2=0
cc_261 N_C_c_276_n N_A_232_162#_c_352_n 0.0116105f $X=1.16 $Y=1.515 $X2=0 $Y2=0
cc_262 N_C_M1018_g N_A_232_162#_c_359_n 0.0032756f $X=1.175 $Y=2.16 $X2=0 $Y2=0
cc_263 N_C_c_270_n N_A_232_162#_c_359_n 0.0050076f $X=2.095 $Y=1.425 $X2=0 $Y2=0
cc_264 N_C_M1000_g N_A_232_162#_c_359_n 0.0012964f $X=2.185 $Y=2.39 $X2=0 $Y2=0
cc_265 N_C_c_276_n N_A_232_162#_c_359_n 4.37201e-19 $X=1.16 $Y=1.515 $X2=0 $Y2=0
cc_266 N_C_c_270_n N_A_232_162#_c_353_n 0.0165956f $X=2.095 $Y=1.425 $X2=0 $Y2=0
cc_267 N_C_c_271_n N_A_232_162#_c_353_n 0.00282714f $X=2.185 $Y=1.59 $X2=0 $Y2=0
cc_268 N_C_c_274_n N_A_232_162#_c_353_n 0.00179145f $X=1.16 $Y=1.425 $X2=0 $Y2=0
cc_269 N_C_c_275_n N_A_232_162#_c_353_n 0.00429029f $X=1.16 $Y=1.35 $X2=0 $Y2=0
cc_270 N_C_c_276_n N_A_232_162#_c_353_n 0.0166868f $X=1.16 $Y=1.515 $X2=0 $Y2=0
cc_271 N_C_M1018_g N_A_232_162#_c_360_n 0.00573469f $X=1.175 $Y=2.16 $X2=0 $Y2=0
cc_272 N_C_M1000_g N_A_232_162#_c_360_n 0.00528648f $X=2.185 $Y=2.39 $X2=0 $Y2=0
cc_273 N_C_c_276_n N_A_232_162#_c_360_n 0.00234061f $X=1.16 $Y=1.515 $X2=0 $Y2=0
cc_274 N_C_M1018_g N_A_232_162#_c_354_n 4.74074e-19 $X=1.175 $Y=2.16 $X2=0 $Y2=0
cc_275 N_C_c_274_n N_A_232_162#_c_354_n 0.00232957f $X=1.16 $Y=1.425 $X2=0 $Y2=0
cc_276 N_C_c_276_n N_A_232_162#_c_354_n 0.0146247f $X=1.16 $Y=1.515 $X2=0 $Y2=0
cc_277 N_C_c_271_n N_A_232_162#_c_355_n 6.70353e-19 $X=2.185 $Y=1.59 $X2=0 $Y2=0
cc_278 N_C_M1000_g N_A_232_162#_c_355_n 3.89547e-19 $X=2.185 $Y=2.39 $X2=0 $Y2=0
cc_279 N_C_c_271_n N_A_232_162#_c_356_n 0.0174697f $X=2.185 $Y=1.59 $X2=0 $Y2=0
cc_280 N_C_c_270_n N_A_232_162#_c_357_n 0.0126387f $X=2.095 $Y=1.425 $X2=0 $Y2=0
cc_281 N_C_c_271_n N_A_232_162#_c_357_n 0.0027142f $X=2.185 $Y=1.59 $X2=0 $Y2=0
cc_282 N_C_M1000_g N_A_232_162#_c_357_n 0.0125626f $X=2.185 $Y=2.39 $X2=0 $Y2=0
cc_283 N_C_M1018_g N_VPWR_c_880_n 9.65328e-19 $X=1.175 $Y=2.16 $X2=0 $Y2=0
cc_284 N_C_M1018_g N_VPWR_c_884_n 2.1643e-19 $X=1.175 $Y=2.16 $X2=0 $Y2=0
cc_285 N_C_M1000_g N_VPWR_c_884_n 8.10111e-19 $X=2.185 $Y=2.39 $X2=0 $Y2=0
cc_286 N_C_M1000_g N_A_363_394#_c_961_n 0.0106523f $X=2.185 $Y=2.39 $X2=0 $Y2=0
cc_287 N_C_M1000_g N_A_363_394#_c_962_n 0.0122408f $X=2.185 $Y=2.39 $X2=0 $Y2=0
cc_288 N_C_M1018_g N_A_363_394#_c_970_n 0.00290352f $X=1.175 $Y=2.16 $X2=0 $Y2=0
cc_289 N_C_M1000_g N_A_363_394#_c_970_n 0.00483343f $X=2.185 $Y=2.39 $X2=0 $Y2=0
cc_290 N_C_c_271_n N_A_371_74#_c_1086_n 0.00333638f $X=2.185 $Y=1.59 $X2=0 $Y2=0
cc_291 N_C_c_273_n N_A_371_74#_c_1086_n 0.0083827f $X=2.215 $Y=1.085 $X2=0 $Y2=0
cc_292 N_C_c_275_n N_A_371_74#_c_1086_n 0.00307068f $X=1.16 $Y=1.35 $X2=0 $Y2=0
cc_293 N_C_c_271_n N_A_371_74#_c_1087_n 0.00273799f $X=2.185 $Y=1.59 $X2=0 $Y2=0
cc_294 N_C_M1000_g N_A_371_74#_c_1098_n 7.51826e-19 $X=2.185 $Y=2.39 $X2=0 $Y2=0
cc_295 N_C_c_270_n N_A_371_74#_c_1092_n 6.37321e-19 $X=2.095 $Y=1.425 $X2=0
+ $Y2=0
cc_296 N_C_c_271_n N_A_371_74#_c_1092_n 0.00142091f $X=2.185 $Y=1.59 $X2=0 $Y2=0
cc_297 N_C_c_270_n N_A_371_74#_c_1094_n 0.00800485f $X=2.095 $Y=1.425 $X2=0
+ $Y2=0
cc_298 N_C_c_271_n N_A_371_74#_c_1094_n 0.01602f $X=2.185 $Y=1.59 $X2=0 $Y2=0
cc_299 N_C_c_273_n N_VGND_c_1331_n 0.00278271f $X=2.215 $Y=1.085 $X2=0 $Y2=0
cc_300 N_C_c_275_n N_VGND_c_1331_n 5.51389e-19 $X=1.16 $Y=1.35 $X2=0 $Y2=0
cc_301 N_C_c_273_n N_VGND_c_1334_n 0.00359139f $X=2.215 $Y=1.085 $X2=0 $Y2=0
cc_302 N_A_232_162#_M1019_g N_VPWR_c_881_n 0.00606038f $X=2.79 $Y=2.39 $X2=0
+ $Y2=0
cc_303 N_A_232_162#_M1019_g N_VPWR_c_884_n 0.00570207f $X=2.79 $Y=2.39 $X2=0
+ $Y2=0
cc_304 N_A_232_162#_M1019_g N_VPWR_c_879_n 0.00599321f $X=2.79 $Y=2.39 $X2=0
+ $Y2=0
cc_305 N_A_232_162#_M1019_g N_A_363_394#_c_961_n 0.00188086f $X=2.79 $Y=2.39
+ $X2=0 $Y2=0
cc_306 N_A_232_162#_c_359_n N_A_363_394#_c_961_n 0.0289958f $X=1.49 $Y=2.125
+ $X2=0 $Y2=0
cc_307 N_A_232_162#_c_357_n N_A_363_394#_c_961_n 0.0180255f $X=2.515 $Y=1.645
+ $X2=0 $Y2=0
cc_308 N_A_232_162#_M1019_g N_A_363_394#_c_962_n 0.0178883f $X=2.79 $Y=2.39
+ $X2=0 $Y2=0
cc_309 N_A_232_162#_c_355_n N_A_363_394#_c_962_n 0.00840336f $X=2.68 $Y=1.645
+ $X2=0 $Y2=0
cc_310 N_A_232_162#_c_356_n N_A_363_394#_c_962_n 0.00305432f $X=2.68 $Y=1.645
+ $X2=0 $Y2=0
cc_311 N_A_232_162#_c_357_n N_A_363_394#_c_962_n 0.00964131f $X=2.515 $Y=1.645
+ $X2=0 $Y2=0
cc_312 N_A_232_162#_M1019_g N_A_363_394#_c_970_n 7.68714e-19 $X=2.79 $Y=2.39
+ $X2=0 $Y2=0
cc_313 N_A_232_162#_c_359_n N_A_363_394#_c_970_n 0.00971033f $X=1.49 $Y=2.125
+ $X2=0 $Y2=0
cc_314 N_A_232_162#_M1006_g N_A_363_394#_c_955_n 0.0045144f $X=2.715 $Y=0.69
+ $X2=0 $Y2=0
cc_315 N_A_232_162#_M1019_g N_A_363_394#_c_955_n 0.00290623f $X=2.79 $Y=2.39
+ $X2=0 $Y2=0
cc_316 N_A_232_162#_M1006_g N_A_363_394#_c_956_n 0.00549115f $X=2.715 $Y=0.69
+ $X2=0 $Y2=0
cc_317 N_A_232_162#_M1006_g N_A_371_74#_c_1086_n 7.04872e-19 $X=2.715 $Y=0.69
+ $X2=0 $Y2=0
cc_318 N_A_232_162#_c_352_n N_A_371_74#_c_1086_n 0.0147639f $X=1.495 $Y=1.085
+ $X2=0 $Y2=0
cc_319 N_A_232_162#_M1006_g N_A_371_74#_c_1087_n 0.0153345f $X=2.715 $Y=0.69
+ $X2=0 $Y2=0
cc_320 N_A_232_162#_c_355_n N_A_371_74#_c_1087_n 0.0210253f $X=2.68 $Y=1.645
+ $X2=0 $Y2=0
cc_321 N_A_232_162#_c_356_n N_A_371_74#_c_1087_n 0.00549164f $X=2.68 $Y=1.645
+ $X2=0 $Y2=0
cc_322 N_A_232_162#_c_357_n N_A_371_74#_c_1087_n 0.00974989f $X=2.515 $Y=1.645
+ $X2=0 $Y2=0
cc_323 N_A_232_162#_M1006_g N_A_371_74#_c_1088_n 0.00503563f $X=2.715 $Y=0.69
+ $X2=0 $Y2=0
cc_324 N_A_232_162#_c_355_n N_A_371_74#_c_1088_n 0.0255178f $X=2.68 $Y=1.645
+ $X2=0 $Y2=0
cc_325 N_A_232_162#_c_356_n N_A_371_74#_c_1088_n 0.0147692f $X=2.68 $Y=1.645
+ $X2=0 $Y2=0
cc_326 N_A_232_162#_M1019_g N_A_371_74#_c_1098_n 0.00523852f $X=2.79 $Y=2.39
+ $X2=0 $Y2=0
cc_327 N_A_232_162#_M1006_g N_A_371_74#_c_1091_n 0.00257359f $X=2.715 $Y=0.69
+ $X2=0 $Y2=0
cc_328 N_A_232_162#_c_355_n N_A_371_74#_c_1091_n 0.00827532f $X=2.68 $Y=1.645
+ $X2=0 $Y2=0
cc_329 N_A_232_162#_c_356_n N_A_371_74#_c_1091_n 0.00570681f $X=2.68 $Y=1.645
+ $X2=0 $Y2=0
cc_330 N_A_232_162#_c_357_n N_A_371_74#_c_1091_n 0.00531172f $X=2.515 $Y=1.645
+ $X2=0 $Y2=0
cc_331 N_A_232_162#_M1006_g N_A_371_74#_c_1092_n 6.38547e-19 $X=2.715 $Y=0.69
+ $X2=0 $Y2=0
cc_332 N_A_232_162#_c_353_n N_A_371_74#_c_1092_n 0.00109031f $X=1.58 $Y=1.58
+ $X2=0 $Y2=0
cc_333 N_A_232_162#_c_357_n N_A_371_74#_c_1092_n 0.00281376f $X=2.515 $Y=1.645
+ $X2=0 $Y2=0
cc_334 N_A_232_162#_M1006_g N_A_371_74#_c_1094_n 0.00147437f $X=2.715 $Y=0.69
+ $X2=0 $Y2=0
cc_335 N_A_232_162#_c_353_n N_A_371_74#_c_1094_n 0.0179576f $X=1.58 $Y=1.58
+ $X2=0 $Y2=0
cc_336 N_A_232_162#_c_357_n N_A_371_74#_c_1094_n 0.0303395f $X=2.515 $Y=1.645
+ $X2=0 $Y2=0
cc_337 N_A_232_162#_M1006_g N_VGND_c_1328_n 0.00277695f $X=2.715 $Y=0.69 $X2=0
+ $Y2=0
cc_338 N_A_232_162#_M1006_g N_VGND_c_1331_n 0.00430908f $X=2.715 $Y=0.69 $X2=0
+ $Y2=0
cc_339 N_A_232_162#_M1006_g N_VGND_c_1334_n 0.00822378f $X=2.715 $Y=0.69 $X2=0
+ $Y2=0
cc_340 N_A_786_100#_c_452_n N_B_M1002_g 0.00514817f $X=4.545 $Y=2.075 $X2=0
+ $Y2=0
cc_341 N_A_786_100#_c_446_n N_B_c_561_n 0.00333872f $X=4.545 $Y=1.095 $X2=0
+ $Y2=0
cc_342 N_A_786_100#_c_447_n N_B_c_561_n 0.00192933f $X=4.63 $Y=1.355 $X2=0 $Y2=0
cc_343 N_A_786_100#_M1009_g N_B_c_568_n 0.0288554f $X=4.955 $Y=2.285 $X2=0 $Y2=0
cc_344 N_A_786_100#_c_452_n N_B_c_568_n 0.0150487f $X=4.545 $Y=2.075 $X2=0 $Y2=0
cc_345 N_A_786_100#_c_453_n N_B_c_568_n 0.00484464f $X=4.63 $Y=1.95 $X2=0 $Y2=0
cc_346 N_A_786_100#_M1009_g N_B_c_569_n 0.00885431f $X=4.955 $Y=2.285 $X2=0
+ $Y2=0
cc_347 N_A_786_100#_M1012_g N_B_M1010_g 0.0213094f $X=5.94 $Y=2.235 $X2=0 $Y2=0
cc_348 N_A_786_100#_M1007_g N_B_M1004_g 0.0345711f $X=4.97 $Y=0.925 $X2=0 $Y2=0
cc_349 N_A_786_100#_c_441_n N_B_M1004_g 0.00976806f $X=6.02 $Y=0.19 $X2=0 $Y2=0
cc_350 N_A_786_100#_M1021_g N_B_M1004_g 0.0194751f $X=6.095 $Y=1.035 $X2=0 $Y2=0
cc_351 N_A_786_100#_c_445_n N_B_M1004_g 0.013752f $X=6.095 $Y=1.395 $X2=0 $Y2=0
cc_352 N_A_786_100#_c_448_n N_B_M1004_g 3.9608e-19 $X=4.88 $Y=1.52 $X2=0 $Y2=0
cc_353 N_A_786_100#_M1012_g N_B_c_573_n 0.00453622f $X=5.94 $Y=2.235 $X2=0 $Y2=0
cc_354 N_A_786_100#_M1012_g N_B_c_574_n 0.0176707f $X=5.94 $Y=2.235 $X2=0 $Y2=0
cc_355 N_A_786_100#_M1012_g N_B_M1014_g 0.00437779f $X=5.94 $Y=2.235 $X2=0 $Y2=0
cc_356 N_A_786_100#_M1021_g N_B_M1014_g 0.0269381f $X=6.095 $Y=1.035 $X2=0 $Y2=0
cc_357 N_A_786_100#_c_446_n N_B_c_564_n 0.00296978f $X=4.545 $Y=1.095 $X2=0
+ $Y2=0
cc_358 N_A_786_100#_c_446_n N_B_c_565_n 0.00238963f $X=4.545 $Y=1.095 $X2=0
+ $Y2=0
cc_359 N_A_786_100#_c_452_n N_B_c_565_n 9.25649e-19 $X=4.545 $Y=2.075 $X2=0
+ $Y2=0
cc_360 N_A_786_100#_c_448_n N_B_c_565_n 0.00277533f $X=4.88 $Y=1.52 $X2=0 $Y2=0
cc_361 N_A_786_100#_c_449_n N_B_c_565_n 0.0156257f $X=4.88 $Y=1.52 $X2=0 $Y2=0
cc_362 N_A_786_100#_M1009_g N_B_c_579_n 0.0239375f $X=4.955 $Y=2.285 $X2=0 $Y2=0
cc_363 N_A_786_100#_M1012_g N_B_c_579_n 0.013752f $X=5.94 $Y=2.235 $X2=0 $Y2=0
cc_364 N_A_786_100#_c_446_n N_B_c_566_n 0.0272396f $X=4.545 $Y=1.095 $X2=0 $Y2=0
cc_365 N_A_786_100#_c_452_n N_B_c_566_n 0.0336771f $X=4.545 $Y=2.075 $X2=0 $Y2=0
cc_366 N_A_786_100#_c_447_n N_B_c_566_n 3.40445e-19 $X=4.63 $Y=1.355 $X2=0 $Y2=0
cc_367 N_A_786_100#_c_453_n N_B_c_566_n 0.00754671f $X=4.63 $Y=1.95 $X2=0 $Y2=0
cc_368 N_A_786_100#_c_448_n N_B_c_566_n 0.0281881f $X=4.88 $Y=1.52 $X2=0 $Y2=0
cc_369 N_A_786_100#_c_449_n N_B_c_566_n 2.82342e-19 $X=4.88 $Y=1.52 $X2=0 $Y2=0
cc_370 N_A_786_100#_c_446_n N_A_897_54#_M1007_s 0.00713947f $X=4.545 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_371 N_A_786_100#_c_447_n N_A_897_54#_M1007_s 0.00190522f $X=4.63 $Y=1.355
+ $X2=-0.19 $Y2=-0.245
cc_372 N_A_786_100#_c_452_n N_A_897_54#_M1009_s 0.00657014f $X=4.545 $Y=2.075
+ $X2=0 $Y2=0
cc_373 N_A_786_100#_c_453_n N_A_897_54#_M1009_s 0.00223036f $X=4.63 $Y=1.95
+ $X2=0 $Y2=0
cc_374 N_A_786_100#_M1009_g N_A_897_54#_c_742_n 0.00185504f $X=4.955 $Y=2.285
+ $X2=0 $Y2=0
cc_375 N_A_786_100#_M1012_g N_A_897_54#_c_742_n 5.48752e-19 $X=5.94 $Y=2.235
+ $X2=0 $Y2=0
cc_376 N_A_786_100#_M1007_g N_A_897_54#_c_734_n 0.0118793f $X=4.97 $Y=0.925
+ $X2=0 $Y2=0
cc_377 N_A_786_100#_c_441_n N_A_897_54#_c_734_n 0.0227936f $X=6.02 $Y=0.19 $X2=0
+ $Y2=0
cc_378 N_A_786_100#_c_442_n N_A_897_54#_c_734_n 0.00158085f $X=5.045 $Y=0.19
+ $X2=0 $Y2=0
cc_379 N_A_786_100#_M1021_g N_A_897_54#_c_734_n 0.0118974f $X=6.095 $Y=1.035
+ $X2=0 $Y2=0
cc_380 N_A_786_100#_M1021_g N_A_897_54#_c_735_n 0.00150595f $X=6.095 $Y=1.035
+ $X2=0 $Y2=0
cc_381 N_A_786_100#_M1007_g N_A_897_54#_c_738_n 0.00316796f $X=4.97 $Y=0.925
+ $X2=0 $Y2=0
cc_382 N_A_786_100#_M1009_g N_A_897_54#_c_745_n 0.00368534f $X=4.955 $Y=2.285
+ $X2=0 $Y2=0
cc_383 N_A_786_100#_c_446_n N_A_363_394#_c_955_n 0.00707775f $X=4.545 $Y=1.095
+ $X2=0 $Y2=0
cc_384 N_A_786_100#_c_452_n N_A_363_394#_c_955_n 0.0101325f $X=4.545 $Y=2.075
+ $X2=0 $Y2=0
cc_385 N_A_786_100#_M1002_d N_A_363_394#_c_964_n 0.00625031f $X=3.95 $Y=1.84
+ $X2=0 $Y2=0
cc_386 N_A_786_100#_M1009_g N_A_363_394#_c_964_n 0.0155514f $X=4.955 $Y=2.285
+ $X2=0 $Y2=0
cc_387 N_A_786_100#_c_452_n N_A_363_394#_c_964_n 0.0553716f $X=4.545 $Y=2.075
+ $X2=0 $Y2=0
cc_388 N_A_786_100#_c_449_n N_A_363_394#_c_964_n 0.00273546f $X=4.88 $Y=1.52
+ $X2=0 $Y2=0
cc_389 N_A_786_100#_M1009_g N_A_363_394#_c_965_n 0.00893761f $X=4.955 $Y=2.285
+ $X2=0 $Y2=0
cc_390 N_A_786_100#_c_452_n N_A_363_394#_c_965_n 0.0130957f $X=4.545 $Y=2.075
+ $X2=0 $Y2=0
cc_391 N_A_786_100#_c_453_n N_A_363_394#_c_965_n 0.00443076f $X=4.63 $Y=1.95
+ $X2=0 $Y2=0
cc_392 N_A_786_100#_c_448_n N_A_363_394#_c_965_n 0.00223621f $X=4.88 $Y=1.52
+ $X2=0 $Y2=0
cc_393 N_A_786_100#_c_441_n N_A_363_394#_c_957_n 0.0016693f $X=6.02 $Y=0.19
+ $X2=0 $Y2=0
cc_394 N_A_786_100#_M1021_g N_A_363_394#_c_957_n 0.0125058f $X=6.095 $Y=1.035
+ $X2=0 $Y2=0
cc_395 N_A_786_100#_c_445_n N_A_363_394#_c_957_n 5.29597e-19 $X=6.095 $Y=1.395
+ $X2=0 $Y2=0
cc_396 N_A_786_100#_M1021_g N_A_363_394#_c_958_n 0.00652313f $X=6.095 $Y=1.035
+ $X2=0 $Y2=0
cc_397 N_A_786_100#_M1001_d N_A_363_394#_c_959_n 0.00718532f $X=3.93 $Y=0.5
+ $X2=0 $Y2=0
cc_398 N_A_786_100#_M1007_g N_A_363_394#_c_959_n 0.0104707f $X=4.97 $Y=0.925
+ $X2=0 $Y2=0
cc_399 N_A_786_100#_c_446_n N_A_363_394#_c_959_n 0.0530741f $X=4.545 $Y=1.095
+ $X2=0 $Y2=0
cc_400 N_A_786_100#_c_448_n N_A_363_394#_c_959_n 0.00420626f $X=4.88 $Y=1.52
+ $X2=0 $Y2=0
cc_401 N_A_786_100#_c_449_n N_A_363_394#_c_959_n 0.00186709f $X=4.88 $Y=1.52
+ $X2=0 $Y2=0
cc_402 N_A_786_100#_M1007_g N_A_363_394#_c_960_n 0.00855512f $X=4.97 $Y=0.925
+ $X2=0 $Y2=0
cc_403 N_A_786_100#_c_441_n N_A_363_394#_c_960_n 0.00158035f $X=6.02 $Y=0.19
+ $X2=0 $Y2=0
cc_404 N_A_786_100#_M1007_g N_A_371_74#_c_1134_n 0.00559226f $X=4.97 $Y=0.925
+ $X2=0 $Y2=0
cc_405 N_A_786_100#_c_446_n N_A_371_74#_c_1134_n 0.00887711f $X=4.545 $Y=1.095
+ $X2=0 $Y2=0
cc_406 N_A_786_100#_c_448_n N_A_371_74#_c_1134_n 0.00147344f $X=4.88 $Y=1.52
+ $X2=0 $Y2=0
cc_407 N_A_786_100#_M1007_g N_A_371_74#_c_1089_n 0.0013539f $X=4.97 $Y=0.925
+ $X2=0 $Y2=0
cc_408 N_A_786_100#_c_447_n N_A_371_74#_c_1089_n 0.0033787f $X=4.63 $Y=1.355
+ $X2=0 $Y2=0
cc_409 N_A_786_100#_c_448_n N_A_371_74#_c_1089_n 0.00263929f $X=4.88 $Y=1.52
+ $X2=0 $Y2=0
cc_410 N_A_786_100#_c_449_n N_A_371_74#_c_1089_n 2.10143e-19 $X=4.88 $Y=1.52
+ $X2=0 $Y2=0
cc_411 N_A_786_100#_M1009_g N_A_371_74#_c_1090_n 4.25321e-19 $X=4.955 $Y=2.285
+ $X2=0 $Y2=0
cc_412 N_A_786_100#_M1012_g N_A_371_74#_c_1090_n 0.00110998f $X=5.94 $Y=2.235
+ $X2=0 $Y2=0
cc_413 N_A_786_100#_c_445_n N_A_371_74#_c_1090_n 2.04704e-19 $X=6.095 $Y=1.395
+ $X2=0 $Y2=0
cc_414 N_A_786_100#_c_448_n N_A_371_74#_c_1090_n 0.0114271f $X=4.88 $Y=1.52
+ $X2=0 $Y2=0
cc_415 N_A_786_100#_c_449_n N_A_371_74#_c_1090_n 0.00111824f $X=4.88 $Y=1.52
+ $X2=0 $Y2=0
cc_416 N_A_786_100#_M1012_g N_A_371_74#_c_1097_n 0.0137687f $X=5.94 $Y=2.235
+ $X2=0 $Y2=0
cc_417 N_A_786_100#_c_445_n N_A_371_74#_c_1097_n 7.82653e-19 $X=6.095 $Y=1.395
+ $X2=0 $Y2=0
cc_418 N_A_786_100#_M1009_g N_A_371_74#_c_1148_n 5.31738e-19 $X=4.955 $Y=2.285
+ $X2=0 $Y2=0
cc_419 N_A_786_100#_M1001_d N_A_371_74#_c_1091_n 0.00209695f $X=3.93 $Y=0.5
+ $X2=0 $Y2=0
cc_420 N_A_786_100#_M1007_g N_A_371_74#_c_1091_n 0.0049795f $X=4.97 $Y=0.925
+ $X2=0 $Y2=0
cc_421 N_A_786_100#_c_446_n N_A_371_74#_c_1091_n 0.0222819f $X=4.545 $Y=1.095
+ $X2=0 $Y2=0
cc_422 N_A_786_100#_c_452_n N_A_371_74#_c_1091_n 0.00652339f $X=4.545 $Y=2.075
+ $X2=0 $Y2=0
cc_423 N_A_786_100#_c_447_n N_A_371_74#_c_1091_n 0.0123134f $X=4.63 $Y=1.355
+ $X2=0 $Y2=0
cc_424 N_A_786_100#_c_453_n N_A_371_74#_c_1091_n 5.40026e-19 $X=4.63 $Y=1.95
+ $X2=0 $Y2=0
cc_425 N_A_786_100#_c_448_n N_A_371_74#_c_1091_n 0.0219425f $X=4.88 $Y=1.52
+ $X2=0 $Y2=0
cc_426 N_A_786_100#_c_449_n N_A_371_74#_c_1091_n 0.0019248f $X=4.88 $Y=1.52
+ $X2=0 $Y2=0
cc_427 N_A_786_100#_c_448_n N_A_371_74#_c_1093_n 2.88257e-19 $X=4.88 $Y=1.52
+ $X2=0 $Y2=0
cc_428 N_A_786_100#_M1012_g N_A_1116_383#_c_1227_n 0.0083658f $X=5.94 $Y=2.235
+ $X2=0 $Y2=0
cc_429 N_A_786_100#_M1012_g N_A_1116_383#_c_1221_n 0.00884366f $X=5.94 $Y=2.235
+ $X2=0 $Y2=0
cc_430 N_A_786_100#_M1009_g N_A_1116_383#_c_1222_n 6.61361e-19 $X=4.955 $Y=2.285
+ $X2=0 $Y2=0
cc_431 N_A_786_100#_M1012_g N_A_1116_383#_c_1222_n 0.00190631f $X=5.94 $Y=2.235
+ $X2=0 $Y2=0
cc_432 N_A_786_100#_c_445_n N_A_1116_383#_c_1212_n 0.00441754f $X=6.095 $Y=1.395
+ $X2=0 $Y2=0
cc_433 N_A_786_100#_M1012_g N_A_1116_383#_c_1213_n 0.00739982f $X=5.94 $Y=2.235
+ $X2=0 $Y2=0
cc_434 N_A_786_100#_c_445_n N_A_1116_383#_c_1213_n 0.00211835f $X=6.095 $Y=1.395
+ $X2=0 $Y2=0
cc_435 N_A_786_100#_M1012_g N_A_1116_383#_c_1214_n 0.00527609f $X=5.94 $Y=2.235
+ $X2=0 $Y2=0
cc_436 N_A_786_100#_M1021_g N_A_1116_383#_c_1217_n 0.00100578f $X=6.095 $Y=1.035
+ $X2=0 $Y2=0
cc_437 N_A_786_100#_c_445_n N_A_1116_383#_c_1217_n 5.09731e-19 $X=6.095 $Y=1.395
+ $X2=0 $Y2=0
cc_438 N_A_786_100#_M1021_g N_A_1116_383#_c_1237_n 0.00119336f $X=6.095 $Y=1.035
+ $X2=0 $Y2=0
cc_439 N_A_786_100#_c_445_n N_A_1116_383#_c_1237_n 0.00120579f $X=6.095 $Y=1.395
+ $X2=0 $Y2=0
cc_440 N_A_786_100#_M1021_g N_A_1116_383#_c_1220_n 0.00758454f $X=6.095 $Y=1.035
+ $X2=0 $Y2=0
cc_441 N_A_786_100#_c_445_n N_A_1116_383#_c_1220_n 0.00826216f $X=6.095 $Y=1.395
+ $X2=0 $Y2=0
cc_442 N_A_786_100#_c_442_n N_VGND_c_1332_n 0.0269013f $X=5.045 $Y=0.19 $X2=0
+ $Y2=0
cc_443 N_A_786_100#_c_441_n N_VGND_c_1334_n 0.0289061f $X=6.02 $Y=0.19 $X2=0
+ $Y2=0
cc_444 N_A_786_100#_c_442_n N_VGND_c_1334_n 0.00589078f $X=5.045 $Y=0.19 $X2=0
+ $Y2=0
cc_445 N_B_M1014_g N_A_M1017_g 0.0195015f $X=6.59 $Y=0.925 $X2=0 $Y2=0
cc_446 N_B_c_574_n N_A_M1020_g 0.0261275f $X=6.575 $Y=1.78 $X2=0 $Y2=0
cc_447 N_B_M1014_g A 0.00224111f $X=6.59 $Y=0.925 $X2=0 $Y2=0
cc_448 N_B_M1014_g N_A_c_691_n 0.0195721f $X=6.59 $Y=0.925 $X2=0 $Y2=0
cc_449 N_B_c_569_n N_A_897_54#_c_742_n 0.00858512f $X=5.4 $Y=3.15 $X2=0 $Y2=0
cc_450 N_B_M1010_g N_A_897_54#_c_742_n 0.0193961f $X=5.49 $Y=2.235 $X2=0 $Y2=0
cc_451 N_B_c_573_n N_A_897_54#_c_742_n 0.0144892f $X=6.485 $Y=3.15 $X2=0 $Y2=0
cc_452 N_B_M1015_g N_A_897_54#_c_742_n 0.0158143f $X=6.575 $Y=2.335 $X2=0 $Y2=0
cc_453 N_B_M1004_g N_A_897_54#_c_734_n 0.00112634f $X=5.535 $Y=0.925 $X2=0 $Y2=0
cc_454 N_B_M1014_g N_A_897_54#_c_734_n 0.00675742f $X=6.59 $Y=0.925 $X2=0 $Y2=0
cc_455 N_B_M1014_g N_A_897_54#_c_735_n 0.00599706f $X=6.59 $Y=0.925 $X2=0 $Y2=0
cc_456 N_B_M1015_g N_A_897_54#_c_767_n 0.00146039f $X=6.575 $Y=2.335 $X2=0 $Y2=0
cc_457 N_B_M1015_g N_A_897_54#_c_743_n 0.0094779f $X=6.575 $Y=2.335 $X2=0 $Y2=0
cc_458 N_B_M1014_g N_A_897_54#_c_737_n 0.00103773f $X=6.59 $Y=0.925 $X2=0 $Y2=0
cc_459 N_B_c_561_n N_A_897_54#_c_738_n 0.00345214f $X=3.855 $Y=1.35 $X2=0 $Y2=0
cc_460 N_B_c_568_n N_A_897_54#_c_745_n 0.0138382f $X=4.37 $Y=3.075 $X2=0 $Y2=0
cc_461 N_B_c_569_n N_A_897_54#_c_745_n 0.00878911f $X=5.4 $Y=3.15 $X2=0 $Y2=0
cc_462 N_B_M1010_g N_A_897_54#_c_745_n 0.00235329f $X=5.49 $Y=2.235 $X2=0 $Y2=0
cc_463 N_B_M1002_g N_VPWR_c_881_n 0.01062f $X=3.86 $Y=2.4 $X2=0 $Y2=0
cc_464 N_B_c_568_n N_VPWR_c_881_n 0.00283118f $X=4.37 $Y=3.075 $X2=0 $Y2=0
cc_465 N_B_c_573_n N_VPWR_c_882_n 0.00234767f $X=6.485 $Y=3.15 $X2=0 $Y2=0
cc_466 N_B_M1002_g N_VPWR_c_885_n 0.00553757f $X=3.86 $Y=2.4 $X2=0 $Y2=0
cc_467 N_B_c_570_n N_VPWR_c_885_n 0.0538526f $X=4.445 $Y=3.15 $X2=0 $Y2=0
cc_468 N_B_M1002_g N_VPWR_c_879_n 0.0054573f $X=3.86 $Y=2.4 $X2=0 $Y2=0
cc_469 N_B_c_569_n N_VPWR_c_879_n 0.022748f $X=5.4 $Y=3.15 $X2=0 $Y2=0
cc_470 N_B_c_570_n N_VPWR_c_879_n 0.00698515f $X=4.445 $Y=3.15 $X2=0 $Y2=0
cc_471 N_B_c_573_n N_VPWR_c_879_n 0.0280817f $X=6.485 $Y=3.15 $X2=0 $Y2=0
cc_472 N_B_c_580_n N_VPWR_c_879_n 0.00445015f $X=5.49 $Y=3.15 $X2=0 $Y2=0
cc_473 N_B_M1002_g N_A_363_394#_c_955_n 0.0166339f $X=3.86 $Y=2.4 $X2=0 $Y2=0
cc_474 N_B_c_561_n N_A_363_394#_c_955_n 0.00884203f $X=3.855 $Y=1.35 $X2=0 $Y2=0
cc_475 N_B_c_564_n N_A_363_394#_c_955_n 0.00851193f $X=3.827 $Y=1.515 $X2=0
+ $Y2=0
cc_476 N_B_c_566_n N_A_363_394#_c_955_n 0.0329945f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_477 N_B_c_561_n N_A_363_394#_c_956_n 0.0090312f $X=3.855 $Y=1.35 $X2=0 $Y2=0
cc_478 N_B_M1002_g N_A_363_394#_c_964_n 0.0177051f $X=3.86 $Y=2.4 $X2=0 $Y2=0
cc_479 N_B_c_568_n N_A_363_394#_c_964_n 0.0130658f $X=4.37 $Y=3.075 $X2=0 $Y2=0
cc_480 N_B_c_569_n N_A_363_394#_c_964_n 9.2662e-19 $X=5.4 $Y=3.15 $X2=0 $Y2=0
cc_481 N_B_M1010_g N_A_363_394#_c_964_n 0.00197533f $X=5.49 $Y=2.235 $X2=0 $Y2=0
cc_482 N_B_c_566_n N_A_363_394#_c_964_n 0.00519529f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_483 N_B_c_568_n N_A_363_394#_c_965_n 9.68017e-19 $X=4.37 $Y=3.075 $X2=0 $Y2=0
cc_484 N_B_M1010_g N_A_363_394#_c_965_n 0.00699929f $X=5.49 $Y=2.235 $X2=0 $Y2=0
cc_485 N_B_M1004_g N_A_363_394#_c_957_n 0.0118759f $X=5.535 $Y=0.925 $X2=0 $Y2=0
cc_486 N_B_M1014_g N_A_363_394#_c_957_n 0.00419855f $X=6.59 $Y=0.925 $X2=0 $Y2=0
cc_487 N_B_M1014_g N_A_363_394#_c_958_n 0.00559764f $X=6.59 $Y=0.925 $X2=0 $Y2=0
cc_488 N_B_c_561_n N_A_363_394#_c_959_n 0.0169531f $X=3.855 $Y=1.35 $X2=0 $Y2=0
cc_489 N_B_c_564_n N_A_363_394#_c_959_n 2.19057e-19 $X=3.827 $Y=1.515 $X2=0
+ $Y2=0
cc_490 N_B_c_566_n N_A_363_394#_c_959_n 0.00256354f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_491 N_B_M1004_g N_A_363_394#_c_960_n 0.00187562f $X=5.535 $Y=0.925 $X2=0
+ $Y2=0
cc_492 N_B_M1004_g N_A_371_74#_c_1089_n 0.0127113f $X=5.535 $Y=0.925 $X2=0 $Y2=0
cc_493 N_B_c_579_n N_A_371_74#_c_1089_n 0.00119047f $X=5.505 $Y=1.84 $X2=0 $Y2=0
cc_494 N_B_M1004_g N_A_371_74#_c_1090_n 0.00754317f $X=5.535 $Y=0.925 $X2=0
+ $Y2=0
cc_495 N_B_c_579_n N_A_371_74#_c_1090_n 0.00371189f $X=5.505 $Y=1.84 $X2=0 $Y2=0
cc_496 N_B_c_574_n N_A_371_74#_c_1097_n 6.52488e-19 $X=6.575 $Y=1.78 $X2=0 $Y2=0
cc_497 N_B_c_579_n N_A_371_74#_c_1097_n 7.85122e-19 $X=5.505 $Y=1.84 $X2=0 $Y2=0
cc_498 N_B_M1010_g N_A_371_74#_c_1148_n 0.00946299f $X=5.49 $Y=2.235 $X2=0 $Y2=0
cc_499 N_B_c_579_n N_A_371_74#_c_1148_n 0.00286139f $X=5.505 $Y=1.84 $X2=0 $Y2=0
cc_500 N_B_M1015_g N_A_371_74#_c_1166_n 0.00141949f $X=6.575 $Y=2.335 $X2=0
+ $Y2=0
cc_501 N_B_c_561_n N_A_371_74#_c_1091_n 0.00556825f $X=3.855 $Y=1.35 $X2=0 $Y2=0
cc_502 N_B_c_564_n N_A_371_74#_c_1091_n 0.00120724f $X=3.827 $Y=1.515 $X2=0
+ $Y2=0
cc_503 N_B_c_565_n N_A_371_74#_c_1091_n 0.00615324f $X=4.295 $Y=1.515 $X2=0
+ $Y2=0
cc_504 N_B_c_566_n N_A_371_74#_c_1091_n 0.0258294f $X=4.21 $Y=1.515 $X2=0 $Y2=0
cc_505 N_B_M1004_g N_A_371_74#_c_1093_n 0.00194376f $X=5.535 $Y=0.925 $X2=0
+ $Y2=0
cc_506 N_B_M1010_g N_A_1116_383#_c_1227_n 0.00796356f $X=5.49 $Y=2.235 $X2=0
+ $Y2=0
cc_507 N_B_M1015_g N_A_1116_383#_c_1227_n 2.17451e-19 $X=6.575 $Y=2.335 $X2=0
+ $Y2=0
cc_508 N_B_M1015_g N_A_1116_383#_c_1221_n 0.0075086f $X=6.575 $Y=2.335 $X2=0
+ $Y2=0
cc_509 N_B_M1010_g N_A_1116_383#_c_1222_n 0.00666049f $X=5.49 $Y=2.235 $X2=0
+ $Y2=0
cc_510 N_B_M1014_g N_A_1116_383#_c_1212_n 0.0066208f $X=6.59 $Y=0.925 $X2=0
+ $Y2=0
cc_511 N_B_M1004_g N_A_1116_383#_c_1213_n 0.00102319f $X=5.535 $Y=0.925 $X2=0
+ $Y2=0
cc_512 N_B_c_574_n N_A_1116_383#_c_1214_n 0.00298078f $X=6.575 $Y=1.78 $X2=0
+ $Y2=0
cc_513 N_B_M1015_g N_A_1116_383#_c_1214_n 0.0209623f $X=6.575 $Y=2.335 $X2=0
+ $Y2=0
cc_514 N_B_M1014_g N_A_1116_383#_c_1214_n 0.00233957f $X=6.59 $Y=0.925 $X2=0
+ $Y2=0
cc_515 N_B_M1014_g N_A_1116_383#_c_1217_n 0.0117925f $X=6.59 $Y=0.925 $X2=0
+ $Y2=0
cc_516 N_B_M1014_g N_A_1116_383#_c_1237_n 2.27589e-19 $X=6.59 $Y=0.925 $X2=0
+ $Y2=0
cc_517 N_B_M1004_g N_A_1116_383#_c_1220_n 0.00483096f $X=5.535 $Y=0.925 $X2=0
+ $Y2=0
cc_518 N_B_M1014_g N_A_1116_383#_c_1220_n 0.00140428f $X=6.59 $Y=0.925 $X2=0
+ $Y2=0
cc_519 N_B_c_561_n N_VGND_c_1328_n 0.00546687f $X=3.855 $Y=1.35 $X2=0 $Y2=0
cc_520 N_B_c_561_n N_VGND_c_1332_n 0.00377304f $X=3.855 $Y=1.35 $X2=0 $Y2=0
cc_521 N_B_c_561_n N_VGND_c_1334_n 0.00505379f $X=3.855 $Y=1.35 $X2=0 $Y2=0
cc_522 N_A_M1020_g N_A_897_54#_M1011_g 0.0269525f $X=7.115 $Y=2.415 $X2=0 $Y2=0
cc_523 N_A_M1017_g N_A_897_54#_M1005_g 0.018076f $X=7.085 $Y=0.925 $X2=0 $Y2=0
cc_524 N_A_M1020_g N_A_897_54#_c_742_n 0.00488111f $X=7.115 $Y=2.415 $X2=0 $Y2=0
cc_525 N_A_M1017_g N_A_897_54#_c_735_n 0.0100072f $X=7.085 $Y=0.925 $X2=0 $Y2=0
cc_526 N_A_M1020_g N_A_897_54#_c_767_n 0.00194944f $X=7.115 $Y=2.415 $X2=0 $Y2=0
cc_527 A N_A_897_54#_c_767_n 0.0178848f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_528 N_A_c_691_n N_A_897_54#_c_767_n 9.43463e-19 $X=7.04 $Y=1.59 $X2=0 $Y2=0
cc_529 N_A_M1020_g N_A_897_54#_c_743_n 0.0146805f $X=7.115 $Y=2.415 $X2=0 $Y2=0
cc_530 N_A_M1017_g N_A_897_54#_c_736_n 0.0108676f $X=7.085 $Y=0.925 $X2=0 $Y2=0
cc_531 A N_A_897_54#_c_736_n 0.0106373f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_532 N_A_c_691_n N_A_897_54#_c_736_n 0.00116518f $X=7.04 $Y=1.59 $X2=0 $Y2=0
cc_533 N_A_M1017_g N_A_897_54#_c_737_n 6.71563e-19 $X=7.085 $Y=0.925 $X2=0 $Y2=0
cc_534 A N_A_897_54#_c_737_n 0.0127015f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_535 N_A_c_691_n N_A_897_54#_c_737_n 0.00301149f $X=7.04 $Y=1.59 $X2=0 $Y2=0
cc_536 N_A_M1020_g N_A_897_54#_c_788_n 0.0107719f $X=7.115 $Y=2.415 $X2=0 $Y2=0
cc_537 A N_A_897_54#_c_788_n 0.00802749f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_538 N_A_M1020_g N_A_897_54#_c_744_n 0.00371028f $X=7.115 $Y=2.415 $X2=0 $Y2=0
cc_539 A N_A_897_54#_c_791_n 0.0221553f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_540 N_A_c_691_n N_A_897_54#_c_791_n 4.17019e-19 $X=7.04 $Y=1.59 $X2=0 $Y2=0
cc_541 A N_A_897_54#_c_739_n 0.0011471f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_542 N_A_c_691_n N_A_897_54#_c_739_n 0.0207694f $X=7.04 $Y=1.59 $X2=0 $Y2=0
cc_543 N_A_M1017_g N_A_897_54#_c_740_n 0.00287145f $X=7.085 $Y=0.925 $X2=0 $Y2=0
cc_544 N_A_M1020_g N_VPWR_c_882_n 0.0044841f $X=7.115 $Y=2.415 $X2=0 $Y2=0
cc_545 N_A_M1020_g N_VPWR_c_885_n 0.00456374f $X=7.115 $Y=2.415 $X2=0 $Y2=0
cc_546 N_A_M1020_g N_VPWR_c_879_n 0.00407483f $X=7.115 $Y=2.415 $X2=0 $Y2=0
cc_547 A N_A_1116_383#_c_1212_n 0.0105608f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_548 N_A_M1020_g N_A_1116_383#_c_1214_n 0.00106063f $X=7.115 $Y=2.415 $X2=0
+ $Y2=0
cc_549 A N_A_1116_383#_c_1214_n 0.0103427f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_550 N_A_M1017_g N_A_1116_383#_c_1217_n 0.00307143f $X=7.085 $Y=0.925 $X2=0
+ $Y2=0
cc_551 A N_A_1116_383#_c_1217_n 0.00974871f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_552 N_A_c_691_n N_A_1116_383#_c_1217_n 0.00481562f $X=7.04 $Y=1.59 $X2=0
+ $Y2=0
cc_553 N_A_M1017_g N_VGND_c_1329_n 0.00317276f $X=7.085 $Y=0.925 $X2=0 $Y2=0
cc_554 N_A_M1017_g N_VGND_c_1332_n 0.00365939f $X=7.085 $Y=0.925 $X2=0 $Y2=0
cc_555 N_A_M1017_g N_VGND_c_1334_n 0.00397505f $X=7.085 $Y=0.925 $X2=0 $Y2=0
cc_556 N_A_897_54#_c_788_n N_VPWR_M1020_d 0.00560843f $X=7.415 $Y=2.035 $X2=0
+ $Y2=0
cc_557 N_A_897_54#_c_744_n N_VPWR_M1020_d 4.15049e-19 $X=7.517 $Y=1.95 $X2=0
+ $Y2=0
cc_558 N_A_897_54#_M1011_g N_VPWR_c_882_n 0.0156702f $X=7.65 $Y=2.415 $X2=0
+ $Y2=0
cc_559 N_A_897_54#_c_742_n N_VPWR_c_882_n 0.0139408f $X=6.76 $Y=2.99 $X2=0 $Y2=0
cc_560 N_A_897_54#_c_788_n N_VPWR_c_882_n 0.0227131f $X=7.415 $Y=2.035 $X2=0
+ $Y2=0
cc_561 N_A_897_54#_c_739_n N_VPWR_c_882_n 4.44487e-19 $X=7.58 $Y=1.59 $X2=0
+ $Y2=0
cc_562 N_A_897_54#_c_742_n N_VPWR_c_885_n 0.147525f $X=6.76 $Y=2.99 $X2=0 $Y2=0
cc_563 N_A_897_54#_c_745_n N_VPWR_c_885_n 0.0213919f $X=4.655 $Y=2.795 $X2=0
+ $Y2=0
cc_564 N_A_897_54#_M1011_g N_VPWR_c_886_n 0.00543803f $X=7.65 $Y=2.415 $X2=0
+ $Y2=0
cc_565 N_A_897_54#_M1011_g N_VPWR_c_879_n 0.00535043f $X=7.65 $Y=2.415 $X2=0
+ $Y2=0
cc_566 N_A_897_54#_c_742_n N_VPWR_c_879_n 0.078121f $X=6.76 $Y=2.99 $X2=0 $Y2=0
cc_567 N_A_897_54#_c_745_n N_VPWR_c_879_n 0.0110564f $X=4.655 $Y=2.795 $X2=0
+ $Y2=0
cc_568 N_A_897_54#_M1009_s N_A_363_394#_c_964_n 0.00699405f $X=4.52 $Y=1.865
+ $X2=0 $Y2=0
cc_569 N_A_897_54#_c_742_n N_A_363_394#_c_964_n 0.0161958f $X=6.76 $Y=2.99 $X2=0
+ $Y2=0
cc_570 N_A_897_54#_c_745_n N_A_363_394#_c_964_n 0.0244309f $X=4.655 $Y=2.795
+ $X2=0 $Y2=0
cc_571 N_A_897_54#_c_734_n N_A_363_394#_c_957_n 0.021871f $X=6.705 $Y=0.34 $X2=0
+ $Y2=0
cc_572 N_A_897_54#_c_735_n N_A_363_394#_c_957_n 0.00753712f $X=6.87 $Y=0.75
+ $X2=0 $Y2=0
cc_573 N_A_897_54#_M1007_s N_A_363_394#_c_959_n 0.0098613f $X=4.485 $Y=0.27
+ $X2=0 $Y2=0
cc_574 N_A_897_54#_c_734_n N_A_363_394#_c_959_n 0.00682298f $X=6.705 $Y=0.34
+ $X2=0 $Y2=0
cc_575 N_A_897_54#_c_738_n N_A_363_394#_c_959_n 0.0267641f $X=4.84 $Y=0.377
+ $X2=0 $Y2=0
cc_576 N_A_897_54#_c_734_n N_A_363_394#_c_960_n 0.0866565f $X=6.705 $Y=0.34
+ $X2=0 $Y2=0
cc_577 N_A_897_54#_M1007_s N_A_371_74#_c_1091_n 0.00228949f $X=4.485 $Y=0.27
+ $X2=0 $Y2=0
cc_578 N_A_897_54#_c_742_n N_A_1116_383#_c_1221_n 0.0481163f $X=6.76 $Y=2.99
+ $X2=0 $Y2=0
cc_579 N_A_897_54#_c_743_n N_A_1116_383#_c_1221_n 0.0140086f $X=6.925 $Y=2.905
+ $X2=0 $Y2=0
cc_580 N_A_897_54#_c_742_n N_A_1116_383#_c_1222_n 0.0256856f $X=6.76 $Y=2.99
+ $X2=0 $Y2=0
cc_581 N_A_897_54#_c_767_n N_A_1116_383#_c_1214_n 0.0134181f $X=6.925 $Y=2.12
+ $X2=0 $Y2=0
cc_582 N_A_897_54#_c_743_n N_A_1116_383#_c_1214_n 0.0328527f $X=6.925 $Y=2.905
+ $X2=0 $Y2=0
cc_583 N_A_897_54#_M1011_g N_A_1116_383#_c_1225_n 7.5409e-19 $X=7.65 $Y=2.415
+ $X2=0 $Y2=0
cc_584 N_A_897_54#_M1005_g N_A_1116_383#_c_1215_n 7.18085e-19 $X=7.665 $Y=0.925
+ $X2=0 $Y2=0
cc_585 N_A_897_54#_c_736_n N_A_1116_383#_c_1216_n 0.00781578f $X=7.415 $Y=1.17
+ $X2=0 $Y2=0
cc_586 N_A_897_54#_M1014_d N_A_1116_383#_c_1217_n 0.00148336f $X=6.665 $Y=0.605
+ $X2=0 $Y2=0
cc_587 N_A_897_54#_M1005_g N_A_1116_383#_c_1217_n 0.00989456f $X=7.665 $Y=0.925
+ $X2=0 $Y2=0
cc_588 N_A_897_54#_c_767_n N_A_1116_383#_c_1217_n 0.00345957f $X=6.925 $Y=2.12
+ $X2=0 $Y2=0
cc_589 N_A_897_54#_c_736_n N_A_1116_383#_c_1217_n 0.0213609f $X=7.415 $Y=1.17
+ $X2=0 $Y2=0
cc_590 N_A_897_54#_c_737_n N_A_1116_383#_c_1217_n 0.0239136f $X=7.035 $Y=1.17
+ $X2=0 $Y2=0
cc_591 N_A_897_54#_c_788_n N_A_1116_383#_c_1217_n 0.00655945f $X=7.415 $Y=2.035
+ $X2=0 $Y2=0
cc_592 N_A_897_54#_c_791_n N_A_1116_383#_c_1217_n 0.0020599f $X=7.58 $Y=1.59
+ $X2=0 $Y2=0
cc_593 N_A_897_54#_c_740_n N_A_1116_383#_c_1217_n 0.0135061f $X=7.54 $Y=1.425
+ $X2=0 $Y2=0
cc_594 N_A_897_54#_c_737_n N_A_1116_383#_c_1237_n 3.64583e-19 $X=7.035 $Y=1.17
+ $X2=0 $Y2=0
cc_595 N_A_897_54#_M1005_g N_A_1116_383#_c_1218_n 0.00116153f $X=7.665 $Y=0.925
+ $X2=0 $Y2=0
cc_596 N_A_897_54#_c_736_n N_A_1116_383#_c_1218_n 0.00133313f $X=7.415 $Y=1.17
+ $X2=0 $Y2=0
cc_597 N_A_897_54#_c_740_n N_A_1116_383#_c_1218_n 0.00132105f $X=7.54 $Y=1.425
+ $X2=0 $Y2=0
cc_598 N_A_897_54#_M1011_g N_A_1116_383#_c_1219_n 0.0103744f $X=7.65 $Y=2.415
+ $X2=0 $Y2=0
cc_599 N_A_897_54#_M1005_g N_A_1116_383#_c_1219_n 0.00324328f $X=7.665 $Y=0.925
+ $X2=0 $Y2=0
cc_600 N_A_897_54#_c_788_n N_A_1116_383#_c_1219_n 0.0114115f $X=7.415 $Y=2.035
+ $X2=0 $Y2=0
cc_601 N_A_897_54#_c_744_n N_A_1116_383#_c_1219_n 0.0120839f $X=7.517 $Y=1.95
+ $X2=0 $Y2=0
cc_602 N_A_897_54#_c_791_n N_A_1116_383#_c_1219_n 0.024951f $X=7.58 $Y=1.59
+ $X2=0 $Y2=0
cc_603 N_A_897_54#_c_739_n N_A_1116_383#_c_1219_n 0.00820404f $X=7.58 $Y=1.59
+ $X2=0 $Y2=0
cc_604 N_A_897_54#_c_740_n N_A_1116_383#_c_1219_n 0.00894219f $X=7.54 $Y=1.425
+ $X2=0 $Y2=0
cc_605 N_A_897_54#_c_737_n N_A_1116_383#_c_1220_n 3.92581e-19 $X=7.035 $Y=1.17
+ $X2=0 $Y2=0
cc_606 N_A_897_54#_c_736_n N_VGND_M1017_d 0.00401601f $X=7.415 $Y=1.17 $X2=0
+ $Y2=0
cc_607 N_A_897_54#_M1005_g N_VGND_c_1329_n 0.0112617f $X=7.665 $Y=0.925 $X2=0
+ $Y2=0
cc_608 N_A_897_54#_c_734_n N_VGND_c_1329_n 0.0152756f $X=6.705 $Y=0.34 $X2=0
+ $Y2=0
cc_609 N_A_897_54#_c_735_n N_VGND_c_1329_n 0.0262473f $X=6.87 $Y=0.75 $X2=0
+ $Y2=0
cc_610 N_A_897_54#_c_736_n N_VGND_c_1329_n 0.0267054f $X=7.415 $Y=1.17 $X2=0
+ $Y2=0
cc_611 N_A_897_54#_c_739_n N_VGND_c_1329_n 5.78471e-19 $X=7.58 $Y=1.59 $X2=0
+ $Y2=0
cc_612 N_A_897_54#_c_734_n N_VGND_c_1332_n 0.0236566f $X=6.705 $Y=0.34 $X2=0
+ $Y2=0
cc_613 N_A_897_54#_c_738_n N_VGND_c_1332_n 0.141098f $X=4.84 $Y=0.377 $X2=0
+ $Y2=0
cc_614 N_A_897_54#_M1005_g N_VGND_c_1333_n 0.00354091f $X=7.665 $Y=0.925 $X2=0
+ $Y2=0
cc_615 N_A_897_54#_M1005_g N_VGND_c_1334_n 0.00398995f $X=7.665 $Y=0.925 $X2=0
+ $Y2=0
cc_616 N_A_897_54#_c_734_n N_VGND_c_1334_n 0.0128296f $X=6.705 $Y=0.34 $X2=0
+ $Y2=0
cc_617 N_A_897_54#_c_738_n N_VGND_c_1334_n 0.0784557f $X=4.84 $Y=0.377 $X2=0
+ $Y2=0
cc_618 N_X_c_862_n N_VPWR_c_880_n 0.0224694f $X=0.27 $Y=2.005 $X2=0 $Y2=0
cc_619 N_X_c_862_n N_VPWR_c_883_n 0.0119584f $X=0.27 $Y=2.005 $X2=0 $Y2=0
cc_620 N_X_c_862_n N_VPWR_c_879_n 0.00989813f $X=0.27 $Y=2.005 $X2=0 $Y2=0
cc_621 X N_VGND_c_1327_n 0.00381405f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_622 X N_VGND_c_1330_n 0.0116428f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_623 X N_VGND_c_1334_n 0.0124588f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_624 N_VPWR_c_879_n N_A_363_394#_c_962_n 0.0257339f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_625 N_VPWR_M1002_s N_A_363_394#_c_955_n 0.00938121f $X=3.425 $Y=1.84 $X2=0
+ $Y2=0
cc_626 N_VPWR_M1002_s N_A_363_394#_c_964_n 0.00953832f $X=3.425 $Y=1.84 $X2=0
+ $Y2=0
cc_627 N_VPWR_c_881_n N_A_363_394#_c_964_n 0.0149016f $X=3.56 $Y=2.875 $X2=0
+ $Y2=0
cc_628 N_VPWR_c_879_n N_A_363_394#_c_964_n 0.0268314f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_629 N_VPWR_M1002_s N_A_363_394#_c_966_n 0.00201704f $X=3.425 $Y=1.84 $X2=0
+ $Y2=0
cc_630 N_VPWR_c_881_n N_A_363_394#_c_966_n 0.0113807f $X=3.56 $Y=2.875 $X2=0
+ $Y2=0
cc_631 N_VPWR_c_879_n N_A_363_394#_c_966_n 0.00217269f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_632 N_VPWR_c_882_n N_A_1116_383#_c_1225_n 0.0215931f $X=7.425 $Y=2.375 $X2=0
+ $Y2=0
cc_633 N_VPWR_c_886_n N_A_1116_383#_c_1225_n 0.0105094f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_634 N_VPWR_c_879_n N_A_1116_383#_c_1225_n 0.010131f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_635 N_A_363_394#_c_957_n N_A_371_74#_M1007_d 0.0031922f $X=6.255 $Y=0.68
+ $X2=0 $Y2=0
cc_636 N_A_363_394#_c_960_n N_A_371_74#_M1007_d 0.00192105f $X=5.18 $Y=0.717
+ $X2=0 $Y2=0
cc_637 N_A_363_394#_c_962_n N_A_371_74#_M1019_d 0.00740053f $X=3.355 $Y=2.455
+ $X2=0 $Y2=0
cc_638 N_A_363_394#_c_955_n N_A_371_74#_c_1087_n 0.0133454f $X=3.44 $Y=2.37
+ $X2=0 $Y2=0
cc_639 N_A_363_394#_c_956_n N_A_371_74#_c_1087_n 0.0274074f $X=3.525 $Y=0.755
+ $X2=0 $Y2=0
cc_640 N_A_363_394#_c_955_n N_A_371_74#_c_1088_n 0.0539191f $X=3.44 $Y=2.37
+ $X2=0 $Y2=0
cc_641 N_A_363_394#_c_965_n N_A_371_74#_c_1134_n 0.00259034f $X=5.18 $Y=2.02
+ $X2=0 $Y2=0
cc_642 N_A_363_394#_c_957_n N_A_371_74#_c_1134_n 0.0066624f $X=6.255 $Y=0.68
+ $X2=0 $Y2=0
cc_643 N_A_363_394#_c_960_n N_A_371_74#_c_1134_n 0.00697655f $X=5.18 $Y=0.717
+ $X2=0 $Y2=0
cc_644 N_A_363_394#_c_957_n N_A_371_74#_c_1089_n 0.00850447f $X=6.255 $Y=0.68
+ $X2=0 $Y2=0
cc_645 N_A_363_394#_c_965_n N_A_371_74#_c_1148_n 0.00647566f $X=5.18 $Y=2.02
+ $X2=0 $Y2=0
cc_646 N_A_363_394#_c_962_n N_A_371_74#_c_1098_n 0.020055f $X=3.355 $Y=2.455
+ $X2=0 $Y2=0
cc_647 N_A_363_394#_c_955_n N_A_371_74#_c_1098_n 0.0133978f $X=3.44 $Y=2.37
+ $X2=0 $Y2=0
cc_648 N_A_363_394#_c_955_n N_A_371_74#_c_1091_n 0.0257254f $X=3.44 $Y=2.37
+ $X2=0 $Y2=0
cc_649 N_A_363_394#_c_956_n N_A_371_74#_c_1091_n 0.0099531f $X=3.525 $Y=0.755
+ $X2=0 $Y2=0
cc_650 N_A_363_394#_c_965_n N_A_371_74#_c_1091_n 0.00535596f $X=5.18 $Y=2.02
+ $X2=0 $Y2=0
cc_651 N_A_363_394#_c_957_n N_A_371_74#_c_1091_n 2.92758e-19 $X=6.255 $Y=0.68
+ $X2=0 $Y2=0
cc_652 N_A_363_394#_c_959_n N_A_371_74#_c_1091_n 0.019754f $X=5.01 $Y=0.717
+ $X2=0 $Y2=0
cc_653 N_A_363_394#_c_957_n N_A_371_74#_c_1093_n 0.0034939f $X=6.255 $Y=0.68
+ $X2=0 $Y2=0
cc_654 N_A_363_394#_c_957_n N_A_1116_383#_M1004_d 0.00548002f $X=6.255 $Y=0.68
+ $X2=-0.19 $Y2=-0.245
cc_655 N_A_363_394#_c_964_n N_A_1116_383#_c_1227_n 0.010696f $X=5.015 $Y=2.455
+ $X2=0 $Y2=0
cc_656 N_A_363_394#_c_965_n N_A_1116_383#_c_1227_n 0.0135225f $X=5.18 $Y=2.02
+ $X2=0 $Y2=0
cc_657 N_A_363_394#_c_964_n N_A_1116_383#_c_1222_n 5.43654e-19 $X=5.015 $Y=2.455
+ $X2=0 $Y2=0
cc_658 N_A_363_394#_c_957_n N_A_1116_383#_c_1212_n 0.00171574f $X=6.255 $Y=0.68
+ $X2=0 $Y2=0
cc_659 N_A_363_394#_c_958_n N_A_1116_383#_c_1212_n 0.0124099f $X=6.375 $Y=1.045
+ $X2=0 $Y2=0
cc_660 N_A_363_394#_M1021_d N_A_1116_383#_c_1217_n 0.00290016f $X=6.17 $Y=0.825
+ $X2=0 $Y2=0
cc_661 N_A_363_394#_c_957_n N_A_1116_383#_c_1217_n 0.00236222f $X=6.255 $Y=0.68
+ $X2=0 $Y2=0
cc_662 N_A_363_394#_c_958_n N_A_1116_383#_c_1217_n 0.0088961f $X=6.375 $Y=1.045
+ $X2=0 $Y2=0
cc_663 N_A_363_394#_c_957_n N_A_1116_383#_c_1237_n 0.00226222f $X=6.255 $Y=0.68
+ $X2=0 $Y2=0
cc_664 N_A_363_394#_c_958_n N_A_1116_383#_c_1237_n 8.11031e-19 $X=6.375 $Y=1.045
+ $X2=0 $Y2=0
cc_665 N_A_363_394#_c_957_n N_A_1116_383#_c_1220_n 0.0214988f $X=6.255 $Y=0.68
+ $X2=0 $Y2=0
cc_666 N_A_363_394#_c_958_n N_A_1116_383#_c_1220_n 0.0205989f $X=6.375 $Y=1.045
+ $X2=0 $Y2=0
cc_667 N_A_363_394#_c_955_n N_VGND_M1001_s 0.00497246f $X=3.44 $Y=2.37 $X2=0
+ $Y2=0
cc_668 N_A_363_394#_c_956_n N_VGND_M1001_s 0.00490689f $X=3.525 $Y=0.755 $X2=0
+ $Y2=0
cc_669 N_A_363_394#_c_959_n N_VGND_M1001_s 0.00590399f $X=5.01 $Y=0.717 $X2=0
+ $Y2=0
cc_670 N_A_363_394#_c_956_n N_VGND_c_1328_n 0.0211907f $X=3.525 $Y=0.755 $X2=0
+ $Y2=0
cc_671 N_A_363_394#_c_959_n N_VGND_c_1328_n 0.015267f $X=5.01 $Y=0.717 $X2=0
+ $Y2=0
cc_672 N_A_363_394#_c_956_n N_VGND_c_1331_n 0.0187385f $X=3.525 $Y=0.755 $X2=0
+ $Y2=0
cc_673 N_A_363_394#_c_959_n N_VGND_c_1332_n 0.011182f $X=5.01 $Y=0.717 $X2=0
+ $Y2=0
cc_674 N_A_363_394#_c_956_n N_VGND_c_1334_n 0.0194089f $X=3.525 $Y=0.755 $X2=0
+ $Y2=0
cc_675 N_A_363_394#_c_959_n N_VGND_c_1334_n 0.022365f $X=5.01 $Y=0.717 $X2=0
+ $Y2=0
cc_676 N_A_371_74#_c_1093_n N_A_1116_383#_M1004_d 9.13166e-19 $X=5.52 $Y=1.295
+ $X2=-0.19 $Y2=-0.245
cc_677 N_A_371_74#_c_1097_n N_A_1116_383#_M1010_d 0.00165831f $X=6.08 $Y=1.85
+ $X2=0 $Y2=0
cc_678 N_A_371_74#_c_1097_n N_A_1116_383#_c_1227_n 0.0147664f $X=6.08 $Y=1.85
+ $X2=0 $Y2=0
cc_679 N_A_371_74#_c_1148_n N_A_1116_383#_c_1227_n 0.00239886f $X=5.605 $Y=1.85
+ $X2=0 $Y2=0
cc_680 N_A_371_74#_M1012_d N_A_1116_383#_c_1221_n 0.00983165f $X=6.03 $Y=1.915
+ $X2=0 $Y2=0
cc_681 N_A_371_74#_c_1097_n N_A_1116_383#_c_1221_n 0.0041687f $X=6.08 $Y=1.85
+ $X2=0 $Y2=0
cc_682 N_A_371_74#_c_1166_n N_A_1116_383#_c_1221_n 0.0134755f $X=6.165 $Y=2.195
+ $X2=0 $Y2=0
cc_683 N_A_371_74#_c_1097_n N_A_1116_383#_c_1212_n 0.013011f $X=6.08 $Y=1.85
+ $X2=0 $Y2=0
cc_684 N_A_371_74#_c_1090_n N_A_1116_383#_c_1213_n 0.0137161f $X=5.52 $Y=1.765
+ $X2=0 $Y2=0
cc_685 N_A_371_74#_c_1097_n N_A_1116_383#_c_1213_n 0.0237352f $X=6.08 $Y=1.85
+ $X2=0 $Y2=0
cc_686 N_A_371_74#_M1012_d N_A_1116_383#_c_1214_n 0.00672686f $X=6.03 $Y=1.915
+ $X2=0 $Y2=0
cc_687 N_A_371_74#_c_1097_n N_A_1116_383#_c_1214_n 0.014294f $X=6.08 $Y=1.85
+ $X2=0 $Y2=0
cc_688 N_A_371_74#_c_1166_n N_A_1116_383#_c_1214_n 0.0333746f $X=6.165 $Y=2.195
+ $X2=0 $Y2=0
cc_689 N_A_371_74#_c_1089_n N_A_1116_383#_c_1237_n 4.22568e-19 $X=5.52 $Y=1.41
+ $X2=0 $Y2=0
cc_690 N_A_371_74#_c_1097_n N_A_1116_383#_c_1237_n 0.00122034f $X=6.08 $Y=1.85
+ $X2=0 $Y2=0
cc_691 N_A_371_74#_c_1093_n N_A_1116_383#_c_1237_n 0.0211316f $X=5.52 $Y=1.295
+ $X2=0 $Y2=0
cc_692 N_A_371_74#_c_1089_n N_A_1116_383#_c_1220_n 0.0237269f $X=5.52 $Y=1.41
+ $X2=0 $Y2=0
cc_693 N_A_371_74#_c_1090_n N_A_1116_383#_c_1220_n 0.00105161f $X=5.52 $Y=1.765
+ $X2=0 $Y2=0
cc_694 N_A_371_74#_c_1093_n N_A_1116_383#_c_1220_n 0.00186944f $X=5.52 $Y=1.295
+ $X2=0 $Y2=0
cc_695 N_A_371_74#_c_1091_n N_VGND_M1001_s 0.00261715f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_696 N_A_1116_383#_c_1215_n N_VGND_c_1329_n 0.0129676f $X=7.88 $Y=0.75 $X2=0
+ $Y2=0
cc_697 N_A_1116_383#_c_1217_n N_VGND_c_1329_n 0.00251679f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_698 N_A_1116_383#_c_1215_n N_VGND_c_1333_n 0.00626724f $X=7.88 $Y=0.75 $X2=0
+ $Y2=0
cc_699 N_A_1116_383#_c_1215_n N_VGND_c_1334_n 0.00875025f $X=7.88 $Y=0.75 $X2=0
+ $Y2=0

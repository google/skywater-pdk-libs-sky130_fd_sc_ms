* File: sky130_fd_sc_ms__a41o_2.spice
* Created: Wed Sep  2 11:56:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a41o_2.pex.spice"
.subckt sky130_fd_sc_ms__a41o_2  VNB VPB A4 A3 A2 A1 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* VPB	VPB
* VNB	VNB
MM1005 A_121_74# N_A4_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.2 SB=75004
+ A=0.111 P=1.78 MULT=1
MM1004 A_199_74# N_A3_M1004_g A_121_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.0888 PD=1.16 PS=0.98 NRD=25.128 NRS=10.536 M=1 R=4.93333 SA=75000.6
+ SB=75003.6 A=0.111 P=1.78 MULT=1
MM1006 A_313_74# N_A2_M1006_g A_199_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1813
+ AS=0.1554 PD=1.23 PS=1.16 NRD=30.804 NRS=25.128 M=1 R=4.93333 SA=75001.2
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1007 N_A_441_74#_M1007_d N_A1_M1007_g A_313_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.1813 PD=1.13 PS=1.23 NRD=8.1 NRS=30.804 M=1 R=4.93333
+ SA=75001.8 SB=75002.4 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_B1_M1003_g N_A_441_74#_M1007_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1591 AS=0.1443 PD=1.17 PS=1.13 NRD=11.34 NRS=9.72 M=1 R=4.93333
+ SA=75002.4 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1009 N_X_M1009_d N_A_441_74#_M1009_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1517 AS=0.1591 PD=1.15 PS=1.17 NRD=13.776 NRS=12.972 M=1 R=4.93333
+ SA=75002.9 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1012 N_X_M1009_d N_A_441_74#_M1012_g N_VGND_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1517 AS=0.5772 PD=1.15 PS=3.04 NRD=7.296 NRS=4.044 M=1 R=4.93333
+ SA=75003.5 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1002 N_VPWR_M1002_d N_A4_M1002_g N_A_27_392#_M1002_s VPB PSHORT L=0.18 W=1
+ AD=0.185 AS=0.28 PD=1.37 PS=2.56 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90002.4 A=0.18 P=2.36 MULT=1
MM1008 N_A_27_392#_M1008_d N_A3_M1008_g N_VPWR_M1002_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.185 PD=1.27 PS=1.37 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90000.7
+ SB=90001.9 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1010_d N_A2_M1010_g N_A_27_392#_M1008_d VPB PSHORT L=0.18 W=1
+ AD=0.275 AS=0.135 PD=1.55 PS=1.27 NRD=26.5753 NRS=0 M=1 R=5.55556 SA=90001.2
+ SB=90001.4 A=0.18 P=2.36 MULT=1
MM1013 N_A_27_392#_M1013_d N_A1_M1013_g N_VPWR_M1010_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.275 PD=1.27 PS=1.55 NRD=0 NRS=26.5753 M=1 R=5.55556 SA=90001.9
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1001 N_A_441_74#_M1001_d N_B1_M1001_g N_A_27_392#_M1013_d VPB PSHORT L=0.18
+ W=1 AD=0.33 AS=0.135 PD=2.66 PS=1.27 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90002.4
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_A_441_74#_M1000_g N_X_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3696 AS=0.1512 PD=2.9 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1011 N_VPWR_M1011_d N_A_441_74#_M1011_g N_X_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3696 AS=0.1512 PD=2.9 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90000.7
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_ms__a41o_2.pxi.spice"
*
.ends
*
*

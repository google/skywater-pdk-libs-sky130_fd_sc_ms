* File: sky130_fd_sc_ms__a311oi_4.pxi.spice
* Created: Fri Aug 28 17:06:28 2020
* 
x_PM_SKY130_FD_SC_MS__A311OI_4%A3 N_A3_M1028_g N_A3_M1010_g N_A3_M1029_g
+ N_A3_M1023_g N_A3_M1031_g N_A3_M1026_g N_A3_M1027_g N_A3_M1034_g A3 A3 A3
+ N_A3_c_163_n N_A3_c_158_n PM_SKY130_FD_SC_MS__A311OI_4%A3
x_PM_SKY130_FD_SC_MS__A311OI_4%A2 N_A2_M1002_g N_A2_M1000_g N_A2_M1003_g
+ N_A2_M1005_g N_A2_M1007_g N_A2_M1008_g N_A2_M1018_g N_A2_M1012_g A2 A2 A2 A2
+ N_A2_c_232_n PM_SKY130_FD_SC_MS__A311OI_4%A2
x_PM_SKY130_FD_SC_MS__A311OI_4%A1 N_A1_M1016_g N_A1_c_307_n N_A1_c_308_n
+ N_A1_M1020_g N_A1_M1004_g N_A1_M1022_g N_A1_M1015_g N_A1_M1030_g N_A1_M1019_g
+ N_A1_M1025_g A1 A1 N_A1_c_314_n PM_SKY130_FD_SC_MS__A311OI_4%A1
x_PM_SKY130_FD_SC_MS__A311OI_4%B1 N_B1_M1001_g N_B1_M1017_g N_B1_M1006_g
+ N_B1_M1032_g N_B1_M1024_g N_B1_M1035_g B1 B1 N_B1_c_396_n N_B1_c_397_n
+ PM_SKY130_FD_SC_MS__A311OI_4%B1
x_PM_SKY130_FD_SC_MS__A311OI_4%C1 N_C1_c_469_n N_C1_M1011_g N_C1_M1009_g
+ N_C1_c_471_n N_C1_M1033_g N_C1_M1013_g N_C1_M1014_g N_C1_c_474_n N_C1_M1021_g
+ C1 C1 N_C1_c_476_n N_C1_c_477_n N_C1_c_478_n C1
+ PM_SKY130_FD_SC_MS__A311OI_4%C1
x_PM_SKY130_FD_SC_MS__A311OI_4%VPWR N_VPWR_M1028_s N_VPWR_M1029_s N_VPWR_M1034_s
+ N_VPWR_M1005_s N_VPWR_M1012_s N_VPWR_M1020_s N_VPWR_M1030_s N_VPWR_c_546_n
+ N_VPWR_c_547_n N_VPWR_c_548_n N_VPWR_c_549_n N_VPWR_c_550_n N_VPWR_c_551_n
+ N_VPWR_c_552_n N_VPWR_c_553_n N_VPWR_c_554_n N_VPWR_c_555_n N_VPWR_c_556_n
+ N_VPWR_c_557_n N_VPWR_c_558_n N_VPWR_c_559_n N_VPWR_c_560_n N_VPWR_c_561_n
+ N_VPWR_c_562_n VPWR N_VPWR_c_563_n N_VPWR_c_564_n N_VPWR_c_545_n
+ N_VPWR_c_566_n N_VPWR_c_567_n PM_SKY130_FD_SC_MS__A311OI_4%VPWR
x_PM_SKY130_FD_SC_MS__A311OI_4%A_117_368# N_A_117_368#_M1028_d
+ N_A_117_368#_M1031_d N_A_117_368#_M1000_d N_A_117_368#_M1008_d
+ N_A_117_368#_M1016_d N_A_117_368#_M1022_d N_A_117_368#_M1001_d
+ N_A_117_368#_M1032_d N_A_117_368#_c_697_n N_A_117_368#_c_686_n
+ N_A_117_368#_c_701_n N_A_117_368#_c_687_n N_A_117_368#_c_705_n
+ N_A_117_368#_c_688_n N_A_117_368#_c_711_n N_A_117_368#_c_689_n
+ N_A_117_368#_c_715_n N_A_117_368#_c_690_n N_A_117_368#_c_724_n
+ N_A_117_368#_c_691_n N_A_117_368#_c_692_n N_A_117_368#_c_789_p
+ N_A_117_368#_c_693_n N_A_117_368#_c_694_n N_A_117_368#_c_792_p
+ N_A_117_368#_c_707_n N_A_117_368#_c_717_n N_A_117_368#_c_719_n
+ N_A_117_368#_c_695_n N_A_117_368#_c_736_n N_A_117_368#_c_696_n
+ PM_SKY130_FD_SC_MS__A311OI_4%A_117_368#
x_PM_SKY130_FD_SC_MS__A311OI_4%A_1213_368# N_A_1213_368#_M1001_s
+ N_A_1213_368#_M1006_s N_A_1213_368#_M1035_s N_A_1213_368#_M1013_s
+ N_A_1213_368#_M1021_s N_A_1213_368#_c_794_n N_A_1213_368#_c_795_n
+ N_A_1213_368#_c_796_n N_A_1213_368#_c_811_n N_A_1213_368#_c_797_n
+ N_A_1213_368#_c_798_n N_A_1213_368#_c_799_n N_A_1213_368#_c_828_n
+ N_A_1213_368#_c_800_n N_A_1213_368#_c_801_n N_A_1213_368#_c_802_n
+ N_A_1213_368#_c_803_n N_A_1213_368#_c_804_n
+ PM_SKY130_FD_SC_MS__A311OI_4%A_1213_368#
x_PM_SKY130_FD_SC_MS__A311OI_4%Y N_Y_M1004_d N_Y_M1015_d N_Y_M1025_d N_Y_M1024_s
+ N_Y_M1033_d N_Y_M1009_d N_Y_M1014_d N_Y_c_874_n N_Y_c_875_n N_Y_c_897_n
+ N_Y_c_876_n N_Y_c_933_n N_Y_c_882_n N_Y_c_883_n N_Y_c_877_n N_Y_c_937_n
+ N_Y_c_878_n N_Y_c_879_n N_Y_c_905_n N_Y_c_885_n Y Y Y N_Y_c_923_n Y
+ N_Y_c_881_n PM_SKY130_FD_SC_MS__A311OI_4%Y
x_PM_SKY130_FD_SC_MS__A311OI_4%A_34_74# N_A_34_74#_M1010_s N_A_34_74#_M1023_s
+ N_A_34_74#_M1027_s N_A_34_74#_M1003_s N_A_34_74#_M1018_s N_A_34_74#_c_965_n
+ N_A_34_74#_c_966_n N_A_34_74#_c_967_n N_A_34_74#_c_968_n N_A_34_74#_c_969_n
+ N_A_34_74#_c_970_n N_A_34_74#_c_971_n N_A_34_74#_c_972_n N_A_34_74#_c_973_n
+ N_A_34_74#_c_974_n N_A_34_74#_c_975_n N_A_34_74#_c_976_n
+ PM_SKY130_FD_SC_MS__A311OI_4%A_34_74#
x_PM_SKY130_FD_SC_MS__A311OI_4%VGND N_VGND_M1010_d N_VGND_M1026_d N_VGND_M1017_d
+ N_VGND_M1011_s N_VGND_c_1039_n N_VGND_c_1040_n N_VGND_c_1041_n VGND
+ N_VGND_c_1042_n N_VGND_c_1043_n N_VGND_c_1044_n N_VGND_c_1045_n
+ N_VGND_c_1046_n N_VGND_c_1047_n N_VGND_c_1048_n N_VGND_c_1049_n
+ N_VGND_c_1050_n N_VGND_c_1051_n PM_SKY130_FD_SC_MS__A311OI_4%VGND
x_PM_SKY130_FD_SC_MS__A311OI_4%A_465_74# N_A_465_74#_M1002_d N_A_465_74#_M1007_d
+ N_A_465_74#_M1004_s N_A_465_74#_M1019_s N_A_465_74#_c_1128_n
+ N_A_465_74#_c_1129_n N_A_465_74#_c_1130_n N_A_465_74#_c_1131_n
+ N_A_465_74#_c_1132_n PM_SKY130_FD_SC_MS__A311OI_4%A_465_74#
cc_1 VNB N_A3_M1010_g 0.0318708f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_2 VNB N_A3_M1023_g 0.0230578f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_3 VNB N_A3_M1026_g 0.0224931f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=0.74
cc_4 VNB N_A3_M1027_g 0.0229868f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=0.74
cc_5 VNB N_A3_c_158_n 0.0829948f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.515
cc_6 VNB N_A2_M1002_g 0.0236065f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_7 VNB N_A2_M1003_g 0.0230075f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_8 VNB N_A2_M1007_g 0.0230075f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.4
cc_9 VNB N_A2_M1018_g 0.0325857f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=0.74
cc_10 VNB A2 0.00306242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A2_c_232_n 0.07883f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.515
cc_12 VNB N_A1_c_307_n 0.0148673f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.35
cc_13 VNB N_A1_c_308_n 0.0149665f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_14 VNB N_A1_M1004_g 0.0337355f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.35
cc_15 VNB N_A1_M1015_g 0.0234256f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=1.35
cc_16 VNB N_A1_M1019_g 0.0234256f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.68
cc_17 VNB N_A1_M1025_g 0.0240737f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_18 VNB A1 0.0109081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_314_n 0.0721086f $X=-0.19 $Y=-0.245 $X2=1.71 $Y2=1.515
cc_20 VNB N_B1_M1001_g 4.86581e-19 $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_21 VNB N_B1_M1017_g 0.0261425f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_22 VNB N_B1_M1006_g 4.7877e-19 $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=2.4
cc_23 VNB N_B1_M1032_g 4.78866e-19 $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_24 VNB N_B1_M1024_g 0.0259064f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.4
cc_25 VNB N_B1_M1035_g 4.95336e-19 $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=0.74
cc_26 VNB B1 0.00573161f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=0.74
cc_27 VNB N_B1_c_396_n 0.100477f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_28 VNB N_B1_c_397_n 0.00679545f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.515
cc_29 VNB N_C1_c_469_n 0.0168861f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.68
cc_30 VNB N_C1_M1009_g 0.00598807f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=0.74
cc_31 VNB N_C1_c_471_n 0.0210077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_C1_M1013_g 0.00579577f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.35
cc_33 VNB N_C1_M1014_g 0.0057674f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=1.68
cc_34 VNB N_C1_c_474_n 0.0422752f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.4
cc_35 VNB N_C1_M1021_g 0.0158274f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=0.74
cc_36 VNB N_C1_c_476_n 0.0046005f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_37 VNB N_C1_c_477_n 0.0705361f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.515
cc_38 VNB N_C1_c_478_n 0.00623501f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.515
cc_39 VNB N_VPWR_c_545_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Y_c_874_n 0.00842476f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=0.74
cc_41 VNB N_Y_c_875_n 0.00206055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_Y_c_876_n 0.00206768f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_43 VNB N_Y_c_877_n 0.0137919f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.515
cc_44 VNB N_Y_c_878_n 0.00967636f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.515
cc_45 VNB N_Y_c_879_n 0.00828779f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.565
cc_46 VNB Y 0.0381136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_Y_c_881_n 0.0357019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_34_74#_c_965_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.4
cc_49 VNB N_A_34_74#_c_966_n 0.00273425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_34_74#_c_967_n 0.0126474f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=1.35
cc_51 VNB N_A_34_74#_c_968_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_34_74#_c_969_n 0.0036153f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=0.74
cc_53 VNB N_A_34_74#_c_970_n 0.00178301f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_54 VNB N_A_34_74#_c_971_n 0.00226168f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_55 VNB N_A_34_74#_c_972_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_34_74#_c_973_n 0.0045734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_34_74#_c_974_n 0.00275936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_34_74#_c_975_n 0.00228886f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.515
cc_59 VNB N_A_34_74#_c_976_n 0.0156582f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.515
cc_60 VNB N_VGND_c_1039_n 0.00481913f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=0.74
cc_61 VNB N_VGND_c_1040_n 0.00334323f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.4
cc_62 VNB N_VGND_c_1041_n 0.00332936f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=0.74
cc_63 VNB N_VGND_c_1042_n 0.0185047f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=0.74
cc_64 VNB N_VGND_c_1043_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1044_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.515
cc_66 VNB N_VGND_c_1045_n 0.0418428f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.565
cc_67 VNB N_VGND_c_1046_n 0.525006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1047_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_69 VNB N_VGND_c_1048_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1049_n 0.12018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1050_n 0.0364641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1051_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_465_74#_c_1128_n 0.00199246f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=0.74
cc_74 VNB N_A_465_74#_c_1129_n 0.00310413f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=1.35
cc_75 VNB N_A_465_74#_c_1130_n 0.00161093f $X=-0.19 $Y=-0.245 $X2=1.82 $Y2=0.74
cc_76 VNB N_A_465_74#_c_1131_n 0.002374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_465_74#_c_1132_n 0.0338474f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.68
cc_78 VPB N_A3_M1028_g 0.0260117f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_79 VPB N_A3_M1029_g 0.0198948f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_80 VPB N_A3_M1031_g 0.0198928f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_81 VPB N_A3_M1034_g 0.020575f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_82 VPB N_A3_c_163_n 0.00755402f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.515
cc_83 VPB N_A3_c_158_n 0.0124572f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.515
cc_84 VPB N_A2_M1000_g 0.0200213f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=0.74
cc_85 VPB N_A2_M1005_g 0.0198928f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=0.74
cc_86 VPB N_A2_M1008_g 0.0198928f $X=-0.19 $Y=1.66 $X2=1.39 $Y2=0.74
cc_87 VPB N_A2_M1012_g 0.0206032f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_88 VPB A2 0.00976107f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A2_c_232_n 0.0116067f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.515
cc_90 VPB N_A1_M1016_g 0.0209894f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_91 VPB N_A1_c_307_n 0.00254267f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=1.35
cc_92 VPB N_A1_c_308_n 7.71944e-19 $X=-0.19 $Y=1.66 $X2=0.53 $Y2=0.74
cc_93 VPB N_A1_M1020_g 0.0202975f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.68
cc_94 VPB N_A1_M1022_g 0.0204946f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.68
cc_95 VPB N_A1_M1030_g 0.0253603f $X=-0.19 $Y=1.66 $X2=1.82 $Y2=1.35
cc_96 VPB A1 0.0118438f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A1_c_314_n 0.0242035f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.515
cc_98 VPB N_B1_M1001_g 0.0260074f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_99 VPB N_B1_M1006_g 0.0213675f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_100 VPB N_B1_M1032_g 0.0213688f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=0.74
cc_101 VPB N_B1_M1035_g 0.021786f $X=-0.19 $Y=1.66 $X2=1.39 $Y2=0.74
cc_102 VPB N_C1_M1009_g 0.0217605f $X=-0.19 $Y=1.66 $X2=0.53 $Y2=0.74
cc_103 VPB N_C1_M1013_g 0.0205117f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.35
cc_104 VPB N_C1_M1014_g 0.0204961f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.68
cc_105 VPB N_C1_M1021_g 0.0288769f $X=-0.19 $Y=1.66 $X2=1.39 $Y2=0.74
cc_106 VPB N_VPWR_c_546_n 0.0103331f $X=-0.19 $Y=1.66 $X2=1.39 $Y2=0.74
cc_107 VPB N_VPWR_c_547_n 0.0598916f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_548_n 0.00271781f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_109 VPB N_VPWR_c_549_n 0.00261791f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_110 VPB N_VPWR_c_550_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_551_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.515
cc_112 VPB N_VPWR_c_552_n 0.00417807f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.515
cc_113 VPB N_VPWR_c_553_n 0.0185253f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.515
cc_114 VPB N_VPWR_c_554_n 0.0121609f $X=-0.19 $Y=1.66 $X2=1.82 $Y2=1.515
cc_115 VPB N_VPWR_c_555_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.565
cc_116 VPB N_VPWR_c_556_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_557_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_558_n 0.00601644f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_119 VPB N_VPWR_c_559_n 0.0164465f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.565
cc_120 VPB N_VPWR_c_560_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_561_n 0.0164465f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.565
cc_122 VPB N_VPWR_c_562_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_563_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_564_n 0.0991002f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_545_n 0.104411f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_566_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_567_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_117_368#_c_686_n 0.00202354f $X=-0.19 $Y=1.66 $X2=1.82 $Y2=0.74
cc_129 VPB N_A_117_368#_c_687_n 0.00179594f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_130 VPB N_A_117_368#_c_688_n 0.00179594f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.515
cc_131 VPB N_A_117_368#_c_689_n 0.00179594f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.515
cc_132 VPB N_A_117_368#_c_690_n 0.00179594f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.515
cc_133 VPB N_A_117_368#_c_691_n 0.00202354f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_134 VPB N_A_117_368#_c_692_n 0.0107168f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_135 VPB N_A_117_368#_c_693_n 0.00310387f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_117_368#_c_694_n 0.00199716f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_117_368#_c_695_n 0.00460758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_117_368#_c_696_n 0.00747115f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_1213_368#_c_794_n 0.00552465f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_140 VPB N_A_1213_368#_c_795_n 0.00192243f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_1213_368#_c_796_n 0.00405878f $X=-0.19 $Y=1.66 $X2=1.39 $Y2=1.35
cc_142 VPB N_A_1213_368#_c_797_n 0.00192243f $X=-0.19 $Y=1.66 $X2=1.82 $Y2=0.74
cc_143 VPB N_A_1213_368#_c_798_n 0.00900487f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_144 VPB N_A_1213_368#_c_799_n 0.00192243f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_145 VPB N_A_1213_368#_c_800_n 0.0115811f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_1213_368#_c_801_n 0.0534124f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.515
cc_147 VPB N_A_1213_368#_c_802_n 0.00196551f $X=-0.19 $Y=1.66 $X2=1.395
+ $Y2=1.515
cc_148 VPB N_A_1213_368#_c_803_n 0.00196551f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.515
cc_149 VPB N_A_1213_368#_c_804_n 0.00196551f $X=-0.19 $Y=1.66 $X2=1.71 $Y2=1.515
cc_150 VPB N_Y_c_882_n 0.00432775f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.515
cc_151 VPB N_Y_c_883_n 0.00265801f $X=-0.19 $Y=1.66 $X2=0.69 $Y2=1.515
cc_152 VPB N_Y_c_877_n 0.00115545f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=1.515
cc_153 VPB N_Y_c_885_n 0.00137054f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_154 N_A3_M1027_g N_A2_M1002_g 0.0195801f $X=1.82 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A3_M1034_g N_A2_M1000_g 0.0212565f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A3_c_163_n A2 0.0381127f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_157 N_A3_c_158_n A2 0.00347669f $X=1.845 $Y=1.515 $X2=0 $Y2=0
cc_158 N_A3_c_163_n N_A2_c_232_n 3.7423e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_159 N_A3_c_158_n N_A2_c_232_n 0.029605f $X=1.845 $Y=1.515 $X2=0 $Y2=0
cc_160 N_A3_M1028_g N_VPWR_c_547_n 0.00551672f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_161 N_A3_M1028_g N_VPWR_c_548_n 5.60169e-19 $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_162 N_A3_M1029_g N_VPWR_c_548_n 0.0129122f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_163 N_A3_M1031_g N_VPWR_c_548_n 0.0127835f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_164 N_A3_M1034_g N_VPWR_c_548_n 5.41206e-19 $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_165 N_A3_M1031_g N_VPWR_c_549_n 5.41206e-19 $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_166 N_A3_M1034_g N_VPWR_c_549_n 0.0127537f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_167 N_A3_M1031_g N_VPWR_c_555_n 0.00460063f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_168 N_A3_M1034_g N_VPWR_c_555_n 0.00460063f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_169 N_A3_M1028_g N_VPWR_c_563_n 0.005209f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_170 N_A3_M1029_g N_VPWR_c_563_n 0.00460063f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_171 N_A3_M1028_g N_VPWR_c_545_n 0.00985972f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_172 N_A3_M1029_g N_VPWR_c_545_n 0.00908554f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_173 N_A3_M1031_g N_VPWR_c_545_n 0.00908554f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_174 N_A3_M1034_g N_VPWR_c_545_n 0.00908554f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_175 N_A3_M1028_g N_A_117_368#_c_697_n 0.0025567f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_176 N_A3_c_163_n N_A_117_368#_c_697_n 0.0189743f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_177 N_A3_c_158_n N_A_117_368#_c_697_n 5.53363e-19 $X=1.845 $Y=1.515 $X2=0
+ $Y2=0
cc_178 N_A3_M1028_g N_A_117_368#_c_686_n 0.0112102f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_179 N_A3_M1029_g N_A_117_368#_c_701_n 0.0142562f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_180 N_A3_M1031_g N_A_117_368#_c_701_n 0.0142562f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A3_c_163_n N_A_117_368#_c_701_n 0.0478981f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_182 N_A3_c_158_n N_A_117_368#_c_701_n 4.90767e-19 $X=1.845 $Y=1.515 $X2=0
+ $Y2=0
cc_183 N_A3_M1034_g N_A_117_368#_c_705_n 0.0159794f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_184 N_A3_c_163_n N_A_117_368#_c_705_n 0.0108884f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_185 N_A3_c_163_n N_A_117_368#_c_707_n 0.0143992f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_186 N_A3_c_158_n N_A_117_368#_c_707_n 5.5407e-19 $X=1.845 $Y=1.515 $X2=0
+ $Y2=0
cc_187 N_A3_M1010_g N_A_34_74#_c_965_n 0.00159319f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_188 N_A3_M1010_g N_A_34_74#_c_966_n 0.0157914f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A3_M1023_g N_A_34_74#_c_966_n 0.01115f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A3_c_163_n N_A_34_74#_c_966_n 0.0364045f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_191 N_A3_c_158_n N_A_34_74#_c_966_n 0.00443556f $X=1.845 $Y=1.515 $X2=0 $Y2=0
cc_192 N_A3_M1010_g N_A_34_74#_c_968_n 6.58468e-19 $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_193 N_A3_M1023_g N_A_34_74#_c_968_n 0.00918302f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A3_M1026_g N_A_34_74#_c_968_n 3.97481e-19 $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A3_M1026_g N_A_34_74#_c_969_n 0.0130918f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A3_M1027_g N_A_34_74#_c_969_n 0.0136838f $X=1.82 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A3_c_163_n N_A_34_74#_c_969_n 0.0460928f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_198 N_A3_c_158_n N_A_34_74#_c_969_n 0.0039811f $X=1.845 $Y=1.515 $X2=0 $Y2=0
cc_199 N_A3_M1027_g N_A_34_74#_c_970_n 3.92313e-19 $X=1.82 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A3_M1023_g N_A_34_74#_c_972_n 0.00157732f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A3_c_163_n N_A_34_74#_c_972_n 0.0213626f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_202 N_A3_c_158_n N_A_34_74#_c_972_n 0.00236901f $X=1.845 $Y=1.515 $X2=0 $Y2=0
cc_203 N_A3_M1010_g N_VGND_c_1039_n 0.0128874f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A3_M1023_g N_VGND_c_1039_n 0.00204878f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A3_M1023_g N_VGND_c_1040_n 5.19194e-19 $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A3_M1026_g N_VGND_c_1040_n 0.0108127f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A3_M1027_g N_VGND_c_1040_n 0.0107959f $X=1.82 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A3_M1010_g N_VGND_c_1042_n 0.00383152f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A3_M1023_g N_VGND_c_1043_n 0.00434272f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A3_M1026_g N_VGND_c_1043_n 0.00383152f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A3_M1010_g N_VGND_c_1046_n 0.00761312f $X=0.53 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A3_M1023_g N_VGND_c_1046_n 0.00820284f $X=0.96 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A3_M1026_g N_VGND_c_1046_n 0.0075754f $X=1.39 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A3_M1027_g N_VGND_c_1046_n 0.00757637f $X=1.82 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A3_M1027_g N_VGND_c_1049_n 0.00383152f $X=1.82 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A2_M1012_g N_A1_M1016_g 0.0213375f $X=3.645 $Y=2.4 $X2=0 $Y2=0
cc_217 A2 N_A1_c_308_n 0.00166304f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_218 N_A2_c_232_n N_A1_c_308_n 0.0213375f $X=3.54 $Y=1.515 $X2=0 $Y2=0
cc_219 N_A2_M1000_g N_VPWR_c_549_n 0.0127537f $X=2.295 $Y=2.4 $X2=0 $Y2=0
cc_220 N_A2_M1005_g N_VPWR_c_549_n 5.41206e-19 $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_221 N_A2_M1000_g N_VPWR_c_550_n 5.41206e-19 $X=2.295 $Y=2.4 $X2=0 $Y2=0
cc_222 N_A2_M1005_g N_VPWR_c_550_n 0.0127835f $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_223 N_A2_M1008_g N_VPWR_c_550_n 0.0127835f $X=3.195 $Y=2.4 $X2=0 $Y2=0
cc_224 N_A2_M1012_g N_VPWR_c_550_n 5.41206e-19 $X=3.645 $Y=2.4 $X2=0 $Y2=0
cc_225 N_A2_M1008_g N_VPWR_c_551_n 5.41206e-19 $X=3.195 $Y=2.4 $X2=0 $Y2=0
cc_226 N_A2_M1012_g N_VPWR_c_551_n 0.0127537f $X=3.645 $Y=2.4 $X2=0 $Y2=0
cc_227 N_A2_M1000_g N_VPWR_c_557_n 0.00460063f $X=2.295 $Y=2.4 $X2=0 $Y2=0
cc_228 N_A2_M1005_g N_VPWR_c_557_n 0.00460063f $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_229 N_A2_M1008_g N_VPWR_c_559_n 0.00460063f $X=3.195 $Y=2.4 $X2=0 $Y2=0
cc_230 N_A2_M1012_g N_VPWR_c_559_n 0.00460063f $X=3.645 $Y=2.4 $X2=0 $Y2=0
cc_231 N_A2_M1000_g N_VPWR_c_545_n 0.00908554f $X=2.295 $Y=2.4 $X2=0 $Y2=0
cc_232 N_A2_M1005_g N_VPWR_c_545_n 0.00908554f $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_233 N_A2_M1008_g N_VPWR_c_545_n 0.00908554f $X=3.195 $Y=2.4 $X2=0 $Y2=0
cc_234 N_A2_M1012_g N_VPWR_c_545_n 0.00908554f $X=3.645 $Y=2.4 $X2=0 $Y2=0
cc_235 N_A2_M1000_g N_A_117_368#_c_705_n 0.0142175f $X=2.295 $Y=2.4 $X2=0 $Y2=0
cc_236 A2 N_A_117_368#_c_705_n 0.0259404f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_237 N_A2_M1005_g N_A_117_368#_c_711_n 0.0142562f $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_238 N_A2_M1008_g N_A_117_368#_c_711_n 0.0142562f $X=3.195 $Y=2.4 $X2=0 $Y2=0
cc_239 A2 N_A_117_368#_c_711_n 0.0478981f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_240 N_A2_c_232_n N_A_117_368#_c_711_n 4.8583e-19 $X=3.54 $Y=1.515 $X2=0 $Y2=0
cc_241 N_A2_M1012_g N_A_117_368#_c_715_n 0.014793f $X=3.645 $Y=2.4 $X2=0 $Y2=0
cc_242 A2 N_A_117_368#_c_715_n 0.013807f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_243 A2 N_A_117_368#_c_717_n 0.0143992f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_244 N_A2_c_232_n N_A_117_368#_c_717_n 5.51241e-19 $X=3.54 $Y=1.515 $X2=0
+ $Y2=0
cc_245 A2 N_A_117_368#_c_719_n 0.0143992f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_246 N_A2_c_232_n N_A_117_368#_c_719_n 5.48413e-19 $X=3.54 $Y=1.515 $X2=0
+ $Y2=0
cc_247 N_A2_M1002_g N_A_34_74#_c_970_n 4.08775e-19 $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_248 N_A2_M1007_g N_A_34_74#_c_971_n 0.00914581f $X=3.11 $Y=0.74 $X2=0 $Y2=0
cc_249 N_A2_M1018_g N_A_34_74#_c_971_n 0.00983999f $X=3.54 $Y=0.74 $X2=0 $Y2=0
cc_250 N_A2_c_232_n N_A_34_74#_c_971_n 0.00264573f $X=3.54 $Y=1.515 $X2=0 $Y2=0
cc_251 A2 N_A_34_74#_c_973_n 0.00676262f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_252 N_A2_M1002_g N_A_34_74#_c_974_n 0.0142123f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A2_M1003_g N_A_34_74#_c_974_n 0.00913639f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_254 A2 N_A_34_74#_c_974_n 0.11368f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_255 N_A2_c_232_n N_A_34_74#_c_974_n 0.00248813f $X=3.54 $Y=1.515 $X2=0 $Y2=0
cc_256 N_A2_M1002_g N_A_34_74#_c_975_n 6.21182e-19 $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_257 N_A2_M1003_g N_A_34_74#_c_975_n 0.0058f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_258 N_A2_M1007_g N_A_34_74#_c_975_n 0.00554487f $X=3.11 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A2_M1018_g N_A_34_74#_c_975_n 6.0146e-19 $X=3.54 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A2_c_232_n N_A_34_74#_c_975_n 0.00260647f $X=3.54 $Y=1.515 $X2=0 $Y2=0
cc_261 N_A2_M1007_g N_A_34_74#_c_976_n 7.02574e-19 $X=3.11 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A2_M1018_g N_A_34_74#_c_976_n 0.00667962f $X=3.54 $Y=0.74 $X2=0 $Y2=0
cc_263 A2 N_A_34_74#_c_976_n 0.0101258f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_264 N_A2_c_232_n N_A_34_74#_c_976_n 0.00359664f $X=3.54 $Y=1.515 $X2=0 $Y2=0
cc_265 N_A2_M1002_g N_VGND_c_1040_n 6.96792e-19 $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_266 N_A2_M1002_g N_VGND_c_1046_n 0.00817716f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_267 N_A2_M1003_g N_VGND_c_1046_n 0.00359121f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_268 N_A2_M1007_g N_VGND_c_1046_n 0.00359121f $X=3.11 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A2_M1018_g N_VGND_c_1046_n 0.0036412f $X=3.54 $Y=0.74 $X2=0 $Y2=0
cc_270 N_A2_M1002_g N_VGND_c_1049_n 0.00433162f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_271 N_A2_M1003_g N_VGND_c_1049_n 0.00291649f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_272 N_A2_M1007_g N_VGND_c_1049_n 0.00291649f $X=3.11 $Y=0.74 $X2=0 $Y2=0
cc_273 N_A2_M1018_g N_VGND_c_1049_n 0.00291649f $X=3.54 $Y=0.74 $X2=0 $Y2=0
cc_274 N_A2_M1002_g N_A_465_74#_c_1128_n 0.00432482f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_275 N_A2_M1003_g N_A_465_74#_c_1129_n 0.0111551f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_276 N_A2_M1007_g N_A_465_74#_c_1129_n 0.0111551f $X=3.11 $Y=0.74 $X2=0 $Y2=0
cc_277 N_A2_M1018_g N_A_465_74#_c_1132_n 0.0141524f $X=3.54 $Y=0.74 $X2=0 $Y2=0
cc_278 N_A1_c_314_n N_B1_M1001_g 0.00966869f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_279 N_A1_M1025_g N_B1_M1017_g 0.0184495f $X=6 $Y=0.74 $X2=0 $Y2=0
cc_280 N_A1_M1025_g N_B1_c_396_n 0.00966869f $X=6 $Y=0.74 $X2=0 $Y2=0
cc_281 A1 N_B1_c_396_n 0.00868173f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_282 A1 N_B1_c_397_n 0.0093478f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_283 N_A1_M1016_g N_VPWR_c_551_n 0.0127537f $X=4.095 $Y=2.4 $X2=0 $Y2=0
cc_284 N_A1_M1020_g N_VPWR_c_551_n 5.41206e-19 $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_285 N_A1_M1016_g N_VPWR_c_552_n 5.43099e-19 $X=4.095 $Y=2.4 $X2=0 $Y2=0
cc_286 N_A1_M1020_g N_VPWR_c_552_n 0.0124151f $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_287 N_A1_M1022_g N_VPWR_c_552_n 0.00166074f $X=4.995 $Y=2.4 $X2=0 $Y2=0
cc_288 N_A1_M1022_g N_VPWR_c_553_n 0.005209f $X=4.995 $Y=2.4 $X2=0 $Y2=0
cc_289 N_A1_M1030_g N_VPWR_c_553_n 0.00460063f $X=5.445 $Y=2.4 $X2=0 $Y2=0
cc_290 N_A1_M1022_g N_VPWR_c_554_n 5.60169e-19 $X=4.995 $Y=2.4 $X2=0 $Y2=0
cc_291 N_A1_M1030_g N_VPWR_c_554_n 0.0140137f $X=5.445 $Y=2.4 $X2=0 $Y2=0
cc_292 N_A1_M1016_g N_VPWR_c_561_n 0.00460063f $X=4.095 $Y=2.4 $X2=0 $Y2=0
cc_293 N_A1_M1020_g N_VPWR_c_561_n 0.00460063f $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_294 N_A1_M1016_g N_VPWR_c_545_n 0.00908554f $X=4.095 $Y=2.4 $X2=0 $Y2=0
cc_295 N_A1_M1020_g N_VPWR_c_545_n 0.00908554f $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_296 N_A1_M1022_g N_VPWR_c_545_n 0.00982266f $X=4.995 $Y=2.4 $X2=0 $Y2=0
cc_297 N_A1_M1030_g N_VPWR_c_545_n 0.00908554f $X=5.445 $Y=2.4 $X2=0 $Y2=0
cc_298 N_A1_M1016_g N_A_117_368#_c_715_n 0.0191313f $X=4.095 $Y=2.4 $X2=0 $Y2=0
cc_299 N_A1_M1016_g N_A_117_368#_c_690_n 3.62369e-19 $X=4.095 $Y=2.4 $X2=0 $Y2=0
cc_300 N_A1_M1020_g N_A_117_368#_c_690_n 3.62369e-19 $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_301 N_A1_M1020_g N_A_117_368#_c_724_n 0.01917f $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_302 N_A1_M1022_g N_A_117_368#_c_724_n 0.012931f $X=4.995 $Y=2.4 $X2=0 $Y2=0
cc_303 A1 N_A_117_368#_c_724_n 0.0282763f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_304 N_A1_c_314_n N_A_117_368#_c_724_n 4.84419e-19 $X=5.91 $Y=1.515 $X2=0
+ $Y2=0
cc_305 N_A1_M1020_g N_A_117_368#_c_691_n 6.76823e-19 $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_306 N_A1_M1022_g N_A_117_368#_c_691_n 0.0120823f $X=4.995 $Y=2.4 $X2=0 $Y2=0
cc_307 N_A1_M1030_g N_A_117_368#_c_692_n 0.0163793f $X=5.445 $Y=2.4 $X2=0 $Y2=0
cc_308 A1 N_A_117_368#_c_692_n 0.0597519f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_309 N_A1_c_314_n N_A_117_368#_c_692_n 0.00281062f $X=5.91 $Y=1.515 $X2=0
+ $Y2=0
cc_310 N_A1_M1016_g N_A_117_368#_c_695_n 4.63009e-19 $X=4.095 $Y=2.4 $X2=0 $Y2=0
cc_311 N_A1_c_307_n N_A_117_368#_c_695_n 0.00382195f $X=4.455 $Y=1.605 $X2=0
+ $Y2=0
cc_312 N_A1_M1020_g N_A_117_368#_c_695_n 4.63009e-19 $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_313 N_A1_M1022_g N_A_117_368#_c_736_n 8.84614e-19 $X=4.995 $Y=2.4 $X2=0 $Y2=0
cc_314 A1 N_A_117_368#_c_736_n 0.0189743f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_315 N_A1_c_314_n N_A_117_368#_c_736_n 5.48413e-19 $X=5.91 $Y=1.515 $X2=0
+ $Y2=0
cc_316 N_A1_M1030_g N_A_1213_368#_c_796_n 5.89323e-19 $X=5.445 $Y=2.4 $X2=0
+ $Y2=0
cc_317 N_A1_M1004_g N_Y_c_874_n 0.0106768f $X=4.71 $Y=0.74 $X2=0 $Y2=0
cc_318 N_A1_M1015_g N_Y_c_874_n 0.0123927f $X=5.14 $Y=0.74 $X2=0 $Y2=0
cc_319 N_A1_M1019_g N_Y_c_874_n 0.0123136f $X=5.57 $Y=0.74 $X2=0 $Y2=0
cc_320 N_A1_M1025_g N_Y_c_874_n 0.0132419f $X=6 $Y=0.74 $X2=0 $Y2=0
cc_321 N_A1_c_314_n N_Y_c_874_n 0.00734485f $X=5.91 $Y=1.515 $X2=0 $Y2=0
cc_322 N_A1_M1025_g N_Y_c_875_n 4.15473e-19 $X=6 $Y=0.74 $X2=0 $Y2=0
cc_323 N_A1_c_307_n N_Y_c_878_n 0.010486f $X=4.455 $Y=1.605 $X2=0 $Y2=0
cc_324 N_A1_M1004_g N_Y_c_878_n 0.00318903f $X=4.71 $Y=0.74 $X2=0 $Y2=0
cc_325 N_A1_M1015_g N_Y_c_878_n 3.85913e-19 $X=5.14 $Y=0.74 $X2=0 $Y2=0
cc_326 A1 N_Y_c_878_n 0.0949302f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_327 N_A1_M1004_g N_VGND_c_1046_n 0.0036412f $X=4.71 $Y=0.74 $X2=0 $Y2=0
cc_328 N_A1_M1015_g N_VGND_c_1046_n 0.00359121f $X=5.14 $Y=0.74 $X2=0 $Y2=0
cc_329 N_A1_M1019_g N_VGND_c_1046_n 0.00359121f $X=5.57 $Y=0.74 $X2=0 $Y2=0
cc_330 N_A1_M1025_g N_VGND_c_1046_n 0.00449183f $X=6 $Y=0.74 $X2=0 $Y2=0
cc_331 N_A1_M1004_g N_VGND_c_1049_n 0.00291649f $X=4.71 $Y=0.74 $X2=0 $Y2=0
cc_332 N_A1_M1015_g N_VGND_c_1049_n 0.00291649f $X=5.14 $Y=0.74 $X2=0 $Y2=0
cc_333 N_A1_M1019_g N_VGND_c_1049_n 0.00291649f $X=5.57 $Y=0.74 $X2=0 $Y2=0
cc_334 N_A1_M1025_g N_VGND_c_1049_n 0.00433162f $X=6 $Y=0.74 $X2=0 $Y2=0
cc_335 N_A1_M1015_g N_A_465_74#_c_1131_n 3.85913e-19 $X=5.14 $Y=0.74 $X2=0 $Y2=0
cc_336 N_A1_M1019_g N_A_465_74#_c_1131_n 0.00281528f $X=5.57 $Y=0.74 $X2=0 $Y2=0
cc_337 N_A1_M1025_g N_A_465_74#_c_1131_n 0.00420713f $X=6 $Y=0.74 $X2=0 $Y2=0
cc_338 N_A1_M1004_g N_A_465_74#_c_1132_n 0.0136253f $X=4.71 $Y=0.74 $X2=0 $Y2=0
cc_339 N_A1_M1015_g N_A_465_74#_c_1132_n 0.0106927f $X=5.14 $Y=0.74 $X2=0 $Y2=0
cc_340 N_A1_M1019_g N_A_465_74#_c_1132_n 0.00920696f $X=5.57 $Y=0.74 $X2=0 $Y2=0
cc_341 N_B1_M1024_g N_C1_c_469_n 0.0122583f $X=7.71 $Y=0.74 $X2=-0.19 $Y2=-0.245
cc_342 B1 N_C1_M1009_g 5.47575e-19 $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_343 N_B1_c_396_n N_C1_M1009_g 0.0236751f $X=7.71 $Y=1.485 $X2=0 $Y2=0
cc_344 B1 N_C1_c_477_n 2.83059e-19 $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_345 N_B1_c_396_n N_C1_c_477_n 0.0156072f $X=7.71 $Y=1.485 $X2=0 $Y2=0
cc_346 N_B1_M1024_g N_C1_c_478_n 3.74992e-19 $X=7.71 $Y=0.74 $X2=0 $Y2=0
cc_347 B1 N_C1_c_478_n 0.0168871f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_348 N_B1_c_396_n N_C1_c_478_n 4.37969e-19 $X=7.71 $Y=1.485 $X2=0 $Y2=0
cc_349 N_B1_M1001_g N_VPWR_c_554_n 0.0018525f $X=6.415 $Y=2.4 $X2=0 $Y2=0
cc_350 N_B1_M1001_g N_VPWR_c_564_n 0.00333896f $X=6.415 $Y=2.4 $X2=0 $Y2=0
cc_351 N_B1_M1006_g N_VPWR_c_564_n 0.00333896f $X=6.865 $Y=2.4 $X2=0 $Y2=0
cc_352 N_B1_M1032_g N_VPWR_c_564_n 0.00333896f $X=7.315 $Y=2.4 $X2=0 $Y2=0
cc_353 N_B1_M1035_g N_VPWR_c_564_n 0.00333896f $X=7.765 $Y=2.4 $X2=0 $Y2=0
cc_354 N_B1_M1001_g N_VPWR_c_545_n 0.00427818f $X=6.415 $Y=2.4 $X2=0 $Y2=0
cc_355 N_B1_M1006_g N_VPWR_c_545_n 0.00422685f $X=6.865 $Y=2.4 $X2=0 $Y2=0
cc_356 N_B1_M1032_g N_VPWR_c_545_n 0.00422685f $X=7.315 $Y=2.4 $X2=0 $Y2=0
cc_357 N_B1_M1035_g N_VPWR_c_545_n 0.00422796f $X=7.765 $Y=2.4 $X2=0 $Y2=0
cc_358 N_B1_M1001_g N_A_117_368#_c_692_n 0.0187057f $X=6.415 $Y=2.4 $X2=0 $Y2=0
cc_359 N_B1_M1006_g N_A_117_368#_c_693_n 0.0195653f $X=6.865 $Y=2.4 $X2=0 $Y2=0
cc_360 N_B1_M1032_g N_A_117_368#_c_693_n 0.0195966f $X=7.315 $Y=2.4 $X2=0 $Y2=0
cc_361 B1 N_A_117_368#_c_693_n 0.0081802f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_362 N_B1_c_396_n N_A_117_368#_c_693_n 0.00205041f $X=7.71 $Y=1.485 $X2=0
+ $Y2=0
cc_363 N_B1_c_397_n N_A_117_368#_c_693_n 0.0431052f $X=7.32 $Y=1.415 $X2=0 $Y2=0
cc_364 B1 N_A_117_368#_c_694_n 0.0197666f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_365 N_B1_c_396_n N_A_117_368#_c_694_n 7.08547e-19 $X=7.71 $Y=1.485 $X2=0
+ $Y2=0
cc_366 N_B1_M1001_g N_A_117_368#_c_696_n 0.011167f $X=6.415 $Y=2.4 $X2=0 $Y2=0
cc_367 N_B1_c_396_n N_A_117_368#_c_696_n 0.00399972f $X=7.71 $Y=1.485 $X2=0
+ $Y2=0
cc_368 N_B1_M1001_g N_A_1213_368#_c_794_n 0.00872426f $X=6.415 $Y=2.4 $X2=0
+ $Y2=0
cc_369 N_B1_M1006_g N_A_1213_368#_c_794_n 5.45116e-19 $X=6.865 $Y=2.4 $X2=0
+ $Y2=0
cc_370 N_B1_M1001_g N_A_1213_368#_c_795_n 0.0116345f $X=6.415 $Y=2.4 $X2=0 $Y2=0
cc_371 N_B1_M1006_g N_A_1213_368#_c_795_n 0.0116345f $X=6.865 $Y=2.4 $X2=0 $Y2=0
cc_372 N_B1_M1001_g N_A_1213_368#_c_796_n 0.00291744f $X=6.415 $Y=2.4 $X2=0
+ $Y2=0
cc_373 N_B1_M1001_g N_A_1213_368#_c_811_n 5.45116e-19 $X=6.415 $Y=2.4 $X2=0
+ $Y2=0
cc_374 N_B1_M1006_g N_A_1213_368#_c_811_n 0.0085173f $X=6.865 $Y=2.4 $X2=0 $Y2=0
cc_375 N_B1_M1032_g N_A_1213_368#_c_811_n 0.0085173f $X=7.315 $Y=2.4 $X2=0 $Y2=0
cc_376 N_B1_M1035_g N_A_1213_368#_c_811_n 5.45116e-19 $X=7.765 $Y=2.4 $X2=0
+ $Y2=0
cc_377 N_B1_M1032_g N_A_1213_368#_c_797_n 0.0116345f $X=7.315 $Y=2.4 $X2=0 $Y2=0
cc_378 N_B1_M1035_g N_A_1213_368#_c_797_n 0.0116345f $X=7.765 $Y=2.4 $X2=0 $Y2=0
cc_379 N_B1_M1032_g N_A_1213_368#_c_798_n 6.88212e-19 $X=7.315 $Y=2.4 $X2=0
+ $Y2=0
cc_380 N_B1_M1035_g N_A_1213_368#_c_798_n 0.0156019f $X=7.765 $Y=2.4 $X2=0 $Y2=0
cc_381 N_B1_M1006_g N_A_1213_368#_c_802_n 0.00194226f $X=6.865 $Y=2.4 $X2=0
+ $Y2=0
cc_382 N_B1_M1032_g N_A_1213_368#_c_802_n 0.00194226f $X=7.315 $Y=2.4 $X2=0
+ $Y2=0
cc_383 N_B1_M1035_g N_A_1213_368#_c_803_n 0.001916f $X=7.765 $Y=2.4 $X2=0 $Y2=0
cc_384 N_B1_M1017_g N_Y_c_875_n 0.0114845f $X=6.43 $Y=0.74 $X2=0 $Y2=0
cc_385 N_B1_M1017_g N_Y_c_897_n 0.0143576f $X=6.43 $Y=0.74 $X2=0 $Y2=0
cc_386 N_B1_M1024_g N_Y_c_897_n 0.0112203f $X=7.71 $Y=0.74 $X2=0 $Y2=0
cc_387 B1 N_Y_c_897_n 0.0268604f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_388 N_B1_c_396_n N_Y_c_897_n 0.00994673f $X=7.71 $Y=1.485 $X2=0 $Y2=0
cc_389 N_B1_c_397_n N_Y_c_897_n 0.0436852f $X=7.32 $Y=1.415 $X2=0 $Y2=0
cc_390 N_B1_M1024_g N_Y_c_876_n 0.0109447f $X=7.71 $Y=0.74 $X2=0 $Y2=0
cc_391 N_B1_M1017_g N_Y_c_879_n 0.00755467f $X=6.43 $Y=0.74 $X2=0 $Y2=0
cc_392 N_B1_c_396_n N_Y_c_879_n 0.00142058f $X=7.71 $Y=1.485 $X2=0 $Y2=0
cc_393 N_B1_M1024_g N_Y_c_905_n 0.0024979f $X=7.71 $Y=0.74 $X2=0 $Y2=0
cc_394 B1 N_Y_c_905_n 0.00135505f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_395 N_B1_c_396_n N_Y_c_905_n 0.0014934f $X=7.71 $Y=1.485 $X2=0 $Y2=0
cc_396 N_B1_M1024_g N_VGND_c_1041_n 4.39708e-19 $X=7.71 $Y=0.74 $X2=0 $Y2=0
cc_397 N_B1_M1024_g N_VGND_c_1044_n 0.00434272f $X=7.71 $Y=0.74 $X2=0 $Y2=0
cc_398 N_B1_M1017_g N_VGND_c_1046_n 0.00449911f $X=6.43 $Y=0.74 $X2=0 $Y2=0
cc_399 N_B1_M1024_g N_VGND_c_1046_n 0.00449911f $X=7.71 $Y=0.74 $X2=0 $Y2=0
cc_400 N_B1_M1017_g N_VGND_c_1049_n 0.00434272f $X=6.43 $Y=0.74 $X2=0 $Y2=0
cc_401 N_B1_M1017_g N_VGND_c_1050_n 0.0113932f $X=6.43 $Y=0.74 $X2=0 $Y2=0
cc_402 N_B1_M1024_g N_VGND_c_1050_n 0.00963538f $X=7.71 $Y=0.74 $X2=0 $Y2=0
cc_403 N_C1_M1009_g N_VPWR_c_564_n 0.00333896f $X=8.215 $Y=2.4 $X2=0 $Y2=0
cc_404 N_C1_M1013_g N_VPWR_c_564_n 0.00333896f $X=8.665 $Y=2.4 $X2=0 $Y2=0
cc_405 N_C1_M1014_g N_VPWR_c_564_n 0.00333896f $X=9.115 $Y=2.4 $X2=0 $Y2=0
cc_406 N_C1_M1021_g N_VPWR_c_564_n 0.00333896f $X=9.565 $Y=2.4 $X2=0 $Y2=0
cc_407 N_C1_M1009_g N_VPWR_c_545_n 0.00422796f $X=8.215 $Y=2.4 $X2=0 $Y2=0
cc_408 N_C1_M1013_g N_VPWR_c_545_n 0.00422685f $X=8.665 $Y=2.4 $X2=0 $Y2=0
cc_409 N_C1_M1014_g N_VPWR_c_545_n 0.00422685f $X=9.115 $Y=2.4 $X2=0 $Y2=0
cc_410 N_C1_M1021_g N_VPWR_c_545_n 0.00426461f $X=9.565 $Y=2.4 $X2=0 $Y2=0
cc_411 N_C1_M1009_g N_A_1213_368#_c_798_n 0.0154197f $X=8.215 $Y=2.4 $X2=0 $Y2=0
cc_412 N_C1_M1013_g N_A_1213_368#_c_798_n 7.29961e-19 $X=8.665 $Y=2.4 $X2=0
+ $Y2=0
cc_413 N_C1_c_477_n N_A_1213_368#_c_798_n 4.44665e-19 $X=9.205 $Y=1.385 $X2=0
+ $Y2=0
cc_414 N_C1_c_478_n N_A_1213_368#_c_798_n 0.00519847f $X=8.47 $Y=1.365 $X2=0
+ $Y2=0
cc_415 N_C1_M1009_g N_A_1213_368#_c_799_n 0.0116345f $X=8.215 $Y=2.4 $X2=0 $Y2=0
cc_416 N_C1_M1013_g N_A_1213_368#_c_799_n 0.0116345f $X=8.665 $Y=2.4 $X2=0 $Y2=0
cc_417 N_C1_M1009_g N_A_1213_368#_c_828_n 6.45773e-19 $X=8.215 $Y=2.4 $X2=0
+ $Y2=0
cc_418 N_C1_M1013_g N_A_1213_368#_c_828_n 0.0139917f $X=8.665 $Y=2.4 $X2=0 $Y2=0
cc_419 N_C1_M1014_g N_A_1213_368#_c_828_n 0.0139917f $X=9.115 $Y=2.4 $X2=0 $Y2=0
cc_420 N_C1_M1021_g N_A_1213_368#_c_828_n 6.45773e-19 $X=9.565 $Y=2.4 $X2=0
+ $Y2=0
cc_421 N_C1_M1014_g N_A_1213_368#_c_800_n 0.0116345f $X=9.115 $Y=2.4 $X2=0 $Y2=0
cc_422 N_C1_M1021_g N_A_1213_368#_c_800_n 0.014552f $X=9.565 $Y=2.4 $X2=0 $Y2=0
cc_423 N_C1_M1014_g N_A_1213_368#_c_801_n 7.29961e-19 $X=9.115 $Y=2.4 $X2=0
+ $Y2=0
cc_424 N_C1_M1021_g N_A_1213_368#_c_801_n 0.0169226f $X=9.565 $Y=2.4 $X2=0 $Y2=0
cc_425 N_C1_M1009_g N_A_1213_368#_c_803_n 0.001916f $X=8.215 $Y=2.4 $X2=0 $Y2=0
cc_426 N_C1_M1013_g N_A_1213_368#_c_804_n 0.00194226f $X=8.665 $Y=2.4 $X2=0
+ $Y2=0
cc_427 N_C1_M1014_g N_A_1213_368#_c_804_n 0.00194226f $X=9.115 $Y=2.4 $X2=0
+ $Y2=0
cc_428 N_C1_M1013_g N_Y_c_882_n 0.0152733f $X=8.665 $Y=2.4 $X2=0 $Y2=0
cc_429 N_C1_M1014_g N_Y_c_882_n 0.0189242f $X=9.115 $Y=2.4 $X2=0 $Y2=0
cc_430 N_C1_c_476_n N_Y_c_882_n 0.0408056f $X=8.91 $Y=1.385 $X2=0 $Y2=0
cc_431 N_C1_c_477_n N_Y_c_882_n 0.00201785f $X=9.205 $Y=1.385 $X2=0 $Y2=0
cc_432 N_C1_M1009_g N_Y_c_883_n 0.00336f $X=8.215 $Y=2.4 $X2=0 $Y2=0
cc_433 N_C1_c_476_n N_Y_c_883_n 0.00463739f $X=8.91 $Y=1.385 $X2=0 $Y2=0
cc_434 N_C1_c_477_n N_Y_c_883_n 9.96062e-19 $X=9.205 $Y=1.385 $X2=0 $Y2=0
cc_435 N_C1_c_478_n N_Y_c_883_n 0.00982302f $X=8.47 $Y=1.365 $X2=0 $Y2=0
cc_436 N_C1_c_471_n N_Y_c_877_n 0.00275313f $X=8.57 $Y=1.22 $X2=0 $Y2=0
cc_437 N_C1_c_474_n N_Y_c_877_n 0.0226183f $X=9.475 $Y=1.345 $X2=0 $Y2=0
cc_438 N_C1_M1021_g N_Y_c_877_n 0.00599051f $X=9.565 $Y=2.4 $X2=0 $Y2=0
cc_439 N_C1_c_476_n N_Y_c_877_n 0.0273925f $X=8.91 $Y=1.385 $X2=0 $Y2=0
cc_440 N_C1_c_477_n N_Y_c_877_n 0.00478936f $X=9.205 $Y=1.385 $X2=0 $Y2=0
cc_441 N_C1_M1021_g N_Y_c_885_n 0.00336f $X=9.565 $Y=2.4 $X2=0 $Y2=0
cc_442 N_C1_c_474_n Y 0.00681241f $X=9.475 $Y=1.345 $X2=0 $Y2=0
cc_443 N_C1_c_469_n N_Y_c_923_n 0.00985057f $X=8.14 $Y=1.22 $X2=0 $Y2=0
cc_444 N_C1_c_471_n N_Y_c_923_n 0.00961729f $X=8.57 $Y=1.22 $X2=0 $Y2=0
cc_445 N_C1_c_476_n N_Y_c_923_n 0.046849f $X=8.91 $Y=1.385 $X2=0 $Y2=0
cc_446 N_C1_c_477_n N_Y_c_923_n 6.22937e-19 $X=9.205 $Y=1.385 $X2=0 $Y2=0
cc_447 N_C1_c_478_n N_Y_c_923_n 0.0251469f $X=8.47 $Y=1.365 $X2=0 $Y2=0
cc_448 N_C1_c_471_n N_Y_c_881_n 8.21094e-19 $X=8.57 $Y=1.22 $X2=0 $Y2=0
cc_449 N_C1_c_474_n N_Y_c_881_n 7.19437e-19 $X=9.475 $Y=1.345 $X2=0 $Y2=0
cc_450 N_C1_c_477_n N_Y_c_881_n 0.0111192f $X=9.205 $Y=1.385 $X2=0 $Y2=0
cc_451 N_C1_c_469_n N_VGND_c_1041_n 0.00769352f $X=8.14 $Y=1.22 $X2=0 $Y2=0
cc_452 N_C1_c_471_n N_VGND_c_1041_n 0.0105522f $X=8.57 $Y=1.22 $X2=0 $Y2=0
cc_453 N_C1_c_469_n N_VGND_c_1044_n 0.00383152f $X=8.14 $Y=1.22 $X2=0 $Y2=0
cc_454 N_C1_c_471_n N_VGND_c_1045_n 0.00383152f $X=8.57 $Y=1.22 $X2=0 $Y2=0
cc_455 N_C1_c_469_n N_VGND_c_1046_n 0.00384065f $X=8.14 $Y=1.22 $X2=0 $Y2=0
cc_456 N_C1_c_471_n N_VGND_c_1046_n 0.00388966f $X=8.57 $Y=1.22 $X2=0 $Y2=0
cc_457 N_VPWR_c_547_n N_A_117_368#_c_686_n 0.0277973f $X=0.27 $Y=1.985 $X2=0
+ $Y2=0
cc_458 N_VPWR_c_548_n N_A_117_368#_c_686_n 0.0234083f $X=1.17 $Y=2.455 $X2=0
+ $Y2=0
cc_459 N_VPWR_c_563_n N_A_117_368#_c_686_n 0.0109793f $X=1.005 $Y=3.33 $X2=0
+ $Y2=0
cc_460 N_VPWR_c_545_n N_A_117_368#_c_686_n 0.00901959f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_461 N_VPWR_M1029_s N_A_117_368#_c_701_n 0.00314376f $X=1.035 $Y=1.84 $X2=0
+ $Y2=0
cc_462 N_VPWR_c_548_n N_A_117_368#_c_701_n 0.0170259f $X=1.17 $Y=2.455 $X2=0
+ $Y2=0
cc_463 N_VPWR_c_548_n N_A_117_368#_c_687_n 0.0233699f $X=1.17 $Y=2.455 $X2=0
+ $Y2=0
cc_464 N_VPWR_c_549_n N_A_117_368#_c_687_n 0.0233699f $X=2.07 $Y=2.455 $X2=0
+ $Y2=0
cc_465 N_VPWR_c_555_n N_A_117_368#_c_687_n 0.00749631f $X=1.905 $Y=3.33 $X2=0
+ $Y2=0
cc_466 N_VPWR_c_545_n N_A_117_368#_c_687_n 0.0062048f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_467 N_VPWR_M1034_s N_A_117_368#_c_705_n 0.00477813f $X=1.935 $Y=1.84 $X2=0
+ $Y2=0
cc_468 N_VPWR_c_549_n N_A_117_368#_c_705_n 0.0170259f $X=2.07 $Y=2.455 $X2=0
+ $Y2=0
cc_469 N_VPWR_c_549_n N_A_117_368#_c_688_n 0.0233699f $X=2.07 $Y=2.455 $X2=0
+ $Y2=0
cc_470 N_VPWR_c_550_n N_A_117_368#_c_688_n 0.0233699f $X=2.97 $Y=2.455 $X2=0
+ $Y2=0
cc_471 N_VPWR_c_557_n N_A_117_368#_c_688_n 0.00749631f $X=2.805 $Y=3.33 $X2=0
+ $Y2=0
cc_472 N_VPWR_c_545_n N_A_117_368#_c_688_n 0.0062048f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_473 N_VPWR_M1005_s N_A_117_368#_c_711_n 0.00314376f $X=2.835 $Y=1.84 $X2=0
+ $Y2=0
cc_474 N_VPWR_c_550_n N_A_117_368#_c_711_n 0.0170259f $X=2.97 $Y=2.455 $X2=0
+ $Y2=0
cc_475 N_VPWR_c_550_n N_A_117_368#_c_689_n 0.0233699f $X=2.97 $Y=2.455 $X2=0
+ $Y2=0
cc_476 N_VPWR_c_551_n N_A_117_368#_c_689_n 0.0233699f $X=3.87 $Y=2.455 $X2=0
+ $Y2=0
cc_477 N_VPWR_c_559_n N_A_117_368#_c_689_n 0.00749631f $X=3.705 $Y=3.33 $X2=0
+ $Y2=0
cc_478 N_VPWR_c_545_n N_A_117_368#_c_689_n 0.0062048f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_479 N_VPWR_M1012_s N_A_117_368#_c_715_n 0.00761058f $X=3.735 $Y=1.84 $X2=0
+ $Y2=0
cc_480 N_VPWR_c_551_n N_A_117_368#_c_715_n 0.0170259f $X=3.87 $Y=2.455 $X2=0
+ $Y2=0
cc_481 N_VPWR_c_551_n N_A_117_368#_c_690_n 0.0233699f $X=3.87 $Y=2.455 $X2=0
+ $Y2=0
cc_482 N_VPWR_c_552_n N_A_117_368#_c_690_n 0.022423f $X=4.77 $Y=2.455 $X2=0
+ $Y2=0
cc_483 N_VPWR_c_561_n N_A_117_368#_c_690_n 0.00749631f $X=4.605 $Y=3.33 $X2=0
+ $Y2=0
cc_484 N_VPWR_c_545_n N_A_117_368#_c_690_n 0.0062048f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_485 N_VPWR_M1020_s N_A_117_368#_c_724_n 0.00314376f $X=4.635 $Y=1.84 $X2=0
+ $Y2=0
cc_486 N_VPWR_c_552_n N_A_117_368#_c_724_n 0.0148589f $X=4.77 $Y=2.455 $X2=0
+ $Y2=0
cc_487 N_VPWR_c_552_n N_A_117_368#_c_691_n 0.0224614f $X=4.77 $Y=2.455 $X2=0
+ $Y2=0
cc_488 N_VPWR_c_553_n N_A_117_368#_c_691_n 0.0109793f $X=5.505 $Y=3.33 $X2=0
+ $Y2=0
cc_489 N_VPWR_c_554_n N_A_117_368#_c_691_n 0.0234083f $X=5.67 $Y=2.455 $X2=0
+ $Y2=0
cc_490 N_VPWR_c_545_n N_A_117_368#_c_691_n 0.00901959f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_491 N_VPWR_M1030_s N_A_117_368#_c_692_n 0.00466601f $X=5.535 $Y=1.84 $X2=0
+ $Y2=0
cc_492 N_VPWR_c_554_n N_A_117_368#_c_692_n 0.0219767f $X=5.67 $Y=2.455 $X2=0
+ $Y2=0
cc_493 N_VPWR_c_554_n N_A_1213_368#_c_794_n 0.0450078f $X=5.67 $Y=2.455 $X2=0
+ $Y2=0
cc_494 N_VPWR_c_564_n N_A_1213_368#_c_795_n 0.0357927f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_495 N_VPWR_c_545_n N_A_1213_368#_c_795_n 0.0200586f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_496 N_VPWR_c_554_n N_A_1213_368#_c_796_n 0.0139f $X=5.67 $Y=2.455 $X2=0 $Y2=0
cc_497 N_VPWR_c_564_n N_A_1213_368#_c_796_n 0.0235512f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_498 N_VPWR_c_545_n N_A_1213_368#_c_796_n 0.0126924f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_499 N_VPWR_c_564_n N_A_1213_368#_c_797_n 0.0357927f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_500 N_VPWR_c_545_n N_A_1213_368#_c_797_n 0.0200586f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_501 N_VPWR_c_564_n N_A_1213_368#_c_799_n 0.0357927f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_502 N_VPWR_c_545_n N_A_1213_368#_c_799_n 0.0200586f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_503 N_VPWR_c_564_n N_A_1213_368#_c_800_n 0.0593439f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_504 N_VPWR_c_545_n N_A_1213_368#_c_800_n 0.032751f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_505 N_VPWR_c_564_n N_A_1213_368#_c_802_n 0.0234458f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_506 N_VPWR_c_545_n N_A_1213_368#_c_802_n 0.0125551f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_507 N_VPWR_c_564_n N_A_1213_368#_c_803_n 0.0234458f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_508 N_VPWR_c_545_n N_A_1213_368#_c_803_n 0.0125551f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_509 N_VPWR_c_564_n N_A_1213_368#_c_804_n 0.0234458f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_510 N_VPWR_c_545_n N_A_1213_368#_c_804_n 0.0125551f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_511 N_VPWR_c_547_n N_A_34_74#_c_967_n 0.00754091f $X=0.27 $Y=1.985 $X2=0
+ $Y2=0
cc_512 N_A_117_368#_c_692_n N_A_1213_368#_M1001_s 0.00940859f $X=6.475 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_513 N_A_117_368#_c_693_n N_A_1213_368#_M1006_s 0.00169251f $X=7.425 $Y=1.985
+ $X2=0 $Y2=0
cc_514 N_A_117_368#_c_692_n N_A_1213_368#_c_794_n 0.0194698f $X=6.475 $Y=2.035
+ $X2=0 $Y2=0
cc_515 N_A_117_368#_M1001_d N_A_1213_368#_c_795_n 0.00165831f $X=6.505 $Y=1.84
+ $X2=0 $Y2=0
cc_516 N_A_117_368#_c_789_p N_A_1213_368#_c_795_n 0.0118736f $X=6.64 $Y=2.57
+ $X2=0 $Y2=0
cc_517 N_A_117_368#_c_693_n N_A_1213_368#_c_811_n 0.0178311f $X=7.425 $Y=1.985
+ $X2=0 $Y2=0
cc_518 N_A_117_368#_M1032_d N_A_1213_368#_c_797_n 0.00165831f $X=7.405 $Y=1.84
+ $X2=0 $Y2=0
cc_519 N_A_117_368#_c_792_p N_A_1213_368#_c_797_n 0.0118736f $X=7.54 $Y=2.57
+ $X2=0 $Y2=0
cc_520 N_A_117_368#_c_694_n N_A_1213_368#_c_798_n 0.0133269f $X=7.54 $Y=2.15
+ $X2=0 $Y2=0
cc_521 N_A_1213_368#_c_799_n N_Y_M1009_d 0.00165831f $X=8.725 $Y=2.99 $X2=0
+ $Y2=0
cc_522 N_A_1213_368#_c_800_n N_Y_M1014_d 0.00165831f $X=9.625 $Y=2.99 $X2=0
+ $Y2=0
cc_523 N_A_1213_368#_c_799_n N_Y_c_933_n 0.0118736f $X=8.725 $Y=2.99 $X2=0 $Y2=0
cc_524 N_A_1213_368#_M1013_s N_Y_c_882_n 0.00165831f $X=8.755 $Y=1.84 $X2=0
+ $Y2=0
cc_525 N_A_1213_368#_c_828_n N_Y_c_882_n 0.0170259f $X=8.89 $Y=2.225 $X2=0 $Y2=0
cc_526 N_A_1213_368#_c_798_n N_Y_c_883_n 0.00310493f $X=7.99 $Y=1.985 $X2=0
+ $Y2=0
cc_527 N_A_1213_368#_c_800_n N_Y_c_937_n 0.0118736f $X=9.625 $Y=2.99 $X2=0 $Y2=0
cc_528 N_A_1213_368#_c_801_n N_Y_c_885_n 0.00310493f $X=9.79 $Y=1.985 $X2=0
+ $Y2=0
cc_529 N_Y_c_878_n N_A_34_74#_c_976_n 0.0169912f $X=4.66 $Y=0.95 $X2=0 $Y2=0
cc_530 N_Y_c_897_n N_VGND_M1017_d 0.0286593f $X=7.76 $Y=0.925 $X2=0 $Y2=0
cc_531 N_Y_c_923_n N_VGND_M1011_s 0.00330259f $X=8.7 $Y=0.68 $X2=0 $Y2=0
cc_532 N_Y_c_876_n N_VGND_c_1041_n 0.0121972f $X=7.925 $Y=0.515 $X2=0 $Y2=0
cc_533 N_Y_c_923_n N_VGND_c_1041_n 0.0167019f $X=8.7 $Y=0.68 $X2=0 $Y2=0
cc_534 N_Y_c_881_n N_VGND_c_1041_n 0.0122903f $X=9.425 $Y=0.68 $X2=0 $Y2=0
cc_535 N_Y_c_876_n N_VGND_c_1044_n 0.0110175f $X=7.925 $Y=0.515 $X2=0 $Y2=0
cc_536 N_Y_c_881_n N_VGND_c_1045_n 0.0544421f $X=9.425 $Y=0.68 $X2=0 $Y2=0
cc_537 N_Y_c_874_n N_VGND_c_1046_n 0.00789134f $X=6.13 $Y=0.99 $X2=0 $Y2=0
cc_538 N_Y_c_875_n N_VGND_c_1046_n 0.00904371f $X=6.215 $Y=0.515 $X2=0 $Y2=0
cc_539 N_Y_c_897_n N_VGND_c_1046_n 0.0132757f $X=7.76 $Y=0.925 $X2=0 $Y2=0
cc_540 N_Y_c_876_n N_VGND_c_1046_n 0.0090528f $X=7.925 $Y=0.515 $X2=0 $Y2=0
cc_541 N_Y_c_923_n N_VGND_c_1046_n 0.0116543f $X=8.7 $Y=0.68 $X2=0 $Y2=0
cc_542 N_Y_c_881_n N_VGND_c_1046_n 0.0458137f $X=9.425 $Y=0.68 $X2=0 $Y2=0
cc_543 N_Y_c_875_n N_VGND_c_1049_n 0.0109942f $X=6.215 $Y=0.515 $X2=0 $Y2=0
cc_544 N_Y_c_875_n N_VGND_c_1050_n 0.0124113f $X=6.215 $Y=0.515 $X2=0 $Y2=0
cc_545 N_Y_c_897_n N_VGND_c_1050_n 0.0804627f $X=7.76 $Y=0.925 $X2=0 $Y2=0
cc_546 N_Y_c_876_n N_VGND_c_1050_n 0.0124113f $X=7.925 $Y=0.515 $X2=0 $Y2=0
cc_547 N_Y_c_874_n N_A_465_74#_M1004_s 0.00209854f $X=6.13 $Y=0.99 $X2=0 $Y2=0
cc_548 N_Y_c_874_n N_A_465_74#_M1019_s 0.00177318f $X=6.13 $Y=0.99 $X2=0 $Y2=0
cc_549 N_Y_c_874_n N_A_465_74#_c_1131_n 0.0163856f $X=6.13 $Y=0.99 $X2=0 $Y2=0
cc_550 N_Y_c_875_n N_A_465_74#_c_1131_n 0.0135554f $X=6.215 $Y=0.515 $X2=0 $Y2=0
cc_551 N_Y_M1004_d N_A_465_74#_c_1132_n 0.00332037f $X=4.37 $Y=0.37 $X2=0 $Y2=0
cc_552 N_Y_M1015_d N_A_465_74#_c_1132_n 0.00212678f $X=5.215 $Y=0.37 $X2=0 $Y2=0
cc_553 N_Y_c_874_n N_A_465_74#_c_1132_n 0.0379865f $X=6.13 $Y=0.99 $X2=0 $Y2=0
cc_554 N_Y_c_878_n N_A_465_74#_c_1132_n 0.0208358f $X=4.66 $Y=0.95 $X2=0 $Y2=0
cc_555 N_A_34_74#_c_966_n N_VGND_M1010_d 0.00176461f $X=1.01 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_556 N_A_34_74#_c_969_n N_VGND_M1026_d 0.00176461f $X=1.95 $Y=1.095 $X2=0
+ $Y2=0
cc_557 N_A_34_74#_c_965_n N_VGND_c_1039_n 0.0175587f $X=0.315 $Y=0.515 $X2=0
+ $Y2=0
cc_558 N_A_34_74#_c_966_n N_VGND_c_1039_n 0.0152916f $X=1.01 $Y=1.095 $X2=0
+ $Y2=0
cc_559 N_A_34_74#_c_968_n N_VGND_c_1039_n 0.0175587f $X=1.175 $Y=0.515 $X2=0
+ $Y2=0
cc_560 N_A_34_74#_c_968_n N_VGND_c_1040_n 0.0182902f $X=1.175 $Y=0.515 $X2=0
+ $Y2=0
cc_561 N_A_34_74#_c_969_n N_VGND_c_1040_n 0.0170777f $X=1.95 $Y=1.095 $X2=0
+ $Y2=0
cc_562 N_A_34_74#_c_970_n N_VGND_c_1040_n 0.0182488f $X=2.035 $Y=0.515 $X2=0
+ $Y2=0
cc_563 N_A_34_74#_c_965_n N_VGND_c_1042_n 0.011066f $X=0.315 $Y=0.515 $X2=0
+ $Y2=0
cc_564 N_A_34_74#_c_968_n N_VGND_c_1043_n 0.0109942f $X=1.175 $Y=0.515 $X2=0
+ $Y2=0
cc_565 N_A_34_74#_c_965_n N_VGND_c_1046_n 0.00915947f $X=0.315 $Y=0.515 $X2=0
+ $Y2=0
cc_566 N_A_34_74#_c_968_n N_VGND_c_1046_n 0.00904371f $X=1.175 $Y=0.515 $X2=0
+ $Y2=0
cc_567 N_A_34_74#_c_970_n N_VGND_c_1046_n 0.0062048f $X=2.035 $Y=0.515 $X2=0
+ $Y2=0
cc_568 N_A_34_74#_c_970_n N_VGND_c_1049_n 0.00749631f $X=2.035 $Y=0.515 $X2=0
+ $Y2=0
cc_569 N_A_34_74#_c_974_n N_A_465_74#_M1002_d 0.00229137f $X=2.73 $Y=0.975
+ $X2=-0.19 $Y2=-0.245
cc_570 N_A_34_74#_c_971_n N_A_465_74#_M1007_d 0.00229137f $X=3.59 $Y=1.077 $X2=0
+ $Y2=0
cc_571 N_A_34_74#_c_970_n N_A_465_74#_c_1128_n 0.0134146f $X=2.035 $Y=0.515
+ $X2=0 $Y2=0
cc_572 N_A_34_74#_c_974_n N_A_465_74#_c_1128_n 0.00971408f $X=2.73 $Y=0.975
+ $X2=0 $Y2=0
cc_573 N_A_34_74#_M1003_s N_A_465_74#_c_1129_n 0.00179007f $X=2.755 $Y=0.37
+ $X2=0 $Y2=0
cc_574 N_A_34_74#_c_971_n N_A_465_74#_c_1129_n 0.00465091f $X=3.59 $Y=1.077
+ $X2=0 $Y2=0
cc_575 N_A_34_74#_c_974_n N_A_465_74#_c_1129_n 0.00465091f $X=2.73 $Y=0.975
+ $X2=0 $Y2=0
cc_576 N_A_34_74#_c_975_n N_A_465_74#_c_1129_n 0.0163588f $X=3.06 $Y=0.975 $X2=0
+ $Y2=0
cc_577 N_A_34_74#_c_971_n N_A_465_74#_c_1130_n 0.00857327f $X=3.59 $Y=1.077
+ $X2=0 $Y2=0
cc_578 N_A_34_74#_M1018_s N_A_465_74#_c_1132_n 0.0033149f $X=3.615 $Y=0.37 $X2=0
+ $Y2=0
cc_579 N_A_34_74#_c_971_n N_A_465_74#_c_1132_n 0.00466938f $X=3.59 $Y=1.077
+ $X2=0 $Y2=0
cc_580 N_A_34_74#_c_976_n N_A_465_74#_c_1132_n 0.0209951f $X=3.755 $Y=0.95 $X2=0
+ $Y2=0
cc_581 N_VGND_c_1046_n N_A_465_74#_c_1128_n 0.126157f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_582 N_VGND_c_1049_n N_A_465_74#_c_1128_n 0.149195f $X=6.55 $Y=0.292 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__o22a_4.spice
* Created: Wed Sep  2 12:23:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o22a_4.pex.spice"
.subckt sky130_fd_sc_ms__o22a_4  VNB VPB A2 A1 B2 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* B2	B2
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1016 N_A_27_136#_M1016_d N_A1_M1016_g N_VGND_M1016_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.112 PD=1.85 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75000.2
+ SB=75003.6 A=0.096 P=1.58 MULT=1
MM1013 N_A_27_136#_M1013_d N_A2_M1013_g N_VGND_M1016_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.112 PD=0.92 PS=0.99 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.7
+ SB=75003.1 A=0.096 P=1.58 MULT=1
MM1014 N_A_27_136#_M1013_d N_A2_M1014_g N_VGND_M1014_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1248 PD=0.92 PS=1.03 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75001.1
+ SB=75002.6 A=0.096 P=1.58 MULT=1
MM1017 N_A_27_136#_M1017_d N_A1_M1017_g N_VGND_M1014_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.12 AS=0.1248 PD=1.015 PS=1.03 NRD=5.616 NRS=7.488 M=1 R=4.26667
+ SA=75001.7 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1005 N_A_27_136#_M1017_d N_B1_M1005_g N_A_209_392#_M1005_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.12 AS=0.0912 PD=1.015 PS=0.925 NRD=12.18 NRS=0.936 M=1 R=4.26667
+ SA=75002.2 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1010 N_A_209_392#_M1005_s N_B2_M1010_g N_A_27_136#_M1010_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0912 AS=0.1136 PD=0.925 PS=0.995 NRD=0 NRS=6.552 M=1 R=4.26667
+ SA=75002.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1012 N_A_209_392#_M1012_d N_B2_M1012_g N_A_27_136#_M1010_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1136 PD=0.92 PS=0.995 NRD=0 NRS=7.488 M=1 R=4.26667
+ SA=75003.1 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1020 N_A_27_136#_M1020_d N_B1_M1020_g N_A_209_392#_M1012_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75003.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1006_d N_A_209_392#_M1006_g N_X_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2991 AS=0.1036 PD=2.41 PS=1.02 NRD=13.776 NRS=0 M=1 R=4.93333 SA=75000.3
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_A_209_392#_M1008_g N_X_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1011 N_VGND_M1008_d N_A_209_392#_M1011_g N_X_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1018_d N_A_209_392#_M1018_g N_X_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2146 AS=0.1036 PD=2.06 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g N_A_119_392#_M1000_s VPB PSHORT L=0.18 W=1
+ AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90005.9 A=0.18 P=2.36 MULT=1
MM1001 N_A_119_392#_M1000_s N_A2_M1001_g N_A_209_392#_M1001_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.16 PD=1.27 PS=1.32 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90000.6
+ SB=90005.4 A=0.18 P=2.36 MULT=1
MM1003 N_A_119_392#_M1003_d N_A2_M1003_g N_A_209_392#_M1001_s VPB PSHORT L=0.18
+ W=1 AD=0.16 AS=0.16 PD=1.32 PS=1.32 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90001.1
+ SB=90004.9 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_119_392#_M1003_d VPB PSHORT L=0.18 W=1
+ AD=0.185 AS=0.16 PD=1.37 PS=1.32 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90001.6
+ SB=90004.4 A=0.18 P=2.36 MULT=1
MM1019 N_A_519_392#_M1019_d N_B1_M1019_g N_VPWR_M1002_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.185 PD=1.27 PS=1.37 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90002.2
+ SB=90003.9 A=0.18 P=2.36 MULT=1
MM1022 N_A_519_392#_M1019_d N_B2_M1022_g N_A_209_392#_M1022_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.16 PD=1.27 PS=1.32 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90002.6
+ SB=90003.4 A=0.18 P=2.36 MULT=1
MM1023 N_A_519_392#_M1023_d N_B2_M1023_g N_A_209_392#_M1022_s VPB PSHORT L=0.18
+ W=1 AD=0.16 AS=0.16 PD=1.32 PS=1.32 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90003.1
+ SB=90002.9 A=0.18 P=2.36 MULT=1
MM1021 N_A_519_392#_M1023_d N_B1_M1021_g N_VPWR_M1021_s VPB PSHORT L=0.18 W=1
+ AD=0.16 AS=0.191226 PD=1.32 PS=1.40566 NRD=0 NRS=16.0752 M=1 R=5.55556
+ SA=90003.6 SB=90002.4 A=0.18 P=2.36 MULT=1
MM1004 N_X_M1004_d N_A_209_392#_M1004_g N_VPWR_M1021_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1708 AS=0.214174 PD=1.425 PS=1.57434 NRD=5.2599 NRS=1.7533 M=1 R=6.22222
+ SA=90003.8 SB=90001.9 A=0.2016 P=2.6 MULT=1
MM1007 N_X_M1004_d N_A_209_392#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1708 AS=0.3052 PD=1.425 PS=1.665 NRD=0 NRS=25.4918 M=1 R=6.22222
+ SA=90004.2 SB=90001.4 A=0.2016 P=2.6 MULT=1
MM1009 N_X_M1009_d N_A_209_392#_M1009_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3052 PD=1.39 PS=1.665 NRD=0 NRS=21.0987 M=1 R=6.22222 SA=90005
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1015 N_X_M1009_d N_A_209_392#_M1015_g N_VPWR_M1015_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90005.4
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX24_noxref VNB VPB NWDIODE A=13.206 P=17.92
c_112 VPB 0 1.20589e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__o22a_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__dlxtn_1.spice
* Created: Fri Aug 28 17:29:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dlxtn_1.pex.spice"
.subckt sky130_fd_sc_ms__dlxtn_1  VNB VPB D GATE_N VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_D_M1005_g N_A_27_115#_M1005_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.171896 AS=0.15675 PD=1.33876 PS=1.67 NRD=56.184 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1009 N_A_220_419#_M1009_d N_GATE_N_M1009_g N_VGND_M1005_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.231279 PD=2.05 PS=1.80124 NRD=0 NRS=41.76 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A_220_419#_M1003_g N_A_369_392#_M1003_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.251922 AS=0.2109 PD=1.53899 PS=2.05 NRD=66.48 NRS=0 M=1
+ R=4.93333 SA=75000.2 SB=75002 A=0.111 P=1.78 MULT=1
MM1016 A_655_79# N_A_27_115#_M1016_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.217878 PD=0.88 PS=1.33101 NRD=12.18 NRS=0.936 M=1 R=4.26667
+ SA=75001.1 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1017 N_A_672_392#_M1017_d N_A_220_419#_M1017_g A_655_79# VNB NLOWVT L=0.15
+ W=0.64 AD=0.168211 AS=0.0768 PD=1.52151 PS=0.88 NRD=25.308 NRS=12.18 M=1
+ R=4.26667 SA=75001.4 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1007 A_871_139# N_A_369_392#_M1007_g N_A_672_392#_M1017_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.110389 PD=0.66 PS=0.998491 NRD=18.564 NRS=35.712 M=1
+ R=2.8 SA=75001.8 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_A_863_441#_M1012_g A_871_139# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0930736 AS=0.0504 PD=0.832075 PS=0.66 NRD=37.848 NRS=18.564 M=1 R=2.8
+ SA=75002.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1013 N_A_863_441#_M1013_d N_A_672_392#_M1013_g N_VGND_M1012_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.141826 PD=1.85 PS=1.26792 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75001.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_Q_M1001_d N_A_863_441#_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2146 AS=0.2109 PD=2.06 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1014 N_VPWR_M1014_d N_D_M1014_g N_A_27_115#_M1014_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1344 AS=0.2352 PD=1.16 PS=2.24 NRD=10.5395 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1011 N_A_220_419#_M1011_d N_GATE_N_M1011_g N_VPWR_M1014_d VPB PSHORT L=0.18
+ W=0.84 AD=0.3066 AS=0.1344 PD=2.41 PS=1.16 NRD=18.7544 NRS=0 M=1 R=4.66667
+ SA=90000.7 SB=90000.3 A=0.1512 P=2.04 MULT=1
MM1015 N_VPWR_M1015_d N_A_220_419#_M1015_g N_A_369_392#_M1015_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.22034 AS=0.2352 PD=1.44717 PS=2.24 NRD=48.5999 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90002 A=0.1512 P=2.04 MULT=1
MM1004 A_588_392# N_A_27_115#_M1004_g N_VPWR_M1015_d VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.26231 PD=1.24 PS=1.72283 NRD=12.7853 NRS=18.6953 M=1 R=5.55556
+ SA=90000.7 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1008 N_A_672_392#_M1008_d N_A_369_392#_M1008_g A_588_392# VPB PSHORT L=0.18
+ W=1 AD=0.346127 AS=0.12 PD=2.16197 PS=1.24 NRD=16.7253 NRS=12.7853 M=1
+ R=5.55556 SA=90001.2 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1000 A_815_508# N_A_220_419#_M1000_g N_A_672_392#_M1008_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.145373 PD=0.66 PS=0.908028 NRD=30.4759 NRS=82.0702 M=1
+ R=2.33333 SA=90001.8 SB=90001.4 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1010_d N_A_863_441#_M1010_g A_815_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.125054 AS=0.0504 PD=0.95831 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.33333
+ SA=90002.2 SB=90001 A=0.0756 P=1.2 MULT=1
MM1006 N_A_863_441#_M1006_d N_A_672_392#_M1006_g N_VPWR_M1010_d VPB PSHORT
+ L=0.18 W=1 AD=0.28 AS=0.297746 PD=2.56 PS=2.28169 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90001.4 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1002 N_Q_M1002_d N_A_863_441#_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.3136 PD=2.8 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX18_noxref VNB VPB NWDIODE A=13.206 P=17.92
c_73 VNB 0 4.76483e-20 $X=0 $Y=0
c_920 A_655_79# 0 3.15497e-20 $X=3.275 $Y=0.395
*
.include "sky130_fd_sc_ms__dlxtn_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__nor4_4.pex.spice
* Created: Fri Aug 28 17:49:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NOR4_4%D 3 7 11 15 19 23 25 26 27 40 41
c62 23 0 9.97624e-20 $X=1.955 $Y=2.4
r63 39 41 22.8076 $w=3.17e-07 $l=1.5e-07 $layer=POLY_cond $X=1.71 $Y=1.515
+ $X2=1.86 $Y2=1.515
r64 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.71
+ $Y=1.515 $X2=1.71 $Y2=1.515
r65 37 39 38.7729 $w=3.17e-07 $l=2.55e-07 $layer=POLY_cond $X=1.455 $Y=1.515
+ $X2=1.71 $Y2=1.515
r66 36 37 68.4227 $w=3.17e-07 $l=4.5e-07 $layer=POLY_cond $X=1.005 $Y=1.515
+ $X2=1.455 $Y2=1.515
r67 34 36 47.8959 $w=3.17e-07 $l=3.15e-07 $layer=POLY_cond $X=0.69 $Y=1.515
+ $X2=1.005 $Y2=1.515
r68 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.69
+ $Y=1.515 $X2=0.69 $Y2=1.515
r69 32 34 20.5268 $w=3.17e-07 $l=1.35e-07 $layer=POLY_cond $X=0.555 $Y=1.515
+ $X2=0.69 $Y2=1.515
r70 31 32 2.28076 $w=3.17e-07 $l=1.5e-08 $layer=POLY_cond $X=0.54 $Y=1.515
+ $X2=0.555 $Y2=1.515
r71 27 40 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=1.68 $Y=1.565 $X2=1.71
+ $Y2=1.565
r72 26 27 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.68 $Y2=1.565
r73 25 26 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r74 25 35 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=0.72 $Y=1.565 $X2=0.69
+ $Y2=1.565
r75 21 41 14.4448 $w=3.17e-07 $l=2.07123e-07 $layer=POLY_cond $X=1.955 $Y=1.68
+ $X2=1.86 $Y2=1.515
r76 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.955 $Y=1.68
+ $X2=1.955 $Y2=2.4
r77 17 41 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.86 $Y=1.35
+ $X2=1.86 $Y2=1.515
r78 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.86 $Y=1.35
+ $X2=1.86 $Y2=0.74
r79 13 37 15.9969 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.455 $Y=1.68
+ $X2=1.455 $Y2=1.515
r80 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.455 $Y=1.68
+ $X2=1.455 $Y2=2.4
r81 9 36 15.9969 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.68
+ $X2=1.005 $Y2=1.515
r82 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.005 $Y=1.68
+ $X2=1.005 $Y2=2.4
r83 5 32 15.9969 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.68
+ $X2=0.555 $Y2=1.515
r84 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.555 $Y=1.68
+ $X2=0.555 $Y2=2.4
r85 1 31 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.35 $X2=0.54
+ $Y2=1.515
r86 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.54 $Y=1.35 $X2=0.54
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4_4%C 3 7 11 15 19 23 25 26 27 40 41
c69 19 0 1.56424e-19 $X=3.71 $Y=0.74
r70 41 42 6.71517 $w=3.23e-07 $l=4.5e-08 $layer=POLY_cond $X=3.71 $Y=1.515
+ $X2=3.755 $Y2=1.515
r71 39 41 13.4303 $w=3.23e-07 $l=9e-08 $layer=POLY_cond $X=3.62 $Y=1.515
+ $X2=3.71 $Y2=1.515
r72 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.62
+ $Y=1.515 $X2=3.62 $Y2=1.515
r73 37 39 47.0062 $w=3.23e-07 $l=3.15e-07 $layer=POLY_cond $X=3.305 $Y=1.515
+ $X2=3.62 $Y2=1.515
r74 36 37 67.1517 $w=3.23e-07 $l=4.5e-07 $layer=POLY_cond $X=2.855 $Y=1.515
+ $X2=3.305 $Y2=1.515
r75 34 36 38.0526 $w=3.23e-07 $l=2.55e-07 $layer=POLY_cond $X=2.6 $Y=1.515
+ $X2=2.855 $Y2=1.515
r76 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.6
+ $Y=1.515 $X2=2.6 $Y2=1.515
r77 32 34 29.0991 $w=3.23e-07 $l=1.95e-07 $layer=POLY_cond $X=2.405 $Y=1.515
+ $X2=2.6 $Y2=1.515
r78 31 32 6.71517 $w=3.23e-07 $l=4.5e-08 $layer=POLY_cond $X=2.36 $Y=1.515
+ $X2=2.405 $Y2=1.515
r79 27 40 0.53602 $w=4.28e-07 $l=2e-08 $layer=LI1_cond $X=3.6 $Y=1.565 $X2=3.62
+ $Y2=1.565
r80 26 27 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.6 $Y2=1.565
r81 25 26 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.12 $Y2=1.565
r82 25 35 1.07204 $w=4.28e-07 $l=4e-08 $layer=LI1_cond $X=2.64 $Y=1.565 $X2=2.6
+ $Y2=1.565
r83 21 42 16.4327 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.755 $Y=1.68
+ $X2=3.755 $Y2=1.515
r84 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.755 $Y=1.68
+ $X2=3.755 $Y2=2.4
r85 17 41 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.71 $Y=1.35
+ $X2=3.71 $Y2=1.515
r86 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.71 $Y=1.35
+ $X2=3.71 $Y2=0.74
r87 13 37 16.4327 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.305 $Y=1.68
+ $X2=3.305 $Y2=1.515
r88 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.305 $Y=1.68
+ $X2=3.305 $Y2=2.4
r89 9 36 16.4327 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.855 $Y=1.68
+ $X2=2.855 $Y2=1.515
r90 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.855 $Y=1.68
+ $X2=2.855 $Y2=2.4
r91 5 32 16.4327 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.405 $Y=1.68
+ $X2=2.405 $Y2=1.515
r92 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.405 $Y=1.68
+ $X2=2.405 $Y2=2.4
r93 1 31 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.36 $Y=1.35
+ $X2=2.36 $Y2=1.515
r94 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.36 $Y=1.35 $X2=2.36
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4_4%B 3 7 11 15 19 23 25 26 27 28 29 30 51
c75 51 0 6.09347e-20 $X=6.135 $Y=1.515
r76 49 51 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6 $Y=1.515
+ $X2=6.135 $Y2=1.515
r77 47 49 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=5.685 $Y=1.515
+ $X2=6 $Y2=1.515
r78 46 47 82.1848 $w=3.3e-07 $l=4.7e-07 $layer=POLY_cond $X=5.215 $Y=1.515
+ $X2=5.685 $Y2=1.515
r79 44 46 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=4.98 $Y=1.515
+ $X2=5.215 $Y2=1.515
r80 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.98
+ $Y=1.515 $X2=4.98 $Y2=1.515
r81 42 44 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=4.765 $Y=1.515
+ $X2=4.98 $Y2=1.515
r82 41 45 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=4.64 $Y=1.565
+ $X2=4.98 $Y2=1.565
r83 40 42 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=4.64 $Y=1.515
+ $X2=4.765 $Y2=1.515
r84 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.64
+ $Y=1.515 $X2=4.64 $Y2=1.515
r85 37 40 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.21 $Y=1.515
+ $X2=4.64 $Y2=1.515
r86 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6 $Y=1.565 $X2=6.48
+ $Y2=1.565
r87 29 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6 $Y=1.515
+ $X2=6 $Y2=1.515
r88 28 29 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.52 $Y=1.565 $X2=6
+ $Y2=1.565
r89 27 28 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.52 $Y2=1.565
r90 27 45 1.60806 $w=4.28e-07 $l=6e-08 $layer=LI1_cond $X=5.04 $Y=1.565 $X2=4.98
+ $Y2=1.565
r91 26 41 2.14408 $w=4.28e-07 $l=8e-08 $layer=LI1_cond $X=4.56 $Y=1.565 $X2=4.64
+ $Y2=1.565
r92 25 26 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=4.56 $Y2=1.565
r93 21 51 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.135 $Y=1.68
+ $X2=6.135 $Y2=1.515
r94 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.135 $Y=1.68
+ $X2=6.135 $Y2=2.4
r95 17 47 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.685 $Y=1.68
+ $X2=5.685 $Y2=1.515
r96 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.685 $Y=1.68
+ $X2=5.685 $Y2=2.4
r97 13 46 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.215 $Y=1.68
+ $X2=5.215 $Y2=1.515
r98 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.215 $Y=1.68
+ $X2=5.215 $Y2=2.4
r99 9 42 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.765 $Y=1.68
+ $X2=4.765 $Y2=1.515
r100 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.765 $Y=1.68
+ $X2=4.765 $Y2=2.4
r101 5 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.64 $Y=1.35
+ $X2=4.64 $Y2=1.515
r102 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.64 $Y=1.35 $X2=4.64
+ $Y2=0.74
r103 1 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.21 $Y=1.35
+ $X2=4.21 $Y2=1.515
r104 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.21 $Y=1.35 $X2=4.21
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4_4%A 3 5 6 9 13 17 21 25 32 33 43 45 50
r76 42 50 3.13269 $w=4.48e-07 $l=8.5e-08 $layer=LI1_cond $X=7.89 $Y=1.405
+ $X2=7.805 $Y2=1.405
r77 41 43 14.2697 $w=3.04e-07 $l=9e-08 $layer=POLY_cond $X=7.89 $Y=1.465
+ $X2=7.98 $Y2=1.465
r78 41 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.89
+ $Y=1.465 $X2=7.89 $Y2=1.465
r79 39 41 48.3586 $w=3.04e-07 $l=3.05e-07 $layer=POLY_cond $X=7.585 $Y=1.465
+ $X2=7.89 $Y2=1.465
r80 36 37 2.37829 $w=3.04e-07 $l=1.5e-08 $layer=POLY_cond $X=7.12 $Y=1.465
+ $X2=7.135 $Y2=1.465
r81 33 45 9.83442 $w=4.48e-07 $l=3.7e-07 $layer=LI1_cond $X=8.4 $Y=1.405
+ $X2=8.03 $Y2=1.405
r82 32 45 2.92375 $w=4.48e-07 $l=1.1e-07 $layer=LI1_cond $X=7.92 $Y=1.405
+ $X2=8.03 $Y2=1.405
r83 32 42 0.797386 $w=4.48e-07 $l=3e-08 $layer=LI1_cond $X=7.92 $Y=1.405
+ $X2=7.89 $Y2=1.405
r84 30 39 59.4572 $w=3.04e-07 $l=3.75e-07 $layer=POLY_cond $X=7.21 $Y=1.465
+ $X2=7.585 $Y2=1.465
r85 30 37 11.8914 $w=3.04e-07 $l=7.5e-08 $layer=POLY_cond $X=7.21 $Y=1.465
+ $X2=7.135 $Y2=1.465
r86 29 50 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=7.21 $Y=1.465
+ $X2=7.805 $Y2=1.465
r87 29 30 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.21
+ $Y=1.465 $X2=7.21 $Y2=1.465
r88 23 43 24.5757 $w=3.04e-07 $l=2.29783e-07 $layer=POLY_cond $X=8.135 $Y=1.63
+ $X2=7.98 $Y2=1.465
r89 23 25 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=8.135 $Y=1.63
+ $X2=8.135 $Y2=2.4
r90 19 43 19.2802 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.98 $Y=1.3
+ $X2=7.98 $Y2=1.465
r91 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.98 $Y=1.3 $X2=7.98
+ $Y2=0.74
r92 15 39 15.0262 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.585 $Y=1.63
+ $X2=7.585 $Y2=1.465
r93 15 17 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=7.585 $Y=1.63
+ $X2=7.585 $Y2=2.4
r94 11 37 15.0262 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.135 $Y=1.63
+ $X2=7.135 $Y2=1.465
r95 11 13 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=7.135 $Y=1.63
+ $X2=7.135 $Y2=2.4
r96 7 36 19.2802 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.12 $Y=1.3 $X2=7.12
+ $Y2=1.465
r97 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.12 $Y=1.3 $X2=7.12
+ $Y2=0.74
r98 5 36 24.2693 $w=3.04e-07 $l=1.21861e-07 $layer=POLY_cond $X=7.045 $Y=1.555
+ $X2=7.12 $Y2=1.465
r99 5 6 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.045 $Y=1.555
+ $X2=6.675 $Y2=1.555
r100 1 6 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.585 $Y=1.63
+ $X2=6.675 $Y2=1.555
r101 1 3 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=6.585 $Y=1.63
+ $X2=6.585 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4_4%A_27_368# 1 2 3 4 5 18 20 21 24 26 28 32 36
+ 38 42 46 48
c59 48 0 6.09347e-20 $X=3.98 $Y=2.115
r60 39 46 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.19 $Y=2.035
+ $X2=3.08 $Y2=2.035
r61 38 48 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.895 $Y=2.035
+ $X2=4.02 $Y2=2.035
r62 38 39 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=3.895 $Y=2.035
+ $X2=3.19 $Y2=2.035
r63 34 46 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.12
+ $X2=3.08 $Y2=2.035
r64 34 36 23.5727 $w=2.18e-07 $l=4.5e-07 $layer=LI1_cond $X=3.08 $Y=2.12
+ $X2=3.08 $Y2=2.57
r65 33 44 3.40825 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=2.265 $Y=2.035
+ $X2=2.18 $Y2=1.97
r66 32 46 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.97 $Y=2.035
+ $X2=3.08 $Y2=2.035
r67 32 33 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.97 $Y=2.035
+ $X2=2.265 $Y2=2.035
r68 29 31 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.18 $Y=2.905
+ $X2=2.18 $Y2=2.4
r69 28 44 3.40825 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.18 $Y=2.12 $X2=2.18
+ $Y2=1.97
r70 28 31 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.18 $Y=2.12
+ $X2=2.18 $Y2=2.4
r71 27 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.395 $Y=2.99
+ $X2=1.27 $Y2=2.99
r72 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.095 $Y=2.99
+ $X2=2.18 $Y2=2.905
r73 26 27 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.095 $Y=2.99
+ $X2=1.395 $Y2=2.99
r74 22 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=2.905
+ $X2=1.27 $Y2=2.99
r75 22 24 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=1.27 $Y=2.905
+ $X2=1.27 $Y2=2.455
r76 20 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.145 $Y=2.99
+ $X2=1.27 $Y2=2.99
r77 20 21 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.145 $Y=2.99
+ $X2=0.445 $Y2=2.99
r78 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.445 $Y2=2.99
r79 16 18 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.28 $Y2=2.455
r80 5 48 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=3.845
+ $Y=1.84 $X2=3.98 $Y2=2.115
r81 4 46 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=2.945
+ $Y=1.84 $X2=3.08 $Y2=2.035
r82 4 36 600 $w=1.7e-07 $l=7.94638e-07 $layer=licon1_PDIFF $count=1 $X=2.945
+ $Y=1.84 $X2=3.08 $Y2=2.57
r83 3 44 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.84 $X2=2.18 $Y2=1.985
r84 3 31 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=2.045
+ $Y=1.84 $X2=2.18 $Y2=2.4
r85 2 24 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.095
+ $Y=1.84 $X2=1.23 $Y2=2.455
r86 1 18 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4_4%Y 1 2 3 4 5 6 20 21 22 25 31 35 37 43 46 48
+ 50 53 56 57 61 63
c102 57 0 1.56424e-19 $X=4.425 $Y=1.07
r103 61 62 1.69739 $w=5.75e-07 $l=8e-08 $layer=LI1_cond $X=7.55 $Y=0.965
+ $X2=7.55 $Y2=1.045
r104 59 61 9.54783 $w=5.75e-07 $l=4.5e-07 $layer=LI1_cond $X=7.55 $Y=0.515
+ $X2=7.55 $Y2=0.965
r105 55 56 10.6082 $w=8.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.495 $Y=0.765
+ $X2=3.59 $Y2=0.765
r106 52 55 13.2577 $w=8.28e-07 $l=9.2e-07 $layer=LI1_cond $X=2.575 $Y=0.765
+ $X2=3.495 $Y2=0.765
r107 52 53 11.617 $w=8.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=0.765
+ $X2=2.41 $Y2=0.765
r108 46 53 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.74 $Y=1.095
+ $X2=2.41 $Y2=1.095
r109 45 46 10.6082 $w=8.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.645 $Y=0.765
+ $X2=1.74 $Y2=0.765
r110 42 45 12.8254 $w=8.28e-07 $l=8.9e-07 $layer=LI1_cond $X=0.755 $Y=0.765
+ $X2=1.645 $Y2=0.765
r111 42 43 11.2567 $w=8.28e-07 $l=1.4e-07 $layer=LI1_cond $X=0.755 $Y=0.765
+ $X2=0.615 $Y2=0.765
r112 40 63 32.8196 $w=2.28e-07 $l=6.55e-07 $layer=LI1_cond $X=0.24 $Y=1.95
+ $X2=0.24 $Y2=1.295
r113 39 63 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.24 $Y=1.18
+ $X2=0.24 $Y2=1.295
r114 38 57 8.61065 $w=1.7e-07 $l=1.77059e-07 $layer=LI1_cond $X=4.59 $Y=1.045
+ $X2=4.425 $Y2=1.07
r115 37 62 8.04321 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=7.24 $Y=1.045
+ $X2=7.55 $Y2=1.045
r116 37 38 172.888 $w=1.68e-07 $l=2.65e-06 $layer=LI1_cond $X=7.24 $Y=1.045
+ $X2=4.59 $Y2=1.045
r117 33 57 0.89609 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.425 $Y=0.96
+ $X2=4.425 $Y2=1.07
r118 33 35 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=4.425 $Y=0.96
+ $X2=4.425 $Y2=0.515
r119 31 57 8.61065 $w=1.7e-07 $l=1.77059e-07 $layer=LI1_cond $X=4.26 $Y=1.095
+ $X2=4.425 $Y2=1.07
r120 31 56 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.26 $Y=1.095
+ $X2=3.59 $Y2=1.095
r121 26 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=2.035
+ $X2=0.78 $Y2=2.035
r122 25 50 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.565 $Y=2.035
+ $X2=1.73 $Y2=2.035
r123 25 26 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.565 $Y=2.035
+ $X2=0.945 $Y2=2.035
r124 22 40 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=2.035
+ $X2=0.24 $Y2=1.95
r125 21 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=2.035
+ $X2=0.78 $Y2=2.035
r126 21 22 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.615 $Y=2.035
+ $X2=0.355 $Y2=2.035
r127 20 39 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.095
+ $X2=0.24 $Y2=1.18
r128 20 43 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.355 $Y=1.095
+ $X2=0.615 $Y2=1.095
r129 6 50 300 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.84 $X2=1.73 $Y2=2.115
r130 5 48 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=0.645
+ $Y=1.84 $X2=0.78 $Y2=2.115
r131 4 61 91 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=2 $X=7.195
+ $Y=0.37 $X2=7.335 $Y2=0.965
r132 4 59 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.195
+ $Y=0.37 $X2=7.335 $Y2=0.515
r133 3 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.285
+ $Y=0.37 $X2=4.425 $Y2=0.515
r134 2 55 60.6667 $w=1.7e-07 $l=1.13018e-06 $layer=licon1_NDIFF $count=3
+ $X=2.435 $Y=0.37 $X2=3.495 $Y2=0.515
r135 2 52 60.6667 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=3
+ $X=2.435 $Y=0.37 $X2=2.575 $Y2=0.515
r136 1 45 60.6667 $w=1.7e-07 $l=1.10011e-06 $layer=licon1_NDIFF $count=3
+ $X=0.615 $Y=0.37 $X2=1.645 $Y2=0.515
r137 1 42 60.6667 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=3
+ $X=0.615 $Y=0.37 $X2=0.755 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4_4%A_499_368# 1 2 3 4 15 17 18 21 23 27 29 33 35
+ 36
c63 18 0 9.97624e-20 $X=2.795 $Y=2.99
r64 31 33 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=5.91 $Y=2.905
+ $X2=5.91 $Y2=2.385
r65 30 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.155 $Y=2.99
+ $X2=4.99 $Y2=2.99
r66 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.745 $Y=2.99
+ $X2=5.91 $Y2=2.905
r67 29 30 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.745 $Y=2.99
+ $X2=5.155 $Y2=2.99
r68 25 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.99 $Y=2.905
+ $X2=4.99 $Y2=2.99
r69 25 27 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=4.99 $Y=2.905
+ $X2=4.99 $Y2=2.385
r70 24 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.695 $Y=2.99
+ $X2=3.53 $Y2=2.99
r71 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.825 $Y=2.99
+ $X2=4.99 $Y2=2.99
r72 23 24 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=4.825 $Y=2.99
+ $X2=3.695 $Y2=2.99
r73 19 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.53 $Y=2.905
+ $X2=3.53 $Y2=2.99
r74 19 21 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=3.53 $Y=2.905
+ $X2=3.53 $Y2=2.375
r75 17 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=2.99
+ $X2=3.53 $Y2=2.99
r76 17 18 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.365 $Y=2.99
+ $X2=2.795 $Y2=2.99
r77 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.63 $Y=2.905
+ $X2=2.795 $Y2=2.99
r78 13 15 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=2.63 $Y=2.905
+ $X2=2.63 $Y2=2.375
r79 4 33 300 $w=1.7e-07 $l=6.08769e-07 $layer=licon1_PDIFF $count=2 $X=5.775
+ $Y=1.84 $X2=5.91 $Y2=2.385
r80 3 27 300 $w=1.7e-07 $l=6.08769e-07 $layer=licon1_PDIFF $count=2 $X=4.855
+ $Y=1.84 $X2=4.99 $Y2=2.385
r81 2 21 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=3.395
+ $Y=1.84 $X2=3.53 $Y2=2.375
r82 1 15 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=2.495
+ $Y=1.84 $X2=2.63 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4_4%A_879_368# 1 2 3 4 5 16 18 20 24 26 30 32 36
+ 38 40 42 47 49 51
r70 40 53 3.0656 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=8.36 $Y=2.12 $X2=8.36
+ $Y2=1.97
r71 40 42 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=8.36 $Y=2.12
+ $X2=8.36 $Y2=2.815
r72 39 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.525 $Y=2.035
+ $X2=7.36 $Y2=2.035
r73 38 53 4.70058 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=8.195 $Y=2.035
+ $X2=8.36 $Y2=1.97
r74 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.195 $Y=2.035
+ $X2=7.525 $Y2=2.035
r75 34 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=2.12 $X2=7.36
+ $Y2=2.035
r76 34 36 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=7.36 $Y=2.12
+ $X2=7.36 $Y2=2.815
r77 33 49 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.525 $Y=2.035
+ $X2=6.39 $Y2=2.035
r78 32 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.195 $Y=2.035
+ $X2=7.36 $Y2=2.035
r79 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.195 $Y=2.035
+ $X2=6.525 $Y2=2.035
r80 28 49 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.39 $Y=2.12
+ $X2=6.39 $Y2=2.035
r81 28 30 13.872 $w=2.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.39 $Y=2.12
+ $X2=6.39 $Y2=2.445
r82 27 47 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=5.56 $Y=2.035
+ $X2=5.45 $Y2=2.035
r83 26 49 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.255 $Y=2.035
+ $X2=6.39 $Y2=2.035
r84 26 27 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.255 $Y=2.035
+ $X2=5.56 $Y2=2.035
r85 22 47 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=5.45 $Y=2.12
+ $X2=5.45 $Y2=2.035
r86 22 24 23.5727 $w=2.18e-07 $l=4.5e-07 $layer=LI1_cond $X=5.45 $Y=2.12
+ $X2=5.45 $Y2=2.57
r87 21 45 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.625 $Y=2.035
+ $X2=4.5 $Y2=2.035
r88 20 47 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=5.34 $Y=2.035
+ $X2=5.45 $Y2=2.035
r89 20 21 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=5.34 $Y=2.035
+ $X2=4.625 $Y2=2.035
r90 16 45 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.5 $Y=2.12 $X2=4.5
+ $Y2=2.035
r91 16 18 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=4.5 $Y=2.12 $X2=4.5
+ $Y2=2.57
r92 5 53 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.225
+ $Y=1.84 $X2=8.36 $Y2=1.985
r93 5 42 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.225
+ $Y=1.84 $X2=8.36 $Y2=2.815
r94 4 51 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=7.225
+ $Y=1.84 $X2=7.36 $Y2=2.035
r95 4 36 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.225
+ $Y=1.84 $X2=7.36 $Y2=2.815
r96 3 49 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=6.225
+ $Y=1.84 $X2=6.36 $Y2=2.035
r97 3 30 300 $w=1.7e-07 $l=6.69104e-07 $layer=licon1_PDIFF $count=2 $X=6.225
+ $Y=1.84 $X2=6.36 $Y2=2.445
r98 2 47 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=5.305
+ $Y=1.84 $X2=5.45 $Y2=2.035
r99 2 24 600 $w=1.7e-07 $l=7.99218e-07 $layer=licon1_PDIFF $count=1 $X=5.305
+ $Y=1.84 $X2=5.45 $Y2=2.57
r100 1 45 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.84 $X2=4.54 $Y2=2.035
r101 1 18 600 $w=1.7e-07 $l=7.99218e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.84 $X2=4.54 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4_4%VPWR 1 2 9 13 16 17 18 27 33 34 37
r80 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r81 34 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r82 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r83 31 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=7.86 $Y2=3.33
r84 31 33 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=8.4 $Y2=3.33
r85 30 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r86 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r87 27 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.695 $Y=3.33
+ $X2=7.86 $Y2=3.33
r88 27 29 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.695 $Y=3.33
+ $X2=7.44 $Y2=3.33
r89 26 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r90 25 26 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r91 21 25 407.102 $w=1.68e-07 $l=6.24e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=6.48 $Y2=3.33
r92 21 22 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r93 18 26 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=6.48 $Y2=3.33
r94 18 22 1.13724 $w=4.9e-07 $l=4.08e-06 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=0.24 $Y2=3.33
r95 16 25 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.695 $Y=3.33
+ $X2=6.48 $Y2=3.33
r96 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.695 $Y=3.33
+ $X2=6.86 $Y2=3.33
r97 15 29 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=7.025 $Y=3.33
+ $X2=7.44 $Y2=3.33
r98 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.025 $Y=3.33
+ $X2=6.86 $Y2=3.33
r99 11 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.86 $Y=3.245
+ $X2=7.86 $Y2=3.33
r100 11 13 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=7.86 $Y=3.245
+ $X2=7.86 $Y2=2.375
r101 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.86 $Y=3.245
+ $X2=6.86 $Y2=3.33
r102 7 9 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=6.86 $Y=3.245
+ $X2=6.86 $Y2=2.375
r103 2 13 300 $w=1.7e-07 $l=6.20645e-07 $layer=licon1_PDIFF $count=2 $X=7.675
+ $Y=1.84 $X2=7.86 $Y2=2.375
r104 1 9 300 $w=1.7e-07 $l=6.20645e-07 $layer=licon1_PDIFF $count=2 $X=6.675
+ $Y=1.84 $X2=6.86 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4_4%VGND 1 2 3 4 5 16 18 22 26 28 29 32 35 36 37
+ 38 39 40 42 64 69 73 82
r69 80 82 11.3568 $w=8.73e-07 $l=1.1e-07 $layer=LI1_cond $X=6.96 $Y=0.352
+ $X2=7.07 $Y2=0.352
r70 80 81 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r71 78 80 0.766857 $w=8.73e-07 $l=5.5e-08 $layer=LI1_cond $X=6.905 $Y=0.352
+ $X2=6.96 $Y2=0.352
r72 76 81 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=6.96
+ $Y2=0
r73 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r74 72 75 2.57943 $w=8.73e-07 $l=1.85e-07 $layer=LI1_cond $X=4.855 $Y=0.352
+ $X2=5.04 $Y2=0.352
r75 72 73 11.1477 $w=8.73e-07 $l=9.5e-08 $layer=LI1_cond $X=4.855 $Y=0.352
+ $X2=4.76 $Y2=0.352
r76 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r77 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r78 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r79 61 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r80 61 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=6.96
+ $Y2=0
r81 60 82 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=7.92 $Y=0 $X2=7.07
+ $Y2=0
r82 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r83 57 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r84 56 73 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=4.76
+ $Y2=0
r85 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r86 53 70 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.16
+ $Y2=0
r87 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r88 50 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=0 $X2=2.075
+ $Y2=0
r89 50 52 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.24 $Y=0 $X2=3.6
+ $Y2=0
r90 49 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r91 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r92 46 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r93 46 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r94 45 48 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r95 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r96 43 66 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r97 43 45 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r98 42 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.91 $Y=0 $X2=2.075
+ $Y2=0
r99 42 48 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.91 $Y=0 $X2=1.68
+ $Y2=0
r100 40 57 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.56 $Y2=0
r101 40 53 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.32 $Y=0 $X2=3.6
+ $Y2=0
r102 38 60 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=8.03 $Y=0 $X2=7.92
+ $Y2=0
r103 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.03 $Y=0 $X2=8.195
+ $Y2=0
r104 37 63 2.87059 $w=1.7e-07 $l=4e-08 $layer=LI1_cond $X=8.36 $Y=0 $X2=8.4
+ $Y2=0
r105 37 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.36 $Y=0 $X2=8.195
+ $Y2=0
r106 35 52 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.6
+ $Y2=0
r107 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.925
+ $Y2=0
r108 34 56 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=4.09 $Y=0 $X2=4.56
+ $Y2=0
r109 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.09 $Y=0 $X2=3.925
+ $Y2=0
r110 30 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.195 $Y=0.085
+ $X2=8.195 $Y2=0
r111 30 32 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.195 $Y=0.085
+ $X2=8.195 $Y2=0.515
r112 29 75 8.296 $w=8.73e-07 $l=5.95e-07 $layer=LI1_cond $X=5.635 $Y=0.352
+ $X2=5.04 $Y2=0.352
r113 28 78 3.79246 $w=8.73e-07 $l=2.72e-07 $layer=LI1_cond $X=6.633 $Y=0.352
+ $X2=6.905 $Y2=0.352
r114 28 29 13.915 $w=8.73e-07 $l=9.98e-07 $layer=LI1_cond $X=6.633 $Y=0.352
+ $X2=5.635 $Y2=0.352
r115 24 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.925 $Y=0.085
+ $X2=3.925 $Y2=0
r116 24 26 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=3.925 $Y=0.085
+ $X2=3.925 $Y2=0.675
r117 20 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=0.085
+ $X2=2.075 $Y2=0
r118 20 22 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=2.075 $Y=0.085
+ $X2=2.075 $Y2=0.675
r119 16 66 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r120 16 18 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.675
r121 5 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.055
+ $Y=0.37 $X2=8.195 $Y2=0.515
r122 4 78 60.6667 $w=1.7e-07 $l=2.31399e-06 $layer=licon1_NDIFF $count=3
+ $X=4.715 $Y=0.37 $X2=6.905 $Y2=0.625
r123 4 72 60.6667 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=3
+ $X=4.715 $Y=0.37 $X2=4.855 $Y2=0.625
r124 3 26 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=3.785
+ $Y=0.37 $X2=3.925 $Y2=0.675
r125 2 22 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.935
+ $Y=0.37 $X2=2.075 $Y2=0.675
r126 1 18 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.675
.ends


* File: sky130_fd_sc_ms__or4bb_1.pxi.spice
* Created: Wed Sep  2 12:29:31 2020
* 
x_PM_SKY130_FD_SC_MS__OR4BB_1%C_N N_C_N_M1005_g N_C_N_M1004_g C_N N_C_N_c_95_n
+ N_C_N_c_96_n PM_SKY130_FD_SC_MS__OR4BB_1%C_N
x_PM_SKY130_FD_SC_MS__OR4BB_1%D_N N_D_N_c_121_n N_D_N_M1003_g N_D_N_M1008_g
+ N_D_N_c_123_n D_N N_D_N_c_125_n PM_SKY130_FD_SC_MS__OR4BB_1%D_N
x_PM_SKY130_FD_SC_MS__OR4BB_1%A_219_424# N_A_219_424#_M1008_d
+ N_A_219_424#_M1003_d N_A_219_424#_c_169_n N_A_219_424#_M1000_g
+ N_A_219_424#_c_170_n N_A_219_424#_M1012_g N_A_219_424#_c_178_n
+ N_A_219_424#_c_171_n N_A_219_424#_c_179_n N_A_219_424#_c_172_n
+ N_A_219_424#_c_173_n N_A_219_424#_c_174_n N_A_219_424#_c_175_n
+ PM_SKY130_FD_SC_MS__OR4BB_1%A_219_424#
x_PM_SKY130_FD_SC_MS__OR4BB_1%A_27_424# N_A_27_424#_M1004_s N_A_27_424#_M1005_s
+ N_A_27_424#_M1002_g N_A_27_424#_M1013_g N_A_27_424#_c_237_n
+ N_A_27_424#_c_238_n N_A_27_424#_c_262_n N_A_27_424#_c_277_n
+ N_A_27_424#_c_244_n N_A_27_424#_c_245_n N_A_27_424#_c_239_n
+ N_A_27_424#_c_240_n N_A_27_424#_c_247_n N_A_27_424#_c_248_n
+ N_A_27_424#_c_241_n PM_SKY130_FD_SC_MS__OR4BB_1%A_27_424#
x_PM_SKY130_FD_SC_MS__OR4BB_1%B N_B_M1001_g N_B_M1010_g B B B B N_B_c_333_n
+ N_B_c_334_n PM_SKY130_FD_SC_MS__OR4BB_1%B
x_PM_SKY130_FD_SC_MS__OR4BB_1%A N_A_M1006_g N_A_M1009_g A N_A_c_371_n
+ N_A_c_372_n PM_SKY130_FD_SC_MS__OR4BB_1%A
x_PM_SKY130_FD_SC_MS__OR4BB_1%A_357_378# N_A_357_378#_M1000_d
+ N_A_357_378#_M1010_d N_A_357_378#_M1012_s N_A_357_378#_M1007_g
+ N_A_357_378#_M1011_g N_A_357_378#_c_411_n N_A_357_378#_c_412_n
+ N_A_357_378#_c_413_n N_A_357_378#_c_414_n N_A_357_378#_c_420_n
+ N_A_357_378#_c_415_n N_A_357_378#_c_416_n N_A_357_378#_c_417_n
+ N_A_357_378#_c_418_n PM_SKY130_FD_SC_MS__OR4BB_1%A_357_378#
x_PM_SKY130_FD_SC_MS__OR4BB_1%VPWR N_VPWR_M1005_d N_VPWR_M1006_d N_VPWR_c_504_n
+ N_VPWR_c_505_n N_VPWR_c_506_n N_VPWR_c_507_n VPWR N_VPWR_c_508_n
+ N_VPWR_c_509_n N_VPWR_c_503_n N_VPWR_c_511_n PM_SKY130_FD_SC_MS__OR4BB_1%VPWR
x_PM_SKY130_FD_SC_MS__OR4BB_1%X N_X_M1011_d N_X_M1007_d N_X_c_555_n N_X_c_556_n
+ N_X_c_552_n X X X PM_SKY130_FD_SC_MS__OR4BB_1%X
x_PM_SKY130_FD_SC_MS__OR4BB_1%VGND N_VGND_M1004_d N_VGND_M1000_s N_VGND_M1013_d
+ N_VGND_M1009_d N_VGND_c_577_n N_VGND_c_578_n N_VGND_c_579_n N_VGND_c_580_n
+ N_VGND_c_581_n N_VGND_c_582_n N_VGND_c_583_n N_VGND_c_584_n N_VGND_c_585_n
+ N_VGND_c_586_n VGND N_VGND_c_587_n N_VGND_c_588_n N_VGND_c_589_n
+ PM_SKY130_FD_SC_MS__OR4BB_1%VGND
cc_1 VNB N_C_N_M1005_g 0.00197312f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_2 VNB N_C_N_M1004_g 0.0429909f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.645
cc_3 VNB N_C_N_c_95_n 0.00450233f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_4 VNB N_C_N_c_96_n 0.0581652f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.465
cc_5 VNB N_D_N_c_121_n 0.0214468f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_6 VNB N_D_N_M1008_g 0.0224232f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_D_N_c_123_n 0.00968085f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_8 VNB D_N 0.00727485f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_9 VNB N_D_N_c_125_n 0.0206515f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_10 VNB N_A_219_424#_c_169_n 0.0197534f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.645
cc_11 VNB N_A_219_424#_c_170_n 0.0737865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_219_424#_c_171_n 0.0015275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_219_424#_c_172_n 0.0143397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_219_424#_c_173_n 0.00934204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_219_424#_c_174_n 0.00350886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_219_424#_c_175_n 0.00104708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_424#_M1002_g 0.00642098f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_18 VNB N_A_27_424#_M1013_g 0.0279099f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_19 VNB N_A_27_424#_c_237_n 0.0266401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_424#_c_238_n 0.00925967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_424#_c_239_n 0.00347813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_424#_c_240_n 0.0327815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_424#_c_241_n 0.0163689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B_M1010_g 0.0368875f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.645
cc_25 VNB N_B_c_333_n 0.0267189f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_26 VNB N_B_c_334_n 0.00217439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_M1009_g 0.036966f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.645
cc_28 VNB N_A_c_371_n 0.0243228f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_29 VNB N_A_c_372_n 0.00381166f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_30 VNB N_A_357_378#_M1007_g 0.00178608f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_31 VNB N_A_357_378#_M1011_g 0.0291041f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.465
cc_32 VNB N_A_357_378#_c_411_n 0.00279725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_357_378#_c_412_n 0.0100047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_357_378#_c_413_n 0.00280455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_357_378#_c_414_n 0.0218818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_357_378#_c_415_n 0.00472238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_357_378#_c_416_n 0.00807754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_357_378#_c_417_n 0.00974512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_357_378#_c_418_n 0.0339301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VPWR_c_503_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_552_n 0.024833f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_42 VNB X 0.0267746f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.465
cc_43 VNB X 0.0144258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_577_n 0.0097033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_578_n 0.00587375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_579_n 0.0058484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_580_n 0.00909064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_581_n 0.0231289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_582_n 0.004633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_583_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_584_n 0.00740817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_585_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_586_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_587_n 0.020271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_588_n 0.279887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_589_n 0.0262945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VPB N_C_N_M1005_g 0.0542902f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_58 VPB N_C_N_c_95_n 0.00793086f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_59 VPB N_D_N_M1003_g 0.0386386f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.3
cc_60 VPB N_D_N_c_123_n 0.0104816f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_61 VPB D_N 0.00287267f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_62 VPB N_A_219_424#_c_170_n 0.0184734f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_219_424#_M1012_g 0.0252172f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_64 VPB N_A_219_424#_c_178_n 0.0179844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_219_424#_c_179_n 0.00386631f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_219_424#_c_175_n 0.00855473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_27_424#_M1002_g 0.021177f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_68 VPB N_A_27_424#_c_238_n 0.00919125f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_27_424#_c_244_n 0.0368694f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_27_424#_c_245_n 0.00259308f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_27_424#_c_239_n 0.00324761f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_27_424#_c_247_n 0.0216643f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_27_424#_c_248_n 0.020611f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_B_M1001_g 0.0242254f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_75 VPB N_B_c_333_n 0.00568825f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_76 VPB N_B_c_334_n 0.00273691f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_M1006_g 0.0255964f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_78 VPB N_A_c_371_n 0.0055319f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_79 VPB N_A_c_372_n 0.00568995f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_80 VPB N_A_357_378#_M1007_g 0.0304722f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_81 VPB N_A_357_378#_c_420_n 0.00239436f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_504_n 0.00635773f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_83 VPB N_VPWR_c_505_n 0.01236f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_84 VPB N_VPWR_c_506_n 0.071143f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_85 VPB N_VPWR_c_507_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_508_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_509_n 0.0216783f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_503_n 0.0914716f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_511_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_X_c_555_n 0.0454029f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_91 VPB N_X_c_556_n 0.0183426f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_X_c_552_n 0.00785975f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_93 N_C_N_c_96_n N_D_N_c_121_n 0.0188536f $X=0.52 $Y=1.465 $X2=0 $Y2=0
cc_94 N_C_N_M1004_g N_D_N_M1008_g 0.0172328f $X=0.52 $Y=0.645 $X2=0 $Y2=0
cc_95 N_C_N_M1005_g N_D_N_c_123_n 0.0188536f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_96 N_C_N_M1004_g D_N 2.57477e-19 $X=0.52 $Y=0.645 $X2=0 $Y2=0
cc_97 N_C_N_M1004_g N_D_N_c_125_n 0.0188536f $X=0.52 $Y=0.645 $X2=0 $Y2=0
cc_98 N_C_N_M1004_g N_A_219_424#_c_172_n 3.64366e-19 $X=0.52 $Y=0.645 $X2=0
+ $Y2=0
cc_99 N_C_N_M1004_g N_A_27_424#_c_237_n 0.012764f $X=0.52 $Y=0.645 $X2=0 $Y2=0
cc_100 N_C_N_M1004_g N_A_27_424#_c_238_n 0.0167165f $X=0.52 $Y=0.645 $X2=0 $Y2=0
cc_101 N_C_N_c_95_n N_A_27_424#_c_238_n 0.0360322f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_102 N_C_N_M1005_g N_A_27_424#_c_247_n 0.0108644f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_103 N_C_N_M1005_g N_A_27_424#_c_248_n 0.0229487f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_104 N_C_N_c_95_n N_A_27_424#_c_248_n 0.0180285f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_105 N_C_N_c_96_n N_A_27_424#_c_248_n 0.00147466f $X=0.52 $Y=1.465 $X2=0 $Y2=0
cc_106 N_C_N_M1004_g N_A_27_424#_c_241_n 0.0195374f $X=0.52 $Y=0.645 $X2=0 $Y2=0
cc_107 N_C_N_c_95_n N_A_27_424#_c_241_n 0.0243771f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_108 N_C_N_c_96_n N_A_27_424#_c_241_n 0.00214727f $X=0.52 $Y=1.465 $X2=0 $Y2=0
cc_109 N_C_N_M1005_g N_VPWR_c_504_n 0.00334717f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_110 N_C_N_M1005_g N_VPWR_c_508_n 0.005209f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_111 N_C_N_M1005_g N_VPWR_c_503_n 0.00540713f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_112 N_C_N_M1004_g N_VGND_c_577_n 0.00592235f $X=0.52 $Y=0.645 $X2=0 $Y2=0
cc_113 N_C_N_M1004_g N_VGND_c_588_n 0.00825053f $X=0.52 $Y=0.645 $X2=0 $Y2=0
cc_114 N_C_N_M1004_g N_VGND_c_589_n 0.00434272f $X=0.52 $Y=0.645 $X2=0 $Y2=0
cc_115 N_D_N_M1008_g N_A_219_424#_c_170_n 4.84394e-19 $X=1.09 $Y=0.645 $X2=0
+ $Y2=0
cc_116 D_N N_A_219_424#_c_170_n 0.00185735f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_117 N_D_N_c_125_n N_A_219_424#_c_170_n 0.0295782f $X=1.13 $Y=1.215 $X2=0
+ $Y2=0
cc_118 N_D_N_M1003_g N_A_219_424#_c_178_n 0.00653743f $X=1.005 $Y=2.54 $X2=0
+ $Y2=0
cc_119 N_D_N_c_123_n N_A_219_424#_c_178_n 0.00103904f $X=1.105 $Y=1.72 $X2=0
+ $Y2=0
cc_120 D_N N_A_219_424#_c_178_n 0.0135506f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_121 N_D_N_c_121_n N_A_219_424#_c_171_n 7.94903e-19 $X=1.105 $Y=1.53 $X2=0
+ $Y2=0
cc_122 N_D_N_M1003_g N_A_219_424#_c_179_n 0.00467887f $X=1.005 $Y=2.54 $X2=0
+ $Y2=0
cc_123 N_D_N_M1008_g N_A_219_424#_c_172_n 0.0100789f $X=1.09 $Y=0.645 $X2=0
+ $Y2=0
cc_124 D_N N_A_219_424#_c_172_n 0.0123892f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_125 N_D_N_c_125_n N_A_219_424#_c_172_n 8.2849e-19 $X=1.13 $Y=1.215 $X2=0
+ $Y2=0
cc_126 D_N N_A_219_424#_c_173_n 0.0568245f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_127 N_D_N_c_125_n N_A_219_424#_c_173_n 7.94903e-19 $X=1.13 $Y=1.215 $X2=0
+ $Y2=0
cc_128 N_D_N_M1008_g N_A_219_424#_c_174_n 0.00479241f $X=1.09 $Y=0.645 $X2=0
+ $Y2=0
cc_129 N_D_N_c_123_n N_A_219_424#_c_175_n 7.94903e-19 $X=1.105 $Y=1.72 $X2=0
+ $Y2=0
cc_130 N_D_N_M1008_g N_A_27_424#_c_237_n 7.35629e-19 $X=1.09 $Y=0.645 $X2=0
+ $Y2=0
cc_131 D_N N_A_27_424#_c_238_n 0.0444641f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_132 N_D_N_c_125_n N_A_27_424#_c_238_n 0.0101911f $X=1.13 $Y=1.215 $X2=0 $Y2=0
cc_133 N_D_N_M1003_g N_A_27_424#_c_262_n 0.017754f $X=1.005 $Y=2.54 $X2=0 $Y2=0
cc_134 N_D_N_c_123_n N_A_27_424#_c_262_n 2.56605e-19 $X=1.105 $Y=1.72 $X2=0
+ $Y2=0
cc_135 D_N N_A_27_424#_c_262_n 0.00380095f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_136 N_D_N_M1003_g N_A_27_424#_c_245_n 0.00400653f $X=1.005 $Y=2.54 $X2=0
+ $Y2=0
cc_137 N_D_N_M1003_g N_A_27_424#_c_247_n 5.42655e-19 $X=1.005 $Y=2.54 $X2=0
+ $Y2=0
cc_138 N_D_N_M1003_g N_A_27_424#_c_248_n 0.00546037f $X=1.005 $Y=2.54 $X2=0
+ $Y2=0
cc_139 N_D_N_M1008_g N_A_27_424#_c_241_n 0.00237818f $X=1.09 $Y=0.645 $X2=0
+ $Y2=0
cc_140 D_N N_A_27_424#_c_241_n 0.00666811f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_141 N_D_N_c_125_n N_A_27_424#_c_241_n 6.66462e-19 $X=1.13 $Y=1.215 $X2=0
+ $Y2=0
cc_142 N_D_N_M1003_g N_VPWR_c_504_n 0.00800896f $X=1.005 $Y=2.54 $X2=0 $Y2=0
cc_143 N_D_N_M1003_g N_VPWR_c_506_n 0.00460063f $X=1.005 $Y=2.54 $X2=0 $Y2=0
cc_144 N_D_N_M1003_g N_VPWR_c_503_n 0.00468499f $X=1.005 $Y=2.54 $X2=0 $Y2=0
cc_145 N_D_N_M1008_g N_VGND_c_577_n 0.00594187f $X=1.09 $Y=0.645 $X2=0 $Y2=0
cc_146 N_D_N_c_125_n N_VGND_c_577_n 0.00206489f $X=1.13 $Y=1.215 $X2=0 $Y2=0
cc_147 N_D_N_M1008_g N_VGND_c_578_n 0.00280116f $X=1.09 $Y=0.645 $X2=0 $Y2=0
cc_148 N_D_N_M1008_g N_VGND_c_581_n 0.00433162f $X=1.09 $Y=0.645 $X2=0 $Y2=0
cc_149 N_D_N_M1008_g N_VGND_c_588_n 0.0082266f $X=1.09 $Y=0.645 $X2=0 $Y2=0
cc_150 N_A_219_424#_c_170_n N_A_27_424#_M1002_g 0.0758432f $X=2.155 $Y=1.7 $X2=0
+ $Y2=0
cc_151 N_A_219_424#_c_169_n N_A_27_424#_M1013_g 0.0187971f $X=2.14 $Y=1.03 $X2=0
+ $Y2=0
cc_152 N_A_219_424#_c_172_n N_A_27_424#_c_237_n 0.00219986f $X=1.57 $Y=0.615
+ $X2=0 $Y2=0
cc_153 N_A_219_424#_c_178_n N_A_27_424#_c_238_n 0.0102899f $X=1.485 $Y=2.015
+ $X2=0 $Y2=0
cc_154 N_A_219_424#_M1003_d N_A_27_424#_c_262_n 0.00486011f $X=1.095 $Y=2.12
+ $X2=0 $Y2=0
cc_155 N_A_219_424#_c_178_n N_A_27_424#_c_262_n 0.0111092f $X=1.485 $Y=2.015
+ $X2=0 $Y2=0
cc_156 N_A_219_424#_M1003_d N_A_27_424#_c_277_n 0.0132011f $X=1.095 $Y=2.12
+ $X2=0 $Y2=0
cc_157 N_A_219_424#_M1003_d N_A_27_424#_c_244_n 0.00942208f $X=1.095 $Y=2.12
+ $X2=0 $Y2=0
cc_158 N_A_219_424#_M1012_g N_A_27_424#_c_244_n 0.0110217f $X=2.155 $Y=2.39
+ $X2=0 $Y2=0
cc_159 N_A_219_424#_M1003_d N_A_27_424#_c_245_n 4.04887e-19 $X=1.095 $Y=2.12
+ $X2=0 $Y2=0
cc_160 N_A_219_424#_c_170_n N_A_27_424#_c_239_n 0.0107976f $X=2.155 $Y=1.7 $X2=0
+ $Y2=0
cc_161 N_A_219_424#_c_170_n N_A_27_424#_c_240_n 0.0207341f $X=2.155 $Y=1.7 $X2=0
+ $Y2=0
cc_162 N_A_219_424#_c_178_n N_A_27_424#_c_248_n 0.00150688f $X=1.485 $Y=2.015
+ $X2=0 $Y2=0
cc_163 N_A_219_424#_c_169_n N_A_357_378#_c_411_n 6.34612e-19 $X=2.14 $Y=1.03
+ $X2=0 $Y2=0
cc_164 N_A_219_424#_c_170_n N_A_357_378#_c_420_n 0.00818071f $X=2.155 $Y=1.7
+ $X2=0 $Y2=0
cc_165 N_A_219_424#_M1012_g N_A_357_378#_c_420_n 0.0245235f $X=2.155 $Y=2.39
+ $X2=0 $Y2=0
cc_166 N_A_219_424#_c_178_n N_A_357_378#_c_420_n 0.0198115f $X=1.485 $Y=2.015
+ $X2=0 $Y2=0
cc_167 N_A_219_424#_c_179_n N_A_357_378#_c_420_n 0.00145426f $X=1.57 $Y=1.89
+ $X2=0 $Y2=0
cc_168 N_A_219_424#_c_175_n N_A_357_378#_c_420_n 0.00516543f $X=1.695 $Y=1.7
+ $X2=0 $Y2=0
cc_169 N_A_219_424#_c_169_n N_A_357_378#_c_415_n 2.37676e-19 $X=2.14 $Y=1.03
+ $X2=0 $Y2=0
cc_170 N_A_219_424#_c_170_n N_A_357_378#_c_415_n 0.0209758f $X=2.155 $Y=1.7
+ $X2=0 $Y2=0
cc_171 N_A_219_424#_M1012_g N_A_357_378#_c_415_n 0.00535413f $X=2.155 $Y=2.39
+ $X2=0 $Y2=0
cc_172 N_A_219_424#_c_179_n N_A_357_378#_c_415_n 0.00614623f $X=1.57 $Y=1.89
+ $X2=0 $Y2=0
cc_173 N_A_219_424#_c_173_n N_A_357_378#_c_415_n 0.0487135f $X=1.74 $Y=1.195
+ $X2=0 $Y2=0
cc_174 N_A_219_424#_c_174_n N_A_357_378#_c_415_n 3.11856e-19 $X=1.695 $Y=1.03
+ $X2=0 $Y2=0
cc_175 N_A_219_424#_c_169_n N_A_357_378#_c_416_n 0.0102787f $X=2.14 $Y=1.03
+ $X2=0 $Y2=0
cc_176 N_A_219_424#_c_172_n N_A_357_378#_c_416_n 0.00128152f $X=1.57 $Y=0.615
+ $X2=0 $Y2=0
cc_177 N_A_219_424#_c_174_n N_A_357_378#_c_416_n 0.00565738f $X=1.695 $Y=1.03
+ $X2=0 $Y2=0
cc_178 N_A_219_424#_M1012_g N_VPWR_c_506_n 9.93465e-19 $X=2.155 $Y=2.39 $X2=0
+ $Y2=0
cc_179 N_A_219_424#_c_172_n N_VGND_c_577_n 0.0184787f $X=1.57 $Y=0.615 $X2=0
+ $Y2=0
cc_180 N_A_219_424#_c_169_n N_VGND_c_578_n 0.0081515f $X=2.14 $Y=1.03 $X2=0
+ $Y2=0
cc_181 N_A_219_424#_c_170_n N_VGND_c_578_n 0.0058001f $X=2.155 $Y=1.7 $X2=0
+ $Y2=0
cc_182 N_A_219_424#_c_172_n N_VGND_c_578_n 0.0274617f $X=1.57 $Y=0.615 $X2=0
+ $Y2=0
cc_183 N_A_219_424#_c_173_n N_VGND_c_578_n 0.00389507f $X=1.74 $Y=1.195 $X2=0
+ $Y2=0
cc_184 N_A_219_424#_c_172_n N_VGND_c_581_n 0.0224005f $X=1.57 $Y=0.615 $X2=0
+ $Y2=0
cc_185 N_A_219_424#_c_169_n N_VGND_c_583_n 0.00429299f $X=2.14 $Y=1.03 $X2=0
+ $Y2=0
cc_186 N_A_219_424#_c_169_n N_VGND_c_588_n 0.00430505f $X=2.14 $Y=1.03 $X2=0
+ $Y2=0
cc_187 N_A_219_424#_c_172_n N_VGND_c_588_n 0.0187278f $X=1.57 $Y=0.615 $X2=0
+ $Y2=0
cc_188 N_A_27_424#_c_244_n N_B_M1001_g 0.00305974f $X=2.425 $Y=2.99 $X2=0 $Y2=0
cc_189 N_A_27_424#_M1013_g N_B_M1010_g 0.0197521f $X=2.625 $Y=0.645 $X2=0 $Y2=0
cc_190 N_A_27_424#_c_239_n N_B_M1010_g 9.42171e-19 $X=2.59 $Y=1.355 $X2=0 $Y2=0
cc_191 N_A_27_424#_c_240_n N_B_M1010_g 0.00587031f $X=2.59 $Y=1.355 $X2=0 $Y2=0
cc_192 N_A_27_424#_M1002_g N_B_c_333_n 0.0569234f $X=2.575 $Y=2.39 $X2=0 $Y2=0
cc_193 N_A_27_424#_c_239_n N_B_c_333_n 0.00961701f $X=2.59 $Y=1.355 $X2=0 $Y2=0
cc_194 N_A_27_424#_c_240_n N_B_c_333_n 0.0103599f $X=2.59 $Y=1.355 $X2=0 $Y2=0
cc_195 N_A_27_424#_M1002_g N_B_c_334_n 0.00152963f $X=2.575 $Y=2.39 $X2=0 $Y2=0
cc_196 N_A_27_424#_c_239_n N_B_c_334_n 0.101728f $X=2.59 $Y=1.355 $X2=0 $Y2=0
cc_197 N_A_27_424#_c_240_n N_B_c_334_n 5.92094e-19 $X=2.59 $Y=1.355 $X2=0 $Y2=0
cc_198 N_A_27_424#_M1013_g N_A_357_378#_c_411_n 0.00835034f $X=2.625 $Y=0.645
+ $X2=0 $Y2=0
cc_199 N_A_27_424#_M1013_g N_A_357_378#_c_412_n 0.00918056f $X=2.625 $Y=0.645
+ $X2=0 $Y2=0
cc_200 N_A_27_424#_c_239_n N_A_357_378#_c_412_n 0.0138033f $X=2.59 $Y=1.355
+ $X2=0 $Y2=0
cc_201 N_A_27_424#_c_240_n N_A_357_378#_c_412_n 3.80672e-19 $X=2.59 $Y=1.355
+ $X2=0 $Y2=0
cc_202 N_A_27_424#_c_262_n N_A_357_378#_c_420_n 0.00602388f $X=1.115 $Y=2.395
+ $X2=0 $Y2=0
cc_203 N_A_27_424#_c_277_n N_A_357_378#_c_420_n 0.00812965f $X=1.2 $Y=2.905
+ $X2=0 $Y2=0
cc_204 N_A_27_424#_c_244_n N_A_357_378#_c_420_n 0.0274179f $X=2.425 $Y=2.99
+ $X2=0 $Y2=0
cc_205 N_A_27_424#_M1002_g N_A_357_378#_c_415_n 0.0016086f $X=2.575 $Y=2.39
+ $X2=0 $Y2=0
cc_206 N_A_27_424#_M1013_g N_A_357_378#_c_415_n 0.00305033f $X=2.625 $Y=0.645
+ $X2=0 $Y2=0
cc_207 N_A_27_424#_c_239_n N_A_357_378#_c_415_n 0.114711f $X=2.59 $Y=1.355 $X2=0
+ $Y2=0
cc_208 N_A_27_424#_c_240_n N_A_357_378#_c_415_n 0.00174446f $X=2.59 $Y=1.355
+ $X2=0 $Y2=0
cc_209 N_A_27_424#_M1013_g N_A_357_378#_c_416_n 0.00303744f $X=2.625 $Y=0.645
+ $X2=0 $Y2=0
cc_210 N_A_27_424#_c_239_n N_A_357_378#_c_416_n 0.0131562f $X=2.59 $Y=1.355
+ $X2=0 $Y2=0
cc_211 N_A_27_424#_c_240_n N_A_357_378#_c_416_n 9.69167e-19 $X=2.59 $Y=1.355
+ $X2=0 $Y2=0
cc_212 N_A_27_424#_c_262_n N_VPWR_M1005_d 0.00301626f $X=1.115 $Y=2.395
+ $X2=-0.19 $Y2=-0.245
cc_213 N_A_27_424#_c_248_n N_VPWR_M1005_d 0.00403508f $X=0.795 $Y=2.29 $X2=-0.19
+ $Y2=-0.245
cc_214 N_A_27_424#_c_245_n N_VPWR_c_504_n 0.0117236f $X=1.285 $Y=2.99 $X2=0
+ $Y2=0
cc_215 N_A_27_424#_c_247_n N_VPWR_c_504_n 0.0131729f $X=0.28 $Y=2.265 $X2=0
+ $Y2=0
cc_216 N_A_27_424#_c_248_n N_VPWR_c_504_n 0.0191275f $X=0.795 $Y=2.29 $X2=0
+ $Y2=0
cc_217 N_A_27_424#_M1002_g N_VPWR_c_506_n 9.92001e-19 $X=2.575 $Y=2.39 $X2=0
+ $Y2=0
cc_218 N_A_27_424#_c_244_n N_VPWR_c_506_n 0.0969628f $X=2.425 $Y=2.99 $X2=0
+ $Y2=0
cc_219 N_A_27_424#_c_245_n N_VPWR_c_506_n 0.0121867f $X=1.285 $Y=2.99 $X2=0
+ $Y2=0
cc_220 N_A_27_424#_c_247_n N_VPWR_c_508_n 0.014231f $X=0.28 $Y=2.265 $X2=0 $Y2=0
cc_221 N_A_27_424#_c_262_n N_VPWR_c_503_n 0.00476311f $X=1.115 $Y=2.395 $X2=0
+ $Y2=0
cc_222 N_A_27_424#_c_244_n N_VPWR_c_503_n 0.0556725f $X=2.425 $Y=2.99 $X2=0
+ $Y2=0
cc_223 N_A_27_424#_c_245_n N_VPWR_c_503_n 0.00660921f $X=1.285 $Y=2.99 $X2=0
+ $Y2=0
cc_224 N_A_27_424#_c_247_n N_VPWR_c_503_n 0.0118508f $X=0.28 $Y=2.265 $X2=0
+ $Y2=0
cc_225 N_A_27_424#_c_248_n N_VPWR_c_503_n 0.00632514f $X=0.795 $Y=2.29 $X2=0
+ $Y2=0
cc_226 N_A_27_424#_c_239_n A_449_378# 0.00936201f $X=2.59 $Y=1.355 $X2=-0.19
+ $Y2=-0.245
cc_227 N_A_27_424#_c_239_n A_533_378# 0.00940914f $X=2.59 $Y=1.355 $X2=-0.19
+ $Y2=-0.245
cc_228 N_A_27_424#_c_237_n N_VGND_c_577_n 0.0173003f $X=0.305 $Y=0.645 $X2=0
+ $Y2=0
cc_229 N_A_27_424#_c_241_n N_VGND_c_577_n 0.0122405f $X=0.71 $Y=1.045 $X2=0
+ $Y2=0
cc_230 N_A_27_424#_M1013_g N_VGND_c_578_n 4.5999e-19 $X=2.625 $Y=0.645 $X2=0
+ $Y2=0
cc_231 N_A_27_424#_M1013_g N_VGND_c_579_n 0.003896f $X=2.625 $Y=0.645 $X2=0
+ $Y2=0
cc_232 N_A_27_424#_M1013_g N_VGND_c_583_n 0.00434272f $X=2.625 $Y=0.645 $X2=0
+ $Y2=0
cc_233 N_A_27_424#_M1013_g N_VGND_c_588_n 0.00448714f $X=2.625 $Y=0.645 $X2=0
+ $Y2=0
cc_234 N_A_27_424#_c_237_n N_VGND_c_588_n 0.0119539f $X=0.305 $Y=0.645 $X2=0
+ $Y2=0
cc_235 N_A_27_424#_c_237_n N_VGND_c_589_n 0.0144497f $X=0.305 $Y=0.645 $X2=0
+ $Y2=0
cc_236 N_B_M1001_g N_A_M1006_g 0.0405557f $X=3.055 $Y=2.39 $X2=0 $Y2=0
cc_237 N_B_c_334_n N_A_M1006_g 0.0133405f $X=3.13 $Y=1.515 $X2=0 $Y2=0
cc_238 N_B_M1010_g N_A_M1009_g 0.0290513f $X=3.19 $Y=0.645 $X2=0 $Y2=0
cc_239 N_B_c_333_n N_A_c_371_n 0.0206935f $X=3.13 $Y=1.515 $X2=0 $Y2=0
cc_240 N_B_c_334_n N_A_c_371_n 3.99347e-19 $X=3.13 $Y=1.515 $X2=0 $Y2=0
cc_241 N_B_M1001_g N_A_c_372_n 2.74716e-19 $X=3.055 $Y=2.39 $X2=0 $Y2=0
cc_242 N_B_c_333_n N_A_c_372_n 0.00188716f $X=3.13 $Y=1.515 $X2=0 $Y2=0
cc_243 N_B_c_334_n N_A_c_372_n 0.0318723f $X=3.13 $Y=1.515 $X2=0 $Y2=0
cc_244 N_B_M1010_g N_A_357_378#_c_411_n 7.77907e-19 $X=3.19 $Y=0.645 $X2=0 $Y2=0
cc_245 N_B_M1010_g N_A_357_378#_c_412_n 0.0122106f $X=3.19 $Y=0.645 $X2=0 $Y2=0
cc_246 N_B_c_333_n N_A_357_378#_c_412_n 0.00107986f $X=3.13 $Y=1.515 $X2=0 $Y2=0
cc_247 N_B_c_334_n N_A_357_378#_c_412_n 0.0153396f $X=3.13 $Y=1.515 $X2=0 $Y2=0
cc_248 N_B_M1010_g N_A_357_378#_c_413_n 0.00267454f $X=3.19 $Y=0.645 $X2=0 $Y2=0
cc_249 N_B_M1010_g N_A_357_378#_c_417_n 0.00501298f $X=3.19 $Y=0.645 $X2=0 $Y2=0
cc_250 N_B_M1001_g N_VPWR_c_506_n 0.00462979f $X=3.055 $Y=2.39 $X2=0 $Y2=0
cc_251 N_B_c_334_n N_VPWR_c_506_n 0.00925382f $X=3.13 $Y=1.515 $X2=0 $Y2=0
cc_252 N_B_M1001_g N_VPWR_c_503_n 0.00628405f $X=3.055 $Y=2.39 $X2=0 $Y2=0
cc_253 N_B_c_334_n N_VPWR_c_503_n 0.0112615f $X=3.13 $Y=1.515 $X2=0 $Y2=0
cc_254 N_B_c_334_n A_629_378# 0.0142703f $X=3.13 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_255 N_B_M1010_g N_VGND_c_579_n 0.00821058f $X=3.19 $Y=0.645 $X2=0 $Y2=0
cc_256 N_B_M1010_g N_VGND_c_585_n 0.00383152f $X=3.19 $Y=0.645 $X2=0 $Y2=0
cc_257 N_B_M1010_g N_VGND_c_588_n 0.0038677f $X=3.19 $Y=0.645 $X2=0 $Y2=0
cc_258 N_A_M1006_g N_A_357_378#_M1007_g 0.0192909f $X=3.595 $Y=2.39 $X2=0 $Y2=0
cc_259 N_A_c_371_n N_A_357_378#_M1007_g 0.0026314f $X=3.67 $Y=1.515 $X2=0 $Y2=0
cc_260 N_A_c_372_n N_A_357_378#_M1007_g 0.00260095f $X=3.67 $Y=1.515 $X2=0 $Y2=0
cc_261 N_A_M1009_g N_A_357_378#_M1011_g 0.0194182f $X=3.69 $Y=0.645 $X2=0 $Y2=0
cc_262 N_A_M1009_g N_A_357_378#_c_413_n 0.00681697f $X=3.69 $Y=0.645 $X2=0 $Y2=0
cc_263 N_A_M1009_g N_A_357_378#_c_414_n 0.0158774f $X=3.69 $Y=0.645 $X2=0 $Y2=0
cc_264 N_A_c_371_n N_A_357_378#_c_414_n 0.00208332f $X=3.67 $Y=1.515 $X2=0 $Y2=0
cc_265 N_A_c_372_n N_A_357_378#_c_414_n 0.0370526f $X=3.67 $Y=1.515 $X2=0 $Y2=0
cc_266 N_A_M1009_g N_A_357_378#_c_417_n 0.00857454f $X=3.69 $Y=0.645 $X2=0 $Y2=0
cc_267 N_A_c_371_n N_A_357_378#_c_417_n 8.60229e-19 $X=3.67 $Y=1.515 $X2=0 $Y2=0
cc_268 N_A_c_372_n N_A_357_378#_c_417_n 0.0131775f $X=3.67 $Y=1.515 $X2=0 $Y2=0
cc_269 N_A_M1009_g N_A_357_378#_c_418_n 0.00204771f $X=3.69 $Y=0.645 $X2=0 $Y2=0
cc_270 N_A_c_371_n N_A_357_378#_c_418_n 0.0175012f $X=3.67 $Y=1.515 $X2=0 $Y2=0
cc_271 N_A_c_372_n N_A_357_378#_c_418_n 3.21988e-19 $X=3.67 $Y=1.515 $X2=0 $Y2=0
cc_272 N_A_M1006_g N_VPWR_c_505_n 0.00939623f $X=3.595 $Y=2.39 $X2=0 $Y2=0
cc_273 N_A_c_371_n N_VPWR_c_505_n 5.67795e-19 $X=3.67 $Y=1.515 $X2=0 $Y2=0
cc_274 N_A_c_372_n N_VPWR_c_505_n 0.0082142f $X=3.67 $Y=1.515 $X2=0 $Y2=0
cc_275 N_A_M1006_g N_VPWR_c_506_n 0.00632934f $X=3.595 $Y=2.39 $X2=0 $Y2=0
cc_276 N_A_M1006_g N_VPWR_c_503_n 0.00628405f $X=3.595 $Y=2.39 $X2=0 $Y2=0
cc_277 N_A_M1006_g N_X_c_556_n 7.82083e-19 $X=3.595 $Y=2.39 $X2=0 $Y2=0
cc_278 N_A_M1009_g X 8.67829e-19 $X=3.69 $Y=0.645 $X2=0 $Y2=0
cc_279 N_A_M1009_g N_VGND_c_579_n 4.70105e-19 $X=3.69 $Y=0.645 $X2=0 $Y2=0
cc_280 N_A_M1009_g N_VGND_c_580_n 0.00509005f $X=3.69 $Y=0.645 $X2=0 $Y2=0
cc_281 N_A_M1009_g N_VGND_c_585_n 0.00434272f $X=3.69 $Y=0.645 $X2=0 $Y2=0
cc_282 N_A_M1009_g N_VGND_c_588_n 0.00822269f $X=3.69 $Y=0.645 $X2=0 $Y2=0
cc_283 N_A_357_378#_M1007_g N_VPWR_c_505_n 0.00448829f $X=4.18 $Y=2.4 $X2=0
+ $Y2=0
cc_284 N_A_357_378#_c_414_n N_VPWR_c_505_n 0.00257846f $X=4.005 $Y=1.095 $X2=0
+ $Y2=0
cc_285 N_A_357_378#_M1007_g N_VPWR_c_509_n 0.005209f $X=4.18 $Y=2.4 $X2=0 $Y2=0
cc_286 N_A_357_378#_M1007_g N_VPWR_c_503_n 0.00990807f $X=4.18 $Y=2.4 $X2=0
+ $Y2=0
cc_287 N_A_357_378#_M1007_g N_X_c_555_n 0.012313f $X=4.18 $Y=2.4 $X2=0 $Y2=0
cc_288 N_A_357_378#_M1007_g N_X_c_556_n 0.004933f $X=4.18 $Y=2.4 $X2=0 $Y2=0
cc_289 N_A_357_378#_c_414_n N_X_c_556_n 0.0103068f $X=4.005 $Y=1.095 $X2=0 $Y2=0
cc_290 N_A_357_378#_c_418_n N_X_c_556_n 8.10431e-19 $X=4.21 $Y=1.465 $X2=0 $Y2=0
cc_291 N_A_357_378#_M1007_g N_X_c_552_n 0.00435745f $X=4.18 $Y=2.4 $X2=0 $Y2=0
cc_292 N_A_357_378#_M1011_g N_X_c_552_n 0.00252147f $X=4.295 $Y=0.74 $X2=0 $Y2=0
cc_293 N_A_357_378#_c_414_n N_X_c_552_n 0.0304153f $X=4.005 $Y=1.095 $X2=0 $Y2=0
cc_294 N_A_357_378#_c_418_n N_X_c_552_n 0.00232633f $X=4.21 $Y=1.465 $X2=0 $Y2=0
cc_295 N_A_357_378#_M1011_g X 0.00957241f $X=4.295 $Y=0.74 $X2=0 $Y2=0
cc_296 N_A_357_378#_M1011_g X 0.00334896f $X=4.295 $Y=0.74 $X2=0 $Y2=0
cc_297 N_A_357_378#_c_414_n X 0.0078079f $X=4.005 $Y=1.095 $X2=0 $Y2=0
cc_298 N_A_357_378#_c_412_n N_VGND_M1013_d 0.00336868f $X=3.31 $Y=0.935 $X2=0
+ $Y2=0
cc_299 N_A_357_378#_c_414_n N_VGND_M1009_d 0.00397172f $X=4.005 $Y=1.095 $X2=0
+ $Y2=0
cc_300 N_A_357_378#_c_411_n N_VGND_c_578_n 0.0126571f $X=2.41 $Y=0.645 $X2=0
+ $Y2=0
cc_301 N_A_357_378#_c_411_n N_VGND_c_579_n 0.0131947f $X=2.41 $Y=0.645 $X2=0
+ $Y2=0
cc_302 N_A_357_378#_c_412_n N_VGND_c_579_n 0.0257202f $X=3.31 $Y=0.935 $X2=0
+ $Y2=0
cc_303 N_A_357_378#_c_413_n N_VGND_c_579_n 0.0135183f $X=3.475 $Y=0.645 $X2=0
+ $Y2=0
cc_304 N_A_357_378#_M1011_g N_VGND_c_580_n 0.00783466f $X=4.295 $Y=0.74 $X2=0
+ $Y2=0
cc_305 N_A_357_378#_c_413_n N_VGND_c_580_n 0.0191765f $X=3.475 $Y=0.645 $X2=0
+ $Y2=0
cc_306 N_A_357_378#_c_414_n N_VGND_c_580_n 0.0274645f $X=4.005 $Y=1.095 $X2=0
+ $Y2=0
cc_307 N_A_357_378#_c_418_n N_VGND_c_580_n 3.94089e-19 $X=4.21 $Y=1.465 $X2=0
+ $Y2=0
cc_308 N_A_357_378#_c_411_n N_VGND_c_583_n 0.0145482f $X=2.41 $Y=0.645 $X2=0
+ $Y2=0
cc_309 N_A_357_378#_c_413_n N_VGND_c_585_n 0.0145639f $X=3.475 $Y=0.645 $X2=0
+ $Y2=0
cc_310 N_A_357_378#_M1011_g N_VGND_c_587_n 0.00434272f $X=4.295 $Y=0.74 $X2=0
+ $Y2=0
cc_311 N_A_357_378#_M1011_g N_VGND_c_588_n 0.00826034f $X=4.295 $Y=0.74 $X2=0
+ $Y2=0
cc_312 N_A_357_378#_c_411_n N_VGND_c_588_n 0.0119922f $X=2.41 $Y=0.645 $X2=0
+ $Y2=0
cc_313 N_A_357_378#_c_412_n N_VGND_c_588_n 0.0111284f $X=3.31 $Y=0.935 $X2=0
+ $Y2=0
cc_314 N_A_357_378#_c_413_n N_VGND_c_588_n 0.0119984f $X=3.475 $Y=0.645 $X2=0
+ $Y2=0
cc_315 N_A_357_378#_c_416_n N_VGND_c_588_n 0.00554827f $X=2.325 $Y=0.935 $X2=0
+ $Y2=0
cc_316 N_VPWR_c_509_n N_X_c_555_n 0.021019f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_317 N_VPWR_c_503_n N_X_c_555_n 0.0173296f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_318 N_VPWR_c_505_n N_X_c_556_n 0.041613f $X=3.905 $Y=2.115 $X2=0 $Y2=0
cc_319 X N_VGND_c_580_n 0.0332442f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_320 X N_VGND_c_587_n 0.0163488f $X=4.475 $Y=0.47 $X2=0 $Y2=0
cc_321 X N_VGND_c_588_n 0.0134757f $X=4.475 $Y=0.47 $X2=0 $Y2=0

* NGSPICE file created from sky130_fd_sc_ms__mux4_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
M1000 VPWR A1 a_540_341# VPB pshort w=1e+06u l=180000u
+  ad=1.87058e+12p pd=1.254e+07u as=3.3e+11p ps=2.66e+06u
M1001 VGND A1 a_450_74# VNB nlowvt w=640000u l=150000u
+  ad=1.2058e+12p pd=9.01e+06u as=4.8e+11p ps=2.78e+06u
M1002 a_766_341# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=3.6525e+11p pd=3.11e+06u as=0p ps=0u
M1003 a_979_74# S0 a_846_74# VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=7.84075e+11p ps=5.5e+06u
M1004 a_1338_125# S1 a_846_74# VNB nlowvt w=640000u l=150000u
+  ad=1.856e+11p pd=1.86e+06u as=0p ps=0u
M1005 a_1068_387# a_27_74# a_846_74# VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=1.155e+12p ps=6.31e+06u
M1006 a_846_74# a_1396_99# a_1338_125# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.2e+11p ps=2.64e+06u
M1007 a_1338_125# S1 a_342_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=5.5e+11p ps=5.1e+06u
M1008 a_846_74# S0 a_766_341# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR S0 a_27_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1010 a_342_74# S0 a_258_341# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=7.8e+11p ps=3.56e+06u
M1011 VGND S1 a_1396_99# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1012 VPWR A3 a_1068_387# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_540_341# a_27_74# a_342_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_264_74# A0 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1015 a_342_74# a_27_74# a_264_74# VNB nlowvt w=640000u l=150000u
+  ad=4.32e+11p pd=3.91e+06u as=0p ps=0u
M1016 VPWR S1 a_1396_99# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.3e+11p ps=2.66e+06u
M1017 X a_1338_125# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1018 X a_1338_125# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.304e+11p pd=2.83e+06u as=0p ps=0u
M1019 a_450_74# S0 a_342_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_258_341# A0 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND S0 a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1022 a_846_74# a_27_74# a_768_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1023 a_768_74# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_342_74# a_1396_99# a_1338_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND A3 a_979_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__einvp_8.spice
* Created: Fri Aug 28 17:34:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__einvp_8.pex.spice"
.subckt sky130_fd_sc_ms__einvp_8  VNB VPB A TE Z VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Z	Z
* TE	TE
* A	A
* VPB	VPB
* VNB	VNB
MM1005 N_A_27_74#_M1005_d N_A_M1005_g N_Z_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75007.2 A=0.111 P=1.78 MULT=1
MM1006 N_A_27_74#_M1006_d N_A_M1006_g N_Z_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75006.8 A=0.111 P=1.78 MULT=1
MM1008 N_A_27_74#_M1006_d N_A_M1008_g N_Z_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75006.3 A=0.111 P=1.78 MULT=1
MM1014 N_A_27_74#_M1014_d N_A_M1014_g N_Z_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75005.8 A=0.111 P=1.78 MULT=1
MM1019 N_A_27_74#_M1014_d N_A_M1019_g N_Z_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.1
+ SB=75005.3 A=0.111 P=1.78 MULT=1
MM1022 N_A_27_74#_M1022_d N_A_M1022_g N_Z_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.6
+ SB=75004.8 A=0.111 P=1.78 MULT=1
MM1028 N_A_27_74#_M1022_d N_A_M1028_g N_Z_M1028_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003.1
+ SB=75004.3 A=0.111 P=1.78 MULT=1
MM1029 N_A_27_74#_M1029_d N_A_M1029_g N_Z_M1028_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.6
+ SB=75003.8 A=0.111 P=1.78 MULT=1
MM1004 N_A_27_74#_M1029_d N_TE_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.1
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1007 N_A_27_74#_M1007_d N_TE_M1007_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75004.6
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1011 N_A_27_74#_M1007_d N_TE_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75005
+ SB=75002.4 A=0.111 P=1.78 MULT=1
MM1015 N_A_27_74#_M1015_d N_TE_M1015_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.4
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1026 N_A_27_74#_M1015_d N_TE_M1026_g N_VGND_M1026_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.9
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1030 N_A_27_74#_M1030_d N_TE_M1030_g N_VGND_M1026_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75006.3
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1031 N_A_27_74#_M1030_d N_TE_M1031_g N_VGND_M1031_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75006.7
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1033 N_A_27_74#_M1033_d N_TE_M1033_g N_VGND_M1031_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75007.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_TE_M1001_g N_A_802_323#_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.2146 PD=2.05 PS=2.06 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_A_27_368#_M1009_d N_A_M1009_g N_Z_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.308 AS=0.1512 PD=2.79 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90006.9 A=0.2016 P=2.6 MULT=1
MM1012 N_A_27_368#_M1012_d N_A_M1012_g N_Z_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90006.5 A=0.2016 P=2.6 MULT=1
MM1016 N_A_27_368#_M1012_d N_A_M1016_g N_Z_M1016_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90006 A=0.2016 P=2.6 MULT=1
MM1017 N_A_27_368#_M1017_d N_A_M1017_g N_Z_M1016_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90005.6 A=0.2016 P=2.6 MULT=1
MM1020 N_A_27_368#_M1017_d N_A_M1020_g N_Z_M1020_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90005.1 A=0.2016 P=2.6 MULT=1
MM1023 N_A_27_368#_M1023_d N_A_M1023_g N_Z_M1020_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.4
+ SB=90004.7 A=0.2016 P=2.6 MULT=1
MM1027 N_A_27_368#_M1023_d N_A_M1027_g N_Z_M1027_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.9
+ SB=90004.2 A=0.2016 P=2.6 MULT=1
MM1032 N_A_27_368#_M1032_d N_A_M1032_g N_Z_M1027_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.3
+ SB=90003.8 A=0.2016 P=2.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_802_323#_M1000_g N_A_27_368#_M1032_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90003.8 SB=90003.3 A=0.2016 P=2.6 MULT=1
MM1002 N_VPWR_M1000_d N_A_802_323#_M1002_g N_A_27_368#_M1002_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90004.2 SB=90002.9 A=0.2016 P=2.6 MULT=1
MM1003 N_VPWR_M1003_d N_A_802_323#_M1003_g N_A_27_368#_M1002_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90004.7 SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1010 N_VPWR_M1003_d N_A_802_323#_M1010_g N_A_27_368#_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90005.1 SB=90002 A=0.2016 P=2.6 MULT=1
MM1013 N_VPWR_M1013_d N_A_802_323#_M1013_g N_A_27_368#_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90005.6 SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1018 N_VPWR_M1013_d N_A_802_323#_M1018_g N_A_27_368#_M1018_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90006
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1021 N_VPWR_M1021_d N_A_802_323#_M1021_g N_A_27_368#_M1018_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90006.5 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1024 N_VPWR_M1021_d N_A_802_323#_M1024_g N_A_27_368#_M1024_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.308 PD=1.39 PS=2.79 NRD=0 NRS=0 M=1 R=6.22222 SA=90006.9
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1025 N_VPWR_M1025_d N_TE_M1025_g N_A_802_323#_M1025_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3024 AS=0.3024 PD=2.78 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX34_noxref VNB VPB NWDIODE A=17.67 P=22.72
*
.include "sky130_fd_sc_ms__einvp_8.pxi.spice"
*
.ends
*
*

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__clkdlyinv5sd3_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__clkdlyinv5sd3_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.264600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.190000 0.730000 1.860000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  0.408100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.830000 0.355000 5.190000 0.755000 ;
        RECT 4.830000 1.900000 5.190000 3.060000 ;
        RECT 4.925000 0.755000 5.190000 1.900000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.280000 0.085000 ;
        RECT 0.585000  0.085000 0.915000 0.650000 ;
        RECT 1.915000  0.085000 2.265000 0.745000 ;
        RECT 4.330000  0.085000 4.660000 0.670000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 5.280000 3.415000 ;
        RECT 0.575000 2.380000 0.905000 3.245000 ;
        RECT 1.915000 1.940000 2.265000 3.245000 ;
        RECT 4.330000 1.900000 4.660000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 0.305000 0.410000 0.820000 ;
      RECT 0.095000 0.820000 1.305000 1.020000 ;
      RECT 0.095000 2.030000 1.305000 2.205000 ;
      RECT 0.095000 2.205000 0.400000 2.725000 ;
      RECT 0.975000 1.020000 1.305000 2.030000 ;
      RECT 1.415000 2.650000 1.745000 2.900000 ;
      RECT 1.475000 0.305000 1.720000 1.140000 ;
      RECT 1.475000 1.140000 2.510000 1.470000 ;
      RECT 1.475000 1.470000 1.745000 2.650000 ;
      RECT 2.800000 0.415000 2.970000 1.220000 ;
      RECT 2.800000 1.220000 4.005000 1.390000 ;
      RECT 2.800000 1.390000 2.970000 2.980000 ;
      RECT 3.370000 0.400000 3.700000 0.880000 ;
      RECT 3.370000 0.880000 4.700000 0.925000 ;
      RECT 3.370000 0.925000 4.755000 1.050000 ;
      RECT 3.415000 1.560000 4.755000 1.730000 ;
      RECT 3.415000 1.730000 3.655000 2.980000 ;
      RECT 4.530000 1.050000 4.755000 1.560000 ;
  END
END sky130_fd_sc_ms__clkdlyinv5sd3_1

* File: sky130_fd_sc_ms__sdfrtp_4.pex.spice
* Created: Wed Sep  2 12:30:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SDFRTP_4%A_27_74# 1 2 7 9 11 14 18 21 24 28 31 33 34
+ 36 37 41
c79 37 0 1.84581e-19 $X=2.53 $Y=1.995
c80 31 0 9.11487e-21 $X=2.375 $Y=2.09
c81 9 0 3.56444e-20 $X=1.485 $Y=0.935
r82 37 47 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.53 $Y=1.995
+ $X2=2.53 $Y2=2.16
r83 36 39 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.54 $Y=1.995
+ $X2=2.54 $Y2=2.09
r84 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.53
+ $Y=1.995 $X2=2.53 $Y2=1.995
r85 32 34 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.09
+ $X2=0.28 $Y2=2.09
r86 31 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=2.09
+ $X2=2.54 $Y2=2.09
r87 31 32 125.914 $w=1.68e-07 $l=1.93e-06 $layer=LI1_cond $X=2.375 $Y=2.09
+ $X2=0.445 $Y2=2.09
r88 29 41 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.975 $Y=1.1 $X2=0.975
+ $Y2=1.01
r89 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.1 $X2=0.975 $Y2=1.1
r90 26 33 0.221902 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=1.1
+ $X2=0.24 $Y2=1.1
r91 26 28 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=0.365 $Y=1.1
+ $X2=0.975 $Y2=1.1
r92 22 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.175
+ $X2=0.28 $Y2=2.09
r93 22 24 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=0.28 $Y=2.175
+ $X2=0.28 $Y2=2.465
r94 21 34 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.2 $Y=2.005
+ $X2=0.28 $Y2=2.09
r95 20 33 7.38875 $w=2.1e-07 $l=1.83916e-07 $layer=LI1_cond $X=0.2 $Y=1.265
+ $X2=0.24 $Y2=1.1
r96 20 21 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.2 $Y=1.265 $X2=0.2
+ $Y2=2.005
r97 16 33 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=0.935
+ $X2=0.24 $Y2=1.1
r98 16 18 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=0.24 $Y=0.935
+ $X2=0.24 $Y2=0.58
r99 14 47 186.581 $w=1.8e-07 $l=4.8e-07 $layer=POLY_cond $X=2.495 $Y=2.64
+ $X2=2.495 $Y2=2.16
r100 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.485 $Y=0.935
+ $X2=1.485 $Y2=0.615
r101 8 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.01
+ $X2=0.975 $Y2=1.01
r102 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.41 $Y=1.01
+ $X2=1.485 $Y2=0.935
r103 7 8 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.41 $Y=1.01 $X2=1.14
+ $Y2=1.01
r104 2 24 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.465
r105 1 18 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_4%SCE 3 7 11 13 15 18 19 20 23 28 29 30 42 51
+ 53
c78 20 0 1.84581e-19 $X=2.405 $Y=1.575
c79 13 0 2.86058e-19 $X=2.7 $Y=1.05
r80 42 51 1.90404 $w=3.43e-07 $l=5.7e-08 $layer=LI1_cond $X=1.623 $Y=1.662
+ $X2=1.68 $Y2=1.662
r81 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.45
+ $Y=1.67 $X2=1.45 $Y2=1.67
r82 36 39 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=0.77 $Y=1.67
+ $X2=1.45 $Y2=1.67
r83 30 53 6.34154 $w=3.43e-07 $l=1.01e-07 $layer=LI1_cond $X=1.694 $Y=1.662
+ $X2=1.795 $Y2=1.662
r84 30 51 0.467658 $w=3.43e-07 $l=1.4e-08 $layer=LI1_cond $X=1.694 $Y=1.662
+ $X2=1.68 $Y2=1.662
r85 30 42 0.467658 $w=3.43e-07 $l=1.4e-08 $layer=LI1_cond $X=1.609 $Y=1.662
+ $X2=1.623 $Y2=1.662
r86 30 40 5.31126 $w=3.43e-07 $l=1.59e-07 $layer=LI1_cond $X=1.609 $Y=1.662
+ $X2=1.45 $Y2=1.662
r87 29 40 8.35104 $w=3.43e-07 $l=2.5e-07 $layer=LI1_cond $X=1.2 $Y=1.662
+ $X2=1.45 $Y2=1.662
r88 28 29 16.034 $w=3.43e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.662 $X2=1.2
+ $Y2=1.662
r89 28 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.77
+ $Y=1.67 $X2=0.77 $Y2=1.67
r90 23 26 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.57 $Y=1.425
+ $X2=2.57 $Y2=1.575
r91 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.53
+ $Y=1.425 $X2=2.53 $Y2=1.425
r92 20 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.405 $Y=1.575
+ $X2=2.57 $Y2=1.575
r93 20 53 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.405 $Y=1.575
+ $X2=1.795 $Y2=1.575
r94 19 39 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=1.535 $Y=1.67
+ $X2=1.45 $Y2=1.67
r95 17 36 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=0.595 $Y=1.67
+ $X2=0.77 $Y2=1.67
r96 17 18 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.595 $Y=1.67
+ $X2=0.505 $Y2=1.67
r97 13 24 74.5963 $w=2.82e-07 $l=4.35172e-07 $layer=POLY_cond $X=2.7 $Y=1.05
+ $X2=2.57 $Y2=1.425
r98 13 15 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.7 $Y=1.05 $X2=2.7
+ $Y2=0.615
r99 9 19 30.0773 $w=3.3e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.625 $Y=1.835
+ $X2=1.535 $Y2=1.67
r100 9 11 312.911 $w=1.8e-07 $l=8.05e-07 $layer=POLY_cond $X=1.625 $Y=1.835
+ $X2=1.625 $Y2=2.64
r101 5 18 34.7346 $w=1.65e-07 $l=1.69926e-07 $layer=POLY_cond $X=0.495 $Y=1.505
+ $X2=0.505 $Y2=1.67
r102 5 7 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.495 $Y=1.505
+ $X2=0.495 $Y2=0.58
r103 1 18 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.835
+ $X2=0.505 $Y2=1.67
r104 1 3 312.911 $w=1.8e-07 $l=8.05e-07 $layer=POLY_cond $X=0.505 $Y=1.835
+ $X2=0.505 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_4%D 3 6 8 11 12 13
r42 11 14 40.9207 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.952 $Y=1.1
+ $X2=1.952 $Y2=1.265
r43 11 13 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.952 $Y=1.1
+ $X2=1.952 $Y2=0.935
r44 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.1 $X2=1.935 $Y2=1.1
r45 8 12 6.7033 $w=4.53e-07 $l=2.55e-07 $layer=LI1_cond $X=1.68 $Y=1.037
+ $X2=1.935 $Y2=1.037
r46 6 14 534.476 $w=1.8e-07 $l=1.375e-06 $layer=POLY_cond $X=2.045 $Y=2.64
+ $X2=2.045 $Y2=1.265
r47 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2 $Y=0.615 $X2=2
+ $Y2=0.935
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_4%SCD 3 6 10 11 12 13 17
c41 12 0 1.64252e-19 $X=3.12 $Y=1.665
c42 11 0 1.34001e-19 $X=3.07 $Y=2.245
r43 12 13 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.11 $Y=1.605
+ $X2=3.11 $Y2=2.035
r44 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.07
+ $Y=1.605 $X2=3.07 $Y2=1.605
r45 10 17 83.0591 $w=3.3e-07 $l=4.75e-07 $layer=POLY_cond $X=3.07 $Y=2.08
+ $X2=3.07 $Y2=1.605
r46 10 11 35.4289 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.07 $Y=2.08
+ $X2=3.07 $Y2=2.245
r47 9 17 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.07 $Y=1.44
+ $X2=3.07 $Y2=1.605
r48 6 9 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=3.06 $Y=0.615
+ $X2=3.06 $Y2=1.44
r49 3 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.055 $Y=2.64
+ $X2=3.055 $Y2=2.245
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_4%CLK 1 3 6 8
c53 1 0 1.55667e-19 $X=4.595 $Y=1.41
r54 11 12 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.99
+ $Y=1.445 $X2=3.99 $Y2=1.445
r55 8 12 3.0298 $w=6.04e-07 $l=1.5e-07 $layer=LI1_cond $X=4.212 $Y=1.295
+ $X2=4.212 $Y2=1.445
r56 4 14 16.7902 $w=1.8e-07 $l=2.48e-07 $layer=POLY_cond $X=4.645 $Y=1.775
+ $X2=4.645 $Y2=1.527
r57 4 6 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.645 $Y=1.775
+ $X2=4.645 $Y2=2.495
r58 1 14 7.34756 $w=3.28e-07 $l=5e-08 $layer=POLY_cond $X=4.595 $Y=1.527
+ $X2=4.645 $Y2=1.527
r59 1 11 88.9055 $w=3.28e-07 $l=6.05e-07 $layer=POLY_cond $X=4.595 $Y=1.527
+ $X2=3.99 $Y2=1.527
r60 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.595 $Y=1.41
+ $X2=4.595 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_4%A_1037_387# 1 2 9 11 15 17 19 20 21 24 29
+ 31 32 33 34 36 39 42 43 44 46 48 49 51 52 57 58 66 67 69
c226 69 0 1.684e-19 $X=6.065 $Y=1.66
c227 67 0 1.40436e-19 $X=9.33 $Y=1.07
c228 66 0 1.39722e-19 $X=9.25 $Y=1.07
c229 57 0 4.31597e-20 $X=5.412 $Y=1.275
c230 15 0 8.28381e-20 $X=6.52 $Y=0.9
r231 66 75 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.25 $Y=1.07 $X2=9.25
+ $Y2=1.16
r232 65 67 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=9.25 $Y=1.07 $X2=9.33
+ $Y2=1.07
r233 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.25
+ $Y=1.07 $X2=9.25 $Y2=1.07
r234 62 65 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.91 $Y=1.07
+ $X2=9.25 $Y2=1.07
r235 58 60 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=7.14 $Y=0.415
+ $X2=7.14 $Y2=0.665
r236 52 79 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.79 $Y=2.215
+ $X2=9.79 $Y2=2.38
r237 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.79
+ $Y=2.215 $X2=9.79 $Y2=2.215
r238 49 51 13.7196 $w=3.13e-07 $l=3.75e-07 $layer=LI1_cond $X=9.415 $Y=2.222
+ $X2=9.79 $Y2=2.222
r239 48 49 7.64049 $w=3.15e-07 $l=1.94921e-07 $layer=LI1_cond $X=9.33 $Y=2.065
+ $X2=9.415 $Y2=2.222
r240 47 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.33 $Y=1.235
+ $X2=9.33 $Y2=1.07
r241 47 48 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=9.33 $Y=1.235
+ $X2=9.33 $Y2=2.065
r242 46 62 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.91 $Y=0.905
+ $X2=8.91 $Y2=1.07
r243 45 46 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=8.91 $Y=0.425
+ $X2=8.91 $Y2=0.905
r244 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.825 $Y=0.34
+ $X2=8.91 $Y2=0.425
r245 43 44 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=8.825 $Y=0.34
+ $X2=8.1 $Y2=0.34
r246 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.015 $Y=0.425
+ $X2=8.1 $Y2=0.34
r247 41 42 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=8.015 $Y=0.425
+ $X2=8.015 $Y2=0.58
r248 40 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.225 $Y=0.665
+ $X2=7.14 $Y2=0.665
r249 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.93 $Y=0.665
+ $X2=8.015 $Y2=0.58
r250 39 40 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=7.93 $Y=0.665
+ $X2=7.225 $Y2=0.665
r251 37 72 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.065 $Y=1.75
+ $X2=6.065 $Y2=1.915
r252 37 69 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.065 $Y=1.75
+ $X2=6.065 $Y2=1.66
r253 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.065
+ $Y=1.75 $X2=6.065 $Y2=1.75
r254 34 56 13.4746 $w=3.35e-07 $l=5.17214e-07 $layer=LI1_cond $X=5.655 $Y=1.75
+ $X2=5.302 $Y2=2.12
r255 34 36 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=5.655 $Y=1.75
+ $X2=6.065 $Y2=1.75
r256 32 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.055 $Y=0.415
+ $X2=7.14 $Y2=0.415
r257 32 33 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=7.055 $Y=0.415
+ $X2=5.62 $Y2=0.415
r258 31 34 8.96243 $w=3.35e-07 $l=2.16852e-07 $layer=LI1_cond $X=5.535 $Y=1.585
+ $X2=5.655 $Y2=1.75
r259 31 57 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.535 $Y=1.585
+ $X2=5.535 $Y2=1.275
r260 27 57 9.87967 $w=4.13e-07 $l=2.07e-07 $layer=LI1_cond $X=5.412 $Y=1.068
+ $X2=5.412 $Y2=1.275
r261 27 29 9.10847 $w=4.13e-07 $l=3.28e-07 $layer=LI1_cond $X=5.412 $Y=1.068
+ $X2=5.412 $Y2=0.74
r262 26 33 8.50155 $w=1.7e-07 $l=2.46868e-07 $layer=LI1_cond $X=5.412 $Y=0.5
+ $X2=5.62 $Y2=0.415
r263 26 29 6.66473 $w=4.13e-07 $l=2.4e-07 $layer=LI1_cond $X=5.412 $Y=0.5
+ $X2=5.412 $Y2=0.74
r264 24 79 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=9.835 $Y=2.75
+ $X2=9.835 $Y2=2.38
r265 20 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.085 $Y=1.16
+ $X2=9.25 $Y2=1.16
r266 20 21 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=9.085 $Y=1.16
+ $X2=8.725 $Y2=1.16
r267 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.65 $Y=1.085
+ $X2=8.725 $Y2=1.16
r268 17 19 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.65 $Y=1.085
+ $X2=8.65 $Y2=0.69
r269 13 15 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=6.52 $Y=1.585
+ $X2=6.52 $Y2=0.9
r270 12 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.23 $Y=1.66
+ $X2=6.065 $Y2=1.66
r271 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.445 $Y=1.66
+ $X2=6.52 $Y2=1.585
r272 11 12 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=6.445 $Y=1.66
+ $X2=6.23 $Y2=1.66
r273 9 72 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=6.135 $Y=2.525
+ $X2=6.135 $Y2=1.915
r274 2 56 600 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=1 $X=5.185
+ $Y=1.935 $X2=5.32 $Y2=2.12
r275 1 29 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.22
+ $Y=0.595 $X2=5.355 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_4%A_1367_112# 1 2 9 13 17 18 21 23 24 26 32
+ 33
c103 33 0 2.99465e-19 $X=8.57 $Y=0.842
c104 21 0 1.09068e-19 $X=7.325 $Y=1.005
c105 17 0 2.34069e-19 $X=7.19 $Y=1.78
c106 9 0 1.59809e-19 $X=6.91 $Y=0.9
r107 39 41 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=6.91 $Y=1.78
+ $X2=7.025 $Y2=1.78
r108 31 33 3.26203 $w=4.93e-07 $l=1.35e-07 $layer=LI1_cond $X=8.435 $Y=0.842
+ $X2=8.57 $Y2=0.842
r109 31 32 9.48656 $w=4.93e-07 $l=1.65e-07 $layer=LI1_cond $X=8.435 $Y=0.842
+ $X2=8.27 $Y2=0.842
r110 26 28 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=8.9 $Y=1.88 $X2=8.9
+ $Y2=2.59
r111 24 35 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.9 $Y=1.49
+ $X2=8.57 $Y2=1.49
r112 24 26 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=8.9 $Y=1.575
+ $X2=8.9 $Y2=1.88
r113 23 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.57 $Y=1.405
+ $X2=8.57 $Y2=1.49
r114 22 33 7.09362 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=8.57 $Y=1.09
+ $X2=8.57 $Y2=0.842
r115 22 23 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.57 $Y=1.09
+ $X2=8.57 $Y2=1.405
r116 21 32 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=7.325 $Y=1.005
+ $X2=8.27 $Y2=1.005
r117 18 41 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.19 $Y=1.78
+ $X2=7.025 $Y2=1.78
r118 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.19
+ $Y=1.78 $X2=7.19 $Y2=1.78
r119 15 21 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=7.19 $Y=1.09
+ $X2=7.325 $Y2=1.005
r120 15 17 29.4513 $w=2.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.19 $Y=1.09
+ $X2=7.19 $Y2=1.78
r121 11 41 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.025 $Y=1.945
+ $X2=7.025 $Y2=1.78
r122 11 13 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=7.025 $Y=1.945
+ $X2=7.025 $Y2=2.525
r123 7 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.91 $Y=1.615
+ $X2=6.91 $Y2=1.78
r124 7 9 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=6.91 $Y=1.615
+ $X2=6.91 $Y2=0.9
r125 2 28 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=8.765
+ $Y=1.735 $X2=8.9 $Y2=2.59
r126 2 26 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.765
+ $Y=1.735 $X2=8.9 $Y2=1.88
r127 1 31 182 $w=1.7e-07 $l=5.24404e-07 $layer=licon1_NDIFF $count=1 $X=8.25
+ $Y=0.37 $X2=8.435 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_4%RESET_B 4 7 8 9 10 11 15 16 17 19 22 26 30
+ 34 35 36 37 38 45 46 50 55 62 63
c215 8 0 1.09068e-19 $X=7.225 $Y=0.18
c216 4 0 1.46183e-19 $X=3.54 $Y=0.615
r217 61 63 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=10.75 $Y=1.985
+ $X2=10.94 $Y2=1.985
r218 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.75
+ $Y=1.985 $X2=10.75 $Y2=1.985
r219 58 61 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=10.63 $Y=1.985
+ $X2=10.75 $Y2=1.985
r220 53 55 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=7.665 $Y=1.985
+ $X2=7.98 $Y2=1.985
r221 51 53 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=7.66 $Y=1.985
+ $X2=7.665 $Y2=1.985
r222 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.995 $X2=3.95 $Y2=1.995
r223 46 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=2.035
+ $X2=10.8 $Y2=2.035
r224 45 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.98
+ $Y=1.985 $X2=7.98 $Y2=1.985
r225 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r226 40 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=2.035
+ $X2=4.08 $Y2=2.035
r227 38 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.065 $Y=2.035
+ $X2=7.92 $Y2=2.035
r228 37 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=10.8 $Y2=2.035
r229 37 38 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=8.065 $Y2=2.035
r230 36 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=2.035
+ $X2=4.08 $Y2=2.035
r231 35 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r232 35 36 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=4.225 $Y2=2.035
r233 28 63 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.94 $Y=2.15
+ $X2=10.94 $Y2=1.985
r234 28 30 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=10.94 $Y=2.15
+ $X2=10.94 $Y2=2.75
r235 24 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.63 $Y=1.82
+ $X2=10.63 $Y2=1.985
r236 24 26 635.83 $w=1.5e-07 $l=1.24e-06 $layer=POLY_cond $X=10.63 $Y=1.82
+ $X2=10.63 $Y2=0.58
r237 20 53 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.665 $Y=2.15
+ $X2=7.665 $Y2=1.985
r238 20 22 145.766 $w=1.8e-07 $l=3.75e-07 $layer=POLY_cond $X=7.665 $Y=2.15
+ $X2=7.665 $Y2=2.525
r239 19 51 18.2676 $w=1.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.66 $Y=1.82
+ $X2=7.66 $Y2=1.985
r240 18 19 205.061 $w=1.7e-07 $l=4.85e-07 $layer=POLY_cond $X=7.66 $Y=1.335
+ $X2=7.66 $Y2=1.82
r241 16 18 27.0678 $w=1.5e-07 $l=1.16619e-07 $layer=POLY_cond $X=7.575 $Y=1.26
+ $X2=7.66 $Y2=1.335
r242 16 17 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=7.575 $Y=1.26
+ $X2=7.375 $Y2=1.26
r243 13 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.3 $Y=1.185
+ $X2=7.375 $Y2=1.26
r244 13 15 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.3 $Y=1.185
+ $X2=7.3 $Y2=0.9
r245 12 15 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=7.3 $Y=0.255
+ $X2=7.3 $Y2=0.9
r246 11 34 67.0835 $w=2.5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.59 $Y=1.995
+ $X2=3.59 $Y2=2.245
r247 11 33 50.8559 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.59 $Y=1.995
+ $X2=3.59 $Y2=1.83
r248 10 49 2.92121 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.93 $Y=1.995
+ $X2=3.95 $Y2=1.995
r249 10 11 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=3.93 $Y=1.995
+ $X2=3.715 $Y2=1.995
r250 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.225 $Y=0.18
+ $X2=7.3 $Y2=0.255
r251 8 9 1851.09 $w=1.5e-07 $l=3.61e-06 $layer=POLY_cond $X=7.225 $Y=0.18
+ $X2=3.615 $Y2=0.18
r252 7 34 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.625 $Y=2.64
+ $X2=3.625 $Y2=2.245
r253 4 33 623.011 $w=1.5e-07 $l=1.215e-06 $layer=POLY_cond $X=3.54 $Y=0.615
+ $X2=3.54 $Y2=1.83
r254 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.54 $Y=0.255
+ $X2=3.615 $Y2=0.18
r255 1 4 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.54 $Y=0.255
+ $X2=3.54 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_4%A_1233_138# 1 2 3 12 14 18 20 24 27 28 31
+ 32 34 35 38 42
c130 35 0 7.6904e-20 $X=8.15 $Y=1.41
c131 24 0 5.85006e-21 $X=6.715 $Y=0.99
c132 12 0 3.00719e-20 $X=8.175 $Y=0.74
r133 38 40 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=6.305 $Y=0.87
+ $X2=6.305 $Y2=0.99
r134 35 48 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=8.15 $Y=1.41
+ $X2=8.15 $Y2=1.52
r135 35 47 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.15 $Y=1.41
+ $X2=8.15 $Y2=1.245
r136 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.15
+ $Y=1.41 $X2=8.15 $Y2=1.41
r137 32 34 17.744 $w=3.13e-07 $l=4.85e-07 $layer=LI1_cond $X=7.665 $Y=1.417
+ $X2=8.15 $Y2=1.417
r138 31 45 11.6012 $w=3.26e-07 $l=4.04191e-07 $layer=LI1_cond $X=7.58 $Y=2.32
+ $X2=7.89 $Y2=2.537
r139 30 32 7.64049 $w=3.15e-07 $l=1.95944e-07 $layer=LI1_cond $X=7.58 $Y=1.575
+ $X2=7.665 $Y2=1.417
r140 30 31 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=7.58 $Y=1.575
+ $X2=7.58 $Y2=2.32
r141 29 42 3.70735 $w=2.5e-07 $l=1.69245e-07 $layer=LI1_cond $X=6.885 $Y=2.405
+ $X2=6.8 $Y2=2.537
r142 28 31 5.9625 $w=3.26e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.495 $Y=2.405
+ $X2=7.58 $Y2=2.32
r143 28 29 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.495 $Y=2.405
+ $X2=6.885 $Y2=2.405
r144 27 42 2.76166 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=6.8 $Y=2.32 $X2=6.8
+ $Y2=2.537
r145 26 27 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=6.8 $Y=1.075
+ $X2=6.8 $Y2=2.32
r146 25 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.47 $Y=0.99
+ $X2=6.305 $Y2=0.99
r147 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.715 $Y=0.99
+ $X2=6.8 $Y2=1.075
r148 24 25 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.715 $Y=0.99
+ $X2=6.47 $Y2=0.99
r149 20 42 3.70735 $w=2.5e-07 $l=1.08305e-07 $layer=LI1_cond $X=6.715 $Y=2.59
+ $X2=6.8 $Y2=2.537
r150 20 22 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.715 $Y=2.59
+ $X2=6.41 $Y2=2.59
r151 16 18 248.774 $w=1.8e-07 $l=6.4e-07 $layer=POLY_cond $X=8.675 $Y=1.595
+ $X2=8.675 $Y2=2.235
r152 15 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.315 $Y=1.52
+ $X2=8.15 $Y2=1.52
r153 14 16 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.585 $Y=1.52
+ $X2=8.675 $Y2=1.595
r154 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=8.585 $Y=1.52
+ $X2=8.315 $Y2=1.52
r155 12 47 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=8.175 $Y=0.74
+ $X2=8.175 $Y2=1.245
r156 3 45 600 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_PDIFF $count=1 $X=7.755
+ $Y=2.315 $X2=7.89 $Y2=2.535
r157 2 22 600 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=1 $X=6.225
+ $Y=2.315 $X2=6.41 $Y2=2.59
r158 1 38 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=6.165
+ $Y=0.69 $X2=6.305 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_4%A_834_93# 1 2 9 13 14 16 17 18 19 20 22 24
+ 27 29 34 35 36 39 43 45 46 47 49 51 55 58 64 67 68
c189 67 0 1.24672e-19 $X=5.14 $Y=1.502
c190 64 0 3.92595e-20 $X=5.14 $Y=1.61
c191 51 0 1.21102e-19 $X=4.895 $Y=1.945
c192 35 0 1.10364e-19 $X=9.625 $Y=1.585
c193 22 0 5.85006e-21 $X=6.09 $Y=1.225
r194 67 68 33.4466 $w=3.3e-07 $l=9.2e-08 $layer=POLY_cond $X=5.14 $Y=1.502
+ $X2=5.14 $Y2=1.41
r195 65 70 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.14 $Y=1.61
+ $X2=5.14 $Y2=1.775
r196 65 67 18.885 $w=3.3e-07 $l=1.08e-07 $layer=POLY_cond $X=5.14 $Y=1.61
+ $X2=5.14 $Y2=1.502
r197 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.14
+ $Y=1.61 $X2=5.14 $Y2=1.61
r198 58 59 21.5428 $w=2.69e-07 $l=4.75e-07 $layer=LI1_cond $X=4.42 $Y=2.115
+ $X2=4.895 $Y2=2.115
r199 53 55 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=4.32 $Y=0.625
+ $X2=4.45 $Y2=0.625
r200 51 59 3.42229 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.895 $Y=1.945
+ $X2=4.895 $Y2=2.115
r201 50 60 5.0588 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=4.895 $Y=1.8
+ $X2=4.895 $Y2=1.622
r202 50 51 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.895 $Y=1.8
+ $X2=4.895 $Y2=1.945
r203 49 64 7.30422 $w=3.53e-07 $l=2.25e-07 $layer=LI1_cond $X=4.915 $Y=1.622
+ $X2=5.14 $Y2=1.622
r204 49 60 0.649264 $w=3.53e-07 $l=2e-08 $layer=LI1_cond $X=4.915 $Y=1.622
+ $X2=4.895 $Y2=1.622
r205 48 49 18.7489 $w=2.08e-07 $l=3.55e-07 $layer=LI1_cond $X=4.915 $Y=1.09
+ $X2=4.915 $Y2=1.445
r206 46 48 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=4.81 $Y=1.005
+ $X2=4.915 $Y2=1.09
r207 46 47 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.81 $Y=1.005
+ $X2=4.535 $Y2=1.005
r208 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.45 $Y=0.92
+ $X2=4.535 $Y2=1.005
r209 44 55 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.45 $Y=0.75
+ $X2=4.45 $Y2=0.625
r210 44 45 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.45 $Y=0.75
+ $X2=4.45 $Y2=0.92
r211 37 39 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=9.7 $Y=1.51 $X2=9.7
+ $Y2=0.58
r212 35 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.625 $Y=1.585
+ $X2=9.7 $Y2=1.51
r213 35 36 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=9.625 $Y=1.585
+ $X2=9.215 $Y2=1.585
r214 32 34 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=9.125 $Y=3.075
+ $X2=9.125 $Y2=2.235
r215 31 36 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=9.125 $Y=1.66
+ $X2=9.215 $Y2=1.585
r216 31 34 223.508 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.125 $Y=1.66
+ $X2=9.125 $Y2=2.235
r217 30 43 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.725 $Y=3.15
+ $X2=6.635 $Y2=3.15
r218 29 32 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=9.035 $Y=3.15
+ $X2=9.125 $Y2=3.075
r219 29 30 1184.49 $w=1.5e-07 $l=2.31e-06 $layer=POLY_cond $X=9.035 $Y=3.15
+ $X2=6.725 $Y2=3.15
r220 25 43 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=6.635 $Y=3.075
+ $X2=6.635 $Y2=3.15
r221 25 27 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=6.635 $Y=3.075
+ $X2=6.635 $Y2=2.525
r222 22 24 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=6.09 $Y=1.225
+ $X2=6.09 $Y2=0.9
r223 21 41 4.37345 $w=1.5e-07 $l=8.8e-08 $layer=POLY_cond $X=5.715 $Y=1.3
+ $X2=5.627 $Y2=1.3
r224 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.015 $Y=1.3
+ $X2=6.09 $Y2=1.225
r225 20 21 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=6.015 $Y=1.3 $X2=5.715
+ $Y2=1.3
r226 18 43 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.545 $Y=3.15
+ $X2=6.635 $Y2=3.15
r227 18 19 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=6.545 $Y=3.15
+ $X2=5.69 $Y2=3.15
r228 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.615 $Y=3.075
+ $X2=5.69 $Y2=3.15
r229 16 17 758.894 $w=1.5e-07 $l=1.48e-06 $layer=POLY_cond $X=5.615 $Y=1.595
+ $X2=5.615 $Y2=3.075
r230 15 67 16.3672 $w=1.85e-07 $l=1.65e-07 $layer=POLY_cond $X=5.305 $Y=1.502
+ $X2=5.14 $Y2=1.502
r231 14 16 28.2677 $w=1.6e-07 $l=9.8818e-08 $layer=POLY_cond $X=5.627 $Y=1.502
+ $X2=5.615 $Y2=1.595
r232 14 41 60.8525 $w=1.6e-07 $l=2.02e-07 $layer=POLY_cond $X=5.627 $Y=1.502
+ $X2=5.627 $Y2=1.3
r233 14 15 86.8144 $w=1.85e-07 $l=2.35e-07 $layer=POLY_cond $X=5.54 $Y=1.502
+ $X2=5.305 $Y2=1.502
r234 13 68 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.145 $Y=0.965
+ $X2=5.145 $Y2=1.41
r235 9 70 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.095 $Y=2.495
+ $X2=5.095 $Y2=1.775
r236 2 58 600 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=4.275
+ $Y=1.935 $X2=4.42 $Y2=2.12
r237 1 53 182 $w=1.7e-07 $l=2.64575e-07 $layer=licon1_NDIFF $count=1 $X=4.17
+ $Y=0.465 $X2=4.32 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_4%A_2003_48# 1 2 9 13 15 17 24 26 27 32 33 36
c85 24 0 1.05829e-19 $X=11.5 $Y=1.385
r86 35 36 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.245 $Y=1.47
+ $X2=11.5 $Y2=1.47
r87 32 33 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=11.165 $Y=2.75
+ $X2=11.165 $Y2=2.52
r88 27 40 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.18 $Y=1.39
+ $X2=10.18 $Y2=1.555
r89 27 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.18 $Y=1.39
+ $X2=10.18 $Y2=1.225
r90 26 29 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=10.18 $Y=1.39 $X2=10.18
+ $Y2=1.47
r91 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.18
+ $Y=1.39 $X2=10.18 $Y2=1.39
r92 24 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.5 $Y=1.385
+ $X2=11.5 $Y2=1.47
r93 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=11.5 $Y=0.715
+ $X2=11.5 $Y2=1.385
r94 21 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.245 $Y=1.555
+ $X2=11.245 $Y2=1.47
r95 21 33 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=11.245 $Y=1.555
+ $X2=11.245 $Y2=2.52
r96 17 23 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.415 $Y=0.55
+ $X2=11.5 $Y2=0.715
r97 17 19 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=11.415 $Y=0.55
+ $X2=11.24 $Y2=0.55
r98 16 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.345 $Y=1.47
+ $X2=10.18 $Y2=1.47
r99 15 35 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=11.16 $Y=1.47
+ $X2=11.245 $Y2=1.47
r100 15 16 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=11.16 $Y=1.47
+ $X2=10.345 $Y2=1.47
r101 13 40 464.508 $w=1.8e-07 $l=1.195e-06 $layer=POLY_cond $X=10.255 $Y=2.75
+ $X2=10.255 $Y2=1.555
r102 9 39 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=10.09 $Y=0.58
+ $X2=10.09 $Y2=1.225
r103 2 32 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=11.03
+ $Y=2.54 $X2=11.165 $Y2=2.75
r104 1 19 182 $w=1.7e-07 $l=2.52785e-07 $layer=licon1_NDIFF $count=1 $X=11.065
+ $Y=0.37 $X2=11.24 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_4%A_1745_74# 1 2 7 9 12 14 16 18 20 21 23 25
+ 26 28 30 31 32 33 34 38 43 45 46 48 49 51 52 53 63
c158 28 0 1.83478e-19 $X=12.49 $Y=1.765
c159 25 0 1.05829e-19 $X=12.055 $Y=1.615
c160 21 0 1.86508e-19 $X=12.055 $Y=1.185
r161 62 63 35.0294 $w=4.35e-07 $l=7.5e-08 $layer=POLY_cond $X=11.46 $Y=1.117
+ $X2=11.535 $Y2=1.117
r162 57 62 48.5836 $w=4.35e-07 $l=3.8e-07 $layer=POLY_cond $X=11.08 $Y=1.117
+ $X2=11.46 $Y2=1.117
r163 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.08
+ $Y=1.065 $X2=11.08 $Y2=1.065
r164 53 56 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=11.08 $Y=0.97
+ $X2=11.08 $Y2=1.065
r165 50 51 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=10.21 $Y=1.895
+ $X2=10.21 $Y2=2.55
r166 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.125 $Y=1.81
+ $X2=10.21 $Y2=1.895
r167 48 49 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=10.125 $Y=1.81
+ $X2=9.755 $Y2=1.81
r168 47 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.755 $Y=0.97
+ $X2=9.67 $Y2=0.97
r169 46 53 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.915 $Y=0.97
+ $X2=11.08 $Y2=0.97
r170 46 47 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=10.915 $Y=0.97
+ $X2=9.755 $Y2=0.97
r171 45 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.67 $Y=1.725
+ $X2=9.755 $Y2=1.81
r172 44 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.67 $Y=1.055
+ $X2=9.67 $Y2=0.97
r173 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.67 $Y=1.055
+ $X2=9.67 $Y2=1.725
r174 43 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.67 $Y=0.885
+ $X2=9.67 $Y2=0.97
r175 42 43 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=9.67 $Y=0.735
+ $X2=9.67 $Y2=0.885
r176 38 51 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.125 $Y=2.715
+ $X2=10.21 $Y2=2.55
r177 38 40 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=10.125 $Y=2.715
+ $X2=9.52 $Y2=2.715
r178 34 42 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.585 $Y=0.57
+ $X2=9.67 $Y2=0.735
r179 34 36 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=9.585 $Y=0.57
+ $X2=9.405 $Y2=0.57
r180 28 30 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=12.49 $Y=1.765
+ $X2=12.49 $Y2=2.26
r181 27 32 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=12.13 $Y=1.69
+ $X2=12.04 $Y2=1.69
r182 26 28 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=12.4 $Y=1.69
+ $X2=12.49 $Y2=1.765
r183 26 27 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=12.4 $Y=1.69
+ $X2=12.13 $Y2=1.69
r184 25 32 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=12.055
+ $Y=1.615 $X2=12.04 $Y2=1.69
r185 24 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.055 $Y=1.335
+ $X2=12.055 $Y2=1.26
r186 24 25 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=12.055 $Y=1.335
+ $X2=12.055 $Y2=1.615
r187 21 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.055 $Y=1.185
+ $X2=12.055 $Y2=1.26
r188 21 23 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=12.055 $Y=1.185
+ $X2=12.055 $Y2=0.74
r189 18 32 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=12.04 $Y=1.765
+ $X2=12.04 $Y2=1.69
r190 18 20 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=12.04 $Y=1.765
+ $X2=12.04 $Y2=2.26
r191 16 33 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.98 $Y=1.26
+ $X2=12.055 $Y2=1.26
r192 16 63 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=11.98 $Y=1.26
+ $X2=11.535 $Y2=1.26
r193 12 31 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.475 $Y=1.665
+ $X2=11.475 $Y2=1.575
r194 12 14 421.75 $w=1.8e-07 $l=1.085e-06 $layer=POLY_cond $X=11.475 $Y=1.665
+ $X2=11.475 $Y2=2.75
r195 10 62 27.9254 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=11.46 $Y=1.335
+ $X2=11.46 $Y2=1.117
r196 10 31 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=11.46 $Y=1.335
+ $X2=11.46 $Y2=1.575
r197 7 57 11.5066 $w=4.35e-07 $l=9e-08 $layer=POLY_cond $X=10.99 $Y=1.117
+ $X2=11.08 $Y2=1.117
r198 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.99 $Y=0.9
+ $X2=10.99 $Y2=0.58
r199 2 40 600 $w=1.7e-07 $l=1.12219e-06 $layer=licon1_PDIFF $count=1 $X=9.215
+ $Y=1.735 $X2=9.52 $Y2=2.715
r200 1 36 182 $w=1.7e-07 $l=7.73563e-07 $layer=licon1_NDIFF $count=1 $X=8.725
+ $Y=0.37 $X2=9.405 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_4%A_2339_74# 1 2 7 9 10 11 12 14 17 21 25 27
+ 29 32 34 36 39 43 45 50 63
c120 63 0 2.72846e-20 $X=14.375 $Y=1.412
r121 63 64 1.28877 $w=3.74e-07 $l=1e-08 $layer=POLY_cond $X=14.375 $Y=1.412
+ $X2=14.385 $Y2=1.412
r122 62 63 54.1283 $w=3.74e-07 $l=4.2e-07 $layer=POLY_cond $X=13.955 $Y=1.412
+ $X2=14.375 $Y2=1.412
r123 61 62 3.86631 $w=3.74e-07 $l=3e-08 $layer=POLY_cond $X=13.925 $Y=1.412
+ $X2=13.955 $Y2=1.412
r124 58 59 57.9947 $w=3.74e-07 $l=4.5e-07 $layer=POLY_cond $X=13.025 $Y=1.412
+ $X2=13.475 $Y2=1.412
r125 53 55 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=11.84 $Y=1.435
+ $X2=12.265 $Y2=1.435
r126 51 61 30.9305 $w=3.74e-07 $l=2.4e-07 $layer=POLY_cond $X=13.685 $Y=1.412
+ $X2=13.925 $Y2=1.412
r127 51 59 27.0642 $w=3.74e-07 $l=2.1e-07 $layer=POLY_cond $X=13.685 $Y=1.412
+ $X2=13.475 $Y2=1.412
r128 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.685
+ $Y=1.435 $X2=13.685 $Y2=1.435
r129 48 58 2.57754 $w=3.74e-07 $l=2e-08 $layer=POLY_cond $X=13.005 $Y=1.412
+ $X2=13.025 $Y2=1.412
r130 48 56 11.5989 $w=3.74e-07 $l=9e-08 $layer=POLY_cond $X=13.005 $Y=1.412
+ $X2=12.915 $Y2=1.412
r131 47 50 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=13.005 $Y=1.435
+ $X2=13.685 $Y2=1.435
r132 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.005
+ $Y=1.435 $X2=13.005 $Y2=1.435
r133 45 55 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.43 $Y=1.435
+ $X2=12.265 $Y2=1.435
r134 45 47 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=12.43 $Y=1.435
+ $X2=13.005 $Y2=1.435
r135 41 55 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=12.265 $Y=1.6
+ $X2=12.265 $Y2=1.435
r136 41 43 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=12.265 $Y=1.6
+ $X2=12.265 $Y2=1.985
r137 37 53 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.84 $Y=1.27
+ $X2=11.84 $Y2=1.435
r138 37 39 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=11.84 $Y=1.27
+ $X2=11.84 $Y2=0.515
r139 34 64 24.2268 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=14.385 $Y=1.225
+ $X2=14.385 $Y2=1.412
r140 34 36 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=14.385 $Y=1.225
+ $X2=14.385 $Y2=0.74
r141 30 63 19.8678 $w=1.8e-07 $l=1.88e-07 $layer=POLY_cond $X=14.375 $Y=1.6
+ $X2=14.375 $Y2=1.412
r142 30 32 310.968 $w=1.8e-07 $l=8e-07 $layer=POLY_cond $X=14.375 $Y=1.6
+ $X2=14.375 $Y2=2.4
r143 27 62 24.2268 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=13.955 $Y=1.225
+ $X2=13.955 $Y2=1.412
r144 27 29 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=13.955 $Y=1.225
+ $X2=13.955 $Y2=0.74
r145 23 61 19.8678 $w=1.8e-07 $l=1.88e-07 $layer=POLY_cond $X=13.925 $Y=1.6
+ $X2=13.925 $Y2=1.412
r146 23 25 310.968 $w=1.8e-07 $l=8e-07 $layer=POLY_cond $X=13.925 $Y=1.6
+ $X2=13.925 $Y2=2.4
r147 19 59 19.8678 $w=1.8e-07 $l=1.88e-07 $layer=POLY_cond $X=13.475 $Y=1.6
+ $X2=13.475 $Y2=1.412
r148 19 21 310.968 $w=1.8e-07 $l=8e-07 $layer=POLY_cond $X=13.475 $Y=1.6
+ $X2=13.475 $Y2=2.4
r149 15 58 19.8678 $w=1.8e-07 $l=1.88e-07 $layer=POLY_cond $X=13.025 $Y=1.6
+ $X2=13.025 $Y2=1.412
r150 15 17 310.968 $w=1.8e-07 $l=8e-07 $layer=POLY_cond $X=13.025 $Y=1.6
+ $X2=13.025 $Y2=2.4
r151 12 56 24.2268 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=12.915 $Y=1.225
+ $X2=12.915 $Y2=1.412
r152 12 14 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=12.915 $Y=1.225
+ $X2=12.915 $Y2=0.74
r153 10 56 27.5199 $w=3.74e-07 $l=1.4472e-07 $layer=POLY_cond $X=12.84 $Y=1.3
+ $X2=12.915 $Y2=1.412
r154 10 11 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=12.84 $Y=1.3
+ $X2=12.56 $Y2=1.3
r155 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.485 $Y=1.225
+ $X2=12.56 $Y2=1.3
r156 7 9 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=12.485 $Y=1.225
+ $X2=12.485 $Y2=0.74
r157 2 43 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=12.13
+ $Y=1.84 $X2=12.265 $Y2=1.985
r158 1 39 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=11.695
+ $Y=0.37 $X2=11.84 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_4%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 43 47 53
+ 57 61 65 69 71 73 76 77 79 80 81 83 88 100 114 118 123 129 136 139 142 145 148
+ 151 155
c191 3 0 1.21102e-19 $X=4.735 $Y=1.935
r192 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r193 151 152 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r194 149 152 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.68 $Y2=3.33
r195 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r196 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r197 142 143 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r198 136 137 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r199 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r200 129 132 11.1084 $w=9.48e-07 $l=8.65e-07 $layer=LI1_cond $X=1.09 $Y=2.465
+ $X2=1.09 $Y2=3.33
r201 127 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=14.64 $Y2=3.33
r202 127 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.68 $Y2=3.33
r203 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r204 124 151 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.865 $Y=3.33
+ $X2=13.74 $Y2=3.33
r205 124 126 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.865 $Y=3.33
+ $X2=14.16 $Y2=3.33
r206 123 154 4.40486 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=14.47 $Y=3.33
+ $X2=14.675 $Y2=3.33
r207 123 126 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=14.47 $Y=3.33
+ $X2=14.16 $Y2=3.33
r208 122 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r209 122 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r210 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r211 119 145 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.9 $Y=3.33
+ $X2=11.775 $Y2=3.33
r212 119 121 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=11.9 $Y=3.33
+ $X2=12.24 $Y2=3.33
r213 118 148 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.635 $Y=3.33
+ $X2=12.76 $Y2=3.33
r214 118 121 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=12.635 $Y=3.33
+ $X2=12.24 $Y2=3.33
r215 117 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r216 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r217 114 145 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.65 $Y=3.33
+ $X2=11.775 $Y2=3.33
r218 114 116 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=11.65 $Y=3.33
+ $X2=11.28 $Y2=3.33
r219 113 117 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r220 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r221 110 113 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r222 110 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r223 109 112 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r224 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r225 107 142 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.535 $Y=3.33
+ $X2=8.45 $Y2=3.33
r226 107 109 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.535 $Y=3.33
+ $X2=8.88 $Y2=3.33
r227 105 106 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r228 103 106 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r229 102 105 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.96 $Y2=3.33
r230 102 103 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r231 100 139 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=7.17 $Y=3.33
+ $X2=7.345 $Y2=3.33
r232 100 105 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.17 $Y=3.33
+ $X2=6.96 $Y2=3.33
r233 99 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r234 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r235 96 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r236 96 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r237 95 98 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r238 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r239 93 136 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=3.45 $Y=3.33
+ $X2=3.272 $Y2=3.33
r240 93 95 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.45 $Y=3.33 $X2=3.6
+ $Y2=3.33
r241 92 137 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r242 92 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r243 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r244 89 132 11.3727 $w=1.7e-07 $l=4.75e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.09 $Y2=3.33
r245 89 91 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.565 $Y=3.33
+ $X2=1.68 $Y2=3.33
r246 88 136 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=3.272 $Y2=3.33
r247 88 91 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=1.68 $Y2=3.33
r248 86 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r249 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r250 83 132 11.3727 $w=1.7e-07 $l=4.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=1.09 $Y2=3.33
r251 83 85 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r252 81 143 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r253 81 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r254 81 139 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r255 79 112 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=10.465 $Y=3.33
+ $X2=10.32 $Y2=3.33
r256 79 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.465 $Y=3.33
+ $X2=10.63 $Y2=3.33
r257 78 116 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=10.795 $Y=3.33
+ $X2=11.28 $Y2=3.33
r258 78 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.795 $Y=3.33
+ $X2=10.63 $Y2=3.33
r259 76 98 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.56 $Y2=3.33
r260 76 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.87 $Y2=3.33
r261 75 102 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=5.04 $Y2=3.33
r262 75 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=4.87 $Y2=3.33
r263 71 154 3.07266 $w=2.95e-07 $l=1.1025e-07 $layer=LI1_cond $X=14.617 $Y=3.245
+ $X2=14.675 $Y2=3.33
r264 71 73 37.8939 $w=2.93e-07 $l=9.7e-07 $layer=LI1_cond $X=14.617 $Y=3.245
+ $X2=14.617 $Y2=2.275
r265 67 151 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.74 $Y=3.245
+ $X2=13.74 $Y2=3.33
r266 67 69 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=13.74 $Y=3.245
+ $X2=13.74 $Y2=2.275
r267 66 148 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.885 $Y=3.33
+ $X2=12.76 $Y2=3.33
r268 65 151 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.615 $Y=3.33
+ $X2=13.74 $Y2=3.33
r269 65 66 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=13.615 $Y=3.33
+ $X2=12.885 $Y2=3.33
r270 61 64 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=12.76 $Y=1.985
+ $X2=12.76 $Y2=2.815
r271 59 148 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.76 $Y=3.245
+ $X2=12.76 $Y2=3.33
r272 59 64 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=12.76 $Y=3.245
+ $X2=12.76 $Y2=2.815
r273 55 145 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.775 $Y=3.245
+ $X2=11.775 $Y2=3.33
r274 55 57 58.0831 $w=2.48e-07 $l=1.26e-06 $layer=LI1_cond $X=11.775 $Y=3.245
+ $X2=11.775 $Y2=1.985
r275 51 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.63 $Y=3.245
+ $X2=10.63 $Y2=3.33
r276 51 53 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.63 $Y=3.245
+ $X2=10.63 $Y2=2.75
r277 47 50 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.45 $Y=1.91
+ $X2=8.45 $Y2=2.59
r278 45 142 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.45 $Y=3.245
+ $X2=8.45 $Y2=3.33
r279 45 50 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=8.45 $Y=3.245
+ $X2=8.45 $Y2=2.59
r280 44 139 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=7.52 $Y=3.33
+ $X2=7.345 $Y2=3.33
r281 43 142 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.365 $Y=3.33
+ $X2=8.45 $Y2=3.33
r282 43 44 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=8.365 $Y=3.33
+ $X2=7.52 $Y2=3.33
r283 39 139 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.345 $Y=3.245
+ $X2=7.345 $Y2=3.33
r284 39 41 13.8293 $w=3.48e-07 $l=4.2e-07 $layer=LI1_cond $X=7.345 $Y=3.245
+ $X2=7.345 $Y2=2.825
r285 35 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=3.33
r286 35 37 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=4.87 $Y=3.245
+ $X2=4.87 $Y2=2.88
r287 31 136 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=3.272 $Y=3.245
+ $X2=3.272 $Y2=3.33
r288 31 33 14.7707 $w=3.53e-07 $l=4.55e-07 $layer=LI1_cond $X=3.272 $Y=3.245
+ $X2=3.272 $Y2=2.79
r289 10 73 300 $w=1.7e-07 $l=4.97946e-07 $layer=licon1_PDIFF $count=2 $X=14.465
+ $Y=1.84 $X2=14.6 $Y2=2.275
r290 9 69 300 $w=1.7e-07 $l=4.97946e-07 $layer=licon1_PDIFF $count=2 $X=13.565
+ $Y=1.84 $X2=13.7 $Y2=2.275
r291 8 64 600 $w=1.7e-07 $l=1.07941e-06 $layer=licon1_PDIFF $count=1 $X=12.58
+ $Y=1.84 $X2=12.8 $Y2=2.815
r292 8 61 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=12.58
+ $Y=1.84 $X2=12.8 $Y2=1.985
r293 7 57 300 $w=1.7e-07 $l=6.68412e-07 $layer=licon1_PDIFF $count=2 $X=11.565
+ $Y=2.54 $X2=11.815 $Y2=1.985
r294 6 53 600 $w=1.7e-07 $l=3.756e-07 $layer=licon1_PDIFF $count=1 $X=10.345
+ $Y=2.54 $X2=10.63 $Y2=2.75
r295 5 50 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=8.305
+ $Y=1.735 $X2=8.45 $Y2=2.59
r296 5 47 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=8.305
+ $Y=1.735 $X2=8.45 $Y2=1.91
r297 4 41 600 $w=1.7e-07 $l=6.14329e-07 $layer=licon1_PDIFF $count=1 $X=7.115
+ $Y=2.315 $X2=7.345 $Y2=2.825
r298 3 37 600 $w=1.7e-07 $l=1.01025e-06 $layer=licon1_PDIFF $count=1 $X=4.735
+ $Y=1.935 $X2=4.87 $Y2=2.88
r299 2 33 600 $w=1.7e-07 $l=5.35444e-07 $layer=licon1_PDIFF $count=1 $X=3.145
+ $Y=2.32 $X2=3.285 $Y2=2.79
r300 1 129 150 $w=1.7e-07 $l=8.745e-07 $layer=licon1_PDIFF $count=4 $X=0.595
+ $Y=2.32 $X2=1.4 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_4%A_415_81# 1 2 3 4 5 18 20 23 26 30 33 34 35
+ 36 37 39 41 43 48
c144 48 0 1.34001e-19 $X=3.732 $Y=2.54
c145 36 0 1.2914e-19 $X=6.375 $Y=2.17
c146 34 0 1.59809e-19 $X=6.375 $Y=1.33
c147 30 0 8.28381e-20 $X=5.875 $Y=0.9
c148 26 0 1.12508e-19 $X=5.825 $Y=2.54
r149 47 48 1.8083 $w=5.06e-07 $l=7.5e-08 $layer=LI1_cond $X=3.732 $Y=2.465
+ $X2=3.732 $Y2=2.54
r150 45 47 0.843874 $w=5.06e-07 $l=3.5e-08 $layer=LI1_cond $X=3.732 $Y=2.43
+ $X2=3.732 $Y2=2.465
r151 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.46 $Y=1.415
+ $X2=6.46 $Y2=2.085
r152 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.375 $Y=2.17
+ $X2=6.46 $Y2=2.085
r153 36 37 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.375 $Y=2.17
+ $X2=6.075 $Y2=2.17
r154 34 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.375 $Y=1.33
+ $X2=6.46 $Y2=1.415
r155 34 35 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.375 $Y=1.33
+ $X2=5.96 $Y2=1.33
r156 33 50 3.11073 $w=2.5e-07 $l=1.35e-07 $layer=LI1_cond $X=5.95 $Y=2.455
+ $X2=5.95 $Y2=2.59
r157 32 37 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.95 $Y=2.255
+ $X2=6.075 $Y2=2.17
r158 32 33 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=5.95 $Y=2.255
+ $X2=5.95 $Y2=2.455
r159 28 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.875 $Y=1.245
+ $X2=5.96 $Y2=1.33
r160 28 30 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.875 $Y=1.245
+ $X2=5.875 $Y2=0.9
r161 27 48 7.23163 $w=1.7e-07 $l=2.88e-07 $layer=LI1_cond $X=4.02 $Y=2.54
+ $X2=3.732 $Y2=2.54
r162 26 50 4.03243 $w=1.7e-07 $l=1.47902e-07 $layer=LI1_cond $X=5.825 $Y=2.54
+ $X2=5.95 $Y2=2.59
r163 26 27 117.759 $w=1.68e-07 $l=1.805e-06 $layer=LI1_cond $X=5.825 $Y=2.54
+ $X2=4.02 $Y2=2.54
r164 23 45 7.81629 $w=5.06e-07 $l=2.40778e-07 $layer=LI1_cond $X=3.53 $Y=2.345
+ $X2=3.732 $Y2=2.43
r165 22 23 81.877 $w=1.68e-07 $l=1.255e-06 $layer=LI1_cond $X=3.53 $Y=1.09
+ $X2=3.53 $Y2=2.345
r166 21 43 13.5324 $w=2.93e-07 $l=4.16203e-07 $layer=LI1_cond $X=2.735 $Y=1.005
+ $X2=2.527 $Y2=0.68
r167 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.445 $Y=1.005
+ $X2=3.53 $Y2=1.09
r168 20 21 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.445 $Y=1.005
+ $X2=2.735 $Y2=1.005
r169 19 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.435 $Y=2.43
+ $X2=2.27 $Y2=2.43
r170 18 45 7.23163 $w=1.7e-07 $l=2.87e-07 $layer=LI1_cond $X=3.445 $Y=2.43
+ $X2=3.732 $Y2=2.43
r171 18 19 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.445 $Y=2.43
+ $X2=2.435 $Y2=2.43
r172 5 50 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=5.765
+ $Y=2.315 $X2=5.91 $Y2=2.525
r173 4 47 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.715
+ $Y=2.32 $X2=3.855 $Y2=2.465
r174 3 41 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.135
+ $Y=2.32 $X2=2.27 $Y2=2.465
r175 2 30 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=5.75
+ $Y=0.69 $X2=5.875 $Y2=0.9
r176 1 43 182 $w=1.7e-07 $l=5.29953e-07 $layer=licon1_NDIFF $count=1 $X=2.075
+ $Y=0.405 $X2=2.485 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_4%Q 1 2 3 4 15 17 18 21 25 26 29 35 38 40
c68 26 0 1.83478e-19 $X=13.415 $Y=1.855
c69 15 0 1.86508e-19 $X=12.7 $Y=0.515
r70 42 43 0.0389776 $w=6.26e-07 $l=2e-09 $layer=LI1_cond $X=14.17 $Y=1.62
+ $X2=14.172 $Y2=1.62
r71 40 43 9.12077 $w=6.26e-07 $l=4.68e-07 $layer=LI1_cond $X=14.64 $Y=1.62
+ $X2=14.172 $Y2=1.62
r72 38 42 8.59112 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=14.17 $Y=1.3
+ $X2=14.17 $Y2=1.62
r73 37 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.17 $Y=1.1
+ $X2=14.17 $Y2=1.015
r74 37 38 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=14.17 $Y=1.1 $X2=14.17
+ $Y2=1.3
r75 33 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.17 $Y=0.93
+ $X2=14.17 $Y2=1.015
r76 33 35 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=14.17 $Y=0.93
+ $X2=14.17 $Y2=0.515
r77 29 31 44.4897 $w=2.13e-07 $l=8.3e-07 $layer=LI1_cond $X=14.172 $Y=1.985
+ $X2=14.172 $Y2=2.815
r78 27 43 7.10307 $w=2.15e-07 $l=3.2e-07 $layer=LI1_cond $X=14.172 $Y=1.94
+ $X2=14.172 $Y2=1.62
r79 27 29 2.41209 $w=2.13e-07 $l=4.5e-08 $layer=LI1_cond $X=14.172 $Y=1.94
+ $X2=14.172 $Y2=1.985
r80 25 42 9.36281 $w=6.26e-07 $l=2.82666e-07 $layer=LI1_cond $X=14.065 $Y=1.855
+ $X2=14.17 $Y2=1.62
r81 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=14.065 $Y=1.855
+ $X2=13.415 $Y2=1.855
r82 21 23 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=13.25 $Y=1.985
+ $X2=13.25 $Y2=2.815
r83 19 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=13.25 $Y=1.94
+ $X2=13.415 $Y2=1.855
r84 19 21 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=13.25 $Y=1.94
+ $X2=13.25 $Y2=1.985
r85 17 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.085 $Y=1.015
+ $X2=14.17 $Y2=1.015
r86 17 18 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=14.085 $Y=1.015
+ $X2=12.865 $Y2=1.015
r87 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.7 $Y=0.93
+ $X2=12.865 $Y2=1.015
r88 13 15 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=12.7 $Y=0.93
+ $X2=12.7 $Y2=0.515
r89 4 31 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=14.015
+ $Y=1.84 $X2=14.15 $Y2=2.815
r90 4 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=14.015
+ $Y=1.84 $X2=14.15 $Y2=1.985
r91 3 23 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=13.115
+ $Y=1.84 $X2=13.25 $Y2=2.815
r92 3 21 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=13.115
+ $Y=1.84 $X2=13.25 $Y2=1.985
r93 2 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.03
+ $Y=0.37 $X2=14.17 $Y2=0.515
r94 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.56
+ $Y=0.37 $X2=12.7 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_4%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 45 47
+ 50 51 53 54 55 57 72 76 84 97 103 107 113 116 121 127 130
c145 130 0 3.56444e-20 $X=14.64 $Y=0
c146 47 0 2.72846e-20 $X=14.6 $Y=0.515
c147 35 0 1.24672e-19 $X=4.87 $Y=0.665
r148 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r149 126 127 11.7074 $w=8.43e-07 $l=1.65e-07 $layer=LI1_cond $X=13.74 $Y=0.337
+ $X2=13.905 $Y2=0.337
r150 123 126 0.849286 $w=8.43e-07 $l=6e-08 $layer=LI1_cond $X=13.68 $Y=0.337
+ $X2=13.74 $Y2=0.337
r151 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r152 120 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=13.68 $Y2=0
r153 119 123 6.79429 $w=8.43e-07 $l=4.8e-07 $layer=LI1_cond $X=13.2 $Y=0.337
+ $X2=13.68 $Y2=0.337
r154 119 121 11.7074 $w=8.43e-07 $l=1.65e-07 $layer=LI1_cond $X=13.2 $Y=0.337
+ $X2=13.035 $Y2=0.337
r155 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r156 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r157 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r158 107 110 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=7.595 $Y=0
+ $X2=7.595 $Y2=0.325
r159 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r160 101 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=14.64 $Y2=0
r161 101 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=13.68 $Y2=0
r162 100 127 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=14.16 $Y=0
+ $X2=13.905 $Y2=0
r163 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r164 97 129 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=14.435 $Y=0
+ $X2=14.657 $Y2=0
r165 97 100 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=14.435 $Y=0
+ $X2=14.16 $Y2=0
r166 96 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r167 96 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r168 95 121 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.72 $Y=0
+ $X2=13.035 $Y2=0
r169 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r170 93 116 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=12.365 $Y=0
+ $X2=12.235 $Y2=0
r171 93 95 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=12.365 $Y=0
+ $X2=12.72 $Y2=0
r172 91 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r173 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r174 88 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.76 $Y2=0
r175 88 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r176 87 90 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=10.8 $Y=0 $X2=11.76
+ $Y2=0
r177 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r178 85 113 10.4332 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=10.58 $Y=0
+ $X2=10.36 $Y2=0
r179 85 87 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=10.58 $Y=0 $X2=10.8
+ $Y2=0
r180 84 116 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=12.105 $Y=0
+ $X2=12.235 $Y2=0
r181 84 90 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=12.105 $Y=0
+ $X2=11.76 $Y2=0
r182 83 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r183 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r184 80 83 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=9.84 $Y2=0
r185 79 82 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=7.92 $Y=0 $X2=9.84
+ $Y2=0
r186 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r187 77 107 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.76 $Y=0
+ $X2=7.595 $Y2=0
r188 77 79 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.76 $Y=0 $X2=7.92
+ $Y2=0
r189 76 113 10.4332 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=10.14 $Y=0
+ $X2=10.36 $Y2=0
r190 76 82 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=10.14 $Y=0 $X2=9.84
+ $Y2=0
r191 74 75 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r192 72 107 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.43 $Y=0
+ $X2=7.595 $Y2=0
r193 72 74 155.925 $w=1.68e-07 $l=2.39e-06 $layer=LI1_cond $X=7.43 $Y=0 $X2=5.04
+ $Y2=0
r194 71 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r195 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r196 68 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r197 67 68 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r198 65 68 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r199 65 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r200 64 67 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r201 64 65 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r202 62 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0
+ $X2=0.71 $Y2=0
r203 62 64 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r204 60 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r205 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r206 57 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.71 $Y2=0
r207 57 59 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r208 55 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r209 55 75 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=7.44 $Y=0 $X2=5.04
+ $Y2=0
r210 55 107 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r211 53 70 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=0
+ $X2=4.56 $Y2=0
r212 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=0 $X2=4.87
+ $Y2=0
r213 52 74 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=0 $X2=5.04
+ $Y2=0
r214 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=0 $X2=4.87
+ $Y2=0
r215 50 67 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=3.64 $Y=0 $X2=3.6
+ $Y2=0
r216 50 51 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.64 $Y=0 $X2=3.79
+ $Y2=0
r217 49 70 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.94 $Y=0 $X2=4.56
+ $Y2=0
r218 49 51 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.94 $Y=0 $X2=3.79
+ $Y2=0
r219 45 129 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=14.6 $Y=0.085
+ $X2=14.657 $Y2=0
r220 45 47 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=14.6 $Y=0.085
+ $X2=14.6 $Y2=0.515
r221 41 116 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=12.235 $Y=0.085
+ $X2=12.235 $Y2=0
r222 41 43 19.0596 $w=2.58e-07 $l=4.3e-07 $layer=LI1_cond $X=12.235 $Y=0.085
+ $X2=12.235 $Y2=0.515
r223 37 113 1.73497 $w=4.4e-07 $l=8.5e-08 $layer=LI1_cond $X=10.36 $Y=0.085
+ $X2=10.36 $Y2=0
r224 37 39 11.2625 $w=4.38e-07 $l=4.3e-07 $layer=LI1_cond $X=10.36 $Y=0.085
+ $X2=10.36 $Y2=0.515
r225 33 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=0.085
+ $X2=4.87 $Y2=0
r226 33 35 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=4.87 $Y=0.085
+ $X2=4.87 $Y2=0.665
r227 29 51 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.79 $Y=0.085
+ $X2=3.79 $Y2=0
r228 29 31 19.2074 $w=2.98e-07 $l=5e-07 $layer=LI1_cond $X=3.79 $Y=0.085
+ $X2=3.79 $Y2=0.585
r229 25 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r230 25 27 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.555
r231 8 47 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.46
+ $Y=0.37 $X2=14.6 $Y2=0.515
r232 7 126 91 $w=1.7e-07 $l=8.55132e-07 $layer=licon1_NDIFF $count=2 $X=12.99
+ $Y=0.37 $X2=13.74 $Y2=0.595
r233 6 43 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.13
+ $Y=0.37 $X2=12.27 $Y2=0.515
r234 5 39 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=10.165
+ $Y=0.37 $X2=10.36 $Y2=0.515
r235 4 110 182 $w=1.7e-07 $l=4.62088e-07 $layer=licon1_NDIFF $count=1 $X=7.375
+ $Y=0.69 $X2=7.595 $Y2=0.325
r236 3 35 182 $w=1.7e-07 $l=2.32379e-07 $layer=licon1_NDIFF $count=1 $X=4.67
+ $Y=0.595 $X2=4.87 $Y2=0.665
r237 2 31 182 $w=1.7e-07 $l=2.47386e-07 $layer=licon1_NDIFF $count=1 $X=3.615
+ $Y=0.405 $X2=3.775 $Y2=0.585
r238 1 27 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTP_4%noxref_24 1 2 7 9 14
c30 7 0 2.58874e-19 $X=3.14 $Y=0.34
r31 14 17 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=3.305 $Y=0.34
+ $X2=3.305 $Y2=0.565
r32 9 12 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.27 $Y=0.34 $X2=1.27
+ $Y2=0.55
r33 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.435 $Y=0.34 $X2=1.27
+ $Y2=0.34
r34 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=0.34
+ $X2=3.305 $Y2=0.34
r35 7 8 111.235 $w=1.68e-07 $l=1.705e-06 $layer=LI1_cond $X=3.14 $Y=0.34
+ $X2=1.435 $Y2=0.34
r36 2 17 182 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_NDIFF $count=1 $X=3.135
+ $Y=0.405 $X2=3.305 $Y2=0.565
r37 1 12 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.405 $X2=1.27 $Y2=0.55
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__or3_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.280000 0.435000 1.110000 ;
        RECT 0.105000 1.110000 3.055000 1.280000 ;
        RECT 0.105000 1.280000 0.435000 1.630000 ;
        RECT 2.755000 1.280000 3.055000 1.550000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.450000 2.545000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.270000 1.380000 0.940000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  1.090100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.565000 0.350000 3.735000 0.960000 ;
        RECT 3.565000 0.960000 5.155000 1.130000 ;
        RECT 3.565000 1.800000 5.155000 1.970000 ;
        RECT 3.565000 1.970000 3.735000 2.980000 ;
        RECT 4.385000 1.970000 4.715000 2.980000 ;
        RECT 4.405000 0.350000 4.655000 0.960000 ;
        RECT 4.925000 1.130000 5.155000 1.800000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.115000  1.920000 0.365000 3.245000 ;
      RECT 0.565000  1.950000 0.815000 2.370000 ;
      RECT 0.565000  2.370000 2.830000 2.540000 ;
      RECT 0.565000  2.540000 0.815000 2.960000 ;
      RECT 1.015000  2.710000 2.330000 2.960000 ;
      RECT 1.495000  1.950000 3.395000 2.120000 ;
      RECT 1.495000  2.120000 1.825000 2.200000 ;
      RECT 1.550000  0.350000 1.880000 0.770000 ;
      RECT 1.550000  0.770000 3.395000 0.940000 ;
      RECT 2.050000  0.085000 2.380000 0.600000 ;
      RECT 2.500000  2.290000 2.830000 2.370000 ;
      RECT 2.500000  2.540000 2.830000 2.960000 ;
      RECT 2.550000  0.350000 2.880000 0.770000 ;
      RECT 3.035000  2.290000 3.365000 3.245000 ;
      RECT 3.050000  0.085000 3.380000 0.600000 ;
      RECT 3.225000  0.940000 3.395000 1.300000 ;
      RECT 3.225000  1.300000 4.685000 1.630000 ;
      RECT 3.225000  1.630000 3.395000 1.950000 ;
      RECT 3.915000  0.085000 4.165000 0.790000 ;
      RECT 3.935000  2.140000 4.185000 3.245000 ;
      RECT 4.835000  0.085000 5.165000 0.790000 ;
      RECT 4.915000  2.140000 5.165000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_ms__or3_4
END LIBRARY

* File: sky130_fd_sc_ms__mux4_2.pex.spice
* Created: Fri Aug 28 17:40:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__MUX4_2%S0 3 6 10 14 18 21 24 25 26 28 31 32 34 36 40
+ 41 44 47 48 49 53 55 59 61 70
c171 70 0 9.37441e-20 $X=4.56 $Y=1.22
c172 59 0 1.77444e-19 $X=0.6 $Y=1.385
c173 53 0 4.5023e-20 $X=4.56 $Y=1.385
c174 49 0 2.33726e-19 $X=4.56 $Y=1.195
c175 44 0 1.72582e-19 $X=1.485 $Y=1.195
c176 31 0 1.35612e-19 $X=2.94 $Y=1.615
c177 14 0 2.47412e-19 $X=3.015 $Y=2.46
r178 59 62 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.6 $Y=1.385
+ $X2=0.6 $Y2=1.55
r179 59 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.6 $Y=1.385
+ $X2=0.6 $Y2=1.22
r180 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.385 $X2=0.6 $Y2=1.385
r181 55 60 3.24852 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=0.62 $Y=1.295
+ $X2=0.62 $Y2=1.385
r182 55 77 3.60947 $w=3.38e-07 $l=1e-07 $layer=LI1_cond $X=0.62 $Y=1.295
+ $X2=0.62 $Y2=1.195
r183 55 77 4.76605 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.805 $Y=1.195
+ $X2=0.62 $Y2=1.195
r184 53 70 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.56 $Y=1.385
+ $X2=4.56 $Y2=1.22
r185 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.56
+ $Y=1.385 $X2=4.56 $Y2=1.385
r186 49 52 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.56 $Y=1.195
+ $X2=4.56 $Y2=1.385
r187 47 64 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=1.425
+ $X2=1.68 $Y2=1.26
r188 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.425 $X2=1.68 $Y2=1.425
r189 44 55 33.6483 $w=2.38e-07 $l=6.8e-07 $layer=LI1_cond $X=1.485 $Y=1.195
+ $X2=0.805 $Y2=1.195
r190 44 46 9.35333 $w=3e-07 $l=3.07083e-07 $layer=LI1_cond $X=1.485 $Y=1.195
+ $X2=1.665 $Y2=1.425
r191 41 74 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.64 $Y=1.585
+ $X2=5.64 $Y2=1.75
r192 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.64
+ $Y=1.585 $X2=5.64 $Y2=1.585
r193 38 40 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.61 $Y=1.28
+ $X2=5.61 $Y2=1.585
r194 37 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.725 $Y=1.195
+ $X2=4.56 $Y2=1.195
r195 36 38 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=5.475 $Y=1.195
+ $X2=5.61 $Y2=1.28
r196 36 37 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=5.475 $Y=1.195
+ $X2=4.725 $Y2=1.195
r197 35 48 3.05049 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.105 $Y=1.195
+ $X2=2.97 $Y2=1.195
r198 34 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.395 $Y=1.195
+ $X2=4.56 $Y2=1.195
r199 34 35 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=4.395 $Y=1.195
+ $X2=3.105 $Y2=1.195
r200 32 68 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.94 $Y=1.615
+ $X2=2.94 $Y2=1.78
r201 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.94
+ $Y=1.615 $X2=2.94 $Y2=1.615
r202 29 48 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=1.28
+ $X2=2.97 $Y2=1.195
r203 29 31 14.2988 $w=2.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.97 $Y=1.28
+ $X2=2.97 $Y2=1.615
r204 28 48 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=1.11
+ $X2=2.97 $Y2=1.195
r205 27 28 22.1952 $w=2.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.97 $Y=0.59
+ $X2=2.97 $Y2=1.11
r206 25 27 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.835 $Y=0.505
+ $X2=2.97 $Y2=0.59
r207 25 26 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=2.835 $Y=0.505
+ $X2=1.655 $Y2=0.505
r208 24 44 5.72868 $w=3e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.57 $Y=1.11
+ $X2=1.485 $Y2=1.195
r209 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.57 $Y=0.59
+ $X2=1.655 $Y2=0.505
r210 23 24 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.57 $Y=0.59
+ $X2=1.57 $Y2=1.11
r211 21 74 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=5.685 $Y=2.46
+ $X2=5.685 $Y2=1.75
r212 18 70 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.47 $Y=0.74
+ $X2=4.47 $Y2=1.22
r213 14 68 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=3.015 $Y=2.46
+ $X2=3.015 $Y2=1.78
r214 10 64 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.59 $Y=0.74
+ $X2=1.59 $Y2=1.26
r215 6 62 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=0.645 $Y=2.46
+ $X2=0.645 $Y2=1.55
r216 3 61 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.515 $Y=0.79
+ $X2=0.515 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_2%A1 3 5 7 9
c34 9 0 1.14029e-19 $X=1.2 $Y=1.665
r35 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=1.615 $X2=1.14 $Y2=1.615
r36 5 12 33.9921 $w=3.34e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.245 $Y=1.78
+ $X2=1.155 $Y2=1.615
r37 5 7 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=1.245 $Y=1.78
+ $X2=1.245 $Y2=2.46
r38 1 12 38.6287 $w=3.34e-07 $l=1.86145e-07 $layer=POLY_cond $X=1.2 $Y=1.45
+ $X2=1.155 $Y2=1.615
r39 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.2 $Y=1.45 $X2=1.2
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_2%A_31_94# 1 2 9 13 15 17 20 26 29 32 33 34 35
+ 38 44 49 50 54 64
c126 50 0 3.08193e-19 $X=2.295 $Y=1.615
c127 49 0 1.67329e-19 $X=2.22 $Y=1.615
c128 34 0 4.5023e-20 $X=4.895 $Y=2.035
c129 15 0 1.11429e-19 $X=4.995 $Y=1.88
r130 66 67 2.37898 $w=4.88e-07 $l=4.5e-08 $layer=LI1_cond $X=0.34 $Y=2.105
+ $X2=0.34 $Y2=2.15
r131 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.1
+ $Y=1.625 $X2=5.1 $Y2=1.625
r132 48 50 13.2418 $w=2.73e-07 $l=7.5e-08 $layer=POLY_cond $X=2.22 $Y=1.615
+ $X2=2.295 $Y2=1.615
r133 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.22
+ $Y=1.615 $X2=2.22 $Y2=1.615
r134 45 54 13.8971 $w=3.38e-07 $l=4.1e-07 $layer=LI1_cond $X=5.095 $Y=2.035
+ $X2=5.095 $Y2=1.625
r135 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=2.035
+ $X2=5.04 $Y2=2.035
r136 42 49 17.2866 $w=2.78e-07 $l=4.2e-07 $layer=LI1_cond $X=2.185 $Y=2.035
+ $X2=2.185 $Y2=1.615
r137 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=2.035
+ $X2=2.16 $Y2=2.035
r138 38 66 1.70868 $w=4.88e-07 $l=7e-08 $layer=LI1_cond $X=0.34 $Y=2.035
+ $X2=0.34 $Y2=2.105
r139 38 64 8.23575 $w=4.88e-07 $l=1.15e-07 $layer=LI1_cond $X=0.34 $Y=2.035
+ $X2=0.34 $Y2=1.92
r140 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=2.035
+ $X2=0.24 $Y2=2.035
r141 35 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=2.035
+ $X2=2.16 $Y2=2.035
r142 34 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=5.04 $Y2=2.035
r143 34 35 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=2.305 $Y2=2.035
r144 33 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.385 $Y=2.035
+ $X2=0.24 $Y2=2.035
r145 32 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.015 $Y=2.035
+ $X2=2.16 $Y2=2.035
r146 32 33 2.01732 $w=1.4e-07 $l=1.63e-06 $layer=MET1_cond $X=2.015 $Y=2.035
+ $X2=0.385 $Y2=2.035
r147 31 64 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=0.18 $Y=1.01
+ $X2=0.18 $Y2=1.92
r148 29 31 11.4978 $w=3.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.28 $Y=0.75
+ $X2=0.28 $Y2=1.01
r149 26 67 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=0.42 $Y=2.815
+ $X2=0.42 $Y2=2.15
r150 18 53 38.5662 $w=2.97e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.16 $Y=1.46
+ $X2=5.085 $Y2=1.625
r151 18 20 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=5.16 $Y=1.46
+ $X2=5.16 $Y2=0.74
r152 15 53 48.8089 $w=2.97e-07 $l=2.96606e-07 $layer=POLY_cond $X=4.995 $Y=1.88
+ $X2=5.085 $Y2=1.625
r153 15 17 155.311 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=4.995 $Y=1.88
+ $X2=4.995 $Y2=2.46
r154 11 50 29.1319 $w=2.73e-07 $l=2.33345e-07 $layer=POLY_cond $X=2.46 $Y=1.45
+ $X2=2.295 $Y2=1.615
r155 11 13 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.46 $Y=1.45
+ $X2=2.46 $Y2=0.74
r156 7 50 12.5437 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=1.78
+ $X2=2.295 $Y2=1.615
r157 7 9 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=2.295 $Y=1.78
+ $X2=2.295 $Y2=2.46
r158 2 66 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.275
+ $Y=1.96 $X2=0.42 $Y2=2.105
r159 2 26 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.275
+ $Y=1.96 $X2=0.42 $Y2=2.815
r160 1 29 182 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_NDIFF $count=1 $X=0.155
+ $Y=0.47 $X2=0.3 $Y2=0.75
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_2%A0 3 5 9 12 15 17
c42 5 0 1.72518e-19 $X=3.48 $Y=1.405
r43 15 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.48 $Y=1.615
+ $X2=3.48 $Y2=1.78
r44 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.48
+ $Y=1.615 $X2=3.48 $Y2=1.615
r45 12 16 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=3.6 $Y=1.615 $X2=3.48
+ $Y2=1.615
r46 9 17 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=3.435 $Y=2.46
+ $X2=3.435 $Y2=1.78
r47 5 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.48 $Y=1.405
+ $X2=3.48 $Y2=1.24
r48 5 15 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=3.48 $Y=1.405
+ $X2=3.48 $Y2=1.615
r49 3 11 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.39 $Y=0.74 $X2=3.39
+ $Y2=1.24
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_2%A3 3 5 7 8
c34 5 0 1.22296e-19 $X=4.125 $Y=1.88
r35 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.02
+ $Y=1.615 $X2=4.02 $Y2=1.615
r36 5 11 50.643 $w=2.94e-07 $l=3.06716e-07 $layer=POLY_cond $X=4.125 $Y=1.88
+ $X2=4.035 $Y2=1.615
r37 5 7 155.311 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=4.125 $Y=1.88
+ $X2=4.125 $Y2=2.46
r38 1 11 38.5845 $w=2.94e-07 $l=1.86145e-07 $layer=POLY_cond $X=4.08 $Y=1.45
+ $X2=4.035 $Y2=1.615
r39 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.08 $Y=1.45 $X2=4.08
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_2%A2 3 6 8 9 13 15
r43 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.18 $Y=1.385
+ $X2=6.18 $Y2=1.55
r44 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.18 $Y=1.385
+ $X2=6.18 $Y2=1.22
r45 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.18
+ $Y=1.385 $X2=6.18 $Y2=1.385
r46 9 14 7.50428 $w=4.28e-07 $l=2.8e-07 $layer=LI1_cond $X=6.13 $Y=1.665
+ $X2=6.13 $Y2=1.385
r47 8 14 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=6.13 $Y=1.295 $X2=6.13
+ $Y2=1.385
r48 6 16 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=6.105 $Y=2.46
+ $X2=6.105 $Y2=1.55
r49 3 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.09 $Y=0.74 $X2=6.09
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_2%A_1500_94# 1 2 7 9 12 15 20 24 27 28
c53 27 0 1.84046e-19 $X=8.23 $Y=1.615
r54 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.23
+ $Y=1.615 $X2=8.23 $Y2=1.615
r55 22 27 6.31733 $w=2.57e-07 $l=1.68953e-07 $layer=LI1_cond $X=8.325 $Y=1.78
+ $X2=8.317 $Y2=1.615
r56 22 24 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=8.325 $Y=1.78
+ $X2=8.325 $Y2=2.155
r57 18 27 6.31733 $w=2.57e-07 $l=1.65e-07 $layer=LI1_cond $X=8.317 $Y=1.45
+ $X2=8.317 $Y2=1.615
r58 18 20 15.2209 $w=2.63e-07 $l=3.5e-07 $layer=LI1_cond $X=8.317 $Y=1.45
+ $X2=8.317 $Y2=1.1
r59 14 28 96.1737 $w=3.3e-07 $l=5.5e-07 $layer=POLY_cond $X=7.68 $Y=1.615
+ $X2=8.23 $Y2=1.615
r60 14 15 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.68 $Y=1.615 $X2=7.59
+ $Y2=1.615
r61 10 15 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=7.59 $Y=1.78
+ $X2=7.59 $Y2=1.615
r62 10 12 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=7.59 $Y=1.78
+ $X2=7.59 $Y2=2.46
r63 7 15 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=7.575 $Y=1.45
+ $X2=7.59 $Y2=1.615
r64 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.575 $Y=1.45 $X2=7.575
+ $Y2=0.97
r65 2 24 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=8.225
+ $Y=1.94 $X2=8.365 $Y2=2.155
r66 1 20 182 $w=1.7e-07 $l=5.70088e-07 $layer=licon1_NDIFF $count=1 $X=8.205
+ $Y=0.6 $X2=8.355 $Y2=1.1
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_2%S1 4 7 9 10 14 15 17 20 23
c77 23 0 1.84046e-19 $X=7.065 $Y=1.615
c78 7 0 6.80408e-20 $X=7.14 $Y=2.46
r79 23 26 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.065 $Y=1.615
+ $X2=7.065 $Y2=1.78
r80 23 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.065 $Y=1.615
+ $X2=7.065 $Y2=1.45
r81 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.065
+ $Y=1.615 $X2=7.065 $Y2=1.615
r82 20 24 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=7.44 $Y=1.615
+ $X2=7.065 $Y2=1.615
r83 15 19 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=8.725 $Y=1.405
+ $X2=8.725 $Y2=1.315
r84 15 17 402.315 $w=1.8e-07 $l=1.035e-06 $layer=POLY_cond $X=8.725 $Y=1.405
+ $X2=8.725 $Y2=2.44
r85 14 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.71 $Y=0.92
+ $X2=8.71 $Y2=1.315
r86 11 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.71 $Y=0.26
+ $X2=8.71 $Y2=0.92
r87 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.635 $Y=0.185
+ $X2=8.71 $Y2=0.26
r88 9 10 764.021 $w=1.5e-07 $l=1.49e-06 $layer=POLY_cond $X=8.635 $Y=0.185
+ $X2=7.145 $Y2=0.185
r89 7 26 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=7.14 $Y=2.46 $X2=7.14
+ $Y2=1.78
r90 4 25 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=7.07 $Y=0.74 $X2=7.07
+ $Y2=1.45
r91 1 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.07 $Y=0.26
+ $X2=7.145 $Y2=0.185
r92 1 4 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.07 $Y=0.26 $X2=7.07
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_2%A_1429_74# 1 2 9 11 13 14 16 19 21 24 26 28
+ 31 33 34 40 47
c102 28 0 6.80408e-20 $X=8.96 $Y=2.99
r103 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.22
+ $Y=1.515 $X2=9.22 $Y2=1.515
r104 44 47 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=9.045 $Y=1.515
+ $X2=9.22 $Y2=1.515
r105 40 42 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=7.365 $Y=2.805
+ $X2=7.365 $Y2=2.99
r106 34 37 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=7.285 $Y=0.34
+ $X2=7.285 $Y2=0.515
r107 32 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.045 $Y=1.68
+ $X2=9.045 $Y2=1.515
r108 32 33 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=9.045 $Y=1.68
+ $X2=9.045 $Y2=2.905
r109 31 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.045 $Y=1.35
+ $X2=9.045 $Y2=1.515
r110 30 31 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=9.045 $Y=0.425
+ $X2=9.045 $Y2=1.35
r111 29 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.53 $Y=2.99
+ $X2=7.365 $Y2=2.99
r112 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.96 $Y=2.99
+ $X2=9.045 $Y2=2.905
r113 28 29 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=8.96 $Y=2.99
+ $X2=7.53 $Y2=2.99
r114 27 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.45 $Y=0.34
+ $X2=7.285 $Y2=0.34
r115 26 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.96 $Y=0.34
+ $X2=9.045 $Y2=0.425
r116 26 27 98.5134 $w=1.68e-07 $l=1.51e-06 $layer=LI1_cond $X=8.96 $Y=0.34
+ $X2=7.45 $Y2=0.34
r117 23 24 68.1616 $w=2.97e-07 $l=4.2e-07 $layer=POLY_cond $X=9.61 $Y=1.515
+ $X2=10.03 $Y2=1.515
r118 22 23 1.6229 $w=2.97e-07 $l=1e-08 $layer=POLY_cond $X=9.6 $Y=1.515 $X2=9.61
+ $Y2=1.515
r119 21 48 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=9.52 $Y=1.515
+ $X2=9.22 $Y2=1.515
r120 21 22 12.2719 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=9.52 $Y=1.515 $X2=9.6
+ $Y2=1.515
r121 17 24 4.86869 $w=2.97e-07 $l=3e-08 $layer=POLY_cond $X=10.06 $Y=1.515
+ $X2=10.03 $Y2=1.515
r122 17 19 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=10.06 $Y=1.65
+ $X2=10.06 $Y2=2.4
r123 14 24 18.7323 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.03 $Y=1.35
+ $X2=10.03 $Y2=1.515
r124 14 16 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=10.03 $Y=1.35
+ $X2=10.03 $Y2=0.87
r125 11 22 18.7323 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.6 $Y=1.35
+ $X2=9.6 $Y2=1.515
r126 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.6 $Y=1.35 $X2=9.6
+ $Y2=0.87
r127 7 23 14.4873 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.61 $Y=1.68
+ $X2=9.61 $Y2=1.515
r128 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=9.61 $Y=1.68 $X2=9.61
+ $Y2=2.4
r129 2 40 600 $w=1.7e-07 $l=9.1e-07 $layer=licon1_PDIFF $count=1 $X=7.23 $Y=1.96
+ $X2=7.365 $Y2=2.805
r130 1 37 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.145
+ $Y=0.37 $X2=7.285 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_2%VPWR 1 2 3 4 5 18 24 28 30 34 38 40 45 46 48
+ 49 50 62 69 75 78 82
c99 18 0 6.34146e-20 $X=0.92 $Y=2.115
r100 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r101 78 79 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r102 76 79 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=9.36 $Y2=3.33
r103 75 76 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r104 73 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r105 73 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r106 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r107 70 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.47 $Y=3.33
+ $X2=9.385 $Y2=3.33
r108 70 72 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.47 $Y=3.33
+ $X2=9.84 $Y2=3.33
r109 69 81 4.01803 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=10.2 $Y=3.33
+ $X2=10.38 $Y2=3.33
r110 69 72 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=10.2 $Y=3.33
+ $X2=9.84 $Y2=3.33
r111 68 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r112 67 68 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r113 64 67 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=3.33 $X2=6
+ $Y2=3.33
r114 64 65 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r115 62 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.165 $Y=3.33
+ $X2=6.33 $Y2=3.33
r116 62 67 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.165 $Y=3.33
+ $X2=6 $Y2=3.33
r117 61 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r118 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r119 58 61 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.6 $Y2=3.33
r120 57 60 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=3.6
+ $Y2=3.33
r121 57 58 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r122 54 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r123 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r124 50 68 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=3.33 $X2=6
+ $Y2=3.33
r125 50 65 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=4.08 $Y2=3.33
r126 48 60 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.615 $Y=3.33
+ $X2=3.6 $Y2=3.33
r127 48 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=3.33
+ $X2=3.78 $Y2=3.33
r128 47 64 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.945 $Y=3.33
+ $X2=4.08 $Y2=3.33
r129 47 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.945 $Y=3.33
+ $X2=3.78 $Y2=3.33
r130 45 53 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=0.755 $Y=3.33
+ $X2=0.72 $Y2=3.33
r131 45 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.755 $Y=3.33
+ $X2=0.92 $Y2=3.33
r132 44 57 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=1.2 $Y2=3.33
r133 44 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.085 $Y=3.33
+ $X2=0.92 $Y2=3.33
r134 40 43 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=10.325 $Y=1.985
+ $X2=10.325 $Y2=2.815
r135 38 81 3.12513 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=10.325 $Y=3.245
+ $X2=10.38 $Y2=3.33
r136 38 43 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.325 $Y=3.245
+ $X2=10.325 $Y2=2.815
r137 34 37 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=9.385 $Y=2.015
+ $X2=9.385 $Y2=2.795
r138 32 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.385 $Y=3.245
+ $X2=9.385 $Y2=3.33
r139 32 37 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=9.385 $Y=3.245
+ $X2=9.385 $Y2=2.795
r140 31 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.495 $Y=3.33
+ $X2=6.33 $Y2=3.33
r141 30 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.3 $Y=3.33
+ $X2=9.385 $Y2=3.33
r142 30 31 183 $w=1.68e-07 $l=2.805e-06 $layer=LI1_cond $X=9.3 $Y=3.33 $X2=6.495
+ $Y2=3.33
r143 26 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.33 $Y=3.245
+ $X2=6.33 $Y2=3.33
r144 26 28 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=6.33 $Y=3.245
+ $X2=6.33 $Y2=2.805
r145 22 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.78 $Y=3.245
+ $X2=3.78 $Y2=3.33
r146 22 24 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=3.78 $Y=3.245
+ $X2=3.78 $Y2=2.455
r147 18 21 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.92 $Y=2.115
+ $X2=0.92 $Y2=2.815
r148 16 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.92 $Y=3.245
+ $X2=0.92 $Y2=3.33
r149 16 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.92 $Y=3.245
+ $X2=0.92 $Y2=2.815
r150 5 43 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.15
+ $Y=1.84 $X2=10.285 $Y2=2.815
r151 5 40 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.15
+ $Y=1.84 $X2=10.285 $Y2=1.985
r152 4 37 400 $w=1.7e-07 $l=1.1038e-06 $layer=licon1_PDIFF $count=1 $X=8.815
+ $Y=1.94 $X2=9.385 $Y2=2.795
r153 4 34 400 $w=1.7e-07 $l=6.06341e-07 $layer=licon1_PDIFF $count=1 $X=8.815
+ $Y=1.94 $X2=9.385 $Y2=2.015
r154 3 28 600 $w=1.7e-07 $l=9.1e-07 $layer=licon1_PDIFF $count=1 $X=6.195
+ $Y=1.96 $X2=6.33 $Y2=2.805
r155 2 24 300 $w=1.7e-07 $l=6.09303e-07 $layer=licon1_PDIFF $count=2 $X=3.525
+ $Y=1.96 $X2=3.78 $Y2=2.455
r156 1 21 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=0.735
+ $Y=1.96 $X2=0.92 $Y2=2.815
r157 1 18 400 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_PDIFF $count=1 $X=0.735
+ $Y=1.96 $X2=0.92 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_2%A_333_74# 1 2 3 4 13 19 22 23 24 25 26 28 29
+ 31 35 37 38 48
c135 38 0 3.59869e-19 $X=2.97 $Y=1.95
c136 29 0 1.65994e-19 $X=6.73 $Y=1.195
c137 19 0 8.00829e-20 $X=4.115 $Y=2.035
r138 40 42 8.98947 $w=9.48e-07 $l=7e-07 $layer=LI1_cond $X=2.97 $Y=2.115
+ $X2=2.97 $Y2=2.815
r139 37 40 1.02737 $w=9.48e-07 $l=8e-08 $layer=LI1_cond $X=2.97 $Y=2.035
+ $X2=2.97 $Y2=2.115
r140 37 38 11.5385 $w=9.48e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=2.035
+ $X2=2.97 $Y2=1.95
r141 33 48 3.77418 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=6.73 $Y=2.075
+ $X2=6.645 $Y2=2.075
r142 33 35 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=6.73 $Y=2.075
+ $X2=6.9 $Y2=2.075
r143 29 31 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=6.73 $Y=1.195
+ $X2=7.79 $Y2=1.195
r144 28 48 2.68609 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.645 $Y=1.95
+ $X2=6.645 $Y2=2.075
r145 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.645 $Y=1.28
+ $X2=6.73 $Y2=1.195
r146 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.645 $Y=1.28
+ $X2=6.645 $Y2=1.95
r147 26 46 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.52 $Y=2.08
+ $X2=5.52 $Y2=2.405
r148 25 48 3.77418 $w=2.45e-07 $l=8.74643e-08 $layer=LI1_cond $X=6.56 $Y=2.08
+ $X2=6.645 $Y2=2.075
r149 25 26 45.8576 $w=2.38e-07 $l=9.55e-07 $layer=LI1_cond $X=6.56 $Y=2.08
+ $X2=5.605 $Y2=2.08
r150 23 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.435 $Y=2.405
+ $X2=5.52 $Y2=2.405
r151 23 24 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=5.435 $Y=2.405
+ $X2=4.285 $Y2=2.405
r152 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.2 $Y=2.32
+ $X2=4.285 $Y2=2.405
r153 21 22 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.2 $Y=2.12 $X2=4.2
+ $Y2=2.32
r154 20 37 11.3727 $w=1.7e-07 $l=4.75e-07 $layer=LI1_cond $X=3.445 $Y=2.035
+ $X2=2.97 $Y2=2.035
r155 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.115 $Y=2.035
+ $X2=4.2 $Y2=2.12
r156 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.115 $Y=2.035
+ $X2=3.445 $Y2=2.035
r157 17 38 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2.58 $Y=1.09
+ $X2=2.58 $Y2=1.95
r158 13 17 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.495 $Y=0.925
+ $X2=2.58 $Y2=1.09
r159 13 15 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=2.495 $Y=0.925
+ $X2=2.08 $Y2=0.925
r160 4 35 600 $w=1.7e-07 $l=2.19203e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.96 $X2=6.9 $Y2=2.115
r161 3 42 400 $w=1.7e-07 $l=9.82929e-07 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=1.96 $X2=2.66 $Y2=2.815
r162 3 40 400 $w=1.7e-07 $l=3.43875e-07 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=1.96 $X2=2.66 $Y2=2.115
r163 2 31 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=7.65
+ $Y=0.6 $X2=7.79 $Y2=1.195
r164 1 15 182 $w=1.7e-07 $l=7.33723e-07 $layer=licon1_NDIFF $count=1 $X=1.665
+ $Y=0.37 $X2=2.08 $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_2%A_909_74# 1 2 3 4 13 17 19 23 25 29 31 33 36
+ 38 42 47 48 50
c128 17 0 9.37441e-20 $X=6.69 $Y=0.855
c129 2 0 1.65994e-19 $X=6.715 $Y=0.37
r130 50 52 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=7.93 $Y=0.68
+ $X2=7.93 $Y2=0.855
r131 48 49 9.75 $w=2.44e-07 $l=1.95e-07 $layer=LI1_cond $X=7.815 $Y=2.455
+ $X2=7.815 $Y2=2.65
r132 38 40 7.07246 $w=5.73e-07 $l=3.4e-07 $layer=LI1_cond $X=4.817 $Y=0.515
+ $X2=4.817 $Y2=0.855
r133 35 36 117.433 $w=1.68e-07 $l=1.8e-06 $layer=LI1_cond $X=8.705 $Y=0.765
+ $X2=8.705 $Y2=2.565
r134 34 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.015 $Y=0.68
+ $X2=7.93 $Y2=0.68
r135 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.62 $Y=0.68
+ $X2=8.705 $Y2=0.765
r136 33 34 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=8.62 $Y=0.68
+ $X2=8.015 $Y2=0.68
r137 32 49 2.85362 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.98 $Y=2.65
+ $X2=7.815 $Y2=2.65
r138 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.62 $Y=2.65
+ $X2=8.705 $Y2=2.565
r139 31 32 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=8.62 $Y=2.65
+ $X2=7.98 $Y2=2.65
r140 27 48 3.99587 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=2.37
+ $X2=7.815 $Y2=2.455
r141 27 29 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=7.815 $Y=2.37
+ $X2=7.815 $Y2=2.115
r142 26 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.94 $Y=0.855
+ $X2=6.815 $Y2=0.855
r143 25 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.845 $Y=0.855
+ $X2=7.93 $Y2=0.855
r144 25 26 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=7.845 $Y=0.855
+ $X2=6.94 $Y2=0.855
r145 21 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.815 $Y=0.77
+ $X2=6.815 $Y2=0.855
r146 21 23 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=6.815 $Y=0.77
+ $X2=6.815 $Y2=0.515
r147 20 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.945 $Y=2.455
+ $X2=5.86 $Y2=2.455
r148 19 48 2.85362 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.65 $Y=2.455
+ $X2=7.815 $Y2=2.455
r149 19 20 111.235 $w=1.68e-07 $l=1.705e-06 $layer=LI1_cond $X=7.65 $Y=2.455
+ $X2=5.945 $Y2=2.455
r150 18 40 8.04321 $w=1.7e-07 $l=2.88e-07 $layer=LI1_cond $X=5.105 $Y=0.855
+ $X2=4.817 $Y2=0.855
r151 17 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.69 $Y=0.855
+ $X2=6.815 $Y2=0.855
r152 17 18 103.406 $w=1.68e-07 $l=1.585e-06 $layer=LI1_cond $X=6.69 $Y=0.855
+ $X2=5.105 $Y2=0.855
r153 13 42 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=5.86 $Y=2.785
+ $X2=5.86 $Y2=2.455
r154 13 15 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=5.775 $Y=2.785
+ $X2=5.34 $Y2=2.785
r155 4 29 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=7.68
+ $Y=1.96 $X2=7.815 $Y2=2.115
r156 3 15 600 $w=1.7e-07 $l=9.03549e-07 $layer=licon1_PDIFF $count=1 $X=5.085
+ $Y=1.96 $X2=5.34 $Y2=2.745
r157 2 47 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=6.715
+ $Y=0.37 $X2=6.855 $Y2=0.855
r158 2 23 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.715
+ $Y=0.37 $X2=6.855 $Y2=0.515
r159 1 38 91 $w=1.7e-07 $l=3.75566e-07 $layer=licon1_NDIFF $count=2 $X=4.545
+ $Y=0.37 $X2=4.855 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_2%X 1 2 7 8 9 10 11 12 13 36
r22 34 36 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=9.825 $Y=1.995
+ $X2=9.825 $Y2=2.035
r23 12 13 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=9.825 $Y=2.405
+ $X2=9.825 $Y2=2.775
r24 11 34 0.75732 $w=3.48e-07 $l=2.3e-08 $layer=LI1_cond $X=9.825 $Y=1.972
+ $X2=9.825 $Y2=1.995
r25 11 45 5.05604 $w=3.48e-07 $l=1.52e-07 $layer=LI1_cond $X=9.825 $Y=1.972
+ $X2=9.825 $Y2=1.82
r26 11 12 11.4586 $w=3.48e-07 $l=3.48e-07 $layer=LI1_cond $X=9.825 $Y=2.057
+ $X2=9.825 $Y2=2.405
r27 11 36 0.724393 $w=3.48e-07 $l=2.2e-08 $layer=LI1_cond $X=9.825 $Y=2.057
+ $X2=9.825 $Y2=2.035
r28 10 45 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=9.815 $Y=1.665
+ $X2=9.815 $Y2=1.82
r29 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=9.815 $Y=1.295
+ $X2=9.815 $Y2=1.665
r30 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=9.815 $Y=0.925
+ $X2=9.815 $Y2=1.295
r31 8 27 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=9.815 $Y=0.925
+ $X2=9.815 $Y2=0.645
r32 7 27 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=9.815 $Y=0.555
+ $X2=9.815 $Y2=0.645
r33 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.7
+ $Y=1.84 $X2=9.835 $Y2=1.985
r34 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.7
+ $Y=1.84 $X2=9.835 $Y2=2.815
r35 1 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.675
+ $Y=0.5 $X2=9.815 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_2%VGND 1 2 3 4 5 18 24 28 32 34 36 39 40 42 43
+ 44 50 64 68 74 77 81
r91 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0 $X2=10.32
+ $Y2=0
r92 77 78 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r93 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r94 72 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=10.32
+ $Y2=0
r95 72 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r96 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r97 69 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.47 $Y=0 $X2=9.385
+ $Y2=0
r98 69 71 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.47 $Y=0 $X2=9.84
+ $Y2=0
r99 68 80 3.96842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=10.16 $Y=0 $X2=10.36
+ $Y2=0
r100 68 71 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=10.16 $Y=0 $X2=9.84
+ $Y2=0
r101 67 78 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=9.36 $Y2=0
r102 66 67 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r103 64 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.3 $Y=0 $X2=9.385
+ $Y2=0
r104 64 66 183.979 $w=1.68e-07 $l=2.82e-06 $layer=LI1_cond $X=9.3 $Y=0 $X2=6.48
+ $Y2=0
r105 63 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r106 62 63 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r107 60 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r108 59 62 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r109 59 60 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r110 57 74 11.015 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=3.925 $Y=0 $X2=3.685
+ $Y2=0
r111 57 59 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.925 $Y=0
+ $X2=4.08 $Y2=0
r112 56 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r113 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r114 53 56 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r115 52 55 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r116 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r117 50 74 11.015 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=3.445 $Y=0 $X2=3.685
+ $Y2=0
r118 50 55 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.445 $Y=0
+ $X2=3.12 $Y2=0
r119 48 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r120 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r121 44 63 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=0 $X2=6
+ $Y2=0
r122 44 60 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=5.28 $Y=0 $X2=4.08
+ $Y2=0
r123 42 62 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.14 $Y=0 $X2=6
+ $Y2=0
r124 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.14 $Y=0 $X2=6.305
+ $Y2=0
r125 41 66 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=6.47 $Y=0 $X2=6.48
+ $Y2=0
r126 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.47 $Y=0 $X2=6.305
+ $Y2=0
r127 39 47 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=0.72
+ $Y2=0
r128 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=0.985
+ $Y2=0
r129 38 52 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=1.15 $Y=0 $X2=1.2
+ $Y2=0
r130 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=0.985
+ $Y2=0
r131 34 80 3.17474 $w=2.5e-07 $l=1.16619e-07 $layer=LI1_cond $X=10.285 $Y=0.085
+ $X2=10.36 $Y2=0
r132 34 36 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=10.285 $Y=0.085
+ $X2=10.285 $Y2=0.645
r133 30 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.385 $Y=0.085
+ $X2=9.385 $Y2=0
r134 30 32 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=9.385 $Y=0.085
+ $X2=9.385 $Y2=0.675
r135 26 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.305 $Y=0.085
+ $X2=6.305 $Y2=0
r136 26 28 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.305 $Y=0.085
+ $X2=6.305 $Y2=0.515
r137 22 74 1.96841 $w=4.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=0.085
+ $X2=3.685 $Y2=0
r138 22 24 10.7149 $w=4.78e-07 $l=4.3e-07 $layer=LI1_cond $X=3.685 $Y=0.085
+ $X2=3.685 $Y2=0.515
r139 18 20 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.985 $Y=0.515
+ $X2=0.985 $Y2=0.855
r140 16 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.985 $Y=0.085
+ $X2=0.985 $Y2=0
r141 16 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.985 $Y=0.085
+ $X2=0.985 $Y2=0.515
r142 5 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.105
+ $Y=0.5 $X2=10.245 $Y2=0.645
r143 4 32 91 $w=1.7e-07 $l=6.36396e-07 $layer=licon1_NDIFF $count=2 $X=8.785
+ $Y=0.6 $X2=9.385 $Y2=0.675
r144 3 28 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.165
+ $Y=0.37 $X2=6.305 $Y2=0.515
r145 2 24 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=3.465
+ $Y=0.37 $X2=3.65 $Y2=0.515
r146 1 20 182 $w=1.7e-07 $l=5.55068e-07 $layer=licon1_NDIFF $count=1 $X=0.59
+ $Y=0.47 $X2=0.985 $Y2=0.855
r147 1 18 182 $w=1.7e-07 $l=4.16893e-07 $layer=licon1_NDIFF $count=1 $X=0.59
+ $Y=0.47 $X2=0.985 $Y2=0.515
.ends


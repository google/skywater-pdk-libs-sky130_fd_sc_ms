* File: sky130_fd_sc_ms__xnor3_4.pxi.spice
* Created: Fri Aug 28 18:18:40 2020
* 
x_PM_SKY130_FD_SC_MS__XNOR3_4%A_75_227# N_A_75_227#_M1003_d N_A_75_227#_M1009_d
+ N_A_75_227#_M1018_d N_A_75_227#_M1000_d N_A_75_227#_M1020_g
+ N_A_75_227#_M1016_g N_A_75_227#_c_188_n N_A_75_227#_c_189_n
+ N_A_75_227#_c_202_p N_A_75_227#_c_256_p N_A_75_227#_c_203_p
+ N_A_75_227#_c_198_n N_A_75_227#_c_207_p N_A_75_227#_c_199_n
+ N_A_75_227#_c_200_n N_A_75_227#_c_190_n N_A_75_227#_c_191_n
+ N_A_75_227#_c_192_n N_A_75_227#_c_193_n N_A_75_227#_c_194_n
+ N_A_75_227#_c_201_n N_A_75_227#_c_195_n PM_SKY130_FD_SC_MS__XNOR3_4%A_75_227#
x_PM_SKY130_FD_SC_MS__XNOR3_4%A N_A_M1018_g N_A_M1003_g A N_A_c_319_n
+ N_A_c_320_n PM_SKY130_FD_SC_MS__XNOR3_4%A
x_PM_SKY130_FD_SC_MS__XNOR3_4%A_386_23# N_A_386_23#_M1022_s N_A_386_23#_M1007_s
+ N_A_386_23#_M1006_g N_A_386_23#_c_363_n N_A_386_23#_c_364_n
+ N_A_386_23#_c_365_n N_A_386_23#_M1014_g N_A_386_23#_M1009_g
+ N_A_386_23#_M1000_g N_A_386_23#_c_368_n N_A_386_23#_c_369_n
+ N_A_386_23#_c_370_n N_A_386_23#_c_378_n N_A_386_23#_c_371_n
+ N_A_386_23#_c_372_n N_A_386_23#_c_379_n N_A_386_23#_c_380_n
+ N_A_386_23#_c_373_n PM_SKY130_FD_SC_MS__XNOR3_4%A_386_23#
x_PM_SKY130_FD_SC_MS__XNOR3_4%B N_B_M1024_g N_B_c_488_n N_B_M1025_g N_B_c_496_n
+ N_B_c_497_n N_B_M1005_g N_B_M1015_g N_B_c_499_n N_B_c_500_n N_B_M1022_g
+ N_B_M1007_g N_B_c_491_n N_B_c_503_n B N_B_c_492_n N_B_c_493_n
+ PM_SKY130_FD_SC_MS__XNOR3_4%B
x_PM_SKY130_FD_SC_MS__XNOR3_4%A_1024_300# N_A_1024_300#_M1017_s
+ N_A_1024_300#_M1012_s N_A_1024_300#_M1027_g N_A_1024_300#_M1021_g
+ N_A_1024_300#_c_621_n N_A_1024_300#_c_622_n N_A_1024_300#_c_629_n
+ N_A_1024_300#_c_623_n N_A_1024_300#_c_624_n N_A_1024_300#_c_625_n
+ N_A_1024_300#_c_626_n N_A_1024_300#_c_633_n
+ PM_SKY130_FD_SC_MS__XNOR3_4%A_1024_300#
x_PM_SKY130_FD_SC_MS__XNOR3_4%C N_C_M1010_g N_C_M1019_g N_C_c_708_n N_C_c_709_n
+ N_C_M1017_g N_C_M1012_g C N_C_c_710_n N_C_c_711_n N_C_c_712_n
+ PM_SKY130_FD_SC_MS__XNOR3_4%C
x_PM_SKY130_FD_SC_MS__XNOR3_4%A_1057_74# N_A_1057_74#_M1027_d
+ N_A_1057_74#_M1021_d N_A_1057_74#_M1002_g N_A_1057_74#_c_782_n
+ N_A_1057_74#_M1001_g N_A_1057_74#_M1008_g N_A_1057_74#_c_783_n
+ N_A_1057_74#_M1004_g N_A_1057_74#_M1023_g N_A_1057_74#_c_784_n
+ N_A_1057_74#_M1011_g N_A_1057_74#_c_785_n N_A_1057_74#_M1026_g
+ N_A_1057_74#_c_786_n N_A_1057_74#_M1013_g N_A_1057_74#_c_787_n
+ N_A_1057_74#_c_788_n N_A_1057_74#_c_789_n N_A_1057_74#_c_801_n
+ N_A_1057_74#_c_790_n N_A_1057_74#_c_791_n N_A_1057_74#_c_792_n
+ N_A_1057_74#_c_908_p N_A_1057_74#_c_822_n N_A_1057_74#_c_824_n
+ N_A_1057_74#_c_802_n N_A_1057_74#_c_793_n N_A_1057_74#_c_803_n
+ N_A_1057_74#_c_842_p N_A_1057_74#_c_804_n N_A_1057_74#_c_837_p
+ N_A_1057_74#_c_794_n N_A_1057_74#_c_795_n
+ PM_SKY130_FD_SC_MS__XNOR3_4%A_1057_74#
x_PM_SKY130_FD_SC_MS__XNOR3_4%A_27_373# N_A_27_373#_M1016_s N_A_27_373#_M1006_d
+ N_A_27_373#_M1020_s N_A_27_373#_M1014_d N_A_27_373#_c_941_n
+ N_A_27_373#_c_947_n N_A_27_373#_c_948_n N_A_27_373#_c_942_n
+ N_A_27_373#_c_949_n N_A_27_373#_c_943_n N_A_27_373#_c_944_n
+ N_A_27_373#_c_945_n N_A_27_373#_c_951_n N_A_27_373#_c_971_n
+ N_A_27_373#_c_978_n N_A_27_373#_c_981_n N_A_27_373#_c_946_n
+ N_A_27_373#_c_953_n PM_SKY130_FD_SC_MS__XNOR3_4%A_27_373#
x_PM_SKY130_FD_SC_MS__XNOR3_4%VPWR N_VPWR_M1020_d N_VPWR_M1007_d N_VPWR_M1012_d
+ N_VPWR_M1008_s N_VPWR_M1026_s N_VPWR_c_1049_n N_VPWR_c_1050_n N_VPWR_c_1051_n
+ N_VPWR_c_1052_n N_VPWR_c_1053_n N_VPWR_c_1054_n N_VPWR_c_1055_n
+ N_VPWR_c_1056_n N_VPWR_c_1118_n VPWR N_VPWR_c_1057_n N_VPWR_c_1058_n
+ N_VPWR_c_1059_n N_VPWR_c_1060_n N_VPWR_c_1061_n N_VPWR_c_1062_n
+ N_VPWR_c_1063_n N_VPWR_c_1064_n N_VPWR_c_1048_n
+ PM_SKY130_FD_SC_MS__XNOR3_4%VPWR
x_PM_SKY130_FD_SC_MS__XNOR3_4%A_327_373# N_A_327_373#_M1005_d
+ N_A_327_373#_M1010_d N_A_327_373#_M1025_d N_A_327_373#_M1021_s
+ N_A_327_373#_c_1163_n N_A_327_373#_c_1155_n N_A_327_373#_c_1156_n
+ N_A_327_373#_c_1157_n N_A_327_373#_c_1158_n N_A_327_373#_c_1159_n
+ N_A_327_373#_c_1160_n N_A_327_373#_c_1161_n N_A_327_373#_c_1180_n
+ N_A_327_373#_c_1162_n N_A_327_373#_c_1166_n N_A_327_373#_c_1190_n
+ N_A_327_373#_c_1167_n N_A_327_373#_c_1168_n N_A_327_373#_c_1191_n
+ PM_SKY130_FD_SC_MS__XNOR3_4%A_327_373#
x_PM_SKY130_FD_SC_MS__XNOR3_4%A_321_77# N_A_321_77#_M1024_d N_A_321_77#_M1027_s
+ N_A_321_77#_M1015_d N_A_321_77#_M1019_d N_A_321_77#_c_1283_n
+ N_A_321_77#_c_1310_n N_A_321_77#_c_1289_n N_A_321_77#_c_1300_n
+ N_A_321_77#_c_1284_n N_A_321_77#_c_1291_n N_A_321_77#_c_1292_n
+ N_A_321_77#_c_1285_n N_A_321_77#_c_1286_n N_A_321_77#_c_1287_n
+ N_A_321_77#_c_1288_n N_A_321_77#_c_1357_n
+ PM_SKY130_FD_SC_MS__XNOR3_4%A_321_77#
x_PM_SKY130_FD_SC_MS__XNOR3_4%X N_X_M1001_d N_X_M1011_d N_X_M1002_d N_X_M1023_d
+ N_X_c_1416_n N_X_c_1413_n N_X_c_1414_n N_X_c_1429_n N_X_c_1417_n N_X_c_1418_n
+ N_X_c_1439_n N_X_c_1442_n X X X X X X X X PM_SKY130_FD_SC_MS__XNOR3_4%X
x_PM_SKY130_FD_SC_MS__XNOR3_4%VGND N_VGND_M1016_d N_VGND_M1022_d N_VGND_M1017_d
+ N_VGND_M1004_s N_VGND_M1013_s N_VGND_c_1471_n N_VGND_c_1472_n N_VGND_c_1473_n
+ N_VGND_c_1523_n N_VGND_c_1474_n N_VGND_c_1475_n N_VGND_c_1476_n
+ N_VGND_c_1477_n N_VGND_c_1478_n VGND N_VGND_c_1479_n N_VGND_c_1480_n
+ N_VGND_c_1481_n N_VGND_c_1482_n N_VGND_c_1483_n N_VGND_c_1484_n
+ PM_SKY130_FD_SC_MS__XNOR3_4%VGND
cc_1 VNB N_A_75_227#_M1020_g 0.0109153f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.365
cc_2 VNB N_A_75_227#_c_188_n 0.00126892f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.95
cc_3 VNB N_A_75_227#_c_189_n 0.0202598f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=1.12
cc_4 VNB N_A_75_227#_c_190_n 0.00307726f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.34
cc_5 VNB N_A_75_227#_c_191_n 0.00348554f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.12
cc_6 VNB N_A_75_227#_c_192_n 0.0344865f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.3
cc_7 VNB N_A_75_227#_c_193_n 0.00538013f $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=0.36
cc_8 VNB N_A_75_227#_c_194_n 0.0120995f $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=0.35
cc_9 VNB N_A_75_227#_c_195_n 0.0210495f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.135
cc_10 VNB N_A_M1003_g 0.0285621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_c_319_n 0.0235519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_c_320_n 0.00424938f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_13 VNB N_A_386_23#_M1006_g 0.0336344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_386_23#_c_363_n 0.076486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_386_23#_c_364_n 0.0126012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_386_23#_c_365_n 0.0246406f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_17 VNB N_A_386_23#_M1014_g 0.00984973f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.365
cc_18 VNB N_A_386_23#_M1009_g 0.0355421f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.465
cc_19 VNB N_A_386_23#_c_368_n 0.00697882f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.72
cc_20 VNB N_A_386_23#_c_369_n 0.0259534f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=0.53
cc_21 VNB N_A_386_23#_c_370_n 0.00682553f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=2.99
cc_22 VNB N_A_386_23#_c_371_n 0.00457202f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.12
cc_23 VNB N_A_386_23#_c_372_n 2.44385e-19 $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.3
cc_24 VNB N_A_386_23#_c_373_n 9.51668e-19 $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=0.35
cc_25 VNB N_B_M1024_g 0.0423531f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.865
cc_26 VNB N_B_c_488_n 0.00197711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B_M1005_g 0.0281997f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_28 VNB N_B_M1022_g 0.0230134f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.035
cc_29 VNB N_B_c_491_n 0.00367469f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=0.53
cc_30 VNB N_B_c_492_n 0.00212715f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.3
cc_31 VNB N_B_c_493_n 0.0521732f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.3
cc_32 VNB N_A_1024_300#_M1027_g 0.0461186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_1024_300#_c_621_n 0.00616832f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.365
cc_34 VNB N_A_1024_300#_c_622_n 0.00342923f $X=-0.19 $Y=-0.245 $X2=0.545
+ $Y2=0.705
cc_35 VNB N_A_1024_300#_c_623_n 0.0175061f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.12
cc_36 VNB N_A_1024_300#_c_624_n 8.68163e-19 $X=-0.19 $Y=-0.245 $X2=0.705
+ $Y2=2.035
cc_37 VNB N_A_1024_300#_c_625_n 0.00169209f $X=-0.19 $Y=-0.245 $X2=1.23
+ $Y2=2.905
cc_38 VNB N_A_1024_300#_c_626_n 6.55071e-19 $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=0.425
cc_39 VNB N_C_M1010_g 0.0354923f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.865
cc_40 VNB N_C_M1019_g 0.0101334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_C_c_708_n 0.017148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_C_c_709_n 0.0214513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_C_c_710_n 0.04531f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.035
cc_44 VNB N_C_c_711_n 0.00271543f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.905
cc_45 VNB N_C_c_712_n 0.0308389f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.72
cc_46 VNB N_A_1057_74#_c_782_n 0.0199489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1057_74#_c_783_n 0.0157326f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.705
cc_48 VNB N_A_1057_74#_c_784_n 0.0156085f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.035
cc_49 VNB N_A_1057_74#_c_785_n 0.0816966f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.72
cc_50 VNB N_A_1057_74#_c_786_n 0.0188693f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=0.53
cc_51 VNB N_A_1057_74#_c_787_n 0.00252995f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.34
cc_52 VNB N_A_1057_74#_c_788_n 0.0159551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1057_74#_c_789_n 0.00425762f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.3
cc_54 VNB N_A_1057_74#_c_790_n 0.010379f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.035
cc_55 VNB N_A_1057_74#_c_791_n 0.00552332f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.035
cc_56 VNB N_A_1057_74#_c_792_n 0.00330549f $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=0.35
cc_57 VNB N_A_1057_74#_c_793_n 0.00511152f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1057_74#_c_794_n 0.00222251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1057_74#_c_795_n 0.0537622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_27_373#_c_941_n 0.00716946f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.365
cc_61 VNB N_A_27_373#_c_942_n 0.0244142f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.465
cc_62 VNB N_A_27_373#_c_943_n 0.0368156f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.035
cc_63 VNB N_A_27_373#_c_944_n 0.00352767f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.035
cc_64 VNB N_A_27_373#_c_945_n 0.00265022f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.72
cc_65 VNB N_A_27_373#_c_946_n 0.00139242f $X=-0.19 $Y=-0.245 $X2=3.365 $Y2=0.35
cc_66 VNB N_VPWR_c_1048_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_327_373#_c_1155_n 0.00693911f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.365
cc_68 VNB N_A_327_373#_c_1156_n 0.00253978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_327_373#_c_1157_n 0.00224367f $X=-0.19 $Y=-0.245 $X2=0.545
+ $Y2=0.705
cc_70 VNB N_A_327_373#_c_1158_n 0.00579396f $X=-0.19 $Y=-0.245 $X2=0.62
+ $Y2=1.465
cc_71 VNB N_A_327_373#_c_1159_n 0.00395107f $X=-0.19 $Y=-0.245 $X2=1.175
+ $Y2=1.12
cc_72 VNB N_A_327_373#_c_1160_n 0.00883735f $X=-0.19 $Y=-0.245 $X2=0.705
+ $Y2=1.12
cc_73 VNB N_A_327_373#_c_1161_n 0.00776468f $X=-0.19 $Y=-0.245 $X2=0.705
+ $Y2=2.035
cc_74 VNB N_A_327_373#_c_1162_n 0.00689628f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=0.53
cc_75 VNB N_A_321_77#_c_1283_n 0.0080413f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.365
cc_76 VNB N_A_321_77#_c_1284_n 0.0120329f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.035
cc_77 VNB N_A_321_77#_c_1285_n 6.15911e-19 $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=1.035
cc_78 VNB N_A_321_77#_c_1286_n 0.00292969f $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=0.34
cc_79 VNB N_A_321_77#_c_1287_n 2.71919e-19 $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.34
cc_80 VNB N_A_321_77#_c_1288_n 0.0234999f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.12
cc_81 VNB N_X_c_1413_n 0.00292847f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.705
cc_82 VNB N_X_c_1414_n 0.0010385f $X=-0.19 $Y=-0.245 $X2=1.175 $Y2=1.12
cc_83 VNB X 0.00279061f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=0.53
cc_84 VNB N_VGND_c_1471_n 0.00734311f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.465
cc_85 VNB N_VGND_c_1472_n 0.0123225f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.035
cc_86 VNB N_VGND_c_1473_n 0.0566559f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.12
cc_87 VNB N_VGND_c_1474_n 0.0198695f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=0.53
cc_88 VNB N_VGND_c_1475_n 0.043087f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=0.53
cc_89 VNB N_VGND_c_1476_n 0.0181352f $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=0.34
cc_90 VNB N_VGND_c_1477_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.12
cc_91 VNB N_VGND_c_1478_n 0.0540788f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.3
cc_92 VNB N_VGND_c_1479_n 0.0779513f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=2.035
cc_93 VNB N_VGND_c_1480_n 0.0197463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1481_n 0.0264817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1482_n 0.00631318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1483_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1484_n 0.537672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VPB N_A_75_227#_M1020_g 0.026576f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.365
cc_99 VPB N_A_75_227#_c_188_n 0.00162476f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.95
cc_100 VPB N_A_75_227#_c_198_n 0.00184277f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.72
cc_101 VPB N_A_75_227#_c_199_n 0.033478f $X=-0.19 $Y=1.66 $X2=3.35 $Y2=2.99
cc_102 VPB N_A_75_227#_c_200_n 0.00315353f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.99
cc_103 VPB N_A_75_227#_c_201_n 0.00854348f $X=-0.19 $Y=1.66 $X2=3.515 $Y2=2.795
cc_104 VPB N_A_M1018_g 0.0215752f $X=-0.19 $Y=1.66 $X2=1.095 $Y2=1.865
cc_105 VPB N_A_c_319_n 0.00725831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_c_320_n 0.00248131f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_107 VPB N_A_386_23#_M1014_g 0.0220735f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.365
cc_108 VPB N_A_386_23#_M1000_g 0.0218908f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.12
cc_109 VPB N_A_386_23#_c_368_n 0.00410146f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.72
cc_110 VPB N_A_386_23#_c_369_n 0.00696907f $X=-0.19 $Y=1.66 $X2=1.3 $Y2=0.53
cc_111 VPB N_A_386_23#_c_378_n 0.00170319f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.34
cc_112 VPB N_A_386_23#_c_379_n 7.04287e-19 $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.3
cc_113 VPB N_A_386_23#_c_380_n 0.00288617f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.035
cc_114 VPB N_B_c_488_n 0.00405898f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_B_M1025_g 0.0371456f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_B_c_496_n 0.0653192f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_B_c_497_n 0.0140967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_B_M1015_g 0.0466349f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=0.705
cc_119 VPB N_B_c_499_n 0.0773091f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=0.705
cc_120 VPB N_B_c_500_n 0.077957f $X=-0.19 $Y=1.66 $X2=1.175 $Y2=1.12
cc_121 VPB N_B_M1007_g 0.0251936f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.72
cc_122 VPB N_B_c_491_n 0.00987388f $X=-0.19 $Y=1.66 $X2=1.26 $Y2=0.53
cc_123 VPB N_B_c_503_n 0.00898883f $X=-0.19 $Y=1.66 $X2=3.35 $Y2=2.99
cc_124 VPB N_B_c_492_n 0.00285555f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.3
cc_125 VPB N_B_c_493_n 0.00742445f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.3
cc_126 VPB N_A_1024_300#_M1021_g 0.0255238f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_127 VPB N_A_1024_300#_c_621_n 0.0138344f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.365
cc_128 VPB N_A_1024_300#_c_629_n 0.00775309f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.465
cc_129 VPB N_A_1024_300#_c_623_n 0.0176763f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.12
cc_130 VPB N_A_1024_300#_c_624_n 0.0017048f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=2.035
cc_131 VPB N_A_1024_300#_c_626_n 0.00270666f $X=-0.19 $Y=1.66 $X2=1.3 $Y2=0.425
cc_132 VPB N_A_1024_300#_c_633_n 0.0145545f $X=-0.19 $Y=1.66 $X2=3.35 $Y2=2.99
cc_133 VPB N_C_M1019_g 0.0383915f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_C_M1012_g 0.0255442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_C_c_711_n 0.00242482f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.905
cc_136 VPB N_C_c_712_n 0.00858732f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.72
cc_137 VPB N_A_1057_74#_M1002_g 0.0249418f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_1057_74#_M1008_g 0.0211049f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_1057_74#_M1023_g 0.0211102f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.12
cc_140 VPB N_A_1057_74#_c_785_n 0.00888143f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.72
cc_141 VPB N_A_1057_74#_M1026_g 0.0266931f $X=-0.19 $Y=1.66 $X2=1.3 $Y2=0.425
cc_142 VPB N_A_1057_74#_c_801_n 0.0369347f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.3
cc_143 VPB N_A_1057_74#_c_802_n 0.0180252f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_1057_74#_c_803_n 0.00375044f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.135
cc_145 VPB N_A_1057_74#_c_804_n 0.00949407f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_1057_74#_c_795_n 0.0234566f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_27_373#_c_947_n 0.00835493f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.135
cc_148 VPB N_A_27_373#_c_948_n 9.77141e-19 $X=-0.19 $Y=1.66 $X2=0.545 $Y2=0.705
cc_149 VPB N_A_27_373#_c_949_n 0.00885838f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.12
cc_150 VPB N_A_27_373#_c_943_n 0.00903108f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=2.035
cc_151 VPB N_A_27_373#_c_951_n 0.00221377f $X=-0.19 $Y=1.66 $X2=3.35 $Y2=2.99
cc_152 VPB N_A_27_373#_c_946_n 0.00139038f $X=-0.19 $Y=1.66 $X2=3.365 $Y2=0.35
cc_153 VPB N_A_27_373#_c_953_n 0.0375448f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_1049_n 0.0110249f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=0.705
cc_155 VPB N_VPWR_c_1050_n 0.0135657f $X=-0.19 $Y=1.66 $X2=1.175 $Y2=1.12
cc_156 VPB N_VPWR_c_1051_n 0.0133031f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=2.035
cc_157 VPB N_VPWR_c_1052_n 0.0023761f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.72
cc_158 VPB N_VPWR_c_1053_n 0.0194151f $X=-0.19 $Y=1.66 $X2=1.3 $Y2=0.425
cc_159 VPB N_VPWR_c_1054_n 0.00959073f $X=-0.19 $Y=1.66 $X2=3.35 $Y2=2.99
cc_160 VPB N_VPWR_c_1055_n 0.0108116f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.12
cc_161 VPB N_VPWR_c_1056_n 0.0585007f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.3
cc_162 VPB N_VPWR_c_1057_n 0.0183206f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_1058_n 0.0861107f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_1059_n 0.0707383f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_1060_n 0.0204088f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_1061_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_1062_n 0.00612764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_1063_n 0.0119958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_1064_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_1048_n 0.106873f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_327_373#_c_1163_n 0.00150059f $X=-0.19 $Y=1.66 $X2=0.505
+ $Y2=2.365
cc_172 VPB N_A_327_373#_c_1155_n 0.00266963f $X=-0.19 $Y=1.66 $X2=0.505
+ $Y2=2.365
cc_173 VPB N_A_327_373#_c_1158_n 0.00644473f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.465
cc_174 VPB N_A_327_373#_c_1166_n 0.00346709f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.99
cc_175 VPB N_A_327_373#_c_1167_n 0.0028292f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.3
cc_176 VPB N_A_327_373#_c_1168_n 0.00746117f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.465
cc_177 VPB N_A_321_77#_c_1289_n 0.00349116f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.95
cc_178 VPB N_A_321_77#_c_1284_n 0.00361177f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=2.035
cc_179 VPB N_A_321_77#_c_1291_n 0.00837164f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=2.035
cc_180 VPB N_A_321_77#_c_1292_n 0.00198231f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.72
cc_181 VPB N_X_c_1416_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.365
cc_182 VPB N_X_c_1417_n 0.00112685f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.72
cc_183 VPB N_X_c_1418_n 0.00161134f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=2.72
cc_184 VPB X 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 N_A_75_227#_c_202_p N_A_M1018_g 0.0131143f $X=1.065 $Y=2.035 $X2=0 $Y2=0
cc_186 N_A_75_227#_c_203_p N_A_M1018_g 8.8334e-19 $X=1.23 $Y=2.12 $X2=0 $Y2=0
cc_187 N_A_75_227#_c_198_n N_A_M1018_g 0.0107347f $X=1.23 $Y=2.72 $X2=0 $Y2=0
cc_188 N_A_75_227#_c_200_n N_A_M1018_g 0.00278284f $X=1.395 $Y=2.99 $X2=0 $Y2=0
cc_189 N_A_75_227#_c_189_n N_A_M1003_g 0.0141792f $X=1.175 $Y=1.12 $X2=0 $Y2=0
cc_190 N_A_75_227#_c_207_p N_A_M1003_g 2.2106e-19 $X=1.26 $Y=0.53 $X2=0 $Y2=0
cc_191 N_A_75_227#_c_190_n N_A_M1003_g 0.00116563f $X=1.425 $Y=0.34 $X2=0 $Y2=0
cc_192 N_A_75_227#_c_191_n N_A_M1003_g 0.00121602f $X=0.58 $Y=1.12 $X2=0 $Y2=0
cc_193 N_A_75_227#_c_192_n N_A_M1003_g 0.0119439f $X=0.54 $Y=1.3 $X2=0 $Y2=0
cc_194 N_A_75_227#_c_195_n N_A_M1003_g 0.0203508f $X=0.54 $Y=1.135 $X2=0 $Y2=0
cc_195 N_A_75_227#_M1020_g N_A_c_319_n 0.0301445f $X=0.505 $Y=2.365 $X2=0 $Y2=0
cc_196 N_A_75_227#_c_188_n N_A_c_319_n 0.0054657f $X=0.62 $Y=1.95 $X2=0 $Y2=0
cc_197 N_A_75_227#_c_189_n N_A_c_319_n 0.00131516f $X=1.175 $Y=1.12 $X2=0 $Y2=0
cc_198 N_A_75_227#_c_203_p N_A_c_319_n 8.26292e-19 $X=1.23 $Y=2.12 $X2=0 $Y2=0
cc_199 N_A_75_227#_c_191_n N_A_c_319_n 3.13863e-19 $X=0.58 $Y=1.12 $X2=0 $Y2=0
cc_200 N_A_75_227#_c_192_n N_A_c_319_n 0.00548466f $X=0.54 $Y=1.3 $X2=0 $Y2=0
cc_201 N_A_75_227#_M1020_g N_A_c_320_n 3.40775e-19 $X=0.505 $Y=2.365 $X2=0 $Y2=0
cc_202 N_A_75_227#_c_189_n N_A_c_320_n 0.031511f $X=1.175 $Y=1.12 $X2=0 $Y2=0
cc_203 N_A_75_227#_c_202_p N_A_c_320_n 0.00978347f $X=1.065 $Y=2.035 $X2=0 $Y2=0
cc_204 N_A_75_227#_c_203_p N_A_c_320_n 0.0172715f $X=1.23 $Y=2.12 $X2=0 $Y2=0
cc_205 N_A_75_227#_c_191_n N_A_c_320_n 0.0261065f $X=0.58 $Y=1.12 $X2=0 $Y2=0
cc_206 N_A_75_227#_c_192_n N_A_c_320_n 3.13185e-19 $X=0.54 $Y=1.3 $X2=0 $Y2=0
cc_207 N_A_75_227#_c_194_n N_A_386_23#_M1006_g 0.00804191f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_208 N_A_75_227#_c_194_n N_A_386_23#_c_363_n 0.0211522f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_209 N_A_75_227#_c_194_n N_A_386_23#_c_364_n 0.00150581f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_210 N_A_75_227#_c_199_n N_A_386_23#_M1014_g 4.96104e-19 $X=3.35 $Y=2.99 $X2=0
+ $Y2=0
cc_211 N_A_75_227#_c_193_n N_A_386_23#_M1009_g 8.00488e-19 $X=3.365 $Y=0.36
+ $X2=0 $Y2=0
cc_212 N_A_75_227#_c_194_n N_A_386_23#_M1009_g 0.0115799f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_213 N_A_75_227#_c_199_n N_A_386_23#_M1000_g 0.00186626f $X=3.35 $Y=2.99 $X2=0
+ $Y2=0
cc_214 N_A_75_227#_c_201_n N_A_386_23#_M1000_g 0.00333964f $X=3.515 $Y=2.795
+ $X2=0 $Y2=0
cc_215 N_A_75_227#_M1000_d N_A_386_23#_c_378_n 0.00112074f $X=3.295 $Y=1.865
+ $X2=0 $Y2=0
cc_216 N_A_75_227#_M1000_d N_A_386_23#_c_379_n 0.00366545f $X=3.295 $Y=1.865
+ $X2=0 $Y2=0
cc_217 N_A_75_227#_c_189_n N_B_M1024_g 0.00470939f $X=1.175 $Y=1.12 $X2=0 $Y2=0
cc_218 N_A_75_227#_c_207_p N_B_M1024_g 2.28462e-19 $X=1.26 $Y=0.53 $X2=0 $Y2=0
cc_219 N_A_75_227#_c_194_n N_B_M1024_g 0.013294f $X=3.2 $Y=0.35 $X2=0 $Y2=0
cc_220 N_A_75_227#_c_203_p N_B_M1025_g 0.00130325f $X=1.23 $Y=2.12 $X2=0 $Y2=0
cc_221 N_A_75_227#_c_198_n N_B_M1025_g 0.0100498f $X=1.23 $Y=2.72 $X2=0 $Y2=0
cc_222 N_A_75_227#_c_199_n N_B_M1025_g 0.0172287f $X=3.35 $Y=2.99 $X2=0 $Y2=0
cc_223 N_A_75_227#_c_199_n N_B_c_496_n 0.0161324f $X=3.35 $Y=2.99 $X2=0 $Y2=0
cc_224 N_A_75_227#_c_194_n N_B_M1005_g 0.00112634f $X=3.2 $Y=0.35 $X2=0 $Y2=0
cc_225 N_A_75_227#_c_199_n N_B_M1015_g 0.0166569f $X=3.35 $Y=2.99 $X2=0 $Y2=0
cc_226 N_A_75_227#_c_201_n N_B_M1015_g 0.00237761f $X=3.515 $Y=2.795 $X2=0 $Y2=0
cc_227 N_A_75_227#_c_199_n N_B_c_499_n 0.00823287f $X=3.35 $Y=2.99 $X2=0 $Y2=0
cc_228 N_A_75_227#_c_201_n N_B_c_499_n 0.00899965f $X=3.515 $Y=2.795 $X2=0 $Y2=0
cc_229 N_A_75_227#_c_201_n N_B_c_500_n 0.0137088f $X=3.515 $Y=2.795 $X2=0 $Y2=0
cc_230 N_A_75_227#_c_193_n N_B_M1022_g 0.00356999f $X=3.365 $Y=0.36 $X2=0 $Y2=0
cc_231 N_A_75_227#_c_199_n N_A_27_373#_c_947_n 0.0382278f $X=3.35 $Y=2.99 $X2=0
+ $Y2=0
cc_232 N_A_75_227#_c_198_n N_A_27_373#_c_948_n 0.0140535f $X=1.23 $Y=2.72 $X2=0
+ $Y2=0
cc_233 N_A_75_227#_c_199_n N_A_27_373#_c_948_n 0.0151801f $X=3.35 $Y=2.99 $X2=0
+ $Y2=0
cc_234 N_A_75_227#_c_191_n N_A_27_373#_c_942_n 0.00252896f $X=0.58 $Y=1.12 $X2=0
+ $Y2=0
cc_235 N_A_75_227#_c_192_n N_A_27_373#_c_942_n 0.00237876f $X=0.54 $Y=1.3 $X2=0
+ $Y2=0
cc_236 N_A_75_227#_c_195_n N_A_27_373#_c_942_n 0.00804959f $X=0.54 $Y=1.135
+ $X2=0 $Y2=0
cc_237 N_A_75_227#_M1020_g N_A_27_373#_c_949_n 0.00145377f $X=0.505 $Y=2.365
+ $X2=0 $Y2=0
cc_238 N_A_75_227#_c_188_n N_A_27_373#_c_949_n 0.00464001f $X=0.62 $Y=1.95 $X2=0
+ $Y2=0
cc_239 N_A_75_227#_c_256_p N_A_27_373#_c_949_n 0.00868849f $X=0.705 $Y=2.035
+ $X2=0 $Y2=0
cc_240 N_A_75_227#_M1020_g N_A_27_373#_c_943_n 0.00829975f $X=0.505 $Y=2.365
+ $X2=0 $Y2=0
cc_241 N_A_75_227#_c_188_n N_A_27_373#_c_943_n 0.0206035f $X=0.62 $Y=1.95 $X2=0
+ $Y2=0
cc_242 N_A_75_227#_c_191_n N_A_27_373#_c_943_n 0.0324438f $X=0.58 $Y=1.12 $X2=0
+ $Y2=0
cc_243 N_A_75_227#_c_192_n N_A_27_373#_c_943_n 0.00816612f $X=0.54 $Y=1.3 $X2=0
+ $Y2=0
cc_244 N_A_75_227#_c_195_n N_A_27_373#_c_943_n 0.00650851f $X=0.54 $Y=1.135
+ $X2=0 $Y2=0
cc_245 N_A_75_227#_c_189_n N_A_27_373#_c_944_n 0.00352449f $X=1.175 $Y=1.12
+ $X2=0 $Y2=0
cc_246 N_A_75_227#_c_199_n N_A_27_373#_c_951_n 0.0310638f $X=3.35 $Y=2.99 $X2=0
+ $Y2=0
cc_247 N_A_75_227#_c_201_n N_A_27_373#_c_951_n 7.42656e-19 $X=3.515 $Y=2.795
+ $X2=0 $Y2=0
cc_248 N_A_75_227#_M1018_d N_A_27_373#_c_971_n 0.00456419f $X=1.095 $Y=1.865
+ $X2=0 $Y2=0
cc_249 N_A_75_227#_M1020_g N_A_27_373#_c_971_n 0.00758101f $X=0.505 $Y=2.365
+ $X2=0 $Y2=0
cc_250 N_A_75_227#_c_202_p N_A_27_373#_c_971_n 0.0252686f $X=1.065 $Y=2.035
+ $X2=0 $Y2=0
cc_251 N_A_75_227#_c_256_p N_A_27_373#_c_971_n 0.0131098f $X=0.705 $Y=2.035
+ $X2=0 $Y2=0
cc_252 N_A_75_227#_c_203_p N_A_27_373#_c_971_n 0.0302905f $X=1.23 $Y=2.12 $X2=0
+ $Y2=0
cc_253 N_A_75_227#_c_191_n N_A_27_373#_c_971_n 0.00231569f $X=0.58 $Y=1.12 $X2=0
+ $Y2=0
cc_254 N_A_75_227#_c_192_n N_A_27_373#_c_971_n 5.79437e-19 $X=0.54 $Y=1.3 $X2=0
+ $Y2=0
cc_255 N_A_75_227#_c_188_n N_A_27_373#_c_978_n 8.60777e-19 $X=0.62 $Y=1.95 $X2=0
+ $Y2=0
cc_256 N_A_75_227#_c_256_p N_A_27_373#_c_978_n 8.91026e-19 $X=0.705 $Y=2.035
+ $X2=0 $Y2=0
cc_257 N_A_75_227#_c_192_n N_A_27_373#_c_978_n 2.18873e-19 $X=0.54 $Y=1.3 $X2=0
+ $Y2=0
cc_258 N_A_75_227#_c_203_p N_A_27_373#_c_981_n 8.00194e-19 $X=1.23 $Y=2.12 $X2=0
+ $Y2=0
cc_259 N_A_75_227#_c_198_n N_A_27_373#_c_981_n 7.80159e-19 $X=1.23 $Y=2.72 $X2=0
+ $Y2=0
cc_260 N_A_75_227#_c_203_p N_A_27_373#_c_946_n 0.0116148f $X=1.23 $Y=2.12 $X2=0
+ $Y2=0
cc_261 N_A_75_227#_c_198_n N_A_27_373#_c_946_n 0.0329333f $X=1.23 $Y=2.72 $X2=0
+ $Y2=0
cc_262 N_A_75_227#_c_188_n N_VPWR_M1020_d 0.00100244f $X=0.62 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_263 N_A_75_227#_c_202_p N_VPWR_M1020_d 0.00741543f $X=1.065 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_264 N_A_75_227#_c_256_p N_VPWR_M1020_d 5.75445e-19 $X=0.705 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_265 N_A_75_227#_M1020_g N_VPWR_c_1049_n 0.0147945f $X=0.505 $Y=2.365 $X2=0
+ $Y2=0
cc_266 N_A_75_227#_c_202_p N_VPWR_c_1049_n 0.0111605f $X=1.065 $Y=2.035 $X2=0
+ $Y2=0
cc_267 N_A_75_227#_c_256_p N_VPWR_c_1049_n 0.0065014f $X=0.705 $Y=2.035 $X2=0
+ $Y2=0
cc_268 N_A_75_227#_c_198_n N_VPWR_c_1049_n 0.0246613f $X=1.23 $Y=2.72 $X2=0
+ $Y2=0
cc_269 N_A_75_227#_c_200_n N_VPWR_c_1049_n 0.0146281f $X=1.395 $Y=2.99 $X2=0
+ $Y2=0
cc_270 N_A_75_227#_M1020_g N_VPWR_c_1057_n 0.00509252f $X=0.505 $Y=2.365 $X2=0
+ $Y2=0
cc_271 N_A_75_227#_c_199_n N_VPWR_c_1058_n 0.124833f $X=3.35 $Y=2.99 $X2=0 $Y2=0
cc_272 N_A_75_227#_c_200_n N_VPWR_c_1058_n 0.0236566f $X=1.395 $Y=2.99 $X2=0
+ $Y2=0
cc_273 N_A_75_227#_c_201_n N_VPWR_c_1058_n 0.0213919f $X=3.515 $Y=2.795 $X2=0
+ $Y2=0
cc_274 N_A_75_227#_M1020_g N_VPWR_c_1048_n 0.00519404f $X=0.505 $Y=2.365 $X2=0
+ $Y2=0
cc_275 N_A_75_227#_c_199_n N_VPWR_c_1048_n 0.0656561f $X=3.35 $Y=2.99 $X2=0
+ $Y2=0
cc_276 N_A_75_227#_c_200_n N_VPWR_c_1048_n 0.0128296f $X=1.395 $Y=2.99 $X2=0
+ $Y2=0
cc_277 N_A_75_227#_c_201_n N_VPWR_c_1048_n 0.0110564f $X=3.515 $Y=2.795 $X2=0
+ $Y2=0
cc_278 N_A_75_227#_M1000_d N_A_327_373#_c_1166_n 0.00548304f $X=3.295 $Y=1.865
+ $X2=0 $Y2=0
cc_279 N_A_75_227#_c_194_n N_A_321_77#_M1024_d 0.00205163f $X=3.2 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_280 N_A_75_227#_M1009_d N_A_321_77#_c_1283_n 0.0106006f $X=3.145 $Y=0.605
+ $X2=0 $Y2=0
cc_281 N_A_75_227#_c_193_n N_A_321_77#_c_1283_n 0.0228577f $X=3.365 $Y=0.36
+ $X2=0 $Y2=0
cc_282 N_A_75_227#_c_194_n N_A_321_77#_c_1283_n 0.0252875f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_283 N_A_75_227#_M1000_d N_A_321_77#_c_1289_n 0.00868909f $X=3.295 $Y=1.865
+ $X2=0 $Y2=0
cc_284 N_A_75_227#_c_199_n N_A_321_77#_c_1289_n 0.00653918f $X=3.35 $Y=2.99
+ $X2=0 $Y2=0
cc_285 N_A_75_227#_c_201_n N_A_321_77#_c_1289_n 0.0240938f $X=3.515 $Y=2.795
+ $X2=0 $Y2=0
cc_286 N_A_75_227#_c_199_n N_A_321_77#_c_1300_n 0.00918631f $X=3.35 $Y=2.99
+ $X2=0 $Y2=0
cc_287 N_A_75_227#_c_194_n N_A_321_77#_c_1285_n 0.0214403f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_288 N_A_75_227#_c_194_n N_A_321_77#_c_1286_n 0.0532333f $X=3.2 $Y=0.35 $X2=0
+ $Y2=0
cc_289 N_A_75_227#_c_189_n N_VGND_c_1471_n 0.0211827f $X=1.175 $Y=1.12 $X2=0
+ $Y2=0
cc_290 N_A_75_227#_c_190_n N_VGND_c_1471_n 0.0118948f $X=1.425 $Y=0.34 $X2=0
+ $Y2=0
cc_291 N_A_75_227#_c_191_n N_VGND_c_1471_n 0.00299742f $X=0.58 $Y=1.12 $X2=0
+ $Y2=0
cc_292 N_A_75_227#_c_192_n N_VGND_c_1471_n 2.06276e-19 $X=0.54 $Y=1.3 $X2=0
+ $Y2=0
cc_293 N_A_75_227#_c_195_n N_VGND_c_1471_n 0.00578941f $X=0.54 $Y=1.135 $X2=0
+ $Y2=0
cc_294 N_A_75_227#_c_190_n N_VGND_c_1479_n 0.0179217f $X=1.425 $Y=0.34 $X2=0
+ $Y2=0
cc_295 N_A_75_227#_c_194_n N_VGND_c_1479_n 0.131374f $X=3.2 $Y=0.35 $X2=0 $Y2=0
cc_296 N_A_75_227#_c_195_n N_VGND_c_1481_n 0.00540915f $X=0.54 $Y=1.135 $X2=0
+ $Y2=0
cc_297 N_A_75_227#_M1009_d N_VGND_c_1484_n 0.00251887f $X=3.145 $Y=0.605 $X2=0
+ $Y2=0
cc_298 N_A_75_227#_c_190_n N_VGND_c_1484_n 0.00971942f $X=1.425 $Y=0.34 $X2=0
+ $Y2=0
cc_299 N_A_75_227#_c_194_n N_VGND_c_1484_n 0.0734849f $X=3.2 $Y=0.35 $X2=0 $Y2=0
cc_300 N_A_75_227#_c_195_n N_VGND_c_1484_n 0.0054106f $X=0.54 $Y=1.135 $X2=0
+ $Y2=0
cc_301 N_A_M1003_g N_B_M1024_g 0.0160975f $X=1.045 $Y=0.705 $X2=0 $Y2=0
cc_302 N_A_c_319_n N_B_M1024_g 0.0194584f $X=1.08 $Y=1.54 $X2=0 $Y2=0
cc_303 N_A_c_320_n N_B_M1024_g 0.00287638f $X=1.08 $Y=1.54 $X2=0 $Y2=0
cc_304 N_A_M1018_g N_B_c_488_n 0.0233156f $X=1.005 $Y=2.365 $X2=0 $Y2=0
cc_305 N_A_M1003_g N_A_27_373#_c_944_n 8.13749e-19 $X=1.045 $Y=0.705 $X2=0 $Y2=0
cc_306 N_A_c_320_n N_A_27_373#_c_944_n 0.00584677f $X=1.08 $Y=1.54 $X2=0 $Y2=0
cc_307 N_A_c_320_n N_A_27_373#_c_971_n 0.00309875f $X=1.08 $Y=1.54 $X2=0 $Y2=0
cc_308 N_A_M1018_g N_A_27_373#_c_946_n 7.76325e-19 $X=1.005 $Y=2.365 $X2=0 $Y2=0
cc_309 N_A_c_319_n N_A_27_373#_c_946_n 2.1885e-19 $X=1.08 $Y=1.54 $X2=0 $Y2=0
cc_310 N_A_c_320_n N_A_27_373#_c_946_n 0.0176914f $X=1.08 $Y=1.54 $X2=0 $Y2=0
cc_311 N_A_M1018_g N_VPWR_c_1049_n 0.00113744f $X=1.005 $Y=2.365 $X2=0 $Y2=0
cc_312 N_A_M1018_g N_VPWR_c_1058_n 0.00525897f $X=1.005 $Y=2.365 $X2=0 $Y2=0
cc_313 N_A_M1018_g N_VPWR_c_1048_n 0.00515964f $X=1.005 $Y=2.365 $X2=0 $Y2=0
cc_314 N_A_M1003_g N_VGND_c_1471_n 0.00984806f $X=1.045 $Y=0.705 $X2=0 $Y2=0
cc_315 N_A_M1003_g N_VGND_c_1479_n 0.00471276f $X=1.045 $Y=0.705 $X2=0 $Y2=0
cc_316 N_A_M1003_g N_VGND_c_1484_n 0.0045449f $X=1.045 $Y=0.705 $X2=0 $Y2=0
cc_317 N_A_386_23#_c_364_n N_B_M1024_g 0.0305639f $X=2.08 $Y=0.19 $X2=0 $Y2=0
cc_318 N_A_386_23#_M1014_g N_B_M1024_g 0.00272004f $X=2.245 $Y=2.185 $X2=0 $Y2=0
cc_319 N_A_386_23#_M1014_g N_B_c_488_n 0.0147746f $X=2.245 $Y=2.185 $X2=0 $Y2=0
cc_320 N_A_386_23#_M1014_g N_B_c_496_n 0.00376558f $X=2.245 $Y=2.185 $X2=0 $Y2=0
cc_321 N_A_386_23#_M1006_g N_B_M1005_g 0.017105f $X=2.005 $Y=0.815 $X2=0 $Y2=0
cc_322 N_A_386_23#_c_363_n N_B_M1005_g 0.00976806f $X=2.995 $Y=0.19 $X2=0 $Y2=0
cc_323 N_A_386_23#_c_365_n N_B_M1005_g 0.0149589f $X=2.245 $Y=1.47 $X2=0 $Y2=0
cc_324 N_A_386_23#_M1009_g N_B_M1005_g 0.0325534f $X=3.07 $Y=0.925 $X2=0 $Y2=0
cc_325 N_A_386_23#_c_368_n N_B_M1005_g 3.10708e-19 $X=3.6 $Y=1.54 $X2=0 $Y2=0
cc_326 N_A_386_23#_M1014_g N_B_M1015_g 0.025379f $X=2.245 $Y=2.185 $X2=0 $Y2=0
cc_327 N_A_386_23#_M1000_g N_B_c_499_n 0.00885431f $X=3.205 $Y=2.285 $X2=0 $Y2=0
cc_328 N_A_386_23#_M1000_g N_B_c_500_n 0.0287371f $X=3.205 $Y=2.285 $X2=0 $Y2=0
cc_329 N_A_386_23#_c_378_n N_B_c_500_n 0.00680454f $X=3.685 $Y=1.95 $X2=0 $Y2=0
cc_330 N_A_386_23#_c_379_n N_B_c_500_n 0.00388903f $X=3.77 $Y=2.075 $X2=0 $Y2=0
cc_331 N_A_386_23#_c_380_n N_B_c_500_n 0.0127273f $X=4.105 $Y=2.115 $X2=0 $Y2=0
cc_332 N_A_386_23#_c_373_n N_B_c_500_n 6.38429e-19 $X=3.685 $Y=1.54 $X2=0 $Y2=0
cc_333 N_A_386_23#_c_370_n N_B_M1022_g 0.00370096f $X=3.685 $Y=1.375 $X2=0 $Y2=0
cc_334 N_A_386_23#_c_372_n N_B_M1022_g 0.00328266f $X=3.925 $Y=1.04 $X2=0 $Y2=0
cc_335 N_A_386_23#_c_378_n N_B_M1007_g 5.41419e-19 $X=3.685 $Y=1.95 $X2=0 $Y2=0
cc_336 N_A_386_23#_c_380_n N_B_M1007_g 0.00319938f $X=4.105 $Y=2.115 $X2=0 $Y2=0
cc_337 N_A_386_23#_M1014_g N_B_c_491_n 0.0149589f $X=2.245 $Y=2.185 $X2=0 $Y2=0
cc_338 N_A_386_23#_M1000_g N_B_c_491_n 0.0186813f $X=3.205 $Y=2.285 $X2=0 $Y2=0
cc_339 N_A_386_23#_c_368_n N_B_c_491_n 3.16617e-19 $X=3.6 $Y=1.54 $X2=0 $Y2=0
cc_340 N_A_386_23#_c_369_n N_B_c_491_n 0.0040067f $X=3.16 $Y=1.54 $X2=0 $Y2=0
cc_341 N_A_386_23#_c_370_n N_B_c_492_n 0.00184128f $X=3.685 $Y=1.375 $X2=0 $Y2=0
cc_342 N_A_386_23#_c_378_n N_B_c_492_n 0.00562831f $X=3.685 $Y=1.95 $X2=0 $Y2=0
cc_343 N_A_386_23#_c_372_n N_B_c_492_n 0.00730998f $X=3.925 $Y=1.04 $X2=0 $Y2=0
cc_344 N_A_386_23#_c_380_n N_B_c_492_n 0.0219714f $X=4.105 $Y=2.115 $X2=0 $Y2=0
cc_345 N_A_386_23#_c_373_n N_B_c_492_n 0.0271008f $X=3.685 $Y=1.54 $X2=0 $Y2=0
cc_346 N_A_386_23#_c_369_n N_B_c_493_n 0.00670177f $X=3.16 $Y=1.54 $X2=0 $Y2=0
cc_347 N_A_386_23#_c_370_n N_B_c_493_n 6.03443e-19 $X=3.685 $Y=1.375 $X2=0 $Y2=0
cc_348 N_A_386_23#_c_372_n N_B_c_493_n 0.00616553f $X=3.925 $Y=1.04 $X2=0 $Y2=0
cc_349 N_A_386_23#_c_380_n N_B_c_493_n 9.75753e-19 $X=4.105 $Y=2.115 $X2=0 $Y2=0
cc_350 N_A_386_23#_c_373_n N_B_c_493_n 0.00765257f $X=3.685 $Y=1.54 $X2=0 $Y2=0
cc_351 N_A_386_23#_M1006_g N_A_27_373#_c_941_n 0.00779425f $X=2.005 $Y=0.815
+ $X2=0 $Y2=0
cc_352 N_A_386_23#_c_365_n N_A_27_373#_c_941_n 0.00339009f $X=2.245 $Y=1.47
+ $X2=0 $Y2=0
cc_353 N_A_386_23#_M1014_g N_A_27_373#_c_947_n 0.00705621f $X=2.245 $Y=2.185
+ $X2=0 $Y2=0
cc_354 N_A_386_23#_c_365_n N_A_27_373#_c_944_n 0.00307815f $X=2.245 $Y=1.47
+ $X2=0 $Y2=0
cc_355 N_A_386_23#_M1006_g N_A_27_373#_c_945_n 0.0046962f $X=2.005 $Y=0.815
+ $X2=0 $Y2=0
cc_356 N_A_386_23#_c_365_n N_A_27_373#_c_945_n 0.00729644f $X=2.245 $Y=1.47
+ $X2=0 $Y2=0
cc_357 N_A_386_23#_M1014_g N_A_27_373#_c_951_n 0.00828963f $X=2.245 $Y=2.185
+ $X2=0 $Y2=0
cc_358 N_A_386_23#_M1000_g N_A_27_373#_c_951_n 9.113e-19 $X=3.205 $Y=2.285 $X2=0
+ $Y2=0
cc_359 N_A_386_23#_M1014_g N_A_27_373#_c_946_n 0.00629315f $X=2.245 $Y=2.185
+ $X2=0 $Y2=0
cc_360 N_A_386_23#_M1014_g N_A_327_373#_c_1163_n 0.00909372f $X=2.245 $Y=2.185
+ $X2=0 $Y2=0
cc_361 N_A_386_23#_M1014_g N_A_327_373#_c_1155_n 0.00586623f $X=2.245 $Y=2.185
+ $X2=0 $Y2=0
cc_362 N_A_386_23#_c_368_n N_A_327_373#_c_1155_n 0.0115248f $X=3.6 $Y=1.54 $X2=0
+ $Y2=0
cc_363 N_A_386_23#_c_369_n N_A_327_373#_c_1155_n 6.38604e-19 $X=3.16 $Y=1.54
+ $X2=0 $Y2=0
cc_364 N_A_386_23#_c_365_n N_A_327_373#_c_1156_n 0.00642326f $X=2.245 $Y=1.47
+ $X2=0 $Y2=0
cc_365 N_A_386_23#_M1014_g N_A_327_373#_c_1156_n 0.00506743f $X=2.245 $Y=2.185
+ $X2=0 $Y2=0
cc_366 N_A_386_23#_c_365_n N_A_327_373#_c_1157_n 0.0012074f $X=2.245 $Y=1.47
+ $X2=0 $Y2=0
cc_367 N_A_386_23#_M1009_g N_A_327_373#_c_1157_n 0.00329076f $X=3.07 $Y=0.925
+ $X2=0 $Y2=0
cc_368 N_A_386_23#_c_368_n N_A_327_373#_c_1157_n 0.00801193f $X=3.6 $Y=1.54
+ $X2=0 $Y2=0
cc_369 N_A_386_23#_c_369_n N_A_327_373#_c_1157_n 4.48181e-19 $X=3.16 $Y=1.54
+ $X2=0 $Y2=0
cc_370 N_A_386_23#_M1009_g N_A_327_373#_c_1180_n 0.00577182f $X=3.07 $Y=0.925
+ $X2=0 $Y2=0
cc_371 N_A_386_23#_c_368_n N_A_327_373#_c_1180_n 0.00180109f $X=3.6 $Y=1.54
+ $X2=0 $Y2=0
cc_372 N_A_386_23#_c_370_n N_A_327_373#_c_1180_n 0.00238919f $X=3.685 $Y=1.375
+ $X2=0 $Y2=0
cc_373 N_A_386_23#_c_371_n N_A_327_373#_c_1180_n 0.00562748f $X=3.77 $Y=1.04
+ $X2=0 $Y2=0
cc_374 N_A_386_23#_M1014_g N_A_327_373#_c_1166_n 0.00139773f $X=2.245 $Y=2.185
+ $X2=0 $Y2=0
cc_375 N_A_386_23#_M1000_g N_A_327_373#_c_1166_n 0.00456556f $X=3.205 $Y=2.285
+ $X2=0 $Y2=0
cc_376 N_A_386_23#_c_368_n N_A_327_373#_c_1166_n 0.013588f $X=3.6 $Y=1.54 $X2=0
+ $Y2=0
cc_377 N_A_386_23#_c_369_n N_A_327_373#_c_1166_n 6.86671e-19 $X=3.16 $Y=1.54
+ $X2=0 $Y2=0
cc_378 N_A_386_23#_c_379_n N_A_327_373#_c_1166_n 0.0167115f $X=3.77 $Y=2.075
+ $X2=0 $Y2=0
cc_379 N_A_386_23#_c_380_n N_A_327_373#_c_1166_n 0.0259468f $X=4.105 $Y=2.115
+ $X2=0 $Y2=0
cc_380 N_A_386_23#_M1014_g N_A_327_373#_c_1190_n 0.0035026f $X=2.245 $Y=2.185
+ $X2=0 $Y2=0
cc_381 N_A_386_23#_M1014_g N_A_327_373#_c_1191_n 0.0045785f $X=2.245 $Y=2.185
+ $X2=0 $Y2=0
cc_382 N_A_386_23#_M1022_s N_A_321_77#_c_1283_n 0.00721616f $X=3.78 $Y=0.445
+ $X2=0 $Y2=0
cc_383 N_A_386_23#_c_363_n N_A_321_77#_c_1283_n 8.21484e-19 $X=2.995 $Y=0.19
+ $X2=0 $Y2=0
cc_384 N_A_386_23#_M1009_g N_A_321_77#_c_1283_n 0.0143626f $X=3.07 $Y=0.925
+ $X2=0 $Y2=0
cc_385 N_A_386_23#_c_368_n N_A_321_77#_c_1283_n 0.0162608f $X=3.6 $Y=1.54 $X2=0
+ $Y2=0
cc_386 N_A_386_23#_c_369_n N_A_321_77#_c_1283_n 0.00312277f $X=3.16 $Y=1.54
+ $X2=0 $Y2=0
cc_387 N_A_386_23#_c_371_n N_A_321_77#_c_1283_n 0.0143583f $X=3.77 $Y=1.04 $X2=0
+ $Y2=0
cc_388 N_A_386_23#_c_372_n N_A_321_77#_c_1283_n 0.0189364f $X=3.925 $Y=1.04
+ $X2=0 $Y2=0
cc_389 N_A_386_23#_M1000_g N_A_321_77#_c_1310_n 0.00906853f $X=3.205 $Y=2.285
+ $X2=0 $Y2=0
cc_390 N_A_386_23#_c_368_n N_A_321_77#_c_1310_n 0.00876312f $X=3.6 $Y=1.54 $X2=0
+ $Y2=0
cc_391 N_A_386_23#_c_369_n N_A_321_77#_c_1310_n 0.00309197f $X=3.16 $Y=1.54
+ $X2=0 $Y2=0
cc_392 N_A_386_23#_c_378_n N_A_321_77#_c_1310_n 0.00251211f $X=3.685 $Y=1.95
+ $X2=0 $Y2=0
cc_393 N_A_386_23#_c_379_n N_A_321_77#_c_1310_n 0.00707159f $X=3.77 $Y=2.075
+ $X2=0 $Y2=0
cc_394 N_A_386_23#_M1007_s N_A_321_77#_c_1289_n 0.00639138f $X=3.96 $Y=1.84
+ $X2=0 $Y2=0
cc_395 N_A_386_23#_M1000_g N_A_321_77#_c_1289_n 0.0113388f $X=3.205 $Y=2.285
+ $X2=0 $Y2=0
cc_396 N_A_386_23#_c_368_n N_A_321_77#_c_1289_n 0.00438203f $X=3.6 $Y=1.54 $X2=0
+ $Y2=0
cc_397 N_A_386_23#_c_379_n N_A_321_77#_c_1289_n 0.0129068f $X=3.77 $Y=2.075
+ $X2=0 $Y2=0
cc_398 N_A_386_23#_c_380_n N_A_321_77#_c_1289_n 0.03012f $X=4.105 $Y=2.115 $X2=0
+ $Y2=0
cc_399 N_A_386_23#_M1000_g N_A_321_77#_c_1300_n 0.00100437f $X=3.205 $Y=2.285
+ $X2=0 $Y2=0
cc_400 N_A_386_23#_c_370_n N_A_321_77#_c_1284_n 0.00632457f $X=3.685 $Y=1.375
+ $X2=0 $Y2=0
cc_401 N_A_386_23#_c_378_n N_A_321_77#_c_1284_n 0.00265176f $X=3.685 $Y=1.95
+ $X2=0 $Y2=0
cc_402 N_A_386_23#_c_372_n N_A_321_77#_c_1284_n 0.00409526f $X=3.925 $Y=1.04
+ $X2=0 $Y2=0
cc_403 N_A_386_23#_c_380_n N_A_321_77#_c_1284_n 0.0116478f $X=4.105 $Y=2.115
+ $X2=0 $Y2=0
cc_404 N_A_386_23#_M1006_g N_A_321_77#_c_1285_n 0.00590709f $X=2.005 $Y=0.815
+ $X2=0 $Y2=0
cc_405 N_A_386_23#_M1006_g N_A_321_77#_c_1286_n 0.00973001f $X=2.005 $Y=0.815
+ $X2=0 $Y2=0
cc_406 N_A_386_23#_c_363_n N_A_321_77#_c_1286_n 0.00193544f $X=2.995 $Y=0.19
+ $X2=0 $Y2=0
cc_407 N_A_386_23#_c_365_n N_A_321_77#_c_1286_n 6.20408e-19 $X=2.245 $Y=1.47
+ $X2=0 $Y2=0
cc_408 N_A_386_23#_M1009_g N_A_321_77#_c_1287_n 2.29766e-19 $X=3.07 $Y=0.925
+ $X2=0 $Y2=0
cc_409 N_A_386_23#_c_372_n N_A_321_77#_c_1288_n 0.00363019f $X=3.925 $Y=1.04
+ $X2=0 $Y2=0
cc_410 N_A_386_23#_c_364_n N_VGND_c_1479_n 0.0257161f $X=2.08 $Y=0.19 $X2=0
+ $Y2=0
cc_411 N_A_386_23#_c_363_n N_VGND_c_1484_n 0.0275023f $X=2.995 $Y=0.19 $X2=0
+ $Y2=0
cc_412 N_A_386_23#_c_364_n N_VGND_c_1484_n 0.00588169f $X=2.08 $Y=0.19 $X2=0
+ $Y2=0
cc_413 N_B_c_493_n N_A_1024_300#_M1027_g 0.00132172f $X=4.14 $Y=1.515 $X2=0
+ $Y2=0
cc_414 N_B_c_493_n N_A_1024_300#_c_623_n 0.00311263f $X=4.14 $Y=1.515 $X2=0
+ $Y2=0
cc_415 N_B_M1015_g N_A_27_373#_c_947_n 3.84395e-19 $X=2.695 $Y=2.185 $X2=0 $Y2=0
cc_416 N_B_M1025_g N_A_27_373#_c_948_n 0.00700455f $X=1.545 $Y=2.285 $X2=0 $Y2=0
cc_417 N_B_M1024_g N_A_27_373#_c_944_n 0.0103289f $X=1.53 $Y=0.705 $X2=0 $Y2=0
cc_418 N_B_M1005_g N_A_27_373#_c_945_n 0.00447538f $X=2.62 $Y=0.925 $X2=0 $Y2=0
cc_419 N_B_M1025_g N_A_27_373#_c_951_n 4.55728e-19 $X=1.545 $Y=2.285 $X2=0 $Y2=0
cc_420 N_B_M1015_g N_A_27_373#_c_951_n 0.0177308f $X=2.695 $Y=2.185 $X2=0 $Y2=0
cc_421 N_B_c_491_n N_A_27_373#_c_951_n 0.00104103f $X=2.665 $Y=1.79 $X2=0 $Y2=0
cc_422 N_B_M1025_g N_A_27_373#_c_971_n 0.00757288f $X=1.545 $Y=2.285 $X2=0 $Y2=0
cc_423 N_B_M1025_g N_A_27_373#_c_981_n 0.00367312f $X=1.545 $Y=2.285 $X2=0 $Y2=0
cc_424 N_B_M1024_g N_A_27_373#_c_946_n 0.00413342f $X=1.53 $Y=0.705 $X2=0 $Y2=0
cc_425 N_B_c_488_n N_A_27_373#_c_946_n 0.00310984f $X=1.545 $Y=1.73 $X2=0 $Y2=0
cc_426 N_B_M1025_g N_A_27_373#_c_946_n 0.0221464f $X=1.545 $Y=2.285 $X2=0 $Y2=0
cc_427 N_B_M1025_g N_VPWR_c_1049_n 2.98118e-19 $X=1.545 $Y=2.285 $X2=0 $Y2=0
cc_428 N_B_c_497_n N_VPWR_c_1049_n 0.00248898f $X=1.635 $Y=3.15 $X2=0 $Y2=0
cc_429 N_B_c_499_n N_VPWR_c_1050_n 0.00232909f $X=3.735 $Y=3.15 $X2=0 $Y2=0
cc_430 N_B_c_500_n N_VPWR_c_1050_n 0.00164526f $X=3.81 $Y=3.075 $X2=0 $Y2=0
cc_431 N_B_M1007_g N_VPWR_c_1050_n 0.0109706f $X=4.33 $Y=2.4 $X2=0 $Y2=0
cc_432 N_B_c_497_n N_VPWR_c_1058_n 0.0552122f $X=1.635 $Y=3.15 $X2=0 $Y2=0
cc_433 N_B_M1007_g N_VPWR_c_1058_n 0.00460063f $X=4.33 $Y=2.4 $X2=0 $Y2=0
cc_434 N_B_c_496_n N_VPWR_c_1048_n 0.0228018f $X=2.605 $Y=3.15 $X2=0 $Y2=0
cc_435 N_B_c_497_n N_VPWR_c_1048_n 0.00678686f $X=1.635 $Y=3.15 $X2=0 $Y2=0
cc_436 N_B_c_499_n N_VPWR_c_1048_n 0.0296833f $X=3.735 $Y=3.15 $X2=0 $Y2=0
cc_437 N_B_M1007_g N_VPWR_c_1048_n 0.0044909f $X=4.33 $Y=2.4 $X2=0 $Y2=0
cc_438 N_B_c_503_n N_VPWR_c_1048_n 0.00445015f $X=2.695 $Y=3.15 $X2=0 $Y2=0
cc_439 N_B_c_488_n N_A_327_373#_c_1163_n 8.6743e-19 $X=1.545 $Y=1.73 $X2=0 $Y2=0
cc_440 N_B_M1015_g N_A_327_373#_c_1163_n 8.15169e-19 $X=2.695 $Y=2.185 $X2=0
+ $Y2=0
cc_441 N_B_c_491_n N_A_327_373#_c_1163_n 6.44081e-19 $X=2.665 $Y=1.79 $X2=0
+ $Y2=0
cc_442 N_B_M1005_g N_A_327_373#_c_1155_n 0.00418594f $X=2.62 $Y=0.925 $X2=0
+ $Y2=0
cc_443 N_B_c_491_n N_A_327_373#_c_1155_n 0.00730111f $X=2.665 $Y=1.79 $X2=0
+ $Y2=0
cc_444 N_B_M1024_g N_A_327_373#_c_1156_n 4.38234e-19 $X=1.53 $Y=0.705 $X2=0
+ $Y2=0
cc_445 N_B_M1005_g N_A_327_373#_c_1157_n 0.00852261f $X=2.62 $Y=0.925 $X2=0
+ $Y2=0
cc_446 N_B_M1005_g N_A_327_373#_c_1180_n 0.00689469f $X=2.62 $Y=0.925 $X2=0
+ $Y2=0
cc_447 N_B_c_491_n N_A_327_373#_c_1180_n 0.00114318f $X=2.665 $Y=1.79 $X2=0
+ $Y2=0
cc_448 N_B_M1015_g N_A_327_373#_c_1166_n 0.00806577f $X=2.695 $Y=2.185 $X2=0
+ $Y2=0
cc_449 N_B_M1007_g N_A_327_373#_c_1166_n 0.00992633f $X=4.33 $Y=2.4 $X2=0 $Y2=0
cc_450 N_B_c_491_n N_A_327_373#_c_1166_n 0.00166648f $X=2.665 $Y=1.79 $X2=0
+ $Y2=0
cc_451 N_B_c_492_n N_A_327_373#_c_1166_n 0.00263253f $X=4.105 $Y=1.515 $X2=0
+ $Y2=0
cc_452 N_B_M1015_g N_A_327_373#_c_1190_n 4.65092e-19 $X=2.695 $Y=2.185 $X2=0
+ $Y2=0
cc_453 N_B_M1025_g N_A_327_373#_c_1191_n 5.64871e-19 $X=1.545 $Y=2.285 $X2=0
+ $Y2=0
cc_454 N_B_M1015_g N_A_327_373#_c_1191_n 6.29986e-19 $X=2.695 $Y=2.185 $X2=0
+ $Y2=0
cc_455 N_B_M1022_g N_A_321_77#_c_1283_n 0.017085f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_456 N_B_c_492_n N_A_321_77#_c_1283_n 0.00418899f $X=4.105 $Y=1.515 $X2=0
+ $Y2=0
cc_457 N_B_c_493_n N_A_321_77#_c_1283_n 0.00411871f $X=4.14 $Y=1.515 $X2=0 $Y2=0
cc_458 N_B_c_500_n N_A_321_77#_c_1310_n 0.00110103f $X=3.81 $Y=3.075 $X2=0 $Y2=0
cc_459 N_B_c_499_n N_A_321_77#_c_1289_n 9.70855e-19 $X=3.735 $Y=3.15 $X2=0 $Y2=0
cc_460 N_B_c_500_n N_A_321_77#_c_1289_n 0.0129906f $X=3.81 $Y=3.075 $X2=0 $Y2=0
cc_461 N_B_M1007_g N_A_321_77#_c_1289_n 0.0159308f $X=4.33 $Y=2.4 $X2=0 $Y2=0
cc_462 N_B_M1015_g N_A_321_77#_c_1300_n 7.80042e-19 $X=2.695 $Y=2.185 $X2=0
+ $Y2=0
cc_463 N_B_M1022_g N_A_321_77#_c_1284_n 0.00689761f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_464 N_B_c_492_n N_A_321_77#_c_1284_n 0.0322749f $X=4.105 $Y=1.515 $X2=0 $Y2=0
cc_465 N_B_c_493_n N_A_321_77#_c_1284_n 0.0185639f $X=4.14 $Y=1.515 $X2=0 $Y2=0
cc_466 N_B_M1005_g N_A_321_77#_c_1285_n 8.232e-19 $X=2.62 $Y=0.925 $X2=0 $Y2=0
cc_467 N_B_M1005_g N_A_321_77#_c_1286_n 0.00343798f $X=2.62 $Y=0.925 $X2=0 $Y2=0
cc_468 N_B_M1005_g N_A_321_77#_c_1287_n 0.00788426f $X=2.62 $Y=0.925 $X2=0 $Y2=0
cc_469 N_B_M1022_g N_A_321_77#_c_1288_n 0.0123212f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_470 N_B_M1022_g N_VGND_c_1472_n 0.00546687f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_471 N_B_M1024_g N_VGND_c_1479_n 0.00388395f $X=1.53 $Y=0.705 $X2=0 $Y2=0
cc_472 N_B_M1022_g N_VGND_c_1479_n 0.00399972f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_473 N_B_M1024_g N_VGND_c_1484_n 0.0054106f $X=1.53 $Y=0.705 $X2=0 $Y2=0
cc_474 N_B_M1022_g N_VGND_c_1484_n 0.0052212f $X=4.14 $Y=0.815 $X2=0 $Y2=0
cc_475 N_A_1024_300#_M1027_g N_C_M1010_g 0.025185f $X=5.21 $Y=0.69 $X2=0 $Y2=0
cc_476 N_A_1024_300#_c_622_n N_C_M1010_g 6.18081e-19 $X=6.5 $Y=1.55 $X2=0 $Y2=0
cc_477 N_A_1024_300#_c_625_n N_C_M1010_g 6.75097e-19 $X=6.555 $Y=1.085 $X2=0
+ $Y2=0
cc_478 N_A_1024_300#_M1021_g N_C_M1019_g 0.0294248f $X=5.34 $Y=2.41 $X2=0 $Y2=0
cc_479 N_A_1024_300#_c_621_n N_C_M1019_g 0.0161722f $X=6.39 $Y=1.635 $X2=0 $Y2=0
cc_480 N_A_1024_300#_c_622_n N_C_M1019_g 0.00100646f $X=6.5 $Y=1.55 $X2=0 $Y2=0
cc_481 N_A_1024_300#_c_629_n N_C_M1019_g 0.0069934f $X=6.525 $Y=1.99 $X2=0 $Y2=0
cc_482 N_A_1024_300#_c_623_n N_C_M1019_g 0.00967896f $X=5.285 $Y=1.665 $X2=0
+ $Y2=0
cc_483 N_A_1024_300#_c_624_n N_C_M1019_g 3.42292e-19 $X=5.45 $Y=1.665 $X2=0
+ $Y2=0
cc_484 N_A_1024_300#_c_633_n N_C_M1019_g 0.00107461f $X=6.795 $Y=2.235 $X2=0
+ $Y2=0
cc_485 N_A_1024_300#_c_621_n N_C_c_708_n 0.00546398f $X=6.39 $Y=1.635 $X2=0
+ $Y2=0
cc_486 N_A_1024_300#_c_622_n N_C_c_709_n 0.00567584f $X=6.5 $Y=1.55 $X2=0 $Y2=0
cc_487 N_A_1024_300#_c_625_n N_C_c_709_n 0.00308441f $X=6.555 $Y=1.085 $X2=0
+ $Y2=0
cc_488 N_A_1024_300#_c_629_n N_C_M1012_g 0.0061466f $X=6.525 $Y=1.99 $X2=0 $Y2=0
cc_489 N_A_1024_300#_c_626_n N_C_M1012_g 2.19982e-19 $X=6.5 $Y=1.635 $X2=0 $Y2=0
cc_490 N_A_1024_300#_c_633_n N_C_M1012_g 0.00953209f $X=6.795 $Y=2.235 $X2=0
+ $Y2=0
cc_491 N_A_1024_300#_c_621_n N_C_c_710_n 0.0113645f $X=6.39 $Y=1.635 $X2=0 $Y2=0
cc_492 N_A_1024_300#_c_622_n N_C_c_710_n 0.0202007f $X=6.5 $Y=1.55 $X2=0 $Y2=0
cc_493 N_A_1024_300#_c_633_n N_C_c_710_n 0.00325694f $X=6.795 $Y=2.235 $X2=0
+ $Y2=0
cc_494 N_A_1024_300#_c_622_n N_C_c_711_n 0.0147109f $X=6.5 $Y=1.55 $X2=0 $Y2=0
cc_495 N_A_1024_300#_c_629_n N_C_c_711_n 0.0047192f $X=6.525 $Y=1.99 $X2=0 $Y2=0
cc_496 N_A_1024_300#_c_626_n N_C_c_711_n 0.0145003f $X=6.5 $Y=1.635 $X2=0 $Y2=0
cc_497 N_A_1024_300#_c_633_n N_C_c_711_n 0.0109838f $X=6.795 $Y=2.235 $X2=0
+ $Y2=0
cc_498 N_A_1024_300#_c_622_n N_C_c_712_n 6.32325e-19 $X=6.5 $Y=1.55 $X2=0 $Y2=0
cc_499 N_A_1024_300#_c_626_n N_C_c_712_n 0.00176488f $X=6.5 $Y=1.635 $X2=0 $Y2=0
cc_500 N_A_1024_300#_c_633_n N_C_c_712_n 0.00417286f $X=6.795 $Y=2.235 $X2=0
+ $Y2=0
cc_501 N_A_1024_300#_M1027_g N_A_1057_74#_c_789_n 0.00371279f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_502 N_A_1024_300#_c_633_n N_A_1057_74#_c_801_n 0.0197165f $X=6.795 $Y=2.235
+ $X2=0 $Y2=0
cc_503 N_A_1024_300#_M1017_s N_A_1057_74#_c_791_n 0.00131178f $X=6.41 $Y=0.81
+ $X2=0 $Y2=0
cc_504 N_A_1024_300#_c_625_n N_A_1057_74#_c_791_n 0.0125593f $X=6.555 $Y=1.085
+ $X2=0 $Y2=0
cc_505 N_A_1024_300#_M1017_s N_A_1057_74#_c_792_n 9.85725e-19 $X=6.41 $Y=0.81
+ $X2=0 $Y2=0
cc_506 N_A_1024_300#_c_625_n N_A_1057_74#_c_792_n 0.00979215f $X=6.555 $Y=1.085
+ $X2=0 $Y2=0
cc_507 N_A_1024_300#_c_633_n N_A_1057_74#_c_802_n 0.0160153f $X=6.795 $Y=2.235
+ $X2=0 $Y2=0
cc_508 N_A_1024_300#_M1021_g N_A_1057_74#_c_804_n 0.00443659f $X=5.34 $Y=2.41
+ $X2=0 $Y2=0
cc_509 N_A_1024_300#_M1021_g N_VPWR_c_1050_n 0.0059693f $X=5.34 $Y=2.41 $X2=0
+ $Y2=0
cc_510 N_A_1024_300#_M1021_g N_VPWR_c_1059_n 0.00585197f $X=5.34 $Y=2.41 $X2=0
+ $Y2=0
cc_511 N_A_1024_300#_M1021_g N_VPWR_c_1048_n 0.00606454f $X=5.34 $Y=2.41 $X2=0
+ $Y2=0
cc_512 N_A_1024_300#_M1027_g N_A_327_373#_c_1158_n 0.00287206f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_513 N_A_1024_300#_M1021_g N_A_327_373#_c_1158_n 0.00350805f $X=5.34 $Y=2.41
+ $X2=0 $Y2=0
cc_514 N_A_1024_300#_c_623_n N_A_327_373#_c_1158_n 0.00360941f $X=5.285 $Y=1.665
+ $X2=0 $Y2=0
cc_515 N_A_1024_300#_c_624_n N_A_327_373#_c_1158_n 0.0179619f $X=5.45 $Y=1.665
+ $X2=0 $Y2=0
cc_516 N_A_1024_300#_M1027_g N_A_327_373#_c_1160_n 8.88219e-19 $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_517 N_A_1024_300#_c_621_n N_A_327_373#_c_1160_n 0.0375039f $X=6.39 $Y=1.635
+ $X2=0 $Y2=0
cc_518 N_A_1024_300#_c_622_n N_A_327_373#_c_1160_n 0.0135138f $X=6.5 $Y=1.55
+ $X2=0 $Y2=0
cc_519 N_A_1024_300#_M1027_g N_A_327_373#_c_1161_n 8.1639e-19 $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_520 N_A_1024_300#_c_625_n N_A_327_373#_c_1161_n 0.0120836f $X=6.555 $Y=1.085
+ $X2=0 $Y2=0
cc_521 N_A_1024_300#_M1027_g N_A_327_373#_c_1162_n 0.0163205f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_522 N_A_1024_300#_c_623_n N_A_327_373#_c_1162_n 0.00488549f $X=5.285 $Y=1.665
+ $X2=0 $Y2=0
cc_523 N_A_1024_300#_c_624_n N_A_327_373#_c_1162_n 0.0375039f $X=5.45 $Y=1.665
+ $X2=0 $Y2=0
cc_524 N_A_1024_300#_M1021_g N_A_327_373#_c_1167_n 8.06492e-19 $X=5.34 $Y=2.41
+ $X2=0 $Y2=0
cc_525 N_A_1024_300#_c_623_n N_A_327_373#_c_1167_n 0.00195829f $X=5.285 $Y=1.665
+ $X2=0 $Y2=0
cc_526 N_A_1024_300#_c_624_n N_A_327_373#_c_1167_n 0.00182723f $X=5.45 $Y=1.665
+ $X2=0 $Y2=0
cc_527 N_A_1024_300#_M1021_g N_A_327_373#_c_1168_n 0.00775196f $X=5.34 $Y=2.41
+ $X2=0 $Y2=0
cc_528 N_A_1024_300#_c_623_n N_A_327_373#_c_1168_n 0.00356588f $X=5.285 $Y=1.665
+ $X2=0 $Y2=0
cc_529 N_A_1024_300#_c_624_n N_A_327_373#_c_1168_n 0.0112608f $X=5.45 $Y=1.665
+ $X2=0 $Y2=0
cc_530 N_A_1024_300#_M1027_g N_A_321_77#_c_1284_n 0.00491664f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_531 N_A_1024_300#_M1021_g N_A_321_77#_c_1284_n 0.00243364f $X=5.34 $Y=2.41
+ $X2=0 $Y2=0
cc_532 N_A_1024_300#_M1021_g N_A_321_77#_c_1291_n 0.0187297f $X=5.34 $Y=2.41
+ $X2=0 $Y2=0
cc_533 N_A_1024_300#_c_621_n N_A_321_77#_c_1291_n 0.0134861f $X=6.39 $Y=1.635
+ $X2=0 $Y2=0
cc_534 N_A_1024_300#_c_624_n N_A_321_77#_c_1291_n 0.00385886f $X=5.45 $Y=1.665
+ $X2=0 $Y2=0
cc_535 N_A_1024_300#_c_633_n N_A_321_77#_c_1291_n 0.00981818f $X=6.795 $Y=2.235
+ $X2=0 $Y2=0
cc_536 N_A_1024_300#_M1021_g N_A_321_77#_c_1292_n 0.00186716f $X=5.34 $Y=2.41
+ $X2=0 $Y2=0
cc_537 N_A_1024_300#_c_621_n N_A_321_77#_c_1292_n 0.0157392f $X=6.39 $Y=1.635
+ $X2=0 $Y2=0
cc_538 N_A_1024_300#_c_629_n N_A_321_77#_c_1292_n 0.00155138f $X=6.525 $Y=1.99
+ $X2=0 $Y2=0
cc_539 N_A_1024_300#_c_633_n N_A_321_77#_c_1292_n 0.0332585f $X=6.795 $Y=2.235
+ $X2=0 $Y2=0
cc_540 N_A_1024_300#_M1027_g N_A_321_77#_c_1288_n 0.00867986f $X=5.21 $Y=0.69
+ $X2=0 $Y2=0
cc_541 N_A_1024_300#_M1021_g N_A_321_77#_c_1357_n 5.14561e-19 $X=5.34 $Y=2.41
+ $X2=0 $Y2=0
cc_542 N_A_1024_300#_M1027_g N_VGND_c_1472_n 0.00294228f $X=5.21 $Y=0.69 $X2=0
+ $Y2=0
cc_543 N_A_1024_300#_M1027_g N_VGND_c_1473_n 0.00433139f $X=5.21 $Y=0.69 $X2=0
+ $Y2=0
cc_544 N_A_1024_300#_M1027_g N_VGND_c_1484_n 0.00823742f $X=5.21 $Y=0.69 $X2=0
+ $Y2=0
cc_545 N_C_M1010_g N_A_1057_74#_c_788_n 0.014965f $X=5.765 $Y=0.69 $X2=0 $Y2=0
cc_546 N_C_M1019_g N_A_1057_74#_c_801_n 0.00906351f $X=5.96 $Y=2.41 $X2=0 $Y2=0
cc_547 N_C_M1012_g N_A_1057_74#_c_801_n 0.00619452f $X=7.02 $Y=2.16 $X2=0 $Y2=0
cc_548 N_C_M1010_g N_A_1057_74#_c_790_n 0.00287215f $X=5.765 $Y=0.69 $X2=0 $Y2=0
cc_549 N_C_c_709_n N_A_1057_74#_c_791_n 0.0148447f $X=6.77 $Y=1.35 $X2=0 $Y2=0
cc_550 N_C_c_710_n N_A_1057_74#_c_791_n 3.54962e-19 $X=6.695 $Y=1.515 $X2=0
+ $Y2=0
cc_551 N_C_c_711_n N_A_1057_74#_c_791_n 0.00258247f $X=6.945 $Y=1.515 $X2=0
+ $Y2=0
cc_552 N_C_c_710_n N_A_1057_74#_c_792_n 0.00209722f $X=6.695 $Y=1.515 $X2=0
+ $Y2=0
cc_553 N_C_c_711_n N_A_1057_74#_c_822_n 0.00367584f $X=6.945 $Y=1.515 $X2=0
+ $Y2=0
cc_554 N_C_c_712_n N_A_1057_74#_c_822_n 3.38629e-19 $X=7.02 $Y=1.515 $X2=0 $Y2=0
cc_555 N_C_c_711_n N_A_1057_74#_c_824_n 0.0135553f $X=6.945 $Y=1.515 $X2=0 $Y2=0
cc_556 N_C_c_712_n N_A_1057_74#_c_824_n 0.0012626f $X=7.02 $Y=1.515 $X2=0 $Y2=0
cc_557 N_C_M1012_g N_A_1057_74#_c_802_n 0.012537f $X=7.02 $Y=2.16 $X2=0 $Y2=0
cc_558 N_C_c_709_n N_A_1057_74#_c_793_n 0.00395023f $X=6.77 $Y=1.35 $X2=0 $Y2=0
cc_559 N_C_c_711_n N_A_1057_74#_c_803_n 0.00699102f $X=6.945 $Y=1.515 $X2=0
+ $Y2=0
cc_560 N_C_c_712_n N_A_1057_74#_c_803_n 0.00783455f $X=7.02 $Y=1.515 $X2=0 $Y2=0
cc_561 N_C_M1019_g N_A_1057_74#_c_804_n 0.00300819f $X=5.96 $Y=2.41 $X2=0 $Y2=0
cc_562 N_C_c_711_n N_A_1057_74#_c_794_n 0.0215512f $X=6.945 $Y=1.515 $X2=0 $Y2=0
cc_563 N_C_c_712_n N_A_1057_74#_c_794_n 0.00122161f $X=7.02 $Y=1.515 $X2=0 $Y2=0
cc_564 N_C_c_711_n N_A_1057_74#_c_795_n 4.00288e-19 $X=6.945 $Y=1.515 $X2=0
+ $Y2=0
cc_565 N_C_c_712_n N_A_1057_74#_c_795_n 0.0209673f $X=7.02 $Y=1.515 $X2=0 $Y2=0
cc_566 N_C_M1012_g N_VPWR_c_1052_n 9.08989e-19 $X=7.02 $Y=2.16 $X2=0 $Y2=0
cc_567 N_C_M1019_g N_VPWR_c_1059_n 8.50192e-19 $X=5.96 $Y=2.41 $X2=0 $Y2=0
cc_568 N_C_M1010_g N_A_327_373#_c_1160_n 0.0147025f $X=5.765 $Y=0.69 $X2=0 $Y2=0
cc_569 N_C_c_708_n N_A_327_373#_c_1160_n 0.00755929f $X=6.05 $Y=1.425 $X2=0
+ $Y2=0
cc_570 N_C_c_710_n N_A_327_373#_c_1160_n 0.00362102f $X=6.695 $Y=1.515 $X2=0
+ $Y2=0
cc_571 N_C_M1010_g N_A_327_373#_c_1161_n 0.0112653f $X=5.765 $Y=0.69 $X2=0 $Y2=0
cc_572 N_C_c_708_n N_A_327_373#_c_1161_n 0.00111695f $X=6.05 $Y=1.425 $X2=0
+ $Y2=0
cc_573 N_C_c_709_n N_A_327_373#_c_1161_n 0.0035702f $X=6.77 $Y=1.35 $X2=0 $Y2=0
cc_574 N_C_M1019_g N_A_327_373#_c_1168_n 0.00118539f $X=5.96 $Y=2.41 $X2=0 $Y2=0
cc_575 N_C_M1019_g N_A_321_77#_c_1291_n 0.0169042f $X=5.96 $Y=2.41 $X2=0 $Y2=0
cc_576 N_C_M1012_g N_A_321_77#_c_1291_n 0.0029046f $X=7.02 $Y=2.16 $X2=0 $Y2=0
cc_577 N_C_M1019_g N_A_321_77#_c_1292_n 0.0105431f $X=5.96 $Y=2.41 $X2=0 $Y2=0
cc_578 N_C_M1012_g N_A_321_77#_c_1292_n 5.24833e-19 $X=7.02 $Y=2.16 $X2=0 $Y2=0
cc_579 N_C_M1010_g N_A_321_77#_c_1288_n 2.05732e-19 $X=5.765 $Y=0.69 $X2=0 $Y2=0
cc_580 N_C_M1010_g N_VGND_c_1473_n 0.00278271f $X=5.765 $Y=0.69 $X2=0 $Y2=0
cc_581 N_C_c_709_n N_VGND_c_1473_n 5.51389e-19 $X=6.77 $Y=1.35 $X2=0 $Y2=0
cc_582 N_C_c_709_n N_VGND_c_1475_n 7.66361e-19 $X=6.77 $Y=1.35 $X2=0 $Y2=0
cc_583 N_C_M1010_g N_VGND_c_1484_n 0.00359569f $X=5.765 $Y=0.69 $X2=0 $Y2=0
cc_584 N_A_1057_74#_c_802_n N_VPWR_M1012_d 0.0080194f $X=7.222 $Y=2.905 $X2=0
+ $Y2=0
cc_585 N_A_1057_74#_c_803_n N_VPWR_M1012_d 0.00388318f $X=7.405 $Y=1.95 $X2=0
+ $Y2=0
cc_586 N_A_1057_74#_c_837_p N_VPWR_M1012_d 0.0181363f $X=7.405 $Y=2.035 $X2=0
+ $Y2=0
cc_587 N_A_1057_74#_M1002_g N_VPWR_c_1051_n 0.0138522f $X=8.22 $Y=2.4 $X2=0
+ $Y2=0
cc_588 N_A_1057_74#_c_801_n N_VPWR_c_1051_n 0.0156625f $X=7.13 $Y=2.99 $X2=0
+ $Y2=0
cc_589 N_A_1057_74#_c_802_n N_VPWR_c_1052_n 0.00750252f $X=7.222 $Y=2.905 $X2=0
+ $Y2=0
cc_590 N_A_1057_74#_c_803_n N_VPWR_c_1052_n 0.00774637f $X=7.405 $Y=1.95 $X2=0
+ $Y2=0
cc_591 N_A_1057_74#_c_842_p N_VPWR_c_1052_n 0.0333159f $X=8.165 $Y=1.505 $X2=0
+ $Y2=0
cc_592 N_A_1057_74#_c_837_p N_VPWR_c_1052_n 0.0125379f $X=7.405 $Y=2.035 $X2=0
+ $Y2=0
cc_593 N_A_1057_74#_c_795_n N_VPWR_c_1052_n 0.00974437f $X=8.13 $Y=1.505 $X2=0
+ $Y2=0
cc_594 N_A_1057_74#_M1002_g N_VPWR_c_1053_n 0.005209f $X=8.22 $Y=2.4 $X2=0 $Y2=0
cc_595 N_A_1057_74#_M1008_g N_VPWR_c_1053_n 0.0048691f $X=8.67 $Y=2.4 $X2=0
+ $Y2=0
cc_596 N_A_1057_74#_M1008_g N_VPWR_c_1054_n 0.00312167f $X=8.67 $Y=2.4 $X2=0
+ $Y2=0
cc_597 N_A_1057_74#_M1023_g N_VPWR_c_1054_n 0.00313866f $X=9.12 $Y=2.4 $X2=0
+ $Y2=0
cc_598 N_A_1057_74#_c_785_n N_VPWR_c_1054_n 0.00234748f $X=9.57 $Y=1.665 $X2=0
+ $Y2=0
cc_599 N_A_1057_74#_M1026_g N_VPWR_c_1056_n 0.0064767f $X=9.57 $Y=2.4 $X2=0
+ $Y2=0
cc_600 N_A_1057_74#_c_802_n N_VPWR_c_1118_n 0.0502413f $X=7.222 $Y=2.905 $X2=0
+ $Y2=0
cc_601 N_A_1057_74#_c_842_p N_VPWR_c_1118_n 0.00580119f $X=8.165 $Y=1.505 $X2=0
+ $Y2=0
cc_602 N_A_1057_74#_c_795_n N_VPWR_c_1118_n 0.00332899f $X=8.13 $Y=1.505 $X2=0
+ $Y2=0
cc_603 N_A_1057_74#_c_801_n N_VPWR_c_1059_n 0.097943f $X=7.13 $Y=2.99 $X2=0
+ $Y2=0
cc_604 N_A_1057_74#_c_804_n N_VPWR_c_1059_n 0.0223614f $X=5.65 $Y=2.895 $X2=0
+ $Y2=0
cc_605 N_A_1057_74#_M1023_g N_VPWR_c_1060_n 0.005209f $X=9.12 $Y=2.4 $X2=0 $Y2=0
cc_606 N_A_1057_74#_M1026_g N_VPWR_c_1060_n 0.00492575f $X=9.57 $Y=2.4 $X2=0
+ $Y2=0
cc_607 N_A_1057_74#_M1002_g N_VPWR_c_1048_n 0.00986727f $X=8.22 $Y=2.4 $X2=0
+ $Y2=0
cc_608 N_A_1057_74#_M1008_g N_VPWR_c_1048_n 0.00872205f $X=8.67 $Y=2.4 $X2=0
+ $Y2=0
cc_609 N_A_1057_74#_M1023_g N_VPWR_c_1048_n 0.00982266f $X=9.12 $Y=2.4 $X2=0
+ $Y2=0
cc_610 N_A_1057_74#_M1026_g N_VPWR_c_1048_n 0.00894308f $X=9.57 $Y=2.4 $X2=0
+ $Y2=0
cc_611 N_A_1057_74#_c_801_n N_VPWR_c_1048_n 0.0566295f $X=7.13 $Y=2.99 $X2=0
+ $Y2=0
cc_612 N_A_1057_74#_c_804_n N_VPWR_c_1048_n 0.0125377f $X=5.65 $Y=2.895 $X2=0
+ $Y2=0
cc_613 N_A_1057_74#_c_788_n N_A_327_373#_M1010_d 0.00294181f $X=6.33 $Y=0.34
+ $X2=0 $Y2=0
cc_614 N_A_1057_74#_c_787_n N_A_327_373#_c_1160_n 0.0200764f $X=5.495 $Y=0.515
+ $X2=0 $Y2=0
cc_615 N_A_1057_74#_c_788_n N_A_327_373#_c_1161_n 0.0204002f $X=6.33 $Y=0.34
+ $X2=0 $Y2=0
cc_616 N_A_1057_74#_c_790_n N_A_327_373#_c_1161_n 0.00511586f $X=6.415 $Y=0.66
+ $X2=0 $Y2=0
cc_617 N_A_1057_74#_c_792_n N_A_327_373#_c_1161_n 0.0150383f $X=6.5 $Y=0.745
+ $X2=0 $Y2=0
cc_618 N_A_1057_74#_c_787_n N_A_327_373#_c_1162_n 0.00496574f $X=5.495 $Y=0.515
+ $X2=0 $Y2=0
cc_619 N_A_1057_74#_M1021_d N_A_321_77#_c_1291_n 0.0110211f $X=5.43 $Y=1.99
+ $X2=0 $Y2=0
cc_620 N_A_1057_74#_c_801_n N_A_321_77#_c_1291_n 0.0231171f $X=7.13 $Y=2.99
+ $X2=0 $Y2=0
cc_621 N_A_1057_74#_c_804_n N_A_321_77#_c_1291_n 0.0243659f $X=5.65 $Y=2.895
+ $X2=0 $Y2=0
cc_622 N_A_1057_74#_c_789_n N_A_321_77#_c_1288_n 0.00373319f $X=5.66 $Y=0.34
+ $X2=0 $Y2=0
cc_623 N_A_1057_74#_M1002_g N_X_c_1416_n 0.0121191f $X=8.22 $Y=2.4 $X2=0 $Y2=0
cc_624 N_A_1057_74#_M1008_g N_X_c_1416_n 0.0138639f $X=8.67 $Y=2.4 $X2=0 $Y2=0
cc_625 N_A_1057_74#_c_782_n N_X_c_1413_n 0.0063516f $X=8.295 $Y=1.34 $X2=0 $Y2=0
cc_626 N_A_1057_74#_c_783_n N_X_c_1413_n 0.00605329f $X=8.725 $Y=1.34 $X2=0
+ $Y2=0
cc_627 N_A_1057_74#_c_784_n N_X_c_1413_n 4.95297e-19 $X=9.155 $Y=1.34 $X2=0
+ $Y2=0
cc_628 N_A_1057_74#_c_782_n N_X_c_1414_n 0.00383504f $X=8.295 $Y=1.34 $X2=0
+ $Y2=0
cc_629 N_A_1057_74#_c_783_n N_X_c_1414_n 0.00350884f $X=8.725 $Y=1.34 $X2=0
+ $Y2=0
cc_630 N_A_1057_74#_c_785_n N_X_c_1414_n 0.00677107f $X=9.57 $Y=1.665 $X2=0
+ $Y2=0
cc_631 N_A_1057_74#_c_842_p N_X_c_1414_n 0.00606139f $X=8.165 $Y=1.505 $X2=0
+ $Y2=0
cc_632 N_A_1057_74#_c_785_n N_X_c_1429_n 0.0433288f $X=9.57 $Y=1.665 $X2=0 $Y2=0
cc_633 N_A_1057_74#_M1002_g N_X_c_1417_n 0.00285641f $X=8.22 $Y=2.4 $X2=0 $Y2=0
cc_634 N_A_1057_74#_M1008_g N_X_c_1417_n 0.00238576f $X=8.67 $Y=2.4 $X2=0 $Y2=0
cc_635 N_A_1057_74#_c_785_n N_X_c_1417_n 0.0023482f $X=9.57 $Y=1.665 $X2=0 $Y2=0
cc_636 N_A_1057_74#_c_842_p N_X_c_1417_n 0.00151667f $X=8.165 $Y=1.505 $X2=0
+ $Y2=0
cc_637 N_A_1057_74#_M1002_g N_X_c_1418_n 0.00353963f $X=8.22 $Y=2.4 $X2=0 $Y2=0
cc_638 N_A_1057_74#_M1008_g N_X_c_1418_n 0.00438312f $X=8.67 $Y=2.4 $X2=0 $Y2=0
cc_639 N_A_1057_74#_M1023_g N_X_c_1418_n 7.99417e-19 $X=9.12 $Y=2.4 $X2=0 $Y2=0
cc_640 N_A_1057_74#_c_785_n N_X_c_1418_n 0.00285477f $X=9.57 $Y=1.665 $X2=0
+ $Y2=0
cc_641 N_A_1057_74#_c_842_p N_X_c_1418_n 0.00331766f $X=8.165 $Y=1.505 $X2=0
+ $Y2=0
cc_642 N_A_1057_74#_c_782_n N_X_c_1439_n 0.00245314f $X=8.295 $Y=1.34 $X2=0
+ $Y2=0
cc_643 N_A_1057_74#_c_783_n N_X_c_1439_n 0.0017052f $X=8.725 $Y=1.34 $X2=0 $Y2=0
cc_644 N_A_1057_74#_c_785_n N_X_c_1439_n 3.01015e-19 $X=9.57 $Y=1.665 $X2=0
+ $Y2=0
cc_645 N_A_1057_74#_c_785_n N_X_c_1442_n 0.00868505f $X=9.57 $Y=1.665 $X2=0
+ $Y2=0
cc_646 N_A_1057_74#_c_842_p N_X_c_1442_n 0.0173534f $X=8.165 $Y=1.505 $X2=0
+ $Y2=0
cc_647 N_A_1057_74#_c_783_n X 5.03719e-19 $X=8.725 $Y=1.34 $X2=0 $Y2=0
cc_648 N_A_1057_74#_c_784_n X 0.0128066f $X=9.155 $Y=1.34 $X2=0 $Y2=0
cc_649 N_A_1057_74#_c_785_n X 0.0101295f $X=9.57 $Y=1.665 $X2=0 $Y2=0
cc_650 N_A_1057_74#_c_786_n X 0.015578f $X=9.585 $Y=1.34 $X2=0 $Y2=0
cc_651 N_A_1057_74#_c_785_n X 0.0173378f $X=9.57 $Y=1.665 $X2=0 $Y2=0
cc_652 N_A_1057_74#_M1008_g X 7.96096e-19 $X=8.67 $Y=2.4 $X2=0 $Y2=0
cc_653 N_A_1057_74#_M1023_g X 0.0196086f $X=9.12 $Y=2.4 $X2=0 $Y2=0
cc_654 N_A_1057_74#_c_785_n X 0.00631655f $X=9.57 $Y=1.665 $X2=0 $Y2=0
cc_655 N_A_1057_74#_M1026_g X 0.0262568f $X=9.57 $Y=2.4 $X2=0 $Y2=0
cc_656 N_A_1057_74#_c_791_n N_VGND_M1017_d 0.00369417f $X=6.89 $Y=0.745 $X2=0
+ $Y2=0
cc_657 N_A_1057_74#_c_908_p N_VGND_M1017_d 0.00687894f $X=6.975 $Y=1.01 $X2=0
+ $Y2=0
cc_658 N_A_1057_74#_c_822_n N_VGND_M1017_d 0.0211435f $X=7.32 $Y=1.095 $X2=0
+ $Y2=0
cc_659 N_A_1057_74#_c_824_n N_VGND_M1017_d 0.00276146f $X=7.06 $Y=1.095 $X2=0
+ $Y2=0
cc_660 N_A_1057_74#_c_793_n N_VGND_M1017_d 0.00260794f $X=7.405 $Y=1.34 $X2=0
+ $Y2=0
cc_661 N_A_1057_74#_c_788_n N_VGND_c_1473_n 0.0546988f $X=6.33 $Y=0.34 $X2=0
+ $Y2=0
cc_662 N_A_1057_74#_c_789_n N_VGND_c_1473_n 0.0236566f $X=5.66 $Y=0.34 $X2=0
+ $Y2=0
cc_663 N_A_1057_74#_c_791_n N_VGND_c_1473_n 0.00691154f $X=6.89 $Y=0.745 $X2=0
+ $Y2=0
cc_664 N_A_1057_74#_c_822_n N_VGND_c_1523_n 0.00671835f $X=7.32 $Y=1.095 $X2=0
+ $Y2=0
cc_665 N_A_1057_74#_c_842_p N_VGND_c_1523_n 0.0203974f $X=8.165 $Y=1.505 $X2=0
+ $Y2=0
cc_666 N_A_1057_74#_c_795_n N_VGND_c_1523_n 0.00588813f $X=8.13 $Y=1.505 $X2=0
+ $Y2=0
cc_667 N_A_1057_74#_c_782_n N_VGND_c_1474_n 0.00473385f $X=8.295 $Y=1.34 $X2=0
+ $Y2=0
cc_668 N_A_1057_74#_c_783_n N_VGND_c_1474_n 0.00473385f $X=8.725 $Y=1.34 $X2=0
+ $Y2=0
cc_669 N_A_1057_74#_c_782_n N_VGND_c_1475_n 0.00558707f $X=8.295 $Y=1.34 $X2=0
+ $Y2=0
cc_670 N_A_1057_74#_c_788_n N_VGND_c_1475_n 0.00877697f $X=6.33 $Y=0.34 $X2=0
+ $Y2=0
cc_671 N_A_1057_74#_c_790_n N_VGND_c_1475_n 0.00301164f $X=6.415 $Y=0.66 $X2=0
+ $Y2=0
cc_672 N_A_1057_74#_c_791_n N_VGND_c_1475_n 0.028714f $X=6.89 $Y=0.745 $X2=0
+ $Y2=0
cc_673 N_A_1057_74#_c_908_p N_VGND_c_1475_n 7.77107e-19 $X=6.975 $Y=1.01 $X2=0
+ $Y2=0
cc_674 N_A_1057_74#_c_822_n N_VGND_c_1475_n 0.0285331f $X=7.32 $Y=1.095 $X2=0
+ $Y2=0
cc_675 N_A_1057_74#_c_842_p N_VGND_c_1475_n 0.0151658f $X=8.165 $Y=1.505 $X2=0
+ $Y2=0
cc_676 N_A_1057_74#_c_795_n N_VGND_c_1475_n 0.00862364f $X=8.13 $Y=1.505 $X2=0
+ $Y2=0
cc_677 N_A_1057_74#_c_783_n N_VGND_c_1476_n 0.0031573f $X=8.725 $Y=1.34 $X2=0
+ $Y2=0
cc_678 N_A_1057_74#_c_784_n N_VGND_c_1476_n 0.00265542f $X=9.155 $Y=1.34 $X2=0
+ $Y2=0
cc_679 N_A_1057_74#_c_785_n N_VGND_c_1476_n 0.00278273f $X=9.57 $Y=1.665 $X2=0
+ $Y2=0
cc_680 N_A_1057_74#_c_786_n N_VGND_c_1478_n 0.00595876f $X=9.585 $Y=1.34 $X2=0
+ $Y2=0
cc_681 N_A_1057_74#_c_784_n N_VGND_c_1480_n 0.00472938f $X=9.155 $Y=1.34 $X2=0
+ $Y2=0
cc_682 N_A_1057_74#_c_786_n N_VGND_c_1480_n 0.00472938f $X=9.585 $Y=1.34 $X2=0
+ $Y2=0
cc_683 N_A_1057_74#_c_782_n N_VGND_c_1484_n 0.00508379f $X=8.295 $Y=1.34 $X2=0
+ $Y2=0
cc_684 N_A_1057_74#_c_783_n N_VGND_c_1484_n 0.00508379f $X=8.725 $Y=1.34 $X2=0
+ $Y2=0
cc_685 N_A_1057_74#_c_784_n N_VGND_c_1484_n 0.00508379f $X=9.155 $Y=1.34 $X2=0
+ $Y2=0
cc_686 N_A_1057_74#_c_786_n N_VGND_c_1484_n 0.00508379f $X=9.585 $Y=1.34 $X2=0
+ $Y2=0
cc_687 N_A_1057_74#_c_788_n N_VGND_c_1484_n 0.0310803f $X=6.33 $Y=0.34 $X2=0
+ $Y2=0
cc_688 N_A_1057_74#_c_789_n N_VGND_c_1484_n 0.0128296f $X=5.66 $Y=0.34 $X2=0
+ $Y2=0
cc_689 N_A_1057_74#_c_791_n N_VGND_c_1484_n 0.0119702f $X=6.89 $Y=0.745 $X2=0
+ $Y2=0
cc_690 N_A_27_373#_c_971_n N_VPWR_c_1049_n 0.0027218f $X=1.535 $Y=2.035 $X2=0
+ $Y2=0
cc_691 N_A_27_373#_c_953_n N_VPWR_c_1049_n 0.0202902f $X=0.28 $Y=2.01 $X2=0
+ $Y2=0
cc_692 N_A_27_373#_c_953_n N_VPWR_c_1057_n 0.00895579f $X=0.28 $Y=2.01 $X2=0
+ $Y2=0
cc_693 N_A_27_373#_c_953_n N_VPWR_c_1048_n 0.0096603f $X=0.28 $Y=2.01 $X2=0
+ $Y2=0
cc_694 N_A_27_373#_c_947_n N_A_327_373#_M1025_d 0.00382627f $X=2.305 $Y=2.65
+ $X2=0 $Y2=0
cc_695 N_A_27_373#_c_981_n N_A_327_373#_M1025_d 0.00254092f $X=1.68 $Y=2.035
+ $X2=0 $Y2=0
cc_696 N_A_27_373#_c_946_n N_A_327_373#_M1025_d 0.007385f $X=1.68 $Y=2.035 $X2=0
+ $Y2=0
cc_697 N_A_27_373#_c_981_n N_A_327_373#_c_1163_n 3.43164e-19 $X=1.68 $Y=2.035
+ $X2=0 $Y2=0
cc_698 N_A_27_373#_c_946_n N_A_327_373#_c_1163_n 0.022295f $X=1.68 $Y=2.035
+ $X2=0 $Y2=0
cc_699 N_A_27_373#_c_945_n N_A_327_373#_c_1155_n 0.0103721f $X=2.3 $Y=1.1 $X2=0
+ $Y2=0
cc_700 N_A_27_373#_c_951_n N_A_327_373#_c_1155_n 0.00421424f $X=2.47 $Y=2.38
+ $X2=0 $Y2=0
cc_701 N_A_27_373#_c_941_n N_A_327_373#_c_1156_n 0.0158636f $X=2.135 $Y=1.25
+ $X2=0 $Y2=0
cc_702 N_A_27_373#_c_945_n N_A_327_373#_c_1156_n 0.00867013f $X=2.3 $Y=1.1 $X2=0
+ $Y2=0
cc_703 N_A_27_373#_c_946_n N_A_327_373#_c_1156_n 0.0145177f $X=1.68 $Y=2.035
+ $X2=0 $Y2=0
cc_704 N_A_27_373#_c_945_n N_A_327_373#_c_1157_n 0.0096475f $X=2.3 $Y=1.1 $X2=0
+ $Y2=0
cc_705 N_A_27_373#_c_945_n N_A_327_373#_c_1180_n 0.0194434f $X=2.3 $Y=1.1 $X2=0
+ $Y2=0
cc_706 N_A_27_373#_M1014_d N_A_327_373#_c_1166_n 0.00499831f $X=2.335 $Y=1.865
+ $X2=0 $Y2=0
cc_707 N_A_27_373#_c_951_n N_A_327_373#_c_1166_n 0.0127573f $X=2.47 $Y=2.38
+ $X2=0 $Y2=0
cc_708 N_A_27_373#_c_941_n N_A_327_373#_c_1190_n 3.65365e-19 $X=2.135 $Y=1.25
+ $X2=0 $Y2=0
cc_709 N_A_27_373#_c_947_n N_A_327_373#_c_1190_n 0.00479203f $X=2.305 $Y=2.65
+ $X2=0 $Y2=0
cc_710 N_A_27_373#_c_945_n N_A_327_373#_c_1190_n 4.49084e-19 $X=2.3 $Y=1.1 $X2=0
+ $Y2=0
cc_711 N_A_27_373#_c_981_n N_A_327_373#_c_1190_n 0.0210157f $X=1.68 $Y=2.035
+ $X2=0 $Y2=0
cc_712 N_A_27_373#_c_946_n N_A_327_373#_c_1190_n 2.03155e-19 $X=1.68 $Y=2.035
+ $X2=0 $Y2=0
cc_713 N_A_27_373#_c_947_n N_A_327_373#_c_1191_n 0.00904187f $X=2.305 $Y=2.65
+ $X2=0 $Y2=0
cc_714 N_A_27_373#_c_981_n N_A_327_373#_c_1191_n 0.00151832f $X=1.68 $Y=2.035
+ $X2=0 $Y2=0
cc_715 N_A_27_373#_c_946_n N_A_327_373#_c_1191_n 0.0126015f $X=1.68 $Y=2.035
+ $X2=0 $Y2=0
cc_716 N_A_27_373#_c_951_n N_A_321_77#_c_1310_n 0.00615404f $X=2.47 $Y=2.38
+ $X2=0 $Y2=0
cc_717 N_A_27_373#_c_951_n N_A_321_77#_c_1300_n 0.0146685f $X=2.47 $Y=2.38 $X2=0
+ $Y2=0
cc_718 N_A_27_373#_c_941_n N_A_321_77#_c_1285_n 0.0124306f $X=2.135 $Y=1.25
+ $X2=0 $Y2=0
cc_719 N_A_27_373#_c_944_n N_A_321_77#_c_1285_n 0.0108039f $X=1.665 $Y=1.475
+ $X2=0 $Y2=0
cc_720 N_A_27_373#_M1006_d N_A_321_77#_c_1286_n 0.00731496f $X=2.08 $Y=0.605
+ $X2=0 $Y2=0
cc_721 N_A_27_373#_c_941_n N_A_321_77#_c_1286_n 0.00539878f $X=2.135 $Y=1.25
+ $X2=0 $Y2=0
cc_722 N_A_27_373#_c_945_n N_A_321_77#_c_1286_n 0.0192566f $X=2.3 $Y=1.1 $X2=0
+ $Y2=0
cc_723 N_A_27_373#_c_942_n N_VGND_c_1471_n 0.0201853f $X=0.33 $Y=0.615 $X2=0
+ $Y2=0
cc_724 N_A_27_373#_c_942_n N_VGND_c_1481_n 0.016911f $X=0.33 $Y=0.615 $X2=0
+ $Y2=0
cc_725 N_A_27_373#_c_942_n N_VGND_c_1484_n 0.0148316f $X=0.33 $Y=0.615 $X2=0
+ $Y2=0
cc_726 N_VPWR_M1007_d N_A_327_373#_c_1166_n 0.00516574f $X=4.42 $Y=1.84 $X2=0
+ $Y2=0
cc_727 N_VPWR_c_1050_n N_A_321_77#_c_1289_n 0.00191073f $X=4.555 $Y=2.815 $X2=0
+ $Y2=0
cc_728 N_VPWR_c_1048_n N_A_321_77#_c_1289_n 0.0245273f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_729 N_VPWR_M1007_d N_A_321_77#_c_1284_n 0.00819394f $X=4.42 $Y=1.84 $X2=0
+ $Y2=0
cc_730 N_VPWR_M1007_d N_A_321_77#_c_1291_n 0.00305933f $X=4.42 $Y=1.84 $X2=0
+ $Y2=0
cc_731 N_VPWR_c_1050_n N_A_321_77#_c_1291_n 0.0086438f $X=4.555 $Y=2.815 $X2=0
+ $Y2=0
cc_732 N_VPWR_c_1048_n N_A_321_77#_c_1291_n 0.0290398f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_733 N_VPWR_M1007_d N_A_321_77#_c_1357_n 0.00194601f $X=4.42 $Y=1.84 $X2=0
+ $Y2=0
cc_734 N_VPWR_c_1050_n N_A_321_77#_c_1357_n 0.0115793f $X=4.555 $Y=2.815 $X2=0
+ $Y2=0
cc_735 N_VPWR_c_1048_n N_A_321_77#_c_1357_n 6.84279e-19 $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_736 N_VPWR_c_1053_n N_X_c_1416_n 0.0157112f $X=8.81 $Y=3.33 $X2=0 $Y2=0
cc_737 N_VPWR_c_1048_n N_X_c_1416_n 0.0127977f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_738 N_VPWR_c_1054_n N_X_c_1429_n 0.0123826f $X=8.895 $Y=1.985 $X2=0 $Y2=0
cc_739 N_VPWR_c_1051_n N_X_c_1417_n 0.0441815f $X=7.797 $Y=3.245 $X2=0 $Y2=0
cc_740 N_VPWR_c_1054_n N_X_c_1418_n 0.0453846f $X=8.895 $Y=1.985 $X2=0 $Y2=0
cc_741 N_VPWR_c_1054_n X 0.0399213f $X=8.895 $Y=1.985 $X2=0 $Y2=0
cc_742 N_VPWR_c_1056_n X 0.0444885f $X=9.795 $Y=1.985 $X2=0 $Y2=0
cc_743 N_VPWR_c_1060_n X 0.0155031f $X=9.71 $Y=3.33 $X2=0 $Y2=0
cc_744 N_VPWR_c_1048_n X 0.0126371f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_745 N_VPWR_c_1056_n N_VGND_c_1478_n 0.00977564f $X=9.795 $Y=1.985 $X2=0 $Y2=0
cc_746 N_A_327_373#_c_1166_n N_A_321_77#_M1015_d 0.00836769f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_747 N_A_327_373#_M1005_d N_A_321_77#_c_1283_n 0.00368186f $X=2.695 $Y=0.605
+ $X2=0 $Y2=0
cc_748 N_A_327_373#_c_1163_n N_A_321_77#_c_1310_n 0.00170948f $X=2.09 $Y=1.965
+ $X2=0 $Y2=0
cc_749 N_A_327_373#_c_1180_n N_A_321_77#_c_1310_n 0.00214892f $X=2.845 $Y=1.04
+ $X2=0 $Y2=0
cc_750 N_A_327_373#_c_1166_n N_A_321_77#_c_1310_n 0.0281991f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_751 N_A_327_373#_c_1190_n N_A_321_77#_c_1310_n 0.0020436f $X=2.305 $Y=2.035
+ $X2=0 $Y2=0
cc_752 N_A_327_373#_c_1191_n N_A_321_77#_c_1310_n 0.00169502f $X=2.02 $Y=1.99
+ $X2=0 $Y2=0
cc_753 N_A_327_373#_c_1166_n N_A_321_77#_c_1289_n 0.0220158f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_754 N_A_327_373#_c_1158_n N_A_321_77#_c_1284_n 0.0425791f $X=4.865 $Y=1.95
+ $X2=0 $Y2=0
cc_755 N_A_327_373#_c_1159_n N_A_321_77#_c_1284_n 0.014358f $X=4.95 $Y=1.295
+ $X2=0 $Y2=0
cc_756 N_A_327_373#_c_1166_n N_A_321_77#_c_1284_n 0.0225247f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_757 N_A_327_373#_c_1167_n N_A_321_77#_c_1284_n 5.02359e-19 $X=5.04 $Y=2.035
+ $X2=0 $Y2=0
cc_758 N_A_327_373#_c_1168_n N_A_321_77#_c_1284_n 0.0200577f $X=5.04 $Y=2.035
+ $X2=0 $Y2=0
cc_759 N_A_327_373#_M1021_s N_A_321_77#_c_1291_n 0.00728035f $X=4.97 $Y=1.99
+ $X2=0 $Y2=0
cc_760 N_A_327_373#_c_1166_n N_A_321_77#_c_1291_n 0.00753536f $X=4.895 $Y=2.035
+ $X2=0 $Y2=0
cc_761 N_A_327_373#_c_1167_n N_A_321_77#_c_1291_n 0.00183698f $X=5.04 $Y=2.035
+ $X2=0 $Y2=0
cc_762 N_A_327_373#_c_1168_n N_A_321_77#_c_1291_n 0.031299f $X=5.04 $Y=2.035
+ $X2=0 $Y2=0
cc_763 N_A_327_373#_c_1180_n N_A_321_77#_c_1287_n 0.0254466f $X=2.845 $Y=1.04
+ $X2=0 $Y2=0
cc_764 N_A_327_373#_c_1159_n N_A_321_77#_c_1288_n 0.015131f $X=4.95 $Y=1.295
+ $X2=0 $Y2=0
cc_765 N_A_327_373#_c_1161_n N_A_321_77#_c_1288_n 5.07708e-19 $X=5.995 $Y=0.81
+ $X2=0 $Y2=0
cc_766 N_A_327_373#_c_1162_n N_A_321_77#_c_1288_n 0.0167867f $X=5.405 $Y=1.28
+ $X2=0 $Y2=0
cc_767 N_A_321_77#_c_1283_n N_VGND_M1022_d 0.00524428f $X=4.44 $Y=0.7 $X2=0
+ $Y2=0
cc_768 N_A_321_77#_c_1284_n N_VGND_M1022_d 0.00315635f $X=4.525 $Y=2.37 $X2=0
+ $Y2=0
cc_769 N_A_321_77#_c_1288_n N_VGND_M1022_d 0.00804534f $X=4.525 $Y=0.69 $X2=0
+ $Y2=0
cc_770 N_A_321_77#_c_1283_n N_VGND_c_1472_n 0.0127357f $X=4.44 $Y=0.7 $X2=0
+ $Y2=0
cc_771 N_A_321_77#_c_1288_n N_VGND_c_1472_n 0.0197889f $X=4.525 $Y=0.69 $X2=0
+ $Y2=0
cc_772 N_A_321_77#_c_1288_n N_VGND_c_1473_n 0.019328f $X=4.525 $Y=0.69 $X2=0
+ $Y2=0
cc_773 N_A_321_77#_c_1283_n N_VGND_c_1479_n 0.0126356f $X=4.44 $Y=0.7 $X2=0
+ $Y2=0
cc_774 N_A_321_77#_c_1283_n N_VGND_c_1484_n 0.0238176f $X=4.44 $Y=0.7 $X2=0
+ $Y2=0
cc_775 N_A_321_77#_c_1288_n N_VGND_c_1484_n 0.0198891f $X=4.525 $Y=0.69 $X2=0
+ $Y2=0
cc_776 N_X_c_1413_n N_VGND_c_1474_n 0.00971834f $X=8.51 $Y=0.635 $X2=0 $Y2=0
cc_777 N_X_c_1413_n N_VGND_c_1475_n 0.0141711f $X=8.51 $Y=0.635 $X2=0 $Y2=0
cc_778 N_X_c_1413_n N_VGND_c_1476_n 0.0290583f $X=8.51 $Y=0.635 $X2=0 $Y2=0
cc_779 N_X_c_1429_n N_VGND_c_1476_n 0.0137224f $X=9.18 $Y=1.522 $X2=0 $Y2=0
cc_780 X N_VGND_c_1476_n 0.0314886f $X=9.275 $Y=0.47 $X2=0 $Y2=0
cc_781 X N_VGND_c_1478_n 0.0316368f $X=9.275 $Y=0.47 $X2=0 $Y2=0
cc_782 X N_VGND_c_1480_n 0.0105983f $X=9.275 $Y=0.47 $X2=0 $Y2=0
cc_783 N_X_c_1413_n N_VGND_c_1484_n 0.0111609f $X=8.51 $Y=0.635 $X2=0 $Y2=0
cc_784 X N_VGND_c_1484_n 0.0113894f $X=9.275 $Y=0.47 $X2=0 $Y2=0

* NGSPICE file created from sky130_fd_sc_ms__nand3_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__nand3_1 A B C VGND VNB VPB VPWR Y
M1000 Y A a_233_74# VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=3.108e+11p ps=2.32e+06u
M1001 a_233_74# B a_155_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1002 a_155_74# C VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1003 Y C VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.16e+11p pd=5.58e+06u as=8.4e+11p ps=5.98e+06u
M1004 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR B Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__dlygate4sd2_1.pex.spice
* Created: Wed Sep  2 12:06:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%A 3 7 9 10 14
c33 9 0 1.89038e-19 $X=0.24 $Y=1.295
r34 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.57 $Y=1.355
+ $X2=0.57 $Y2=1.52
r35 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.57 $Y=1.355
+ $X2=0.57 $Y2=1.19
r36 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.57
+ $Y=1.355 $X2=0.57 $Y2=1.355
r37 10 15 5.88547 $w=6.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.415 $Y=1.665
+ $X2=0.415 $Y2=1.355
r38 9 15 1.13912 $w=6.28e-07 $l=6e-08 $layer=LI1_cond $X=0.415 $Y=1.295
+ $X2=0.415 $Y2=1.355
r39 7 17 398.427 $w=1.8e-07 $l=1.025e-06 $layer=POLY_cond $X=0.495 $Y=2.545
+ $X2=0.495 $Y2=1.52
r40 3 16 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.48 $Y=0.58 $X2=0.48
+ $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%A_28_74# 1 2 9 13 17 21 23 24 25 26 30
+ 31
c60 9 0 1.89038e-19 $X=1.32 $Y=2.46
r61 31 34 67.4048 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.195 $Y=1.295
+ $X2=1.195 $Y2=1.8
r62 31 33 40.7881 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.195 $Y=1.295
+ $X2=1.195 $Y2=1.13
r63 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.14
+ $Y=1.295 $X2=1.14 $Y2=1.295
r64 28 30 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=1.14 $Y=2.03
+ $X2=1.14 $Y2=1.295
r65 27 30 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.14 $Y=1.02
+ $X2=1.14 $Y2=1.295
r66 25 27 7.36389 $w=2e-07 $l=2.09105e-07 $layer=LI1_cond $X=0.975 $Y=0.92
+ $X2=1.14 $Y2=1.02
r67 25 26 31.3318 $w=1.98e-07 $l=5.65e-07 $layer=LI1_cond $X=0.975 $Y=0.92
+ $X2=0.41 $Y2=0.92
r68 23 28 7.68689 $w=1.75e-07 $l=2.03912e-07 $layer=LI1_cond $X=0.975 $Y=2.117
+ $X2=1.14 $Y2=2.03
r69 23 24 36.4416 $w=1.73e-07 $l=5.75e-07 $layer=LI1_cond $X=0.975 $Y=2.117
+ $X2=0.4 $Y2=2.117
r70 19 24 7.48781 $w=1.75e-07 $l=1.92023e-07 $layer=LI1_cond $X=0.247 $Y=2.205
+ $X2=0.4 $Y2=2.117
r71 19 21 13.4137 $w=3.03e-07 $l=3.55e-07 $layer=LI1_cond $X=0.247 $Y=2.205
+ $X2=0.247 $Y2=2.56
r72 15 26 7.26812 $w=2e-07 $l=2.01901e-07 $layer=LI1_cond $X=0.252 $Y=0.82
+ $X2=0.41 $Y2=0.92
r73 15 17 8.78052 $w=3.13e-07 $l=2.4e-07 $layer=LI1_cond $X=0.252 $Y=0.82
+ $X2=0.252 $Y2=0.58
r74 13 33 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=1.35 $Y=0.58 $X2=1.35
+ $Y2=1.13
r75 9 34 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.32 $Y=2.46 $X2=1.32
+ $Y2=1.8
r76 2 21 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=2.335 $X2=0.265 $Y2=2.56
r77 1 17 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.37 $X2=0.265 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%A_288_74# 1 2 11 15 17 18 23 24 29 30
+ 32
c57 24 0 5.479e-19 $X=2.575 $Y=1.465
r58 29 30 6.71392 $w=3.03e-07 $l=1.65e-07 $layer=LI1_cond $X=1.567 $Y=2.56
+ $X2=1.567 $Y2=2.395
r59 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.575
+ $Y=1.465 $X2=2.575 $Y2=1.465
r60 21 32 1.57103 $w=2.3e-07 $l=1.23e-07 $layer=LI1_cond $X=1.72 $Y=1.495
+ $X2=1.597 $Y2=1.495
r61 21 23 42.8408 $w=2.28e-07 $l=8.55e-07 $layer=LI1_cond $X=1.72 $Y=1.495
+ $X2=2.575 $Y2=1.495
r62 19 32 4.89986 $w=2.45e-07 $l=1.15e-07 $layer=LI1_cond $X=1.597 $Y=1.61
+ $X2=1.597 $Y2=1.495
r63 19 30 36.9252 $w=2.43e-07 $l=7.85e-07 $layer=LI1_cond $X=1.597 $Y=1.61
+ $X2=1.597 $Y2=2.395
r64 18 32 4.89986 $w=2.45e-07 $l=1.15e-07 $layer=LI1_cond $X=1.597 $Y=1.38
+ $X2=1.597 $Y2=1.495
r65 17 27 2.70749 $w=3.05e-07 $l=5.5e-08 $layer=LI1_cond $X=1.597 $Y=0.635
+ $X2=1.597 $Y2=0.58
r66 17 18 35.0437 $w=2.43e-07 $l=7.45e-07 $layer=LI1_cond $X=1.597 $Y=0.635
+ $X2=1.597 $Y2=1.38
r67 13 24 28.6811 $w=2.15e-07 $l=1.80748e-07 $layer=POLY_cond $X=2.695 $Y=1.3
+ $X2=2.662 $Y2=1.465
r68 13 15 155.484 $w=1.8e-07 $l=4e-07 $layer=POLY_cond $X=2.695 $Y=1.3 $X2=2.695
+ $Y2=0.9
r69 9 24 28.6811 $w=2.15e-07 $l=1.65997e-07 $layer=POLY_cond $X=2.66 $Y=1.63
+ $X2=2.662 $Y2=1.465
r70 9 11 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.66 $Y=1.63 $X2=2.66
+ $Y2=2.34
r71 2 29 600 $w=1.7e-07 $l=6.64078e-07 $layer=licon1_PDIFF $count=1 $X=1.445
+ $Y=1.96 $X2=1.58 $Y2=2.56
r72 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.44
+ $Y=0.37 $X2=1.58 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%A_405_138# 1 2 9 13 15 17 19 20 22 26
+ 34
c60 20 0 1.10523e-19 $X=3.032 $Y=1.825
c61 17 0 1.30285e-19 $X=2.91 $Y=1.91
c62 15 0 1.49037e-19 $X=2.91 $Y=1.125
c63 9 0 1.58057e-19 $X=3.215 $Y=2.4
r64 34 37 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=1.46
+ $X2=3.165 $Y2=1.625
r65 34 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=1.46
+ $X2=3.165 $Y2=1.295
r66 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.165
+ $Y=1.46 $X2=3.165 $Y2=1.46
r67 31 33 12.9746 $w=3.15e-07 $l=3.35e-07 $layer=LI1_cond $X=3.095 $Y=1.125
+ $X2=3.095 $Y2=1.46
r68 26 29 3.68142 $w=3.58e-07 $l=1.15e-07 $layer=LI1_cond $X=2.165 $Y=1.91
+ $X2=2.165 $Y2=2.025
r69 22 24 8.00308 $w=3.58e-07 $l=2.5e-07 $layer=LI1_cond $X=2.165 $Y=0.875
+ $X2=2.165 $Y2=1.125
r70 19 33 7.02551 $w=3.15e-07 $l=1.93959e-07 $layer=LI1_cond $X=3.032 $Y=1.625
+ $X2=3.095 $Y2=1.46
r71 19 20 9.4077 $w=2.43e-07 $l=2e-07 $layer=LI1_cond $X=3.032 $Y=1.625
+ $X2=3.032 $Y2=1.825
r72 18 26 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.345 $Y=1.91
+ $X2=2.165 $Y2=1.91
r73 17 20 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=2.91 $Y=1.91
+ $X2=3.032 $Y2=1.825
r74 17 18 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.91 $Y=1.91
+ $X2=2.345 $Y2=1.91
r75 16 24 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.345 $Y=1.125
+ $X2=2.165 $Y2=1.125
r76 15 31 4.34843 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.91 $Y=1.125
+ $X2=3.095 $Y2=1.125
r77 15 16 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.91 $Y=1.125
+ $X2=2.345 $Y2=1.125
r78 13 36 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.205 $Y=0.74
+ $X2=3.205 $Y2=1.295
r79 9 37 301.25 $w=1.8e-07 $l=7.75e-07 $layer=POLY_cond $X=3.215 $Y=2.4
+ $X2=3.215 $Y2=1.625
r80 2 29 600 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_PDIFF $count=1 $X=2.025
+ $Y=1.84 $X2=2.15 $Y2=2.025
r81 1 22 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.69 $X2=2.15 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%VPWR 1 2 9 13 18 19 20 22 35 36 39
r35 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r36 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r37 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r38 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r39 30 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 29 32 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r42 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=0.74 $Y2=3.33
r43 27 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=1.2 $Y2=3.33
r44 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r46 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.74 $Y2=3.33
r47 22 24 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 20 33 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 20 30 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 18 32 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.825 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.825 $Y=3.33
+ $X2=2.99 $Y2=3.33
r52 17 35 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.155 $Y=3.33
+ $X2=3.6 $Y2=3.33
r53 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=3.33
+ $X2=2.99 $Y2=3.33
r54 13 16 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=2.99 $Y=2.27
+ $X2=2.99 $Y2=2.81
r55 11 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=3.245
+ $X2=2.99 $Y2=3.33
r56 11 16 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=2.99 $Y=3.245
+ $X2=2.99 $Y2=2.81
r57 7 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=3.245 $X2=0.74
+ $Y2=3.33
r58 7 9 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.74 $Y=3.245 $X2=0.74
+ $Y2=2.545
r59 2 16 600 $w=1.7e-07 $l=1.06759e-06 $layer=licon1_PDIFF $count=1 $X=2.785
+ $Y=1.84 $X2=2.99 $Y2=2.81
r60 2 13 600 $w=1.7e-07 $l=5.22542e-07 $layer=licon1_PDIFF $count=1 $X=2.785
+ $Y=1.84 $X2=2.99 $Y2=2.27
r61 1 9 600 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.335 $X2=0.74 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%X 1 2 7 8 9 10 11 12 13 25 38 48 52
r22 52 53 5.77907 $w=4.13e-07 $l=1.7e-07 $layer=LI1_cond $X=3.532 $Y=1.985
+ $X2=3.532 $Y2=1.815
r23 36 38 0.361006 $w=4.13e-07 $l=1.3e-08 $layer=LI1_cond $X=3.532 $Y=2.022
+ $X2=3.532 $Y2=2.035
r24 23 48 0.333237 $w=4.13e-07 $l=1.2e-08 $layer=LI1_cond $X=3.532 $Y=0.913
+ $X2=3.532 $Y2=0.925
r25 13 45 0.97194 $w=4.13e-07 $l=3.5e-08 $layer=LI1_cond $X=3.532 $Y=2.775
+ $X2=3.532 $Y2=2.81
r26 12 13 10.2748 $w=4.13e-07 $l=3.7e-07 $layer=LI1_cond $X=3.532 $Y=2.405
+ $X2=3.532 $Y2=2.775
r27 11 36 0.99971 $w=4.13e-07 $l=3.6e-08 $layer=LI1_cond $X=3.532 $Y=1.986
+ $X2=3.532 $Y2=2.022
r28 11 52 0.0277697 $w=4.13e-07 $l=1e-09 $layer=LI1_cond $X=3.532 $Y=1.986
+ $X2=3.532 $Y2=1.985
r29 11 12 9.27508 $w=4.13e-07 $l=3.34e-07 $layer=LI1_cond $X=3.532 $Y=2.071
+ $X2=3.532 $Y2=2.405
r30 11 38 0.99971 $w=4.13e-07 $l=3.6e-08 $layer=LI1_cond $X=3.532 $Y=2.071
+ $X2=3.532 $Y2=2.035
r31 10 53 5.96091 $w=2.88e-07 $l=1.5e-07 $layer=LI1_cond $X=3.595 $Y=1.665
+ $X2=3.595 $Y2=1.815
r32 9 10 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=3.595 $Y=1.295
+ $X2=3.595 $Y2=1.665
r33 9 50 6.9544 $w=2.88e-07 $l=1.75e-07 $layer=LI1_cond $X=3.595 $Y=1.295
+ $X2=3.595 $Y2=1.12
r34 8 50 5.4736 $w=4.13e-07 $l=1.59e-07 $layer=LI1_cond $X=3.532 $Y=0.961
+ $X2=3.532 $Y2=1.12
r35 8 48 0.99971 $w=4.13e-07 $l=3.6e-08 $layer=LI1_cond $X=3.532 $Y=0.961
+ $X2=3.532 $Y2=0.925
r36 8 23 1.02748 $w=4.13e-07 $l=3.7e-08 $layer=LI1_cond $X=3.532 $Y=0.876
+ $X2=3.532 $Y2=0.913
r37 7 8 8.91408 $w=4.13e-07 $l=3.21e-07 $layer=LI1_cond $X=3.532 $Y=0.555
+ $X2=3.532 $Y2=0.876
r38 7 25 0.97194 $w=4.13e-07 $l=3.5e-08 $layer=LI1_cond $X=3.532 $Y=0.555
+ $X2=3.532 $Y2=0.52
r39 2 52 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.305
+ $Y=1.84 $X2=3.445 $Y2=1.985
r40 2 45 400 $w=1.7e-07 $l=1.03764e-06 $layer=licon1_PDIFF $count=1 $X=3.305
+ $Y=1.84 $X2=3.445 $Y2=2.81
r41 1 25 91 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=2 $X=3.28
+ $Y=0.37 $X2=3.42 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_MS__DLYGATE4SD2_1%VGND 1 2 9 13 16 17 18 20 33 34 37
r38 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r39 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r40 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r41 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r42 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r43 27 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r44 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r45 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.75
+ $Y2=0
r46 25 27 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.2
+ $Y2=0
r47 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r48 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r49 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.75
+ $Y2=0
r50 20 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r51 18 31 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r52 18 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r53 16 30 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.825 $Y=0 $X2=2.64
+ $Y2=0
r54 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.825 $Y=0 $X2=2.99
+ $Y2=0
r55 15 33 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.155 $Y=0 $X2=3.6
+ $Y2=0
r56 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=0 $X2=2.99
+ $Y2=0
r57 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=0.085
+ $X2=2.99 $Y2=0
r58 11 13 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=2.99 $Y=0.085
+ $X2=2.99 $Y2=0.62
r59 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085 $X2=0.75
+ $Y2=0
r60 7 9 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.75 $Y=0.085 $X2=0.75
+ $Y2=0.565
r61 2 13 182 $w=1.7e-07 $l=2.37434e-07 $layer=licon1_NDIFF $count=1 $X=2.785
+ $Y=0.69 $X2=2.99 $Y2=0.62
r62 1 9 182 $w=1.7e-07 $l=2.75772e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.37 $X2=0.75 $Y2=0.565
.ends


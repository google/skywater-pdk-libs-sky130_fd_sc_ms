# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__a22oi_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 5.635000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 1.350000 7.465000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.265000 1.350000 3.275000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.116000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.350000 1.955000 1.780000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  2.172800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635000 1.950000 3.615000 2.120000 ;
        RECT 0.635000 2.120000 0.885000 2.735000 ;
        RECT 1.615000 2.120000 1.785000 2.735000 ;
        RECT 2.350000 0.595000 2.680000 1.010000 ;
        RECT 2.350000 1.010000 5.780000 1.130000 ;
        RECT 2.350000 1.130000 4.195000 1.180000 ;
        RECT 2.515000 2.120000 2.685000 2.735000 ;
        RECT 3.210000 0.770000 3.990000 0.850000 ;
        RECT 3.210000 0.850000 5.780000 1.010000 ;
        RECT 3.415000 2.120000 3.615000 2.735000 ;
        RECT 3.445000 1.180000 4.195000 1.520000 ;
        RECT 3.445000 1.520000 3.615000 1.950000 ;
        RECT 5.450000 0.770000 5.780000 0.850000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.185000  1.820000 0.435000 2.905000 ;
      RECT 0.185000  2.905000 4.035000 3.075000 ;
      RECT 0.200000  0.350000 0.450000 1.010000 ;
      RECT 0.200000  1.010000 2.170000 1.180000 ;
      RECT 0.630000  0.085000 0.880000 0.840000 ;
      RECT 1.060000  0.350000 1.310000 1.010000 ;
      RECT 1.085000  2.290000 1.415000 2.905000 ;
      RECT 1.490000  0.085000 1.820000 0.840000 ;
      RECT 1.985000  2.290000 2.315000 2.905000 ;
      RECT 2.000000  0.255000 3.970000 0.425000 ;
      RECT 2.000000  0.425000 2.170000 1.010000 ;
      RECT 2.860000  0.425000 3.970000 0.600000 ;
      RECT 2.860000  0.600000 3.030000 0.840000 ;
      RECT 2.885000  2.290000 3.215000 2.905000 ;
      RECT 3.785000  1.820000 4.035000 1.950000 ;
      RECT 3.785000  1.950000 7.945000 2.120000 ;
      RECT 3.785000  2.120000 4.035000 2.905000 ;
      RECT 4.160000  0.350000 6.130000 0.600000 ;
      RECT 4.160000  0.600000 4.490000 0.680000 ;
      RECT 4.235000  2.290000 4.565000 3.245000 ;
      RECT 4.765000  2.120000 5.015000 2.980000 ;
      RECT 5.185000  2.290000 5.645000 3.245000 ;
      RECT 5.815000  2.120000 6.065000 2.980000 ;
      RECT 5.960000  0.600000 6.130000 1.010000 ;
      RECT 5.960000  1.010000 7.930000 1.180000 ;
      RECT 6.265000  2.290000 6.595000 3.245000 ;
      RECT 6.310000  0.085000 6.560000 0.840000 ;
      RECT 6.740000  0.350000 6.990000 1.010000 ;
      RECT 6.795000  2.120000 6.965000 2.980000 ;
      RECT 7.165000  2.290000 7.495000 3.245000 ;
      RECT 7.170000  0.085000 7.420000 0.840000 ;
      RECT 7.600000  0.350000 7.930000 1.010000 ;
      RECT 7.695000  1.820000 7.945000 1.950000 ;
      RECT 7.695000  2.120000 7.945000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_ms__a22oi_4

* File: sky130_fd_sc_ms__nand4_4.pex.spice
* Created: Wed Sep  2 12:14:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NAND4_4%D 3 7 9 13 17 21 25 27 28 29 30 31 32 33 34
+ 52
c74 21 0 7.27676e-20 $X=2.195 $Y=0.74
r75 51 52 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=2.195 $Y=1.515
+ $X2=2.26 $Y2=1.515
r76 49 51 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.105 $Y=1.515
+ $X2=2.195 $Y2=1.515
r77 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.105
+ $Y=1.515 $X2=2.105 $Y2=1.515
r78 47 49 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=1.76 $Y=1.515
+ $X2=2.105 $Y2=1.515
r79 46 47 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=1.495 $Y=1.515
+ $X2=1.76 $Y2=1.515
r80 44 46 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=1.425 $Y=1.515
+ $X2=1.495 $Y2=1.515
r81 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.425
+ $Y=1.515 $X2=1.425 $Y2=1.515
r82 41 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.745
+ $Y=1.515 $X2=0.745 $Y2=1.515
r83 34 50 1.47406 $w=4.28e-07 $l=5.5e-08 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.105 $Y2=1.565
r84 33 50 11.3904 $w=4.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=2.105 $Y2=1.565
r85 33 45 6.83426 $w=4.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.425 $Y2=1.565
r86 32 45 6.03022 $w=4.28e-07 $l=2.25e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.425 $Y2=1.565
r87 32 42 12.1945 $w=4.28e-07 $l=4.55e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=0.745 $Y2=1.565
r88 31 42 0.670025 $w=4.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.745 $Y2=1.565
r89 30 31 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.72 $Y2=1.565
r90 28 41 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=0.92 $Y=1.515
+ $X2=0.745 $Y2=1.515
r91 28 29 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.92 $Y=1.515
+ $X2=0.995 $Y2=1.515
r92 27 41 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=0.57 $Y=1.515
+ $X2=0.745 $Y2=1.515
r93 23 52 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=1.68
+ $X2=2.26 $Y2=1.515
r94 23 25 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.26 $Y=1.68
+ $X2=2.26 $Y2=2.4
r95 19 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.35
+ $X2=2.195 $Y2=1.515
r96 19 21 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.195 $Y=1.35
+ $X2=2.195 $Y2=0.74
r97 15 47 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.76 $Y=1.68
+ $X2=1.76 $Y2=1.515
r98 15 17 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.76 $Y=1.68
+ $X2=1.76 $Y2=2.4
r99 11 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.495 $Y=1.35
+ $X2=1.495 $Y2=1.515
r100 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.495 $Y=1.35
+ $X2=1.495 $Y2=0.74
r101 10 29 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.07 $Y=1.515
+ $X2=0.995 $Y2=1.515
r102 9 44 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=1.42 $Y=1.515
+ $X2=1.425 $Y2=1.515
r103 9 10 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=1.42 $Y=1.515
+ $X2=1.07 $Y2=1.515
r104 5 29 16.9349 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=1.515
r105 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=0.74
r106 1 27 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.57 $Y2=1.515
r107 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4_4%C 3 7 11 15 19 23 25 26 27 28 48
r58 46 48 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=3.805 $Y=1.515
+ $X2=3.985 $Y2=1.515
r59 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.805
+ $Y=1.515 $X2=3.805 $Y2=1.515
r60 44 46 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.555 $Y=1.515
+ $X2=3.805 $Y2=1.515
r61 43 44 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.54 $Y=1.515
+ $X2=3.555 $Y2=1.515
r62 41 43 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.465 $Y=1.515
+ $X2=3.54 $Y2=1.515
r63 41 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.465
+ $Y=1.515 $X2=3.465 $Y2=1.515
r64 39 41 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.125 $Y=1.515
+ $X2=3.465 $Y2=1.515
r65 37 39 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.785 $Y=1.515
+ $X2=3.125 $Y2=1.515
r66 37 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.785
+ $Y=1.515 $X2=2.785 $Y2=1.515
r67 35 37 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.71 $Y=1.515
+ $X2=2.785 $Y2=1.515
r68 33 35 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.695 $Y=1.515
+ $X2=2.71 $Y2=1.515
r69 28 47 7.37028 $w=4.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=3.805 $Y2=1.565
r70 27 47 5.4942 $w=4.28e-07 $l=2.05e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.805 $Y2=1.565
r71 27 42 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.465 $Y2=1.565
r72 26 42 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.465 $Y2=1.565
r73 26 38 8.97834 $w=4.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=2.785 $Y2=1.565
r74 25 38 3.88615 $w=4.28e-07 $l=1.45e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.785 $Y2=1.565
r75 21 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.985 $Y=1.35
+ $X2=3.985 $Y2=1.515
r76 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.985 $Y=1.35
+ $X2=3.985 $Y2=0.74
r77 17 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.555 $Y=1.35
+ $X2=3.555 $Y2=1.515
r78 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.555 $Y=1.35
+ $X2=3.555 $Y2=0.74
r79 13 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.54 $Y=1.68
+ $X2=3.54 $Y2=1.515
r80 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.54 $Y=1.68
+ $X2=3.54 $Y2=2.4
r81 9 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.125 $Y=1.35
+ $X2=3.125 $Y2=1.515
r82 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.125 $Y=1.35
+ $X2=3.125 $Y2=0.74
r83 5 35 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.68
+ $X2=2.71 $Y2=1.515
r84 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.71 $Y=1.68 $X2=2.71
+ $Y2=2.4
r85 1 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.695 $Y=1.35
+ $X2=2.695 $Y2=1.515
r86 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.695 $Y=1.35
+ $X2=2.695 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4_4%B 3 7 11 15 19 23 25 26 27 28 48
r65 46 48 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=5.995 $Y=1.515
+ $X2=6.265 $Y2=1.515
r66 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.995
+ $Y=1.515 $X2=5.995 $Y2=1.515
r67 44 46 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=5.835 $Y=1.515
+ $X2=5.995 $Y2=1.515
r68 43 44 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=5.405 $Y=1.515
+ $X2=5.835 $Y2=1.515
r69 42 43 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.39 $Y=1.515
+ $X2=5.405 $Y2=1.515
r70 40 42 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.315 $Y=1.515
+ $X2=5.39 $Y2=1.515
r71 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.315
+ $Y=1.515 $X2=5.315 $Y2=1.515
r72 38 40 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.975 $Y=1.515
+ $X2=5.315 $Y2=1.515
r73 36 38 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.635 $Y=1.515
+ $X2=4.975 $Y2=1.515
r74 36 37 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.635
+ $Y=1.515 $X2=4.635 $Y2=1.515
r75 33 36 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.56 $Y=1.515
+ $X2=4.635 $Y2=1.515
r76 28 47 0.134005 $w=4.28e-07 $l=5e-09 $layer=LI1_cond $X=6 $Y=1.565 $X2=5.995
+ $Y2=1.565
r77 27 47 12.7305 $w=4.28e-07 $l=4.75e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.995 $Y2=1.565
r78 27 41 5.4942 $w=4.28e-07 $l=2.05e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.315 $Y2=1.565
r79 26 41 7.37028 $w=4.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.315 $Y2=1.565
r80 26 37 10.8544 $w=4.28e-07 $l=4.05e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=4.635 $Y2=1.565
r81 25 37 2.01008 $w=4.28e-07 $l=7.5e-08 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.635 $Y2=1.565
r82 21 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.265 $Y=1.35
+ $X2=6.265 $Y2=1.515
r83 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.265 $Y=1.35
+ $X2=6.265 $Y2=0.74
r84 17 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.835 $Y=1.35
+ $X2=5.835 $Y2=1.515
r85 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.835 $Y=1.35
+ $X2=5.835 $Y2=0.74
r86 13 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.405 $Y=1.35
+ $X2=5.405 $Y2=1.515
r87 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.405 $Y=1.35
+ $X2=5.405 $Y2=0.74
r88 9 42 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.39 $Y=1.68
+ $X2=5.39 $Y2=1.515
r89 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.39 $Y=1.68 $X2=5.39
+ $Y2=2.4
r90 5 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.975 $Y=1.35
+ $X2=4.975 $Y2=1.515
r91 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.975 $Y=1.35
+ $X2=4.975 $Y2=0.74
r92 1 33 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.56 $Y=1.68
+ $X2=4.56 $Y2=1.515
r93 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.56 $Y=1.68 $X2=4.56
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4_4%A 3 7 11 15 19 23 25 26 27 28 29 33
r67 45 47 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=7.24 $Y=1.515
+ $X2=7.555 $Y2=1.515
r68 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.24
+ $Y=1.515 $X2=7.24 $Y2=1.515
r69 43 45 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=7.2 $Y=1.515 $X2=7.24
+ $Y2=1.515
r70 42 43 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.125 $Y=1.515
+ $X2=7.2 $Y2=1.515
r71 40 42 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=6.9 $Y=1.515
+ $X2=7.125 $Y2=1.515
r72 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.9
+ $Y=1.515 $X2=6.9 $Y2=1.515
r73 37 40 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=6.695 $Y=1.515
+ $X2=6.9 $Y2=1.515
r74 33 47 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.63 $Y=1.515
+ $X2=7.555 $Y2=1.515
r75 33 35 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=7.63 $Y=1.515
+ $X2=7.92 $Y2=1.515
r76 29 35 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.92
+ $Y=1.515 $X2=7.92 $Y2=1.515
r77 28 29 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.92 $Y2=1.565
r78 28 46 5.3602 $w=4.28e-07 $l=2e-07 $layer=LI1_cond $X=7.44 $Y=1.565 $X2=7.24
+ $Y2=1.565
r79 27 46 7.50428 $w=4.28e-07 $l=2.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.24 $Y2=1.565
r80 27 41 1.60806 $w=4.28e-07 $l=6e-08 $layer=LI1_cond $X=6.96 $Y=1.565 $X2=6.9
+ $Y2=1.565
r81 25 35 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=8.04 $Y=1.515
+ $X2=7.92 $Y2=1.515
r82 25 26 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.04 $Y=1.515 $X2=8.13
+ $Y2=1.515
r83 21 26 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=8.145 $Y=1.35
+ $X2=8.13 $Y2=1.515
r84 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.145 $Y=1.35
+ $X2=8.145 $Y2=0.74
r85 17 26 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=8.13 $Y=1.68
+ $X2=8.13 $Y2=1.515
r86 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.13 $Y=1.68
+ $X2=8.13 $Y2=2.4
r87 13 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.555 $Y=1.35
+ $X2=7.555 $Y2=1.515
r88 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.555 $Y=1.35
+ $X2=7.555 $Y2=0.74
r89 9 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.2 $Y=1.68 $X2=7.2
+ $Y2=1.515
r90 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.2 $Y=1.68 $X2=7.2
+ $Y2=2.4
r91 5 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.125 $Y=1.35
+ $X2=7.125 $Y2=1.515
r92 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.125 $Y=1.35
+ $X2=7.125 $Y2=0.74
r93 1 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.695 $Y=1.35
+ $X2=6.695 $Y2=1.515
r94 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.695 $Y=1.35
+ $X2=6.695 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4_4%VPWR 1 2 3 4 5 18 20 24 26 28 30 32 33 42 61
+ 64 71 82 85
r66 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r67 81 82 13.5255 $w=1.123e-06 $l=1.65e-07 $layer=LI1_cond $X=6.975 $Y=2.852
+ $X2=7.14 $Y2=2.852
r68 78 81 0.162667 $w=1.123e-06 $l=1.5e-08 $layer=LI1_cond $X=6.96 $Y=2.852
+ $X2=6.975 $Y2=2.852
r69 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r70 76 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r71 75 78 10.4107 $w=1.123e-06 $l=9.6e-07 $layer=LI1_cond $X=6 $Y=2.852 $X2=6.96
+ $Y2=2.852
r72 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r73 73 75 4.17511 $w=1.123e-06 $l=3.85e-07 $layer=LI1_cond $X=5.615 $Y=2.852
+ $X2=6 $Y2=2.852
r74 70 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r75 69 73 1.03022 $w=1.123e-06 $l=9.5e-08 $layer=LI1_cond $X=5.52 $Y=2.852
+ $X2=5.615 $Y2=2.852
r76 69 71 12.4953 $w=1.123e-06 $l=7e-08 $layer=LI1_cond $X=5.52 $Y=2.852
+ $X2=5.45 $Y2=2.852
r77 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r78 65 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r79 64 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r80 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r81 62 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r82 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r83 56 59 2.93013 $w=1.374e-06 $l=3.3e-07 $layer=LI1_cond $X=1.2 $Y=2.682
+ $X2=1.53 $Y2=2.682
r84 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r85 53 56 4.21761 $w=1.374e-06 $l=4.75e-07 $layer=LI1_cond $X=0.725 $Y=2.682
+ $X2=1.2 $Y2=2.682
r86 51 53 3.55167 $w=1.374e-06 $l=4e-07 $layer=LI1_cond $X=0.325 $Y=2.682
+ $X2=0.725 $Y2=2.682
r87 49 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r88 48 51 0.754731 $w=1.374e-06 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.682
+ $X2=0.325 $Y2=2.682
r89 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r90 46 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r91 46 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=6.96 $Y2=3.33
r92 45 82 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=7.92 $Y=3.33
+ $X2=7.14 $Y2=3.33
r93 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r94 42 84 4.72267 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=8.19 $Y=3.33
+ $X2=8.415 $Y2=3.33
r95 42 45 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.19 $Y=3.33 $X2=7.92
+ $Y2=3.33
r96 41 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r97 40 71 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=5.45 $Y2=3.33
r98 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r99 38 64 15.5046 $w=1.7e-07 $l=4.5e-07 $layer=LI1_cond $X=4.5 $Y=3.33 $X2=4.05
+ $Y2=3.33
r100 38 40 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=4.5 $Y=3.33 $X2=4.56
+ $Y2=3.33
r101 36 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r102 36 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r103 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r104 33 59 14.335 $w=1.374e-06 $l=7.05453e-07 $layer=LI1_cond $X=1.65 $Y=3.33
+ $X2=1.53 $Y2=2.682
r105 33 35 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.65 $Y=3.33
+ $X2=2.16 $Y2=3.33
r106 32 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.32 $Y=3.33
+ $X2=2.485 $Y2=3.33
r107 32 35 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.32 $Y=3.33
+ $X2=2.16 $Y2=3.33
r108 30 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r109 30 65 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r110 26 84 3.0435 $w=3.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=8.355 $Y=3.245
+ $X2=8.415 $Y2=3.33
r111 26 28 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=8.355 $Y=3.245
+ $X2=8.355 $Y2=2.415
r112 22 64 3.34993 $w=9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.05 $Y=3.245 $X2=4.05
+ $Y2=3.33
r113 22 24 11.2511 $w=8.98e-07 $l=8.3e-07 $layer=LI1_cond $X=4.05 $Y=3.245
+ $X2=4.05 $Y2=2.415
r114 21 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.65 $Y=3.33
+ $X2=2.485 $Y2=3.33
r115 20 64 15.5046 $w=1.7e-07 $l=4.5e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.05
+ $Y2=3.33
r116 20 21 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=2.65 $Y2=3.33
r117 16 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.485 $Y=3.245
+ $X2=2.485 $Y2=3.33
r118 16 18 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.485 $Y=3.245
+ $X2=2.485 $Y2=2.455
r119 5 28 300 $w=1.7e-07 $l=6.38944e-07 $layer=licon1_PDIFF $count=2 $X=8.22
+ $Y=1.84 $X2=8.355 $Y2=2.415
r120 4 81 120 $w=1.7e-07 $l=1.75916e-06 $layer=licon1_PDIFF $count=5 $X=5.48
+ $Y=1.84 $X2=6.975 $Y2=2.415
r121 4 73 120 $w=1.7e-07 $l=6.38944e-07 $layer=licon1_PDIFF $count=5 $X=5.48
+ $Y=1.84 $X2=5.615 $Y2=2.415
r122 3 24 150 $w=1.7e-07 $l=9.49947e-07 $layer=licon1_PDIFF $count=4 $X=3.63
+ $Y=1.84 $X2=4.335 $Y2=2.415
r123 2 18 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=2.35
+ $Y=1.84 $X2=2.485 $Y2=2.455
r124 1 59 200 $w=1.7e-07 $l=1.6745e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=1.84 $X2=1.53 $Y2=2.455
r125 1 53 200 $w=1.7e-07 $l=1.23526e-06 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=1.84 $X2=0.725 $Y2=2.815
r126 1 53 200 $w=1.7e-07 $l=7.14388e-07 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=1.84 $X2=0.725 $Y2=2.115
r127 1 51 200 $w=1.7e-07 $l=7.03616e-07 $layer=licon1_PDIFF $count=3 $X=0.135
+ $Y=1.84 $X2=0.325 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4_4%Y 1 2 3 4 5 6 19 21 23 27 29 33 35 38 41 43
+ 45 50 52 56 59 60 63 64
r96 63 64 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.4 $Y=1.295 $X2=8.4
+ $Y2=1.665
r97 62 64 14.2803 $w=2.28e-07 $l=2.85e-07 $layer=LI1_cond $X=8.4 $Y=1.95 $X2=8.4
+ $Y2=1.665
r98 61 63 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.4 $Y=1.13 $X2=8.4
+ $Y2=1.295
r99 58 60 4.02231 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=7.85 $Y=0.965
+ $X2=7.945 $Y2=0.965
r100 58 59 4.02231 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=7.85 $Y=0.965
+ $X2=7.755 $Y2=0.965
r101 46 56 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=8.01 $Y=2.035
+ $X2=7.665 $Y2=2.035
r102 45 62 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=8.285 $Y=2.035
+ $X2=8.4 $Y2=1.95
r103 45 46 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.285 $Y=2.035
+ $X2=8.01 $Y2=2.035
r104 43 61 6.8319 $w=2.5e-07 $l=1.73205e-07 $layer=LI1_cond $X=8.285 $Y=1.005
+ $X2=8.4 $Y2=1.13
r105 43 60 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=8.285 $Y=1.005
+ $X2=7.945 $Y2=1.005
r106 39 56 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.665 $Y=2.12
+ $X2=7.665 $Y2=2.035
r107 39 41 5.11367 $w=6.88e-07 $l=2.95e-07 $layer=LI1_cond $X=7.665 $Y=2.12
+ $X2=7.665 $Y2=2.415
r108 38 54 4.23145 $w=3.08e-07 $l=1.13248e-07 $layer=LI1_cond $X=7.005 $Y=1.005
+ $X2=6.91 $Y2=0.965
r109 38 59 34.5733 $w=2.48e-07 $l=7.5e-07 $layer=LI1_cond $X=7.005 $Y=1.005
+ $X2=7.755 $Y2=1.005
r110 36 52 12.6759 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=5.28 $Y=2.035
+ $X2=4.975 $Y2=2.035
r111 35 56 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=7.32 $Y=2.035
+ $X2=7.665 $Y2=2.035
r112 35 36 133.091 $w=1.68e-07 $l=2.04e-06 $layer=LI1_cond $X=7.32 $Y=2.035
+ $X2=5.28 $Y2=2.035
r113 31 52 2.55884 $w=6.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.975 $Y=2.12
+ $X2=4.975 $Y2=2.035
r114 31 33 5.78431 $w=6.08e-07 $l=2.95e-07 $layer=LI1_cond $X=4.975 $Y=2.12
+ $X2=4.975 $Y2=2.415
r115 30 50 12.6759 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=3.43 $Y=2.035
+ $X2=3.125 $Y2=2.035
r116 29 52 12.6759 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=4.67 $Y=2.035
+ $X2=4.975 $Y2=2.035
r117 29 30 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=4.67 $Y=2.035
+ $X2=3.43 $Y2=2.035
r118 25 50 2.55884 $w=6.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.125 $Y=2.12
+ $X2=3.125 $Y2=2.035
r119 25 27 5.78431 $w=6.08e-07 $l=2.95e-07 $layer=LI1_cond $X=3.125 $Y=2.12
+ $X2=3.125 $Y2=2.415
r120 24 48 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.15 $Y=2.035
+ $X2=1.985 $Y2=2.035
r121 23 50 12.6759 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=2.82 $Y=2.035
+ $X2=3.125 $Y2=2.035
r122 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.82 $Y=2.035
+ $X2=2.15 $Y2=2.035
r123 19 48 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=2.12
+ $X2=1.985 $Y2=2.035
r124 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.985 $Y=2.12
+ $X2=1.985 $Y2=2.415
r125 6 56 300 $w=1.7e-07 $l=7.05797e-07 $layer=licon1_PDIFF $count=2 $X=7.29
+ $Y=1.84 $X2=7.905 $Y2=2.035
r126 6 41 150 $w=1.7e-07 $l=8.55482e-07 $layer=licon1_PDIFF $count=4 $X=7.29
+ $Y=1.84 $X2=7.905 $Y2=2.415
r127 5 52 300 $w=1.7e-07 $l=6.0469e-07 $layer=licon1_PDIFF $count=2 $X=4.65
+ $Y=1.84 $X2=5.165 $Y2=2.035
r128 5 33 150 $w=1.7e-07 $l=7.91675e-07 $layer=licon1_PDIFF $count=4 $X=4.65
+ $Y=1.84 $X2=5.165 $Y2=2.415
r129 4 50 300 $w=1.7e-07 $l=6.0469e-07 $layer=licon1_PDIFF $count=2 $X=2.8
+ $Y=1.84 $X2=3.315 $Y2=2.035
r130 4 27 150 $w=1.7e-07 $l=7.91675e-07 $layer=licon1_PDIFF $count=4 $X=2.8
+ $Y=1.84 $X2=3.315 $Y2=2.415
r131 3 48 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=1.85
+ $Y=1.84 $X2=1.985 $Y2=2.035
r132 3 21 300 $w=1.7e-07 $l=6.38944e-07 $layer=licon1_PDIFF $count=2 $X=1.85
+ $Y=1.84 $X2=1.985 $Y2=2.415
r133 2 58 182 $w=1.7e-07 $l=6.96366e-07 $layer=licon1_NDIFF $count=1 $X=7.63
+ $Y=0.37 $X2=7.85 $Y2=0.965
r134 1 54 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=6.77
+ $Y=0.37 $X2=6.91 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4_4%A_27_74# 1 2 3 4 5 18 20 21 24 26 28 31 36
+ 38
r62 34 36 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=3.34 $Y=0.515
+ $X2=4.2 $Y2=0.515
r63 32 40 3.40825 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=0.515
+ $X2=2.41 $Y2=0.515
r64 32 34 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=2.575 $Y=0.515
+ $X2=3.34 $Y2=0.515
r65 29 31 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=2.41 $Y=1.01
+ $X2=2.41 $Y2=0.965
r66 28 40 3.40825 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.41 $Y=0.68
+ $X2=2.41 $Y2=0.515
r67 28 31 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.41 $Y=0.68
+ $X2=2.41 $Y2=0.965
r68 27 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=1.095
+ $X2=1.28 $Y2=1.095
r69 26 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.245 $Y=1.095
+ $X2=2.41 $Y2=1.01
r70 26 27 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=2.245 $Y=1.095
+ $X2=1.445 $Y2=1.095
r71 22 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=1.01 $X2=1.28
+ $Y2=1.095
r72 22 24 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.28 $Y=1.01
+ $X2=1.28 $Y2=0.515
r73 20 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=1.095
+ $X2=1.28 $Y2=1.095
r74 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=1.095
+ $X2=0.445 $Y2=1.095
r75 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.445 $Y2=1.095
r76 16 18 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.28 $Y=1.01
+ $X2=0.28 $Y2=0.515
r77 5 36 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.06
+ $Y=0.37 $X2=4.2 $Y2=0.515
r78 4 34 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.2
+ $Y=0.37 $X2=3.34 $Y2=0.515
r79 3 40 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.37 $X2=2.41 $Y2=0.515
r80 3 31 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.37 $X2=2.41 $Y2=0.965
r81 2 24 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.28 $Y2=0.515
r82 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4_4%VGND 1 2 9 11 15 17 19 29 30 33 36
r68 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r69 34 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r70 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r71 29 30 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r72 27 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r73 26 29 407.102 $w=1.68e-07 $l=6.24e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=8.4
+ $Y2=0
r74 26 27 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r75 24 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=1.78
+ $Y2=0
r76 24 26 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=2.16
+ $Y2=0
r77 22 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r78 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r79 19 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r80 19 21 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r81 17 30 1.13724 $w=4.9e-07 $l=4.08e-06 $layer=MET1_cond $X=4.32 $Y=0 $X2=8.4
+ $Y2=0
r82 17 27 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=4.32 $Y=0 $X2=2.16
+ $Y2=0
r83 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0
r84 13 15 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.78 $Y=0.085
+ $X2=1.78 $Y2=0.675
r85 12 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r86 11 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.615 $Y=0 $X2=1.78
+ $Y2=0
r87 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=0 $X2=0.945
+ $Y2=0
r88 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0
r89 7 9 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0.675
r90 2 15 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.37 $X2=1.78 $Y2=0.675
r91 1 9 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4_4%A_554_74# 1 2 3 4 13 21 23 26 27
c40 13 0 7.27676e-20 $X=3.795 $Y=0.99
r41 25 27 4.02231 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=5.19 $Y=0.965
+ $X2=5.285 $Y2=0.965
r42 25 26 4.02231 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=5.19 $Y=0.965
+ $X2=5.095 $Y2=0.965
r43 23 26 53.4734 $w=2.48e-07 $l=1.16e-06 $layer=LI1_cond $X=3.935 $Y=1.005
+ $X2=5.095 $Y2=1.005
r44 21 29 4.23145 $w=3.08e-07 $l=1.13248e-07 $layer=LI1_cond $X=5.955 $Y=1.005
+ $X2=6.05 $Y2=0.965
r45 21 27 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=5.955 $Y=1.005
+ $X2=5.285 $Y2=1.005
r46 15 18 35.3965 $w=2.78e-07 $l=8.6e-07 $layer=LI1_cond $X=2.91 $Y=0.99
+ $X2=3.77 $Y2=0.99
r47 13 23 5.9212 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=3.795 $Y=0.99
+ $X2=3.935 $Y2=0.99
r48 13 18 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=3.795 $Y=0.99
+ $X2=3.77 $Y2=0.99
r49 4 29 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=5.91
+ $Y=0.37 $X2=6.05 $Y2=0.965
r50 3 25 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=5.05
+ $Y=0.37 $X2=5.19 $Y2=0.965
r51 2 18 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=3.63
+ $Y=0.37 $X2=3.77 $Y2=0.95
r52 1 15 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=2.77
+ $Y=0.37 $X2=2.91 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4_4%A_923_74# 1 2 3 4 5 22 24 31 32 35 36 39 40
+ 41
r62 41 44 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=8.36 $Y=0.435
+ $X2=8.36 $Y2=0.545
r63 38 40 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=7.34 $Y=0.53
+ $X2=7.505 $Y2=0.53
r64 38 39 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=7.34 $Y=0.53
+ $X2=7.175 $Y2=0.53
r65 36 39 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.645 $Y=0.435
+ $X2=7.175 $Y2=0.435
r66 34 36 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=6.48 $Y=0.53
+ $X2=6.645 $Y2=0.53
r67 34 35 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=6.48 $Y=0.53
+ $X2=6.315 $Y2=0.53
r68 32 35 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.785 $Y=0.435
+ $X2=6.315 $Y2=0.435
r69 30 32 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.62 $Y=0.53
+ $X2=5.785 $Y2=0.53
r70 30 31 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.62 $Y=0.53
+ $X2=5.455 $Y2=0.53
r71 24 27 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=4.76 $Y=0.435
+ $X2=4.76 $Y2=0.545
r72 22 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.195 $Y=0.435
+ $X2=8.36 $Y2=0.435
r73 22 40 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.195 $Y=0.435
+ $X2=7.505 $Y2=0.435
r74 17 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.925 $Y=0.435
+ $X2=4.76 $Y2=0.435
r75 17 31 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.925 $Y=0.435
+ $X2=5.455 $Y2=0.435
r76 5 44 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=8.22
+ $Y=0.37 $X2=8.36 $Y2=0.545
r77 4 38 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=7.2
+ $Y=0.37 $X2=7.34 $Y2=0.545
r78 3 34 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=6.34
+ $Y=0.37 $X2=6.48 $Y2=0.545
r79 2 30 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=5.48
+ $Y=0.37 $X2=5.62 $Y2=0.545
r80 1 27 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=4.615
+ $Y=0.37 $X2=4.76 $Y2=0.545
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__dlclkp_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__dlclkp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN GATE
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.530000 1.430000 1.800000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  1.036000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.795000 1.550000 8.515000 1.720000 ;
        RECT 6.795000 1.720000 7.125000 2.980000 ;
        RECT 6.835000 0.350000 7.165000 1.210000 ;
        RECT 6.835000 1.210000 8.015000 1.380000 ;
        RECT 7.745000 1.720000 8.515000 1.780000 ;
        RECT 7.745000 1.780000 7.995000 2.980000 ;
        RECT 7.765000 0.350000 8.015000 1.210000 ;
        RECT 7.805000 1.380000 8.015000 1.550000 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.574800 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.400000 1.360000 5.070000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.640000 0.085000 ;
        RECT 0.550000  0.085000 0.925000 0.680000 ;
        RECT 3.315000  0.085000 3.645000 0.850000 ;
        RECT 4.780000  0.085000 5.110000 0.850000 ;
        RECT 6.160000  0.085000 6.655000 0.500000 ;
        RECT 7.335000  0.085000 7.585000 1.040000 ;
        RECT 8.195000  0.085000 8.525000 1.040000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 8.640000 3.415000 ;
        RECT 0.785000 2.310000 1.160000 3.245000 ;
        RECT 3.110000 2.860000 3.440000 3.245000 ;
        RECT 4.740000 2.090000 5.070000 3.245000 ;
        RECT 5.740000 2.160000 6.625000 3.245000 ;
        RECT 7.295000 1.890000 7.545000 3.245000 ;
        RECT 8.195000 1.950000 8.525000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.115000 0.350000 0.365000 0.850000 ;
      RECT 0.115000 0.850000 1.265000 1.020000 ;
      RECT 0.115000 1.020000 0.365000 1.820000 ;
      RECT 0.115000 1.820000 0.540000 2.980000 ;
      RECT 0.535000 1.190000 1.605000 1.360000 ;
      RECT 0.535000 1.360000 0.880000 1.550000 ;
      RECT 0.710000 1.550000 0.880000 1.970000 ;
      RECT 0.710000 1.970000 1.605000 2.140000 ;
      RECT 1.095000 0.255000 3.145000 0.425000 ;
      RECT 1.095000 0.425000 1.265000 0.850000 ;
      RECT 1.435000 0.650000 2.330000 0.980000 ;
      RECT 1.435000 0.980000 1.605000 1.190000 ;
      RECT 1.435000 2.140000 1.605000 2.520000 ;
      RECT 1.435000 2.520000 2.485000 2.850000 ;
      RECT 1.775000 1.150000 2.065000 2.050000 ;
      RECT 1.775000 2.050000 3.475000 2.350000 ;
      RECT 2.305000 1.360000 4.155000 1.530000 ;
      RECT 2.305000 1.530000 2.635000 1.805000 ;
      RECT 2.815000 0.425000 3.145000 1.020000 ;
      RECT 2.815000 1.020000 5.430000 1.190000 ;
      RECT 3.305000 1.700000 3.655000 1.960000 ;
      RECT 3.305000 1.960000 3.475000 2.050000 ;
      RECT 3.305000 2.350000 3.475000 2.520000 ;
      RECT 3.305000 2.520000 4.535000 2.690000 ;
      RECT 3.645000 2.180000 3.995000 2.350000 ;
      RECT 3.815000 0.255000 4.610000 0.515000 ;
      RECT 3.825000 1.530000 4.155000 1.610000 ;
      RECT 3.825000 1.610000 3.995000 2.180000 ;
      RECT 4.205000 2.090000 4.535000 2.520000 ;
      RECT 4.205000 2.690000 4.535000 2.970000 ;
      RECT 4.280000 0.515000 4.610000 0.850000 ;
      RECT 5.240000 1.820000 6.350000 1.990000 ;
      RECT 5.240000 1.990000 5.570000 2.980000 ;
      RECT 5.260000 1.190000 5.430000 1.300000 ;
      RECT 5.260000 1.300000 5.805000 1.630000 ;
      RECT 5.600000 0.350000 5.975000 0.670000 ;
      RECT 5.600000 0.670000 6.350000 1.130000 ;
      RECT 5.975000 1.130000 6.350000 1.820000 ;
  END
END sky130_fd_sc_ms__dlclkp_4

* File: sky130_fd_sc_ms__mux2i_4.pxi.spice
* Created: Fri Aug 28 17:40:42 2020
* 
x_PM_SKY130_FD_SC_MS__MUX2I_4%A1 N_A1_M1008_g N_A1_M1000_g N_A1_M1005_g
+ N_A1_M1009_g N_A1_M1022_g N_A1_M1011_g N_A1_M1015_g N_A1_M1023_g A1 A1 A1
+ N_A1_c_141_n N_A1_c_136_n PM_SKY130_FD_SC_MS__MUX2I_4%A1
x_PM_SKY130_FD_SC_MS__MUX2I_4%A0 N_A0_M1007_g N_A0_M1001_g N_A0_M1016_g
+ N_A0_M1030_g N_A0_M1031_g N_A0_M1018_g N_A0_c_219_n N_A0_M1034_g N_A0_M1019_g
+ N_A0_c_222_n A0 A0 N_A0_c_224_n PM_SKY130_FD_SC_MS__MUX2I_4%A0
x_PM_SKY130_FD_SC_MS__MUX2I_4%A_1030_268# N_A_1030_268#_M1024_d
+ N_A_1030_268#_M1027_d N_A_1030_268#_M1002_g N_A_1030_268#_c_299_n
+ N_A_1030_268#_M1013_g N_A_1030_268#_M1012_g N_A_1030_268#_c_300_n
+ N_A_1030_268#_M1014_g N_A_1030_268#_M1020_g N_A_1030_268#_M1026_g
+ N_A_1030_268#_M1021_g N_A_1030_268#_M1029_g N_A_1030_268#_c_303_n
+ N_A_1030_268#_c_313_n N_A_1030_268#_c_314_n N_A_1030_268#_c_315_n
+ N_A_1030_268#_c_304_n N_A_1030_268#_c_305_n N_A_1030_268#_c_317_n
+ N_A_1030_268#_c_306_n N_A_1030_268#_c_307_n
+ PM_SKY130_FD_SC_MS__MUX2I_4%A_1030_268#
x_PM_SKY130_FD_SC_MS__MUX2I_4%S N_S_M1003_g N_S_c_429_n N_S_M1010_g N_S_M1004_g
+ N_S_c_431_n N_S_M1017_g N_S_M1006_g N_S_c_433_n N_S_M1025_g N_S_M1032_g
+ N_S_c_435_n N_S_M1028_g N_S_M1027_g N_S_c_437_n N_S_M1024_g N_S_M1033_g S S S
+ S S N_S_c_440_n PM_SKY130_FD_SC_MS__MUX2I_4%S
x_PM_SKY130_FD_SC_MS__MUX2I_4%Y N_Y_M1000_d N_Y_M1005_d N_Y_M1023_d N_Y_M1030_s
+ N_Y_M1034_s N_Y_M1008_s N_Y_M1009_s N_Y_M1015_s N_Y_M1016_s N_Y_M1019_s
+ N_Y_c_543_n N_Y_c_553_n N_Y_c_554_n N_Y_c_544_n N_Y_c_545_n N_Y_c_564_n
+ N_Y_c_646_p N_Y_c_620_p N_Y_c_546_n N_Y_c_572_n N_Y_c_576_n N_Y_c_588_n
+ N_Y_c_547_n N_Y_c_600_n N_Y_c_548_n N_Y_c_549_n N_Y_c_550_n N_Y_c_580_n
+ N_Y_c_582_n N_Y_c_551_n N_Y_c_608_n Y N_Y_c_552_n
+ PM_SKY130_FD_SC_MS__MUX2I_4%Y
x_PM_SKY130_FD_SC_MS__MUX2I_4%A_119_368# N_A_119_368#_M1008_d
+ N_A_119_368#_M1011_d N_A_119_368#_M1002_s N_A_119_368#_M1020_s
+ N_A_119_368#_c_670_n N_A_119_368#_c_664_n N_A_119_368#_c_665_n
+ N_A_119_368#_c_677_n N_A_119_368#_c_666_n N_A_119_368#_c_667_n
+ N_A_119_368#_c_668_n N_A_119_368#_c_669_n
+ PM_SKY130_FD_SC_MS__MUX2I_4%A_119_368#
x_PM_SKY130_FD_SC_MS__MUX2I_4%A_481_368# N_A_481_368#_M1001_d
+ N_A_481_368#_M1018_d N_A_481_368#_M1003_d N_A_481_368#_M1006_d
+ N_A_481_368#_c_728_n N_A_481_368#_c_725_n N_A_481_368#_c_736_n
+ N_A_481_368#_c_742_n N_A_481_368#_c_731_n N_A_481_368#_c_733_n
+ N_A_481_368#_c_772_n N_A_481_368#_c_726_n N_A_481_368#_c_727_n
+ PM_SKY130_FD_SC_MS__MUX2I_4%A_481_368#
x_PM_SKY130_FD_SC_MS__MUX2I_4%VPWR N_VPWR_M1002_d N_VPWR_M1012_d N_VPWR_M1021_d
+ N_VPWR_M1004_s N_VPWR_M1032_s N_VPWR_M1033_s N_VPWR_c_799_n N_VPWR_c_838_n
+ N_VPWR_c_800_n N_VPWR_c_801_n N_VPWR_c_845_n N_VPWR_c_802_n N_VPWR_c_803_n
+ N_VPWR_c_804_n N_VPWR_c_849_n VPWR N_VPWR_c_805_n N_VPWR_c_806_n
+ N_VPWR_c_807_n N_VPWR_c_808_n N_VPWR_c_809_n N_VPWR_c_810_n N_VPWR_c_811_n
+ N_VPWR_c_798_n PM_SKY130_FD_SC_MS__MUX2I_4%VPWR
x_PM_SKY130_FD_SC_MS__MUX2I_4%A_114_85# N_A_114_85#_M1000_s N_A_114_85#_M1022_s
+ N_A_114_85#_M1010_d N_A_114_85#_M1025_d N_A_114_85#_c_936_n
+ N_A_114_85#_c_927_n N_A_114_85#_c_928_n N_A_114_85#_c_943_n
+ N_A_114_85#_c_929_n N_A_114_85#_c_930_n N_A_114_85#_c_931_n
+ N_A_114_85#_c_953_n N_A_114_85#_c_964_n N_A_114_85#_c_932_n
+ N_A_114_85#_c_933_n N_A_114_85#_c_934_n N_A_114_85#_c_958_n
+ N_A_114_85#_c_935_n PM_SKY130_FD_SC_MS__MUX2I_4%A_114_85#
x_PM_SKY130_FD_SC_MS__MUX2I_4%A_475_85# N_A_475_85#_M1007_d N_A_475_85#_M1031_d
+ N_A_475_85#_M1013_d N_A_475_85#_M1026_d N_A_475_85#_c_1036_n
+ N_A_475_85#_c_1037_n N_A_475_85#_c_1038_n N_A_475_85#_c_1039_n
+ N_A_475_85#_c_1040_n PM_SKY130_FD_SC_MS__MUX2I_4%A_475_85#
x_PM_SKY130_FD_SC_MS__MUX2I_4%VGND N_VGND_M1013_s N_VGND_M1014_s N_VGND_M1029_s
+ N_VGND_M1017_s N_VGND_M1028_s N_VGND_c_1080_n N_VGND_c_1081_n N_VGND_c_1082_n
+ N_VGND_c_1083_n N_VGND_c_1084_n N_VGND_c_1085_n N_VGND_c_1086_n VGND
+ N_VGND_c_1087_n N_VGND_c_1088_n N_VGND_c_1089_n N_VGND_c_1090_n
+ N_VGND_c_1091_n N_VGND_c_1092_n N_VGND_c_1093_n N_VGND_c_1094_n
+ PM_SKY130_FD_SC_MS__MUX2I_4%VGND
cc_1 VNB N_A1_M1000_g 0.0277082f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.795
cc_2 VNB N_A1_M1005_g 0.0189276f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.795
cc_3 VNB N_A1_M1022_g 0.0199624f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.795
cc_4 VNB N_A1_M1023_g 0.0202873f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.795
cc_5 VNB N_A1_c_136_n 0.0833979f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.515
cc_6 VNB N_A0_M1007_g 0.0201198f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_7 VNB N_A0_M1030_g 0.0203857f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_8 VNB N_A0_M1031_g 0.0195144f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.795
cc_9 VNB N_A0_c_219_n 0.00940195f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.68
cc_10 VNB N_A0_M1034_g 0.0217715f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.35
cc_11 VNB N_A0_M1019_g 0.00981115f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_12 VNB N_A0_c_222_n 0.0109546f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_13 VNB A0 0.00548856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A0_c_224_n 0.0546126f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.515
cc_15 VNB N_A_1030_268#_c_299_n 0.0200837f $X=-0.19 $Y=-0.245 $X2=0.925
+ $Y2=0.795
cc_16 VNB N_A_1030_268#_c_300_n 0.0177417f $X=-0.19 $Y=-0.245 $X2=1.355
+ $Y2=0.795
cc_17 VNB N_A_1030_268#_M1026_g 0.021673f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_18 VNB N_A_1030_268#_M1029_g 0.021686f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_19 VNB N_A_1030_268#_c_303_n 0.0129921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_1030_268#_c_304_n 0.0205803f $X=-0.19 $Y=-0.245 $X2=1.855
+ $Y2=1.515
cc_21 VNB N_A_1030_268#_c_305_n 0.0249886f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.565
cc_22 VNB N_A_1030_268#_c_306_n 0.00626527f $X=-0.19 $Y=-0.245 $X2=1.72
+ $Y2=1.565
cc_23 VNB N_A_1030_268#_c_307_n 0.0865901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_S_M1003_g 0.00370517f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_25 VNB N_S_c_429_n 0.0168573f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_26 VNB N_S_M1004_g 0.0039416f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.795
cc_27 VNB N_S_c_431_n 0.0171169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_S_M1006_g 0.00394217f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.35
cc_29 VNB N_S_c_433_n 0.0171165f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.795
cc_30 VNB N_S_M1032_g 0.00382473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_S_c_435_n 0.0159706f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_32 VNB N_S_M1027_g 0.00382105f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.795
cc_33 VNB N_S_c_437_n 0.0202827f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_34 VNB N_S_M1033_g 0.00447002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB S 0.0239755f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.515
cc_36 VNB N_S_c_440_n 0.148174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_543_n 0.0247969f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_38 VNB N_Y_c_544_n 0.00448175f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_39 VNB N_Y_c_545_n 0.0110245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Y_c_546_n 0.00326111f $X=-0.19 $Y=-0.245 $X2=1.72 $Y2=1.515
cc_41 VNB N_Y_c_547_n 0.0111441f $X=-0.19 $Y=-0.245 $X2=1.72 $Y2=1.565
cc_42 VNB N_Y_c_548_n 0.00303818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_Y_c_549_n 0.0169696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_Y_c_550_n 0.00124931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_Y_c_551_n 0.0111967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_Y_c_552_n 0.0146497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VPWR_c_798_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_114_85#_c_927_n 0.00702435f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.35
cc_49 VNB N_A_114_85#_c_928_n 0.00401069f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.795
cc_50 VNB N_A_114_85#_c_929_n 0.0491073f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_51 VNB N_A_114_85#_c_930_n 0.0102191f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_52 VNB N_A_114_85#_c_931_n 0.00425516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_114_85#_c_932_n 0.00256522f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_54 VNB N_A_114_85#_c_933_n 0.00241303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_114_85#_c_934_n 0.00312303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_114_85#_c_935_n 0.00256522f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.515
cc_57 VNB N_A_475_85#_c_1036_n 0.0127642f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.68
cc_58 VNB N_A_475_85#_c_1037_n 0.0104048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_475_85#_c_1038_n 0.00907981f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_60 VNB N_A_475_85#_c_1039_n 0.00225985f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_61 VNB N_A_475_85#_c_1040_n 0.0178151f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_62 VNB N_VGND_c_1080_n 0.00967703f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.795
cc_63 VNB N_VGND_c_1081_n 0.0185379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1082_n 0.0183334f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_65 VNB N_VGND_c_1083_n 0.012576f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_66 VNB N_VGND_c_1084_n 0.0079491f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.795
cc_67 VNB N_VGND_c_1085_n 0.0188882f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_68 VNB N_VGND_c_1086_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_69 VNB N_VGND_c_1087_n 0.117093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1088_n 0.0186341f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.515
cc_71 VNB N_VGND_c_1089_n 0.0238f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.565
cc_72 VNB N_VGND_c_1090_n 0.556973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1091_n 0.00477852f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_74 VNB N_VGND_c_1092_n 0.0194475f $X=-0.19 $Y=-0.245 $X2=1.72 $Y2=1.565
cc_75 VNB N_VGND_c_1093_n 0.0169988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1094_n 0.0080786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VPB N_A1_M1008_g 0.0283836f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_78 VPB N_A1_M1009_g 0.0196336f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_79 VPB N_A1_M1011_g 0.0196343f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_80 VPB N_A1_M1015_g 0.0204832f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_81 VPB N_A1_c_141_n 0.00755806f $X=-0.19 $Y=1.66 $X2=1.72 $Y2=1.515
cc_82 VPB N_A1_c_136_n 0.012467f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.515
cc_83 VPB N_A0_M1001_g 0.0213204f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.795
cc_84 VPB N_A0_M1016_g 0.0206799f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.795
cc_85 VPB N_A0_M1018_g 0.0211459f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_86 VPB N_A0_M1019_g 0.0256923f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_87 VPB A0 0.00620664f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A0_c_224_n 0.0108414f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.515
cc_89 VPB N_A_1030_268#_M1002_g 0.0283587f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.35
cc_90 VPB N_A_1030_268#_M1012_g 0.0209385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_1030_268#_M1020_g 0.0218913f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_92 VPB N_A_1030_268#_M1021_g 0.0220296f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=0.795
cc_93 VPB N_A_1030_268#_c_303_n 0.00104f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_1030_268#_c_313_n 0.018179f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.515
cc_95 VPB N_A_1030_268#_c_314_n 0.00329898f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.515
cc_96 VPB N_A_1030_268#_c_315_n 0.00581265f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.515
cc_97 VPB N_A_1030_268#_c_305_n 0.00168332f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.565
cc_98 VPB N_A_1030_268#_c_317_n 0.00195024f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_1030_268#_c_307_n 0.0141991f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_S_M1003_g 0.0221567f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_101 VPB N_S_M1004_g 0.0224675f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.795
cc_102 VPB N_S_M1006_g 0.0224688f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=1.35
cc_103 VPB N_S_M1032_g 0.0224211f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_S_M1027_g 0.0215746f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=0.795
cc_105 VPB N_S_M1033_g 0.0249818f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_Y_c_553_n 0.0157543f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_107 VPB N_Y_c_554_n 0.0339588f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_Y_c_552_n 0.0212775f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_119_368#_c_664_n 0.00192243f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=1.35
cc_110 VPB N_A_119_368#_c_665_n 0.00196551f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.795
cc_111 VPB N_A_119_368#_c_666_n 0.00102348f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.68
cc_112 VPB N_A_119_368#_c_667_n 0.0064993f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_113 VPB N_A_119_368#_c_668_n 0.00160153f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.35
cc_114 VPB N_A_119_368#_c_669_n 0.0248357f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_481_368#_c_725_n 0.0121948f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_116 VPB N_A_481_368#_c_726_n 0.0023101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_481_368#_c_727_n 0.0023101f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.515
cc_118 VPB N_VPWR_c_799_n 0.00404197f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.795
cc_119 VPB N_VPWR_c_800_n 0.00565985f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_120 VPB N_VPWR_c_801_n 0.00899828f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=0.795
cc_121 VPB N_VPWR_c_802_n 0.012691f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_803_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_804_n 0.0517059f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.515
cc_124 VPB N_VPWR_c_805_n 0.156339f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.515
cc_125 VPB N_VPWR_c_806_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_807_n 0.0196495f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.565
cc_127 VPB N_VPWR_c_808_n 0.0186201f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_809_n 0.00612764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_810_n 0.00632182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_811_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_798_n 0.0983636f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 N_A1_M1023_g N_A0_M1007_g 0.0208152f $X=1.87 $Y=0.795 $X2=0 $Y2=0
cc_133 N_A1_M1015_g N_A0_M1001_g 0.0208152f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_134 N_A1_c_141_n N_A0_M1001_g 3.53138e-19 $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_135 N_A1_c_141_n A0 0.0190784f $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_136 N_A1_c_136_n A0 0.00153124f $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_137 N_A1_c_141_n N_A0_c_224_n 3.78435e-19 $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_138 N_A1_c_136_n N_A0_c_224_n 0.0208152f $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_139 N_A1_M1000_g N_Y_c_543_n 0.00159289f $X=0.495 $Y=0.795 $X2=0 $Y2=0
cc_140 N_A1_M1008_g N_Y_c_553_n 8.13654e-19 $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_141 N_A1_M1008_g N_Y_c_554_n 0.00147281f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_142 N_A1_M1000_g N_Y_c_544_n 0.0160051f $X=0.495 $Y=0.795 $X2=0 $Y2=0
cc_143 N_A1_M1005_g N_Y_c_544_n 0.0120585f $X=0.925 $Y=0.795 $X2=0 $Y2=0
cc_144 N_A1_c_141_n N_Y_c_544_n 0.0391613f $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_145 N_A1_c_136_n N_Y_c_544_n 0.00254808f $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_146 N_A1_M1000_g N_Y_c_545_n 2.03611e-19 $X=0.495 $Y=0.795 $X2=0 $Y2=0
cc_147 N_A1_M1008_g N_Y_c_564_n 0.0177137f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_148 N_A1_M1009_g N_Y_c_564_n 0.0142562f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_149 N_A1_c_141_n N_Y_c_564_n 0.0370097f $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_150 N_A1_c_136_n N_Y_c_564_n 4.89709e-19 $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_151 N_A1_M1022_g N_Y_c_546_n 0.0125268f $X=1.355 $Y=0.795 $X2=0 $Y2=0
cc_152 N_A1_M1023_g N_Y_c_546_n 0.0105121f $X=1.87 $Y=0.795 $X2=0 $Y2=0
cc_153 N_A1_c_141_n N_Y_c_546_n 0.0496944f $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_154 N_A1_c_136_n N_Y_c_546_n 0.00452209f $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_155 N_A1_M1011_g N_Y_c_572_n 0.0142562f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A1_M1015_g N_Y_c_572_n 0.0138167f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_157 N_A1_c_141_n N_Y_c_572_n 0.0413875f $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_158 N_A1_c_136_n N_Y_c_572_n 4.90767e-19 $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_159 N_A1_M1022_g N_Y_c_576_n 3.72237e-19 $X=1.355 $Y=0.795 $X2=0 $Y2=0
cc_160 N_A1_M1023_g N_Y_c_576_n 0.00475726f $X=1.87 $Y=0.795 $X2=0 $Y2=0
cc_161 N_A1_c_141_n N_Y_c_550_n 0.0144276f $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_162 N_A1_c_136_n N_Y_c_550_n 0.00249296f $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_163 N_A1_c_141_n N_Y_c_580_n 0.0143992f $X=1.72 $Y=1.515 $X2=0 $Y2=0
cc_164 N_A1_c_136_n N_Y_c_580_n 5.52302e-19 $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_165 N_A1_M1011_g N_Y_c_582_n 4.47651e-19 $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_166 N_A1_M1015_g N_Y_c_582_n 0.0127995f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_167 N_A1_M1022_g N_Y_c_551_n 3.49095e-19 $X=1.355 $Y=0.795 $X2=0 $Y2=0
cc_168 N_A1_M1023_g N_Y_c_551_n 0.00335902f $X=1.87 $Y=0.795 $X2=0 $Y2=0
cc_169 N_A1_M1008_g N_A_119_368#_c_670_n 0.00821143f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_170 N_A1_M1009_g N_A_119_368#_c_670_n 0.00904396f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_171 N_A1_M1011_g N_A_119_368#_c_670_n 5.73047e-19 $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_172 N_A1_M1009_g N_A_119_368#_c_664_n 0.0116345f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_173 N_A1_M1011_g N_A_119_368#_c_664_n 0.0116345f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_174 N_A1_M1008_g N_A_119_368#_c_665_n 0.00696959f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_175 N_A1_M1009_g N_A_119_368#_c_665_n 0.00194226f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_176 N_A1_M1009_g N_A_119_368#_c_677_n 5.74986e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_177 N_A1_M1011_g N_A_119_368#_c_677_n 0.00892729f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_178 N_A1_M1011_g N_A_119_368#_c_668_n 0.00194226f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_179 N_A1_M1015_g N_A_119_368#_c_669_n 0.0140436f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_180 N_A1_M1008_g N_VPWR_c_805_n 0.00517089f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A1_M1009_g N_VPWR_c_805_n 0.00333896f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_182 N_A1_M1011_g N_VPWR_c_805_n 0.00333896f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_183 N_A1_M1015_g N_VPWR_c_805_n 0.00333926f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_184 N_A1_M1008_g N_VPWR_c_798_n 0.00982317f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_185 N_A1_M1009_g N_VPWR_c_798_n 0.00422685f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_186 N_A1_M1011_g N_VPWR_c_798_n 0.00422685f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A1_M1015_g N_VPWR_c_798_n 0.00422893f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A1_M1000_g N_A_114_85#_c_936_n 0.00549852f $X=0.495 $Y=0.795 $X2=0
+ $Y2=0
cc_189 N_A1_M1005_g N_A_114_85#_c_936_n 0.00646199f $X=0.925 $Y=0.795 $X2=0
+ $Y2=0
cc_190 N_A1_M1022_g N_A_114_85#_c_936_n 5.7278e-19 $X=1.355 $Y=0.795 $X2=0 $Y2=0
cc_191 N_A1_M1005_g N_A_114_85#_c_927_n 0.00821552f $X=0.925 $Y=0.795 $X2=0
+ $Y2=0
cc_192 N_A1_M1022_g N_A_114_85#_c_927_n 0.00821552f $X=1.355 $Y=0.795 $X2=0
+ $Y2=0
cc_193 N_A1_M1000_g N_A_114_85#_c_928_n 0.00731971f $X=0.495 $Y=0.795 $X2=0
+ $Y2=0
cc_194 N_A1_M1005_g N_A_114_85#_c_928_n 0.00221614f $X=0.925 $Y=0.795 $X2=0
+ $Y2=0
cc_195 N_A1_M1005_g N_A_114_85#_c_943_n 5.7278e-19 $X=0.925 $Y=0.795 $X2=0 $Y2=0
cc_196 N_A1_M1022_g N_A_114_85#_c_943_n 0.00648141f $X=1.355 $Y=0.795 $X2=0
+ $Y2=0
cc_197 N_A1_M1023_g N_A_114_85#_c_943_n 0.00687051f $X=1.87 $Y=0.795 $X2=0 $Y2=0
cc_198 N_A1_M1023_g N_A_114_85#_c_929_n 0.0111339f $X=1.87 $Y=0.795 $X2=0 $Y2=0
cc_199 N_A1_M1022_g N_A_114_85#_c_933_n 0.00257574f $X=1.355 $Y=0.795 $X2=0
+ $Y2=0
cc_200 N_A1_M1000_g N_VGND_c_1087_n 0.00462669f $X=0.495 $Y=0.795 $X2=0 $Y2=0
cc_201 N_A1_M1005_g N_VGND_c_1087_n 8.82278e-19 $X=0.925 $Y=0.795 $X2=0 $Y2=0
cc_202 N_A1_M1022_g N_VGND_c_1087_n 8.82278e-19 $X=1.355 $Y=0.795 $X2=0 $Y2=0
cc_203 N_A1_M1023_g N_VGND_c_1087_n 8.63546e-19 $X=1.87 $Y=0.795 $X2=0 $Y2=0
cc_204 N_A1_M1000_g N_VGND_c_1090_n 0.00440294f $X=0.495 $Y=0.795 $X2=0 $Y2=0
cc_205 N_A0_M1007_g N_Y_c_576_n 0.00532225f $X=2.3 $Y=0.795 $X2=0 $Y2=0
cc_206 N_A0_M1030_g N_Y_c_576_n 5.45614e-19 $X=2.8 $Y=0.795 $X2=0 $Y2=0
cc_207 N_A0_M1001_g N_Y_c_588_n 0.0144699f $X=2.315 $Y=2.4 $X2=0 $Y2=0
cc_208 N_A0_M1016_g N_Y_c_588_n 0.0117097f $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_209 A0 N_Y_c_588_n 0.0398513f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_210 N_A0_c_224_n N_Y_c_588_n 7.36189e-19 $X=3.395 $Y=1.515 $X2=0 $Y2=0
cc_211 N_A0_M1007_g N_Y_c_547_n 0.0111843f $X=2.3 $Y=0.795 $X2=0 $Y2=0
cc_212 N_A0_M1030_g N_Y_c_547_n 0.0112096f $X=2.8 $Y=0.795 $X2=0 $Y2=0
cc_213 N_A0_M1031_g N_Y_c_547_n 0.0143524f $X=3.275 $Y=0.795 $X2=0 $Y2=0
cc_214 N_A0_c_219_n N_Y_c_547_n 0.00312821f $X=3.63 $Y=1.425 $X2=0 $Y2=0
cc_215 N_A0_M1034_g N_Y_c_547_n 0.0115304f $X=3.705 $Y=0.795 $X2=0 $Y2=0
cc_216 N_A0_c_222_n N_Y_c_547_n 0.00332812f $X=3.762 $Y=1.425 $X2=0 $Y2=0
cc_217 A0 N_Y_c_547_n 0.0763715f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_218 N_A0_c_224_n N_Y_c_547_n 0.00227531f $X=3.395 $Y=1.515 $X2=0 $Y2=0
cc_219 N_A0_M1018_g N_Y_c_600_n 0.0152341f $X=3.305 $Y=2.4 $X2=0 $Y2=0
cc_220 N_A0_M1034_g N_Y_c_549_n 0.00600966f $X=3.705 $Y=0.795 $X2=0 $Y2=0
cc_221 N_A0_c_222_n N_Y_c_549_n 0.00935391f $X=3.762 $Y=1.425 $X2=0 $Y2=0
cc_222 N_A0_M1001_g N_Y_c_582_n 0.0107194f $X=2.315 $Y=2.4 $X2=0 $Y2=0
cc_223 N_A0_M1016_g N_Y_c_582_n 5.87286e-19 $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_224 A0 N_Y_c_582_n 0.00107584f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_225 N_A0_M1007_g N_Y_c_551_n 0.00106304f $X=2.3 $Y=0.795 $X2=0 $Y2=0
cc_226 A0 N_Y_c_551_n 0.00198303f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_227 N_A0_M1018_g N_Y_c_608_n 0.00778103f $X=3.305 $Y=2.4 $X2=0 $Y2=0
cc_228 N_A0_M1019_g N_Y_c_608_n 5.33487e-19 $X=3.805 $Y=2.4 $X2=0 $Y2=0
cc_229 A0 N_Y_c_608_n 0.0233787f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_230 N_A0_c_224_n N_Y_c_608_n 8.23691e-19 $X=3.395 $Y=1.515 $X2=0 $Y2=0
cc_231 N_A0_c_219_n N_Y_c_552_n 0.00443588f $X=3.63 $Y=1.425 $X2=0 $Y2=0
cc_232 N_A0_M1019_g N_Y_c_552_n 0.029069f $X=3.805 $Y=2.4 $X2=0 $Y2=0
cc_233 A0 N_Y_c_552_n 0.015321f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_234 N_A0_c_224_n N_Y_c_552_n 0.00771179f $X=3.395 $Y=1.515 $X2=0 $Y2=0
cc_235 N_A0_M1001_g N_A_119_368#_c_669_n 0.0152753f $X=2.315 $Y=2.4 $X2=0 $Y2=0
cc_236 N_A0_M1016_g N_A_119_368#_c_669_n 0.0106187f $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_237 N_A0_M1018_g N_A_119_368#_c_669_n 0.0106897f $X=3.305 $Y=2.4 $X2=0 $Y2=0
cc_238 N_A0_M1019_g N_A_119_368#_c_669_n 0.0125017f $X=3.805 $Y=2.4 $X2=0 $Y2=0
cc_239 N_A0_M1016_g N_A_481_368#_c_728_n 0.0105718f $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_240 N_A0_M1018_g N_A_481_368#_c_728_n 0.0117357f $X=3.305 $Y=2.4 $X2=0 $Y2=0
cc_241 N_A0_M1019_g N_A_481_368#_c_725_n 0.0124441f $X=3.805 $Y=2.4 $X2=0 $Y2=0
cc_242 N_A0_M1016_g N_A_481_368#_c_731_n 0.00747184f $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_243 N_A0_M1018_g N_A_481_368#_c_731_n 5.3106e-19 $X=3.305 $Y=2.4 $X2=0 $Y2=0
cc_244 N_A0_M1019_g N_A_481_368#_c_733_n 0.0115124f $X=3.805 $Y=2.4 $X2=0 $Y2=0
cc_245 N_A0_M1001_g N_VPWR_c_805_n 0.00333926f $X=2.315 $Y=2.4 $X2=0 $Y2=0
cc_246 N_A0_M1016_g N_VPWR_c_805_n 0.00333926f $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_247 N_A0_M1018_g N_VPWR_c_805_n 0.00333926f $X=3.305 $Y=2.4 $X2=0 $Y2=0
cc_248 N_A0_M1019_g N_VPWR_c_805_n 0.00333926f $X=3.805 $Y=2.4 $X2=0 $Y2=0
cc_249 N_A0_M1001_g N_VPWR_c_798_n 0.00423287f $X=2.315 $Y=2.4 $X2=0 $Y2=0
cc_250 N_A0_M1016_g N_VPWR_c_798_n 0.00422661f $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_251 N_A0_M1018_g N_VPWR_c_798_n 0.00423664f $X=3.305 $Y=2.4 $X2=0 $Y2=0
cc_252 N_A0_M1019_g N_VPWR_c_798_n 0.004274f $X=3.805 $Y=2.4 $X2=0 $Y2=0
cc_253 N_A0_M1007_g N_A_114_85#_c_929_n 0.0108384f $X=2.3 $Y=0.795 $X2=0 $Y2=0
cc_254 N_A0_M1030_g N_A_114_85#_c_929_n 0.0096715f $X=2.8 $Y=0.795 $X2=0 $Y2=0
cc_255 N_A0_M1031_g N_A_114_85#_c_929_n 0.00936954f $X=3.275 $Y=0.795 $X2=0
+ $Y2=0
cc_256 N_A0_M1034_g N_A_114_85#_c_929_n 0.0107358f $X=3.705 $Y=0.795 $X2=0 $Y2=0
cc_257 N_A0_M1030_g N_A_475_85#_c_1036_n 0.0086729f $X=2.8 $Y=0.795 $X2=0 $Y2=0
cc_258 N_A0_M1031_g N_A_475_85#_c_1036_n 0.0086729f $X=3.275 $Y=0.795 $X2=0
+ $Y2=0
cc_259 N_A0_M1034_g N_A_475_85#_c_1036_n 0.0103582f $X=3.705 $Y=0.795 $X2=0
+ $Y2=0
cc_260 N_A0_M1034_g N_A_475_85#_c_1037_n 0.00286364f $X=3.705 $Y=0.795 $X2=0
+ $Y2=0
cc_261 N_A0_M1034_g N_A_475_85#_c_1038_n 3.04488e-19 $X=3.705 $Y=0.795 $X2=0
+ $Y2=0
cc_262 N_A0_M1007_g N_VGND_c_1087_n 8.63546e-19 $X=2.3 $Y=0.795 $X2=0 $Y2=0
cc_263 N_A0_M1030_g N_VGND_c_1087_n 8.63546e-19 $X=2.8 $Y=0.795 $X2=0 $Y2=0
cc_264 N_A0_M1031_g N_VGND_c_1087_n 8.63546e-19 $X=3.275 $Y=0.795 $X2=0 $Y2=0
cc_265 N_A0_M1034_g N_VGND_c_1087_n 8.63546e-19 $X=3.705 $Y=0.795 $X2=0 $Y2=0
cc_266 N_A_1030_268#_M1021_g N_S_M1003_g 0.0433825f $X=6.67 $Y=2.4 $X2=0 $Y2=0
cc_267 N_A_1030_268#_c_303_n N_S_M1003_g 9.43084e-19 $X=6.67 $Y=1.505 $X2=0
+ $Y2=0
cc_268 N_A_1030_268#_c_313_n N_S_M1003_g 0.0114442f $X=9.185 $Y=1.795 $X2=0
+ $Y2=0
cc_269 N_A_1030_268#_c_307_n N_S_M1003_g 0.0117717f $X=6.765 $Y=1.505 $X2=0
+ $Y2=0
cc_270 N_A_1030_268#_M1029_g N_S_c_429_n 0.0249132f $X=6.765 $Y=0.78 $X2=0 $Y2=0
cc_271 N_A_1030_268#_c_313_n N_S_M1004_g 0.01218f $X=9.185 $Y=1.795 $X2=0 $Y2=0
cc_272 N_A_1030_268#_c_313_n N_S_M1006_g 0.0122187f $X=9.185 $Y=1.795 $X2=0
+ $Y2=0
cc_273 N_A_1030_268#_c_313_n N_S_M1032_g 0.0119872f $X=9.185 $Y=1.795 $X2=0
+ $Y2=0
cc_274 N_A_1030_268#_c_314_n N_S_M1032_g 5.42017e-19 $X=9.35 $Y=1.985 $X2=0
+ $Y2=0
cc_275 N_A_1030_268#_c_313_n N_S_M1027_g 0.0132546f $X=9.185 $Y=1.795 $X2=0
+ $Y2=0
cc_276 N_A_1030_268#_c_314_n N_S_M1027_g 0.012805f $X=9.35 $Y=1.985 $X2=0 $Y2=0
cc_277 N_A_1030_268#_c_305_n N_S_M1027_g 5.48653e-19 $X=9.74 $Y=1.71 $X2=0 $Y2=0
cc_278 N_A_1030_268#_c_317_n N_S_M1027_g 0.00237445f $X=9.32 $Y=1.795 $X2=0
+ $Y2=0
cc_279 N_A_1030_268#_c_304_n N_S_c_437_n 0.0120705f $X=9.66 $Y=0.555 $X2=0 $Y2=0
cc_280 N_A_1030_268#_c_305_n N_S_c_437_n 0.00729166f $X=9.74 $Y=1.71 $X2=0 $Y2=0
cc_281 N_A_1030_268#_c_314_n N_S_M1033_g 8.71028e-19 $X=9.35 $Y=1.985 $X2=0
+ $Y2=0
cc_282 N_A_1030_268#_c_315_n N_S_M1033_g 0.0210257f $X=9.655 $Y=1.795 $X2=0
+ $Y2=0
cc_283 N_A_1030_268#_c_305_n N_S_M1033_g 0.00401145f $X=9.74 $Y=1.71 $X2=0 $Y2=0
cc_284 N_A_1030_268#_M1029_g S 0.00347612f $X=6.765 $Y=0.78 $X2=0 $Y2=0
cc_285 N_A_1030_268#_c_303_n S 0.0114918f $X=6.67 $Y=1.505 $X2=0 $Y2=0
cc_286 N_A_1030_268#_c_313_n S 0.155982f $X=9.185 $Y=1.795 $X2=0 $Y2=0
cc_287 N_A_1030_268#_c_315_n S 0.00147587f $X=9.655 $Y=1.795 $X2=0 $Y2=0
cc_288 N_A_1030_268#_c_305_n S 0.0282041f $X=9.74 $Y=1.71 $X2=0 $Y2=0
cc_289 N_A_1030_268#_c_317_n S 0.0227736f $X=9.32 $Y=1.795 $X2=0 $Y2=0
cc_290 N_A_1030_268#_M1029_g N_S_c_440_n 0.0117717f $X=6.765 $Y=0.78 $X2=0 $Y2=0
cc_291 N_A_1030_268#_c_303_n N_S_c_440_n 0.00117342f $X=6.67 $Y=1.505 $X2=0
+ $Y2=0
cc_292 N_A_1030_268#_c_313_n N_S_c_440_n 0.0142231f $X=9.185 $Y=1.795 $X2=0
+ $Y2=0
cc_293 N_A_1030_268#_c_305_n N_S_c_440_n 0.00663373f $X=9.74 $Y=1.71 $X2=0 $Y2=0
cc_294 N_A_1030_268#_c_317_n N_S_c_440_n 0.00260214f $X=9.32 $Y=1.795 $X2=0
+ $Y2=0
cc_295 N_A_1030_268#_c_306_n N_S_c_440_n 0.00555289f $X=9.66 $Y=1.01 $X2=0 $Y2=0
cc_296 N_A_1030_268#_M1002_g N_A_119_368#_c_666_n 0.0106709f $X=5.24 $Y=2.4
+ $X2=0 $Y2=0
cc_297 N_A_1030_268#_M1012_g N_A_119_368#_c_667_n 0.0144936f $X=5.69 $Y=2.4
+ $X2=0 $Y2=0
cc_298 N_A_1030_268#_M1020_g N_A_119_368#_c_667_n 0.0145871f $X=6.14 $Y=2.4
+ $X2=0 $Y2=0
cc_299 N_A_1030_268#_M1021_g N_A_119_368#_c_667_n 0.0024369f $X=6.67 $Y=2.4
+ $X2=0 $Y2=0
cc_300 N_A_1030_268#_M1002_g N_A_119_368#_c_669_n 0.0101684f $X=5.24 $Y=2.4
+ $X2=0 $Y2=0
cc_301 N_A_1030_268#_c_313_n N_A_481_368#_M1003_d 0.00166235f $X=9.185 $Y=1.795
+ $X2=0 $Y2=0
cc_302 N_A_1030_268#_c_313_n N_A_481_368#_M1006_d 0.00166235f $X=9.185 $Y=1.795
+ $X2=0 $Y2=0
cc_303 N_A_1030_268#_M1002_g N_A_481_368#_c_736_n 0.0130461f $X=5.24 $Y=2.4
+ $X2=0 $Y2=0
cc_304 N_A_1030_268#_M1012_g N_A_481_368#_c_736_n 0.0116133f $X=5.69 $Y=2.4
+ $X2=0 $Y2=0
cc_305 N_A_1030_268#_M1020_g N_A_481_368#_c_736_n 0.0121077f $X=6.14 $Y=2.4
+ $X2=0 $Y2=0
cc_306 N_A_1030_268#_M1021_g N_A_481_368#_c_736_n 0.0135408f $X=6.67 $Y=2.4
+ $X2=0 $Y2=0
cc_307 N_A_1030_268#_M1021_g N_A_481_368#_c_726_n 6.10943e-19 $X=6.67 $Y=2.4
+ $X2=0 $Y2=0
cc_308 N_A_1030_268#_c_303_n N_VPWR_M1021_d 3.38829e-19 $X=6.67 $Y=1.505 $X2=0
+ $Y2=0
cc_309 N_A_1030_268#_c_313_n N_VPWR_M1021_d 0.00204228f $X=9.185 $Y=1.795 $X2=0
+ $Y2=0
cc_310 N_A_1030_268#_c_313_n N_VPWR_M1004_s 0.00274955f $X=9.185 $Y=1.795 $X2=0
+ $Y2=0
cc_311 N_A_1030_268#_c_313_n N_VPWR_M1032_s 0.00224297f $X=9.185 $Y=1.795 $X2=0
+ $Y2=0
cc_312 N_A_1030_268#_c_315_n N_VPWR_M1033_s 0.00294424f $X=9.655 $Y=1.795 $X2=0
+ $Y2=0
cc_313 N_A_1030_268#_M1002_g N_VPWR_c_799_n 0.0162865f $X=5.24 $Y=2.4 $X2=0
+ $Y2=0
cc_314 N_A_1030_268#_M1012_g N_VPWR_c_799_n 0.0158206f $X=5.69 $Y=2.4 $X2=0
+ $Y2=0
cc_315 N_A_1030_268#_c_303_n N_VPWR_c_799_n 0.0624716f $X=6.67 $Y=1.505 $X2=0
+ $Y2=0
cc_316 N_A_1030_268#_c_307_n N_VPWR_c_799_n 0.0045073f $X=6.765 $Y=1.505 $X2=0
+ $Y2=0
cc_317 N_A_1030_268#_M1020_g N_VPWR_c_838_n 0.00996518f $X=6.14 $Y=2.4 $X2=0
+ $Y2=0
cc_318 N_A_1030_268#_M1021_g N_VPWR_c_838_n 0.0130312f $X=6.67 $Y=2.4 $X2=0
+ $Y2=0
cc_319 N_A_1030_268#_c_303_n N_VPWR_c_838_n 0.0289854f $X=6.67 $Y=1.505 $X2=0
+ $Y2=0
cc_320 N_A_1030_268#_c_313_n N_VPWR_c_838_n 0.103316f $X=9.185 $Y=1.795 $X2=0
+ $Y2=0
cc_321 N_A_1030_268#_c_307_n N_VPWR_c_838_n 0.00406181f $X=6.765 $Y=1.505 $X2=0
+ $Y2=0
cc_322 N_A_1030_268#_M1020_g N_VPWR_c_800_n 2.09622e-19 $X=6.14 $Y=2.4 $X2=0
+ $Y2=0
cc_323 N_A_1030_268#_M1021_g N_VPWR_c_800_n 0.00668035f $X=6.67 $Y=2.4 $X2=0
+ $Y2=0
cc_324 N_A_1030_268#_c_313_n N_VPWR_c_845_n 0.0171666f $X=9.185 $Y=1.795 $X2=0
+ $Y2=0
cc_325 N_A_1030_268#_c_314_n N_VPWR_c_802_n 0.0178065f $X=9.35 $Y=1.985 $X2=0
+ $Y2=0
cc_326 N_A_1030_268#_c_314_n N_VPWR_c_804_n 0.0240333f $X=9.35 $Y=1.985 $X2=0
+ $Y2=0
cc_327 N_A_1030_268#_c_315_n N_VPWR_c_804_n 0.0114618f $X=9.655 $Y=1.795 $X2=0
+ $Y2=0
cc_328 N_A_1030_268#_M1020_g N_VPWR_c_849_n 0.00578758f $X=6.14 $Y=2.4 $X2=0
+ $Y2=0
cc_329 N_A_1030_268#_M1021_g N_VPWR_c_849_n 8.96733e-19 $X=6.67 $Y=2.4 $X2=0
+ $Y2=0
cc_330 N_A_1030_268#_c_303_n N_VPWR_c_849_n 0.00105934f $X=6.67 $Y=1.505 $X2=0
+ $Y2=0
cc_331 N_A_1030_268#_M1002_g N_VPWR_c_805_n 0.00333926f $X=5.24 $Y=2.4 $X2=0
+ $Y2=0
cc_332 N_A_1030_268#_M1012_g N_VPWR_c_805_n 0.00333926f $X=5.69 $Y=2.4 $X2=0
+ $Y2=0
cc_333 N_A_1030_268#_M1020_g N_VPWR_c_805_n 0.00333926f $X=6.14 $Y=2.4 $X2=0
+ $Y2=0
cc_334 N_A_1030_268#_M1021_g N_VPWR_c_805_n 0.00460063f $X=6.67 $Y=2.4 $X2=0
+ $Y2=0
cc_335 N_A_1030_268#_c_314_n N_VPWR_c_808_n 0.00541659f $X=9.35 $Y=1.985 $X2=0
+ $Y2=0
cc_336 N_A_1030_268#_M1002_g N_VPWR_c_798_n 0.0042782f $X=5.24 $Y=2.4 $X2=0
+ $Y2=0
cc_337 N_A_1030_268#_M1012_g N_VPWR_c_798_n 0.00422687f $X=5.69 $Y=2.4 $X2=0
+ $Y2=0
cc_338 N_A_1030_268#_M1020_g N_VPWR_c_798_n 0.00423447f $X=6.14 $Y=2.4 $X2=0
+ $Y2=0
cc_339 N_A_1030_268#_M1021_g N_VPWR_c_798_n 0.00444006f $X=6.67 $Y=2.4 $X2=0
+ $Y2=0
cc_340 N_A_1030_268#_c_314_n N_VPWR_c_798_n 0.00812781f $X=9.35 $Y=1.985 $X2=0
+ $Y2=0
cc_341 N_A_1030_268#_c_299_n N_A_114_85#_c_930_n 0.00360488f $X=5.315 $Y=1.34
+ $X2=0 $Y2=0
cc_342 N_A_1030_268#_c_300_n N_A_114_85#_c_953_n 0.0123654f $X=5.745 $Y=1.34
+ $X2=0 $Y2=0
cc_343 N_A_1030_268#_M1026_g N_A_114_85#_c_953_n 0.0124889f $X=6.335 $Y=0.78
+ $X2=0 $Y2=0
cc_344 N_A_1030_268#_M1029_g N_A_114_85#_c_953_n 0.0136654f $X=6.765 $Y=0.78
+ $X2=0 $Y2=0
cc_345 N_A_1030_268#_c_303_n N_A_114_85#_c_953_n 0.00330535f $X=6.67 $Y=1.505
+ $X2=0 $Y2=0
cc_346 N_A_1030_268#_c_299_n N_A_114_85#_c_934_n 0.00968689f $X=5.315 $Y=1.34
+ $X2=0 $Y2=0
cc_347 N_A_1030_268#_c_299_n N_A_114_85#_c_958_n 0.00594482f $X=5.315 $Y=1.34
+ $X2=0 $Y2=0
cc_348 N_A_1030_268#_c_300_n N_A_114_85#_c_958_n 0.00224136f $X=5.745 $Y=1.34
+ $X2=0 $Y2=0
cc_349 N_A_1030_268#_M1029_g N_A_114_85#_c_935_n 0.00203198f $X=6.765 $Y=0.78
+ $X2=0 $Y2=0
cc_350 N_A_1030_268#_c_300_n N_A_475_85#_c_1039_n 3.5725e-19 $X=5.745 $Y=1.34
+ $X2=0 $Y2=0
cc_351 N_A_1030_268#_M1026_g N_A_475_85#_c_1039_n 0.00291974f $X=6.335 $Y=0.78
+ $X2=0 $Y2=0
cc_352 N_A_1030_268#_M1029_g N_A_475_85#_c_1039_n 0.00631778f $X=6.765 $Y=0.78
+ $X2=0 $Y2=0
cc_353 N_A_1030_268#_c_303_n N_A_475_85#_c_1039_n 0.00345449f $X=6.67 $Y=1.505
+ $X2=0 $Y2=0
cc_354 N_A_1030_268#_c_307_n N_A_475_85#_c_1039_n 0.00265643f $X=6.765 $Y=1.505
+ $X2=0 $Y2=0
cc_355 N_A_1030_268#_c_299_n N_A_475_85#_c_1040_n 0.0104833f $X=5.315 $Y=1.34
+ $X2=0 $Y2=0
cc_356 N_A_1030_268#_c_300_n N_A_475_85#_c_1040_n 0.00971056f $X=5.745 $Y=1.34
+ $X2=0 $Y2=0
cc_357 N_A_1030_268#_M1026_g N_A_475_85#_c_1040_n 0.00855243f $X=6.335 $Y=0.78
+ $X2=0 $Y2=0
cc_358 N_A_1030_268#_c_303_n N_A_475_85#_c_1040_n 0.104f $X=6.67 $Y=1.505 $X2=0
+ $Y2=0
cc_359 N_A_1030_268#_c_307_n N_A_475_85#_c_1040_n 0.011422f $X=6.765 $Y=1.505
+ $X2=0 $Y2=0
cc_360 N_A_1030_268#_c_299_n N_VGND_c_1080_n 0.00528295f $X=5.315 $Y=1.34 $X2=0
+ $Y2=0
cc_361 N_A_1030_268#_M1026_g N_VGND_c_1081_n 0.00414982f $X=6.335 $Y=0.78 $X2=0
+ $Y2=0
cc_362 N_A_1030_268#_M1029_g N_VGND_c_1081_n 0.00414982f $X=6.765 $Y=0.78 $X2=0
+ $Y2=0
cc_363 N_A_1030_268#_c_304_n N_VGND_c_1084_n 0.0240544f $X=9.66 $Y=0.555 $X2=0
+ $Y2=0
cc_364 N_A_1030_268#_c_299_n N_VGND_c_1088_n 0.00379795f $X=5.315 $Y=1.34 $X2=0
+ $Y2=0
cc_365 N_A_1030_268#_c_300_n N_VGND_c_1088_n 0.00374721f $X=5.745 $Y=1.34 $X2=0
+ $Y2=0
cc_366 N_A_1030_268#_c_304_n N_VGND_c_1089_n 0.0125646f $X=9.66 $Y=0.555 $X2=0
+ $Y2=0
cc_367 N_A_1030_268#_c_299_n N_VGND_c_1090_n 0.00508379f $X=5.315 $Y=1.34 $X2=0
+ $Y2=0
cc_368 N_A_1030_268#_c_300_n N_VGND_c_1090_n 0.00508379f $X=5.745 $Y=1.34 $X2=0
+ $Y2=0
cc_369 N_A_1030_268#_M1026_g N_VGND_c_1090_n 0.00533081f $X=6.335 $Y=0.78 $X2=0
+ $Y2=0
cc_370 N_A_1030_268#_M1029_g N_VGND_c_1090_n 0.00533081f $X=6.765 $Y=0.78 $X2=0
+ $Y2=0
cc_371 N_A_1030_268#_c_304_n N_VGND_c_1090_n 0.0117982f $X=9.66 $Y=0.555 $X2=0
+ $Y2=0
cc_372 N_A_1030_268#_c_300_n N_VGND_c_1092_n 0.0014541f $X=5.745 $Y=1.34 $X2=0
+ $Y2=0
cc_373 N_A_1030_268#_M1026_g N_VGND_c_1092_n 0.00481833f $X=6.335 $Y=0.78 $X2=0
+ $Y2=0
cc_374 N_A_1030_268#_M1029_g N_VGND_c_1093_n 0.00378066f $X=6.765 $Y=0.78 $X2=0
+ $Y2=0
cc_375 N_S_M1003_g N_A_481_368#_c_736_n 0.0097893f $X=7.17 $Y=2.4 $X2=0 $Y2=0
cc_376 N_S_M1004_g N_A_481_368#_c_742_n 0.0100971f $X=7.62 $Y=2.4 $X2=0 $Y2=0
cc_377 N_S_M1006_g N_A_481_368#_c_742_n 0.0100971f $X=8.17 $Y=2.4 $X2=0 $Y2=0
cc_378 N_S_M1003_g N_A_481_368#_c_726_n 0.00753492f $X=7.17 $Y=2.4 $X2=0 $Y2=0
cc_379 N_S_M1004_g N_A_481_368#_c_726_n 0.0077957f $X=7.62 $Y=2.4 $X2=0 $Y2=0
cc_380 N_S_M1006_g N_A_481_368#_c_726_n 3.16734e-19 $X=8.17 $Y=2.4 $X2=0 $Y2=0
cc_381 N_S_M1004_g N_A_481_368#_c_727_n 3.16734e-19 $X=7.62 $Y=2.4 $X2=0 $Y2=0
cc_382 N_S_M1006_g N_A_481_368#_c_727_n 0.0077957f $X=8.17 $Y=2.4 $X2=0 $Y2=0
cc_383 N_S_M1032_g N_A_481_368#_c_727_n 0.00806773f $X=8.62 $Y=2.4 $X2=0 $Y2=0
cc_384 N_S_M1003_g N_VPWR_c_838_n 0.0119096f $X=7.17 $Y=2.4 $X2=0 $Y2=0
cc_385 N_S_M1004_g N_VPWR_c_838_n 0.0122174f $X=7.62 $Y=2.4 $X2=0 $Y2=0
cc_386 N_S_M1006_g N_VPWR_c_838_n 0.0122174f $X=8.17 $Y=2.4 $X2=0 $Y2=0
cc_387 N_S_M1032_g N_VPWR_c_838_n 0.0142256f $X=8.62 $Y=2.4 $X2=0 $Y2=0
cc_388 N_S_M1003_g N_VPWR_c_800_n 0.00194999f $X=7.17 $Y=2.4 $X2=0 $Y2=0
cc_389 N_S_M1004_g N_VPWR_c_801_n 0.00203999f $X=7.62 $Y=2.4 $X2=0 $Y2=0
cc_390 N_S_M1006_g N_VPWR_c_801_n 0.00343717f $X=8.17 $Y=2.4 $X2=0 $Y2=0
cc_391 N_S_M1032_g N_VPWR_c_802_n 0.00848516f $X=8.62 $Y=2.4 $X2=0 $Y2=0
cc_392 N_S_M1027_g N_VPWR_c_802_n 0.00198124f $X=9.125 $Y=2.26 $X2=0 $Y2=0
cc_393 N_S_M1027_g N_VPWR_c_804_n 5.9032e-19 $X=9.125 $Y=2.26 $X2=0 $Y2=0
cc_394 N_S_M1033_g N_VPWR_c_804_n 0.0132893f $X=9.575 $Y=2.26 $X2=0 $Y2=0
cc_395 N_S_M1003_g N_VPWR_c_806_n 0.005209f $X=7.17 $Y=2.4 $X2=0 $Y2=0
cc_396 N_S_M1004_g N_VPWR_c_806_n 0.005209f $X=7.62 $Y=2.4 $X2=0 $Y2=0
cc_397 N_S_M1006_g N_VPWR_c_807_n 0.005209f $X=8.17 $Y=2.4 $X2=0 $Y2=0
cc_398 N_S_M1032_g N_VPWR_c_807_n 0.005209f $X=8.62 $Y=2.4 $X2=0 $Y2=0
cc_399 N_S_M1027_g N_VPWR_c_808_n 0.00465228f $X=9.125 $Y=2.26 $X2=0 $Y2=0
cc_400 N_S_M1033_g N_VPWR_c_808_n 0.00401533f $X=9.575 $Y=2.26 $X2=0 $Y2=0
cc_401 N_S_M1003_g N_VPWR_c_798_n 0.00515319f $X=7.17 $Y=2.4 $X2=0 $Y2=0
cc_402 N_S_M1004_g N_VPWR_c_798_n 0.00515684f $X=7.62 $Y=2.4 $X2=0 $Y2=0
cc_403 N_S_M1006_g N_VPWR_c_798_n 0.00515684f $X=8.17 $Y=2.4 $X2=0 $Y2=0
cc_404 N_S_M1032_g N_VPWR_c_798_n 0.00987399f $X=8.62 $Y=2.4 $X2=0 $Y2=0
cc_405 N_S_M1027_g N_VPWR_c_798_n 0.00555093f $X=9.125 $Y=2.26 $X2=0 $Y2=0
cc_406 N_S_M1033_g N_VPWR_c_798_n 0.00465661f $X=9.575 $Y=2.26 $X2=0 $Y2=0
cc_407 N_S_c_429_n N_A_114_85#_c_953_n 0.0109174f $X=7.355 $Y=1.26 $X2=0 $Y2=0
cc_408 S N_A_114_85#_c_953_n 0.0113104f $X=9.275 $Y=1.21 $X2=0 $Y2=0
cc_409 N_S_c_440_n N_A_114_85#_c_953_n 8.30163e-19 $X=9.375 $Y=1.425 $X2=0 $Y2=0
cc_410 N_S_c_431_n N_A_114_85#_c_964_n 0.0105974f $X=7.785 $Y=1.26 $X2=0 $Y2=0
cc_411 N_S_c_433_n N_A_114_85#_c_964_n 0.0102857f $X=8.445 $Y=1.26 $X2=0 $Y2=0
cc_412 N_S_c_435_n N_A_114_85#_c_964_n 0.00207683f $X=8.875 $Y=1.26 $X2=0 $Y2=0
cc_413 S N_A_114_85#_c_964_n 0.076957f $X=9.275 $Y=1.21 $X2=0 $Y2=0
cc_414 N_S_c_440_n N_A_114_85#_c_964_n 0.0024933f $X=9.375 $Y=1.425 $X2=0 $Y2=0
cc_415 N_S_c_431_n N_A_114_85#_c_932_n 9.07055e-19 $X=7.785 $Y=1.26 $X2=0 $Y2=0
cc_416 N_S_c_433_n N_A_114_85#_c_932_n 0.00741284f $X=8.445 $Y=1.26 $X2=0 $Y2=0
cc_417 N_S_c_435_n N_A_114_85#_c_932_n 0.00507642f $X=8.875 $Y=1.26 $X2=0 $Y2=0
cc_418 N_S_c_429_n N_A_114_85#_c_935_n 0.0108387f $X=7.355 $Y=1.26 $X2=0 $Y2=0
cc_419 N_S_c_431_n N_A_114_85#_c_935_n 0.00867525f $X=7.785 $Y=1.26 $X2=0 $Y2=0
cc_420 N_S_c_433_n N_A_114_85#_c_935_n 9.88713e-19 $X=8.445 $Y=1.26 $X2=0 $Y2=0
cc_421 S N_A_114_85#_c_935_n 0.022955f $X=9.275 $Y=1.21 $X2=0 $Y2=0
cc_422 N_S_c_440_n N_A_114_85#_c_935_n 6.29182e-19 $X=9.375 $Y=1.425 $X2=0 $Y2=0
cc_423 N_S_c_429_n N_A_475_85#_c_1039_n 0.00111481f $X=7.355 $Y=1.26 $X2=0 $Y2=0
cc_424 N_S_c_429_n N_VGND_c_1082_n 0.00412495f $X=7.355 $Y=1.26 $X2=0 $Y2=0
cc_425 N_S_c_431_n N_VGND_c_1082_n 0.00523933f $X=7.785 $Y=1.26 $X2=0 $Y2=0
cc_426 N_S_c_431_n N_VGND_c_1083_n 0.00531504f $X=7.785 $Y=1.26 $X2=0 $Y2=0
cc_427 N_S_c_433_n N_VGND_c_1083_n 0.00384096f $X=8.445 $Y=1.26 $X2=0 $Y2=0
cc_428 N_S_c_435_n N_VGND_c_1084_n 0.00502021f $X=8.875 $Y=1.26 $X2=0 $Y2=0
cc_429 N_S_c_437_n N_VGND_c_1084_n 0.0137136f $X=9.375 $Y=1.26 $X2=0 $Y2=0
cc_430 S N_VGND_c_1084_n 0.025356f $X=9.275 $Y=1.21 $X2=0 $Y2=0
cc_431 N_S_c_440_n N_VGND_c_1084_n 0.00108447f $X=9.375 $Y=1.425 $X2=0 $Y2=0
cc_432 N_S_c_433_n N_VGND_c_1085_n 0.00523933f $X=8.445 $Y=1.26 $X2=0 $Y2=0
cc_433 N_S_c_435_n N_VGND_c_1085_n 0.00523933f $X=8.875 $Y=1.26 $X2=0 $Y2=0
cc_434 N_S_c_437_n N_VGND_c_1089_n 0.00455951f $X=9.375 $Y=1.26 $X2=0 $Y2=0
cc_435 N_S_c_429_n N_VGND_c_1090_n 0.00533081f $X=7.355 $Y=1.26 $X2=0 $Y2=0
cc_436 N_S_c_431_n N_VGND_c_1090_n 0.00533081f $X=7.785 $Y=1.26 $X2=0 $Y2=0
cc_437 N_S_c_433_n N_VGND_c_1090_n 0.00533081f $X=8.445 $Y=1.26 $X2=0 $Y2=0
cc_438 N_S_c_435_n N_VGND_c_1090_n 0.00533081f $X=8.875 $Y=1.26 $X2=0 $Y2=0
cc_439 N_S_c_437_n N_VGND_c_1090_n 0.00447788f $X=9.375 $Y=1.26 $X2=0 $Y2=0
cc_440 N_S_c_429_n N_VGND_c_1093_n 0.00339091f $X=7.355 $Y=1.26 $X2=0 $Y2=0
cc_441 N_Y_c_564_n N_A_119_368#_M1008_d 0.00314376f $X=1.095 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_442 N_Y_c_572_n N_A_119_368#_M1011_d 0.00314376f $X=1.915 $Y=2.035 $X2=0
+ $Y2=0
cc_443 N_Y_c_564_n N_A_119_368#_c_670_n 0.0170259f $X=1.095 $Y=2.035 $X2=0 $Y2=0
cc_444 N_Y_M1009_s N_A_119_368#_c_664_n 0.00165831f $X=1.045 $Y=1.84 $X2=0 $Y2=0
cc_445 N_Y_c_620_p N_A_119_368#_c_664_n 0.0118736f $X=1.18 $Y=2.57 $X2=0 $Y2=0
cc_446 N_Y_c_554_n N_A_119_368#_c_665_n 0.00345031f $X=0.28 $Y=2.4 $X2=0 $Y2=0
cc_447 N_Y_c_572_n N_A_119_368#_c_677_n 0.0148589f $X=1.915 $Y=2.035 $X2=0 $Y2=0
cc_448 N_Y_M1015_s N_A_119_368#_c_669_n 0.00176461f $X=1.945 $Y=1.84 $X2=0 $Y2=0
cc_449 N_Y_M1016_s N_A_119_368#_c_669_n 0.00219516f $X=2.895 $Y=1.84 $X2=0 $Y2=0
cc_450 N_Y_M1019_s N_A_119_368#_c_669_n 0.00335745f $X=3.895 $Y=1.84 $X2=0 $Y2=0
cc_451 N_Y_c_582_n N_A_119_368#_c_669_n 0.0159805f $X=2.08 $Y=2.035 $X2=0 $Y2=0
cc_452 N_Y_c_588_n N_A_481_368#_M1001_d 0.00404817f $X=2.915 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_453 N_Y_c_600_n N_A_481_368#_M1018_d 0.00156114f $X=3.485 $Y=2.035 $X2=0
+ $Y2=0
cc_454 N_Y_c_552_n N_A_481_368#_M1018_d 0.00334856f $X=4.08 $Y=1.965 $X2=0 $Y2=0
cc_455 N_Y_M1016_s N_A_481_368#_c_728_n 0.00428212f $X=2.895 $Y=1.84 $X2=0 $Y2=0
cc_456 N_Y_c_588_n N_A_481_368#_c_728_n 0.00464895f $X=2.915 $Y=2.035 $X2=0
+ $Y2=0
cc_457 N_Y_c_600_n N_A_481_368#_c_728_n 0.00464895f $X=3.485 $Y=2.035 $X2=0
+ $Y2=0
cc_458 N_Y_c_608_n N_A_481_368#_c_728_n 0.0182896f $X=3.08 $Y=2.035 $X2=0 $Y2=0
cc_459 N_Y_M1019_s N_A_481_368#_c_725_n 0.00706967f $X=3.895 $Y=1.84 $X2=0 $Y2=0
cc_460 N_Y_c_552_n N_A_481_368#_c_725_n 0.0290322f $X=4.08 $Y=1.965 $X2=0 $Y2=0
cc_461 N_Y_c_588_n N_A_481_368#_c_731_n 0.0175034f $X=2.915 $Y=2.035 $X2=0 $Y2=0
cc_462 N_Y_c_600_n N_A_481_368#_c_733_n 0.00255808f $X=3.485 $Y=2.035 $X2=0
+ $Y2=0
cc_463 N_Y_c_552_n N_A_481_368#_c_733_n 0.0172271f $X=4.08 $Y=1.965 $X2=0 $Y2=0
cc_464 N_Y_c_552_n N_VPWR_c_799_n 0.0282236f $X=4.08 $Y=1.965 $X2=0 $Y2=0
cc_465 N_Y_c_554_n N_VPWR_c_805_n 0.011066f $X=0.28 $Y=2.4 $X2=0 $Y2=0
cc_466 N_Y_c_554_n N_VPWR_c_798_n 0.00915947f $X=0.28 $Y=2.4 $X2=0 $Y2=0
cc_467 N_Y_c_544_n N_A_114_85#_M1000_s 0.00176461f $X=1.055 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_468 N_Y_c_546_n N_A_114_85#_M1022_s 0.00266828f $X=1.92 $Y=1.095 $X2=0 $Y2=0
cc_469 N_Y_c_544_n N_A_114_85#_c_936_n 0.0168694f $X=1.055 $Y=1.095 $X2=0 $Y2=0
cc_470 N_Y_c_544_n N_A_114_85#_c_927_n 0.00390898f $X=1.055 $Y=1.095 $X2=0 $Y2=0
cc_471 N_Y_c_646_p N_A_114_85#_c_927_n 0.0127861f $X=1.14 $Y=0.82 $X2=0 $Y2=0
cc_472 N_Y_c_546_n N_A_114_85#_c_927_n 0.00390898f $X=1.92 $Y=1.095 $X2=0 $Y2=0
cc_473 N_Y_c_543_n N_A_114_85#_c_928_n 0.00153535f $X=0.28 $Y=0.57 $X2=0 $Y2=0
cc_474 N_Y_c_546_n N_A_114_85#_c_943_n 0.021615f $X=1.92 $Y=1.095 $X2=0 $Y2=0
cc_475 N_Y_c_576_n N_A_114_85#_c_943_n 0.0178172f $X=2.085 $Y=0.68 $X2=0 $Y2=0
cc_476 N_Y_c_546_n N_A_114_85#_c_929_n 0.00402835f $X=1.92 $Y=1.095 $X2=0 $Y2=0
cc_477 N_Y_c_576_n N_A_114_85#_c_929_n 0.0203275f $X=2.085 $Y=0.68 $X2=0 $Y2=0
cc_478 N_Y_c_547_n N_A_114_85#_c_929_n 0.00433239f $X=3.915 $Y=1.057 $X2=0 $Y2=0
cc_479 N_Y_c_547_n N_A_475_85#_M1007_d 0.00254333f $X=3.915 $Y=1.057 $X2=-0.19
+ $Y2=-0.245
cc_480 N_Y_c_547_n N_A_475_85#_M1031_d 0.00178895f $X=3.915 $Y=1.057 $X2=0 $Y2=0
cc_481 N_Y_M1030_s N_A_475_85#_c_1036_n 0.00425377f $X=2.875 $Y=0.425 $X2=0
+ $Y2=0
cc_482 N_Y_M1034_s N_A_475_85#_c_1036_n 0.00566273f $X=3.78 $Y=0.425 $X2=0 $Y2=0
cc_483 N_Y_c_547_n N_A_475_85#_c_1036_n 0.0827364f $X=3.915 $Y=1.057 $X2=0 $Y2=0
cc_484 N_Y_c_548_n N_A_475_85#_c_1036_n 0.013893f $X=4 $Y=1.18 $X2=0 $Y2=0
cc_485 N_Y_c_548_n N_A_475_85#_c_1037_n 0.00545207f $X=4 $Y=1.18 $X2=0 $Y2=0
cc_486 N_Y_c_548_n N_A_475_85#_c_1038_n 0.0159284f $X=4 $Y=1.18 $X2=0 $Y2=0
cc_487 N_Y_c_543_n N_VGND_c_1087_n 0.00905681f $X=0.28 $Y=0.57 $X2=0 $Y2=0
cc_488 N_Y_c_543_n N_VGND_c_1090_n 0.00884938f $X=0.28 $Y=0.57 $X2=0 $Y2=0
cc_489 N_A_119_368#_c_669_n N_A_481_368#_M1001_d 0.00208352f $X=5.3 $Y=2.902
+ $X2=-0.19 $Y2=1.66
cc_490 N_A_119_368#_c_669_n N_A_481_368#_M1018_d 0.00218982f $X=5.3 $Y=2.902
+ $X2=0 $Y2=0
cc_491 N_A_119_368#_c_669_n N_A_481_368#_c_728_n 0.035128f $X=5.3 $Y=2.902 $X2=0
+ $Y2=0
cc_492 N_A_119_368#_c_669_n N_A_481_368#_c_725_n 0.0791409f $X=5.3 $Y=2.902
+ $X2=0 $Y2=0
cc_493 N_A_119_368#_M1002_s N_A_481_368#_c_736_n 0.00329181f $X=5.33 $Y=1.84
+ $X2=0 $Y2=0
cc_494 N_A_119_368#_M1020_s N_A_481_368#_c_736_n 0.00497992f $X=6.23 $Y=1.84
+ $X2=0 $Y2=0
cc_495 N_A_119_368#_c_666_n N_A_481_368#_c_736_n 0.0676826f $X=5.472 $Y=2.902
+ $X2=0 $Y2=0
cc_496 N_A_119_368#_c_669_n N_A_481_368#_c_736_n 0.00500376f $X=5.3 $Y=2.902
+ $X2=0 $Y2=0
cc_497 N_A_119_368#_c_669_n N_A_481_368#_c_731_n 0.0164435f $X=5.3 $Y=2.902
+ $X2=0 $Y2=0
cc_498 N_A_119_368#_c_669_n N_A_481_368#_c_733_n 0.0171805f $X=5.3 $Y=2.902
+ $X2=0 $Y2=0
cc_499 N_A_119_368#_c_669_n N_A_481_368#_c_772_n 0.009546f $X=5.3 $Y=2.902 $X2=0
+ $Y2=0
cc_500 N_A_119_368#_c_669_n N_VPWR_M1002_d 0.00777801f $X=5.3 $Y=2.902 $X2=-0.19
+ $Y2=1.66
cc_501 N_A_119_368#_c_667_n N_VPWR_M1012_d 0.00169896f $X=6.38 $Y=2.815 $X2=0
+ $Y2=0
cc_502 N_A_119_368#_M1002_s N_VPWR_c_799_n 0.00319704f $X=5.33 $Y=1.84 $X2=0
+ $Y2=0
cc_503 N_A_119_368#_M1020_s N_VPWR_c_838_n 0.0057207f $X=6.23 $Y=1.84 $X2=0
+ $Y2=0
cc_504 N_A_119_368#_c_667_n N_VPWR_c_800_n 0.0181992f $X=6.38 $Y=2.815 $X2=0
+ $Y2=0
cc_505 N_A_119_368#_c_664_n N_VPWR_c_805_n 0.0357927f $X=1.465 $Y=2.99 $X2=0
+ $Y2=0
cc_506 N_A_119_368#_c_665_n N_VPWR_c_805_n 0.0234458f $X=0.895 $Y=2.99 $X2=0
+ $Y2=0
cc_507 N_A_119_368#_c_668_n N_VPWR_c_805_n 0.0178163f $X=1.59 $Y=2.99 $X2=0
+ $Y2=0
cc_508 N_A_119_368#_c_669_n N_VPWR_c_805_n 0.311874f $X=5.3 $Y=2.902 $X2=0 $Y2=0
cc_509 N_A_119_368#_c_664_n N_VPWR_c_798_n 0.0200586f $X=1.465 $Y=2.99 $X2=0
+ $Y2=0
cc_510 N_A_119_368#_c_665_n N_VPWR_c_798_n 0.0125551f $X=0.895 $Y=2.99 $X2=0
+ $Y2=0
cc_511 N_A_119_368#_c_668_n N_VPWR_c_798_n 0.00958215f $X=1.59 $Y=2.99 $X2=0
+ $Y2=0
cc_512 N_A_119_368#_c_669_n N_VPWR_c_798_n 0.176347f $X=5.3 $Y=2.902 $X2=0 $Y2=0
cc_513 N_A_481_368#_c_725_n N_VPWR_M1002_d 0.0163552f $X=4.96 $Y=2.65 $X2=-0.19
+ $Y2=1.66
cc_514 N_A_481_368#_c_772_n N_VPWR_M1002_d 0.0101853f $X=5.045 $Y=2.475
+ $X2=-0.19 $Y2=1.66
cc_515 N_A_481_368#_c_736_n N_VPWR_M1012_d 0.00329181f $X=7.23 $Y=2.475 $X2=0
+ $Y2=0
cc_516 N_A_481_368#_c_736_n N_VPWR_M1021_d 0.00432071f $X=7.23 $Y=2.475 $X2=0
+ $Y2=0
cc_517 N_A_481_368#_c_742_n N_VPWR_M1004_s 0.00548861f $X=8.23 $Y=2.475 $X2=0
+ $Y2=0
cc_518 N_A_481_368#_c_725_n N_VPWR_c_799_n 0.022342f $X=4.96 $Y=2.65 $X2=0 $Y2=0
cc_519 N_A_481_368#_c_736_n N_VPWR_c_799_n 0.11666f $X=7.23 $Y=2.475 $X2=0 $Y2=0
cc_520 N_A_481_368#_c_772_n N_VPWR_c_799_n 0.0107875f $X=5.045 $Y=2.475 $X2=0
+ $Y2=0
cc_521 N_A_481_368#_M1003_d N_VPWR_c_838_n 0.00320283f $X=7.26 $Y=1.84 $X2=0
+ $Y2=0
cc_522 N_A_481_368#_M1006_d N_VPWR_c_838_n 0.00320283f $X=8.26 $Y=1.84 $X2=0
+ $Y2=0
cc_523 N_A_481_368#_c_742_n N_VPWR_c_838_n 0.0388605f $X=8.23 $Y=2.475 $X2=0
+ $Y2=0
cc_524 N_A_481_368#_c_726_n N_VPWR_c_838_n 0.0169819f $X=7.395 $Y=2.475 $X2=0
+ $Y2=0
cc_525 N_A_481_368#_c_727_n N_VPWR_c_838_n 0.0169819f $X=8.395 $Y=2.475 $X2=0
+ $Y2=0
cc_526 N_A_481_368#_c_736_n N_VPWR_c_800_n 0.0183185f $X=7.23 $Y=2.475 $X2=0
+ $Y2=0
cc_527 N_A_481_368#_c_726_n N_VPWR_c_800_n 0.0101711f $X=7.395 $Y=2.475 $X2=0
+ $Y2=0
cc_528 N_A_481_368#_c_742_n N_VPWR_c_801_n 0.0202465f $X=8.23 $Y=2.475 $X2=0
+ $Y2=0
cc_529 N_A_481_368#_c_726_n N_VPWR_c_801_n 0.0101711f $X=7.395 $Y=2.475 $X2=0
+ $Y2=0
cc_530 N_A_481_368#_c_727_n N_VPWR_c_801_n 0.0101711f $X=8.395 $Y=2.475 $X2=0
+ $Y2=0
cc_531 N_A_481_368#_c_727_n N_VPWR_c_802_n 0.0144801f $X=8.395 $Y=2.475 $X2=0
+ $Y2=0
cc_532 N_A_481_368#_c_726_n N_VPWR_c_806_n 0.0143153f $X=7.395 $Y=2.475 $X2=0
+ $Y2=0
cc_533 N_A_481_368#_c_727_n N_VPWR_c_807_n 0.0143153f $X=8.395 $Y=2.475 $X2=0
+ $Y2=0
cc_534 N_A_481_368#_c_736_n N_VPWR_c_798_n 0.0138002f $X=7.23 $Y=2.475 $X2=0
+ $Y2=0
cc_535 N_A_481_368#_c_742_n N_VPWR_c_798_n 0.0115311f $X=8.23 $Y=2.475 $X2=0
+ $Y2=0
cc_536 N_A_481_368#_c_726_n N_VPWR_c_798_n 0.0117766f $X=7.395 $Y=2.475 $X2=0
+ $Y2=0
cc_537 N_A_481_368#_c_727_n N_VPWR_c_798_n 0.0117766f $X=8.395 $Y=2.475 $X2=0
+ $Y2=0
cc_538 N_VPWR_c_799_n N_A_475_85#_c_1040_n 0.0183764f $X=5.89 $Y=2.03 $X2=0
+ $Y2=0
cc_539 N_A_114_85#_c_953_n N_A_475_85#_M1013_d 0.00245099f $X=7.405 $Y=0.665
+ $X2=0 $Y2=0
cc_540 N_A_114_85#_c_958_n N_A_475_85#_M1013_d 0.0031412f $X=5.525 $Y=0.705
+ $X2=0 $Y2=0
cc_541 N_A_114_85#_c_953_n N_A_475_85#_M1026_d 0.00437807f $X=7.405 $Y=0.665
+ $X2=0 $Y2=0
cc_542 N_A_114_85#_c_929_n N_A_475_85#_c_1036_n 0.127231f $X=4.595 $Y=0.34 $X2=0
+ $Y2=0
cc_543 N_A_114_85#_c_930_n N_A_475_85#_c_1036_n 0.00545212f $X=4.68 $Y=0.66
+ $X2=0 $Y2=0
cc_544 N_A_114_85#_c_931_n N_A_475_85#_c_1036_n 0.00983825f $X=4.765 $Y=0.745
+ $X2=0 $Y2=0
cc_545 N_A_114_85#_c_931_n N_A_475_85#_c_1037_n 0.00545212f $X=4.765 $Y=0.745
+ $X2=0 $Y2=0
cc_546 N_A_114_85#_c_953_n N_A_475_85#_c_1039_n 0.0158362f $X=7.405 $Y=0.665
+ $X2=0 $Y2=0
cc_547 N_A_114_85#_c_929_n N_A_475_85#_c_1040_n 0.00546133f $X=4.595 $Y=0.34
+ $X2=0 $Y2=0
cc_548 N_A_114_85#_c_931_n N_A_475_85#_c_1040_n 0.0141608f $X=4.765 $Y=0.745
+ $X2=0 $Y2=0
cc_549 N_A_114_85#_c_953_n N_A_475_85#_c_1040_n 0.0362502f $X=7.405 $Y=0.665
+ $X2=0 $Y2=0
cc_550 N_A_114_85#_c_934_n N_A_475_85#_c_1040_n 0.0466221f $X=5.355 $Y=0.705
+ $X2=0 $Y2=0
cc_551 N_A_114_85#_c_934_n N_VGND_M1013_s 0.00857417f $X=5.355 $Y=0.705
+ $X2=-0.19 $Y2=-0.245
cc_552 N_A_114_85#_c_953_n N_VGND_M1014_s 0.00784108f $X=7.405 $Y=0.665 $X2=0
+ $Y2=0
cc_553 N_A_114_85#_c_953_n N_VGND_M1029_s 0.0130597f $X=7.405 $Y=0.665 $X2=0
+ $Y2=0
cc_554 N_A_114_85#_c_964_n N_VGND_M1017_s 0.00938892f $X=8.495 $Y=0.925 $X2=0
+ $Y2=0
cc_555 N_A_114_85#_c_929_n N_VGND_c_1080_n 0.0145007f $X=4.595 $Y=0.34 $X2=0
+ $Y2=0
cc_556 N_A_114_85#_c_930_n N_VGND_c_1080_n 0.00491053f $X=4.68 $Y=0.66 $X2=0
+ $Y2=0
cc_557 N_A_114_85#_c_934_n N_VGND_c_1080_n 0.0190193f $X=5.355 $Y=0.705 $X2=0
+ $Y2=0
cc_558 N_A_114_85#_c_953_n N_VGND_c_1081_n 0.0114147f $X=7.405 $Y=0.665 $X2=0
+ $Y2=0
cc_559 N_A_114_85#_c_953_n N_VGND_c_1082_n 0.0029521f $X=7.405 $Y=0.665 $X2=0
+ $Y2=0
cc_560 N_A_114_85#_c_935_n N_VGND_c_1082_n 0.012388f $X=7.57 $Y=0.555 $X2=0
+ $Y2=0
cc_561 N_A_114_85#_c_964_n N_VGND_c_1083_n 0.0275613f $X=8.495 $Y=0.925 $X2=0
+ $Y2=0
cc_562 N_A_114_85#_c_932_n N_VGND_c_1083_n 0.0102004f $X=8.66 $Y=0.555 $X2=0
+ $Y2=0
cc_563 N_A_114_85#_c_935_n N_VGND_c_1083_n 0.0102004f $X=7.57 $Y=0.555 $X2=0
+ $Y2=0
cc_564 N_A_114_85#_c_932_n N_VGND_c_1084_n 0.017638f $X=8.66 $Y=0.555 $X2=0
+ $Y2=0
cc_565 N_A_114_85#_c_932_n N_VGND_c_1085_n 0.012388f $X=8.66 $Y=0.555 $X2=0
+ $Y2=0
cc_566 N_A_114_85#_c_927_n N_VGND_c_1087_n 0.0340834f $X=1.405 $Y=0.34 $X2=0
+ $Y2=0
cc_567 N_A_114_85#_c_928_n N_VGND_c_1087_n 0.023391f $X=0.875 $Y=0.34 $X2=0
+ $Y2=0
cc_568 N_A_114_85#_c_929_n N_VGND_c_1087_n 0.196212f $X=4.595 $Y=0.34 $X2=0
+ $Y2=0
cc_569 N_A_114_85#_c_933_n N_VGND_c_1087_n 0.023391f $X=1.57 $Y=0.34 $X2=0 $Y2=0
cc_570 N_A_114_85#_c_934_n N_VGND_c_1087_n 0.00287846f $X=5.355 $Y=0.705 $X2=0
+ $Y2=0
cc_571 N_A_114_85#_c_934_n N_VGND_c_1088_n 0.00226196f $X=5.355 $Y=0.705 $X2=0
+ $Y2=0
cc_572 N_A_114_85#_c_958_n N_VGND_c_1088_n 0.00869542f $X=5.525 $Y=0.705 $X2=0
+ $Y2=0
cc_573 N_A_114_85#_c_927_n N_VGND_c_1090_n 0.0199188f $X=1.405 $Y=0.34 $X2=0
+ $Y2=0
cc_574 N_A_114_85#_c_928_n N_VGND_c_1090_n 0.0127797f $X=0.875 $Y=0.34 $X2=0
+ $Y2=0
cc_575 N_A_114_85#_c_929_n N_VGND_c_1090_n 0.114102f $X=4.595 $Y=0.34 $X2=0
+ $Y2=0
cc_576 N_A_114_85#_c_953_n N_VGND_c_1090_n 0.0288944f $X=7.405 $Y=0.665 $X2=0
+ $Y2=0
cc_577 N_A_114_85#_c_964_n N_VGND_c_1090_n 0.0123991f $X=8.495 $Y=0.925 $X2=0
+ $Y2=0
cc_578 N_A_114_85#_c_932_n N_VGND_c_1090_n 0.0117351f $X=8.66 $Y=0.555 $X2=0
+ $Y2=0
cc_579 N_A_114_85#_c_933_n N_VGND_c_1090_n 0.0127797f $X=1.57 $Y=0.34 $X2=0
+ $Y2=0
cc_580 N_A_114_85#_c_934_n N_VGND_c_1090_n 0.010536f $X=5.355 $Y=0.705 $X2=0
+ $Y2=0
cc_581 N_A_114_85#_c_958_n N_VGND_c_1090_n 0.0154249f $X=5.525 $Y=0.705 $X2=0
+ $Y2=0
cc_582 N_A_114_85#_c_935_n N_VGND_c_1090_n 0.0117351f $X=7.57 $Y=0.555 $X2=0
+ $Y2=0
cc_583 N_A_114_85#_c_953_n N_VGND_c_1092_n 0.024515f $X=7.405 $Y=0.665 $X2=0
+ $Y2=0
cc_584 N_A_114_85#_c_953_n N_VGND_c_1093_n 0.0244835f $X=7.405 $Y=0.665 $X2=0
+ $Y2=0
cc_585 N_A_114_85#_c_935_n N_VGND_c_1093_n 0.00151601f $X=7.57 $Y=0.555 $X2=0
+ $Y2=0
cc_586 N_A_475_85#_c_1040_n N_VGND_M1013_s 0.0110424f $X=6.385 $Y=1.045
+ $X2=-0.19 $Y2=-0.245
cc_587 N_A_475_85#_c_1040_n N_VGND_M1014_s 0.00651909f $X=6.385 $Y=1.045 $X2=0
+ $Y2=0

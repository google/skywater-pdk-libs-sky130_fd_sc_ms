* File: sky130_fd_sc_ms__and2_1.pxi.spice
* Created: Fri Aug 28 17:10:38 2020
* 
x_PM_SKY130_FD_SC_MS__AND2_1%A N_A_c_46_n N_A_M1004_g N_A_M1000_g N_A_c_49_n A A
+ N_A_c_51_n PM_SKY130_FD_SC_MS__AND2_1%A
x_PM_SKY130_FD_SC_MS__AND2_1%B N_B_M1003_g N_B_M1001_g B N_B_c_80_n N_B_c_81_n
+ PM_SKY130_FD_SC_MS__AND2_1%B
x_PM_SKY130_FD_SC_MS__AND2_1%A_56_136# N_A_56_136#_M1004_s N_A_56_136#_M1000_d
+ N_A_56_136#_M1002_g N_A_56_136#_M1005_g N_A_56_136#_c_123_n
+ N_A_56_136#_c_129_n N_A_56_136#_c_130_n N_A_56_136#_c_131_n
+ N_A_56_136#_c_132_n N_A_56_136#_c_133_n N_A_56_136#_c_134_n
+ N_A_56_136#_c_124_n N_A_56_136#_c_125_n N_A_56_136#_c_126_n
+ PM_SKY130_FD_SC_MS__AND2_1%A_56_136#
x_PM_SKY130_FD_SC_MS__AND2_1%VPWR N_VPWR_M1000_s N_VPWR_M1001_d N_VPWR_c_191_n
+ N_VPWR_c_192_n N_VPWR_c_193_n N_VPWR_c_194_n N_VPWR_c_195_n N_VPWR_c_196_n
+ VPWR N_VPWR_c_197_n N_VPWR_c_190_n PM_SKY130_FD_SC_MS__AND2_1%VPWR
x_PM_SKY130_FD_SC_MS__AND2_1%X N_X_M1005_d N_X_M1002_d N_X_c_220_n X X X
+ N_X_c_221_n X PM_SKY130_FD_SC_MS__AND2_1%X
x_PM_SKY130_FD_SC_MS__AND2_1%VGND N_VGND_M1003_d N_VGND_c_243_n N_VGND_c_244_n
+ N_VGND_c_245_n VGND N_VGND_c_246_n N_VGND_c_247_n
+ PM_SKY130_FD_SC_MS__AND2_1%VGND
cc_1 VNB N_A_c_46_n 0.02449f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.57
cc_2 VNB N_A_M1004_g 0.0120472f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1
cc_3 VNB N_A_M1000_g 0.00665438f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=2.54
cc_4 VNB N_A_c_49_n 0.0204322f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.545
cc_5 VNB A 0.0358286f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_6 VNB N_A_c_51_n 0.0544958f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.405
cc_7 VNB B 0.00237204f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=2.54
cc_8 VNB N_B_c_80_n 0.0272161f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.395
cc_9 VNB N_B_c_81_n 0.0182698f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_10 VNB N_A_56_136#_c_123_n 0.0335551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_56_136#_c_124_n 0.00556882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_56_136#_c_125_n 0.0290474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_56_136#_c_126_n 0.0216407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_VPWR_c_190_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_X_c_220_n 0.0367857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_X_c_221_n 0.02259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_243_n 0.0186268f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1
cc_18 VNB N_VGND_c_244_n 0.037648f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=2.54
cc_19 VNB N_VGND_c_245_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_246_n 0.0224545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_247_n 0.173493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VPB N_A_M1000_g 0.0457628f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=2.54
cc_23 VPB N_B_M1001_g 0.038269f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1
cc_24 VPB B 0.00138105f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=2.54
cc_25 VPB N_B_c_80_n 0.00562806f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=1.395
cc_26 VPB N_A_56_136#_M1002_g 0.0265323f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=2.54
cc_27 VPB N_A_56_136#_c_123_n 0.0101637f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_28 VPB N_A_56_136#_c_129_n 0.00257779f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.405
cc_29 VPB N_A_56_136#_c_130_n 0.0141715f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.405
cc_30 VPB N_A_56_136#_c_131_n 0.00382904f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_31 VPB N_A_56_136#_c_132_n 0.00402361f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.462
cc_32 VPB N_A_56_136#_c_133_n 0.0018089f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_33 VPB N_A_56_136#_c_134_n 0.00948496f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_A_56_136#_c_124_n 4.76351e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_A_56_136#_c_125_n 0.00665765f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_191_n 0.0394681f $X=-0.19 $Y=1.66 $X2=0.745 $Y2=2.54
cc_37 VPB N_VPWR_c_192_n 0.0063584f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.47
cc_38 VPB N_VPWR_c_193_n 0.013281f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_194_n 0.00622357f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=0.405
cc_40 VPB N_VPWR_c_195_n 0.0195482f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=0.405
cc_41 VPB N_VPWR_c_196_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.462
cc_42 VPB N_VPWR_c_197_n 0.0205542f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_190_n 0.0642224f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB X 0.0535168f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=0.47
cc_45 VPB N_X_c_221_n 0.0090547f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 N_A_M1000_g N_B_M1001_g 0.027694f $X=0.745 $Y=2.54 $X2=0 $Y2=0
cc_47 N_A_M1004_g B 0.00151136f $X=0.64 $Y=1 $X2=0 $Y2=0
cc_48 N_A_c_49_n B 0.00112834f $X=0.7 $Y=1.545 $X2=0 $Y2=0
cc_49 N_A_M1004_g N_B_c_80_n 0.00137655f $X=0.64 $Y=1 $X2=0 $Y2=0
cc_50 N_A_c_49_n N_B_c_80_n 0.0150816f $X=0.7 $Y=1.545 $X2=0 $Y2=0
cc_51 N_A_c_46_n N_B_c_81_n 0.00298419f $X=0.64 $Y=0.57 $X2=0 $Y2=0
cc_52 N_A_M1004_g N_B_c_81_n 0.0210976f $X=0.64 $Y=1 $X2=0 $Y2=0
cc_53 A N_B_c_81_n 0.00194518f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_54 N_A_M1004_g N_A_56_136#_c_123_n 0.014365f $X=0.64 $Y=1 $X2=0 $Y2=0
cc_55 N_A_M1000_g N_A_56_136#_c_123_n 0.0108936f $X=0.745 $Y=2.54 $X2=0 $Y2=0
cc_56 N_A_c_49_n N_A_56_136#_c_123_n 0.00648097f $X=0.7 $Y=1.545 $X2=0 $Y2=0
cc_57 A N_A_56_136#_c_123_n 0.0255901f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_58 N_A_c_51_n N_A_56_136#_c_123_n 0.00172729f $X=0.61 $Y=0.405 $X2=0 $Y2=0
cc_59 N_A_M1000_g N_A_56_136#_c_129_n 0.0233387f $X=0.745 $Y=2.54 $X2=0 $Y2=0
cc_60 N_A_c_49_n N_A_56_136#_c_129_n 0.00232067f $X=0.7 $Y=1.545 $X2=0 $Y2=0
cc_61 N_A_M1000_g N_A_56_136#_c_131_n 0.00416461f $X=0.745 $Y=2.54 $X2=0 $Y2=0
cc_62 N_A_M1000_g N_VPWR_c_191_n 0.0171812f $X=0.745 $Y=2.54 $X2=0 $Y2=0
cc_63 N_A_M1000_g N_VPWR_c_195_n 0.00460063f $X=0.745 $Y=2.54 $X2=0 $Y2=0
cc_64 N_A_M1000_g N_VPWR_c_190_n 0.00909121f $X=0.745 $Y=2.54 $X2=0 $Y2=0
cc_65 N_A_c_46_n N_VGND_c_243_n 0.00157877f $X=0.64 $Y=0.57 $X2=0 $Y2=0
cc_66 A N_VGND_c_243_n 0.015731f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_67 A N_VGND_c_244_n 0.0478766f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_68 N_A_c_51_n N_VGND_c_244_n 0.0116176f $X=0.61 $Y=0.405 $X2=0 $Y2=0
cc_69 N_A_c_46_n N_VGND_c_247_n 0.00487856f $X=0.64 $Y=0.57 $X2=0 $Y2=0
cc_70 A N_VGND_c_247_n 0.0249126f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_71 N_A_c_51_n N_VGND_c_247_n 0.0101636f $X=0.61 $Y=0.405 $X2=0 $Y2=0
cc_72 N_B_M1001_g N_A_56_136#_M1002_g 0.0304724f $X=1.245 $Y=2.54 $X2=0 $Y2=0
cc_73 B N_A_56_136#_c_123_n 0.0171072f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_74 N_B_c_80_n N_A_56_136#_c_123_n 5.35461e-19 $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_75 N_B_c_81_n N_A_56_136#_c_123_n 0.00171729f $X=1.24 $Y=1.35 $X2=0 $Y2=0
cc_76 N_B_M1001_g N_A_56_136#_c_131_n 0.0171513f $X=1.245 $Y=2.54 $X2=0 $Y2=0
cc_77 N_B_M1001_g N_A_56_136#_c_132_n 0.0133513f $X=1.245 $Y=2.54 $X2=0 $Y2=0
cc_78 B N_A_56_136#_c_132_n 0.0164847f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_79 N_B_c_80_n N_A_56_136#_c_132_n 4.86414e-19 $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_80 N_B_M1001_g N_A_56_136#_c_133_n 0.00333279f $X=1.245 $Y=2.54 $X2=0 $Y2=0
cc_81 N_B_M1001_g N_A_56_136#_c_134_n 0.00313133f $X=1.245 $Y=2.54 $X2=0 $Y2=0
cc_82 B N_A_56_136#_c_134_n 0.00937184f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_83 N_B_c_80_n N_A_56_136#_c_134_n 6.23375e-19 $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_84 B N_A_56_136#_c_124_n 0.0258883f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_85 N_B_c_80_n N_A_56_136#_c_124_n 0.00201866f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_86 B N_A_56_136#_c_125_n 3.66423e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_87 N_B_c_80_n N_A_56_136#_c_125_n 0.0174253f $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_88 B N_A_56_136#_c_126_n 0.00358991f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_89 N_B_c_81_n N_A_56_136#_c_126_n 0.0187211f $X=1.24 $Y=1.35 $X2=0 $Y2=0
cc_90 N_B_M1001_g N_VPWR_c_191_n 7.20741e-19 $X=1.245 $Y=2.54 $X2=0 $Y2=0
cc_91 N_B_M1001_g N_VPWR_c_192_n 0.00703269f $X=1.245 $Y=2.54 $X2=0 $Y2=0
cc_92 N_B_M1001_g N_VPWR_c_195_n 0.00520371f $X=1.245 $Y=2.54 $X2=0 $Y2=0
cc_93 N_B_M1001_g N_VPWR_c_190_n 0.00983436f $X=1.245 $Y=2.54 $X2=0 $Y2=0
cc_94 N_B_c_81_n N_X_c_220_n 8.72408e-19 $X=1.24 $Y=1.35 $X2=0 $Y2=0
cc_95 B A_143_136# 8.67896e-19 $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_96 B N_VGND_M1003_d 0.00152312f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_97 B N_VGND_c_243_n 0.00546541f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_98 N_B_c_80_n N_VGND_c_243_n 3.3155e-19 $X=1.24 $Y=1.515 $X2=0 $Y2=0
cc_99 N_B_c_81_n N_VGND_c_243_n 0.0043444f $X=1.24 $Y=1.35 $X2=0 $Y2=0
cc_100 N_B_c_81_n N_VGND_c_244_n 0.00428744f $X=1.24 $Y=1.35 $X2=0 $Y2=0
cc_101 N_B_c_81_n N_VGND_c_247_n 0.00476395f $X=1.24 $Y=1.35 $X2=0 $Y2=0
cc_102 N_A_56_136#_c_132_n N_VPWR_M1001_d 0.00734463f $X=1.58 $Y=1.935 $X2=0
+ $Y2=0
cc_103 N_A_56_136#_c_129_n N_VPWR_c_191_n 0.00494571f $X=0.855 $Y=1.935 $X2=0
+ $Y2=0
cc_104 N_A_56_136#_c_130_n N_VPWR_c_191_n 0.0219579f $X=0.59 $Y=1.935 $X2=0
+ $Y2=0
cc_105 N_A_56_136#_c_131_n N_VPWR_c_191_n 0.0320857f $X=1.02 $Y=2.265 $X2=0
+ $Y2=0
cc_106 N_A_56_136#_M1002_g N_VPWR_c_192_n 0.0180494f $X=1.78 $Y=2.4 $X2=0 $Y2=0
cc_107 N_A_56_136#_c_131_n N_VPWR_c_192_n 0.0275873f $X=1.02 $Y=2.265 $X2=0
+ $Y2=0
cc_108 N_A_56_136#_c_132_n N_VPWR_c_192_n 0.0221548f $X=1.58 $Y=1.935 $X2=0
+ $Y2=0
cc_109 N_A_56_136#_c_131_n N_VPWR_c_195_n 0.0158202f $X=1.02 $Y=2.265 $X2=0
+ $Y2=0
cc_110 N_A_56_136#_M1002_g N_VPWR_c_197_n 0.00460063f $X=1.78 $Y=2.4 $X2=0 $Y2=0
cc_111 N_A_56_136#_M1002_g N_VPWR_c_190_n 0.00912634f $X=1.78 $Y=2.4 $X2=0 $Y2=0
cc_112 N_A_56_136#_c_131_n N_VPWR_c_190_n 0.0121193f $X=1.02 $Y=2.265 $X2=0
+ $Y2=0
cc_113 N_A_56_136#_c_124_n N_X_c_220_n 0.00842104f $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_114 N_A_56_136#_c_125_n N_X_c_220_n 0.00240804f $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_115 N_A_56_136#_c_126_n N_X_c_220_n 0.0106952f $X=1.81 $Y=1.35 $X2=0 $Y2=0
cc_116 N_A_56_136#_M1002_g X 8.78237e-19 $X=1.78 $Y=2.4 $X2=0 $Y2=0
cc_117 N_A_56_136#_c_124_n X 0.00419007f $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_118 N_A_56_136#_c_125_n X 0.00123968f $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_119 N_A_56_136#_M1002_g N_X_c_221_n 0.0023318f $X=1.78 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A_56_136#_c_133_n N_X_c_221_n 0.00456328f $X=1.665 $Y=1.85 $X2=0 $Y2=0
cc_121 N_A_56_136#_c_124_n N_X_c_221_n 0.0251162f $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_122 N_A_56_136#_c_125_n N_X_c_221_n 0.00231223f $X=1.81 $Y=1.515 $X2=0 $Y2=0
cc_123 N_A_56_136#_c_126_n N_X_c_221_n 0.00348686f $X=1.81 $Y=1.35 $X2=0 $Y2=0
cc_124 N_A_56_136#_c_124_n N_VGND_c_243_n 0.00429544f $X=1.81 $Y=1.515 $X2=0
+ $Y2=0
cc_125 N_A_56_136#_c_125_n N_VGND_c_243_n 4.5946e-19 $X=1.81 $Y=1.515 $X2=0
+ $Y2=0
cc_126 N_A_56_136#_c_126_n N_VGND_c_243_n 0.00769141f $X=1.81 $Y=1.35 $X2=0
+ $Y2=0
cc_127 N_A_56_136#_c_126_n N_VGND_c_246_n 0.0046731f $X=1.81 $Y=1.35 $X2=0 $Y2=0
cc_128 N_A_56_136#_c_126_n N_VGND_c_247_n 0.00505379f $X=1.81 $Y=1.35 $X2=0
+ $Y2=0
cc_129 N_VPWR_c_192_n X 0.0267513f $X=1.555 $Y=2.355 $X2=0 $Y2=0
cc_130 N_VPWR_c_197_n X 0.017536f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_131 N_VPWR_c_190_n X 0.0145148f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_132 N_X_c_220_n N_VGND_c_243_n 0.0226294f $X=2.005 $Y=0.645 $X2=0 $Y2=0
cc_133 N_X_c_220_n N_VGND_c_246_n 0.0141483f $X=2.005 $Y=0.645 $X2=0 $Y2=0
cc_134 N_X_c_220_n N_VGND_c_247_n 0.0161522f $X=2.005 $Y=0.645 $X2=0 $Y2=0

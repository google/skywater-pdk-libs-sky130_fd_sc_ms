* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdlclkp_4 CLK GATE SCE VGND VNB VPB VPWR GCLK
X0 a_324_79# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_634_74# a_354_105# a_744_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X2 a_119_143# a_354_105# a_634_74# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X3 VPWR CLK a_1292_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X4 VPWR a_634_74# a_792_48# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 GCLK a_1292_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X6 VGND a_1292_368# GCLK VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_119_143# a_324_79# a_634_74# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X8 VGND a_324_79# a_354_105# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 VPWR SCE a_119_395# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X10 GCLK a_1292_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_119_143# GATE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X12 a_119_395# GATE a_119_143# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X13 a_1292_368# a_792_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X14 GCLK a_1292_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 GCLK a_1292_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 VGND SCE a_119_143# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X17 VPWR a_324_79# a_354_105# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X18 a_324_79# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X19 a_744_74# a_792_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X20 VGND a_1292_368# GCLK VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 a_1292_74# a_792_48# a_1292_368# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 VPWR a_1292_368# GCLK VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X23 VPWR a_1292_368# GCLK VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X24 a_634_74# a_324_79# a_788_455# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X25 VGND CLK a_1292_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 VGND a_634_74# a_792_48# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 a_788_455# a_792_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
.ends

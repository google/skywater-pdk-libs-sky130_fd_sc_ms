* File: sky130_fd_sc_ms__a31oi_1.pxi.spice
* Created: Fri Aug 28 17:07:23 2020
* 
x_PM_SKY130_FD_SC_MS__A31OI_1%A3 N_A3_M1007_g N_A3_c_48_n N_A3_M1006_g
+ N_A3_c_49_n N_A3_c_50_n A3 PM_SKY130_FD_SC_MS__A31OI_1%A3
x_PM_SKY130_FD_SC_MS__A31OI_1%A2 N_A2_M1004_g N_A2_M1000_g A2 A2 N_A2_c_77_n
+ N_A2_c_78_n PM_SKY130_FD_SC_MS__A31OI_1%A2
x_PM_SKY130_FD_SC_MS__A31OI_1%A1 N_A1_M1003_g N_A1_M1001_g A1 N_A1_c_109_n
+ N_A1_c_110_n PM_SKY130_FD_SC_MS__A31OI_1%A1
x_PM_SKY130_FD_SC_MS__A31OI_1%B1 N_B1_c_142_n N_B1_M1005_g N_B1_M1002_g
+ N_B1_c_144_n B1 B1 N_B1_c_146_n PM_SKY130_FD_SC_MS__A31OI_1%B1
x_PM_SKY130_FD_SC_MS__A31OI_1%VPWR N_VPWR_M1007_s N_VPWR_M1000_d N_VPWR_c_168_n
+ N_VPWR_c_169_n N_VPWR_c_170_n N_VPWR_c_171_n N_VPWR_c_172_n VPWR
+ N_VPWR_c_173_n N_VPWR_c_167_n PM_SKY130_FD_SC_MS__A31OI_1%VPWR
x_PM_SKY130_FD_SC_MS__A31OI_1%A_139_368# N_A_139_368#_M1007_d
+ N_A_139_368#_M1001_d N_A_139_368#_c_204_n N_A_139_368#_c_202_n
+ N_A_139_368#_c_208_n N_A_139_368#_c_212_n N_A_139_368#_c_203_n
+ PM_SKY130_FD_SC_MS__A31OI_1%A_139_368#
x_PM_SKY130_FD_SC_MS__A31OI_1%Y N_Y_M1003_d N_Y_M1002_d N_Y_c_232_n N_Y_c_233_n
+ N_Y_c_234_n N_Y_c_237_n N_Y_c_244_n N_Y_c_235_n Y Y Y N_Y_c_238_n
+ PM_SKY130_FD_SC_MS__A31OI_1%Y
x_PM_SKY130_FD_SC_MS__A31OI_1%VGND N_VGND_M1006_s N_VGND_M1005_d N_VGND_c_290_n
+ N_VGND_c_291_n N_VGND_c_292_n N_VGND_c_293_n N_VGND_c_294_n VGND
+ N_VGND_c_295_n N_VGND_c_296_n PM_SKY130_FD_SC_MS__A31OI_1%VGND
cc_1 VNB N_A3_M1007_g 0.00872128f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.4
cc_2 VNB N_A3_c_48_n 0.0193012f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.22
cc_3 VNB N_A3_c_49_n 0.0564055f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.385
cc_4 VNB N_A3_c_50_n 0.0153482f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.385
cc_5 VNB A3 0.00839483f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_A2_M1000_g 0.00688704f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.74
cc_7 VNB A2 0.00485115f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.385
cc_8 VNB N_A2_c_77_n 0.0306907f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_9 VNB N_A2_c_78_n 0.0178222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A1_M1001_g 0.00711974f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.74
cc_11 VNB A1 0.00362176f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.385
cc_12 VNB N_A1_c_109_n 0.0326396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_c_110_n 0.0197655f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_14 VNB N_B1_c_142_n 0.0223503f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.55
cc_15 VNB N_B1_M1002_g 0.00957504f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.74
cc_16 VNB N_B1_c_144_n 0.0109684f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.385
cc_17 VNB B1 0.030738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_c_146_n 0.0528453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_167_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_232_n 0.00369921f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.385
cc_21 VNB N_Y_c_233_n 0.00534354f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.385
cc_22 VNB N_Y_c_234_n 6.00478e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_23 VNB N_Y_c_235_n 0.00306185f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_24 VNB N_VGND_c_290_n 0.0125358f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.74
cc_25 VNB N_VGND_c_291_n 0.0377251f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.385
cc_26 VNB N_VGND_c_292_n 0.0344107f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_27 VNB N_VGND_c_293_n 0.0450666f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_28 VNB N_VGND_c_294_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_295_n 0.0123263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_296_n 0.19226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VPB N_A3_M1007_g 0.0276199f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=2.4
cc_32 VPB N_A2_M1000_g 0.0239457f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=0.74
cc_33 VPB N_A1_M1001_g 0.0245785f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=0.74
cc_34 VPB N_B1_M1002_g 0.0297445f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=0.74
cc_35 VPB N_VPWR_c_168_n 0.0125099f $X=-0.19 $Y=1.66 $X2=0.65 $Y2=0.74
cc_36 VPB N_VPWR_c_169_n 0.0594561f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.385
cc_37 VPB N_VPWR_c_170_n 0.00986613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_171_n 0.0212406f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_172_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.385
cc_40 VPB N_VPWR_c_173_n 0.0384912f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_167_n 0.0626314f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A_139_368#_c_202_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.62 $Y2=1.385
cc_43 VPB N_A_139_368#_c_203_n 0.00275675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_Y_c_232_n 5.66269e-19 $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.385
cc_45 VPB N_Y_c_237_n 0.0339211f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_Y_c_238_n 0.0544117f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 N_A3_M1007_g N_A2_M1000_g 0.0243055f $X=0.605 $Y=2.4 $X2=0 $Y2=0
cc_48 N_A3_c_48_n A2 8.19586e-19 $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_49 N_A3_c_50_n N_A2_c_77_n 0.0337327f $X=0.62 $Y=1.385 $X2=0 $Y2=0
cc_50 N_A3_c_48_n N_A2_c_78_n 0.0337327f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_51 N_A3_M1007_g N_VPWR_c_169_n 0.0353476f $X=0.605 $Y=2.4 $X2=0 $Y2=0
cc_52 N_A3_c_49_n N_VPWR_c_169_n 0.00245403f $X=0.515 $Y=1.385 $X2=0 $Y2=0
cc_53 A3 N_VPWR_c_169_n 0.0198099f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_54 N_A3_M1007_g N_VPWR_c_171_n 0.005209f $X=0.605 $Y=2.4 $X2=0 $Y2=0
cc_55 N_A3_M1007_g N_VPWR_c_167_n 0.00986643f $X=0.605 $Y=2.4 $X2=0 $Y2=0
cc_56 N_A3_M1007_g N_A_139_368#_c_204_n 0.00259983f $X=0.605 $Y=2.4 $X2=0 $Y2=0
cc_57 N_A3_M1007_g N_A_139_368#_c_202_n 0.0100782f $X=0.605 $Y=2.4 $X2=0 $Y2=0
cc_58 N_A3_M1007_g N_Y_c_232_n 0.00844195f $X=0.605 $Y=2.4 $X2=0 $Y2=0
cc_59 N_A3_c_48_n N_Y_c_232_n 0.0191301f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_60 N_A3_c_50_n N_Y_c_232_n 0.009604f $X=0.62 $Y=1.385 $X2=0 $Y2=0
cc_61 A3 N_Y_c_232_n 0.0265523f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_62 N_A3_c_48_n N_Y_c_234_n 0.00539306f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_63 N_A3_M1007_g N_Y_c_244_n 0.0105307f $X=0.605 $Y=2.4 $X2=0 $Y2=0
cc_64 N_A3_c_48_n N_VGND_c_291_n 0.0179036f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_65 N_A3_c_49_n N_VGND_c_291_n 0.00232901f $X=0.515 $Y=1.385 $X2=0 $Y2=0
cc_66 A3 N_VGND_c_291_n 0.0288422f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_67 N_A3_c_48_n N_VGND_c_293_n 0.00348163f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_68 N_A3_c_48_n N_VGND_c_296_n 0.00546242f $X=0.65 $Y=1.22 $X2=0 $Y2=0
cc_69 N_A2_M1000_g N_A1_M1001_g 0.0346013f $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_70 A2 A1 0.0242365f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_71 N_A2_c_77_n A1 4.06701e-19 $X=1.13 $Y=1.385 $X2=0 $Y2=0
cc_72 N_A2_c_77_n N_A1_c_109_n 0.0175474f $X=1.13 $Y=1.385 $X2=0 $Y2=0
cc_73 A2 N_A1_c_110_n 0.00825186f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_74 N_A2_c_78_n N_A1_c_110_n 0.0265239f $X=1.13 $Y=1.22 $X2=0 $Y2=0
cc_75 N_A2_M1000_g N_VPWR_c_170_n 0.00929294f $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_76 N_A2_M1000_g N_VPWR_c_171_n 0.005209f $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_77 N_A2_M1000_g N_VPWR_c_167_n 0.00984243f $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_78 N_A2_M1000_g N_A_139_368#_c_204_n 8.84614e-19 $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_79 N_A2_M1000_g N_A_139_368#_c_202_n 0.0114144f $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_80 N_A2_M1000_g N_A_139_368#_c_208_n 0.0138062f $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_81 N_A2_M1000_g N_A_139_368#_c_203_n 8.71334e-19 $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_82 A2 N_Y_c_232_n 0.0554335f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_83 N_A2_c_78_n N_Y_c_232_n 0.0133143f $X=1.13 $Y=1.22 $X2=0 $Y2=0
cc_84 A2 N_Y_c_233_n 0.013653f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_85 N_A2_c_78_n N_Y_c_233_n 0.0109398f $X=1.13 $Y=1.22 $X2=0 $Y2=0
cc_86 N_A2_M1000_g N_Y_c_237_n 0.0124777f $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_87 A2 N_Y_c_237_n 0.0272275f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_88 N_A2_c_77_n N_Y_c_237_n 0.00105742f $X=1.13 $Y=1.385 $X2=0 $Y2=0
cc_89 N_A2_c_78_n N_VGND_c_293_n 0.00291649f $X=1.13 $Y=1.22 $X2=0 $Y2=0
cc_90 N_A2_c_78_n N_VGND_c_296_n 0.00359136f $X=1.13 $Y=1.22 $X2=0 $Y2=0
cc_91 A2 A_223_74# 0.00606047f $X=1.115 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_92 N_A1_c_110_n N_B1_c_142_n 0.0233894f $X=1.7 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_93 N_A1_M1001_g N_B1_M1002_g 0.0220564f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_94 A1 N_B1_c_144_n 3.68035e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_95 N_A1_c_109_n N_B1_c_144_n 0.0174972f $X=1.7 $Y=1.385 $X2=0 $Y2=0
cc_96 A1 B1 0.029889f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_97 N_A1_c_109_n B1 0.00216087f $X=1.7 $Y=1.385 $X2=0 $Y2=0
cc_98 N_A1_M1001_g N_VPWR_c_170_n 0.0092232f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_99 N_A1_M1001_g N_VPWR_c_173_n 0.005209f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_100 N_A1_M1001_g N_VPWR_c_167_n 0.00984923f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_101 N_A1_M1001_g N_A_139_368#_c_202_n 8.65962e-19 $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_102 N_A1_M1001_g N_A_139_368#_c_208_n 0.0138062f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_103 N_A1_M1001_g N_A_139_368#_c_212_n 8.84614e-19 $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_104 N_A1_M1001_g N_A_139_368#_c_203_n 0.0115643f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_105 A1 N_Y_c_233_n 0.00420927f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_106 N_A1_c_110_n N_Y_c_233_n 0.0131896f $X=1.7 $Y=1.22 $X2=0 $Y2=0
cc_107 N_A1_M1001_g N_Y_c_237_n 0.0127774f $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_108 A1 N_Y_c_237_n 0.024317f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_109 N_A1_c_109_n N_Y_c_237_n 0.00103683f $X=1.7 $Y=1.385 $X2=0 $Y2=0
cc_110 A1 N_Y_c_235_n 0.0111615f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_111 N_A1_c_109_n N_Y_c_235_n 9.02374e-19 $X=1.7 $Y=1.385 $X2=0 $Y2=0
cc_112 N_A1_M1001_g N_Y_c_238_n 7.64188e-19 $X=1.695 $Y=2.4 $X2=0 $Y2=0
cc_113 N_A1_c_110_n N_VGND_c_292_n 7.24629e-19 $X=1.7 $Y=1.22 $X2=0 $Y2=0
cc_114 N_A1_c_110_n N_VGND_c_293_n 0.00291649f $X=1.7 $Y=1.22 $X2=0 $Y2=0
cc_115 N_A1_c_110_n N_VGND_c_296_n 0.00361625f $X=1.7 $Y=1.22 $X2=0 $Y2=0
cc_116 N_B1_M1002_g N_VPWR_c_173_n 0.005209f $X=2.195 $Y=2.4 $X2=0 $Y2=0
cc_117 N_B1_M1002_g N_VPWR_c_167_n 0.00988155f $X=2.195 $Y=2.4 $X2=0 $Y2=0
cc_118 N_B1_M1002_g N_Y_c_237_n 0.0167358f $X=2.195 $Y=2.4 $X2=0 $Y2=0
cc_119 B1 N_Y_c_237_n 0.0579042f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_120 N_B1_c_146_n N_Y_c_237_n 0.0109287f $X=2.61 $Y=1.385 $X2=0 $Y2=0
cc_121 N_B1_c_142_n N_Y_c_235_n 0.00110948f $X=2.18 $Y=1.22 $X2=0 $Y2=0
cc_122 B1 N_Y_c_235_n 7.29591e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_123 N_B1_M1002_g N_Y_c_238_n 0.0156855f $X=2.195 $Y=2.4 $X2=0 $Y2=0
cc_124 N_B1_c_142_n N_VGND_c_292_n 0.0124734f $X=2.18 $Y=1.22 $X2=0 $Y2=0
cc_125 N_B1_c_144_n N_VGND_c_292_n 0.00199599f $X=2.195 $Y=1.385 $X2=0 $Y2=0
cc_126 B1 N_VGND_c_292_n 0.0259403f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_127 N_B1_c_142_n N_VGND_c_293_n 0.00383152f $X=2.18 $Y=1.22 $X2=0 $Y2=0
cc_128 N_B1_c_142_n N_VGND_c_296_n 0.00758792f $X=2.18 $Y=1.22 $X2=0 $Y2=0
cc_129 N_VPWR_c_169_n N_A_139_368#_c_204_n 0.0118923f $X=0.29 $Y=1.985 $X2=0
+ $Y2=0
cc_130 N_VPWR_c_169_n N_A_139_368#_c_202_n 0.0494853f $X=0.29 $Y=1.985 $X2=0
+ $Y2=0
cc_131 N_VPWR_c_170_n N_A_139_368#_c_202_n 0.0383002f $X=1.37 $Y=2.485 $X2=0
+ $Y2=0
cc_132 N_VPWR_c_171_n N_A_139_368#_c_202_n 0.0144436f $X=1.205 $Y=3.33 $X2=0
+ $Y2=0
cc_133 N_VPWR_c_167_n N_A_139_368#_c_202_n 0.0118287f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_134 N_VPWR_M1000_d N_A_139_368#_c_208_n 0.0085164f $X=1.145 $Y=1.84 $X2=0
+ $Y2=0
cc_135 N_VPWR_c_170_n N_A_139_368#_c_208_n 0.0266856f $X=1.37 $Y=2.485 $X2=0
+ $Y2=0
cc_136 N_VPWR_c_170_n N_A_139_368#_c_203_n 0.0369618f $X=1.37 $Y=2.485 $X2=0
+ $Y2=0
cc_137 N_VPWR_c_173_n N_A_139_368#_c_203_n 0.014549f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_138 N_VPWR_c_167_n N_A_139_368#_c_203_n 0.0119743f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_139 N_VPWR_M1000_d N_Y_c_237_n 0.00391561f $X=1.145 $Y=1.84 $X2=0 $Y2=0
cc_140 N_VPWR_c_169_n N_Y_c_244_n 0.00579824f $X=0.29 $Y=1.985 $X2=0 $Y2=0
cc_141 N_VPWR_c_173_n N_Y_c_238_n 0.0221345f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_142 N_VPWR_c_167_n N_Y_c_238_n 0.0182529f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_143 N_A_139_368#_M1007_d N_Y_c_237_n 0.00119058f $X=0.695 $Y=1.84 $X2=0 $Y2=0
cc_144 N_A_139_368#_M1001_d N_Y_c_237_n 0.00218982f $X=1.785 $Y=1.84 $X2=0 $Y2=0
cc_145 N_A_139_368#_c_204_n N_Y_c_237_n 0.0114002f $X=0.83 $Y=2.23 $X2=0 $Y2=0
cc_146 N_A_139_368#_c_208_n N_Y_c_237_n 0.0453975f $X=1.755 $Y=2.145 $X2=0 $Y2=0
cc_147 N_A_139_368#_c_212_n N_Y_c_237_n 0.019003f $X=1.92 $Y=2.23 $X2=0 $Y2=0
cc_148 N_A_139_368#_M1007_d N_Y_c_244_n 4.75848e-19 $X=0.695 $Y=1.84 $X2=0 $Y2=0
cc_149 N_A_139_368#_c_204_n N_Y_c_244_n 0.00637416f $X=0.83 $Y=2.23 $X2=0 $Y2=0
cc_150 N_A_139_368#_c_203_n N_Y_c_238_n 0.0307786f $X=1.92 $Y=2.825 $X2=0 $Y2=0
cc_151 N_Y_c_232_n N_VGND_c_291_n 0.0362227f $X=0.71 $Y=1.72 $X2=0 $Y2=0
cc_152 N_Y_c_234_n N_VGND_c_291_n 0.0140387f $X=0.795 $Y=0.435 $X2=0 $Y2=0
cc_153 N_Y_c_235_n N_VGND_c_292_n 0.00729487f $X=1.895 $Y=0.515 $X2=0 $Y2=0
cc_154 N_Y_c_233_n N_VGND_c_293_n 0.0369511f $X=1.73 $Y=0.435 $X2=0 $Y2=0
cc_155 N_Y_c_234_n N_VGND_c_293_n 0.00728664f $X=0.795 $Y=0.435 $X2=0 $Y2=0
cc_156 N_Y_c_235_n N_VGND_c_293_n 0.014693f $X=1.895 $Y=0.515 $X2=0 $Y2=0
cc_157 N_Y_c_233_n N_VGND_c_296_n 0.0316226f $X=1.73 $Y=0.435 $X2=0 $Y2=0
cc_158 N_Y_c_234_n N_VGND_c_296_n 0.00579633f $X=0.795 $Y=0.435 $X2=0 $Y2=0
cc_159 N_Y_c_235_n N_VGND_c_296_n 0.0121757f $X=1.895 $Y=0.515 $X2=0 $Y2=0
cc_160 N_Y_c_232_n A_145_74# 0.00586266f $X=0.71 $Y=1.72 $X2=-0.19 $Y2=-0.245
cc_161 N_Y_c_233_n A_145_74# 0.00427342f $X=1.73 $Y=0.435 $X2=-0.19 $Y2=-0.245
cc_162 N_Y_c_233_n A_223_74# 0.00868086f $X=1.73 $Y=0.435 $X2=-0.19 $Y2=-0.245

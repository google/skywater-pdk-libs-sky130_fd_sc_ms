* File: sky130_fd_sc_ms__inv_1.pex.spice
* Created: Fri Aug 28 17:37:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__INV_1%A 3 7 9 10 11 15
r21 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.65
+ $Y=1.465 $X2=0.65 $Y2=1.465
r22 11 15 10.2165 $w=4.78e-07 $l=4.1e-07 $layer=LI1_cond $X=0.24 $Y=1.54
+ $X2=0.65 $Y2=1.54
r23 9 14 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=0.835 $Y=1.465
+ $X2=0.65 $Y2=1.465
r24 9 10 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.835 $Y=1.465
+ $X2=0.925 $Y2=1.465
r25 5 10 34.7346 $w=1.65e-07 $l=1.69926e-07 $layer=POLY_cond $X=0.935 $Y=1.3
+ $X2=0.925 $Y2=1.465
r26 5 7 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.935 $Y=1.3 $X2=0.935
+ $Y2=0.74
r27 1 10 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.63
+ $X2=0.925 $Y2=1.465
r28 1 3 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.925 $Y=1.63
+ $X2=0.925 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__INV_1%VPWR 1 6 10 12 19 20 23
r14 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r15 17 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.65 $Y2=3.33
r16 17 19 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=1.2 $Y2=3.33
r17 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r18 12 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.485 $Y=3.33
+ $X2=0.65 $Y2=3.33
r19 12 14 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.485 $Y=3.33
+ $X2=0.24 $Y2=3.33
r20 10 20 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r21 10 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r22 10 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r23 6 9 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.65 $Y=2.115 $X2=0.65
+ $Y2=2.815
r24 4 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.65 $Y=3.245 $X2=0.65
+ $Y2=3.33
r25 4 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.65 $Y=3.245 $X2=0.65
+ $Y2=2.815
r26 1 9 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.505
+ $Y=1.84 $X2=0.65 $Y2=2.815
r27 1 6 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.505
+ $Y=1.84 $X2=0.65 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__INV_1%Y 1 2 7 8 9 10 11 12 13
r12 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=2.405
+ $X2=1.15 $Y2=2.775
r13 11 12 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.15 $Y=1.985
+ $X2=1.15 $Y2=2.405
r14 10 11 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=1.15 $Y=1.665
+ $X2=1.15 $Y2=1.985
r15 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=1.295
+ $X2=1.15 $Y2=1.665
r16 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=0.925 $X2=1.15
+ $Y2=1.295
r17 7 8 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.15 $Y=0.515 $X2=1.15
+ $Y2=0.925
r18 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.015
+ $Y=1.84 $X2=1.15 $Y2=2.815
r19 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.015
+ $Y=1.84 $X2=1.15 $Y2=1.985
r20 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.01
+ $Y=0.37 $X2=1.15 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__INV_1%VGND 1 6 8 10 17 18 21
r13 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r14 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.65
+ $Y2=0
r15 15 17 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=1.2
+ $Y2=0
r16 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r17 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.485 $Y=0 $X2=0.65
+ $Y2=0
r18 10 12 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.485 $Y=0 $X2=0.24
+ $Y2=0
r19 8 18 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r20 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r21 8 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r22 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.65 $Y=0.085 $X2=0.65
+ $Y2=0
r23 4 6 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.65 $Y=0.085 $X2=0.65
+ $Y2=0.515
r24 1 6 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.505
+ $Y=0.37 $X2=0.65 $Y2=0.515
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__clkbuf_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__clkbuf_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.264600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.055000 1.080000 2.455000 1.410000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.856800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.980000 1.750000 1.150000 ;
        RECT 0.535000 1.150000 0.705000 1.920000 ;
        RECT 0.535000 1.920000 1.795000 2.090000 ;
        RECT 0.535000 2.090000 0.815000 2.980000 ;
        RECT 0.560000 0.350000 0.890000 0.980000 ;
        RECT 1.420000 0.350000 1.750000 0.980000 ;
        RECT 1.465000 2.090000 1.795000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.115000  1.820000 0.365000 3.245000 ;
      RECT 0.130000  0.085000 0.380000 0.810000 ;
      RECT 0.875000  1.350000 1.885000 1.580000 ;
      RECT 0.875000  1.580000 2.795000 1.750000 ;
      RECT 1.015000  2.260000 1.265000 3.245000 ;
      RECT 1.070000  0.085000 1.240000 0.810000 ;
      RECT 1.920000  0.085000 2.250000 0.810000 ;
      RECT 1.995000  1.920000 2.245000 3.245000 ;
      RECT 2.415000  1.750000 2.795000 2.980000 ;
      RECT 2.420000  0.480000 2.795000 0.810000 ;
      RECT 2.625000  0.810000 2.795000 1.580000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_ms__clkbuf_4

* File: sky130_fd_sc_ms__o21bai_4.spice
* Created: Fri Aug 28 17:56:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o21bai_4.pex.spice"
.subckt sky130_fd_sc_ms__o21bai_4  VNB VPB A1 A2 B1_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1_N	B1_N
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A1_M1009_g N_A_27_74#_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1221 AS=0.2109 PD=1.07 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75005.4 A=0.111 P=1.78 MULT=1
MM1020 N_VGND_M1009_d N_A1_M1020_g N_A_27_74#_M1020_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1221 AS=0.1036 PD=1.07 PS=1.02 NRD=8.1 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75004.9 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1021_d N_A1_M1021_g N_A_27_74#_M1020_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75004.5 A=0.111 P=1.78 MULT=1
MM1023 N_VGND_M1021_d N_A1_M1023_g N_A_27_74#_M1023_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75004.1 A=0.111 P=1.78 MULT=1
MM1005 N_A_27_74#_M1023_s N_A2_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75003.7 A=0.111 P=1.78 MULT=1
MM1007 N_A_27_74#_M1007_d N_A2_M1007_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.4
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1019 N_A_27_74#_M1007_d N_A2_M1019_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1889 PD=1.02 PS=1.36 NRD=0 NRS=32.472 M=1 R=4.93333 SA=75002.8
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1024 N_A_27_74#_M1024_d N_A2_M1024_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1889 PD=1.09 PS=1.36 NRD=0 NRS=32.472 M=1 R=4.93333 SA=75003.4
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1000 N_Y_M1000_d N_A_828_48#_M1000_g N_A_27_74#_M1024_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75003.9 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1000_d N_A_828_48#_M1001_g N_A_27_74#_M1001_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75004.4 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1006 N_Y_M1006_d N_A_828_48#_M1006_g N_A_27_74#_M1001_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75004.9 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1018 N_Y_M1006_d N_A_828_48#_M1018_g N_A_27_74#_M1018_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.2627 PD=1.09 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75005.4 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_B1_N_M1010_g N_A_828_48#_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_28_368#_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003.4 A=0.2016 P=2.6 MULT=1
MM1003 N_VPWR_M1002_d N_A1_M1003_g N_A_28_368#_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90003 A=0.2016 P=2.6 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g N_A_28_368#_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90002.5 A=0.2016 P=2.6 MULT=1
MM1008 N_VPWR_M1004_d N_A1_M1008_g N_A_28_368#_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90002.1 A=0.2016 P=2.6 MULT=1
MM1011 N_Y_M1011_d N_A2_M1011_g N_A_28_368#_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1014 N_Y_M1011_d N_A2_M1014_g N_A_28_368#_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.4
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1016 N_Y_M1016_d N_A2_M1016_g N_A_28_368#_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90002.9
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1017 N_Y_M1016_d N_A2_M1017_g N_A_28_368#_M1017_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.3696 PD=1.44 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003.4
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1012 N_Y_M1012_d N_A_828_48#_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1596 PD=2.8 PS=1.405 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1022 N_Y_M1022_d N_A_828_48#_M1022_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1596 PD=2.8 PS=1.405 NRD=0 NRS=1.7533 M=1 R=6.22222 SA=90000.7
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1013 N_A_828_48#_M1013_d N_B1_N_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1134 AS=0.2352 PD=1.11 PS=2.24 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90000.6 A=0.1512 P=2.04 MULT=1
MM1015 N_A_828_48#_M1013_d N_B1_N_M1015_g N_VPWR_M1015_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1134 AS=0.2352 PD=1.11 PS=2.24 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90000.6 SB=90000.2 A=0.1512 P=2.04 MULT=1
DX25_noxref VNB VPB NWDIODE A=14.0988 P=18.88
*
.include "sky130_fd_sc_ms__o21bai_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__o41a_1.pex.spice
* Created: Wed Sep  2 12:26:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O41A_1%A_83_270# 1 2 9 13 16 18 19 20 22 23 26 30
c71 18 0 6.43674e-20 $X=0.62 $Y=1.515
r72 28 30 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=1.915 $Y=2.12
+ $X2=1.915 $Y2=2.13
r73 24 26 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=1.34 $Y=1.11
+ $X2=1.34 $Y2=0.515
r74 22 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.75 $Y=2.035
+ $X2=1.915 $Y2=2.12
r75 22 23 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=1.75 $Y=2.035
+ $X2=0.785 $Y2=2.035
r76 21 32 2.6346 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.785 $Y=1.195
+ $X2=0.62 $Y2=1.195
r77 20 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.175 $Y=1.195
+ $X2=1.34 $Y2=1.11
r78 20 21 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.175 $Y=1.195
+ $X2=0.785 $Y2=1.195
r79 19 35 40.9837 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.6 $Y=1.515
+ $X2=0.6 $Y2=1.68
r80 19 34 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.6 $Y=1.515
+ $X2=0.6 $Y2=1.35
r81 18 32 12.8588 $w=3.3e-07 $l=3.2e-07 $layer=LI1_cond $X=0.62 $Y=1.515
+ $X2=0.62 $Y2=1.195
r82 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.62
+ $Y=1.515 $X2=0.62 $Y2=1.515
r83 16 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.62 $Y=1.95
+ $X2=0.785 $Y2=2.035
r84 16 18 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=0.62 $Y=1.95
+ $X2=0.62 $Y2=1.515
r85 13 34 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=0.74
+ $X2=0.495 $Y2=1.35
r86 9 35 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.505 $Y=2.4
+ $X2=0.505 $Y2=1.68
r87 2 30 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=1.695
+ $Y=1.985 $X2=1.915 $Y2=2.13
r88 1 26 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.195
+ $Y=0.37 $X2=1.34 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_1%B1 3 5 7 8 12
c37 5 0 6.43674e-20 $X=1.605 $Y=1.91
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.415
+ $Y=1.615 $X2=1.415 $Y2=1.615
r39 8 12 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=1.415 $Y2=1.615
r40 5 11 50.2893 $w=4.01e-07 $l=3.55331e-07 $layer=POLY_cond $X=1.605 $Y=1.91
+ $X2=1.472 $Y2=1.615
r41 5 7 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=1.605 $Y=1.91
+ $X2=1.605 $Y2=2.405
r42 1 11 39.605 $w=4.01e-07 $l=2.02287e-07 $layer=POLY_cond $X=1.555 $Y=1.45
+ $X2=1.472 $Y2=1.615
r43 1 3 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.555 $Y=1.45
+ $X2=1.555 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_1%A4 3 5 7 9 13
r45 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.035
+ $Y=1.355 $X2=2.035 $Y2=1.355
r46 9 13 8.82117 $w=4.03e-07 $l=3.1e-07 $layer=LI1_cond $X=2.072 $Y=1.665
+ $X2=2.072 $Y2=1.355
r47 5 12 34.0194 $w=3.43e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.14 $Y=1.52
+ $X2=2.05 $Y2=1.355
r48 5 7 342.065 $w=1.8e-07 $l=8.8e-07 $layer=POLY_cond $X=2.14 $Y=1.52 $X2=2.14
+ $Y2=2.4
r49 1 12 38.7084 $w=3.43e-07 $l=1.67481e-07 $layer=POLY_cond $X=2.055 $Y=1.19
+ $X2=2.05 $Y2=1.355
r50 1 3 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.055 $Y=1.19 $X2=2.055
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_1%A3 3 7 9 10 11 12 18 19
r44 18 21 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.635 $Y=1.385
+ $X2=2.635 $Y2=1.55
r45 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.635 $Y=1.385
+ $X2=2.635 $Y2=1.22
r46 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.635
+ $Y=1.385 $X2=2.635 $Y2=1.385
r47 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.635 $Y=2.405
+ $X2=2.635 $Y2=2.775
r48 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.635 $Y=2.035
+ $X2=2.635 $Y2=2.405
r49 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.635 $Y=1.665
+ $X2=2.635 $Y2=2.035
r50 9 19 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=2.635 $Y=1.665
+ $X2=2.635 $Y2=1.385
r51 7 20 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.625 $Y=0.69
+ $X2=2.625 $Y2=1.22
r52 3 21 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.56 $Y=2.4 $X2=2.56
+ $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_1%A2 3 7 9 10 11 12 18 19
r38 18 21 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=1.465
+ $X2=3.205 $Y2=1.63
r39 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=1.465
+ $X2=3.205 $Y2=1.3
r40 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.205
+ $Y=1.465 $X2=3.205 $Y2=1.465
r41 11 12 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=3.187 $Y=2.405
+ $X2=3.187 $Y2=2.775
r42 10 11 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=3.187 $Y=2.035
+ $X2=3.187 $Y2=2.405
r43 9 10 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=3.187 $Y=1.665
+ $X2=3.187 $Y2=2.035
r44 9 19 6.31476 $w=3.63e-07 $l=2e-07 $layer=LI1_cond $X=3.187 $Y=1.665
+ $X2=3.187 $Y2=1.465
r45 7 21 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=3.13 $Y=2.4 $X2=3.13
+ $Y2=1.63
r46 3 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.115 $Y=0.69
+ $X2=3.115 $Y2=1.3
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_1%A1 3 7 9 10 14 15
r28 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.775 $Y=1.515
+ $X2=3.775 $Y2=1.68
r29 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.775 $Y=1.515
+ $X2=3.775 $Y2=1.35
r30 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.775
+ $Y=1.515 $X2=3.775 $Y2=1.515
r31 9 10 7.56494 $w=5.83e-07 $l=3.7e-07 $layer=LI1_cond $X=3.902 $Y=1.665
+ $X2=3.902 $Y2=2.035
r32 9 15 3.06687 $w=5.83e-07 $l=1.5e-07 $layer=LI1_cond $X=3.902 $Y=1.665
+ $X2=3.902 $Y2=1.515
r33 7 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.825 $Y=0.69
+ $X2=3.825 $Y2=1.35
r34 3 17 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.7 $Y=2.4 $X2=3.7
+ $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_1%X 1 2 9 13 14 15 26 28
r21 14 28 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=0.28 $Y=2.455 $X2=0.28
+ $Y2=2.405
r22 14 28 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=0.28 $Y=2.387
+ $X2=0.28 $Y2=2.405
r23 14 26 6.08745 $w=3.28e-07 $l=9.7e-08 $layer=LI1_cond $X=0.28 $Y=2.387
+ $X2=0.28 $Y2=2.29
r24 14 15 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.28 $Y=2.455
+ $X2=0.28 $Y2=2.775
r25 13 26 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=0.2 $Y=1.13 $X2=0.2
+ $Y2=2.29
r26 7 13 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.245 $Y=1 $X2=0.245
+ $Y2=1.13
r27 7 9 21.4975 $w=2.58e-07 $l=4.85e-07 $layer=LI1_cond $X=0.245 $Y=1 $X2=0.245
+ $Y2=0.515
r28 2 14 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.455
r29 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_1%VPWR 1 2 9 12 14 16 18 23 32 36
r45 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r46 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r47 30 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r48 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r49 27 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 26 29 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r51 26 27 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 24 32 15.7083 $w=1.7e-07 $l=4.63e-07 $layer=LI1_cond $X=1.54 $Y=3.33
+ $X2=1.077 $Y2=3.33
r53 24 26 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.54 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 23 35 5.79967 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=3.76 $Y=3.33 $X2=4.04
+ $Y2=3.33
r55 23 29 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.76 $Y=3.33 $X2=3.6
+ $Y2=3.33
r56 21 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r57 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r58 18 32 15.7083 $w=1.7e-07 $l=4.62e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=1.077 $Y2=3.33
r59 18 20 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r60 16 30 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r61 16 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 12 35 2.96198 $w=4.45e-07 $l=1.1025e-07 $layer=LI1_cond $X=3.982 $Y=3.245
+ $X2=4.04 $Y2=3.33
r63 12 14 21.754 $w=4.43e-07 $l=8.4e-07 $layer=LI1_cond $X=3.982 $Y=3.245
+ $X2=3.982 $Y2=2.405
r64 7 32 3.39807 $w=9.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.077 $Y=3.245
+ $X2=1.077 $Y2=3.33
r65 7 9 11.4746 $w=9.23e-07 $l=8.7e-07 $layer=LI1_cond $X=1.077 $Y=3.245
+ $X2=1.077 $Y2=2.375
r66 2 14 300 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=2 $X=3.79
+ $Y=1.84 $X2=3.925 $Y2=2.405
r67 1 9 300 $w=1.7e-07 $l=1.01277e-06 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=1.375 $Y2=2.375
r68 1 9 300 $w=1.7e-07 $l=6.20645e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.78 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_1%VGND 1 2 3 12 16 20 23 24 25 27 39 45 46 49
+ 52
r56 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r57 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r58 46 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r59 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r60 43 52 11.6921 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=3.705 $Y=0 $X2=3.44
+ $Y2=0
r61 43 45 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.705 $Y=0 $X2=4.08
+ $Y2=0
r62 42 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r63 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r64 39 52 11.6921 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=3.175 $Y=0 $X2=3.44
+ $Y2=0
r65 39 41 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.175 $Y=0 $X2=3.12
+ $Y2=0
r66 35 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r67 34 37 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r68 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r69 32 49 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.745
+ $Y2=0
r70 32 34 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r71 30 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r72 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r73 27 49 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.745
+ $Y2=0
r74 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r75 25 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r76 25 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r77 25 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r78 23 37 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.175 $Y=0 $X2=2.16
+ $Y2=0
r79 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.175 $Y=0 $X2=2.34
+ $Y2=0
r80 22 41 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=2.505 $Y=0 $X2=3.12
+ $Y2=0
r81 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=0 $X2=2.34
+ $Y2=0
r82 18 52 2.222 $w=5.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=0.085 $X2=3.44
+ $Y2=0
r83 18 20 9.70403 $w=5.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.44 $Y=0.085
+ $X2=3.44 $Y2=0.515
r84 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=0.085
+ $X2=2.34 $Y2=0
r85 14 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.34 $Y=0.085
+ $X2=2.34 $Y2=0.515
r86 10 49 1.46811 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0
r87 10 12 11.8125 $w=3.98e-07 $l=4.1e-07 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0.495
r88 3 20 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=3.19
+ $Y=0.37 $X2=3.44 $Y2=0.515
r89 2 16 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.13
+ $Y=0.37 $X2=2.34 $Y2=0.515
r90 1 12 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_MS__O41A_1%A_326_74# 1 2 3 12 14 15 18 20 24 26
r52 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.04 $Y=0.85
+ $X2=4.04 $Y2=0.515
r53 21 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.005 $Y=0.935
+ $X2=2.84 $Y2=0.935
r54 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.875 $Y=0.935
+ $X2=4.04 $Y2=0.85
r55 20 21 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=3.875 $Y=0.935
+ $X2=3.005 $Y2=0.935
r56 16 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=0.85 $X2=2.84
+ $Y2=0.935
r57 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.84 $Y=0.85
+ $X2=2.84 $Y2=0.515
r58 14 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.675 $Y=0.935
+ $X2=2.84 $Y2=0.935
r59 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.675 $Y=0.935
+ $X2=2.005 $Y2=0.935
r60 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.84 $Y=0.85
+ $X2=2.005 $Y2=0.935
r61 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.84 $Y=0.85
+ $X2=1.84 $Y2=0.515
r62 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.9
+ $Y=0.37 $X2=4.04 $Y2=0.515
r63 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.7
+ $Y=0.37 $X2=2.84 $Y2=0.515
r64 1 12 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.63
+ $Y=0.37 $X2=1.84 $Y2=0.515
.ends


* File: sky130_fd_sc_ms__o2bb2a_1.pxi.spice
* Created: Fri Aug 28 17:59:28 2020
* 
x_PM_SKY130_FD_SC_MS__O2BB2A_1%A_83_260# N_A_83_260#_M1006_s N_A_83_260#_M1007_d
+ N_A_83_260#_M1002_g N_A_83_260#_M1001_g N_A_83_260#_c_81_n N_A_83_260#_c_82_n
+ N_A_83_260#_c_83_n N_A_83_260#_c_84_n N_A_83_260#_c_85_n N_A_83_260#_c_86_n
+ N_A_83_260#_c_87_n N_A_83_260#_c_92_n N_A_83_260#_c_93_n N_A_83_260#_c_88_n
+ N_A_83_260#_c_89_n N_A_83_260#_c_94_n PM_SKY130_FD_SC_MS__O2BB2A_1%A_83_260#
x_PM_SKY130_FD_SC_MS__O2BB2A_1%A1_N N_A1_N_M1000_g N_A1_N_M1003_g A1_N
+ N_A1_N_c_184_n PM_SKY130_FD_SC_MS__O2BB2A_1%A1_N
x_PM_SKY130_FD_SC_MS__O2BB2A_1%A2_N N_A2_N_M1004_g N_A2_N_M1010_g A2_N
+ N_A2_N_c_223_n PM_SKY130_FD_SC_MS__O2BB2A_1%A2_N
x_PM_SKY130_FD_SC_MS__O2BB2A_1%A_236_384# N_A_236_384#_M1004_d
+ N_A_236_384#_M1000_d N_A_236_384#_c_255_n N_A_236_384#_c_256_n
+ N_A_236_384#_c_257_n N_A_236_384#_M1006_g N_A_236_384#_c_262_n
+ N_A_236_384#_M1007_g N_A_236_384#_c_258_n N_A_236_384#_c_259_n
+ N_A_236_384#_c_279_n N_A_236_384#_c_280_n N_A_236_384#_c_264_n
+ N_A_236_384#_c_260_n N_A_236_384#_c_261_n
+ PM_SKY130_FD_SC_MS__O2BB2A_1%A_236_384#
x_PM_SKY130_FD_SC_MS__O2BB2A_1%B2 N_B2_M1011_g N_B2_M1005_g B2 B2 N_B2_c_323_n
+ PM_SKY130_FD_SC_MS__O2BB2A_1%B2
x_PM_SKY130_FD_SC_MS__O2BB2A_1%B1 N_B1_c_362_n N_B1_M1008_g N_B1_M1009_g
+ N_B1_c_359_n B1 N_B1_c_361_n PM_SKY130_FD_SC_MS__O2BB2A_1%B1
x_PM_SKY130_FD_SC_MS__O2BB2A_1%X N_X_M1001_s N_X_M1002_s N_X_c_385_n N_X_c_386_n
+ X X X X N_X_c_387_n PM_SKY130_FD_SC_MS__O2BB2A_1%X
x_PM_SKY130_FD_SC_MS__O2BB2A_1%VPWR N_VPWR_M1002_d N_VPWR_M1010_d N_VPWR_M1008_d
+ N_VPWR_c_410_n N_VPWR_c_411_n N_VPWR_c_412_n VPWR N_VPWR_c_413_n
+ N_VPWR_c_414_n N_VPWR_c_415_n N_VPWR_c_416_n N_VPWR_c_417_n N_VPWR_c_409_n
+ PM_SKY130_FD_SC_MS__O2BB2A_1%VPWR
x_PM_SKY130_FD_SC_MS__O2BB2A_1%VGND N_VGND_M1001_d N_VGND_M1011_d N_VGND_c_456_n
+ N_VGND_c_457_n VGND N_VGND_c_458_n N_VGND_c_459_n N_VGND_c_460_n
+ N_VGND_c_461_n N_VGND_c_462_n N_VGND_c_463_n PM_SKY130_FD_SC_MS__O2BB2A_1%VGND
x_PM_SKY130_FD_SC_MS__O2BB2A_1%A_588_74# N_A_588_74#_M1006_d N_A_588_74#_M1009_d
+ N_A_588_74#_c_505_n N_A_588_74#_c_506_n N_A_588_74#_c_507_n
+ N_A_588_74#_c_508_n PM_SKY130_FD_SC_MS__O2BB2A_1%A_588_74#
cc_1 VNB N_A_83_260#_M1002_g 0.00185695f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A_83_260#_M1001_g 0.0293121f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.74
cc_3 VNB N_A_83_260#_c_81_n 0.0138399f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.165
cc_4 VNB N_A_83_260#_c_82_n 0.0094333f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.165
cc_5 VNB N_A_83_260#_c_83_n 6.79008e-19 $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=1.08
cc_6 VNB N_A_83_260#_c_84_n 0.0263861f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=0.34
cc_7 VNB N_A_83_260#_c_85_n 0.00270027f $X=-0.19 $Y=-0.245 $X2=1.46 $Y2=0.34
cc_8 VNB N_A_83_260#_c_86_n 0.00910354f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.495
cc_9 VNB N_A_83_260#_c_87_n 0.00580571f $X=-0.19 $Y=-0.245 $X2=2.73 $Y2=1.9
cc_10 VNB N_A_83_260#_c_88_n 0.033478f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.465
cc_11 VNB N_A_83_260#_c_89_n 0.00299619f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.92
cc_12 VNB N_A1_N_M1003_g 0.0235016f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.63
cc_13 VNB A1_N 0.0034197f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_14 VNB N_A1_N_c_184_n 0.0227092f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.74
cc_15 VNB N_A2_N_M1004_g 0.0297096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB A2_N 0.00166191f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_17 VNB N_A2_N_c_223_n 0.0208531f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.74
cc_18 VNB N_A_236_384#_c_255_n 0.0277098f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.63
cc_19 VNB N_A_236_384#_c_256_n 0.0199158f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_20 VNB N_A_236_384#_c_257_n 0.0185273f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_21 VNB N_A_236_384#_c_258_n 0.00526231f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=1.08
cc_22 VNB N_A_236_384#_c_259_n 0.0221028f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=0.34
cc_23 VNB N_A_236_384#_c_260_n 0.0106619f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.465
cc_24 VNB N_A_236_384#_c_261_n 0.0320751f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.465
cc_25 VNB N_B2_M1011_g 0.0219963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B2_M1005_g 0.00895283f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.63
cc_27 VNB B2 0.0175784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B2_c_323_n 0.0288405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B1_M1009_g 0.0297108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B1_c_359_n 0.0121866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB B1 0.00760591f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.3
cc_32 VNB N_B1_c_361_n 0.0575527f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.165
cc_33 VNB N_X_c_385_n 0.0267746f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_34 VNB N_X_c_386_n 0.0141322f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.74
cc_35 VNB N_X_c_387_n 0.0247901f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.465
cc_36 VNB N_VPWR_c_409_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_456_n 0.0101787f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_38 VNB N_VGND_c_457_n 0.00963715f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.74
cc_39 VNB N_VGND_c_458_n 0.0191572f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=0.425
cc_40 VNB N_VGND_c_459_n 0.0565361f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.755
cc_41 VNB N_VGND_c_460_n 0.018414f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.465
cc_42 VNB N_VGND_c_461_n 0.255724f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.465
cc_43 VNB N_VGND_c_462_n 0.00952121f $X=-0.19 $Y=-0.245 $X2=3.155 $Y2=1.985
cc_44 VNB N_VGND_c_463_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.3
cc_45 VNB N_A_588_74#_c_505_n 0.00210896f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_46 VNB N_A_588_74#_c_506_n 0.0085555f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.3
cc_47 VNB N_A_588_74#_c_507_n 0.00180855f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.74
cc_48 VNB N_A_588_74#_c_508_n 0.0208508f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.165
cc_49 VPB N_A_83_260#_M1002_g 0.0302708f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_50 VPB N_A_83_260#_c_87_n 0.00223621f $X=-0.19 $Y=1.66 $X2=2.73 $Y2=1.9
cc_51 VPB N_A_83_260#_c_92_n 6.52718e-19 $X=-0.19 $Y=1.66 $X2=2.99 $Y2=1.985
cc_52 VPB N_A_83_260#_c_93_n 2.22016e-19 $X=-0.19 $Y=1.66 $X2=2.815 $Y2=1.985
cc_53 VPB N_A_83_260#_c_94_n 0.00488472f $X=-0.19 $Y=1.66 $X2=3.155 $Y2=2.065
cc_54 VPB N_A1_N_M1000_g 0.0264606f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB A1_N 0.00391782f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_56 VPB N_A1_N_c_184_n 0.00737466f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=0.74
cc_57 VPB N_A2_N_M1010_g 0.0247671f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.63
cc_58 VPB A2_N 0.0015854f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_59 VPB N_A2_N_c_223_n 0.0113216f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=0.74
cc_60 VPB N_A_236_384#_c_262_n 0.0272195f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_236_384#_c_259_n 0.00497281f $X=-0.19 $Y=1.66 $X2=2.485 $Y2=0.34
cc_62 VPB N_A_236_384#_c_264_n 0.00314957f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_236_384#_c_261_n 0.0167473f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.465
cc_64 VPB N_B2_M1005_g 0.0283493f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.63
cc_65 VPB N_B1_c_362_n 0.0288486f $X=-0.19 $Y=1.66 $X2=2.505 $Y2=0.37
cc_66 VPB N_B1_c_359_n 0.00727927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB X 0.0136968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB X 0.0415472f $X=-0.19 $Y=1.66 $X2=2.65 $Y2=0.495
cc_69 VPB N_X_c_387_n 0.00769959f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.465
cc_70 VPB N_VPWR_c_410_n 0.0172963f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=0.74
cc_71 VPB N_VPWR_c_411_n 0.0123504f $X=-0.19 $Y=1.66 $X2=1.375 $Y2=1.08
cc_72 VPB N_VPWR_c_412_n 0.0546749f $X=-0.19 $Y=1.66 $X2=1.46 $Y2=0.34
cc_73 VPB N_VPWR_c_413_n 0.0189171f $X=-0.19 $Y=1.66 $X2=2.73 $Y2=1.9
cc_74 VPB N_VPWR_c_414_n 0.0316212f $X=-0.19 $Y=1.66 $X2=0.795 $Y2=1.165
cc_75 VPB N_VPWR_c_415_n 0.00632158f $X=-0.19 $Y=1.66 $X2=3.155 $Y2=2.065
cc_76 VPB N_VPWR_c_416_n 0.02253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_417_n 0.0543461f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_409_n 0.0911562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 N_A_83_260#_M1002_g N_A1_N_M1000_g 0.0158552f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_80 N_A_83_260#_M1001_g N_A1_N_M1003_g 0.0102428f $X=0.505 $Y=0.74 $X2=0 $Y2=0
cc_81 N_A_83_260#_c_81_n N_A1_N_M1003_g 0.0149897f $X=1.29 $Y=1.165 $X2=0 $Y2=0
cc_82 N_A_83_260#_c_82_n N_A1_N_M1003_g 0.00200333f $X=0.795 $Y=1.165 $X2=0
+ $Y2=0
cc_83 N_A_83_260#_c_83_n N_A1_N_M1003_g 0.0026876f $X=1.375 $Y=1.08 $X2=0 $Y2=0
cc_84 N_A_83_260#_c_85_n N_A1_N_M1003_g 6.82792e-19 $X=1.46 $Y=0.34 $X2=0 $Y2=0
cc_85 N_A_83_260#_c_88_n N_A1_N_M1003_g 0.00148094f $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_86 N_A_83_260#_M1002_g A1_N 8.28658e-19 $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_87 N_A_83_260#_c_81_n A1_N 0.0261759f $X=1.29 $Y=1.165 $X2=0 $Y2=0
cc_88 N_A_83_260#_c_82_n A1_N 0.0170081f $X=0.795 $Y=1.165 $X2=0 $Y2=0
cc_89 N_A_83_260#_c_88_n A1_N 2.41701e-19 $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_90 N_A_83_260#_M1002_g N_A1_N_c_184_n 0.00234771f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_91 N_A_83_260#_c_81_n N_A1_N_c_184_n 0.00490114f $X=1.29 $Y=1.165 $X2=0 $Y2=0
cc_92 N_A_83_260#_c_82_n N_A1_N_c_184_n 0.00237388f $X=0.795 $Y=1.165 $X2=0
+ $Y2=0
cc_93 N_A_83_260#_c_88_n N_A1_N_c_184_n 0.0180042f $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_94 N_A_83_260#_c_81_n N_A2_N_M1004_g 0.00118344f $X=1.29 $Y=1.165 $X2=0 $Y2=0
cc_95 N_A_83_260#_c_83_n N_A2_N_M1004_g 0.00330892f $X=1.375 $Y=1.08 $X2=0 $Y2=0
cc_96 N_A_83_260#_c_84_n N_A2_N_M1004_g 0.0121086f $X=2.485 $Y=0.34 $X2=0 $Y2=0
cc_97 N_A_83_260#_c_87_n N_A_236_384#_c_255_n 0.00944143f $X=2.73 $Y=1.9 $X2=0
+ $Y2=0
cc_98 N_A_83_260#_c_89_n N_A_236_384#_c_255_n 0.00646708f $X=2.65 $Y=0.92 $X2=0
+ $Y2=0
cc_99 N_A_83_260#_c_84_n N_A_236_384#_c_256_n 0.00825806f $X=2.485 $Y=0.34 $X2=0
+ $Y2=0
cc_100 N_A_83_260#_c_84_n N_A_236_384#_c_257_n 0.00534381f $X=2.485 $Y=0.34
+ $X2=0 $Y2=0
cc_101 N_A_83_260#_c_86_n N_A_236_384#_c_257_n 0.00338973f $X=2.65 $Y=0.495
+ $X2=0 $Y2=0
cc_102 N_A_83_260#_c_87_n N_A_236_384#_c_257_n 0.00361776f $X=2.73 $Y=1.9 $X2=0
+ $Y2=0
cc_103 N_A_83_260#_c_89_n N_A_236_384#_c_257_n 0.00170336f $X=2.65 $Y=0.92 $X2=0
+ $Y2=0
cc_104 N_A_83_260#_c_87_n N_A_236_384#_c_262_n 0.0052021f $X=2.73 $Y=1.9 $X2=0
+ $Y2=0
cc_105 N_A_83_260#_c_92_n N_A_236_384#_c_262_n 0.0158895f $X=2.99 $Y=1.985 $X2=0
+ $Y2=0
cc_106 N_A_83_260#_c_93_n N_A_236_384#_c_262_n 0.00387599f $X=2.815 $Y=1.985
+ $X2=0 $Y2=0
cc_107 N_A_83_260#_c_94_n N_A_236_384#_c_262_n 0.00104557f $X=3.155 $Y=2.065
+ $X2=0 $Y2=0
cc_108 N_A_83_260#_c_87_n N_A_236_384#_c_258_n 0.00216975f $X=2.73 $Y=1.9 $X2=0
+ $Y2=0
cc_109 N_A_83_260#_c_87_n N_A_236_384#_c_259_n 0.0122328f $X=2.73 $Y=1.9 $X2=0
+ $Y2=0
cc_110 N_A_83_260#_c_93_n N_A_236_384#_c_279_n 0.00777292f $X=2.815 $Y=1.985
+ $X2=0 $Y2=0
cc_111 N_A_83_260#_c_84_n N_A_236_384#_c_280_n 0.0164516f $X=2.485 $Y=0.34 $X2=0
+ $Y2=0
cc_112 N_A_83_260#_c_86_n N_A_236_384#_c_280_n 0.0104187f $X=2.65 $Y=0.495 $X2=0
+ $Y2=0
cc_113 N_A_83_260#_c_87_n N_A_236_384#_c_264_n 0.035097f $X=2.73 $Y=1.9 $X2=0
+ $Y2=0
cc_114 N_A_83_260#_c_93_n N_A_236_384#_c_264_n 0.00310584f $X=2.815 $Y=1.985
+ $X2=0 $Y2=0
cc_115 N_A_83_260#_c_81_n N_A_236_384#_c_260_n 0.0132372f $X=1.29 $Y=1.165 $X2=0
+ $Y2=0
cc_116 N_A_83_260#_c_84_n N_A_236_384#_c_260_n 0.0132653f $X=2.485 $Y=0.34 $X2=0
+ $Y2=0
cc_117 N_A_83_260#_c_87_n N_A_236_384#_c_260_n 0.00900461f $X=2.73 $Y=1.9 $X2=0
+ $Y2=0
cc_118 N_A_83_260#_c_87_n N_A_236_384#_c_261_n 0.00379203f $X=2.73 $Y=1.9 $X2=0
+ $Y2=0
cc_119 N_A_83_260#_c_84_n N_B2_M1011_g 2.94862e-19 $X=2.485 $Y=0.34 $X2=0 $Y2=0
cc_120 N_A_83_260#_c_87_n N_B2_M1011_g 8.2968e-19 $X=2.73 $Y=1.9 $X2=0 $Y2=0
cc_121 N_A_83_260#_c_87_n N_B2_M1005_g 0.00185135f $X=2.73 $Y=1.9 $X2=0 $Y2=0
cc_122 N_A_83_260#_c_94_n N_B2_M1005_g 0.0187374f $X=3.155 $Y=2.065 $X2=0 $Y2=0
cc_123 N_A_83_260#_c_87_n B2 0.0244039f $X=2.73 $Y=1.9 $X2=0 $Y2=0
cc_124 N_A_83_260#_c_94_n B2 0.014975f $X=3.155 $Y=2.065 $X2=0 $Y2=0
cc_125 N_A_83_260#_c_87_n N_B2_c_323_n 2.57511e-19 $X=2.73 $Y=1.9 $X2=0 $Y2=0
cc_126 N_A_83_260#_c_94_n N_B2_c_323_n 0.00268889f $X=3.155 $Y=2.065 $X2=0 $Y2=0
cc_127 N_A_83_260#_c_94_n N_B1_c_362_n 0.00245317f $X=3.155 $Y=2.065 $X2=-0.19
+ $Y2=-0.245
cc_128 N_A_83_260#_M1001_g N_X_c_385_n 0.0084877f $X=0.505 $Y=0.74 $X2=0 $Y2=0
cc_129 N_A_83_260#_M1001_g N_X_c_386_n 0.00427425f $X=0.505 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A_83_260#_c_82_n N_X_c_386_n 0.00515361f $X=0.795 $Y=1.165 $X2=0 $Y2=0
cc_131 N_A_83_260#_c_88_n N_X_c_386_n 5.22956e-19 $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_132 N_A_83_260#_M1002_g X 0.0045132f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_133 N_A_83_260#_c_82_n X 0.00139316f $X=0.795 $Y=1.165 $X2=0 $Y2=0
cc_134 N_A_83_260#_M1002_g X 0.0128957f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_135 N_A_83_260#_M1001_g N_X_c_387_n 0.00252147f $X=0.505 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A_83_260#_c_82_n N_X_c_387_n 0.0307714f $X=0.795 $Y=1.165 $X2=0 $Y2=0
cc_137 N_A_83_260#_c_88_n N_X_c_387_n 0.0124571f $X=0.59 $Y=1.465 $X2=0 $Y2=0
cc_138 N_A_83_260#_c_93_n N_VPWR_M1010_d 0.00346975f $X=2.815 $Y=1.985 $X2=0
+ $Y2=0
cc_139 N_A_83_260#_M1002_g N_VPWR_c_410_n 0.00541032f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_140 N_A_83_260#_c_82_n N_VPWR_c_410_n 0.00860035f $X=0.795 $Y=1.165 $X2=0
+ $Y2=0
cc_141 N_A_83_260#_c_88_n N_VPWR_c_410_n 8.70386e-19 $X=0.59 $Y=1.465 $X2=0
+ $Y2=0
cc_142 N_A_83_260#_c_94_n N_VPWR_c_412_n 0.0254482f $X=3.155 $Y=2.065 $X2=0
+ $Y2=0
cc_143 N_A_83_260#_M1002_g N_VPWR_c_413_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A_83_260#_c_94_n N_VPWR_c_414_n 0.00707426f $X=3.155 $Y=2.065 $X2=0
+ $Y2=0
cc_145 N_A_83_260#_c_93_n N_VPWR_c_417_n 0.00541727f $X=2.815 $Y=1.985 $X2=0
+ $Y2=0
cc_146 N_A_83_260#_c_94_n N_VPWR_c_417_n 0.0146526f $X=3.155 $Y=2.065 $X2=0
+ $Y2=0
cc_147 N_A_83_260#_M1002_g N_VPWR_c_409_n 0.00990469f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_148 N_A_83_260#_c_94_n N_VPWR_c_409_n 0.010555f $X=3.155 $Y=2.065 $X2=0 $Y2=0
cc_149 N_A_83_260#_c_81_n N_VGND_M1001_d 0.00300823f $X=1.29 $Y=1.165 $X2=-0.19
+ $Y2=-0.245
cc_150 N_A_83_260#_c_82_n N_VGND_M1001_d 0.00199955f $X=0.795 $Y=1.165 $X2=-0.19
+ $Y2=-0.245
cc_151 N_A_83_260#_M1001_g N_VGND_c_456_n 0.00660116f $X=0.505 $Y=0.74 $X2=0
+ $Y2=0
cc_152 N_A_83_260#_c_81_n N_VGND_c_456_n 0.0216234f $X=1.29 $Y=1.165 $X2=0 $Y2=0
cc_153 N_A_83_260#_c_82_n N_VGND_c_456_n 0.0140249f $X=0.795 $Y=1.165 $X2=0
+ $Y2=0
cc_154 N_A_83_260#_c_83_n N_VGND_c_456_n 0.0209803f $X=1.375 $Y=1.08 $X2=0 $Y2=0
cc_155 N_A_83_260#_c_85_n N_VGND_c_456_n 0.0151159f $X=1.46 $Y=0.34 $X2=0 $Y2=0
cc_156 N_A_83_260#_c_88_n N_VGND_c_456_n 5.97302e-19 $X=0.59 $Y=1.465 $X2=0
+ $Y2=0
cc_157 N_A_83_260#_c_84_n N_VGND_c_457_n 0.00270678f $X=2.485 $Y=0.34 $X2=0
+ $Y2=0
cc_158 N_A_83_260#_M1001_g N_VGND_c_458_n 0.00434272f $X=0.505 $Y=0.74 $X2=0
+ $Y2=0
cc_159 N_A_83_260#_c_84_n N_VGND_c_459_n 0.08952f $X=2.485 $Y=0.34 $X2=0 $Y2=0
cc_160 N_A_83_260#_c_85_n N_VGND_c_459_n 0.0121867f $X=1.46 $Y=0.34 $X2=0 $Y2=0
cc_161 N_A_83_260#_M1001_g N_VGND_c_461_n 0.00828751f $X=0.505 $Y=0.74 $X2=0
+ $Y2=0
cc_162 N_A_83_260#_c_84_n N_VGND_c_461_n 0.0512413f $X=2.485 $Y=0.34 $X2=0 $Y2=0
cc_163 N_A_83_260#_c_85_n N_VGND_c_461_n 0.00660921f $X=1.46 $Y=0.34 $X2=0 $Y2=0
cc_164 N_A_83_260#_c_83_n A_253_94# 0.00212313f $X=1.375 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_165 N_A_83_260#_c_84_n N_A_588_74#_c_505_n 0.00453469f $X=2.485 $Y=0.34 $X2=0
+ $Y2=0
cc_166 N_A1_N_M1003_g N_A2_N_M1004_g 0.0466035f $X=1.19 $Y=0.79 $X2=0 $Y2=0
cc_167 A1_N N_A2_N_M1004_g 0.00229262f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_168 N_A1_N_c_184_n N_A2_N_M1004_g 0.0230306f $X=1.13 $Y=1.545 $X2=0 $Y2=0
cc_169 A1_N A2_N 0.0255141f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_170 N_A1_N_c_184_n A2_N 3.38054e-19 $X=1.13 $Y=1.545 $X2=0 $Y2=0
cc_171 N_A1_N_M1000_g N_A2_N_c_223_n 0.0304101f $X=1.09 $Y=2.34 $X2=0 $Y2=0
cc_172 N_A1_N_M1000_g N_A_236_384#_c_279_n 0.00576164f $X=1.09 $Y=2.34 $X2=0
+ $Y2=0
cc_173 A1_N N_A_236_384#_c_279_n 0.0111062f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_174 N_A1_N_c_184_n N_A_236_384#_c_279_n 5.74989e-19 $X=1.13 $Y=1.545 $X2=0
+ $Y2=0
cc_175 N_A1_N_M1003_g N_X_c_385_n 6.5955e-19 $X=1.19 $Y=0.79 $X2=0 $Y2=0
cc_176 N_A1_N_M1000_g X 7.67894e-19 $X=1.09 $Y=2.34 $X2=0 $Y2=0
cc_177 N_A1_N_M1000_g N_VPWR_c_410_n 0.00861351f $X=1.09 $Y=2.34 $X2=0 $Y2=0
cc_178 N_A1_N_M1000_g N_VPWR_c_416_n 0.00534617f $X=1.09 $Y=2.34 $X2=0 $Y2=0
cc_179 N_A1_N_M1000_g N_VPWR_c_417_n 0.00203214f $X=1.09 $Y=2.34 $X2=0 $Y2=0
cc_180 N_A1_N_M1000_g N_VPWR_c_409_n 0.00581878f $X=1.09 $Y=2.34 $X2=0 $Y2=0
cc_181 N_A1_N_M1003_g N_VGND_c_456_n 0.00998285f $X=1.19 $Y=0.79 $X2=0 $Y2=0
cc_182 N_A1_N_M1003_g N_VGND_c_459_n 0.00489033f $X=1.19 $Y=0.79 $X2=0 $Y2=0
cc_183 N_A1_N_M1003_g N_VGND_c_461_n 0.00500719f $X=1.19 $Y=0.79 $X2=0 $Y2=0
cc_184 N_A2_N_M1004_g N_A_236_384#_c_256_n 0.0105126f $X=1.58 $Y=0.79 $X2=0
+ $Y2=0
cc_185 N_A2_N_M1010_g N_A_236_384#_c_279_n 0.0230811f $X=1.595 $Y=2.34 $X2=0
+ $Y2=0
cc_186 A2_N N_A_236_384#_c_279_n 0.0235602f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_187 N_A2_N_c_223_n N_A_236_384#_c_279_n 9.03803e-19 $X=1.67 $Y=1.595 $X2=0
+ $Y2=0
cc_188 N_A2_N_M1004_g N_A_236_384#_c_280_n 0.00735949f $X=1.58 $Y=0.79 $X2=0
+ $Y2=0
cc_189 N_A2_N_M1004_g N_A_236_384#_c_264_n 9.76708e-19 $X=1.58 $Y=0.79 $X2=0
+ $Y2=0
cc_190 N_A2_N_M1010_g N_A_236_384#_c_264_n 0.0053099f $X=1.595 $Y=2.34 $X2=0
+ $Y2=0
cc_191 A2_N N_A_236_384#_c_264_n 0.0219371f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_192 N_A2_N_c_223_n N_A_236_384#_c_264_n 0.00116124f $X=1.67 $Y=1.595 $X2=0
+ $Y2=0
cc_193 N_A2_N_M1004_g N_A_236_384#_c_260_n 0.00474488f $X=1.58 $Y=0.79 $X2=0
+ $Y2=0
cc_194 A2_N N_A_236_384#_c_260_n 0.0153833f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_195 N_A2_N_c_223_n N_A_236_384#_c_260_n 0.00125903f $X=1.67 $Y=1.595 $X2=0
+ $Y2=0
cc_196 A2_N N_A_236_384#_c_261_n 0.00116124f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_197 N_A2_N_c_223_n N_A_236_384#_c_261_n 0.0195426f $X=1.67 $Y=1.595 $X2=0
+ $Y2=0
cc_198 N_A2_N_M1010_g N_VPWR_c_416_n 0.0044453f $X=1.595 $Y=2.34 $X2=0 $Y2=0
cc_199 N_A2_N_M1010_g N_VPWR_c_417_n 0.0136796f $X=1.595 $Y=2.34 $X2=0 $Y2=0
cc_200 N_A2_N_M1010_g N_VPWR_c_409_n 0.00484898f $X=1.595 $Y=2.34 $X2=0 $Y2=0
cc_201 N_A2_N_M1004_g N_VGND_c_456_n 2.05365e-19 $X=1.58 $Y=0.79 $X2=0 $Y2=0
cc_202 N_A2_N_M1004_g N_VGND_c_459_n 7.64118e-19 $X=1.58 $Y=0.79 $X2=0 $Y2=0
cc_203 N_A_236_384#_c_257_n N_B2_M1011_g 0.0137058f $X=2.865 $Y=1.09 $X2=0 $Y2=0
cc_204 N_A_236_384#_c_262_n N_B2_M1005_g 0.0160016f $X=2.88 $Y=1.84 $X2=0 $Y2=0
cc_205 N_A_236_384#_c_259_n N_B2_M1005_g 0.0085276f $X=2.88 $Y=1.75 $X2=0 $Y2=0
cc_206 N_A_236_384#_c_258_n B2 0.0026374f $X=2.865 $Y=1.165 $X2=0 $Y2=0
cc_207 N_A_236_384#_c_258_n N_B2_c_323_n 0.0166018f $X=2.865 $Y=1.165 $X2=0
+ $Y2=0
cc_208 N_A_236_384#_c_279_n N_VPWR_M1010_d 0.030922f $X=2.05 $Y=2.115 $X2=0
+ $Y2=0
cc_209 N_A_236_384#_c_264_n N_VPWR_M1010_d 9.17904e-19 $X=2.215 $Y=1.95 $X2=0
+ $Y2=0
cc_210 N_A_236_384#_c_262_n N_VPWR_c_414_n 0.0044453f $X=2.88 $Y=1.84 $X2=0
+ $Y2=0
cc_211 N_A_236_384#_c_262_n N_VPWR_c_417_n 0.0105526f $X=2.88 $Y=1.84 $X2=0
+ $Y2=0
cc_212 N_A_236_384#_c_279_n N_VPWR_c_417_n 0.0579491f $X=2.05 $Y=2.115 $X2=0
+ $Y2=0
cc_213 N_A_236_384#_c_261_n N_VPWR_c_417_n 9.36276e-19 $X=2.215 $Y=1.255 $X2=0
+ $Y2=0
cc_214 N_A_236_384#_c_262_n N_VPWR_c_409_n 0.00484898f $X=2.88 $Y=1.84 $X2=0
+ $Y2=0
cc_215 N_A_236_384#_c_257_n N_VGND_c_459_n 0.00430908f $X=2.865 $Y=1.09 $X2=0
+ $Y2=0
cc_216 N_A_236_384#_c_257_n N_VGND_c_461_n 0.00821764f $X=2.865 $Y=1.09 $X2=0
+ $Y2=0
cc_217 N_A_236_384#_c_257_n N_A_588_74#_c_505_n 2.18574e-19 $X=2.865 $Y=1.09
+ $X2=0 $Y2=0
cc_218 N_B2_M1005_g N_B1_c_362_n 0.0682545f $X=3.39 $Y=2.42 $X2=-0.19 $Y2=-0.245
cc_219 N_B2_M1011_g N_B1_M1009_g 0.0217086f $X=3.295 $Y=0.69 $X2=0 $Y2=0
cc_220 N_B2_M1005_g N_B1_c_359_n 0.0126967f $X=3.39 $Y=2.42 $X2=0 $Y2=0
cc_221 B2 B1 0.0277564f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_222 N_B2_c_323_n B1 2.37823e-19 $X=3.345 $Y=1.345 $X2=0 $Y2=0
cc_223 B2 N_B1_c_361_n 0.00294527f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_224 N_B2_c_323_n N_B1_c_361_n 0.0175815f $X=3.345 $Y=1.345 $X2=0 $Y2=0
cc_225 N_B2_M1005_g N_VPWR_c_412_n 0.00380326f $X=3.39 $Y=2.42 $X2=0 $Y2=0
cc_226 N_B2_M1005_g N_VPWR_c_414_n 0.00641103f $X=3.39 $Y=2.42 $X2=0 $Y2=0
cc_227 N_B2_M1005_g N_VPWR_c_417_n 0.00527091f $X=3.39 $Y=2.42 $X2=0 $Y2=0
cc_228 N_B2_M1005_g N_VPWR_c_409_n 0.00639697f $X=3.39 $Y=2.42 $X2=0 $Y2=0
cc_229 N_B2_M1011_g N_VGND_c_457_n 0.00363829f $X=3.295 $Y=0.69 $X2=0 $Y2=0
cc_230 N_B2_M1011_g N_VGND_c_459_n 0.00434054f $X=3.295 $Y=0.69 $X2=0 $Y2=0
cc_231 N_B2_M1011_g N_VGND_c_461_n 0.00445726f $X=3.295 $Y=0.69 $X2=0 $Y2=0
cc_232 N_B2_M1011_g N_A_588_74#_c_505_n 0.00711952f $X=3.295 $Y=0.69 $X2=0 $Y2=0
cc_233 N_B2_M1011_g N_A_588_74#_c_506_n 0.0090049f $X=3.295 $Y=0.69 $X2=0 $Y2=0
cc_234 B2 N_A_588_74#_c_506_n 0.0323411f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_235 N_B2_c_323_n N_A_588_74#_c_506_n 0.00344722f $X=3.345 $Y=1.345 $X2=0
+ $Y2=0
cc_236 N_B2_M1011_g N_A_588_74#_c_507_n 7.17385e-19 $X=3.295 $Y=0.69 $X2=0 $Y2=0
cc_237 B2 N_A_588_74#_c_507_n 0.0178517f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_238 N_B1_c_362_n N_VPWR_c_412_n 0.0261686f $X=3.81 $Y=1.84 $X2=0 $Y2=0
cc_239 B1 N_VPWR_c_412_n 0.014201f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_240 N_B1_c_361_n N_VPWR_c_412_n 0.00211705f $X=4.05 $Y=1.345 $X2=0 $Y2=0
cc_241 N_B1_c_362_n N_VPWR_c_414_n 0.00547402f $X=3.81 $Y=1.84 $X2=0 $Y2=0
cc_242 N_B1_c_362_n N_VPWR_c_409_n 0.00536634f $X=3.81 $Y=1.84 $X2=0 $Y2=0
cc_243 N_B1_M1009_g N_VGND_c_457_n 0.00330983f $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_244 N_B1_M1009_g N_VGND_c_460_n 0.00461464f $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_245 N_B1_M1009_g N_VGND_c_461_n 0.00467092f $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_246 N_B1_M1009_g N_A_588_74#_c_505_n 6.85083e-19 $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_247 N_B1_M1009_g N_A_588_74#_c_506_n 0.0144732f $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_248 B1 N_A_588_74#_c_506_n 0.0237154f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_249 N_B1_c_361_n N_A_588_74#_c_506_n 0.00196043f $X=4.05 $Y=1.345 $X2=0 $Y2=0
cc_250 N_B1_M1009_g N_A_588_74#_c_508_n 6.81345e-19 $X=3.825 $Y=0.69 $X2=0 $Y2=0
cc_251 X N_VPWR_c_410_n 0.0399187f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_252 X N_VPWR_c_413_n 0.0158876f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_253 X N_VPWR_c_409_n 0.0130823f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_254 N_X_c_385_n N_VGND_c_456_n 0.0222242f $X=0.29 $Y=0.515 $X2=0 $Y2=0
cc_255 N_X_c_385_n N_VGND_c_458_n 0.0163488f $X=0.29 $Y=0.515 $X2=0 $Y2=0
cc_256 N_X_c_385_n N_VGND_c_461_n 0.0134757f $X=0.29 $Y=0.515 $X2=0 $Y2=0
cc_257 N_VGND_c_457_n N_A_588_74#_c_505_n 0.0130732f $X=3.58 $Y=0.55 $X2=0 $Y2=0
cc_258 N_VGND_c_459_n N_A_588_74#_c_505_n 0.0114427f $X=3.415 $Y=0 $X2=0 $Y2=0
cc_259 N_VGND_c_461_n N_A_588_74#_c_505_n 0.00909435f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_260 N_VGND_M1011_d N_A_588_74#_c_506_n 0.00561113f $X=3.37 $Y=0.37 $X2=0
+ $Y2=0
cc_261 N_VGND_c_457_n N_A_588_74#_c_506_n 0.0211672f $X=3.58 $Y=0.55 $X2=0 $Y2=0
cc_262 N_VGND_c_461_n N_A_588_74#_c_506_n 0.0122262f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_263 N_VGND_c_457_n N_A_588_74#_c_508_n 0.00203724f $X=3.58 $Y=0.55 $X2=0
+ $Y2=0
cc_264 N_VGND_c_460_n N_A_588_74#_c_508_n 0.0115155f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_265 N_VGND_c_461_n N_A_588_74#_c_508_n 0.00920958f $X=4.08 $Y=0 $X2=0 $Y2=0

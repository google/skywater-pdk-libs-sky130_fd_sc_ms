* File: sky130_fd_sc_ms__nor4_2.pxi.spice
* Created: Fri Aug 28 17:49:34 2020
* 
x_PM_SKY130_FD_SC_MS__NOR4_2%C N_C_M1001_g N_C_M1008_g N_C_M1002_g N_C_c_83_n
+ N_C_c_84_n C C N_C_c_85_n N_C_c_86_n C N_C_c_88_n PM_SKY130_FD_SC_MS__NOR4_2%C
x_PM_SKY130_FD_SC_MS__NOR4_2%D N_D_c_152_n N_D_M1004_g N_D_c_153_n N_D_c_154_n
+ N_D_M1006_g N_D_c_156_n N_D_M1005_g D N_D_c_158_n PM_SKY130_FD_SC_MS__NOR4_2%D
x_PM_SKY130_FD_SC_MS__NOR4_2%B N_B_M1003_g N_B_M1009_g N_B_M1011_g N_B_c_218_n
+ N_B_c_211_n N_B_c_212_n B B B B N_B_c_213_n N_B_c_214_n N_B_c_215_n
+ N_B_c_221_n B PM_SKY130_FD_SC_MS__NOR4_2%B
x_PM_SKY130_FD_SC_MS__NOR4_2%A N_A_M1007_g N_A_c_288_n N_A_M1000_g N_A_M1010_g A
+ N_A_c_291_n PM_SKY130_FD_SC_MS__NOR4_2%A
x_PM_SKY130_FD_SC_MS__NOR4_2%A_27_368# N_A_27_368#_M1001_s N_A_27_368#_M1008_s
+ N_A_27_368#_M1011_s N_A_27_368#_c_331_n N_A_27_368#_c_338_n
+ N_A_27_368#_c_332_n N_A_27_368#_c_353_n N_A_27_368#_c_333_n
+ N_A_27_368#_c_334_n N_A_27_368#_c_335_n N_A_27_368#_c_336_n
+ PM_SKY130_FD_SC_MS__NOR4_2%A_27_368#
x_PM_SKY130_FD_SC_MS__NOR4_2%A_119_368# N_A_119_368#_M1001_d
+ N_A_119_368#_M1006_s N_A_119_368#_c_393_n
+ PM_SKY130_FD_SC_MS__NOR4_2%A_119_368#
x_PM_SKY130_FD_SC_MS__NOR4_2%Y N_Y_M1005_d N_Y_M1009_d N_Y_M1004_d N_Y_c_408_n
+ N_Y_c_409_n N_Y_c_410_n N_Y_c_416_n N_Y_c_411_n N_Y_c_412_n N_Y_c_413_n
+ N_Y_c_414_n Y Y N_Y_c_418_n PM_SKY130_FD_SC_MS__NOR4_2%Y
x_PM_SKY130_FD_SC_MS__NOR4_2%A_493_368# N_A_493_368#_M1003_d
+ N_A_493_368#_M1010_s N_A_493_368#_c_492_n N_A_493_368#_c_489_n
+ N_A_493_368#_c_484_n N_A_493_368#_c_485_n
+ PM_SKY130_FD_SC_MS__NOR4_2%A_493_368#
x_PM_SKY130_FD_SC_MS__NOR4_2%VPWR N_VPWR_M1007_d N_VPWR_c_513_n VPWR
+ N_VPWR_c_514_n N_VPWR_c_515_n N_VPWR_c_512_n N_VPWR_c_517_n
+ PM_SKY130_FD_SC_MS__NOR4_2%VPWR
x_PM_SKY130_FD_SC_MS__NOR4_2%VGND N_VGND_M1005_s N_VGND_M1002_d N_VGND_M1000_d
+ N_VGND_c_559_n N_VGND_c_560_n N_VGND_c_561_n VGND N_VGND_c_562_n
+ N_VGND_c_563_n N_VGND_c_564_n N_VGND_c_565_n N_VGND_c_566_n N_VGND_c_567_n
+ N_VGND_c_568_n PM_SKY130_FD_SC_MS__NOR4_2%VGND
cc_1 VNB N_C_M1001_g 0.00985164f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_C_M1008_g 5.18536e-19 $X=-0.19 $Y=-0.245 $X2=1.895 $Y2=2.4
cc_3 VNB N_C_M1002_g 0.0248615f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=0.74
cc_4 VNB N_C_c_83_n 0.00272143f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.335
cc_5 VNB N_C_c_84_n 0.0325028f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.335
cc_6 VNB N_C_c_85_n 0.0271624f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=1.485
cc_7 VNB N_C_c_86_n 0.00590745f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=1.485
cc_8 VNB C 6.99497e-19 $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.665
cc_9 VNB N_C_c_88_n 0.00494578f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.485
cc_10 VNB N_D_c_152_n 0.0378968f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.5
cc_11 VNB N_D_c_153_n 0.018773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_D_c_154_n 0.0466197f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=1.32
cc_13 VNB N_D_M1006_g 0.00743291f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=0.74
cc_14 VNB N_D_c_156_n 0.016723f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.41
cc_15 VNB D 0.00434149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_D_c_158_n 0.0732973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B_M1003_g 4.98563e-19 $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_18 VNB N_B_M1009_g 0.024237f $X=-0.19 $Y=-0.245 $X2=1.895 $Y2=2.4
cc_19 VNB N_B_M1011_g 0.00193177f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=0.74
cc_20 VNB N_B_c_211_n 0.00715627f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.335
cc_21 VNB N_B_c_212_n 0.0276743f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.335
cc_22 VNB N_B_c_213_n 0.163114f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=1.485
cc_23 VNB N_B_c_214_n 0.00361276f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=1.485
cc_24 VNB N_B_c_215_n 0.0392861f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.7
cc_25 VNB N_A_M1007_g 0.00577383f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_26 VNB N_A_c_288_n 0.0200555f $X=-0.19 $Y=-0.245 $X2=1.895 $Y2=1.65
cc_27 VNB N_A_M1010_g 0.00599095f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=0.74
cc_28 VNB A 0.021158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_c_291_n 0.0490677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_408_n 0.0320702f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=0.74
cc_31 VNB N_Y_c_409_n 0.00804079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_410_n 0.00833338f $X=-0.19 $Y=-0.245 $X2=1.565 $Y2=1.41
cc_33 VNB N_Y_c_411_n 0.00280855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_Y_c_412_n 0.00861013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_Y_c_413_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_Y_c_414_n 0.00287885f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.335
cc_37 VNB N_VPWR_c_512_n 0.183584f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_38 VNB N_VGND_c_559_n 0.00830622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_560_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.41
cc_40 VNB N_VGND_c_561_n 0.017069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_562_n 0.0186436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_563_n 0.0291174f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.65
cc_43 VNB N_VGND_c_564_n 0.262723f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.665
cc_44 VNB N_VGND_c_565_n 0.0187181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_566_n 0.0328803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_567_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_568_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VPB N_C_M1001_g 0.0270589f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_49 VPB N_C_M1008_g 0.0238365f $X=-0.19 $Y=1.66 $X2=1.895 $Y2=2.4
cc_50 VPB C 0.00281955f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.665
cc_51 VPB N_D_M1004_g 0.0193942f $X=-0.19 $Y=1.66 $X2=1.895 $Y2=1.65
cc_52 VPB N_D_c_154_n 0.0021862f $X=-0.19 $Y=1.66 $X2=1.93 $Y2=1.32
cc_53 VPB N_D_M1006_g 0.0224353f $X=-0.19 $Y=1.66 $X2=1.93 $Y2=0.74
cc_54 VPB N_B_M1003_g 0.0238907f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_55 VPB N_B_M1011_g 0.0275465f $X=-0.19 $Y=1.66 $X2=1.93 $Y2=0.74
cc_56 VPB N_B_c_218_n 0.0102383f $X=-0.19 $Y=1.66 $X2=1.565 $Y2=1.41
cc_57 VPB N_B_c_211_n 4.90622e-19 $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.335
cc_58 VPB N_B_c_214_n 0.00182616f $X=-0.19 $Y=1.66 $X2=1.91 $Y2=1.485
cc_59 VPB N_B_c_221_n 0.00766629f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_M1007_g 0.0220181f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_61 VPB N_A_M1010_g 0.0209988f $X=-0.19 $Y=1.66 $X2=1.93 $Y2=0.74
cc_62 VPB N_A_27_368#_c_331_n 0.021397f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_27_368#_c_332_n 0.00253248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_27_368#_c_333_n 0.00718969f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.95
cc_65 VPB N_A_27_368#_c_334_n 0.030619f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_27_368#_c_335_n 0.0184043f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_27_368#_c_336_n 0.0041877f $X=-0.19 $Y=1.66 $X2=1.91 $Y2=1.32
cc_68 VPB N_A_119_368#_c_393_n 0.00720268f $X=-0.19 $Y=1.66 $X2=1.93 $Y2=0.74
cc_69 VPB N_Y_c_408_n 4.44592e-19 $X=-0.19 $Y=1.66 $X2=1.93 $Y2=0.74
cc_70 VPB N_Y_c_416_n 0.00926672f $X=-0.19 $Y=1.66 $X2=0.562 $Y2=1.335
cc_71 VPB Y 0.0045771f $X=-0.19 $Y=1.66 $X2=1.91 $Y2=1.32
cc_72 VPB N_Y_c_418_n 0.00397817f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.665
cc_73 VPB N_A_493_368#_c_484_n 0.00210821f $X=-0.19 $Y=1.66 $X2=1.565 $Y2=1.41
cc_74 VPB N_A_493_368#_c_485_n 0.00371622f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.335
cc_75 VPB N_VPWR_c_513_n 0.00396467f $X=-0.19 $Y=1.66 $X2=1.895 $Y2=2.4
cc_76 VPB N_VPWR_c_514_n 0.0801244f $X=-0.19 $Y=1.66 $X2=1.93 $Y2=0.74
cc_77 VPB N_VPWR_c_515_n 0.0302153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_512_n 0.0656222f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_79 VPB N_VPWR_c_517_n 0.00601668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 N_C_c_88_n N_D_c_152_n 0.00105479f $X=1.565 $Y=1.485 $X2=-0.19 $Y2=-0.245
cc_81 N_C_c_83_n N_D_c_153_n 0.00113177f $X=0.535 $Y=1.335 $X2=0 $Y2=0
cc_82 N_C_c_84_n N_D_c_153_n 0.0222163f $X=0.535 $Y=1.335 $X2=0 $Y2=0
cc_83 N_C_M1001_g N_D_c_154_n 0.0528863f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_84 N_C_c_85_n N_D_c_154_n 0.0207003f $X=1.91 $Y=1.485 $X2=0 $Y2=0
cc_85 N_C_c_86_n N_D_c_154_n 0.00443665f $X=1.91 $Y=1.485 $X2=0 $Y2=0
cc_86 N_C_c_88_n N_D_c_154_n 0.0379444f $X=1.565 $Y=1.485 $X2=0 $Y2=0
cc_87 N_C_M1008_g N_D_M1006_g 0.0469122f $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_88 C N_D_M1006_g 0.00324652f $X=1.68 $Y=1.665 $X2=0 $Y2=0
cc_89 N_C_M1002_g N_D_c_156_n 0.0162664f $X=1.93 $Y=0.74 $X2=0 $Y2=0
cc_90 N_C_c_83_n N_D_c_158_n 2.88011e-19 $X=0.535 $Y=1.335 $X2=0 $Y2=0
cc_91 N_C_c_84_n N_D_c_158_n 0.0145155f $X=0.535 $Y=1.335 $X2=0 $Y2=0
cc_92 N_C_M1008_g N_B_M1003_g 0.0149348f $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_93 N_C_M1002_g N_B_M1009_g 0.0254515f $X=1.93 $Y=0.74 $X2=0 $Y2=0
cc_94 N_C_M1008_g N_B_c_211_n 5.10653e-19 $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_95 N_C_c_85_n N_B_c_211_n 4.14781e-19 $X=1.91 $Y=1.485 $X2=0 $Y2=0
cc_96 N_C_c_86_n N_B_c_211_n 0.0220044f $X=1.91 $Y=1.485 $X2=0 $Y2=0
cc_97 C N_B_c_211_n 0.00468098f $X=1.68 $Y=1.665 $X2=0 $Y2=0
cc_98 N_C_c_85_n N_B_c_212_n 0.0214219f $X=1.91 $Y=1.485 $X2=0 $Y2=0
cc_99 N_C_c_86_n N_B_c_212_n 4.11724e-19 $X=1.91 $Y=1.485 $X2=0 $Y2=0
cc_100 N_C_M1001_g N_A_27_368#_c_331_n 0.00132054f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_101 N_C_M1001_g N_A_27_368#_c_338_n 0.0117118f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_102 N_C_M1008_g N_A_27_368#_c_338_n 0.0137577f $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_103 N_C_c_86_n N_A_27_368#_c_338_n 0.00481713f $X=1.91 $Y=1.485 $X2=0 $Y2=0
cc_104 C N_A_27_368#_c_338_n 0.0123798f $X=1.68 $Y=1.665 $X2=0 $Y2=0
cc_105 N_C_M1008_g N_A_27_368#_c_332_n 2.97279e-19 $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_106 N_C_M1001_g N_A_27_368#_c_335_n 0.00695575f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_107 N_C_M1008_g N_A_27_368#_c_336_n 2.91527e-19 $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_108 N_C_c_85_n N_A_27_368#_c_336_n 9.08531e-19 $X=1.91 $Y=1.485 $X2=0 $Y2=0
cc_109 N_C_c_86_n N_A_27_368#_c_336_n 0.003289f $X=1.91 $Y=1.485 $X2=0 $Y2=0
cc_110 C N_A_27_368#_c_336_n 0.00118327f $X=1.68 $Y=1.665 $X2=0 $Y2=0
cc_111 C N_A_119_368#_M1006_s 0.00431345f $X=1.68 $Y=1.665 $X2=0 $Y2=0
cc_112 N_C_M1001_g N_A_119_368#_c_393_n 0.00516813f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_113 N_C_M1008_g N_A_119_368#_c_393_n 0.00472091f $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_114 N_C_M1001_g N_Y_c_408_n 0.0059715f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_115 N_C_c_83_n N_Y_c_408_n 0.0244588f $X=0.535 $Y=1.335 $X2=0 $Y2=0
cc_116 N_C_c_84_n N_Y_c_408_n 0.00789454f $X=0.535 $Y=1.335 $X2=0 $Y2=0
cc_117 N_C_c_83_n N_Y_c_409_n 0.0206189f $X=0.535 $Y=1.335 $X2=0 $Y2=0
cc_118 N_C_c_84_n N_Y_c_409_n 0.00149408f $X=0.535 $Y=1.335 $X2=0 $Y2=0
cc_119 N_C_c_88_n N_Y_c_409_n 0.0358256f $X=1.565 $Y=1.485 $X2=0 $Y2=0
cc_120 N_C_M1002_g N_Y_c_411_n 0.00627366f $X=1.93 $Y=0.74 $X2=0 $Y2=0
cc_121 N_C_M1002_g N_Y_c_412_n 0.0123739f $X=1.93 $Y=0.74 $X2=0 $Y2=0
cc_122 N_C_c_85_n N_Y_c_412_n 0.00156944f $X=1.91 $Y=1.485 $X2=0 $Y2=0
cc_123 N_C_c_86_n N_Y_c_412_n 0.0141875f $X=1.91 $Y=1.485 $X2=0 $Y2=0
cc_124 N_C_M1002_g N_Y_c_413_n 6.22903e-19 $X=1.93 $Y=0.74 $X2=0 $Y2=0
cc_125 N_C_M1002_g N_Y_c_414_n 0.00473451f $X=1.93 $Y=0.74 $X2=0 $Y2=0
cc_126 N_C_c_85_n N_Y_c_414_n 0.00275973f $X=1.91 $Y=1.485 $X2=0 $Y2=0
cc_127 N_C_c_88_n N_Y_c_414_n 0.0282645f $X=1.565 $Y=1.485 $X2=0 $Y2=0
cc_128 C Y 0.0256087f $X=1.68 $Y=1.665 $X2=0 $Y2=0
cc_129 N_C_c_88_n Y 0.0534858f $X=1.565 $Y=1.485 $X2=0 $Y2=0
cc_130 N_C_M1001_g N_Y_c_418_n 0.0149189f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_131 N_C_c_83_n N_Y_c_418_n 0.0204894f $X=0.535 $Y=1.335 $X2=0 $Y2=0
cc_132 N_C_c_84_n N_Y_c_418_n 0.00201086f $X=0.535 $Y=1.335 $X2=0 $Y2=0
cc_133 N_C_M1001_g N_VPWR_c_514_n 0.00519794f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_134 N_C_M1008_g N_VPWR_c_514_n 0.00519794f $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_135 N_C_M1001_g N_VPWR_c_512_n 0.00537282f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_136 N_C_M1008_g N_VPWR_c_512_n 0.00535486f $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_137 N_C_M1002_g N_VGND_c_559_n 0.00466065f $X=1.93 $Y=0.74 $X2=0 $Y2=0
cc_138 N_C_M1002_g N_VGND_c_562_n 0.00434272f $X=1.93 $Y=0.74 $X2=0 $Y2=0
cc_139 N_C_M1002_g N_VGND_c_564_n 0.0082177f $X=1.93 $Y=0.74 $X2=0 $Y2=0
cc_140 N_D_M1004_g N_A_27_368#_c_338_n 0.0118607f $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_141 N_D_M1006_g N_A_27_368#_c_338_n 0.0163522f $X=1.445 $Y=2.4 $X2=0 $Y2=0
cc_142 N_D_M1004_g N_A_27_368#_c_335_n 9.81305e-19 $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_143 N_D_M1004_g N_A_119_368#_c_393_n 0.0140976f $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_144 N_D_M1006_g N_A_119_368#_c_393_n 0.0138367f $X=1.445 $Y=2.4 $X2=0 $Y2=0
cc_145 N_D_c_153_n N_Y_c_408_n 0.00351765f $X=0.985 $Y=1.185 $X2=0 $Y2=0
cc_146 N_D_c_152_n N_Y_c_409_n 0.0167197f $X=0.91 $Y=0.81 $X2=0 $Y2=0
cc_147 N_D_c_153_n N_Y_c_409_n 0.00870161f $X=0.985 $Y=1.185 $X2=0 $Y2=0
cc_148 N_D_c_154_n N_Y_c_409_n 0.00355636f $X=1.445 $Y=1.52 $X2=0 $Y2=0
cc_149 N_D_c_156_n N_Y_c_409_n 0.0109092f $X=1.46 $Y=1.185 $X2=0 $Y2=0
cc_150 D N_Y_c_409_n 0.012611f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_151 N_D_c_158_n N_Y_c_409_n 0.00582959f $X=0.27 $Y=0.495 $X2=0 $Y2=0
cc_152 D N_Y_c_410_n 0.0122776f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_153 N_D_c_158_n N_Y_c_410_n 0.0011793f $X=0.27 $Y=0.495 $X2=0 $Y2=0
cc_154 N_D_c_156_n N_Y_c_411_n 4.77705e-19 $X=1.46 $Y=1.185 $X2=0 $Y2=0
cc_155 N_D_c_156_n N_Y_c_414_n 0.00113886f $X=1.46 $Y=1.185 $X2=0 $Y2=0
cc_156 N_D_M1004_g Y 0.0163525f $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_157 N_D_c_154_n Y 0.00646722f $X=1.445 $Y=1.52 $X2=0 $Y2=0
cc_158 N_D_M1006_g Y 0.00843581f $X=1.445 $Y=2.4 $X2=0 $Y2=0
cc_159 N_D_M1004_g N_VPWR_c_514_n 0.00349978f $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_160 N_D_M1006_g N_VPWR_c_514_n 0.00349978f $X=1.445 $Y=2.4 $X2=0 $Y2=0
cc_161 N_D_M1004_g N_VPWR_c_512_n 0.0043002f $X=0.97 $Y=2.4 $X2=0 $Y2=0
cc_162 N_D_M1006_g N_VPWR_c_512_n 0.00429879f $X=1.445 $Y=2.4 $X2=0 $Y2=0
cc_163 N_D_c_156_n N_VGND_c_562_n 0.00461464f $X=1.46 $Y=1.185 $X2=0 $Y2=0
cc_164 N_D_c_152_n N_VGND_c_564_n 0.00367388f $X=0.91 $Y=0.81 $X2=0 $Y2=0
cc_165 N_D_c_156_n N_VGND_c_564_n 0.00465425f $X=1.46 $Y=1.185 $X2=0 $Y2=0
cc_166 D N_VGND_c_564_n 0.0117407f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_167 N_D_c_152_n N_VGND_c_565_n 0.00272934f $X=0.91 $Y=0.81 $X2=0 $Y2=0
cc_168 D N_VGND_c_565_n 0.01419f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_169 N_D_c_158_n N_VGND_c_565_n 0.0019148f $X=0.27 $Y=0.495 $X2=0 $Y2=0
cc_170 N_D_c_152_n N_VGND_c_566_n 0.011043f $X=0.91 $Y=0.81 $X2=0 $Y2=0
cc_171 N_D_c_156_n N_VGND_c_566_n 0.00417838f $X=1.46 $Y=1.185 $X2=0 $Y2=0
cc_172 D N_VGND_c_566_n 0.0226857f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_173 N_D_c_158_n N_VGND_c_566_n 0.00626653f $X=0.27 $Y=0.495 $X2=0 $Y2=0
cc_174 N_B_M1003_g N_A_M1007_g 0.0261847f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_175 N_B_c_218_n N_A_M1007_g 0.0165486f $X=3.885 $Y=1.795 $X2=0 $Y2=0
cc_176 N_B_M1009_g N_A_c_288_n 0.013405f $X=2.5 $Y=0.74 $X2=0 $Y2=0
cc_177 N_B_c_213_n N_A_c_288_n 0.00834965f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_178 N_B_c_218_n N_A_M1010_g 0.0116248f $X=3.885 $Y=1.795 $X2=0 $Y2=0
cc_179 N_B_c_215_n N_A_M1010_g 0.0288678f $X=4.05 $Y=1.465 $X2=0 $Y2=0
cc_180 N_B_M1009_g A 3.75378e-19 $X=2.5 $Y=0.74 $X2=0 $Y2=0
cc_181 N_B_c_218_n A 0.0473225f $X=3.885 $Y=1.795 $X2=0 $Y2=0
cc_182 N_B_c_211_n A 0.00850511f $X=2.45 $Y=1.485 $X2=0 $Y2=0
cc_183 N_B_c_213_n A 0.00384508f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_184 N_B_c_214_n A 0.0299183f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_185 N_B_M1009_g N_A_c_291_n 0.00591688f $X=2.5 $Y=0.74 $X2=0 $Y2=0
cc_186 N_B_c_218_n N_A_c_291_n 0.00204163f $X=3.885 $Y=1.795 $X2=0 $Y2=0
cc_187 N_B_c_211_n N_A_c_291_n 0.0057799f $X=2.45 $Y=1.485 $X2=0 $Y2=0
cc_188 N_B_c_212_n N_A_c_291_n 0.0211473f $X=2.45 $Y=1.485 $X2=0 $Y2=0
cc_189 N_B_c_213_n N_A_c_291_n 0.0288678f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_190 N_B_c_214_n N_A_c_291_n 0.00100972f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_191 N_B_c_221_n N_A_27_368#_M1011_s 0.00268917f $X=4.05 $Y=1.71 $X2=0 $Y2=0
cc_192 N_B_M1003_g N_A_27_368#_c_332_n 3.01943e-19 $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_193 N_B_M1003_g N_A_27_368#_c_353_n 0.0169762f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_194 N_B_M1011_g N_A_27_368#_c_353_n 0.0141725f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_195 N_B_c_218_n N_A_27_368#_c_353_n 0.0682237f $X=3.885 $Y=1.795 $X2=0 $Y2=0
cc_196 N_B_c_211_n N_A_27_368#_c_353_n 0.0150896f $X=2.45 $Y=1.485 $X2=0 $Y2=0
cc_197 N_B_c_212_n N_A_27_368#_c_353_n 5.36923e-19 $X=2.45 $Y=1.485 $X2=0 $Y2=0
cc_198 N_B_c_221_n N_A_27_368#_c_353_n 0.00144733f $X=4.05 $Y=1.71 $X2=0 $Y2=0
cc_199 N_B_c_215_n N_A_27_368#_c_333_n 0.00114697f $X=4.05 $Y=1.465 $X2=0 $Y2=0
cc_200 N_B_c_221_n N_A_27_368#_c_333_n 0.02198f $X=4.05 $Y=1.71 $X2=0 $Y2=0
cc_201 N_B_M1011_g N_A_27_368#_c_334_n 0.00639412f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_202 N_B_c_211_n N_A_27_368#_c_336_n 0.00489089f $X=2.45 $Y=1.485 $X2=0 $Y2=0
cc_203 N_B_M1009_g N_Y_c_411_n 6.27466e-19 $X=2.5 $Y=0.74 $X2=0 $Y2=0
cc_204 N_B_M1009_g N_Y_c_412_n 0.0129975f $X=2.5 $Y=0.74 $X2=0 $Y2=0
cc_205 N_B_c_218_n N_Y_c_412_n 0.00904733f $X=3.885 $Y=1.795 $X2=0 $Y2=0
cc_206 N_B_c_211_n N_Y_c_412_n 0.0263393f $X=2.45 $Y=1.485 $X2=0 $Y2=0
cc_207 N_B_c_212_n N_Y_c_412_n 0.00129034f $X=2.45 $Y=1.485 $X2=0 $Y2=0
cc_208 N_B_M1009_g N_Y_c_413_n 0.00935132f $X=2.5 $Y=0.74 $X2=0 $Y2=0
cc_209 N_B_c_218_n N_A_493_368#_M1003_d 0.00151317f $X=3.885 $Y=1.795 $X2=-0.19
+ $Y2=-0.245
cc_210 N_B_c_211_n N_A_493_368#_M1003_d 0.00113588f $X=2.45 $Y=1.485 $X2=-0.19
+ $Y2=-0.245
cc_211 N_B_c_218_n N_A_493_368#_M1010_s 0.00166235f $X=3.885 $Y=1.795 $X2=0
+ $Y2=0
cc_212 N_B_M1011_g N_A_493_368#_c_489_n 0.00247387f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_213 N_B_M1011_g N_A_493_368#_c_484_n 0.0065402f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_214 N_B_M1003_g N_A_493_368#_c_485_n 7.9554e-19 $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_215 N_B_c_218_n N_VPWR_M1007_d 0.00166235f $X=3.885 $Y=1.795 $X2=-0.19
+ $Y2=-0.245
cc_216 N_B_M1003_g N_VPWR_c_513_n 4.8273e-19 $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_217 N_B_M1011_g N_VPWR_c_513_n 5.44165e-19 $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_218 N_B_M1003_g N_VPWR_c_514_n 0.00553757f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_219 N_B_M1011_g N_VPWR_c_515_n 0.00520371f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_220 N_B_M1003_g N_VPWR_c_512_n 0.0109105f $X=2.375 $Y=2.4 $X2=0 $Y2=0
cc_221 N_B_M1011_g N_VPWR_c_512_n 0.00986846f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_222 N_B_M1009_g N_VGND_c_559_n 0.00466189f $X=2.5 $Y=0.74 $X2=0 $Y2=0
cc_223 N_B_M1009_g N_VGND_c_560_n 0.00434272f $X=2.5 $Y=0.74 $X2=0 $Y2=0
cc_224 N_B_c_213_n N_VGND_c_561_n 0.00867528f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_225 N_B_c_214_n N_VGND_c_561_n 0.0255316f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_226 N_B_c_213_n N_VGND_c_563_n 0.00793088f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_227 N_B_c_214_n N_VGND_c_563_n 0.0191905f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_228 N_B_M1009_g N_VGND_c_564_n 0.0082141f $X=2.5 $Y=0.74 $X2=0 $Y2=0
cc_229 N_B_c_213_n N_VGND_c_564_n 0.00575727f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_230 N_B_c_214_n N_VGND_c_564_n 0.012382f $X=4.05 $Y=0.445 $X2=0 $Y2=0
cc_231 N_A_M1007_g N_A_27_368#_c_353_n 0.0121142f $X=2.915 $Y=2.4 $X2=0 $Y2=0
cc_232 N_A_M1010_g N_A_27_368#_c_353_n 0.0116248f $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_233 N_A_c_288_n N_Y_c_412_n 0.00807097f $X=2.93 $Y=1.22 $X2=0 $Y2=0
cc_234 N_A_c_291_n N_Y_c_412_n 0.00112261f $X=3.365 $Y=1.385 $X2=0 $Y2=0
cc_235 N_A_c_288_n N_Y_c_413_n 0.00786622f $X=2.93 $Y=1.22 $X2=0 $Y2=0
cc_236 N_A_M1007_g N_A_493_368#_c_492_n 0.0108426f $X=2.915 $Y=2.4 $X2=0 $Y2=0
cc_237 N_A_M1010_g N_A_493_368#_c_492_n 0.0108426f $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_238 N_A_M1010_g N_A_493_368#_c_484_n 3.10483e-19 $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_239 N_A_M1007_g N_A_493_368#_c_485_n 3.70456e-19 $X=2.915 $Y=2.4 $X2=0 $Y2=0
cc_240 N_A_M1007_g N_VPWR_c_513_n 0.00741359f $X=2.915 $Y=2.4 $X2=0 $Y2=0
cc_241 N_A_M1010_g N_VPWR_c_513_n 0.00744566f $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_242 N_A_M1007_g N_VPWR_c_514_n 0.00460063f $X=2.915 $Y=2.4 $X2=0 $Y2=0
cc_243 N_A_M1010_g N_VPWR_c_515_n 0.00460063f $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_244 N_A_M1007_g N_VPWR_c_512_n 0.00444149f $X=2.915 $Y=2.4 $X2=0 $Y2=0
cc_245 N_A_M1010_g N_VPWR_c_512_n 0.00443357f $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_246 N_A_c_288_n N_VGND_c_560_n 0.00434272f $X=2.93 $Y=1.22 $X2=0 $Y2=0
cc_247 N_A_c_288_n N_VGND_c_561_n 0.00279441f $X=2.93 $Y=1.22 $X2=0 $Y2=0
cc_248 A N_VGND_c_561_n 0.0248105f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_249 N_A_c_291_n N_VGND_c_561_n 0.00378911f $X=3.365 $Y=1.385 $X2=0 $Y2=0
cc_250 N_A_c_288_n N_VGND_c_564_n 0.00825157f $X=2.93 $Y=1.22 $X2=0 $Y2=0
cc_251 N_A_27_368#_c_338_n N_A_119_368#_M1001_d 0.0036196f $X=2.035 $Y=2.405
+ $X2=-0.19 $Y2=1.66
cc_252 N_A_27_368#_c_338_n N_A_119_368#_M1006_s 0.00326616f $X=2.035 $Y=2.405
+ $X2=0 $Y2=0
cc_253 N_A_27_368#_c_331_n N_A_119_368#_c_393_n 0.0123956f $X=0.28 $Y=2.495
+ $X2=0 $Y2=0
cc_254 N_A_27_368#_c_338_n N_A_119_368#_c_393_n 0.0668733f $X=2.035 $Y=2.405
+ $X2=0 $Y2=0
cc_255 N_A_27_368#_c_332_n N_A_119_368#_c_393_n 0.0123955f $X=2.12 $Y=2.815
+ $X2=0 $Y2=0
cc_256 N_A_27_368#_c_338_n N_Y_M1004_d 0.00383128f $X=2.035 $Y=2.405 $X2=0 $Y2=0
cc_257 N_A_27_368#_M1001_s N_Y_c_416_n 0.00132795f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_258 N_A_27_368#_c_335_n N_Y_c_416_n 0.0125997f $X=0.28 $Y=2.155 $X2=0 $Y2=0
cc_259 N_A_27_368#_c_336_n N_Y_c_412_n 0.00675162f $X=2.12 $Y=1.985 $X2=0 $Y2=0
cc_260 N_A_27_368#_c_338_n Y 0.0430934f $X=2.035 $Y=2.405 $X2=0 $Y2=0
cc_261 N_A_27_368#_c_338_n N_Y_c_418_n 0.00472017f $X=2.035 $Y=2.405 $X2=0 $Y2=0
cc_262 N_A_27_368#_c_335_n N_Y_c_418_n 0.0127403f $X=0.28 $Y=2.155 $X2=0 $Y2=0
cc_263 N_A_27_368#_c_353_n N_A_493_368#_M1003_d 0.00509402f $X=3.94 $Y=2.135
+ $X2=-0.19 $Y2=1.66
cc_264 N_A_27_368#_c_353_n N_A_493_368#_M1010_s 0.00332066f $X=3.94 $Y=2.135
+ $X2=0 $Y2=0
cc_265 N_A_27_368#_c_353_n N_A_493_368#_c_492_n 0.0356639f $X=3.94 $Y=2.135
+ $X2=0 $Y2=0
cc_266 N_A_27_368#_c_353_n N_A_493_368#_c_489_n 0.0148038f $X=3.94 $Y=2.135
+ $X2=0 $Y2=0
cc_267 N_A_27_368#_c_334_n N_A_493_368#_c_484_n 0.0148001f $X=4.04 $Y=2.815
+ $X2=0 $Y2=0
cc_268 N_A_27_368#_c_332_n N_A_493_368#_c_485_n 0.0152623f $X=2.12 $Y=2.815
+ $X2=0 $Y2=0
cc_269 N_A_27_368#_c_353_n N_A_493_368#_c_485_n 0.0198377f $X=3.94 $Y=2.135
+ $X2=0 $Y2=0
cc_270 N_A_27_368#_c_353_n N_VPWR_M1007_d 0.003218f $X=3.94 $Y=2.135 $X2=-0.19
+ $Y2=1.66
cc_271 N_A_27_368#_c_331_n N_VPWR_c_514_n 0.0120294f $X=0.28 $Y=2.495 $X2=0
+ $Y2=0
cc_272 N_A_27_368#_c_332_n N_VPWR_c_514_n 0.011066f $X=2.12 $Y=2.815 $X2=0 $Y2=0
cc_273 N_A_27_368#_c_334_n N_VPWR_c_515_n 0.0117353f $X=4.04 $Y=2.815 $X2=0
+ $Y2=0
cc_274 N_A_27_368#_c_331_n N_VPWR_c_512_n 0.00926813f $X=0.28 $Y=2.495 $X2=0
+ $Y2=0
cc_275 N_A_27_368#_c_338_n N_VPWR_c_512_n 0.0107436f $X=2.035 $Y=2.405 $X2=0
+ $Y2=0
cc_276 N_A_27_368#_c_332_n N_VPWR_c_512_n 0.00915947f $X=2.12 $Y=2.815 $X2=0
+ $Y2=0
cc_277 N_A_27_368#_c_334_n N_VPWR_c_512_n 0.00971347f $X=4.04 $Y=2.815 $X2=0
+ $Y2=0
cc_278 N_A_27_368#_c_335_n N_VPWR_c_512_n 0.00275594f $X=0.28 $Y=2.155 $X2=0
+ $Y2=0
cc_279 N_A_119_368#_c_393_n N_Y_M1004_d 0.00196669f $X=1.67 $Y=2.78 $X2=0 $Y2=0
cc_280 N_A_119_368#_M1001_d Y 0.00220542f $X=0.595 $Y=1.84 $X2=0 $Y2=0
cc_281 N_A_119_368#_c_393_n N_VPWR_c_514_n 0.0523508f $X=1.67 $Y=2.78 $X2=0
+ $Y2=0
cc_282 N_A_119_368#_c_393_n N_VPWR_c_512_n 0.0437259f $X=1.67 $Y=2.78 $X2=0
+ $Y2=0
cc_283 N_Y_c_409_n N_VGND_M1005_s 0.0045742f $X=1.55 $Y=0.915 $X2=-0.19
+ $Y2=-0.245
cc_284 N_Y_c_412_n N_VGND_M1002_d 0.00368125f $X=2.55 $Y=1.065 $X2=0 $Y2=0
cc_285 N_Y_c_411_n N_VGND_c_559_n 0.0180508f $X=1.715 $Y=0.515 $X2=0 $Y2=0
cc_286 N_Y_c_412_n N_VGND_c_559_n 0.0248957f $X=2.55 $Y=1.065 $X2=0 $Y2=0
cc_287 N_Y_c_413_n N_VGND_c_559_n 0.0180508f $X=2.715 $Y=0.515 $X2=0 $Y2=0
cc_288 N_Y_c_413_n N_VGND_c_560_n 0.0144922f $X=2.715 $Y=0.515 $X2=0 $Y2=0
cc_289 N_Y_c_413_n N_VGND_c_561_n 0.0243921f $X=2.715 $Y=0.515 $X2=0 $Y2=0
cc_290 N_Y_c_411_n N_VGND_c_562_n 0.0145639f $X=1.715 $Y=0.515 $X2=0 $Y2=0
cc_291 N_Y_c_409_n N_VGND_c_564_n 0.0130841f $X=1.55 $Y=0.915 $X2=0 $Y2=0
cc_292 N_Y_c_410_n N_VGND_c_564_n 0.00111297f $X=0.255 $Y=0.915 $X2=0 $Y2=0
cc_293 N_Y_c_411_n N_VGND_c_564_n 0.0119984f $X=1.715 $Y=0.515 $X2=0 $Y2=0
cc_294 N_Y_c_413_n N_VGND_c_564_n 0.0118826f $X=2.715 $Y=0.515 $X2=0 $Y2=0
cc_295 N_Y_c_409_n N_VGND_c_566_n 0.0436524f $X=1.55 $Y=0.915 $X2=0 $Y2=0
cc_296 N_Y_c_411_n N_VGND_c_566_n 0.00167954f $X=1.715 $Y=0.515 $X2=0 $Y2=0
cc_297 N_A_493_368#_c_492_n N_VPWR_M1007_d 0.00328796f $X=3.505 $Y=2.475
+ $X2=-0.19 $Y2=1.66
cc_298 N_A_493_368#_c_492_n N_VPWR_c_513_n 0.0165487f $X=3.505 $Y=2.475 $X2=0
+ $Y2=0
cc_299 N_A_493_368#_c_484_n N_VPWR_c_513_n 0.0102829f $X=3.59 $Y=2.835 $X2=0
+ $Y2=0
cc_300 N_A_493_368#_c_485_n N_VPWR_c_513_n 0.0117536f $X=2.64 $Y=2.495 $X2=0
+ $Y2=0
cc_301 N_A_493_368#_c_485_n N_VPWR_c_514_n 0.0157837f $X=2.64 $Y=2.495 $X2=0
+ $Y2=0
cc_302 N_A_493_368#_c_484_n N_VPWR_c_515_n 0.0118457f $X=3.59 $Y=2.835 $X2=0
+ $Y2=0
cc_303 N_A_493_368#_c_492_n N_VPWR_c_512_n 0.0125347f $X=3.505 $Y=2.475 $X2=0
+ $Y2=0
cc_304 N_A_493_368#_c_484_n N_VPWR_c_512_n 0.00909694f $X=3.59 $Y=2.835 $X2=0
+ $Y2=0
cc_305 N_A_493_368#_c_485_n N_VPWR_c_512_n 0.0122146f $X=2.64 $Y=2.495 $X2=0
+ $Y2=0

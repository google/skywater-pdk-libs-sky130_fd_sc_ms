* File: sky130_fd_sc_ms__sdfrtp_1.pxi.spice
* Created: Wed Sep  2 12:30:33 2020
* 
x_PM_SKY130_FD_SC_MS__SDFRTP_1%SCE N_SCE_M1005_g N_SCE_M1034_g N_SCE_M1002_g
+ N_SCE_M1025_g N_SCE_c_285_n N_SCE_c_286_n N_SCE_c_287_n N_SCE_c_288_n
+ N_SCE_c_289_n SCE SCE SCE N_SCE_c_290_n N_SCE_c_291_n N_SCE_c_292_n SCE
+ N_SCE_c_298_n PM_SKY130_FD_SC_MS__SDFRTP_1%SCE
x_PM_SKY130_FD_SC_MS__SDFRTP_1%A_27_88# N_A_27_88#_M1034_s N_A_27_88#_M1005_s
+ N_A_27_88#_c_374_n N_A_27_88#_M1008_g N_A_27_88#_c_381_n N_A_27_88#_M1016_g
+ N_A_27_88#_c_375_n N_A_27_88#_c_376_n N_A_27_88#_c_384_n N_A_27_88#_c_377_n
+ N_A_27_88#_c_385_n N_A_27_88#_c_386_n N_A_27_88#_c_387_n N_A_27_88#_c_378_n
+ N_A_27_88#_c_388_n N_A_27_88#_c_379_n N_A_27_88#_c_380_n N_A_27_88#_c_389_n
+ PM_SKY130_FD_SC_MS__SDFRTP_1%A_27_88#
x_PM_SKY130_FD_SC_MS__SDFRTP_1%D N_D_c_462_n N_D_M1013_g N_D_c_456_n N_D_c_457_n
+ N_D_M1009_g N_D_c_464_n N_D_c_458_n D N_D_c_459_n N_D_c_460_n N_D_c_461_n
+ PM_SKY130_FD_SC_MS__SDFRTP_1%D
x_PM_SKY130_FD_SC_MS__SDFRTP_1%SCD N_SCD_M1019_g N_SCD_M1015_g N_SCD_c_513_n
+ N_SCD_c_517_n SCD SCD N_SCD_c_515_n PM_SKY130_FD_SC_MS__SDFRTP_1%SCD
x_PM_SKY130_FD_SC_MS__SDFRTP_1%CLK N_CLK_c_553_n N_CLK_M1029_g N_CLK_c_556_n
+ N_CLK_M1018_g CLK PM_SKY130_FD_SC_MS__SDFRTP_1%CLK
x_PM_SKY130_FD_SC_MS__SDFRTP_1%A_1037_387# N_A_1037_387#_M1032_d
+ N_A_1037_387#_M1030_d N_A_1037_387#_M1000_g N_A_1037_387#_c_609_n
+ N_A_1037_387#_M1001_g N_A_1037_387#_c_611_n N_A_1037_387#_M1006_g
+ N_A_1037_387#_c_612_n N_A_1037_387#_M1014_g N_A_1037_387#_c_613_n
+ N_A_1037_387#_c_614_n N_A_1037_387#_c_615_n N_A_1037_387#_c_616_n
+ N_A_1037_387#_c_631_n N_A_1037_387#_c_617_n N_A_1037_387#_c_618_n
+ N_A_1037_387#_c_619_n N_A_1037_387#_c_643_p N_A_1037_387#_c_669_p
+ N_A_1037_387#_c_620_n N_A_1037_387#_c_621_n N_A_1037_387#_c_622_n
+ N_A_1037_387#_c_623_n N_A_1037_387#_c_740_p N_A_1037_387#_c_634_n
+ N_A_1037_387#_c_624_n N_A_1037_387#_c_625_n N_A_1037_387#_c_626_n
+ N_A_1037_387#_c_627_n N_A_1037_387#_c_628_n N_A_1037_387#_c_636_n
+ PM_SKY130_FD_SC_MS__SDFRTP_1%A_1037_387#
x_PM_SKY130_FD_SC_MS__SDFRTP_1%A_1367_93# N_A_1367_93#_M1033_d
+ N_A_1367_93#_M1026_d N_A_1367_93#_M1020_g N_A_1367_93#_M1028_g
+ N_A_1367_93#_c_818_n N_A_1367_93#_c_819_n N_A_1367_93#_c_820_n
+ N_A_1367_93#_c_821_n N_A_1367_93#_c_827_n N_A_1367_93#_c_828_n
+ N_A_1367_93#_c_822_n N_A_1367_93#_c_823_n
+ PM_SKY130_FD_SC_MS__SDFRTP_1%A_1367_93#
x_PM_SKY130_FD_SC_MS__SDFRTP_1%RESET_B N_RESET_B_M1036_g N_RESET_B_M1023_g
+ N_RESET_B_c_922_n N_RESET_B_c_923_n N_RESET_B_c_932_n N_RESET_B_c_933_n
+ N_RESET_B_M1012_g N_RESET_B_c_925_n N_RESET_B_c_926_n N_RESET_B_c_927_n
+ N_RESET_B_M1010_g N_RESET_B_M1038_g N_RESET_B_c_929_n N_RESET_B_M1021_g
+ N_RESET_B_c_938_n N_RESET_B_c_930_n N_RESET_B_c_939_n N_RESET_B_c_940_n
+ N_RESET_B_c_941_n N_RESET_B_c_942_n N_RESET_B_c_943_n RESET_B
+ N_RESET_B_c_945_n N_RESET_B_c_946_n N_RESET_B_c_947_n N_RESET_B_c_948_n
+ PM_SKY130_FD_SC_MS__SDFRTP_1%RESET_B
x_PM_SKY130_FD_SC_MS__SDFRTP_1%A_1234_119# N_A_1234_119#_M1035_d
+ N_A_1234_119#_M1000_d N_A_1234_119#_M1010_d N_A_1234_119#_M1033_g
+ N_A_1234_119#_c_1147_n N_A_1234_119#_M1026_g N_A_1234_119#_c_1157_n
+ N_A_1234_119#_c_1148_n N_A_1234_119#_c_1149_n N_A_1234_119#_c_1190_n
+ N_A_1234_119#_c_1150_n N_A_1234_119#_c_1151_n N_A_1234_119#_c_1152_n
+ N_A_1234_119#_c_1153_n N_A_1234_119#_c_1154_n N_A_1234_119#_c_1161_n
+ PM_SKY130_FD_SC_MS__SDFRTP_1%A_1234_119#
x_PM_SKY130_FD_SC_MS__SDFRTP_1%A_835_93# N_A_835_93#_M1029_s N_A_835_93#_M1018_s
+ N_A_835_93#_c_1287_n N_A_835_93#_M1030_g N_A_835_93#_c_1275_n
+ N_A_835_93#_M1032_g N_A_835_93#_c_1288_n N_A_835_93#_c_1289_n
+ N_A_835_93#_c_1290_n N_A_835_93#_c_1276_n N_A_835_93#_c_1277_n
+ N_A_835_93#_M1035_g N_A_835_93#_M1017_g N_A_835_93#_c_1293_n
+ N_A_835_93#_M1031_g N_A_835_93#_c_1279_n N_A_835_93#_c_1280_n
+ N_A_835_93#_c_1281_n N_A_835_93#_M1004_g N_A_835_93#_c_1297_n
+ N_A_835_93#_c_1283_n N_A_835_93#_c_1305_n N_A_835_93#_c_1306_n
+ N_A_835_93#_c_1308_n N_A_835_93#_c_1310_n N_A_835_93#_c_1284_n
+ N_A_835_93#_c_1298_n N_A_835_93#_c_1285_n N_A_835_93#_c_1317_n
+ N_A_835_93#_c_1286_n PM_SKY130_FD_SC_MS__SDFRTP_1%A_835_93#
x_PM_SKY130_FD_SC_MS__SDFRTP_1%A_1997_272# N_A_1997_272#_M1022_d
+ N_A_1997_272#_M1021_d N_A_1997_272#_M1003_g N_A_1997_272#_c_1465_n
+ N_A_1997_272#_M1037_g N_A_1997_272#_c_1466_n N_A_1997_272#_c_1467_n
+ N_A_1997_272#_c_1468_n N_A_1997_272#_c_1469_n N_A_1997_272#_c_1470_n
+ N_A_1997_272#_c_1471_n N_A_1997_272#_c_1472_n N_A_1997_272#_c_1477_n
+ N_A_1997_272#_c_1473_n N_A_1997_272#_c_1474_n
+ PM_SKY130_FD_SC_MS__SDFRTP_1%A_1997_272#
x_PM_SKY130_FD_SC_MS__SDFRTP_1%A_1745_74# N_A_1745_74#_M1006_d
+ N_A_1745_74#_M1031_d N_A_1745_74#_M1022_g N_A_1745_74#_c_1575_n
+ N_A_1745_74#_M1024_g N_A_1745_74#_c_1576_n N_A_1745_74#_c_1577_n
+ N_A_1745_74#_c_1587_n N_A_1745_74#_M1039_g N_A_1745_74#_M1027_g
+ N_A_1745_74#_c_1589_n N_A_1745_74#_c_1590_n N_A_1745_74#_c_1579_n
+ N_A_1745_74#_c_1580_n N_A_1745_74#_c_1592_n N_A_1745_74#_c_1593_n
+ N_A_1745_74#_c_1594_n N_A_1745_74#_c_1581_n N_A_1745_74#_c_1582_n
+ N_A_1745_74#_c_1583_n N_A_1745_74#_c_1584_n
+ PM_SKY130_FD_SC_MS__SDFRTP_1%A_1745_74#
x_PM_SKY130_FD_SC_MS__SDFRTP_1%A_2402_424# N_A_2402_424#_M1027_d
+ N_A_2402_424#_M1039_d N_A_2402_424#_M1011_g N_A_2402_424#_M1007_g
+ N_A_2402_424#_c_1733_n N_A_2402_424#_c_1734_n N_A_2402_424#_c_1739_n
+ N_A_2402_424#_c_1735_n N_A_2402_424#_c_1757_p N_A_2402_424#_c_1736_n
+ N_A_2402_424#_c_1737_n PM_SKY130_FD_SC_MS__SDFRTP_1%A_2402_424#
x_PM_SKY130_FD_SC_MS__SDFRTP_1%VPWR N_VPWR_M1005_d N_VPWR_M1019_d N_VPWR_M1018_d
+ N_VPWR_M1028_d N_VPWR_M1026_s N_VPWR_M1037_d N_VPWR_M1024_d N_VPWR_M1011_s
+ N_VPWR_c_1777_n N_VPWR_c_1778_n N_VPWR_c_1779_n N_VPWR_c_1780_n
+ N_VPWR_c_1781_n N_VPWR_c_1782_n N_VPWR_c_1783_n N_VPWR_c_1784_n
+ N_VPWR_c_1785_n N_VPWR_c_1786_n N_VPWR_c_1787_n N_VPWR_c_1788_n
+ N_VPWR_c_1789_n N_VPWR_c_1790_n N_VPWR_c_1791_n VPWR N_VPWR_c_1792_n
+ N_VPWR_c_1793_n N_VPWR_c_1794_n N_VPWR_c_1795_n N_VPWR_c_1796_n
+ N_VPWR_c_1776_n N_VPWR_c_1798_n N_VPWR_c_1799_n N_VPWR_c_1800_n
+ N_VPWR_c_1801_n N_VPWR_c_1802_n PM_SKY130_FD_SC_MS__SDFRTP_1%VPWR
x_PM_SKY130_FD_SC_MS__SDFRTP_1%A_303_464# N_A_303_464#_M1009_d
+ N_A_303_464#_M1035_s N_A_303_464#_M1013_d N_A_303_464#_M1023_d
+ N_A_303_464#_M1000_s N_A_303_464#_c_1946_n N_A_303_464#_c_1968_n
+ N_A_303_464#_c_1937_n N_A_303_464#_c_1938_n N_A_303_464#_c_1948_n
+ N_A_303_464#_c_1949_n N_A_303_464#_c_1939_n N_A_303_464#_c_1940_n
+ N_A_303_464#_c_1950_n N_A_303_464#_c_1941_n N_A_303_464#_c_1942_n
+ N_A_303_464#_c_1951_n N_A_303_464#_c_1952_n N_A_303_464#_c_1943_n
+ N_A_303_464#_c_1954_n N_A_303_464#_c_1944_n N_A_303_464#_c_1955_n
+ N_A_303_464#_c_1945_n PM_SKY130_FD_SC_MS__SDFRTP_1%A_303_464#
x_PM_SKY130_FD_SC_MS__SDFRTP_1%Q N_Q_M1007_d N_Q_M1011_d Q Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_MS__SDFRTP_1%Q
x_PM_SKY130_FD_SC_MS__SDFRTP_1%VGND N_VGND_M1034_d N_VGND_M1036_d N_VGND_M1029_d
+ N_VGND_M1012_d N_VGND_M1003_d N_VGND_M1027_s N_VGND_M1007_s N_VGND_c_2120_n
+ N_VGND_c_2121_n N_VGND_c_2122_n N_VGND_c_2123_n N_VGND_c_2124_n
+ N_VGND_c_2125_n N_VGND_c_2126_n N_VGND_c_2127_n VGND N_VGND_c_2128_n
+ N_VGND_c_2129_n N_VGND_c_2130_n N_VGND_c_2131_n N_VGND_c_2132_n
+ N_VGND_c_2133_n N_VGND_c_2134_n N_VGND_c_2135_n N_VGND_c_2136_n
+ N_VGND_c_2137_n N_VGND_c_2138_n N_VGND_c_2139_n N_VGND_c_2140_n
+ N_VGND_c_2141_n PM_SKY130_FD_SC_MS__SDFRTP_1%VGND
x_PM_SKY130_FD_SC_MS__SDFRTP_1%noxref_24 N_noxref_24_M1008_s N_noxref_24_M1015_d
+ N_noxref_24_c_2252_n N_noxref_24_c_2253_n N_noxref_24_c_2254_n
+ PM_SKY130_FD_SC_MS__SDFRTP_1%noxref_24
cc_1 VNB N_SCE_M1034_g 0.062352f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.65
cc_2 VNB N_SCE_c_285_n 0.0148916f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=0.9
cc_3 VNB N_SCE_c_286_n 0.0107474f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=1.05
cc_4 VNB N_SCE_c_287_n 0.0132325f $X=-0.19 $Y=-0.245 $X2=2.345 $Y2=1.575
cc_5 VNB N_SCE_c_288_n 0.00683626f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.425
cc_6 VNB N_SCE_c_289_n 0.0319913f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.425
cc_7 VNB N_SCE_c_290_n 0.0331371f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.67
cc_8 VNB N_SCE_c_291_n 0.0119307f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.26
cc_9 VNB N_SCE_c_292_n 0.0110089f $X=-0.19 $Y=-0.245 $X2=1.623 $Y2=1.662
cc_10 VNB N_A_27_88#_c_374_n 0.0192577f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.65
cc_11 VNB N_A_27_88#_c_375_n 0.0282802f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=0.9
cc_12 VNB N_A_27_88#_c_376_n 0.0187337f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.575
cc_13 VNB N_A_27_88#_c_377_n 0.0167058f $X=-0.19 $Y=-0.245 $X2=2.535 $Y2=1.575
cc_14 VNB N_A_27_88#_c_378_n 0.0130086f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.67
cc_15 VNB N_A_27_88#_c_379_n 0.00840348f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.67
cc_16 VNB N_A_27_88#_c_380_n 0.0522403f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.67
cc_17 VNB N_D_c_456_n 0.00442527f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.505
cc_18 VNB N_D_c_457_n 0.0150551f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.65
cc_19 VNB N_D_c_458_n 0.0209259f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.615
cc_20 VNB N_D_c_459_n 0.0321108f $X=-0.19 $Y=-0.245 $X2=2.535 $Y2=1.425
cc_21 VNB N_D_c_460_n 0.00935279f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.425
cc_22 VNB N_D_c_461_n 0.0161524f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.425
cc_23 VNB N_SCD_M1015_g 0.0413981f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.65
cc_24 VNB N_SCD_c_513_n 0.0128566f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.64
cc_25 VNB SCD 0.00413347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_SCD_c_515_n 0.0155097f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.615
cc_27 VNB N_CLK_c_553_n 0.0945618f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.835
cc_28 VNB CLK 0.01846f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.65
cc_29 VNB N_A_1037_387#_c_609_n 0.0238685f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.64
cc_30 VNB N_A_1037_387#_M1001_g 0.0392232f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.9
cc_31 VNB N_A_1037_387#_c_611_n 0.0161967f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.615
cc_32 VNB N_A_1037_387#_c_612_n 0.00792759f $X=-0.19 $Y=-0.245 $X2=1.795
+ $Y2=1.575
cc_33 VNB N_A_1037_387#_c_613_n 0.0105387f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_34 VNB N_A_1037_387#_c_614_n 6.30651e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_1037_387#_c_615_n 0.0379848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_1037_387#_c_616_n 0.00321642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_1037_387#_c_617_n 0.0017868f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.67
cc_38 VNB N_A_1037_387#_c_618_n 0.00375765f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=1.67
cc_39 VNB N_A_1037_387#_c_619_n 8.10761e-19 $X=-0.19 $Y=-0.245 $X2=2.51
+ $Y2=1.425
cc_40 VNB N_A_1037_387#_c_620_n 0.00889307f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=1.662
cc_41 VNB N_A_1037_387#_c_621_n 0.00224396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1037_387#_c_622_n 0.00270816f $X=-0.19 $Y=-0.245 $X2=0.96
+ $Y2=1.662
cc_43 VNB N_A_1037_387#_c_623_n 0.00419892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1037_387#_c_624_n 8.81729e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1037_387#_c_625_n 0.0363807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_1037_387#_c_626_n 0.00354363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1037_387#_c_627_n 0.0168635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1037_387#_c_628_n 0.0259737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1367_93#_M1020_g 0.0317694f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.835
cc_50 VNB N_A_1367_93#_c_818_n 0.00358202f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.615
cc_51 VNB N_A_1367_93#_c_819_n 0.0300415f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=0.9
cc_52 VNB N_A_1367_93#_c_820_n 0.00667339f $X=-0.19 $Y=-0.245 $X2=2.345
+ $Y2=1.575
cc_53 VNB N_A_1367_93#_c_821_n 4.38526e-19 $X=-0.19 $Y=-0.245 $X2=1.795
+ $Y2=1.575
cc_54 VNB N_A_1367_93#_c_822_n 0.00364646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1367_93#_c_823_n 0.00552017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_RESET_B_M1036_g 0.0600377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_RESET_B_c_922_n 0.272487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_RESET_B_c_923_n 0.012806f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.835
cc_59 VNB N_RESET_B_M1012_g 0.0265319f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.9
cc_60 VNB N_RESET_B_c_925_n 0.0260909f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.615
cc_61 VNB N_RESET_B_c_926_n 0.0069569f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.615
cc_62 VNB N_RESET_B_c_927_n 0.0202613f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=1.05
cc_63 VNB N_RESET_B_M1038_g 0.0378564f $X=-0.19 $Y=-0.245 $X2=2.535 $Y2=1.575
cc_64 VNB N_RESET_B_c_929_n 0.0109809f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_65 VNB N_RESET_B_c_930_n 0.0164222f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.67
cc_66 VNB N_A_1234_119#_M1033_g 0.0268916f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1234_119#_c_1147_n 0.0175816f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.26
cc_68 VNB N_A_1234_119#_c_1148_n 0.00374454f $X=-0.19 $Y=-0.245 $X2=2.51
+ $Y2=1.425
cc_69 VNB N_A_1234_119#_c_1149_n 0.00484689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1234_119#_c_1150_n 4.99311e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1234_119#_c_1151_n 0.00215276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1234_119#_c_1152_n 0.00602363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1234_119#_c_1153_n 0.0279564f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.67
cc_74 VNB N_A_1234_119#_c_1154_n 0.00304106f $X=-0.19 $Y=-0.245 $X2=0.96
+ $Y2=1.67
cc_75 VNB N_A_835_93#_c_1275_n 0.0155098f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.64
cc_76 VNB N_A_835_93#_c_1276_n 0.0283279f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.615
cc_77 VNB N_A_835_93#_c_1277_n 0.0620262f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=0.9
cc_78 VNB N_A_835_93#_M1035_g 0.0198814f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.575
cc_79 VNB N_A_835_93#_c_1279_n 0.0176143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_835_93#_c_1280_n 0.00502237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_835_93#_c_1281_n 0.0208108f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.67
cc_82 VNB N_A_835_93#_M1004_g 0.0235073f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.67
cc_83 VNB N_A_835_93#_c_1283_n 0.0124432f $X=-0.19 $Y=-0.245 $X2=1.623 $Y2=1.662
cc_84 VNB N_A_835_93#_c_1284_n 0.00160997f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.665
cc_85 VNB N_A_835_93#_c_1285_n 0.00359899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_835_93#_c_1286_n 0.00222099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1997_272#_M1003_g 0.0393068f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=1.835
cc_88 VNB N_A_1997_272#_c_1465_n 0.0235946f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=2.64
cc_89 VNB N_A_1997_272#_c_1466_n 0.0152817f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.9
cc_90 VNB N_A_1997_272#_c_1467_n 0.0073172f $X=-0.19 $Y=-0.245 $X2=2.625
+ $Y2=1.05
cc_91 VNB N_A_1997_272#_c_1468_n 0.00658513f $X=-0.19 $Y=-0.245 $X2=2.51
+ $Y2=1.425
cc_92 VNB N_A_1997_272#_c_1469_n 0.00719764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1997_272#_c_1470_n 0.00239418f $X=-0.19 $Y=-0.245 $X2=2.535
+ $Y2=1.575
cc_94 VNB N_A_1997_272#_c_1471_n 0.00890748f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_95 VNB N_A_1997_272#_c_1472_n 0.00132368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1997_272#_c_1473_n 4.91246e-19 $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=1.67
cc_97 VNB N_A_1997_272#_c_1474_n 6.26987e-19 $X=-0.19 $Y=-0.245 $X2=0.96
+ $Y2=1.67
cc_98 VNB N_A_1745_74#_M1022_g 0.0220606f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.835
cc_99 VNB N_A_1745_74#_c_1575_n 0.0178723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1745_74#_c_1576_n 0.0372707f $X=-0.19 $Y=-0.245 $X2=2.65
+ $Y2=0.615
cc_101 VNB N_A_1745_74#_c_1577_n 0.0476514f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=0.9
cc_102 VNB N_A_1745_74#_M1027_g 0.0313727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1745_74#_c_1579_n 0.0027518f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.67
cc_104 VNB N_A_1745_74#_c_1580_n 0.00220477f $X=-0.19 $Y=-0.245 $X2=0.96
+ $Y2=1.67
cc_105 VNB N_A_1745_74#_c_1581_n 0.00284242f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=1.662
cc_106 VNB N_A_1745_74#_c_1582_n 0.00104193f $X=-0.19 $Y=-0.245 $X2=0.96
+ $Y2=1.662
cc_107 VNB N_A_1745_74#_c_1583_n 8.69032e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_1745_74#_c_1584_n 0.0278597f $X=-0.19 $Y=-0.245 $X2=1.68
+ $Y2=1.662
cc_109 VNB N_A_2402_424#_M1011_g 0.00203363f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=1.835
cc_110 VNB N_A_2402_424#_M1007_g 0.0281108f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.05
cc_111 VNB N_A_2402_424#_c_1733_n 0.0717607f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=0.9
cc_112 VNB N_A_2402_424#_c_1734_n 0.0161946f $X=-0.19 $Y=-0.245 $X2=2.65
+ $Y2=0.615
cc_113 VNB N_A_2402_424#_c_1735_n 0.016101f $X=-0.19 $Y=-0.245 $X2=2.51
+ $Y2=1.425
cc_114 VNB N_A_2402_424#_c_1736_n 8.47259e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_2402_424#_c_1737_n 0.00458466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VPWR_c_1776_n 0.561729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_303_464#_c_1937_n 0.022757f $X=-0.19 $Y=-0.245 $X2=2.535
+ $Y2=1.425
cc_118 VNB N_A_303_464#_c_1938_n 0.00554942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_303_464#_c_1939_n 9.90482e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_303_464#_c_1940_n 0.00247329f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.67
cc_121 VNB N_A_303_464#_c_1941_n 0.00526205f $X=-0.19 $Y=-0.245 $X2=0.96
+ $Y2=1.67
cc_122 VNB N_A_303_464#_c_1942_n 0.00155211f $X=-0.19 $Y=-0.245 $X2=0.96
+ $Y2=1.67
cc_123 VNB N_A_303_464#_c_1943_n 0.00311688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_303_464#_c_1944_n 0.00434949f $X=-0.19 $Y=-0.245 $X2=0.96
+ $Y2=1.662
cc_125 VNB N_A_303_464#_c_1945_n 2.70707e-19 $X=-0.19 $Y=-0.245 $X2=1.795
+ $Y2=1.662
cc_126 VNB Q 0.0259999f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.65
cc_127 VNB Q 0.00837931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB Q 0.027119f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.835
cc_129 VNB N_VGND_c_2120_n 0.0181638f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.425
cc_130 VNB N_VGND_c_2121_n 0.0123363f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_131 VNB N_VGND_c_2122_n 0.0126479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2123_n 0.0100142f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.67
cc_133 VNB N_VGND_c_2124_n 0.00854448f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.67
cc_134 VNB N_VGND_c_2125_n 0.0169646f $X=-0.19 $Y=-0.245 $X2=1.623 $Y2=1.662
cc_135 VNB N_VGND_c_2126_n 0.021767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2127_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.662
cc_137 VNB N_VGND_c_2128_n 0.0177976f $X=-0.19 $Y=-0.245 $X2=1.609 $Y2=1.662
cc_138 VNB N_VGND_c_2129_n 0.0636435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2130_n 0.0552549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2131_n 0.0611983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2132_n 0.0297773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2133_n 0.0188435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2134_n 0.0194697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2135_n 0.704864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2136_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2137_n 0.0038619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2138_n 0.0140297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2139_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2140_n 0.00622769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2141_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_noxref_24_c_2252_n 0.0131255f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.65
cc_152 VNB N_noxref_24_c_2253_n 0.00667823f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=1.835
cc_153 VNB N_noxref_24_c_2254_n 0.00408915f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.26
cc_154 VPB N_SCE_M1005_g 0.0472519f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.64
cc_155 VPB N_SCE_M1002_g 0.0401067f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.64
cc_156 VPB N_SCE_c_288_n 0.00175837f $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.425
cc_157 VPB N_SCE_c_290_n 0.0253847f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_158 VPB N_SCE_c_292_n 0.00455267f $X=-0.19 $Y=1.66 $X2=1.623 $Y2=1.662
cc_159 VPB N_SCE_c_298_n 0.00736556f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.662
cc_160 VPB N_A_27_88#_c_381_n 0.0129195f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_27_88#_M1016_g 0.0299187f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=1.26
cc_162 VPB N_A_27_88#_c_376_n 0.0161852f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.575
cc_163 VPB N_A_27_88#_c_384_n 0.0337004f $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.425
cc_164 VPB N_A_27_88#_c_385_n 0.00159951f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_165 VPB N_A_27_88#_c_386_n 0.00570155f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_27_88#_c_387_n 0.0472568f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_27_88#_c_388_n 0.0129728f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.67
cc_168 VPB N_A_27_88#_c_389_n 0.0236923f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_D_c_462_n 0.024605f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.835
cc_170 VPB N_D_c_456_n 0.0247476f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.505
cc_171 VPB N_D_c_464_n 0.0269791f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=1.05
cc_172 VPB N_SCD_c_513_n 0.0225841f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.64
cc_173 VPB N_SCD_c_517_n 0.0321851f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.64
cc_174 VPB SCD 0.00296148f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_CLK_c_553_n 0.0169513f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.835
cc_176 VPB N_CLK_c_556_n 0.0214803f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_1037_387#_M1000_g 0.0366198f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.835
cc_178 VPB N_A_1037_387#_M1014_g 0.0248818f $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.425
cc_179 VPB N_A_1037_387#_c_631_n 0.00148328f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_1037_387#_c_617_n 0.00207438f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.67
cc_181 VPB N_A_1037_387#_c_623_n 0.00116288f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_1037_387#_c_634_n 0.00218598f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.665
cc_183 VPB N_A_1037_387#_c_627_n 0.0121291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_1037_387#_c_636_n 0.0363275f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_1367_93#_M1028_g 0.0441787f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=1.05
cc_186 VPB N_A_1367_93#_c_818_n 0.00197089f $X=-0.19 $Y=1.66 $X2=2.65 $Y2=0.615
cc_187 VPB N_A_1367_93#_c_819_n 0.0187028f $X=-0.19 $Y=1.66 $X2=2.625 $Y2=0.9
cc_188 VPB N_A_1367_93#_c_827_n 0.00177891f $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.425
cc_189 VPB N_A_1367_93#_c_828_n 0.00210098f $X=-0.19 $Y=1.66 $X2=2.535 $Y2=1.575
cc_190 VPB N_A_1367_93#_c_823_n 0.00121812f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_RESET_B_M1036_g 0.0024311f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_RESET_B_c_932_n 0.0399718f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.64
cc_193 VPB N_RESET_B_c_933_n 0.0292448f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.64
cc_194 VPB N_RESET_B_c_927_n 0.010477f $X=-0.19 $Y=1.66 $X2=2.625 $Y2=1.05
cc_195 VPB N_RESET_B_M1010_g 0.0235155f $X=-0.19 $Y=1.66 $X2=2.535 $Y2=1.425
cc_196 VPB N_RESET_B_c_929_n 0.00936563f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_197 VPB N_RESET_B_M1021_g 0.0374057f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_RESET_B_c_938_n 0.0228368f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.67
cc_199 VPB N_RESET_B_c_939_n 0.0233875f $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.425
cc_200 VPB N_RESET_B_c_940_n 0.00176136f $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.26
cc_201 VPB N_RESET_B_c_941_n 0.0217281f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_RESET_B_c_942_n 0.0020849f $X=-0.19 $Y=1.66 $X2=1.623 $Y2=1.662
cc_203 VPB N_RESET_B_c_943_n 0.00627787f $X=-0.19 $Y=1.66 $X2=1.609 $Y2=1.662
cc_204 VPB RESET_B 0.00299651f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.662
cc_205 VPB N_RESET_B_c_945_n 0.00907336f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_RESET_B_c_946_n 0.0531181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_RESET_B_c_947_n 0.00324614f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_RESET_B_c_948_n 0.0327596f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_1234_119#_c_1147_n 0.0103324f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=1.26
cc_210 VPB N_A_1234_119#_M1026_g 0.0217692f $X=-0.19 $Y=1.66 $X2=2.625 $Y2=0.9
cc_211 VPB N_A_1234_119#_c_1157_n 5.6078e-19 $X=-0.19 $Y=1.66 $X2=2.345
+ $Y2=1.575
cc_212 VPB N_A_1234_119#_c_1149_n 0.00675099f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_1234_119#_c_1150_n 0.0123477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_1234_119#_c_1153_n 0.00754174f $X=-0.19 $Y=1.66 $X2=0.495
+ $Y2=1.67
cc_215 VPB N_A_1234_119#_c_1161_n 9.35175e-19 $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.26
cc_216 VPB N_A_835_93#_c_1287_n 0.0186292f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.65
cc_217 VPB N_A_835_93#_c_1288_n 0.0723226f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=1.26
cc_218 VPB N_A_835_93#_c_1289_n 0.0591183f $X=-0.19 $Y=1.66 $X2=2.65 $Y2=0.9
cc_219 VPB N_A_835_93#_c_1290_n 0.0101558f $X=-0.19 $Y=1.66 $X2=2.65 $Y2=0.615
cc_220 VPB N_A_835_93#_c_1277_n 0.0153981f $X=-0.19 $Y=1.66 $X2=2.625 $Y2=0.9
cc_221 VPB N_A_835_93#_M1017_g 0.041698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_835_93#_c_1293_n 0.18662f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_835_93#_M1031_g 0.0287499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_835_93#_c_1279_n 0.0186371f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_835_93#_c_1280_n 0.00404075f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_835_93#_c_1297_n 0.00898883f $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.425
cc_227 VPB N_A_835_93#_c_1298_n 0.00233827f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.662
cc_228 VPB N_A_835_93#_c_1286_n 7.00034e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_1997_272#_c_1465_n 0.0211446f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.64
cc_230 VPB N_A_1997_272#_M1037_g 0.0525607f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=1.05
cc_231 VPB N_A_1997_272#_c_1477_n 0.00870521f $X=-0.19 $Y=1.66 $X2=0.495
+ $Y2=1.67
cc_232 VPB N_A_1997_272#_c_1473_n 0.00704771f $X=-0.19 $Y=1.66 $X2=0.505
+ $Y2=1.67
cc_233 VPB N_A_1745_74#_c_1575_n 0.00901615f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_1745_74#_M1024_g 0.0431356f $X=-0.19 $Y=1.66 $X2=2.65 $Y2=0.9
cc_235 VPB N_A_1745_74#_c_1587_n 0.0323038f $X=-0.19 $Y=1.66 $X2=2.625 $Y2=1.05
cc_236 VPB N_A_1745_74#_M1039_g 0.0234055f $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.425
cc_237 VPB N_A_1745_74#_c_1589_n 0.00552913f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_238 VPB N_A_1745_74#_c_1590_n 0.00177482f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_239 VPB N_A_1745_74#_c_1580_n 0.00223137f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_240 VPB N_A_1745_74#_c_1592_n 0.00730775f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.67
cc_241 VPB N_A_1745_74#_c_1593_n 0.00276148f $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.425
cc_242 VPB N_A_1745_74#_c_1594_n 0.00535671f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_2402_424#_M1011_g 0.0303184f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.835
cc_244 VPB N_A_2402_424#_c_1739_n 0.0135269f $X=-0.19 $Y=1.66 $X2=2.625 $Y2=1.05
cc_245 VPB N_A_2402_424#_c_1736_n 0.0131801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1777_n 0.00635773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1778_n 0.00645734f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1779_n 7.46595e-19 $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.67
cc_249 VPB N_VPWR_c_1780_n 0.0144177f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_250 VPB N_VPWR_c_1781_n 0.02311f $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.425
cc_251 VPB N_VPWR_c_1782_n 0.0144384f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.662
cc_252 VPB N_VPWR_c_1783_n 0.0127787f $X=-0.19 $Y=1.66 $X2=1.609 $Y2=1.662
cc_253 VPB N_VPWR_c_1784_n 0.0180602f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.662
cc_254 VPB N_VPWR_c_1785_n 0.0190424f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1786_n 0.034345f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1787_n 0.00448735f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1788_n 0.0523435f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1789_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1790_n 0.020808f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1791_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1792_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1793_n 0.0596953f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1794_n 0.0597208f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1795_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1796_n 0.0181474f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1776_n 0.120869f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1798_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1799_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1800_n 0.00443527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1801_n 0.00223798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1802_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_A_303_464#_c_1946_n 0.00657677f $X=-0.19 $Y=1.66 $X2=2.65 $Y2=0.615
cc_273 VPB N_A_303_464#_c_1938_n 0.00339097f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_A_303_464#_c_1948_n 0.0119253f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_275 VPB N_A_303_464#_c_1949_n 0.00131949f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_276 VPB N_A_303_464#_c_1950_n 0.00260011f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.67
cc_277 VPB N_A_303_464#_c_1951_n 0.00655688f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.67
cc_278 VPB N_A_303_464#_c_1952_n 0.0019149f $X=-0.19 $Y=1.66 $X2=2.51 $Y2=1.425
cc_279 VPB N_A_303_464#_c_1943_n 0.00493723f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_A_303_464#_c_1954_n 0.00225957f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_A_303_464#_c_1955_n 0.00800072f $X=-0.19 $Y=1.66 $X2=1.694
+ $Y2=1.662
cc_282 VPB Q 0.0544577f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.835
cc_283 N_SCE_M1034_g N_A_27_88#_c_375_n 0.00834942f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_284 N_SCE_M1034_g N_A_27_88#_c_376_n 0.0131974f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_285 N_SCE_c_290_n N_A_27_88#_c_376_n 0.0103131f $X=0.96 $Y=1.67 $X2=0 $Y2=0
cc_286 N_SCE_c_292_n N_A_27_88#_c_376_n 0.0273678f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_287 N_SCE_M1005_g N_A_27_88#_c_384_n 0.0140661f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_288 N_SCE_M1002_g N_A_27_88#_c_384_n 8.96015e-19 $X=1.005 $Y=2.64 $X2=0 $Y2=0
cc_289 N_SCE_M1034_g N_A_27_88#_c_377_n 0.0204376f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_290 N_SCE_c_290_n N_A_27_88#_c_377_n 0.00325047f $X=0.96 $Y=1.67 $X2=0 $Y2=0
cc_291 N_SCE_c_292_n N_A_27_88#_c_377_n 0.0382971f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_292 N_SCE_c_287_n N_A_27_88#_c_385_n 0.0233402f $X=2.345 $Y=1.575 $X2=0 $Y2=0
cc_293 N_SCE_c_288_n N_A_27_88#_c_386_n 0.0291709f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_294 N_SCE_c_289_n N_A_27_88#_c_386_n 3.60884e-19 $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_295 N_SCE_c_287_n N_A_27_88#_c_387_n 0.00644926f $X=2.345 $Y=1.575 $X2=0
+ $Y2=0
cc_296 N_SCE_c_288_n N_A_27_88#_c_387_n 0.00214235f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_297 N_SCE_c_289_n N_A_27_88#_c_387_n 0.0179723f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_298 N_SCE_M1005_g N_A_27_88#_c_388_n 0.00543545f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_299 N_SCE_M1034_g N_A_27_88#_c_379_n 7.61834e-19 $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_300 N_SCE_c_292_n N_A_27_88#_c_379_n 0.0212113f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_301 N_SCE_M1034_g N_A_27_88#_c_380_n 0.00727818f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_302 N_SCE_c_290_n N_A_27_88#_c_380_n 0.00441678f $X=0.96 $Y=1.67 $X2=0 $Y2=0
cc_303 N_SCE_c_292_n N_A_27_88#_c_380_n 0.008287f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_304 N_SCE_M1005_g N_A_27_88#_c_389_n 0.013502f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_305 N_SCE_M1002_g N_A_27_88#_c_389_n 0.0168794f $X=1.005 $Y=2.64 $X2=0 $Y2=0
cc_306 N_SCE_c_287_n N_A_27_88#_c_389_n 0.0109158f $X=2.345 $Y=1.575 $X2=0 $Y2=0
cc_307 N_SCE_c_290_n N_A_27_88#_c_389_n 0.00381149f $X=0.96 $Y=1.67 $X2=0 $Y2=0
cc_308 N_SCE_c_292_n N_A_27_88#_c_389_n 0.101415f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_309 N_SCE_M1002_g N_D_c_456_n 0.0062192f $X=1.005 $Y=2.64 $X2=0 $Y2=0
cc_310 N_SCE_c_292_n N_D_c_456_n 0.00447951f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_311 N_SCE_c_298_n N_D_c_456_n 0.00929488f $X=1.795 $Y=1.662 $X2=0 $Y2=0
cc_312 N_SCE_c_288_n N_D_c_457_n 0.00129438f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_313 N_SCE_c_289_n N_D_c_457_n 0.00957253f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_314 N_SCE_M1002_g N_D_c_464_n 0.0539454f $X=1.005 $Y=2.64 $X2=0 $Y2=0
cc_315 N_SCE_c_292_n N_D_c_464_n 0.00172785f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_316 N_SCE_c_287_n N_D_c_458_n 0.00657898f $X=2.345 $Y=1.575 $X2=0 $Y2=0
cc_317 N_SCE_c_290_n N_D_c_458_n 0.00663484f $X=0.96 $Y=1.67 $X2=0 $Y2=0
cc_318 N_SCE_c_292_n N_D_c_458_n 0.00195725f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_319 N_SCE_c_298_n N_D_c_458_n 0.0037388f $X=1.795 $Y=1.662 $X2=0 $Y2=0
cc_320 N_SCE_c_286_n N_D_c_459_n 0.00800462f $X=2.625 $Y=1.05 $X2=0 $Y2=0
cc_321 N_SCE_c_287_n N_D_c_459_n 0.00281358f $X=2.345 $Y=1.575 $X2=0 $Y2=0
cc_322 N_SCE_c_289_n N_D_c_459_n 3.01001e-19 $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_323 N_SCE_c_285_n N_D_c_460_n 2.00624e-19 $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_324 N_SCE_c_286_n N_D_c_460_n 2.26947e-19 $X=2.625 $Y=1.05 $X2=0 $Y2=0
cc_325 N_SCE_c_291_n N_D_c_460_n 9.5263e-19 $X=2.51 $Y=1.26 $X2=0 $Y2=0
cc_326 N_SCE_c_292_n N_D_c_460_n 0.0338107f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_327 N_SCE_c_285_n N_D_c_461_n 0.00692407f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_328 N_SCE_c_286_n N_D_c_461_n 5.10539e-19 $X=2.625 $Y=1.05 $X2=0 $Y2=0
cc_329 N_SCE_c_285_n N_SCD_M1015_g 0.0408623f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_330 N_SCE_c_288_n N_SCD_M1015_g 0.00402266f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_331 N_SCE_c_291_n N_SCD_M1015_g 0.0171335f $X=2.51 $Y=1.26 $X2=0 $Y2=0
cc_332 N_SCE_c_288_n SCD 0.0144929f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_333 N_SCE_c_288_n N_SCD_c_515_n 0.002632f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_334 N_SCE_c_289_n N_SCD_c_515_n 0.00936322f $X=2.51 $Y=1.425 $X2=0 $Y2=0
cc_335 N_SCE_M1005_g N_VPWR_c_1777_n 0.00334717f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_336 N_SCE_M1002_g N_VPWR_c_1777_n 0.016273f $X=1.005 $Y=2.64 $X2=0 $Y2=0
cc_337 N_SCE_M1005_g N_VPWR_c_1792_n 0.005209f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_338 N_SCE_M1002_g N_VPWR_c_1793_n 0.00460063f $X=1.005 $Y=2.64 $X2=0 $Y2=0
cc_339 N_SCE_M1005_g N_VPWR_c_1776_n 0.00985824f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_340 N_SCE_M1002_g N_VPWR_c_1776_n 0.00908371f $X=1.005 $Y=2.64 $X2=0 $Y2=0
cc_341 N_SCE_M1002_g N_A_303_464#_c_1946_n 0.00178733f $X=1.005 $Y=2.64 $X2=0
+ $Y2=0
cc_342 N_SCE_c_286_n N_A_303_464#_c_1937_n 0.00703396f $X=2.625 $Y=1.05 $X2=0
+ $Y2=0
cc_343 N_SCE_c_288_n N_A_303_464#_c_1937_n 0.00943064f $X=2.51 $Y=1.425 $X2=0
+ $Y2=0
cc_344 N_SCE_c_291_n N_A_303_464#_c_1937_n 0.00186472f $X=2.51 $Y=1.26 $X2=0
+ $Y2=0
cc_345 N_SCE_c_285_n N_A_303_464#_c_1944_n 0.00663897f $X=2.625 $Y=0.9 $X2=0
+ $Y2=0
cc_346 N_SCE_c_286_n N_A_303_464#_c_1944_n 0.00472894f $X=2.625 $Y=1.05 $X2=0
+ $Y2=0
cc_347 N_SCE_c_287_n N_A_303_464#_c_1944_n 0.00336351f $X=2.345 $Y=1.575 $X2=0
+ $Y2=0
cc_348 N_SCE_c_288_n N_A_303_464#_c_1944_n 0.0208536f $X=2.51 $Y=1.425 $X2=0
+ $Y2=0
cc_349 N_SCE_c_289_n N_A_303_464#_c_1944_n 0.0013723f $X=2.51 $Y=1.425 $X2=0
+ $Y2=0
cc_350 N_SCE_c_291_n N_A_303_464#_c_1944_n 0.00193022f $X=2.51 $Y=1.26 $X2=0
+ $Y2=0
cc_351 N_SCE_M1034_g N_VGND_c_2120_n 0.0142996f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_352 N_SCE_M1034_g N_VGND_c_2128_n 0.00438299f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_353 N_SCE_c_285_n N_VGND_c_2129_n 9.15902e-19 $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_354 N_SCE_M1034_g N_VGND_c_2135_n 0.00439883f $X=0.495 $Y=0.65 $X2=0 $Y2=0
cc_355 N_SCE_c_285_n N_noxref_24_c_2252_n 0.0120947f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_356 N_SCE_M1034_g N_noxref_24_c_2253_n 8.90151e-19 $X=0.495 $Y=0.65 $X2=0
+ $Y2=0
cc_357 N_SCE_c_285_n N_noxref_24_c_2254_n 0.001431f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_358 N_A_27_88#_c_385_n N_D_c_456_n 0.00102504f $X=2.207 $Y=2.002 $X2=0 $Y2=0
cc_359 N_A_27_88#_c_387_n N_D_c_456_n 0.0190261f $X=2.51 $Y=1.995 $X2=0 $Y2=0
cc_360 N_A_27_88#_c_389_n N_D_c_456_n 0.00492692f $X=2.035 $Y=2.002 $X2=0 $Y2=0
cc_361 N_A_27_88#_c_389_n N_D_c_464_n 0.0192419f $X=2.035 $Y=2.002 $X2=0 $Y2=0
cc_362 N_A_27_88#_c_389_n N_D_c_458_n 7.9327e-19 $X=2.035 $Y=2.002 $X2=0 $Y2=0
cc_363 N_A_27_88#_c_387_n N_D_c_459_n 0.00133757f $X=2.51 $Y=1.995 $X2=0 $Y2=0
cc_364 N_A_27_88#_c_379_n N_D_c_459_n 2.69613e-19 $X=1.21 $Y=1.1 $X2=0 $Y2=0
cc_365 N_A_27_88#_c_380_n N_D_c_459_n 0.0143534f $X=1.21 $Y=1.1 $X2=0 $Y2=0
cc_366 N_A_27_88#_c_374_n N_D_c_460_n 0.00484268f $X=1.485 $Y=0.935 $X2=0 $Y2=0
cc_367 N_A_27_88#_c_379_n N_D_c_460_n 0.0250153f $X=1.21 $Y=1.1 $X2=0 $Y2=0
cc_368 N_A_27_88#_c_380_n N_D_c_460_n 0.0014755f $X=1.21 $Y=1.1 $X2=0 $Y2=0
cc_369 N_A_27_88#_c_374_n N_D_c_461_n 0.0356736f $X=1.485 $Y=0.935 $X2=0 $Y2=0
cc_370 N_A_27_88#_c_381_n N_SCD_c_513_n 0.0133038f $X=2.585 $Y=2.16 $X2=0 $Y2=0
cc_371 N_A_27_88#_c_386_n N_SCD_c_513_n 0.00290511f $X=2.51 $Y=1.995 $X2=0 $Y2=0
cc_372 N_A_27_88#_M1016_g N_SCD_c_517_n 0.0532358f $X=2.585 $Y=2.64 $X2=0 $Y2=0
cc_373 N_A_27_88#_c_381_n SCD 3.43581e-19 $X=2.585 $Y=2.16 $X2=0 $Y2=0
cc_374 N_A_27_88#_c_386_n SCD 0.0207487f $X=2.51 $Y=1.995 $X2=0 $Y2=0
cc_375 N_A_27_88#_c_384_n N_VPWR_c_1777_n 0.0246172f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_376 N_A_27_88#_c_389_n N_VPWR_c_1777_n 0.0227172f $X=2.035 $Y=2.002 $X2=0
+ $Y2=0
cc_377 N_A_27_88#_M1016_g N_VPWR_c_1778_n 0.00139042f $X=2.585 $Y=2.64 $X2=0
+ $Y2=0
cc_378 N_A_27_88#_c_384_n N_VPWR_c_1792_n 0.014549f $X=0.28 $Y=2.465 $X2=0 $Y2=0
cc_379 N_A_27_88#_M1016_g N_VPWR_c_1793_n 0.00485831f $X=2.585 $Y=2.64 $X2=0
+ $Y2=0
cc_380 N_A_27_88#_M1016_g N_VPWR_c_1776_n 0.00514146f $X=2.585 $Y=2.64 $X2=0
+ $Y2=0
cc_381 N_A_27_88#_c_384_n N_VPWR_c_1776_n 0.0119743f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_382 N_A_27_88#_c_387_n N_A_303_464#_c_1946_n 0.00354002f $X=2.51 $Y=1.995
+ $X2=0 $Y2=0
cc_383 N_A_27_88#_c_389_n N_A_303_464#_c_1946_n 0.0309465f $X=2.035 $Y=2.002
+ $X2=0 $Y2=0
cc_384 N_A_27_88#_M1016_g N_A_303_464#_c_1968_n 0.00809766f $X=2.585 $Y=2.64
+ $X2=0 $Y2=0
cc_385 N_A_27_88#_c_386_n N_A_303_464#_c_1968_n 0.0309465f $X=2.51 $Y=1.995
+ $X2=0 $Y2=0
cc_386 N_A_27_88#_M1016_g N_A_303_464#_c_1954_n 0.0128106f $X=2.585 $Y=2.64
+ $X2=0 $Y2=0
cc_387 N_A_27_88#_c_385_n N_A_303_464#_c_1954_n 0.0309465f $X=2.207 $Y=2.002
+ $X2=0 $Y2=0
cc_388 N_A_27_88#_c_374_n N_VGND_c_2120_n 0.00578639f $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_389 N_A_27_88#_c_375_n N_VGND_c_2120_n 0.0179429f $X=0.28 $Y=0.65 $X2=0 $Y2=0
cc_390 N_A_27_88#_c_377_n N_VGND_c_2120_n 0.0279517f $X=1.045 $Y=1.157 $X2=0
+ $Y2=0
cc_391 N_A_27_88#_c_375_n N_VGND_c_2128_n 0.00862619f $X=0.28 $Y=0.65 $X2=0
+ $Y2=0
cc_392 N_A_27_88#_c_374_n N_VGND_c_2129_n 9.09582e-19 $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_393 N_A_27_88#_c_375_n N_VGND_c_2135_n 0.00876292f $X=0.28 $Y=0.65 $X2=0
+ $Y2=0
cc_394 N_A_27_88#_c_374_n N_noxref_24_c_2252_n 0.0108727f $X=1.485 $Y=0.935
+ $X2=0 $Y2=0
cc_395 N_A_27_88#_c_374_n N_noxref_24_c_2253_n 0.00859442f $X=1.485 $Y=0.935
+ $X2=0 $Y2=0
cc_396 N_A_27_88#_c_379_n N_noxref_24_c_2253_n 0.0133426f $X=1.21 $Y=1.1 $X2=0
+ $Y2=0
cc_397 N_A_27_88#_c_380_n N_noxref_24_c_2253_n 0.0017694f $X=1.21 $Y=1.1 $X2=0
+ $Y2=0
cc_398 N_D_c_462_n N_VPWR_c_1777_n 0.00234685f $X=1.425 $Y=2.225 $X2=0 $Y2=0
cc_399 N_D_c_462_n N_VPWR_c_1793_n 0.00519794f $X=1.425 $Y=2.225 $X2=0 $Y2=0
cc_400 N_D_c_462_n N_VPWR_c_1776_n 0.00984666f $X=1.425 $Y=2.225 $X2=0 $Y2=0
cc_401 N_D_c_460_n N_A_303_464#_M1009_d 0.00160189f $X=1.935 $Y=1.1 $X2=-0.19
+ $Y2=-0.245
cc_402 N_D_c_462_n N_A_303_464#_c_1946_n 0.012911f $X=1.425 $Y=2.225 $X2=0 $Y2=0
cc_403 N_D_c_464_n N_A_303_464#_c_1946_n 0.00624489f $X=1.69 $Y=2.15 $X2=0 $Y2=0
cc_404 N_D_c_459_n N_A_303_464#_c_1944_n 6.08332e-19 $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_405 N_D_c_460_n N_A_303_464#_c_1944_n 0.0234915f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_406 N_D_c_461_n N_A_303_464#_c_1944_n 0.00517774f $X=1.935 $Y=0.935 $X2=0
+ $Y2=0
cc_407 N_D_c_461_n N_VGND_c_2129_n 9.15902e-19 $X=1.935 $Y=0.935 $X2=0 $Y2=0
cc_408 N_D_c_459_n N_noxref_24_c_2252_n 5.66605e-19 $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_409 N_D_c_460_n N_noxref_24_c_2252_n 0.0128576f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_410 N_D_c_461_n N_noxref_24_c_2252_n 0.011902f $X=1.935 $Y=0.935 $X2=0 $Y2=0
cc_411 N_D_c_461_n N_noxref_24_c_2253_n 0.00113655f $X=1.935 $Y=0.935 $X2=0
+ $Y2=0
cc_412 N_D_c_460_n noxref_25 0.00198619f $X=1.935 $Y=1.1 $X2=-0.19 $Y2=-0.245
cc_413 N_SCD_M1015_g N_RESET_B_M1036_g 0.0329664f $X=3.04 $Y=0.615 $X2=0 $Y2=0
cc_414 SCD N_RESET_B_M1036_g 0.00424522f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_415 N_SCD_c_515_n N_RESET_B_M1036_g 0.0255034f $X=3.05 $Y=1.605 $X2=0 $Y2=0
cc_416 N_SCD_c_513_n N_RESET_B_c_933_n 0.0255034f $X=3.05 $Y=2.08 $X2=0 $Y2=0
cc_417 N_SCD_c_517_n N_RESET_B_c_938_n 0.0183737f $X=3.05 $Y=2.245 $X2=0 $Y2=0
cc_418 N_SCD_c_517_n N_VPWR_c_1778_n 0.0102726f $X=3.05 $Y=2.245 $X2=0 $Y2=0
cc_419 N_SCD_c_517_n N_VPWR_c_1793_n 0.00460063f $X=3.05 $Y=2.245 $X2=0 $Y2=0
cc_420 N_SCD_c_517_n N_VPWR_c_1776_n 0.00454691f $X=3.05 $Y=2.245 $X2=0 $Y2=0
cc_421 N_SCD_c_517_n N_A_303_464#_c_1968_n 0.0177692f $X=3.05 $Y=2.245 $X2=0
+ $Y2=0
cc_422 SCD N_A_303_464#_c_1968_n 0.0212141f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_423 N_SCD_M1015_g N_A_303_464#_c_1937_n 0.0123829f $X=3.04 $Y=0.615 $X2=0
+ $Y2=0
cc_424 SCD N_A_303_464#_c_1937_n 0.0149629f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_425 N_SCD_c_515_n N_A_303_464#_c_1937_n 0.00280161f $X=3.05 $Y=1.605 $X2=0
+ $Y2=0
cc_426 N_SCD_M1015_g N_A_303_464#_c_1938_n 0.00207067f $X=3.04 $Y=0.615 $X2=0
+ $Y2=0
cc_427 N_SCD_c_517_n N_A_303_464#_c_1938_n 0.00218868f $X=3.05 $Y=2.245 $X2=0
+ $Y2=0
cc_428 SCD N_A_303_464#_c_1938_n 0.0535746f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_429 N_SCD_c_515_n N_A_303_464#_c_1938_n 7.6448e-19 $X=3.05 $Y=1.605 $X2=0
+ $Y2=0
cc_430 N_SCD_c_517_n N_A_303_464#_c_1949_n 7.47337e-19 $X=3.05 $Y=2.245 $X2=0
+ $Y2=0
cc_431 N_SCD_c_517_n N_A_303_464#_c_1954_n 0.00174599f $X=3.05 $Y=2.245 $X2=0
+ $Y2=0
cc_432 N_SCD_M1015_g N_A_303_464#_c_1944_n 0.00135432f $X=3.04 $Y=0.615 $X2=0
+ $Y2=0
cc_433 N_SCD_M1015_g N_VGND_c_2129_n 9.09315e-19 $X=3.04 $Y=0.615 $X2=0 $Y2=0
cc_434 N_SCD_M1015_g N_noxref_24_c_2252_n 0.00698763f $X=3.04 $Y=0.615 $X2=0
+ $Y2=0
cc_435 N_SCD_M1015_g N_noxref_24_c_2254_n 0.01038f $X=3.04 $Y=0.615 $X2=0 $Y2=0
cc_436 N_CLK_c_553_n N_A_1037_387#_c_613_n 9.62665e-19 $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_437 N_CLK_c_556_n N_A_1037_387#_c_631_n 5.28783e-19 $X=4.645 $Y=1.86 $X2=0
+ $Y2=0
cc_438 N_CLK_c_553_n N_RESET_B_M1036_g 0.0213809f $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_439 CLK N_RESET_B_M1036_g 0.00322884f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_440 N_CLK_c_553_n N_RESET_B_c_922_n 0.0100723f $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_441 CLK N_RESET_B_c_922_n 0.00667701f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_442 N_CLK_c_553_n N_RESET_B_c_932_n 0.0229612f $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_443 N_CLK_c_556_n N_RESET_B_c_932_n 0.00444062f $X=4.645 $Y=1.86 $X2=0 $Y2=0
cc_444 CLK N_RESET_B_c_932_n 0.00124257f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_445 N_CLK_c_553_n N_RESET_B_c_939_n 6.34206e-19 $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_446 CLK N_RESET_B_c_939_n 0.00698533f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_447 N_CLK_c_556_n N_RESET_B_c_940_n 3.98306e-19 $X=4.645 $Y=1.86 $X2=0 $Y2=0
cc_448 CLK N_RESET_B_c_940_n 0.00449516f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_449 N_CLK_c_553_n N_RESET_B_c_945_n 0.00111606f $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_450 N_CLK_c_556_n N_RESET_B_c_945_n 7.01353e-19 $X=4.645 $Y=1.86 $X2=0 $Y2=0
cc_451 CLK N_RESET_B_c_945_n 0.0310766f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_452 CLK N_A_835_93#_M1029_s 0.00709744f $X=3.995 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_453 N_CLK_c_553_n N_A_835_93#_c_1287_n 0.0474507f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_454 N_CLK_c_553_n N_A_835_93#_c_1275_n 0.0210768f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_455 N_CLK_c_553_n N_A_835_93#_c_1277_n 0.0265768f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_456 CLK N_A_835_93#_c_1277_n 3.01982e-19 $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_457 N_CLK_c_553_n N_A_835_93#_c_1305_n 0.00608321f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_458 N_CLK_c_553_n N_A_835_93#_c_1306_n 0.0102663f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_459 CLK N_A_835_93#_c_1306_n 0.00778119f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_460 N_CLK_c_553_n N_A_835_93#_c_1308_n 0.00409385f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_461 CLK N_A_835_93#_c_1308_n 0.0241878f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_462 N_CLK_c_556_n N_A_835_93#_c_1310_n 0.0129999f $X=4.645 $Y=1.86 $X2=0
+ $Y2=0
cc_463 CLK N_A_835_93#_c_1310_n 0.00366247f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_464 N_CLK_c_553_n N_A_835_93#_c_1284_n 0.00345877f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_465 CLK N_A_835_93#_c_1284_n 0.0202553f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_466 N_CLK_c_553_n N_A_835_93#_c_1298_n 0.00216991f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_467 N_CLK_c_553_n N_A_835_93#_c_1285_n 0.00882412f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_468 CLK N_A_835_93#_c_1285_n 0.0112621f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_469 N_CLK_c_553_n N_A_835_93#_c_1317_n 0.00578473f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_470 N_CLK_c_556_n N_A_835_93#_c_1317_n 0.00382572f $X=4.645 $Y=1.86 $X2=0
+ $Y2=0
cc_471 CLK N_A_835_93#_c_1317_n 0.0154577f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_472 N_CLK_c_553_n N_A_835_93#_c_1286_n 0.00320572f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_473 CLK N_A_835_93#_c_1286_n 0.0279373f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_474 N_CLK_c_556_n N_VPWR_c_1779_n 0.0182372f $X=4.645 $Y=1.86 $X2=0 $Y2=0
cc_475 N_CLK_c_556_n N_VPWR_c_1786_n 0.00425118f $X=4.645 $Y=1.86 $X2=0 $Y2=0
cc_476 N_CLK_c_556_n N_VPWR_c_1776_n 0.00633028f $X=4.645 $Y=1.86 $X2=0 $Y2=0
cc_477 CLK N_A_303_464#_c_1937_n 0.0153429f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_478 N_CLK_c_553_n N_A_303_464#_c_1938_n 0.00320931f $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_479 CLK N_A_303_464#_c_1938_n 0.0460205f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_480 N_CLK_c_553_n N_A_303_464#_c_1948_n 3.15997e-19 $X=4.595 $Y=1.41 $X2=0
+ $Y2=0
cc_481 N_CLK_c_556_n N_A_303_464#_c_1948_n 0.0162077f $X=4.645 $Y=1.86 $X2=0
+ $Y2=0
cc_482 N_CLK_c_556_n N_A_303_464#_c_1949_n 0.00181048f $X=4.645 $Y=1.86 $X2=0
+ $Y2=0
cc_483 N_CLK_c_556_n N_A_303_464#_c_1955_n 0.00880061f $X=4.645 $Y=1.86 $X2=0
+ $Y2=0
cc_484 N_CLK_c_553_n N_VGND_c_2121_n 0.00199669f $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_485 CLK N_VGND_c_2121_n 0.00867496f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_486 N_CLK_c_553_n N_VGND_c_2122_n 0.0028517f $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_487 N_CLK_c_553_n N_VGND_c_2135_n 9.39239e-19 $X=4.595 $Y=1.41 $X2=0 $Y2=0
cc_488 N_A_1037_387#_c_620_n N_A_1367_93#_M1033_d 0.00176461f $X=9.065 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_489 N_A_1037_387#_M1001_g N_A_1367_93#_M1020_g 0.0333343f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_490 N_A_1037_387#_c_615_n N_A_1367_93#_M1020_g 0.00311064f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_491 N_A_1037_387#_c_618_n N_A_1367_93#_M1020_g 0.00262964f $X=7.135 $Y=0.58
+ $X2=0 $Y2=0
cc_492 N_A_1037_387#_c_643_p N_A_1367_93#_M1020_g 0.0026982f $X=7.22 $Y=0.665
+ $X2=0 $Y2=0
cc_493 N_A_1037_387#_c_609_n N_A_1367_93#_c_819_n 0.0333343f $X=6.45 $Y=1.65
+ $X2=0 $Y2=0
cc_494 N_A_1037_387#_c_627_n N_A_1367_93#_c_819_n 0.00102464f $X=6.065 $Y=1.65
+ $X2=0 $Y2=0
cc_495 N_A_1037_387#_c_619_n N_A_1367_93#_c_820_n 0.0520186f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_496 N_A_1037_387#_c_620_n N_A_1367_93#_c_820_n 0.00353238f $X=9.065 $Y=0.34
+ $X2=0 $Y2=0
cc_497 N_A_1037_387#_c_619_n N_A_1367_93#_c_821_n 0.00761753f $X=7.93 $Y=0.665
+ $X2=0 $Y2=0
cc_498 N_A_1037_387#_c_643_p N_A_1367_93#_c_821_n 0.0103944f $X=7.22 $Y=0.665
+ $X2=0 $Y2=0
cc_499 N_A_1037_387#_c_623_n N_A_1367_93#_c_827_n 0.00471763f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_500 N_A_1037_387#_c_628_n N_A_1367_93#_c_827_n 0.00323506f $X=9.085 $Y=1.105
+ $X2=0 $Y2=0
cc_501 N_A_1037_387#_c_611_n N_A_1367_93#_c_822_n 0.014712f $X=8.65 $Y=1.085
+ $X2=0 $Y2=0
cc_502 N_A_1037_387#_c_612_n N_A_1367_93#_c_822_n 0.00243289f $X=8.725 $Y=1.16
+ $X2=0 $Y2=0
cc_503 N_A_1037_387#_c_620_n N_A_1367_93#_c_822_n 0.0257761f $X=9.065 $Y=0.34
+ $X2=0 $Y2=0
cc_504 N_A_1037_387#_c_622_n N_A_1367_93#_c_822_n 0.0141828f $X=9.15 $Y=0.94
+ $X2=0 $Y2=0
cc_505 N_A_1037_387#_c_625_n N_A_1367_93#_c_822_n 5.79172e-19 $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_506 N_A_1037_387#_c_626_n N_A_1367_93#_c_822_n 0.0131302f $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_507 N_A_1037_387#_c_628_n N_A_1367_93#_c_822_n 0.00313966f $X=9.085 $Y=1.105
+ $X2=0 $Y2=0
cc_508 N_A_1037_387#_c_623_n N_A_1367_93#_c_823_n 0.0197158f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_509 N_A_1037_387#_c_625_n N_A_1367_93#_c_823_n 2.26254e-19 $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_510 N_A_1037_387#_c_626_n N_A_1367_93#_c_823_n 0.0131446f $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_511 N_A_1037_387#_c_628_n N_A_1367_93#_c_823_n 0.00960948f $X=9.085 $Y=1.105
+ $X2=0 $Y2=0
cc_512 N_A_1037_387#_M1001_g N_RESET_B_c_922_n 0.00882199f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_513 N_A_1037_387#_c_615_n N_RESET_B_c_922_n 0.0294278f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_514 N_A_1037_387#_c_616_n N_RESET_B_c_922_n 0.00992957f $X=5.62 $Y=0.34 $X2=0
+ $Y2=0
cc_515 N_A_1037_387#_c_615_n N_RESET_B_M1012_g 0.00466687f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_516 N_A_1037_387#_c_618_n N_RESET_B_M1012_g 0.00445709f $X=7.135 $Y=0.58
+ $X2=0 $Y2=0
cc_517 N_A_1037_387#_c_619_n N_RESET_B_M1012_g 0.0128143f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_518 N_A_1037_387#_c_669_p N_RESET_B_M1012_g 0.0035287f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_519 N_A_1037_387#_c_621_n N_RESET_B_M1012_g 6.46496e-19 $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_520 N_A_1037_387#_M1030_d N_RESET_B_c_939_n 0.00342297f $X=5.185 $Y=1.935
+ $X2=0 $Y2=0
cc_521 N_A_1037_387#_M1000_g N_RESET_B_c_939_n 0.00340123f $X=6.135 $Y=2.495
+ $X2=0 $Y2=0
cc_522 N_A_1037_387#_c_609_n N_RESET_B_c_939_n 0.00388808f $X=6.45 $Y=1.65 $X2=0
+ $Y2=0
cc_523 N_A_1037_387#_c_631_n N_RESET_B_c_939_n 0.0301466f $X=5.63 $Y=1.71 $X2=0
+ $Y2=0
cc_524 N_A_1037_387#_c_617_n N_RESET_B_c_939_n 0.0163625f $X=6.065 $Y=1.71 $X2=0
+ $Y2=0
cc_525 N_A_1037_387#_c_627_n N_RESET_B_c_939_n 0.00379596f $X=6.065 $Y=1.65
+ $X2=0 $Y2=0
cc_526 N_A_1037_387#_c_623_n N_RESET_B_c_941_n 0.0173785f $X=9.33 $Y=2.125 $X2=0
+ $Y2=0
cc_527 N_A_1037_387#_c_634_n N_RESET_B_c_941_n 0.0197423f $X=9.81 $Y=2.215 $X2=0
+ $Y2=0
cc_528 N_A_1037_387#_c_636_n N_RESET_B_c_941_n 0.00644248f $X=9.89 $Y=2.215
+ $X2=0 $Y2=0
cc_529 N_A_1037_387#_c_611_n N_A_1234_119#_M1033_g 0.0286306f $X=8.65 $Y=1.085
+ $X2=0 $Y2=0
cc_530 N_A_1037_387#_c_620_n N_A_1234_119#_M1033_g 0.0116373f $X=9.065 $Y=0.34
+ $X2=0 $Y2=0
cc_531 N_A_1037_387#_c_612_n N_A_1234_119#_c_1147_n 0.0153032f $X=8.725 $Y=1.16
+ $X2=0 $Y2=0
cc_532 N_A_1037_387#_c_623_n N_A_1234_119#_c_1147_n 4.45025e-19 $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_533 N_A_1037_387#_c_609_n N_A_1234_119#_c_1157_n 7.69506e-19 $X=6.45 $Y=1.65
+ $X2=0 $Y2=0
cc_534 N_A_1037_387#_M1001_g N_A_1234_119#_c_1148_n 0.0102762f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_535 N_A_1037_387#_c_615_n N_A_1234_119#_c_1148_n 0.0118472f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_536 N_A_1037_387#_M1000_g N_A_1234_119#_c_1149_n 9.59875e-19 $X=6.135
+ $Y=2.495 $X2=0 $Y2=0
cc_537 N_A_1037_387#_M1001_g N_A_1234_119#_c_1149_n 0.0068601f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_538 N_A_1037_387#_c_609_n N_A_1234_119#_c_1154_n 4.79797e-19 $X=6.45 $Y=1.65
+ $X2=0 $Y2=0
cc_539 N_A_1037_387#_M1001_g N_A_1234_119#_c_1154_n 0.00636651f $X=6.525
+ $Y=0.805 $X2=0 $Y2=0
cc_540 N_A_1037_387#_c_615_n N_A_1234_119#_c_1154_n 0.019863f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_541 N_A_1037_387#_c_643_p N_A_1234_119#_c_1154_n 0.00486547f $X=7.22 $Y=0.665
+ $X2=0 $Y2=0
cc_542 N_A_1037_387#_c_631_n N_A_835_93#_c_1287_n 0.00556337f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_543 N_A_1037_387#_c_613_n N_A_835_93#_c_1275_n 0.010288f $X=5.36 $Y=0.74
+ $X2=0 $Y2=0
cc_544 N_A_1037_387#_c_614_n N_A_835_93#_c_1275_n 0.00105741f $X=5.54 $Y=1.545
+ $X2=0 $Y2=0
cc_545 N_A_1037_387#_c_624_n N_A_835_93#_c_1275_n 0.00138092f $X=5.422 $Y=1.265
+ $X2=0 $Y2=0
cc_546 N_A_1037_387#_M1000_g N_A_835_93#_c_1288_n 0.024942f $X=6.135 $Y=2.495
+ $X2=0 $Y2=0
cc_547 N_A_1037_387#_c_631_n N_A_835_93#_c_1288_n 0.0145816f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_548 N_A_1037_387#_c_617_n N_A_835_93#_c_1288_n 0.00175916f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_549 N_A_1037_387#_M1000_g N_A_835_93#_c_1289_n 0.0107339f $X=6.135 $Y=2.495
+ $X2=0 $Y2=0
cc_550 N_A_1037_387#_c_617_n N_A_835_93#_c_1276_n 0.00417616f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_551 N_A_1037_387#_c_627_n N_A_835_93#_c_1276_n 0.0173325f $X=6.065 $Y=1.65
+ $X2=0 $Y2=0
cc_552 N_A_1037_387#_c_614_n N_A_835_93#_c_1277_n 0.0146301f $X=5.54 $Y=1.545
+ $X2=0 $Y2=0
cc_553 N_A_1037_387#_c_631_n N_A_835_93#_c_1277_n 0.0169559f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_554 N_A_1037_387#_c_617_n N_A_835_93#_c_1277_n 0.00794502f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_555 N_A_1037_387#_c_624_n N_A_835_93#_c_1277_n 0.0109985f $X=5.422 $Y=1.265
+ $X2=0 $Y2=0
cc_556 N_A_1037_387#_c_627_n N_A_835_93#_c_1277_n 0.0215064f $X=6.065 $Y=1.65
+ $X2=0 $Y2=0
cc_557 N_A_1037_387#_M1001_g N_A_835_93#_M1035_g 0.022001f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_558 N_A_1037_387#_c_613_n N_A_835_93#_M1035_g 0.00479917f $X=5.36 $Y=0.74
+ $X2=0 $Y2=0
cc_559 N_A_1037_387#_c_615_n N_A_835_93#_M1035_g 0.00330666f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_560 N_A_1037_387#_M1000_g N_A_835_93#_M1017_g 0.0117434f $X=6.135 $Y=2.495
+ $X2=0 $Y2=0
cc_561 N_A_1037_387#_c_609_n N_A_835_93#_M1017_g 0.0015696f $X=6.45 $Y=1.65
+ $X2=0 $Y2=0
cc_562 N_A_1037_387#_M1014_g N_A_835_93#_M1031_g 0.0149474f $X=9.89 $Y=2.75
+ $X2=0 $Y2=0
cc_563 N_A_1037_387#_c_623_n N_A_835_93#_M1031_g 0.00903517f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_564 N_A_1037_387#_c_636_n N_A_835_93#_M1031_g 0.00826222f $X=9.89 $Y=2.215
+ $X2=0 $Y2=0
cc_565 N_A_1037_387#_c_623_n N_A_835_93#_c_1279_n 0.0121351f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_566 N_A_1037_387#_c_634_n N_A_835_93#_c_1279_n 0.00479207f $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_567 N_A_1037_387#_c_636_n N_A_835_93#_c_1279_n 0.00418242f $X=9.89 $Y=2.215
+ $X2=0 $Y2=0
cc_568 N_A_1037_387#_c_625_n N_A_835_93#_c_1280_n 0.0191612f $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_569 N_A_1037_387#_c_626_n N_A_835_93#_c_1280_n 0.00166135f $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_570 N_A_1037_387#_c_628_n N_A_835_93#_c_1280_n 0.00150758f $X=9.085 $Y=1.105
+ $X2=0 $Y2=0
cc_571 N_A_1037_387#_c_623_n N_A_835_93#_c_1281_n 0.00153175f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_572 N_A_1037_387#_c_620_n N_A_835_93#_M1004_g 0.00301232f $X=9.065 $Y=0.34
+ $X2=0 $Y2=0
cc_573 N_A_1037_387#_c_622_n N_A_835_93#_M1004_g 0.00129859f $X=9.15 $Y=0.94
+ $X2=0 $Y2=0
cc_574 N_A_1037_387#_c_625_n N_A_835_93#_M1004_g 0.00125371f $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_575 N_A_1037_387#_c_625_n N_A_835_93#_c_1283_n 0.0194128f $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_576 N_A_1037_387#_c_626_n N_A_835_93#_c_1283_n 3.65519e-19 $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_577 N_A_1037_387#_c_631_n N_A_835_93#_c_1310_n 0.00962532f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_578 N_A_1037_387#_c_614_n N_A_835_93#_c_1284_n 0.00570182f $X=5.54 $Y=1.545
+ $X2=0 $Y2=0
cc_579 N_A_1037_387#_c_631_n N_A_835_93#_c_1298_n 0.00517731f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_580 N_A_1037_387#_c_631_n N_A_835_93#_c_1317_n 0.0032297f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_581 N_A_1037_387#_c_614_n N_A_835_93#_c_1286_n 0.00730886f $X=5.54 $Y=1.545
+ $X2=0 $Y2=0
cc_582 N_A_1037_387#_c_631_n N_A_835_93#_c_1286_n 0.0281469f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_583 N_A_1037_387#_c_624_n N_A_835_93#_c_1286_n 0.00257969f $X=5.422 $Y=1.265
+ $X2=0 $Y2=0
cc_584 N_A_1037_387#_c_634_n N_A_1997_272#_M1037_g 2.75671e-19 $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_585 N_A_1037_387#_c_636_n N_A_1997_272#_M1037_g 0.0560328f $X=9.89 $Y=2.215
+ $X2=0 $Y2=0
cc_586 N_A_1037_387#_c_620_n N_A_1745_74#_M1006_d 0.00630965f $X=9.065 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_587 N_A_1037_387#_c_622_n N_A_1745_74#_M1006_d 0.0113887f $X=9.15 $Y=0.94
+ $X2=-0.19 $Y2=-0.245
cc_588 N_A_1037_387#_c_623_n N_A_1745_74#_M1031_d 0.0072549f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_589 N_A_1037_387#_c_740_p N_A_1745_74#_M1031_d 0.00308947f $X=9.415 $Y=2.252
+ $X2=0 $Y2=0
cc_590 N_A_1037_387#_c_634_n N_A_1745_74#_M1031_d 0.00176657f $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_591 N_A_1037_387#_M1014_g N_A_1745_74#_c_1590_n 0.0199621f $X=9.89 $Y=2.75
+ $X2=0 $Y2=0
cc_592 N_A_1037_387#_c_740_p N_A_1745_74#_c_1590_n 0.01001f $X=9.415 $Y=2.252
+ $X2=0 $Y2=0
cc_593 N_A_1037_387#_c_634_n N_A_1745_74#_c_1590_n 0.0389958f $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_594 N_A_1037_387#_c_636_n N_A_1745_74#_c_1590_n 0.00338558f $X=9.89 $Y=2.215
+ $X2=0 $Y2=0
cc_595 N_A_1037_387#_c_622_n N_A_1745_74#_c_1579_n 0.00768735f $X=9.15 $Y=0.94
+ $X2=0 $Y2=0
cc_596 N_A_1037_387#_c_625_n N_A_1745_74#_c_1579_n 4.55554e-19 $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_597 N_A_1037_387#_c_626_n N_A_1745_74#_c_1579_n 0.0116456f $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_598 N_A_1037_387#_c_623_n N_A_1745_74#_c_1580_n 0.0375442f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_599 N_A_1037_387#_c_634_n N_A_1745_74#_c_1592_n 0.0125258f $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_600 N_A_1037_387#_c_636_n N_A_1745_74#_c_1592_n 0.00446735f $X=9.89 $Y=2.215
+ $X2=0 $Y2=0
cc_601 N_A_1037_387#_c_623_n N_A_1745_74#_c_1593_n 0.0141313f $X=9.33 $Y=2.125
+ $X2=0 $Y2=0
cc_602 N_A_1037_387#_c_634_n N_A_1745_74#_c_1593_n 0.0111216f $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_603 N_A_1037_387#_c_636_n N_A_1745_74#_c_1593_n 9.16255e-19 $X=9.89 $Y=2.215
+ $X2=0 $Y2=0
cc_604 N_A_1037_387#_c_634_n N_A_1745_74#_c_1594_n 0.0202186f $X=9.81 $Y=2.215
+ $X2=0 $Y2=0
cc_605 N_A_1037_387#_c_636_n N_A_1745_74#_c_1594_n 0.00627357f $X=9.89 $Y=2.215
+ $X2=0 $Y2=0
cc_606 N_A_1037_387#_c_611_n N_A_1745_74#_c_1581_n 5.77109e-19 $X=8.65 $Y=1.085
+ $X2=0 $Y2=0
cc_607 N_A_1037_387#_c_620_n N_A_1745_74#_c_1581_n 0.00648023f $X=9.065 $Y=0.34
+ $X2=0 $Y2=0
cc_608 N_A_1037_387#_c_622_n N_A_1745_74#_c_1581_n 0.0264512f $X=9.15 $Y=0.94
+ $X2=0 $Y2=0
cc_609 N_A_1037_387#_c_625_n N_A_1745_74#_c_1581_n 2.06488e-19 $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_610 N_A_1037_387#_c_626_n N_A_1745_74#_c_1581_n 7.15367e-19 $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_611 N_A_1037_387#_c_625_n N_A_1745_74#_c_1582_n 6.39686e-19 $X=9.25 $Y=1.105
+ $X2=0 $Y2=0
cc_612 N_A_1037_387#_c_626_n N_A_1745_74#_c_1582_n 0.0144646f $X=9.33 $Y=1.105
+ $X2=0 $Y2=0
cc_613 N_A_1037_387#_M1014_g N_VPWR_c_1788_n 0.00365611f $X=9.89 $Y=2.75 $X2=0
+ $Y2=0
cc_614 N_A_1037_387#_M1000_g N_VPWR_c_1776_n 0.00113998f $X=6.135 $Y=2.495 $X2=0
+ $Y2=0
cc_615 N_A_1037_387#_M1014_g N_VPWR_c_1776_n 0.00449015f $X=9.89 $Y=2.75 $X2=0
+ $Y2=0
cc_616 N_A_1037_387#_M1030_d N_A_303_464#_c_1948_n 0.00628547f $X=5.185 $Y=1.935
+ $X2=0 $Y2=0
cc_617 N_A_1037_387#_c_631_n N_A_303_464#_c_1948_n 0.0307389f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_618 N_A_1037_387#_c_617_n N_A_303_464#_c_1948_n 0.00248787f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_619 N_A_1037_387#_c_613_n N_A_303_464#_c_1939_n 0.0342763f $X=5.36 $Y=0.74
+ $X2=0 $Y2=0
cc_620 N_A_1037_387#_c_615_n N_A_303_464#_c_1939_n 0.013349f $X=7.05 $Y=0.34
+ $X2=0 $Y2=0
cc_621 N_A_1037_387#_c_613_n N_A_303_464#_c_1940_n 0.00574014f $X=5.36 $Y=0.74
+ $X2=0 $Y2=0
cc_622 N_A_1037_387#_c_624_n N_A_303_464#_c_1940_n 0.00712827f $X=5.422 $Y=1.265
+ $X2=0 $Y2=0
cc_623 N_A_1037_387#_M1000_g N_A_303_464#_c_1950_n 0.00897858f $X=6.135 $Y=2.495
+ $X2=0 $Y2=0
cc_624 N_A_1037_387#_c_631_n N_A_303_464#_c_1950_n 0.00500857f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_625 N_A_1037_387#_c_609_n N_A_303_464#_c_1941_n 0.00319576f $X=6.45 $Y=1.65
+ $X2=0 $Y2=0
cc_626 N_A_1037_387#_M1001_g N_A_303_464#_c_1941_n 0.00615688f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_627 N_A_1037_387#_c_617_n N_A_303_464#_c_1941_n 0.0160606f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_628 N_A_1037_387#_c_627_n N_A_303_464#_c_1941_n 0.00280396f $X=6.065 $Y=1.65
+ $X2=0 $Y2=0
cc_629 N_A_1037_387#_c_617_n N_A_303_464#_c_1942_n 0.0144255f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_630 N_A_1037_387#_c_624_n N_A_303_464#_c_1942_n 0.0134292f $X=5.422 $Y=1.265
+ $X2=0 $Y2=0
cc_631 N_A_1037_387#_c_627_n N_A_303_464#_c_1942_n 4.61571e-19 $X=6.065 $Y=1.65
+ $X2=0 $Y2=0
cc_632 N_A_1037_387#_M1000_g N_A_303_464#_c_1951_n 0.0131959f $X=6.135 $Y=2.495
+ $X2=0 $Y2=0
cc_633 N_A_1037_387#_c_609_n N_A_303_464#_c_1951_n 0.00254238f $X=6.45 $Y=1.65
+ $X2=0 $Y2=0
cc_634 N_A_1037_387#_c_617_n N_A_303_464#_c_1951_n 0.00770757f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_635 N_A_1037_387#_M1000_g N_A_303_464#_c_1952_n 0.00250682f $X=6.135 $Y=2.495
+ $X2=0 $Y2=0
cc_636 N_A_1037_387#_c_631_n N_A_303_464#_c_1952_n 0.0123094f $X=5.63 $Y=1.71
+ $X2=0 $Y2=0
cc_637 N_A_1037_387#_c_617_n N_A_303_464#_c_1952_n 0.0168093f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_638 N_A_1037_387#_c_627_n N_A_303_464#_c_1952_n 0.00323248f $X=6.065 $Y=1.65
+ $X2=0 $Y2=0
cc_639 N_A_1037_387#_M1000_g N_A_303_464#_c_1943_n 0.00549102f $X=6.135 $Y=2.495
+ $X2=0 $Y2=0
cc_640 N_A_1037_387#_c_609_n N_A_303_464#_c_1943_n 0.0106696f $X=6.45 $Y=1.65
+ $X2=0 $Y2=0
cc_641 N_A_1037_387#_M1001_g N_A_303_464#_c_1943_n 0.00578983f $X=6.525 $Y=0.805
+ $X2=0 $Y2=0
cc_642 N_A_1037_387#_c_617_n N_A_303_464#_c_1943_n 0.0256508f $X=6.065 $Y=1.71
+ $X2=0 $Y2=0
cc_643 N_A_1037_387#_c_627_n N_A_303_464#_c_1943_n 0.00266104f $X=6.065 $Y=1.65
+ $X2=0 $Y2=0
cc_644 N_A_1037_387#_c_619_n N_VGND_M1012_d 0.0170064f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_645 N_A_1037_387#_c_669_p N_VGND_M1012_d 0.00275919f $X=8.015 $Y=0.58 $X2=0
+ $Y2=0
cc_646 N_A_1037_387#_c_621_n N_VGND_M1012_d 7.93589e-19 $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_647 N_A_1037_387#_c_613_n N_VGND_c_2122_n 0.0189029f $X=5.36 $Y=0.74 $X2=0
+ $Y2=0
cc_648 N_A_1037_387#_c_616_n N_VGND_c_2122_n 0.0144411f $X=5.62 $Y=0.34 $X2=0
+ $Y2=0
cc_649 N_A_1037_387#_c_615_n N_VGND_c_2130_n 0.103356f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_650 N_A_1037_387#_c_616_n N_VGND_c_2130_n 0.0276098f $X=5.62 $Y=0.34 $X2=0
+ $Y2=0
cc_651 N_A_1037_387#_c_619_n N_VGND_c_2130_n 0.00402072f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_652 N_A_1037_387#_c_611_n N_VGND_c_2131_n 0.00278271f $X=8.65 $Y=1.085 $X2=0
+ $Y2=0
cc_653 N_A_1037_387#_c_619_n N_VGND_c_2131_n 0.00335833f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_654 N_A_1037_387#_c_620_n N_VGND_c_2131_n 0.0734255f $X=9.065 $Y=0.34 $X2=0
+ $Y2=0
cc_655 N_A_1037_387#_c_621_n N_VGND_c_2131_n 0.0118998f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_656 N_A_1037_387#_c_611_n N_VGND_c_2135_n 0.00358525f $X=8.65 $Y=1.085 $X2=0
+ $Y2=0
cc_657 N_A_1037_387#_c_615_n N_VGND_c_2135_n 0.0538367f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_658 N_A_1037_387#_c_616_n N_VGND_c_2135_n 0.0138923f $X=5.62 $Y=0.34 $X2=0
+ $Y2=0
cc_659 N_A_1037_387#_c_619_n N_VGND_c_2135_n 0.0122484f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_660 N_A_1037_387#_c_620_n N_VGND_c_2135_n 0.0415191f $X=9.065 $Y=0.34 $X2=0
+ $Y2=0
cc_661 N_A_1037_387#_c_621_n N_VGND_c_2135_n 0.00655543f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_662 N_A_1037_387#_c_615_n N_VGND_c_2138_n 0.0118008f $X=7.05 $Y=0.34 $X2=0
+ $Y2=0
cc_663 N_A_1037_387#_c_619_n N_VGND_c_2138_n 0.0246013f $X=7.93 $Y=0.665 $X2=0
+ $Y2=0
cc_664 N_A_1037_387#_c_621_n N_VGND_c_2138_n 0.0135793f $X=8.1 $Y=0.34 $X2=0
+ $Y2=0
cc_665 N_A_1037_387#_c_643_p A_1397_119# 0.00349303f $X=7.22 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_666 N_A_1367_93#_M1020_g N_RESET_B_c_922_n 0.00882199f $X=6.91 $Y=0.805 $X2=0
+ $Y2=0
cc_667 N_A_1367_93#_c_821_n N_RESET_B_c_922_n 2.57602e-19 $X=7.325 $Y=1.005
+ $X2=0 $Y2=0
cc_668 N_A_1367_93#_M1020_g N_RESET_B_M1012_g 0.0398707f $X=6.91 $Y=0.805 $X2=0
+ $Y2=0
cc_669 N_A_1367_93#_c_818_n N_RESET_B_M1012_g 0.00127951f $X=7.185 $Y=1.64 $X2=0
+ $Y2=0
cc_670 N_A_1367_93#_c_820_n N_RESET_B_M1012_g 0.00681742f $X=8.27 $Y=1.005 $X2=0
+ $Y2=0
cc_671 N_A_1367_93#_c_821_n N_RESET_B_M1012_g 0.00424625f $X=7.325 $Y=1.005
+ $X2=0 $Y2=0
cc_672 N_A_1367_93#_c_820_n N_RESET_B_c_925_n 0.0117401f $X=8.27 $Y=1.005 $X2=0
+ $Y2=0
cc_673 N_A_1367_93#_c_818_n N_RESET_B_c_926_n 0.00932005f $X=7.185 $Y=1.64 $X2=0
+ $Y2=0
cc_674 N_A_1367_93#_c_819_n N_RESET_B_c_926_n 0.0083853f $X=7.185 $Y=1.64 $X2=0
+ $Y2=0
cc_675 N_A_1367_93#_M1020_g N_RESET_B_c_927_n 0.0024449f $X=6.91 $Y=0.805 $X2=0
+ $Y2=0
cc_676 N_A_1367_93#_M1028_g N_RESET_B_c_927_n 0.0244836f $X=7.06 $Y=2.515 $X2=0
+ $Y2=0
cc_677 N_A_1367_93#_c_818_n N_RESET_B_c_927_n 0.00103605f $X=7.185 $Y=1.64 $X2=0
+ $Y2=0
cc_678 N_A_1367_93#_c_819_n N_RESET_B_c_927_n 0.0173421f $X=7.185 $Y=1.64 $X2=0
+ $Y2=0
cc_679 N_A_1367_93#_M1028_g N_RESET_B_c_939_n 0.0101599f $X=7.06 $Y=2.515 $X2=0
+ $Y2=0
cc_680 N_A_1367_93#_c_818_n N_RESET_B_c_939_n 0.00823427f $X=7.185 $Y=1.64 $X2=0
+ $Y2=0
cc_681 N_A_1367_93#_c_819_n N_RESET_B_c_939_n 0.00318126f $X=7.185 $Y=1.64 $X2=0
+ $Y2=0
cc_682 N_A_1367_93#_M1026_d N_RESET_B_c_941_n 0.00365135f $X=8.785 $Y=1.735
+ $X2=0 $Y2=0
cc_683 N_A_1367_93#_c_828_n N_RESET_B_c_941_n 0.0364688f $X=8.92 $Y=1.88 $X2=0
+ $Y2=0
cc_684 N_A_1367_93#_c_820_n N_A_1234_119#_M1033_g 0.01076f $X=8.27 $Y=1.005
+ $X2=0 $Y2=0
cc_685 N_A_1367_93#_c_822_n N_A_1234_119#_M1033_g 0.0114957f $X=8.435 $Y=0.81
+ $X2=0 $Y2=0
cc_686 N_A_1367_93#_c_823_n N_A_1234_119#_M1033_g 9.26224e-19 $X=8.865 $Y=1.715
+ $X2=0 $Y2=0
cc_687 N_A_1367_93#_c_822_n N_A_1234_119#_c_1147_n 0.00717853f $X=8.435 $Y=0.81
+ $X2=0 $Y2=0
cc_688 N_A_1367_93#_c_823_n N_A_1234_119#_c_1147_n 0.00666709f $X=8.865 $Y=1.715
+ $X2=0 $Y2=0
cc_689 N_A_1367_93#_c_827_n N_A_1234_119#_M1026_g 0.00304901f $X=8.865 $Y=1.855
+ $X2=0 $Y2=0
cc_690 N_A_1367_93#_c_828_n N_A_1234_119#_M1026_g 0.0127532f $X=8.92 $Y=1.88
+ $X2=0 $Y2=0
cc_691 N_A_1367_93#_c_823_n N_A_1234_119#_M1026_g 0.00586625f $X=8.865 $Y=1.715
+ $X2=0 $Y2=0
cc_692 N_A_1367_93#_M1020_g N_A_1234_119#_c_1148_n 0.004969f $X=6.91 $Y=0.805
+ $X2=0 $Y2=0
cc_693 N_A_1367_93#_c_821_n N_A_1234_119#_c_1148_n 0.00929856f $X=7.325 $Y=1.005
+ $X2=0 $Y2=0
cc_694 N_A_1367_93#_M1020_g N_A_1234_119#_c_1149_n 0.00772383f $X=6.91 $Y=0.805
+ $X2=0 $Y2=0
cc_695 N_A_1367_93#_M1028_g N_A_1234_119#_c_1149_n 0.0109301f $X=7.06 $Y=2.515
+ $X2=0 $Y2=0
cc_696 N_A_1367_93#_c_818_n N_A_1234_119#_c_1149_n 0.0517809f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_697 N_A_1367_93#_c_819_n N_A_1234_119#_c_1149_n 0.00938542f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_698 N_A_1367_93#_c_821_n N_A_1234_119#_c_1149_n 0.00480628f $X=7.325 $Y=1.005
+ $X2=0 $Y2=0
cc_699 N_A_1367_93#_M1028_g N_A_1234_119#_c_1190_n 0.012749f $X=7.06 $Y=2.515
+ $X2=0 $Y2=0
cc_700 N_A_1367_93#_c_818_n N_A_1234_119#_c_1190_n 0.00338945f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_701 N_A_1367_93#_c_819_n N_A_1234_119#_c_1190_n 0.00333925f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_702 N_A_1367_93#_M1028_g N_A_1234_119#_c_1150_n 0.00485223f $X=7.06 $Y=2.515
+ $X2=0 $Y2=0
cc_703 N_A_1367_93#_c_818_n N_A_1234_119#_c_1150_n 0.0170101f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_704 N_A_1367_93#_c_819_n N_A_1234_119#_c_1150_n 0.00147646f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_705 N_A_1367_93#_c_818_n N_A_1234_119#_c_1151_n 0.0270592f $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_706 N_A_1367_93#_c_819_n N_A_1234_119#_c_1151_n 7.33487e-19 $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_707 N_A_1367_93#_c_820_n N_A_1234_119#_c_1151_n 0.0135416f $X=8.27 $Y=1.005
+ $X2=0 $Y2=0
cc_708 N_A_1367_93#_c_820_n N_A_1234_119#_c_1152_n 0.0457531f $X=8.27 $Y=1.005
+ $X2=0 $Y2=0
cc_709 N_A_1367_93#_c_822_n N_A_1234_119#_c_1152_n 0.00357705f $X=8.435 $Y=0.81
+ $X2=0 $Y2=0
cc_710 N_A_1367_93#_c_823_n N_A_1234_119#_c_1152_n 0.0123924f $X=8.865 $Y=1.715
+ $X2=0 $Y2=0
cc_711 N_A_1367_93#_c_820_n N_A_1234_119#_c_1153_n 0.00365093f $X=8.27 $Y=1.005
+ $X2=0 $Y2=0
cc_712 N_A_1367_93#_c_822_n N_A_1234_119#_c_1153_n 4.74815e-19 $X=8.435 $Y=0.81
+ $X2=0 $Y2=0
cc_713 N_A_1367_93#_c_823_n N_A_1234_119#_c_1153_n 0.00153128f $X=8.865 $Y=1.715
+ $X2=0 $Y2=0
cc_714 N_A_1367_93#_M1020_g N_A_1234_119#_c_1154_n 0.00107029f $X=6.91 $Y=0.805
+ $X2=0 $Y2=0
cc_715 N_A_1367_93#_M1028_g N_A_1234_119#_c_1161_n 0.00559455f $X=7.06 $Y=2.515
+ $X2=0 $Y2=0
cc_716 N_A_1367_93#_M1028_g N_A_835_93#_M1017_g 0.0354987f $X=7.06 $Y=2.515
+ $X2=0 $Y2=0
cc_717 N_A_1367_93#_M1028_g N_A_835_93#_c_1293_n 0.0114392f $X=7.06 $Y=2.515
+ $X2=0 $Y2=0
cc_718 N_A_1367_93#_c_828_n N_A_835_93#_c_1293_n 0.00382437f $X=8.92 $Y=1.88
+ $X2=0 $Y2=0
cc_719 N_A_1367_93#_c_827_n N_A_835_93#_M1031_g 5.91667e-19 $X=8.865 $Y=1.855
+ $X2=0 $Y2=0
cc_720 N_A_1367_93#_c_823_n N_A_835_93#_c_1280_n 0.00176495f $X=8.865 $Y=1.715
+ $X2=0 $Y2=0
cc_721 N_A_1367_93#_c_822_n N_A_1745_74#_M1006_d 0.00295216f $X=8.435 $Y=0.81
+ $X2=-0.19 $Y2=-0.245
cc_722 N_A_1367_93#_c_828_n N_A_1745_74#_c_1590_n 0.00115576f $X=8.92 $Y=1.88
+ $X2=0 $Y2=0
cc_723 N_A_1367_93#_M1028_g N_VPWR_c_1780_n 0.00423282f $X=7.06 $Y=2.515 $X2=0
+ $Y2=0
cc_724 N_A_1367_93#_c_827_n N_VPWR_c_1782_n 0.0395418f $X=8.865 $Y=1.855 $X2=0
+ $Y2=0
cc_725 N_A_1367_93#_c_822_n N_VPWR_c_1782_n 0.0054981f $X=8.435 $Y=0.81 $X2=0
+ $Y2=0
cc_726 N_A_1367_93#_c_828_n N_VPWR_c_1788_n 0.00626239f $X=8.92 $Y=1.88 $X2=0
+ $Y2=0
cc_727 N_A_1367_93#_M1028_g N_VPWR_c_1776_n 0.0011317f $X=7.06 $Y=2.515 $X2=0
+ $Y2=0
cc_728 N_A_1367_93#_c_828_n N_VPWR_c_1776_n 0.00764493f $X=8.92 $Y=1.88 $X2=0
+ $Y2=0
cc_729 N_A_1367_93#_M1020_g N_A_303_464#_c_1943_n 3.24142e-19 $X=6.91 $Y=0.805
+ $X2=0 $Y2=0
cc_730 N_A_1367_93#_c_819_n N_A_303_464#_c_1943_n 2.3169e-19 $X=7.185 $Y=1.64
+ $X2=0 $Y2=0
cc_731 N_A_1367_93#_c_820_n N_VGND_M1012_d 0.00911951f $X=8.27 $Y=1.005 $X2=0
+ $Y2=0
cc_732 N_A_1367_93#_c_821_n A_1397_119# 0.00204263f $X=7.325 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_733 N_RESET_B_c_925_n N_A_1234_119#_M1033_g 0.0052575f $X=7.595 $Y=1.19 $X2=0
+ $Y2=0
cc_734 N_RESET_B_c_941_n N_A_1234_119#_M1026_g 0.00941657f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_735 N_RESET_B_c_939_n N_A_1234_119#_c_1157_n 0.00855554f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_736 N_RESET_B_M1012_g N_A_1234_119#_c_1148_n 3.96747e-19 $X=7.3 $Y=0.805
+ $X2=0 $Y2=0
cc_737 N_RESET_B_c_939_n N_A_1234_119#_c_1149_n 0.023753f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_738 N_RESET_B_c_939_n N_A_1234_119#_c_1190_n 0.0214903f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_739 N_RESET_B_c_927_n N_A_1234_119#_c_1150_n 0.0113497f $X=7.67 $Y=1.815
+ $X2=0 $Y2=0
cc_740 N_RESET_B_M1010_g N_A_1234_119#_c_1150_n 0.0240975f $X=7.685 $Y=2.515
+ $X2=0 $Y2=0
cc_741 N_RESET_B_c_939_n N_A_1234_119#_c_1150_n 0.0272492f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_742 N_RESET_B_c_942_n N_A_1234_119#_c_1150_n 0.0119438f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_743 N_RESET_B_c_943_n N_A_1234_119#_c_1150_n 0.0388968f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_744 N_RESET_B_c_946_n N_A_1234_119#_c_1150_n 0.0115469f $X=8 $Y=1.98 $X2=0
+ $Y2=0
cc_745 N_RESET_B_c_925_n N_A_1234_119#_c_1151_n 0.00404376f $X=7.595 $Y=1.19
+ $X2=0 $Y2=0
cc_746 N_RESET_B_c_927_n N_A_1234_119#_c_1151_n 0.00501753f $X=7.67 $Y=1.815
+ $X2=0 $Y2=0
cc_747 N_RESET_B_c_925_n N_A_1234_119#_c_1152_n 7.39613e-19 $X=7.595 $Y=1.19
+ $X2=0 $Y2=0
cc_748 N_RESET_B_c_927_n N_A_1234_119#_c_1152_n 0.00710493f $X=7.67 $Y=1.815
+ $X2=0 $Y2=0
cc_749 N_RESET_B_c_939_n N_A_1234_119#_c_1152_n 0.00357593f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_750 N_RESET_B_c_941_n N_A_1234_119#_c_1152_n 0.00581394f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_751 N_RESET_B_c_942_n N_A_1234_119#_c_1152_n 0.00371961f $X=8.065 $Y=2.035
+ $X2=0 $Y2=0
cc_752 N_RESET_B_c_943_n N_A_1234_119#_c_1152_n 0.0172409f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_753 N_RESET_B_c_946_n N_A_1234_119#_c_1152_n 0.00739726f $X=8 $Y=1.98 $X2=0
+ $Y2=0
cc_754 N_RESET_B_c_925_n N_A_1234_119#_c_1153_n 0.0182615f $X=7.595 $Y=1.19
+ $X2=0 $Y2=0
cc_755 N_RESET_B_c_927_n N_A_1234_119#_c_1153_n 6.54113e-19 $X=7.67 $Y=1.815
+ $X2=0 $Y2=0
cc_756 N_RESET_B_c_941_n N_A_1234_119#_c_1153_n 0.00590391f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_757 N_RESET_B_c_943_n N_A_1234_119#_c_1153_n 6.74459e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_758 N_RESET_B_c_946_n N_A_1234_119#_c_1153_n 0.0093828f $X=8 $Y=1.98 $X2=0
+ $Y2=0
cc_759 N_RESET_B_c_939_n N_A_835_93#_M1018_s 0.00115526f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_760 N_RESET_B_c_939_n N_A_835_93#_c_1287_n 0.00406718f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_761 N_RESET_B_c_922_n N_A_835_93#_c_1275_n 0.0103973f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_762 N_RESET_B_c_939_n N_A_835_93#_c_1288_n 0.00223435f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_763 N_RESET_B_c_939_n N_A_835_93#_c_1277_n 0.00534227f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_764 N_RESET_B_c_922_n N_A_835_93#_M1035_g 0.00882199f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_765 N_RESET_B_c_939_n N_A_835_93#_M1017_g 0.00413599f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_766 N_RESET_B_M1010_g N_A_835_93#_c_1293_n 0.0113685f $X=7.685 $Y=2.515 $X2=0
+ $Y2=0
cc_767 N_RESET_B_c_941_n N_A_835_93#_M1031_g 0.0161088f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_768 N_RESET_B_c_941_n N_A_835_93#_c_1279_n 0.00354541f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_769 N_RESET_B_c_922_n N_A_835_93#_c_1306_n 0.00127515f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_770 N_RESET_B_c_939_n N_A_835_93#_c_1310_n 0.0225778f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_771 N_RESET_B_c_940_n N_A_835_93#_c_1298_n 6.58602e-19 $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_772 N_RESET_B_c_945_n N_A_835_93#_c_1298_n 0.00327062f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_773 N_RESET_B_c_922_n N_A_835_93#_c_1285_n 0.00782328f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_774 N_RESET_B_c_932_n N_A_835_93#_c_1317_n 6.13411e-19 $X=3.93 $Y=1.995 $X2=0
+ $Y2=0
cc_775 N_RESET_B_c_933_n N_A_835_93#_c_1317_n 0.00153911f $X=3.695 $Y=1.995
+ $X2=0 $Y2=0
cc_776 N_RESET_B_c_939_n N_A_835_93#_c_1317_n 0.01139f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_777 N_RESET_B_c_940_n N_A_835_93#_c_1317_n 0.00185043f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_778 N_RESET_B_c_945_n N_A_835_93#_c_1317_n 0.0195373f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_779 N_RESET_B_c_939_n N_A_835_93#_c_1286_n 0.0088587f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_780 N_RESET_B_M1038_g N_A_1997_272#_M1003_g 0.0312551f $X=10.6 $Y=0.58 $X2=0
+ $Y2=0
cc_781 N_RESET_B_c_929_n N_A_1997_272#_c_1465_n 0.0225363f $X=10.715 $Y=1.82
+ $X2=0 $Y2=0
cc_782 N_RESET_B_c_930_n N_A_1997_272#_c_1465_n 0.00643996f $X=10.715 $Y=1.375
+ $X2=0 $Y2=0
cc_783 N_RESET_B_c_947_n N_A_1997_272#_c_1465_n 0.00119422f $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_784 N_RESET_B_M1021_g N_A_1997_272#_M1037_g 0.0202099f $X=10.885 $Y=2.75
+ $X2=0 $Y2=0
cc_785 N_RESET_B_c_941_n N_A_1997_272#_M1037_g 0.00514751f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_786 N_RESET_B_c_948_n N_A_1997_272#_M1037_g 0.0128577f $X=10.885 $Y=1.985
+ $X2=0 $Y2=0
cc_787 N_RESET_B_c_929_n N_A_1997_272#_c_1466_n 0.00935059f $X=10.715 $Y=1.82
+ $X2=0 $Y2=0
cc_788 N_RESET_B_c_930_n N_A_1997_272#_c_1466_n 0.0053082f $X=10.715 $Y=1.375
+ $X2=0 $Y2=0
cc_789 RESET_B N_A_1997_272#_c_1466_n 0.00164136f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_790 N_RESET_B_c_947_n N_A_1997_272#_c_1466_n 0.0191591f $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_791 N_RESET_B_c_948_n N_A_1997_272#_c_1466_n 0.00143756f $X=10.885 $Y=1.985
+ $X2=0 $Y2=0
cc_792 N_RESET_B_M1038_g N_A_1997_272#_c_1467_n 0.00111706f $X=10.6 $Y=0.58
+ $X2=0 $Y2=0
cc_793 N_RESET_B_M1038_g N_A_1997_272#_c_1470_n 7.22053e-19 $X=10.6 $Y=0.58
+ $X2=0 $Y2=0
cc_794 N_RESET_B_c_941_n N_A_1997_272#_c_1472_n 0.0131744f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_795 N_RESET_B_M1021_g N_A_1997_272#_c_1477_n 0.00756168f $X=10.885 $Y=2.75
+ $X2=0 $Y2=0
cc_796 N_RESET_B_c_947_n N_A_1997_272#_c_1477_n 9.53119e-19 $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_797 N_RESET_B_c_929_n N_A_1997_272#_c_1473_n 0.00366777f $X=10.715 $Y=1.82
+ $X2=0 $Y2=0
cc_798 RESET_B N_A_1997_272#_c_1473_n 0.00158814f $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_799 N_RESET_B_c_947_n N_A_1997_272#_c_1473_n 0.0232461f $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_800 N_RESET_B_c_948_n N_A_1997_272#_c_1473_n 0.00971401f $X=10.885 $Y=1.985
+ $X2=0 $Y2=0
cc_801 N_RESET_B_c_941_n N_A_1745_74#_M1031_d 0.00215383f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_802 N_RESET_B_M1038_g N_A_1745_74#_M1022_g 0.0518692f $X=10.6 $Y=0.58 $X2=0
+ $Y2=0
cc_803 N_RESET_B_c_930_n N_A_1745_74#_c_1575_n 0.0117915f $X=10.715 $Y=1.375
+ $X2=0 $Y2=0
cc_804 N_RESET_B_c_947_n N_A_1745_74#_c_1575_n 3.43698e-19 $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_805 N_RESET_B_c_948_n N_A_1745_74#_c_1575_n 0.0195805f $X=10.885 $Y=1.985
+ $X2=0 $Y2=0
cc_806 N_RESET_B_M1038_g N_A_1745_74#_c_1577_n 0.00646231f $X=10.6 $Y=0.58 $X2=0
+ $Y2=0
cc_807 N_RESET_B_c_930_n N_A_1745_74#_c_1577_n 0.0030434f $X=10.715 $Y=1.375
+ $X2=0 $Y2=0
cc_808 N_RESET_B_M1021_g N_A_1745_74#_c_1589_n 0.0195805f $X=10.885 $Y=2.75
+ $X2=0 $Y2=0
cc_809 N_RESET_B_c_941_n N_A_1745_74#_c_1590_n 0.00559189f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_810 N_RESET_B_c_929_n N_A_1745_74#_c_1592_n 6.20198e-19 $X=10.715 $Y=1.82
+ $X2=0 $Y2=0
cc_811 N_RESET_B_c_941_n N_A_1745_74#_c_1592_n 0.0131083f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_812 RESET_B N_A_1745_74#_c_1592_n 2.51275e-19 $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_813 N_RESET_B_c_947_n N_A_1745_74#_c_1592_n 0.00608543f $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_814 N_RESET_B_c_941_n N_A_1745_74#_c_1593_n 0.0053742f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_815 N_RESET_B_M1021_g N_A_1745_74#_c_1594_n 0.00189085f $X=10.885 $Y=2.75
+ $X2=0 $Y2=0
cc_816 N_RESET_B_c_941_n N_A_1745_74#_c_1594_n 0.020931f $X=10.655 $Y=2.035
+ $X2=0 $Y2=0
cc_817 RESET_B N_A_1745_74#_c_1594_n 3.29892e-19 $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_818 N_RESET_B_c_947_n N_A_1745_74#_c_1594_n 0.00622512f $X=10.805 $Y=1.985
+ $X2=0 $Y2=0
cc_819 N_RESET_B_c_948_n N_A_1745_74#_c_1594_n 6.08738e-19 $X=10.885 $Y=1.985
+ $X2=0 $Y2=0
cc_820 N_RESET_B_M1038_g N_A_1745_74#_c_1584_n 0.015752f $X=10.6 $Y=0.58 $X2=0
+ $Y2=0
cc_821 N_RESET_B_c_930_n N_A_1745_74#_c_1584_n 0.00357206f $X=10.715 $Y=1.375
+ $X2=0 $Y2=0
cc_822 N_RESET_B_c_939_n N_VPWR_M1018_d 4.24275e-19 $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_823 N_RESET_B_c_941_n N_VPWR_M1026_s 0.00596563f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_824 N_RESET_B_c_938_n N_VPWR_c_1778_n 0.00580956f $X=3.56 $Y=2.245 $X2=0
+ $Y2=0
cc_825 N_RESET_B_M1010_g N_VPWR_c_1780_n 0.00386909f $X=7.685 $Y=2.515 $X2=0
+ $Y2=0
cc_826 N_RESET_B_c_939_n N_VPWR_c_1780_n 7.54713e-19 $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_827 N_RESET_B_c_927_n N_VPWR_c_1782_n 0.00146391f $X=7.67 $Y=1.815 $X2=0
+ $Y2=0
cc_828 N_RESET_B_M1010_g N_VPWR_c_1782_n 0.00704456f $X=7.685 $Y=2.515 $X2=0
+ $Y2=0
cc_829 N_RESET_B_c_941_n N_VPWR_c_1782_n 0.0186169f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_830 N_RESET_B_c_942_n N_VPWR_c_1782_n 5.19261e-19 $X=8.065 $Y=2.035 $X2=0
+ $Y2=0
cc_831 N_RESET_B_c_943_n N_VPWR_c_1782_n 0.0183634f $X=7.92 $Y=2.035 $X2=0 $Y2=0
cc_832 N_RESET_B_c_946_n N_VPWR_c_1782_n 0.00112124f $X=8 $Y=1.98 $X2=0 $Y2=0
cc_833 N_RESET_B_M1021_g N_VPWR_c_1783_n 0.00732775f $X=10.885 $Y=2.75 $X2=0
+ $Y2=0
cc_834 N_RESET_B_c_941_n N_VPWR_c_1783_n 0.00652534f $X=10.655 $Y=2.035 $X2=0
+ $Y2=0
cc_835 RESET_B N_VPWR_c_1783_n 6.45709e-19 $X=10.715 $Y=1.95 $X2=0 $Y2=0
cc_836 N_RESET_B_c_947_n N_VPWR_c_1783_n 0.00292772f $X=10.805 $Y=1.985 $X2=0
+ $Y2=0
cc_837 N_RESET_B_c_948_n N_VPWR_c_1783_n 6.5955e-19 $X=10.885 $Y=1.985 $X2=0
+ $Y2=0
cc_838 N_RESET_B_c_938_n N_VPWR_c_1786_n 0.005209f $X=3.56 $Y=2.245 $X2=0 $Y2=0
cc_839 N_RESET_B_M1021_g N_VPWR_c_1790_n 0.005209f $X=10.885 $Y=2.75 $X2=0 $Y2=0
cc_840 N_RESET_B_M1010_g N_VPWR_c_1776_n 0.0011317f $X=7.685 $Y=2.515 $X2=0
+ $Y2=0
cc_841 N_RESET_B_M1021_g N_VPWR_c_1776_n 0.00983777f $X=10.885 $Y=2.75 $X2=0
+ $Y2=0
cc_842 N_RESET_B_c_938_n N_VPWR_c_1776_n 0.00533602f $X=3.56 $Y=2.245 $X2=0
+ $Y2=0
cc_843 N_RESET_B_c_933_n N_A_303_464#_c_1968_n 8.77027e-19 $X=3.695 $Y=1.995
+ $X2=0 $Y2=0
cc_844 N_RESET_B_M1036_g N_A_303_464#_c_1937_n 0.0154538f $X=3.5 $Y=0.615 $X2=0
+ $Y2=0
cc_845 N_RESET_B_M1036_g N_A_303_464#_c_1938_n 0.0210607f $X=3.5 $Y=0.615 $X2=0
+ $Y2=0
cc_846 N_RESET_B_c_933_n N_A_303_464#_c_1938_n 0.0176624f $X=3.695 $Y=1.995
+ $X2=0 $Y2=0
cc_847 N_RESET_B_c_938_n N_A_303_464#_c_1938_n 0.00450975f $X=3.56 $Y=2.245
+ $X2=0 $Y2=0
cc_848 N_RESET_B_c_940_n N_A_303_464#_c_1938_n 0.00108729f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_849 N_RESET_B_c_945_n N_A_303_464#_c_1938_n 0.0258319f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_850 N_RESET_B_c_932_n N_A_303_464#_c_1948_n 6.89121e-19 $X=3.93 $Y=1.995
+ $X2=0 $Y2=0
cc_851 N_RESET_B_c_939_n N_A_303_464#_c_1948_n 0.0185926f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_852 N_RESET_B_c_940_n N_A_303_464#_c_1948_n 0.00357248f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_853 N_RESET_B_c_945_n N_A_303_464#_c_1948_n 0.00973466f $X=3.95 $Y=1.995
+ $X2=0 $Y2=0
cc_854 N_RESET_B_c_932_n N_A_303_464#_c_1949_n 0.00408396f $X=3.93 $Y=1.995
+ $X2=0 $Y2=0
cc_855 N_RESET_B_c_938_n N_A_303_464#_c_1949_n 0.0155999f $X=3.56 $Y=2.245 $X2=0
+ $Y2=0
cc_856 N_RESET_B_c_940_n N_A_303_464#_c_1949_n 4.21578e-19 $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_857 N_RESET_B_c_945_n N_A_303_464#_c_1949_n 0.0149172f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_858 N_RESET_B_c_939_n N_A_303_464#_c_1941_n 0.00360371f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_859 N_RESET_B_c_939_n N_A_303_464#_c_1951_n 0.0179072f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_860 N_RESET_B_c_939_n N_A_303_464#_c_1952_n 0.0167645f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_861 N_RESET_B_c_939_n N_A_303_464#_c_1943_n 0.0094217f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_862 N_RESET_B_c_938_n N_A_303_464#_c_1955_n 0.00564559f $X=3.56 $Y=2.245
+ $X2=0 $Y2=0
cc_863 N_RESET_B_M1036_g N_VGND_c_2121_n 0.00141396f $X=3.5 $Y=0.615 $X2=0 $Y2=0
cc_864 N_RESET_B_c_922_n N_VGND_c_2121_n 0.0211426f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_865 N_RESET_B_c_922_n N_VGND_c_2122_n 0.02563f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_866 N_RESET_B_M1038_g N_VGND_c_2123_n 0.00390833f $X=10.6 $Y=0.58 $X2=0 $Y2=0
cc_867 N_RESET_B_c_922_n N_VGND_c_2126_n 0.0242452f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_868 N_RESET_B_c_923_n N_VGND_c_2129_n 0.0064002f $X=3.575 $Y=0.18 $X2=0 $Y2=0
cc_869 N_RESET_B_c_922_n N_VGND_c_2130_n 0.0512939f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_870 N_RESET_B_M1038_g N_VGND_c_2132_n 0.00460063f $X=10.6 $Y=0.58 $X2=0 $Y2=0
cc_871 N_RESET_B_c_922_n N_VGND_c_2135_n 0.0903551f $X=7.225 $Y=0.18 $X2=0 $Y2=0
cc_872 N_RESET_B_c_923_n N_VGND_c_2135_n 0.0113744f $X=3.575 $Y=0.18 $X2=0 $Y2=0
cc_873 N_RESET_B_M1038_g N_VGND_c_2135_n 0.00906826f $X=10.6 $Y=0.58 $X2=0 $Y2=0
cc_874 N_RESET_B_c_922_n N_VGND_c_2138_n 0.00939536f $X=7.225 $Y=0.18 $X2=0
+ $Y2=0
cc_875 N_RESET_B_M1036_g N_noxref_24_c_2254_n 0.00190559f $X=3.5 $Y=0.615 $X2=0
+ $Y2=0
cc_876 N_A_1234_119#_c_1157_n N_A_835_93#_c_1289_n 0.00396944f $X=6.71 $Y=2.555
+ $X2=0 $Y2=0
cc_877 N_A_1234_119#_c_1154_n N_A_835_93#_M1035_g 0.00566398f $X=6.31 $Y=0.81
+ $X2=0 $Y2=0
cc_878 N_A_1234_119#_c_1157_n N_A_835_93#_M1017_g 0.0107269f $X=6.71 $Y=2.555
+ $X2=0 $Y2=0
cc_879 N_A_1234_119#_c_1149_n N_A_835_93#_M1017_g 0.00388381f $X=6.795 $Y=2.32
+ $X2=0 $Y2=0
cc_880 N_A_1234_119#_c_1161_n N_A_835_93#_M1017_g 0.00560099f $X=6.795 $Y=2.522
+ $X2=0 $Y2=0
cc_881 N_A_1234_119#_M1026_g N_A_835_93#_c_1293_n 0.0122143f $X=8.695 $Y=2.235
+ $X2=0 $Y2=0
cc_882 N_A_1234_119#_c_1190_n N_A_835_93#_c_1293_n 0.00281582f $X=7.495 $Y=2.405
+ $X2=0 $Y2=0
cc_883 N_A_1234_119#_c_1150_n N_A_835_93#_c_1293_n 0.00657047f $X=7.58 $Y=2.32
+ $X2=0 $Y2=0
cc_884 N_A_1234_119#_c_1161_n N_A_835_93#_c_1293_n 0.00119096f $X=6.795 $Y=2.522
+ $X2=0 $Y2=0
cc_885 N_A_1234_119#_M1026_g N_A_835_93#_M1031_g 0.00809731f $X=8.695 $Y=2.235
+ $X2=0 $Y2=0
cc_886 N_A_1234_119#_c_1147_n N_A_835_93#_c_1280_n 0.00809731f $X=8.605 $Y=1.52
+ $X2=0 $Y2=0
cc_887 N_A_1234_119#_c_1190_n N_VPWR_M1028_d 0.00719273f $X=7.495 $Y=2.405 $X2=0
+ $Y2=0
cc_888 N_A_1234_119#_c_1150_n N_VPWR_M1028_d 6.22498e-19 $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_889 N_A_1234_119#_c_1190_n N_VPWR_c_1780_n 0.0221454f $X=7.495 $Y=2.405 $X2=0
+ $Y2=0
cc_890 N_A_1234_119#_c_1150_n N_VPWR_c_1780_n 0.00708775f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_891 N_A_1234_119#_c_1150_n N_VPWR_c_1781_n 0.00710805f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_892 N_A_1234_119#_c_1147_n N_VPWR_c_1782_n 0.00454201f $X=8.605 $Y=1.52 $X2=0
+ $Y2=0
cc_893 N_A_1234_119#_M1026_g N_VPWR_c_1782_n 0.00500542f $X=8.695 $Y=2.235 $X2=0
+ $Y2=0
cc_894 N_A_1234_119#_c_1150_n N_VPWR_c_1782_n 0.0222059f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_895 N_A_1234_119#_c_1157_n N_VPWR_c_1794_n 0.00831318f $X=6.71 $Y=2.555 $X2=0
+ $Y2=0
cc_896 N_A_1234_119#_c_1161_n N_VPWR_c_1794_n 0.00289582f $X=6.795 $Y=2.522
+ $X2=0 $Y2=0
cc_897 N_A_1234_119#_M1026_g N_VPWR_c_1776_n 0.00112709f $X=8.695 $Y=2.235 $X2=0
+ $Y2=0
cc_898 N_A_1234_119#_c_1157_n N_VPWR_c_1776_n 0.0117964f $X=6.71 $Y=2.555 $X2=0
+ $Y2=0
cc_899 N_A_1234_119#_c_1190_n N_VPWR_c_1776_n 0.010332f $X=7.495 $Y=2.405 $X2=0
+ $Y2=0
cc_900 N_A_1234_119#_c_1150_n N_VPWR_c_1776_n 0.0154063f $X=7.58 $Y=2.32 $X2=0
+ $Y2=0
cc_901 N_A_1234_119#_c_1161_n N_VPWR_c_1776_n 0.00455287f $X=6.795 $Y=2.522
+ $X2=0 $Y2=0
cc_902 N_A_1234_119#_c_1157_n N_A_303_464#_c_1950_n 0.0113877f $X=6.71 $Y=2.555
+ $X2=0 $Y2=0
cc_903 N_A_1234_119#_c_1149_n N_A_303_464#_c_1950_n 0.0024271f $X=6.795 $Y=2.32
+ $X2=0 $Y2=0
cc_904 N_A_1234_119#_c_1161_n N_A_303_464#_c_1950_n 0.00169394f $X=6.795
+ $Y=2.522 $X2=0 $Y2=0
cc_905 N_A_1234_119#_c_1148_n N_A_303_464#_c_1941_n 0.00533227f $X=6.71 $Y=0.945
+ $X2=0 $Y2=0
cc_906 N_A_1234_119#_c_1149_n N_A_303_464#_c_1941_n 0.0135847f $X=6.795 $Y=2.32
+ $X2=0 $Y2=0
cc_907 N_A_1234_119#_c_1154_n N_A_303_464#_c_1941_n 0.0268176f $X=6.31 $Y=0.81
+ $X2=0 $Y2=0
cc_908 N_A_1234_119#_c_1157_n N_A_303_464#_c_1951_n 0.0196101f $X=6.71 $Y=2.555
+ $X2=0 $Y2=0
cc_909 N_A_1234_119#_c_1149_n N_A_303_464#_c_1951_n 0.0135339f $X=6.795 $Y=2.32
+ $X2=0 $Y2=0
cc_910 N_A_1234_119#_c_1149_n N_A_303_464#_c_1943_n 0.0490008f $X=6.795 $Y=2.32
+ $X2=0 $Y2=0
cc_911 N_A_1234_119#_c_1154_n N_A_303_464#_c_1945_n 0.0168155f $X=6.31 $Y=0.81
+ $X2=0 $Y2=0
cc_912 N_A_1234_119#_c_1190_n A_1346_461# 4.56836e-19 $X=7.495 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_913 N_A_1234_119#_c_1161_n A_1346_461# 0.00433362f $X=6.795 $Y=2.522
+ $X2=-0.19 $Y2=-0.245
cc_914 N_A_1234_119#_M1033_g N_VGND_c_2131_n 0.00278271f $X=8.22 $Y=0.69 $X2=0
+ $Y2=0
cc_915 N_A_1234_119#_M1033_g N_VGND_c_2135_n 0.00358525f $X=8.22 $Y=0.69 $X2=0
+ $Y2=0
cc_916 N_A_1234_119#_M1033_g N_VGND_c_2138_n 0.00111149f $X=8.22 $Y=0.69 $X2=0
+ $Y2=0
cc_917 N_A_1234_119#_c_1148_n A_1320_119# 0.00177672f $X=6.71 $Y=0.945 $X2=-0.19
+ $Y2=-0.245
cc_918 N_A_835_93#_c_1281_n N_A_1997_272#_M1003_g 0.0100846f $X=9.7 $Y=1.51
+ $X2=0 $Y2=0
cc_919 N_A_835_93#_M1004_g N_A_1997_272#_M1003_g 0.0520068f $X=9.785 $Y=0.58
+ $X2=0 $Y2=0
cc_920 N_A_835_93#_c_1281_n N_A_1997_272#_c_1465_n 0.019486f $X=9.7 $Y=1.51
+ $X2=0 $Y2=0
cc_921 N_A_835_93#_c_1281_n N_A_1997_272#_c_1472_n 6.49074e-19 $X=9.7 $Y=1.51
+ $X2=0 $Y2=0
cc_922 N_A_835_93#_M1031_g N_A_1745_74#_c_1590_n 0.0061022f $X=9.145 $Y=2.235
+ $X2=0 $Y2=0
cc_923 N_A_835_93#_M1004_g N_A_1745_74#_c_1579_n 0.00653104f $X=9.785 $Y=0.58
+ $X2=0 $Y2=0
cc_924 N_A_835_93#_c_1283_n N_A_1745_74#_c_1579_n 0.00549286f $X=9.785 $Y=1.045
+ $X2=0 $Y2=0
cc_925 N_A_835_93#_c_1279_n N_A_1745_74#_c_1580_n 0.0090777f $X=9.625 $Y=1.585
+ $X2=0 $Y2=0
cc_926 N_A_835_93#_c_1281_n N_A_1745_74#_c_1580_n 0.00911046f $X=9.7 $Y=1.51
+ $X2=0 $Y2=0
cc_927 N_A_835_93#_c_1279_n N_A_1745_74#_c_1592_n 2.60059e-19 $X=9.625 $Y=1.585
+ $X2=0 $Y2=0
cc_928 N_A_835_93#_c_1283_n N_A_1745_74#_c_1592_n 3.58986e-19 $X=9.785 $Y=1.045
+ $X2=0 $Y2=0
cc_929 N_A_835_93#_M1004_g N_A_1745_74#_c_1581_n 0.00822927f $X=9.785 $Y=0.58
+ $X2=0 $Y2=0
cc_930 N_A_835_93#_c_1281_n N_A_1745_74#_c_1582_n 0.00212136f $X=9.7 $Y=1.51
+ $X2=0 $Y2=0
cc_931 N_A_835_93#_c_1283_n N_A_1745_74#_c_1582_n 3.68292e-19 $X=9.785 $Y=1.045
+ $X2=0 $Y2=0
cc_932 N_A_835_93#_c_1281_n N_A_1745_74#_c_1584_n 0.00241471f $X=9.7 $Y=1.51
+ $X2=0 $Y2=0
cc_933 N_A_835_93#_c_1283_n N_A_1745_74#_c_1584_n 0.00651625f $X=9.785 $Y=1.045
+ $X2=0 $Y2=0
cc_934 N_A_835_93#_c_1310_n N_VPWR_M1018_d 0.0030475f $X=4.81 $Y=2.06 $X2=0
+ $Y2=0
cc_935 N_A_835_93#_c_1287_n N_VPWR_c_1779_n 0.0114622f $X=5.095 $Y=1.85 $X2=0
+ $Y2=0
cc_936 N_A_835_93#_c_1288_n N_VPWR_c_1779_n 0.00219791f $X=5.615 $Y=3.075 $X2=0
+ $Y2=0
cc_937 N_A_835_93#_M1017_g N_VPWR_c_1780_n 0.00626049f $X=6.64 $Y=2.515 $X2=0
+ $Y2=0
cc_938 N_A_835_93#_c_1293_n N_VPWR_c_1780_n 0.025635f $X=9.055 $Y=3.15 $X2=0
+ $Y2=0
cc_939 N_A_835_93#_c_1293_n N_VPWR_c_1781_n 0.0260958f $X=9.055 $Y=3.15 $X2=0
+ $Y2=0
cc_940 N_A_835_93#_c_1293_n N_VPWR_c_1782_n 0.0170937f $X=9.055 $Y=3.15 $X2=0
+ $Y2=0
cc_941 N_A_835_93#_M1031_g N_VPWR_c_1782_n 0.00538421f $X=9.145 $Y=2.235 $X2=0
+ $Y2=0
cc_942 N_A_835_93#_c_1293_n N_VPWR_c_1788_n 0.0218279f $X=9.055 $Y=3.15 $X2=0
+ $Y2=0
cc_943 N_A_835_93#_c_1287_n N_VPWR_c_1794_n 0.00425118f $X=5.095 $Y=1.85 $X2=0
+ $Y2=0
cc_944 N_A_835_93#_c_1290_n N_VPWR_c_1794_n 0.048387f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_945 N_A_835_93#_c_1287_n N_VPWR_c_1776_n 0.00520454f $X=5.095 $Y=1.85 $X2=0
+ $Y2=0
cc_946 N_A_835_93#_c_1289_n N_VPWR_c_1776_n 0.0247907f $X=6.55 $Y=3.15 $X2=0
+ $Y2=0
cc_947 N_A_835_93#_c_1290_n N_VPWR_c_1776_n 0.00561538f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_948 N_A_835_93#_c_1293_n N_VPWR_c_1776_n 0.0747517f $X=9.055 $Y=3.15 $X2=0
+ $Y2=0
cc_949 N_A_835_93#_c_1297_n N_VPWR_c_1776_n 0.00508716f $X=6.64 $Y=3.15 $X2=0
+ $Y2=0
cc_950 N_A_835_93#_M1018_s N_A_303_464#_c_1948_n 0.00754337f $X=4.275 $Y=1.935
+ $X2=0 $Y2=0
cc_951 N_A_835_93#_c_1287_n N_A_303_464#_c_1948_n 0.0158853f $X=5.095 $Y=1.85
+ $X2=0 $Y2=0
cc_952 N_A_835_93#_c_1288_n N_A_303_464#_c_1948_n 0.0138072f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_953 N_A_835_93#_c_1289_n N_A_303_464#_c_1948_n 7.51694e-19 $X=6.55 $Y=3.15
+ $X2=0 $Y2=0
cc_954 N_A_835_93#_c_1310_n N_A_303_464#_c_1948_n 0.0130343f $X=4.81 $Y=2.06
+ $X2=0 $Y2=0
cc_955 N_A_835_93#_c_1317_n N_A_303_464#_c_1948_n 0.013725f $X=4.46 $Y=2.06
+ $X2=0 $Y2=0
cc_956 N_A_835_93#_c_1286_n N_A_303_464#_c_1948_n 0.00147857f $X=5.115 $Y=1.61
+ $X2=0 $Y2=0
cc_957 N_A_835_93#_c_1276_n N_A_303_464#_c_1940_n 0.00465542f $X=6.02 $Y=1.26
+ $X2=0 $Y2=0
cc_958 N_A_835_93#_c_1288_n N_A_303_464#_c_1950_n 0.00687903f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_959 N_A_835_93#_c_1289_n N_A_303_464#_c_1950_n 0.00443868f $X=6.55 $Y=3.15
+ $X2=0 $Y2=0
cc_960 N_A_835_93#_M1017_g N_A_303_464#_c_1950_n 4.63471e-19 $X=6.64 $Y=2.515
+ $X2=0 $Y2=0
cc_961 N_A_835_93#_c_1276_n N_A_303_464#_c_1941_n 0.0119509f $X=6.02 $Y=1.26
+ $X2=0 $Y2=0
cc_962 N_A_835_93#_c_1276_n N_A_303_464#_c_1942_n 0.0057513f $X=6.02 $Y=1.26
+ $X2=0 $Y2=0
cc_963 N_A_835_93#_c_1277_n N_A_303_464#_c_1942_n 7.71387e-19 $X=5.71 $Y=1.26
+ $X2=0 $Y2=0
cc_964 N_A_835_93#_M1017_g N_A_303_464#_c_1951_n 3.89682e-19 $X=6.64 $Y=2.515
+ $X2=0 $Y2=0
cc_965 N_A_835_93#_c_1288_n N_A_303_464#_c_1952_n 0.00126052f $X=5.615 $Y=3.075
+ $X2=0 $Y2=0
cc_966 N_A_835_93#_c_1277_n N_A_303_464#_c_1943_n 0.00420931f $X=5.71 $Y=1.26
+ $X2=0 $Y2=0
cc_967 N_A_835_93#_M1035_g N_A_303_464#_c_1945_n 0.00697619f $X=6.095 $Y=0.805
+ $X2=0 $Y2=0
cc_968 N_A_835_93#_c_1306_n N_VGND_M1029_d 0.0073489f $X=4.81 $Y=1.005 $X2=0
+ $Y2=0
cc_969 N_A_835_93#_c_1284_n N_VGND_M1029_d 0.00429495f $X=4.927 $Y=1.445 $X2=0
+ $Y2=0
cc_970 N_A_835_93#_c_1285_n N_VGND_c_2121_n 0.0156989f $X=4.45 $Y=0.625 $X2=0
+ $Y2=0
cc_971 N_A_835_93#_c_1275_n N_VGND_c_2122_n 0.0021556f $X=5.145 $Y=1.41 $X2=0
+ $Y2=0
cc_972 N_A_835_93#_c_1277_n N_VGND_c_2122_n 2.25445e-19 $X=5.71 $Y=1.26 $X2=0
+ $Y2=0
cc_973 N_A_835_93#_c_1306_n N_VGND_c_2122_n 0.0246763f $X=4.81 $Y=1.005 $X2=0
+ $Y2=0
cc_974 N_A_835_93#_c_1285_n N_VGND_c_2122_n 0.0135218f $X=4.45 $Y=0.625 $X2=0
+ $Y2=0
cc_975 N_A_835_93#_M1004_g N_VGND_c_2123_n 0.0018065f $X=9.785 $Y=0.58 $X2=0
+ $Y2=0
cc_976 N_A_835_93#_c_1285_n N_VGND_c_2126_n 0.0100041f $X=4.45 $Y=0.625 $X2=0
+ $Y2=0
cc_977 N_A_835_93#_M1004_g N_VGND_c_2131_n 0.00411612f $X=9.785 $Y=0.58 $X2=0
+ $Y2=0
cc_978 N_A_835_93#_c_1275_n N_VGND_c_2135_n 9.10391e-19 $X=5.145 $Y=1.41 $X2=0
+ $Y2=0
cc_979 N_A_835_93#_M1004_g N_VGND_c_2135_n 0.00752295f $X=9.785 $Y=0.58 $X2=0
+ $Y2=0
cc_980 N_A_835_93#_c_1285_n N_VGND_c_2135_n 0.0112422f $X=4.45 $Y=0.625 $X2=0
+ $Y2=0
cc_981 N_A_1997_272#_c_1467_n N_A_1745_74#_M1022_g 0.00755075f $X=11.175 $Y=0.58
+ $X2=0 $Y2=0
cc_982 N_A_1997_272#_c_1470_n N_A_1745_74#_M1022_g 0.00686241f $X=11.34 $Y=0.84
+ $X2=0 $Y2=0
cc_983 N_A_1997_272#_c_1471_n N_A_1745_74#_M1022_g 3.28981e-19 $X=11.65 $Y=1.445
+ $X2=0 $Y2=0
cc_984 N_A_1997_272#_c_1468_n N_A_1745_74#_c_1575_n 0.0096742f $X=11.565 $Y=1.53
+ $X2=0 $Y2=0
cc_985 N_A_1997_272#_c_1473_n N_A_1745_74#_c_1575_n 0.012401f $X=11.127 $Y=2.52
+ $X2=0 $Y2=0
cc_986 N_A_1997_272#_c_1474_n N_A_1745_74#_c_1575_n 0.00480843f $X=11.225
+ $Y=1.53 $X2=0 $Y2=0
cc_987 N_A_1997_272#_c_1477_n N_A_1745_74#_M1024_g 0.00777963f $X=11.11 $Y=2.75
+ $X2=0 $Y2=0
cc_988 N_A_1997_272#_c_1473_n N_A_1745_74#_M1024_g 0.0114263f $X=11.127 $Y=2.52
+ $X2=0 $Y2=0
cc_989 N_A_1997_272#_c_1468_n N_A_1745_74#_c_1576_n 0.00243079f $X=11.565
+ $Y=1.53 $X2=0 $Y2=0
cc_990 N_A_1997_272#_c_1469_n N_A_1745_74#_c_1576_n 0.00158858f $X=11.565
+ $Y=0.84 $X2=0 $Y2=0
cc_991 N_A_1997_272#_c_1471_n N_A_1745_74#_c_1576_n 0.0150077f $X=11.65 $Y=1.445
+ $X2=0 $Y2=0
cc_992 N_A_1997_272#_c_1466_n N_A_1745_74#_c_1577_n 0.00191851f $X=11.14 $Y=1.53
+ $X2=0 $Y2=0
cc_993 N_A_1997_272#_c_1469_n N_A_1745_74#_c_1577_n 0.00173828f $X=11.565
+ $Y=0.84 $X2=0 $Y2=0
cc_994 N_A_1997_272#_c_1470_n N_A_1745_74#_c_1577_n 0.00908089f $X=11.34 $Y=0.84
+ $X2=0 $Y2=0
cc_995 N_A_1997_272#_c_1471_n N_A_1745_74#_c_1577_n 0.00419353f $X=11.65
+ $Y=1.445 $X2=0 $Y2=0
cc_996 N_A_1997_272#_c_1474_n N_A_1745_74#_c_1577_n 0.00279652f $X=11.225
+ $Y=1.53 $X2=0 $Y2=0
cc_997 N_A_1997_272#_c_1468_n N_A_1745_74#_c_1587_n 0.00200907f $X=11.565
+ $Y=1.53 $X2=0 $Y2=0
cc_998 N_A_1997_272#_c_1473_n N_A_1745_74#_M1039_g 7.12087e-19 $X=11.127 $Y=2.52
+ $X2=0 $Y2=0
cc_999 N_A_1997_272#_c_1467_n N_A_1745_74#_M1027_g 0.00345625f $X=11.175 $Y=0.58
+ $X2=0 $Y2=0
cc_1000 N_A_1997_272#_c_1469_n N_A_1745_74#_M1027_g 0.00399686f $X=11.565
+ $Y=0.84 $X2=0 $Y2=0
cc_1001 N_A_1997_272#_c_1471_n N_A_1745_74#_M1027_g 0.00292154f $X=11.65
+ $Y=1.445 $X2=0 $Y2=0
cc_1002 N_A_1997_272#_c_1468_n N_A_1745_74#_c_1589_n 0.00289244f $X=11.565
+ $Y=1.53 $X2=0 $Y2=0
cc_1003 N_A_1997_272#_c_1473_n N_A_1745_74#_c_1589_n 0.00843513f $X=11.127
+ $Y=2.52 $X2=0 $Y2=0
cc_1004 N_A_1997_272#_M1037_g N_A_1745_74#_c_1590_n 0.0099993f $X=10.31 $Y=2.75
+ $X2=0 $Y2=0
cc_1005 N_A_1997_272#_M1003_g N_A_1745_74#_c_1580_n 5.63627e-19 $X=10.145
+ $Y=0.58 $X2=0 $Y2=0
cc_1006 N_A_1997_272#_c_1465_n N_A_1745_74#_c_1580_n 0.00475655f $X=10.31
+ $Y=1.84 $X2=0 $Y2=0
cc_1007 N_A_1997_272#_c_1472_n N_A_1745_74#_c_1580_n 0.0105779f $X=10.315
+ $Y=1.525 $X2=0 $Y2=0
cc_1008 N_A_1997_272#_c_1465_n N_A_1745_74#_c_1592_n 0.0112071f $X=10.31 $Y=1.84
+ $X2=0 $Y2=0
cc_1009 N_A_1997_272#_M1037_g N_A_1745_74#_c_1592_n 0.00484392f $X=10.31 $Y=2.75
+ $X2=0 $Y2=0
cc_1010 N_A_1997_272#_c_1472_n N_A_1745_74#_c_1592_n 0.0232183f $X=10.315
+ $Y=1.525 $X2=0 $Y2=0
cc_1011 N_A_1997_272#_M1037_g N_A_1745_74#_c_1594_n 0.016309f $X=10.31 $Y=2.75
+ $X2=0 $Y2=0
cc_1012 N_A_1997_272#_M1003_g N_A_1745_74#_c_1581_n 0.00279105f $X=10.145
+ $Y=0.58 $X2=0 $Y2=0
cc_1013 N_A_1997_272#_c_1466_n N_A_1745_74#_c_1583_n 0.00534862f $X=11.14
+ $Y=1.53 $X2=0 $Y2=0
cc_1014 N_A_1997_272#_c_1468_n N_A_1745_74#_c_1583_n 0.0057529f $X=11.565
+ $Y=1.53 $X2=0 $Y2=0
cc_1015 N_A_1997_272#_c_1469_n N_A_1745_74#_c_1583_n 0.00391205f $X=11.565
+ $Y=0.84 $X2=0 $Y2=0
cc_1016 N_A_1997_272#_c_1471_n N_A_1745_74#_c_1583_n 0.0139087f $X=11.65
+ $Y=1.445 $X2=0 $Y2=0
cc_1017 N_A_1997_272#_c_1474_n N_A_1745_74#_c_1583_n 0.0134734f $X=11.225
+ $Y=1.53 $X2=0 $Y2=0
cc_1018 N_A_1997_272#_M1003_g N_A_1745_74#_c_1584_n 0.0145056f $X=10.145 $Y=0.58
+ $X2=0 $Y2=0
cc_1019 N_A_1997_272#_c_1465_n N_A_1745_74#_c_1584_n 0.00481612f $X=10.31
+ $Y=1.84 $X2=0 $Y2=0
cc_1020 N_A_1997_272#_c_1466_n N_A_1745_74#_c_1584_n 0.0525955f $X=11.14 $Y=1.53
+ $X2=0 $Y2=0
cc_1021 N_A_1997_272#_c_1470_n N_A_1745_74#_c_1584_n 0.0263803f $X=11.34 $Y=0.84
+ $X2=0 $Y2=0
cc_1022 N_A_1997_272#_c_1472_n N_A_1745_74#_c_1584_n 0.023139f $X=10.315
+ $Y=1.525 $X2=0 $Y2=0
cc_1023 N_A_1997_272#_c_1468_n N_A_2402_424#_c_1733_n 9.19806e-19 $X=11.565
+ $Y=1.53 $X2=0 $Y2=0
cc_1024 N_A_1997_272#_c_1471_n N_A_2402_424#_c_1733_n 4.60428e-19 $X=11.65
+ $Y=1.445 $X2=0 $Y2=0
cc_1025 N_A_1997_272#_c_1469_n N_A_2402_424#_c_1735_n 0.00457908f $X=11.565
+ $Y=0.84 $X2=0 $Y2=0
cc_1026 N_A_1997_272#_c_1471_n N_A_2402_424#_c_1735_n 0.0171651f $X=11.65
+ $Y=1.445 $X2=0 $Y2=0
cc_1027 N_A_1997_272#_c_1468_n N_A_2402_424#_c_1737_n 0.00962353f $X=11.565
+ $Y=1.53 $X2=0 $Y2=0
cc_1028 N_A_1997_272#_c_1471_n N_A_2402_424#_c_1737_n 0.00719431f $X=11.65
+ $Y=1.445 $X2=0 $Y2=0
cc_1029 N_A_1997_272#_M1037_g N_VPWR_c_1783_n 0.00636044f $X=10.31 $Y=2.75 $X2=0
+ $Y2=0
cc_1030 N_A_1997_272#_c_1477_n N_VPWR_c_1783_n 0.0299965f $X=11.11 $Y=2.75 $X2=0
+ $Y2=0
cc_1031 N_A_1997_272#_c_1468_n N_VPWR_c_1784_n 0.0110105f $X=11.565 $Y=1.53
+ $X2=0 $Y2=0
cc_1032 N_A_1997_272#_c_1473_n N_VPWR_c_1784_n 0.0506546f $X=11.127 $Y=2.52
+ $X2=0 $Y2=0
cc_1033 N_A_1997_272#_M1037_g N_VPWR_c_1788_n 0.00454379f $X=10.31 $Y=2.75 $X2=0
+ $Y2=0
cc_1034 N_A_1997_272#_c_1477_n N_VPWR_c_1790_n 0.0156837f $X=11.11 $Y=2.75 $X2=0
+ $Y2=0
cc_1035 N_A_1997_272#_M1037_g N_VPWR_c_1776_n 0.00751043f $X=10.31 $Y=2.75 $X2=0
+ $Y2=0
cc_1036 N_A_1997_272#_c_1477_n N_VPWR_c_1776_n 0.0128663f $X=11.11 $Y=2.75 $X2=0
+ $Y2=0
cc_1037 N_A_1997_272#_c_1469_n N_VGND_M1027_s 0.00480139f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1038 N_A_1997_272#_M1003_g N_VGND_c_2123_n 0.01204f $X=10.145 $Y=0.58 $X2=0
+ $Y2=0
cc_1039 N_A_1997_272#_c_1467_n N_VGND_c_2123_n 0.0142227f $X=11.175 $Y=0.58
+ $X2=0 $Y2=0
cc_1040 N_A_1997_272#_c_1470_n N_VGND_c_2123_n 0.00176365f $X=11.34 $Y=0.84
+ $X2=0 $Y2=0
cc_1041 N_A_1997_272#_c_1467_n N_VGND_c_2124_n 0.0158614f $X=11.175 $Y=0.58
+ $X2=0 $Y2=0
cc_1042 N_A_1997_272#_c_1469_n N_VGND_c_2124_n 0.0143444f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1043 N_A_1997_272#_M1003_g N_VGND_c_2131_n 0.00383152f $X=10.145 $Y=0.58
+ $X2=0 $Y2=0
cc_1044 N_A_1997_272#_c_1467_n N_VGND_c_2132_n 0.0143883f $X=11.175 $Y=0.58
+ $X2=0 $Y2=0
cc_1045 N_A_1997_272#_c_1469_n N_VGND_c_2132_n 0.00329108f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1046 N_A_1997_272#_M1003_g N_VGND_c_2135_n 0.0075694f $X=10.145 $Y=0.58 $X2=0
+ $Y2=0
cc_1047 N_A_1997_272#_c_1467_n N_VGND_c_2135_n 0.0119301f $X=11.175 $Y=0.58
+ $X2=0 $Y2=0
cc_1048 N_A_1997_272#_c_1469_n N_VGND_c_2135_n 0.00670825f $X=11.565 $Y=0.84
+ $X2=0 $Y2=0
cc_1049 N_A_1745_74#_c_1576_n N_A_2402_424#_c_1733_n 0.00328297f $X=11.88
+ $Y=1.275 $X2=0 $Y2=0
cc_1050 N_A_1745_74#_M1039_g N_A_2402_424#_c_1739_n 0.0156493f $X=11.92 $Y=2.54
+ $X2=0 $Y2=0
cc_1051 N_A_1745_74#_M1027_g N_A_2402_424#_c_1735_n 0.0137683f $X=11.955
+ $Y=0.645 $X2=0 $Y2=0
cc_1052 N_A_1745_74#_c_1575_n N_A_2402_424#_c_1736_n 0.00247742f $X=11.32
+ $Y=1.84 $X2=0 $Y2=0
cc_1053 N_A_1745_74#_c_1587_n N_A_2402_424#_c_1736_n 0.0114621f $X=11.83
+ $Y=1.915 $X2=0 $Y2=0
cc_1054 N_A_1745_74#_c_1575_n N_A_2402_424#_c_1737_n 0.00108268f $X=11.32
+ $Y=1.84 $X2=0 $Y2=0
cc_1055 N_A_1745_74#_c_1576_n N_A_2402_424#_c_1737_n 5.99943e-19 $X=11.88
+ $Y=1.275 $X2=0 $Y2=0
cc_1056 N_A_1745_74#_c_1590_n N_VPWR_c_1783_n 0.0266532f $X=10.145 $Y=2.715
+ $X2=0 $Y2=0
cc_1057 N_A_1745_74#_c_1594_n N_VPWR_c_1783_n 0.00216546f $X=10.23 $Y=2.55 $X2=0
+ $Y2=0
cc_1058 N_A_1745_74#_M1024_g N_VPWR_c_1784_n 0.00993345f $X=11.335 $Y=2.75 $X2=0
+ $Y2=0
cc_1059 N_A_1745_74#_c_1587_n N_VPWR_c_1784_n 0.00608623f $X=11.83 $Y=1.915
+ $X2=0 $Y2=0
cc_1060 N_A_1745_74#_M1039_g N_VPWR_c_1784_n 0.00472774f $X=11.92 $Y=2.54 $X2=0
+ $Y2=0
cc_1061 N_A_1745_74#_M1039_g N_VPWR_c_1785_n 0.00478071f $X=11.92 $Y=2.54 $X2=0
+ $Y2=0
cc_1062 N_A_1745_74#_c_1590_n N_VPWR_c_1788_n 0.0274419f $X=10.145 $Y=2.715
+ $X2=0 $Y2=0
cc_1063 N_A_1745_74#_M1024_g N_VPWR_c_1790_n 0.00481245f $X=11.335 $Y=2.75 $X2=0
+ $Y2=0
cc_1064 N_A_1745_74#_M1039_g N_VPWR_c_1795_n 0.005209f $X=11.92 $Y=2.54 $X2=0
+ $Y2=0
cc_1065 N_A_1745_74#_M1024_g N_VPWR_c_1776_n 0.00855303f $X=11.335 $Y=2.75 $X2=0
+ $Y2=0
cc_1066 N_A_1745_74#_M1039_g N_VPWR_c_1776_n 0.00987945f $X=11.92 $Y=2.54 $X2=0
+ $Y2=0
cc_1067 N_A_1745_74#_c_1590_n N_VPWR_c_1776_n 0.0332915f $X=10.145 $Y=2.715
+ $X2=0 $Y2=0
cc_1068 N_A_1745_74#_c_1590_n A_1996_508# 0.00356223f $X=10.145 $Y=2.715
+ $X2=-0.19 $Y2=-0.245
cc_1069 N_A_1745_74#_c_1581_n N_VGND_c_2123_n 0.0159689f $X=9.57 $Y=0.56 $X2=0
+ $Y2=0
cc_1070 N_A_1745_74#_c_1584_n N_VGND_c_2123_n 0.0191133f $X=11.065 $Y=1.185
+ $X2=0 $Y2=0
cc_1071 N_A_1745_74#_M1022_g N_VGND_c_2124_n 0.00322527f $X=10.96 $Y=0.58 $X2=0
+ $Y2=0
cc_1072 N_A_1745_74#_c_1576_n N_VGND_c_2124_n 0.00195495f $X=11.88 $Y=1.275
+ $X2=0 $Y2=0
cc_1073 N_A_1745_74#_M1027_g N_VGND_c_2124_n 0.00927494f $X=11.955 $Y=0.645
+ $X2=0 $Y2=0
cc_1074 N_A_1745_74#_M1027_g N_VGND_c_2125_n 0.00296233f $X=11.955 $Y=0.645
+ $X2=0 $Y2=0
cc_1075 N_A_1745_74#_c_1581_n N_VGND_c_2131_n 0.0151251f $X=9.57 $Y=0.56 $X2=0
+ $Y2=0
cc_1076 N_A_1745_74#_M1022_g N_VGND_c_2132_n 0.00434272f $X=10.96 $Y=0.58 $X2=0
+ $Y2=0
cc_1077 N_A_1745_74#_M1027_g N_VGND_c_2133_n 0.00383152f $X=11.955 $Y=0.645
+ $X2=0 $Y2=0
cc_1078 N_A_1745_74#_M1022_g N_VGND_c_2135_n 0.00825669f $X=10.96 $Y=0.58 $X2=0
+ $Y2=0
cc_1079 N_A_1745_74#_M1027_g N_VGND_c_2135_n 0.00762539f $X=11.955 $Y=0.645
+ $X2=0 $Y2=0
cc_1080 N_A_1745_74#_c_1581_n N_VGND_c_2135_n 0.0125365f $X=9.57 $Y=0.56 $X2=0
+ $Y2=0
cc_1081 N_A_2402_424#_c_1739_n N_VPWR_c_1784_n 0.0345631f $X=12.145 $Y=2.265
+ $X2=0 $Y2=0
cc_1082 N_A_2402_424#_M1011_g N_VPWR_c_1785_n 0.0243126f $X=12.93 $Y=2.4 $X2=0
+ $Y2=0
cc_1083 N_A_2402_424#_c_1733_n N_VPWR_c_1785_n 0.00687596f $X=12.84 $Y=1.465
+ $X2=0 $Y2=0
cc_1084 N_A_2402_424#_c_1757_p N_VPWR_c_1785_n 0.0252753f $X=12.745 $Y=1.465
+ $X2=0 $Y2=0
cc_1085 N_A_2402_424#_c_1736_n N_VPWR_c_1785_n 0.0776078f $X=12.145 $Y=2.1 $X2=0
+ $Y2=0
cc_1086 N_A_2402_424#_c_1739_n N_VPWR_c_1795_n 0.014549f $X=12.145 $Y=2.265
+ $X2=0 $Y2=0
cc_1087 N_A_2402_424#_M1011_g N_VPWR_c_1796_n 0.00460063f $X=12.93 $Y=2.4 $X2=0
+ $Y2=0
cc_1088 N_A_2402_424#_M1011_g N_VPWR_c_1776_n 0.00912313f $X=12.93 $Y=2.4 $X2=0
+ $Y2=0
cc_1089 N_A_2402_424#_c_1739_n N_VPWR_c_1776_n 0.0119743f $X=12.145 $Y=2.265
+ $X2=0 $Y2=0
cc_1090 N_A_2402_424#_M1007_g Q 0.00853833f $X=12.945 $Y=0.74 $X2=0 $Y2=0
cc_1091 N_A_2402_424#_M1007_g Q 0.00343176f $X=12.945 $Y=0.74 $X2=0 $Y2=0
cc_1092 N_A_2402_424#_M1007_g Q 0.0270842f $X=12.945 $Y=0.74 $X2=0 $Y2=0
cc_1093 N_A_2402_424#_c_1757_p Q 0.0238691f $X=12.745 $Y=1.465 $X2=0 $Y2=0
cc_1094 N_A_2402_424#_c_1735_n N_VGND_c_2124_n 0.00917009f $X=12.17 $Y=0.645
+ $X2=0 $Y2=0
cc_1095 N_A_2402_424#_M1007_g N_VGND_c_2125_n 0.00647412f $X=12.945 $Y=0.74
+ $X2=0 $Y2=0
cc_1096 N_A_2402_424#_c_1733_n N_VGND_c_2125_n 0.00577732f $X=12.84 $Y=1.465
+ $X2=0 $Y2=0
cc_1097 N_A_2402_424#_c_1735_n N_VGND_c_2125_n 0.0504216f $X=12.17 $Y=0.645
+ $X2=0 $Y2=0
cc_1098 N_A_2402_424#_c_1757_p N_VGND_c_2125_n 0.0209147f $X=12.745 $Y=1.465
+ $X2=0 $Y2=0
cc_1099 N_A_2402_424#_c_1735_n N_VGND_c_2133_n 0.011066f $X=12.17 $Y=0.645 $X2=0
+ $Y2=0
cc_1100 N_A_2402_424#_M1007_g N_VGND_c_2134_n 0.00434272f $X=12.945 $Y=0.74
+ $X2=0 $Y2=0
cc_1101 N_A_2402_424#_M1007_g N_VGND_c_2135_n 0.00828941f $X=12.945 $Y=0.74
+ $X2=0 $Y2=0
cc_1102 N_A_2402_424#_c_1735_n N_VGND_c_2135_n 0.00915947f $X=12.17 $Y=0.645
+ $X2=0 $Y2=0
cc_1103 N_VPWR_c_1777_n N_A_303_464#_c_1946_n 0.0195189f $X=0.78 $Y=2.465 $X2=0
+ $Y2=0
cc_1104 N_VPWR_c_1793_n N_A_303_464#_c_1946_n 0.0470186f $X=3.095 $Y=3.33 $X2=0
+ $Y2=0
cc_1105 N_VPWR_c_1776_n N_A_303_464#_c_1946_n 0.0389581f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1106 N_VPWR_M1019_d N_A_303_464#_c_1968_n 0.00999698f $X=3.125 $Y=2.32 $X2=0
+ $Y2=0
cc_1107 N_VPWR_c_1778_n N_A_303_464#_c_1968_n 0.0213283f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1108 N_VPWR_c_1776_n N_A_303_464#_c_1968_n 0.018952f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1109 N_VPWR_M1018_d N_A_303_464#_c_1948_n 0.00357521f $X=4.735 $Y=1.935 $X2=0
+ $Y2=0
cc_1110 N_VPWR_c_1779_n N_A_303_464#_c_1948_n 0.0162896f $X=4.87 $Y=2.885 $X2=0
+ $Y2=0
cc_1111 N_VPWR_c_1786_n N_A_303_464#_c_1948_n 0.0104512f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1112 N_VPWR_c_1794_n N_A_303_464#_c_1948_n 0.0114056f $X=7.205 $Y=3.33 $X2=0
+ $Y2=0
cc_1113 N_VPWR_c_1776_n N_A_303_464#_c_1948_n 0.0393494f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1114 N_VPWR_M1019_d N_A_303_464#_c_1949_n 4.92358e-19 $X=3.125 $Y=2.32 $X2=0
+ $Y2=0
cc_1115 N_VPWR_c_1776_n N_A_303_464#_c_1949_n 0.00747731f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1116 N_VPWR_c_1794_n N_A_303_464#_c_1950_n 0.00531602f $X=7.205 $Y=3.33 $X2=0
+ $Y2=0
cc_1117 N_VPWR_c_1776_n N_A_303_464#_c_1950_n 0.00673278f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1118 N_VPWR_c_1778_n N_A_303_464#_c_1954_n 0.00906618f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1119 N_VPWR_c_1778_n N_A_303_464#_c_1955_n 0.0176067f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1120 N_VPWR_c_1786_n N_A_303_464#_c_1955_n 0.0144363f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1121 N_VPWR_c_1776_n N_A_303_464#_c_1955_n 0.0119305f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1122 N_VPWR_c_1785_n Q 0.0395727f $X=12.705 $Y=1.985 $X2=0 $Y2=0
cc_1123 N_VPWR_c_1796_n Q 0.0112891f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1124 N_VPWR_c_1776_n Q 0.00934413f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1125 N_A_303_464#_c_1968_n A_535_464# 0.00890703f $X=3.445 $Y=2.43 $X2=-0.19
+ $Y2=-0.245
cc_1126 N_A_303_464#_M1009_d N_noxref_24_c_2252_n 0.0106902f $X=1.95 $Y=0.405
+ $X2=0 $Y2=0
cc_1127 N_A_303_464#_c_1937_n N_noxref_24_c_2252_n 0.0126305f $X=3.445 $Y=1.005
+ $X2=0 $Y2=0
cc_1128 N_A_303_464#_c_1944_n N_noxref_24_c_2252_n 0.019982f $X=2.435 $Y=0.68
+ $X2=0 $Y2=0
cc_1129 N_A_303_464#_c_1937_n N_noxref_24_c_2254_n 0.0234737f $X=3.445 $Y=1.005
+ $X2=0 $Y2=0
cc_1130 N_A_303_464#_c_1944_n N_noxref_24_c_2254_n 0.00520956f $X=2.435 $Y=0.68
+ $X2=0 $Y2=0
cc_1131 Q N_VGND_c_2125_n 0.0293763f $X=13.115 $Y=0.47 $X2=0 $Y2=0
cc_1132 Q N_VGND_c_2134_n 0.0145639f $X=13.115 $Y=0.47 $X2=0 $Y2=0
cc_1133 Q N_VGND_c_2135_n 0.0119984f $X=13.115 $Y=0.47 $X2=0 $Y2=0
cc_1134 N_VGND_c_2129_n N_noxref_24_c_2252_n 0.10468f $X=3.59 $Y=0 $X2=0 $Y2=0
cc_1135 N_VGND_c_2135_n N_noxref_24_c_2252_n 0.0610965f $X=13.2 $Y=0 $X2=0 $Y2=0
cc_1136 N_VGND_c_2120_n N_noxref_24_c_2253_n 0.0259562f $X=0.71 $Y=0.65 $X2=0
+ $Y2=0
cc_1137 N_VGND_c_2129_n N_noxref_24_c_2253_n 0.0225398f $X=3.59 $Y=0 $X2=0 $Y2=0
cc_1138 N_VGND_c_2135_n N_noxref_24_c_2253_n 0.0125704f $X=13.2 $Y=0 $X2=0 $Y2=0
cc_1139 N_VGND_c_2121_n N_noxref_24_c_2254_n 0.0118481f $X=3.715 $Y=0.565 $X2=0
+ $Y2=0
cc_1140 N_VGND_c_2129_n N_noxref_24_c_2254_n 0.0243596f $X=3.59 $Y=0 $X2=0 $Y2=0
cc_1141 N_VGND_c_2135_n N_noxref_24_c_2254_n 0.0134194f $X=13.2 $Y=0 $X2=0 $Y2=0
cc_1142 N_noxref_24_c_2252_n noxref_25 0.00198134f $X=3.06 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1143 N_noxref_24_c_2252_n noxref_26 0.00226367f $X=3.06 $Y=0.34 $X2=-0.19
+ $Y2=-0.245

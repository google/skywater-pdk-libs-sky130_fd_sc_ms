* File: sky130_fd_sc_ms__a32oi_2.pex.spice
* Created: Wed Sep  2 11:56:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A32OI_2%B2 3 7 11 15 19 22 29 34
r48 28 29 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=0.975 $Y=1.465
+ $X2=1.005 $Y2=1.465
r49 24 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.465
+ $X2=0.51 $Y2=1.465
r50 22 34 4.04332 $w=4.78e-07 $l=1.15e-07 $layer=LI1_cond $X=0.24 $Y=1.54
+ $X2=0.355 $Y2=1.54
r51 20 28 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=0.925 $Y=1.465
+ $X2=0.975 $Y2=1.465
r52 20 26 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=0.925 $Y=1.465
+ $X2=0.51 $Y2=1.465
r53 19 34 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=0.925 $Y=1.465
+ $X2=0.355 $Y2=1.465
r54 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.925
+ $Y=1.465 $X2=0.925 $Y2=1.465
r55 13 29 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.63
+ $X2=1.005 $Y2=1.465
r56 13 15 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.005 $Y=1.63
+ $X2=1.005 $Y2=2.4
r57 9 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.3
+ $X2=0.975 $Y2=1.465
r58 9 11 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.975 $Y=1.3
+ $X2=0.975 $Y2=0.74
r59 5 26 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.63
+ $X2=0.51 $Y2=1.465
r60 5 7 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.51 $Y=1.63 $X2=0.51
+ $Y2=2.4
r61 1 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.465
r62 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_2%B1 1 3 6 8 10 13 15 16 22
c56 13 0 1.72332e-19 $X=2.005 $Y=2.4
c57 8 0 1.33933e-19 $X=1.835 $Y=1.22
c58 1 0 8.87788e-21 $X=1.405 $Y=1.22
r59 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.01
+ $Y=1.385 $X2=2.01 $Y2=1.385
r60 22 24 0.77492 $w=3.11e-07 $l=5e-09 $layer=POLY_cond $X=2.005 $Y=1.385
+ $X2=2.01 $Y2=1.385
r61 21 22 26.3473 $w=3.11e-07 $l=1.7e-07 $layer=POLY_cond $X=1.835 $Y=1.385
+ $X2=2.005 $Y2=1.385
r62 20 21 51.1447 $w=3.11e-07 $l=3.3e-07 $layer=POLY_cond $X=1.505 $Y=1.385
+ $X2=1.835 $Y2=1.385
r63 16 25 4.67207 $w=3.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.16 $Y=1.365
+ $X2=2.01 $Y2=1.365
r64 15 25 10.2785 $w=3.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=2.01 $Y2=1.365
r65 11 22 15.5536 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.005 $Y=1.55
+ $X2=2.005 $Y2=1.385
r66 11 13 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.005 $Y=1.55
+ $X2=2.005 $Y2=2.4
r67 8 21 19.8172 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=1.22
+ $X2=1.835 $Y2=1.385
r68 8 10 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.835 $Y=1.22
+ $X2=1.835 $Y2=0.74
r69 4 20 15.5536 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.505 $Y=1.55
+ $X2=1.505 $Y2=1.385
r70 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.505 $Y=1.55
+ $X2=1.505 $Y2=2.4
r71 1 20 15.4984 $w=3.11e-07 $l=2.09105e-07 $layer=POLY_cond $X=1.405 $Y=1.22
+ $X2=1.505 $Y2=1.385
r72 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.405 $Y=1.22 $X2=1.405
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_2%A1 3 5 7 8 10 13 15 24
c57 15 0 1.33933e-19 $X=2.64 $Y=1.295
c58 13 0 1.57199e-19 $X=3.345 $Y=2.4
r59 23 24 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.325 $Y=1.385
+ $X2=3.345 $Y2=1.385
r60 22 23 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.895 $Y=1.385
+ $X2=3.325 $Y2=1.385
r61 20 22 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=2.61 $Y=1.385
+ $X2=2.895 $Y2=1.385
r62 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.385 $X2=2.61 $Y2=1.385
r63 17 20 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=2.505 $Y=1.385
+ $X2=2.61 $Y2=1.385
r64 15 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.61 $Y=1.295 $X2=2.61
+ $Y2=1.385
r65 11 24 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.345 $Y=1.55
+ $X2=3.345 $Y2=1.385
r66 11 13 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.345 $Y=1.55
+ $X2=3.345 $Y2=2.4
r67 8 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.325 $Y=1.22
+ $X2=3.325 $Y2=1.385
r68 8 10 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.325 $Y=1.22
+ $X2=3.325 $Y2=0.74
r69 5 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.895 $Y=1.22
+ $X2=2.895 $Y2=1.385
r70 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.895 $Y=1.22 $X2=2.895
+ $Y2=0.74
r71 1 17 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.505 $Y=1.55
+ $X2=2.505 $Y2=1.385
r72 1 3 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.505 $Y=1.55
+ $X2=2.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_2%A2 3 7 11 15 18 19 20 21 22 27
c57 27 0 4.79191e-20 $X=4.21 $Y=1.515
c58 18 0 1.39445e-19 $X=3.795 $Y=1.515
c59 11 0 1.89611e-19 $X=4.31 $Y=2.4
c60 3 0 5.89156e-20 $X=3.78 $Y=0.74
r61 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.21
+ $Y=1.515 $X2=4.21 $Y2=1.515
r62 22 27 3.48413 $w=4.28e-07 $l=1.3e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=4.21 $Y2=1.565
r63 21 22 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=4.08 $Y2=1.565
r64 19 26 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=4.22 $Y=1.515 $X2=4.21
+ $Y2=1.515
r65 19 20 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.22 $Y=1.515 $X2=4.31
+ $Y2=1.515
r66 17 26 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=3.885 $Y=1.515
+ $X2=4.21 $Y2=1.515
r67 17 18 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.885 $Y=1.515
+ $X2=3.795 $Y2=1.515
r68 13 20 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=4.325 $Y=1.35
+ $X2=4.31 $Y2=1.515
r69 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.325 $Y=1.35
+ $X2=4.325 $Y2=0.74
r70 9 20 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=4.31 $Y=1.68
+ $X2=4.31 $Y2=1.515
r71 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.31 $Y=1.68 $X2=4.31
+ $Y2=2.4
r72 5 18 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=3.795 $Y=1.68
+ $X2=3.795 $Y2=1.515
r73 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.795 $Y=1.68
+ $X2=3.795 $Y2=2.4
r74 1 18 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=3.78 $Y=1.35
+ $X2=3.795 $Y2=1.515
r75 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.78 $Y=1.35 $X2=3.78
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_2%A3 3 5 7 10 12 14 15 23
c41 3 0 4.79191e-20 $X=4.935 $Y=2.4
r42 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.95
+ $Y=1.385 $X2=5.95 $Y2=1.385
r43 21 23 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=5.745 $Y=1.385
+ $X2=5.95 $Y2=1.385
r44 20 21 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=5.485 $Y=1.385
+ $X2=5.745 $Y2=1.385
r45 19 20 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=5.315 $Y=1.385
+ $X2=5.485 $Y2=1.385
r46 17 19 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=4.935 $Y=1.385
+ $X2=5.315 $Y2=1.385
r47 15 24 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.95 $Y=1.295 $X2=5.95
+ $Y2=1.385
r48 12 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.745 $Y=1.22
+ $X2=5.745 $Y2=1.385
r49 12 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.745 $Y=1.22
+ $X2=5.745 $Y2=0.74
r50 8 20 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.485 $Y=1.55
+ $X2=5.485 $Y2=1.385
r51 8 10 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=5.485 $Y=1.55
+ $X2=5.485 $Y2=2.4
r52 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.315 $Y=1.22
+ $X2=5.315 $Y2=1.385
r53 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.315 $Y=1.22 $X2=5.315
+ $Y2=0.74
r54 1 17 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.935 $Y=1.55
+ $X2=4.935 $Y2=1.385
r55 1 3 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=4.935 $Y=1.55
+ $X2=4.935 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_2%A_27_368# 1 2 3 4 5 6 21 25 26 29 31 33 37
+ 41 43 45 47 49 53 57 60
c85 41 0 3.4681e-19 $X=3.57 $Y=2.465
r86 68 69 1.59269 $w=3.83e-07 $l=5e-08 $layer=LI1_cond $X=4.647 $Y=1.985
+ $X2=4.647 $Y2=2.035
r87 66 68 5.73368 $w=3.83e-07 $l=1.8e-07 $layer=LI1_cond $X=4.647 $Y=1.805
+ $X2=4.647 $Y2=1.985
r88 64 65 3.21434 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=2.145
+ $X2=3.57 $Y2=2.23
r89 63 64 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=3.57 $Y=2.115 $X2=3.57
+ $Y2=2.145
r90 60 63 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.57 $Y=2.035 $X2=3.57
+ $Y2=2.115
r91 53 55 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=5.71 $Y=1.985
+ $X2=5.71 $Y2=2.815
r92 51 53 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=5.71 $Y=1.89
+ $X2=5.71 $Y2=1.985
r93 50 66 5.51523 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=4.875 $Y=1.805
+ $X2=4.647 $Y2=1.805
r94 49 51 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.545 $Y=1.805
+ $X2=5.71 $Y2=1.89
r95 49 50 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.545 $Y=1.805
+ $X2=4.875 $Y2=1.805
r96 45 69 2.6202 $w=4.55e-07 $l=8.5e-08 $layer=LI1_cond $X=4.647 $Y=2.12
+ $X2=4.647 $Y2=2.035
r97 45 47 7.36048 $w=4.53e-07 $l=2.8e-07 $layer=LI1_cond $X=4.647 $Y=2.12
+ $X2=4.647 $Y2=2.4
r98 44 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.735 $Y=2.035
+ $X2=3.57 $Y2=2.035
r99 43 69 5.51523 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=4.42 $Y=2.035
+ $X2=4.647 $Y2=2.035
r100 43 44 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=4.42 $Y=2.035
+ $X2=3.735 $Y2=2.035
r101 41 65 9.5026 $w=2.83e-07 $l=2.35e-07 $layer=LI1_cond $X=3.592 $Y=2.465
+ $X2=3.592 $Y2=2.23
r102 38 59 4.64039 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=2.4 $Y=2.145
+ $X2=2.257 $Y2=2.145
r103 37 64 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=2.145
+ $X2=3.57 $Y2=2.145
r104 37 38 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=3.405 $Y=2.145
+ $X2=2.4 $Y2=2.145
r105 34 36 16.579 $w=2.83e-07 $l=4.1e-07 $layer=LI1_cond $X=2.257 $Y=2.905
+ $X2=2.257 $Y2=2.495
r106 33 59 2.75828 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.257 $Y=2.23
+ $X2=2.257 $Y2=2.145
r107 33 36 10.7157 $w=2.83e-07 $l=2.65e-07 $layer=LI1_cond $X=2.257 $Y=2.23
+ $X2=2.257 $Y2=2.495
r108 32 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=2.99
+ $X2=1.28 $Y2=2.99
r109 31 34 7.39867 $w=1.7e-07 $l=1.79538e-07 $layer=LI1_cond $X=2.115 $Y=2.99
+ $X2=2.257 $Y2=2.905
r110 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.115 $Y=2.99
+ $X2=1.445 $Y2=2.99
r111 27 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=2.905
+ $X2=1.28 $Y2=2.99
r112 27 29 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.28 $Y=2.905
+ $X2=1.28 $Y2=2.27
r113 25 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=2.99
+ $X2=1.28 $Y2=2.99
r114 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=2.99
+ $X2=0.445 $Y2=2.99
r115 21 24 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.28 $Y=2.115
+ $X2=0.28 $Y2=2.815
r116 19 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.445 $Y2=2.99
r117 19 24 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.28 $Y2=2.815
r118 6 55 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.575
+ $Y=1.84 $X2=5.71 $Y2=2.815
r119 6 53 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.575
+ $Y=1.84 $X2=5.71 $Y2=1.985
r120 5 68 600 $w=1.7e-07 $l=3.75566e-07 $layer=licon1_PDIFF $count=1 $X=4.4
+ $Y=1.84 $X2=4.71 $Y2=1.985
r121 5 47 300 $w=1.7e-07 $l=6.4591e-07 $layer=licon1_PDIFF $count=2 $X=4.4
+ $Y=1.84 $X2=4.585 $Y2=2.4
r122 4 63 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=3.435
+ $Y=1.84 $X2=3.57 $Y2=2.115
r123 4 41 300 $w=1.7e-07 $l=6.89202e-07 $layer=licon1_PDIFF $count=2 $X=3.435
+ $Y=1.84 $X2=3.57 $Y2=2.465
r124 3 59 600 $w=1.7e-07 $l=3.86588e-07 $layer=licon1_PDIFF $count=1 $X=2.095
+ $Y=1.84 $X2=2.28 $Y2=2.145
r125 3 36 300 $w=1.7e-07 $l=7.41755e-07 $layer=licon1_PDIFF $count=2 $X=2.095
+ $Y=1.84 $X2=2.28 $Y2=2.495
r126 2 29 300 $w=1.7e-07 $l=5.14247e-07 $layer=licon1_PDIFF $count=2 $X=1.095
+ $Y=1.84 $X2=1.28 $Y2=2.27
r127 1 24 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r128 1 21 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_2%Y 1 2 3 4 13 15 17 23 25 27 29 34 38 42 43
+ 44 47 50
c80 44 0 1.39445e-19 $X=3.035 $Y=1.58
c81 43 0 5.89156e-20 $X=3.12 $Y=1.235
c82 25 0 8.87788e-21 $X=3.005 $Y=0.925
r83 47 50 2.75584 $w=2.28e-07 $l=5.5e-08 $layer=LI1_cond $X=3.12 $Y=1.72
+ $X2=3.12 $Y2=1.665
r84 44 47 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=1.805 $X2=3.12
+ $Y2=1.72
r85 44 50 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.12 $Y=1.65
+ $X2=3.12 $Y2=1.665
r86 42 44 15.0319 $w=2.28e-07 $l=3e-07 $layer=LI1_cond $X=3.12 $Y=1.35 $X2=3.12
+ $Y2=1.65
r87 42 43 5.98911 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=1.35
+ $X2=3.12 $Y2=1.235
r88 40 41 10.3763 $w=1.94e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=0.76
+ $X2=3.105 $Y2=0.925
r89 34 36 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=1.62 $Y=0.8
+ $X2=1.62 $Y2=0.925
r90 29 41 5.185 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.105 $Y=1.01 $X2=3.105
+ $Y2=0.925
r91 29 43 12.4773 $w=1.98e-07 $l=2.25e-07 $layer=LI1_cond $X=3.105 $Y=1.01
+ $X2=3.105 $Y2=1.235
r92 28 38 8.61065 $w=1.7e-07 $l=1.83916e-07 $layer=LI1_cond $X=1.945 $Y=1.805
+ $X2=1.78 $Y2=1.845
r93 27 44 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.005 $Y=1.805
+ $X2=3.12 $Y2=1.805
r94 27 28 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=3.005 $Y=1.805
+ $X2=1.945 $Y2=1.805
r95 26 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=0.925
+ $X2=1.62 $Y2=0.925
r96 25 41 1.50975 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.005 $Y=0.925
+ $X2=3.105 $Y2=0.925
r97 25 26 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=3.005 $Y=0.925
+ $X2=1.785 $Y2=0.925
r98 21 38 0.89609 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=1.78 $Y=1.97
+ $X2=1.78 $Y2=1.845
r99 21 23 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.78 $Y=1.97
+ $X2=1.78 $Y2=2.65
r100 18 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=1.885
+ $X2=0.78 $Y2=1.885
r101 17 38 8.61065 $w=1.7e-07 $l=1.83916e-07 $layer=LI1_cond $X=1.615 $Y=1.885
+ $X2=1.78 $Y2=1.845
r102 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=1.885
+ $X2=0.945 $Y2=1.885
r103 13 32 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=1.97 $X2=0.78
+ $Y2=1.885
r104 13 15 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.78 $Y=1.97
+ $X2=0.78 $Y2=2.645
r105 4 23 400 $w=1.7e-07 $l=8.97747e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.84 $X2=1.78 $Y2=2.65
r106 4 21 400 $w=1.7e-07 $l=2.41402e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.84 $X2=1.78 $Y2=1.97
r107 3 32 400 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.84 $X2=0.78 $Y2=1.965
r108 3 15 400 $w=1.7e-07 $l=8.90463e-07 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.84 $X2=0.78 $Y2=2.645
r109 2 40 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=2.97
+ $Y=0.37 $X2=3.11 $Y2=0.76
r110 1 34 182 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_NDIFF $count=1 $X=1.48
+ $Y=0.37 $X2=1.62 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_2%VPWR 1 2 3 12 16 20 25 26 27 29 34 44 45 48
+ 53
c68 12 0 1.72332e-19 $X=3.115 $Y=2.495
r69 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r70 48 51 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r71 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r72 42 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r73 42 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.08 $Y2=3.33
r74 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r75 39 53 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=4.25 $Y=3.33
+ $X2=4.077 $Y2=3.33
r76 39 41 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.25 $Y=3.33
+ $X2=5.04 $Y2=3.33
r77 38 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r78 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r79 35 48 13.764 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=3.28 $Y=3.33
+ $X2=2.925 $Y2=3.33
r80 35 37 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.28 $Y=3.33 $X2=3.6
+ $Y2=3.33
r81 34 53 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=4.077 $Y2=3.33
r82 34 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=3.6 $Y2=3.33
r83 32 51 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=2.64 $Y2=3.33
r84 31 32 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r85 29 48 13.764 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=2.57 $Y=3.33
+ $X2=2.925 $Y2=3.33
r86 29 31 152.011 $w=1.68e-07 $l=2.33e-06 $layer=LI1_cond $X=2.57 $Y=3.33
+ $X2=0.24 $Y2=3.33
r87 27 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r88 27 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r89 27 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r90 25 41 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.045 $Y=3.33
+ $X2=5.04 $Y2=3.33
r91 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.045 $Y=3.33
+ $X2=5.21 $Y2=3.33
r92 24 44 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=5.375 $Y=3.33 $X2=6
+ $Y2=3.33
r93 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.375 $Y=3.33
+ $X2=5.21 $Y2=3.33
r94 20 23 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.21 $Y=2.155
+ $X2=5.21 $Y2=2.835
r95 18 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.21 $Y=3.245
+ $X2=5.21 $Y2=3.33
r96 18 23 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=5.21 $Y=3.245
+ $X2=5.21 $Y2=2.835
r97 14 53 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=4.077 $Y=3.245
+ $X2=4.077 $Y2=3.33
r98 14 16 29.0616 $w=3.43e-07 $l=8.7e-07 $layer=LI1_cond $X=4.077 $Y=3.245
+ $X2=4.077 $Y2=2.375
r99 10 48 2.89202 $w=7.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=3.245
+ $X2=2.925 $Y2=3.33
r100 10 12 12.6346 $w=7.08e-07 $l=7.5e-07 $layer=LI1_cond $X=2.925 $Y=3.245
+ $X2=2.925 $Y2=2.495
r101 3 23 400 $w=1.7e-07 $l=1.08356e-06 $layer=licon1_PDIFF $count=1 $X=5.025
+ $Y=1.84 $X2=5.21 $Y2=2.835
r102 3 20 400 $w=1.7e-07 $l=3.96863e-07 $layer=licon1_PDIFF $count=1 $X=5.025
+ $Y=1.84 $X2=5.21 $Y2=2.155
r103 2 16 300 $w=1.7e-07 $l=6.22796e-07 $layer=licon1_PDIFF $count=2 $X=3.885
+ $Y=1.84 $X2=4.075 $Y2=2.375
r104 1 12 150 $w=1.7e-07 $l=8.77283e-07 $layer=licon1_PDIFF $count=4 $X=2.595
+ $Y=1.84 $X2=3.115 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_2%A_27_74# 1 2 3 12 14 15 20 21 22
r37 22 25 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.12 $Y=0.34
+ $X2=2.12 $Y2=0.55
r38 20 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=0.34
+ $X2=2.12 $Y2=0.34
r39 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.955 $Y=0.34
+ $X2=1.275 $Y2=0.34
r40 17 19 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.19 $Y=0.96
+ $X2=1.19 $Y2=0.515
r41 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.19 $Y=0.425
+ $X2=1.275 $Y2=0.34
r42 16 19 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.19 $Y=0.425 $X2=1.19
+ $Y2=0.515
r43 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.105 $Y=1.045
+ $X2=1.19 $Y2=0.96
r44 14 15 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.105 $Y=1.045
+ $X2=0.365 $Y2=1.045
r45 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.96
+ $X2=0.365 $Y2=1.045
r46 10 12 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.24 $Y=0.96
+ $X2=0.24 $Y2=0.515
r47 3 25 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=1.91
+ $Y=0.37 $X2=2.12 $Y2=0.55
r48 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.05
+ $Y=0.37 $X2=1.19 $Y2=0.515
r49 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_2%VGND 1 2 3 12 16 18 20 22 24 29 37 43 46 50
r67 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r68 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r69 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r70 41 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r71 41 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r72 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r73 38 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.185 $Y=0 $X2=5.06
+ $Y2=0
r74 38 40 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.185 $Y=0 $X2=5.52
+ $Y2=0
r75 37 49 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=5.795 $Y=0 $X2=6.017
+ $Y2=0
r76 37 40 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.795 $Y=0 $X2=5.52
+ $Y2=0
r77 36 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r78 35 36 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r79 33 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r80 32 35 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=4.56
+ $Y2=0
r81 32 33 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r82 30 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r83 30 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r84 29 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.935 $Y=0 $X2=5.06
+ $Y2=0
r85 29 35 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.935 $Y=0 $X2=4.56
+ $Y2=0
r86 27 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r87 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r88 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r89 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r90 22 36 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.56
+ $Y2=0
r91 22 33 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=1.2
+ $Y2=0
r92 18 49 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.96 $Y=0.085
+ $X2=6.017 $Y2=0
r93 18 20 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.96 $Y=0.085
+ $X2=5.96 $Y2=0.515
r94 14 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.06 $Y=0.085
+ $X2=5.06 $Y2=0
r95 14 16 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=5.06 $Y=0.085
+ $X2=5.06 $Y2=0.675
r96 10 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r97 10 12 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.625
r98 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.82
+ $Y=0.37 $X2=5.96 $Y2=0.515
r99 2 16 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=4.955
+ $Y=0.37 $X2=5.1 $Y2=0.675
r100 1 12 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_2%A_507_74# 1 2 3 10 14 16 20 22 27
r44 22 25 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.68 $Y=0.34
+ $X2=2.68 $Y2=0.55
r45 18 20 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=4.54 $Y=0.425
+ $X2=4.54 $Y2=0.675
r46 17 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=0.34
+ $X2=3.54 $Y2=0.34
r47 16 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.375 $Y=0.34
+ $X2=4.54 $Y2=0.425
r48 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.375 $Y=0.34
+ $X2=3.705 $Y2=0.34
r49 12 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=0.425
+ $X2=3.54 $Y2=0.34
r50 12 14 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.54 $Y=0.425 $X2=3.54
+ $Y2=0.515
r51 11 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.845 $Y=0.34
+ $X2=2.68 $Y2=0.34
r52 10 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=0.34
+ $X2=3.54 $Y2=0.34
r53 10 11 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.375 $Y=0.34
+ $X2=2.845 $Y2=0.34
r54 3 20 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=4.4
+ $Y=0.37 $X2=4.54 $Y2=0.675
r55 2 14 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.4
+ $Y=0.37 $X2=3.54 $Y2=0.515
r56 1 25 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=2.535
+ $Y=0.37 $X2=2.68 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_MS__A32OI_2%A_771_74# 1 2 9 11 12 15
r28 13 15 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=5.49 $Y=1.01
+ $X2=5.49 $Y2=0.515
r29 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.365 $Y=1.095
+ $X2=5.49 $Y2=1.01
r30 11 12 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=5.365 $Y=1.095
+ $X2=4.205 $Y2=1.095
r31 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.04 $Y=1.01
+ $X2=4.205 $Y2=1.095
r32 7 9 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=4.04 $Y=1.01 $X2=4.04
+ $Y2=0.76
r33 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.39
+ $Y=0.37 $X2=5.53 $Y2=0.515
r34 1 9 182 $w=1.7e-07 $l=4.7355e-07 $layer=licon1_NDIFF $count=1 $X=3.855
+ $Y=0.37 $X2=4.04 $Y2=0.76
.ends


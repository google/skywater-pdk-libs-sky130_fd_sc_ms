* File: sky130_fd_sc_ms__dlymetal6s6s_1.spice
* Created: Fri Aug 28 17:31:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dlymetal6s6s_1.pex.spice"
.subckt sky130_fd_sc_ms__dlymetal6s6s_1  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_M1006_g N_A_28_138#_M1006_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0824069 AS=0.1113 PD=0.782069 PS=1.37 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_A_209_74#_M1002_d N_A_28_138#_M1002_g N_VGND_M1006_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1961 AS=0.145193 PD=2.01 PS=1.37793 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_209_74#_M1007_g N_A_316_138#_M1007_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0824069 AS=0.1113 PD=0.782069 PS=1.37 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1008 N_A_497_74#_M1008_d N_A_316_138#_M1008_g N_VGND_M1007_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1961 AS=0.145193 PD=2.01 PS=1.37793 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A_497_74#_M1001_g N_A_604_138#_M1001_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0824069 AS=0.1113 PD=0.782069 PS=1.37 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_604_138#_M1005_g N_VGND_M1001_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.145193 PD=2.01 PS=1.37793 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_28_138#_M1000_s VPB PSHORT L=0.18 W=0.42
+ AD=0.0880091 AS=0.1092 PD=0.793636 PS=1.36 NRD=72.4763 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1003 N_A_209_74#_M1003_d N_A_28_138#_M1003_g N_VPWR_M1000_d VPB PSHORT L=0.18
+ W=1.12 AD=0.2912 AS=0.234691 PD=2.76 PS=2.11636 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.4 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1004 N_VPWR_M1004_d N_A_209_74#_M1004_g N_A_316_138#_M1004_s VPB PSHORT L=0.18
+ W=0.42 AD=0.0880091 AS=0.1092 PD=0.793636 PS=1.36 NRD=72.4763 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1009 N_A_497_74#_M1009_d N_A_316_138#_M1009_g N_VPWR_M1004_d VPB PSHORT L=0.18
+ W=1.12 AD=0.2912 AS=0.234691 PD=2.76 PS=2.11636 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.4 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1010 N_VPWR_M1010_d N_A_497_74#_M1010_g N_A_604_138#_M1010_s VPB PSHORT L=0.18
+ W=0.42 AD=0.0895364 AS=0.1092 PD=0.796364 PS=1.36 NRD=74.1902 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1011 N_X_M1011_d N_A_604_138#_M1011_g N_VPWR_M1010_d VPB PSHORT L=0.18 W=1.12
+ AD=0.2912 AS=0.238764 PD=2.76 PS=2.12364 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.4
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX12_noxref VNB VPB NWDIODE A=9.6348 P=14.08
*
.include "sky130_fd_sc_ms__dlymetal6s6s_1.pxi.spice"
*
.ends
*
*

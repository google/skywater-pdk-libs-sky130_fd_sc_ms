* File: sky130_fd_sc_ms__a2bb2o_4.pxi.spice
* Created: Fri Aug 28 17:04:24 2020
* 
x_PM_SKY130_FD_SC_MS__A2BB2O_4%A_162_48# N_A_162_48#_M1017_d N_A_162_48#_M1001_s
+ N_A_162_48#_M1003_d N_A_162_48#_M1000_g N_A_162_48#_M1012_g
+ N_A_162_48#_M1007_g N_A_162_48#_M1016_g N_A_162_48#_M1010_g
+ N_A_162_48#_M1018_g N_A_162_48#_M1021_g N_A_162_48#_M1020_g
+ N_A_162_48#_c_230_p N_A_162_48#_c_146_n N_A_162_48#_c_147_n
+ N_A_162_48#_c_148_n N_A_162_48#_c_149_n N_A_162_48#_c_150_n
+ N_A_162_48#_c_151_n N_A_162_48#_c_152_n N_A_162_48#_c_153_n
+ N_A_162_48#_c_154_n N_A_162_48#_c_155_n N_A_162_48#_c_156_n
+ N_A_162_48#_c_157_n N_A_162_48#_c_158_n N_A_162_48#_c_159_n
+ PM_SKY130_FD_SC_MS__A2BB2O_4%A_162_48#
x_PM_SKY130_FD_SC_MS__A2BB2O_4%A1_N N_A1_N_M1002_g N_A1_N_M1014_g A1_N
+ N_A1_N_c_305_n N_A1_N_c_306_n PM_SKY130_FD_SC_MS__A2BB2O_4%A1_N
x_PM_SKY130_FD_SC_MS__A2BB2O_4%A2_N N_A2_N_M1006_g N_A2_N_M1022_g A2_N
+ N_A2_N_c_344_n PM_SKY130_FD_SC_MS__A2BB2O_4%A2_N
x_PM_SKY130_FD_SC_MS__A2BB2O_4%A_586_94# N_A_586_94#_M1014_d N_A_586_94#_M1006_d
+ N_A_586_94#_c_380_n N_A_586_94#_M1017_g N_A_586_94#_M1003_g
+ N_A_586_94#_c_382_n N_A_586_94#_M1004_g N_A_586_94#_c_383_n
+ N_A_586_94#_c_408_n N_A_586_94#_c_384_n N_A_586_94#_c_394_n
+ N_A_586_94#_c_395_n N_A_586_94#_c_396_n N_A_586_94#_c_385_n
+ N_A_586_94#_c_386_n N_A_586_94#_c_387_n PM_SKY130_FD_SC_MS__A2BB2O_4%A_586_94#
x_PM_SKY130_FD_SC_MS__A2BB2O_4%B2 N_B2_M1009_g N_B2_M1001_g N_B2_M1013_g
+ N_B2_M1011_g B2 B2 N_B2_c_471_n PM_SKY130_FD_SC_MS__A2BB2O_4%B2
x_PM_SKY130_FD_SC_MS__A2BB2O_4%B1 N_B1_M1015_g N_B1_M1005_g N_B1_M1019_g
+ N_B1_M1008_g B1 B1 N_B1_c_520_n PM_SKY130_FD_SC_MS__A2BB2O_4%B1
x_PM_SKY130_FD_SC_MS__A2BB2O_4%VPWR N_VPWR_M1012_s N_VPWR_M1016_s N_VPWR_M1020_s
+ N_VPWR_M1009_d N_VPWR_M1015_d N_VPWR_c_561_n N_VPWR_c_562_n N_VPWR_c_563_n
+ N_VPWR_c_564_n N_VPWR_c_565_n N_VPWR_c_566_n N_VPWR_c_567_n N_VPWR_c_568_n
+ N_VPWR_c_569_n VPWR N_VPWR_c_570_n N_VPWR_c_571_n N_VPWR_c_572_n
+ N_VPWR_c_573_n N_VPWR_c_560_n N_VPWR_c_575_n N_VPWR_c_576_n N_VPWR_c_577_n
+ PM_SKY130_FD_SC_MS__A2BB2O_4%VPWR
x_PM_SKY130_FD_SC_MS__A2BB2O_4%X N_X_M1000_s N_X_M1010_s N_X_M1012_d N_X_M1018_d
+ N_X_c_651_n N_X_c_647_n N_X_c_648_n N_X_c_653_n N_X_c_649_n N_X_c_654_n
+ N_X_c_650_n N_X_c_655_n N_X_c_656_n X X PM_SKY130_FD_SC_MS__A2BB2O_4%X
x_PM_SKY130_FD_SC_MS__A2BB2O_4%A_820_392# N_A_820_392#_M1003_s
+ N_A_820_392#_M1004_s N_A_820_392#_M1013_s N_A_820_392#_M1019_s
+ N_A_820_392#_c_718_n N_A_820_392#_c_719_n N_A_820_392#_c_720_n
+ N_A_820_392#_c_721_n N_A_820_392#_c_742_n N_A_820_392#_c_722_n
+ N_A_820_392#_c_723_n N_A_820_392#_c_724_n N_A_820_392#_c_725_n
+ N_A_820_392#_c_726_n N_A_820_392#_c_727_n
+ PM_SKY130_FD_SC_MS__A2BB2O_4%A_820_392#
x_PM_SKY130_FD_SC_MS__A2BB2O_4%VGND N_VGND_M1000_d N_VGND_M1007_d N_VGND_M1021_d
+ N_VGND_M1022_d N_VGND_M1005_s N_VGND_c_780_n N_VGND_c_781_n N_VGND_c_782_n
+ N_VGND_c_783_n N_VGND_c_784_n N_VGND_c_785_n N_VGND_c_786_n N_VGND_c_787_n
+ N_VGND_c_788_n N_VGND_c_789_n N_VGND_c_790_n N_VGND_c_791_n N_VGND_c_792_n
+ N_VGND_c_793_n VGND N_VGND_c_794_n N_VGND_c_795_n N_VGND_c_796_n
+ N_VGND_c_797_n PM_SKY130_FD_SC_MS__A2BB2O_4%VGND
x_PM_SKY130_FD_SC_MS__A2BB2O_4%A_1009_74# N_A_1009_74#_M1001_d
+ N_A_1009_74#_M1011_d N_A_1009_74#_M1008_d N_A_1009_74#_c_875_n
+ N_A_1009_74#_c_876_n N_A_1009_74#_c_877_n N_A_1009_74#_c_878_n
+ N_A_1009_74#_c_879_n PM_SKY130_FD_SC_MS__A2BB2O_4%A_1009_74#
cc_1 VNB N_A_162_48#_M1000_g 0.0237255f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.74
cc_2 VNB N_A_162_48#_M1012_g 0.00167398f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.4
cc_3 VNB N_A_162_48#_M1007_g 0.0203596f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=0.74
cc_4 VNB N_A_162_48#_M1016_g 0.00154179f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=2.4
cc_5 VNB N_A_162_48#_M1010_g 0.0209199f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=0.74
cc_6 VNB N_A_162_48#_M1018_g 0.00154258f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=2.4
cc_7 VNB N_A_162_48#_M1021_g 0.0229405f $X=-0.19 $Y=-0.245 $X2=2.175 $Y2=0.74
cc_8 VNB N_A_162_48#_M1020_g 0.00152102f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=2.4
cc_9 VNB N_A_162_48#_c_146_n 0.00750527f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.095
cc_10 VNB N_A_162_48#_c_147_n 2.98445e-19 $X=-0.19 $Y=-0.245 $X2=2.73 $Y2=1.01
cc_11 VNB N_A_162_48#_c_148_n 0.0112066f $X=-0.19 $Y=-0.245 $X2=3.36 $Y2=0.34
cc_12 VNB N_A_162_48#_c_149_n 0.00241579f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=0.34
cc_13 VNB N_A_162_48#_c_150_n 7.35049e-19 $X=-0.19 $Y=-0.245 $X2=3.445 $Y2=1.01
cc_14 VNB N_A_162_48#_c_151_n 0.0132956f $X=-0.19 $Y=-0.245 $X2=4.565 $Y2=1.095
cc_15 VNB N_A_162_48#_c_152_n 0.00142487f $X=-0.19 $Y=-0.245 $X2=3.53 $Y2=1.095
cc_16 VNB N_A_162_48#_c_153_n 0.00278408f $X=-0.19 $Y=-0.245 $X2=4.69 $Y2=0.6
cc_17 VNB N_A_162_48#_c_154_n 0.0046355f $X=-0.19 $Y=-0.245 $X2=4.69 $Y2=1.01
cc_18 VNB N_A_162_48#_c_155_n 0.01106f $X=-0.19 $Y=-0.245 $X2=4.675 $Y2=2.105
cc_19 VNB N_A_162_48#_c_156_n 0.015867f $X=-0.19 $Y=-0.245 $X2=5.6 $Y2=0.515
cc_20 VNB N_A_162_48#_c_157_n 0.00148253f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.095
cc_21 VNB N_A_162_48#_c_158_n 0.00325813f $X=-0.19 $Y=-0.245 $X2=4.69 $Y2=1.095
cc_22 VNB N_A_162_48#_c_159_n 0.0908561f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.465
cc_23 VNB N_A1_N_M1014_g 0.0250245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A1_N_c_305_n 0.0242551f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.74
cc_25 VNB N_A1_N_c_306_n 0.00408011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A2_N_M1022_g 0.0298731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB A2_N 0.00375198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A2_N_c_344_n 0.0325429f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.4
cc_29 VNB N_A_586_94#_c_380_n 0.00596955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_586_94#_M1017_g 0.0530923f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.74
cc_31 VNB N_A_586_94#_c_382_n 0.0183901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_586_94#_c_383_n 0.00116432f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=2.4
cc_33 VNB N_A_586_94#_c_384_n 0.00576653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_586_94#_c_385_n 0.00337719f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=1.63
cc_35 VNB N_A_586_94#_c_386_n 0.0217151f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=2.4
cc_36 VNB N_A_586_94#_c_387_n 0.00170689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_B2_M1009_g 0.00409125f $X=-0.19 $Y=-0.245 $X2=4.54 $Y2=1.96
cc_38 VNB N_B2_M1001_g 0.0300448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_B2_M1013_g 0.00309826f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.74
cc_40 VNB N_B2_M1011_g 0.0240386f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.4
cc_41 VNB B2 0.00542577f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=1.3
cc_42 VNB N_B2_c_471_n 0.0434519f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=0.74
cc_43 VNB N_B1_M1015_g 0.00375404f $X=-0.19 $Y=-0.245 $X2=4.54 $Y2=1.96
cc_44 VNB N_B1_M1005_g 0.0245899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_B1_M1019_g 0.00418093f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.74
cc_46 VNB N_B1_M1008_g 0.0330373f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.4
cc_47 VNB B1 0.0210179f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=1.3
cc_48 VNB N_B1_c_520_n 0.0441015f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=0.74
cc_49 VNB N_VPWR_c_560_n 0.302998f $X=-0.19 $Y=-0.245 $X2=4.69 $Y2=0.475
cc_50 VNB N_X_c_647_n 0.0596433f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.63
cc_51 VNB N_X_c_648_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_X_c_649_n 0.0046653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_X_c_650_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=2.4
cc_54 VNB N_VGND_c_780_n 0.0276293f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=1.3
cc_55 VNB N_VGND_c_781_n 0.00420208f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.63
cc_56 VNB N_VGND_c_782_n 0.00520439f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=1.3
cc_57 VNB N_VGND_c_783_n 0.0126152f $X=-0.19 $Y=-0.245 $X2=1.85 $Y2=1.63
cc_58 VNB N_VGND_c_784_n 0.0182134f $X=-0.19 $Y=-0.245 $X2=2.175 $Y2=0.74
cc_59 VNB N_VGND_c_785_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_786_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=2.4
cc_61 VNB N_VGND_c_787_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=2.3 $Y2=2.4
cc_62 VNB N_VGND_c_788_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=2.215 $Y2=1.465
cc_63 VNB N_VGND_c_789_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.465
cc_64 VNB N_VGND_c_790_n 0.00114005f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.465
cc_65 VNB N_VGND_c_791_n 0.00500927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_792_n 0.054636f $X=-0.19 $Y=-0.245 $X2=2.73 $Y2=0.425
cc_67 VNB N_VGND_c_793_n 0.00311272f $X=-0.19 $Y=-0.245 $X2=2.73 $Y2=1.01
cc_68 VNB N_VGND_c_794_n 0.0306025f $X=-0.19 $Y=-0.245 $X2=4.815 $Y2=0.475
cc_69 VNB N_VGND_c_795_n 0.0170727f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.465
cc_70 VNB N_VGND_c_796_n 0.418406f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.465
cc_71 VNB N_VGND_c_797_n 0.0129863f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=1.465
cc_72 VNB N_A_1009_74#_c_875_n 0.0162311f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=1.3
cc_73 VNB N_A_1009_74#_c_876_n 0.00178301f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.4
cc_74 VNB N_A_1009_74#_c_877_n 0.0161319f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=1.3
cc_75 VNB N_A_1009_74#_c_878_n 0.0237116f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.63
cc_76 VNB N_A_1009_74#_c_879_n 0.00159638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VPB N_A_162_48#_M1012_g 0.0253328f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.4
cc_78 VPB N_A_162_48#_M1016_g 0.0220569f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=2.4
cc_79 VPB N_A_162_48#_M1018_g 0.0220581f $X=-0.19 $Y=1.66 $X2=1.85 $Y2=2.4
cc_80 VPB N_A_162_48#_M1020_g 0.0236381f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=2.4
cc_81 VPB N_A_162_48#_c_155_n 0.00268752f $X=-0.19 $Y=1.66 $X2=4.675 $Y2=2.105
cc_82 VPB N_A1_N_M1002_g 0.021191f $X=-0.19 $Y=1.66 $X2=4.54 $Y2=1.96
cc_83 VPB N_A1_N_c_305_n 0.00552298f $X=-0.19 $Y=1.66 $X2=0.885 $Y2=0.74
cc_84 VPB N_A1_N_c_306_n 0.00303227f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A2_N_M1006_g 0.0253332f $X=-0.19 $Y=1.66 $X2=4.54 $Y2=1.96
cc_86 VPB A2_N 0.00432203f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A2_N_c_344_n 0.00966947f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.4
cc_88 VPB N_A_586_94#_c_380_n 0.00891792f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_586_94#_M1003_g 0.0236077f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.4
cc_90 VPB N_A_586_94#_c_382_n 0.0119758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_586_94#_M1004_g 0.020652f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_586_94#_c_383_n 0.00267445f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=2.4
cc_93 VPB N_A_586_94#_c_384_n 0.00125128f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_586_94#_c_394_n 0.0198168f $X=-0.19 $Y=1.66 $X2=1.85 $Y2=2.4
cc_95 VPB N_A_586_94#_c_395_n 0.0248325f $X=-0.19 $Y=1.66 $X2=2.175 $Y2=1.3
cc_96 VPB N_A_586_94#_c_396_n 6.41458e-19 $X=-0.19 $Y=1.66 $X2=2.175 $Y2=0.74
cc_97 VPB N_A_586_94#_c_385_n 0.00291884f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=1.63
cc_98 VPB N_A_586_94#_c_386_n 0.0176849f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=2.4
cc_99 VPB N_B2_M1009_g 0.0283247f $X=-0.19 $Y=1.66 $X2=4.54 $Y2=1.96
cc_100 VPB N_B2_M1013_g 0.0282176f $X=-0.19 $Y=1.66 $X2=0.885 $Y2=0.74
cc_101 VPB B2 0.00561136f $X=-0.19 $Y=1.66 $X2=1.315 $Y2=1.3
cc_102 VPB N_B1_M1015_g 0.0293486f $X=-0.19 $Y=1.66 $X2=4.54 $Y2=1.96
cc_103 VPB N_B1_M1019_g 0.0386589f $X=-0.19 $Y=1.66 $X2=0.885 $Y2=0.74
cc_104 VPB B1 0.0110874f $X=-0.19 $Y=1.66 $X2=1.315 $Y2=1.3
cc_105 VPB N_VPWR_c_561_n 0.0435224f $X=-0.19 $Y=1.66 $X2=1.315 $Y2=1.3
cc_106 VPB N_VPWR_c_562_n 0.00797179f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.63
cc_107 VPB N_VPWR_c_563_n 0.0067963f $X=-0.19 $Y=1.66 $X2=1.745 $Y2=1.3
cc_108 VPB N_VPWR_c_564_n 0.00554449f $X=-0.19 $Y=1.66 $X2=1.85 $Y2=2.4
cc_109 VPB N_VPWR_c_565_n 0.00797179f $X=-0.19 $Y=1.66 $X2=2.175 $Y2=0.74
cc_110 VPB N_VPWR_c_566_n 0.0206041f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=2.4
cc_111 VPB N_VPWR_c_567_n 0.00324402f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=2.4
cc_112 VPB N_VPWR_c_568_n 0.0206041f $X=-0.19 $Y=1.66 $X2=2.215 $Y2=1.465
cc_113 VPB N_VPWR_c_569_n 0.00324402f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.465
cc_114 VPB N_VPWR_c_570_n 0.0199636f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_571_n 0.0196495f $X=-0.19 $Y=1.66 $X2=4.565 $Y2=1.095
cc_116 VPB N_VPWR_c_572_n 0.0696198f $X=-0.19 $Y=1.66 $X2=4.662 $Y2=1.18
cc_117 VPB N_VPWR_c_573_n 0.0199471f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_560_n 0.122376f $X=-0.19 $Y=1.66 $X2=4.69 $Y2=0.475
cc_119 VPB N_VPWR_c_575_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0.885 $Y2=1.465
cc_120 VPB N_VPWR_c_576_n 0.00689679f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.465
cc_121 VPB N_VPWR_c_577_n 0.00458862f $X=-0.19 $Y=1.66 $X2=1.745 $Y2=1.465
cc_122 VPB N_X_c_651_n 2.14924e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_X_c_647_n 0.0296656f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.63
cc_124 VPB N_X_c_653_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_X_c_654_n 0.00443716f $X=-0.19 $Y=1.66 $X2=1.745 $Y2=0.74
cc_126 VPB N_X_c_655_n 0.00231613f $X=-0.19 $Y=1.66 $X2=2.175 $Y2=0.74
cc_127 VPB N_X_c_656_n 0.00224287f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=2.4
cc_128 VPB N_A_820_392#_c_718_n 0.00964539f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=2.4
cc_129 VPB N_A_820_392#_c_719_n 0.00440264f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_820_392#_c_720_n 0.00769469f $X=-0.19 $Y=1.66 $X2=1.315 $Y2=1.3
cc_131 VPB N_A_820_392#_c_721_n 0.00896004f $X=-0.19 $Y=1.66 $X2=1.315 $Y2=0.74
cc_132 VPB N_A_820_392#_c_722_n 0.00393558f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=2.4
cc_133 VPB N_A_820_392#_c_723_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.745 $Y2=0.74
cc_134 VPB N_A_820_392#_c_724_n 0.00288143f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_820_392#_c_725_n 0.010492f $X=-0.19 $Y=1.66 $X2=1.85 $Y2=2.4
cc_136 VPB N_A_820_392#_c_726_n 0.0358769f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_820_392#_c_727_n 0.0039456f $X=-0.19 $Y=1.66 $X2=2.3 $Y2=1.63
cc_138 N_A_162_48#_M1020_g N_A1_N_M1002_g 0.0241994f $X=2.3 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A_162_48#_M1021_g N_A1_N_M1014_g 0.0130514f $X=2.175 $Y=0.74 $X2=0
+ $Y2=0
cc_140 N_A_162_48#_c_146_n N_A1_N_M1014_g 0.00512257f $X=2.645 $Y=1.095 $X2=0
+ $Y2=0
cc_141 N_A_162_48#_c_147_n N_A1_N_M1014_g 0.0143856f $X=2.73 $Y=1.01 $X2=0 $Y2=0
cc_142 N_A_162_48#_c_148_n N_A1_N_M1014_g 0.00873242f $X=3.36 $Y=0.34 $X2=0
+ $Y2=0
cc_143 N_A_162_48#_c_149_n N_A1_N_M1014_g 0.00182405f $X=2.815 $Y=0.34 $X2=0
+ $Y2=0
cc_144 N_A_162_48#_c_157_n N_A1_N_M1014_g 0.00135656f $X=2.3 $Y=1.095 $X2=0
+ $Y2=0
cc_145 N_A_162_48#_c_159_n N_A1_N_M1014_g 0.00154283f $X=2.3 $Y=1.465 $X2=0
+ $Y2=0
cc_146 N_A_162_48#_c_146_n N_A1_N_c_305_n 0.0013807f $X=2.645 $Y=1.095 $X2=0
+ $Y2=0
cc_147 N_A_162_48#_c_157_n N_A1_N_c_305_n 3.19362e-19 $X=2.3 $Y=1.095 $X2=0
+ $Y2=0
cc_148 N_A_162_48#_c_159_n N_A1_N_c_305_n 0.0215078f $X=2.3 $Y=1.465 $X2=0 $Y2=0
cc_149 N_A_162_48#_c_146_n N_A1_N_c_306_n 0.0215242f $X=2.645 $Y=1.095 $X2=0
+ $Y2=0
cc_150 N_A_162_48#_c_157_n N_A1_N_c_306_n 0.0209458f $X=2.3 $Y=1.095 $X2=0 $Y2=0
cc_151 N_A_162_48#_c_159_n N_A1_N_c_306_n 0.00528487f $X=2.3 $Y=1.465 $X2=0
+ $Y2=0
cc_152 N_A_162_48#_c_147_n N_A2_N_M1022_g 6.37674e-19 $X=2.73 $Y=1.01 $X2=0
+ $Y2=0
cc_153 N_A_162_48#_c_148_n N_A2_N_M1022_g 0.0126063f $X=3.36 $Y=0.34 $X2=0 $Y2=0
cc_154 N_A_162_48#_c_150_n N_A2_N_M1022_g 0.0122699f $X=3.445 $Y=1.01 $X2=0
+ $Y2=0
cc_155 N_A_162_48#_c_152_n N_A2_N_M1022_g 0.00420304f $X=3.53 $Y=1.095 $X2=0
+ $Y2=0
cc_156 N_A_162_48#_c_151_n A2_N 0.0121728f $X=4.565 $Y=1.095 $X2=0 $Y2=0
cc_157 N_A_162_48#_c_152_n A2_N 0.0146015f $X=3.53 $Y=1.095 $X2=0 $Y2=0
cc_158 N_A_162_48#_c_151_n N_A2_N_c_344_n 0.00179145f $X=4.565 $Y=1.095 $X2=0
+ $Y2=0
cc_159 N_A_162_48#_c_152_n N_A2_N_c_344_n 0.00396026f $X=3.53 $Y=1.095 $X2=0
+ $Y2=0
cc_160 N_A_162_48#_c_151_n N_A_586_94#_c_380_n 0.00521975f $X=4.565 $Y=1.095
+ $X2=0 $Y2=0
cc_161 N_A_162_48#_c_151_n N_A_586_94#_M1017_g 0.0202752f $X=4.565 $Y=1.095
+ $X2=0 $Y2=0
cc_162 N_A_162_48#_c_153_n N_A_586_94#_M1017_g 4.60815e-19 $X=4.69 $Y=0.6 $X2=0
+ $Y2=0
cc_163 N_A_162_48#_c_155_n N_A_586_94#_M1017_g 0.0159753f $X=4.675 $Y=2.105
+ $X2=0 $Y2=0
cc_164 N_A_162_48#_c_155_n N_A_586_94#_M1003_g 0.00211741f $X=4.675 $Y=2.105
+ $X2=0 $Y2=0
cc_165 N_A_162_48#_c_155_n N_A_586_94#_c_382_n 0.0158993f $X=4.675 $Y=2.105
+ $X2=0 $Y2=0
cc_166 N_A_162_48#_c_158_n N_A_586_94#_c_382_n 0.00192341f $X=4.69 $Y=1.095
+ $X2=0 $Y2=0
cc_167 N_A_162_48#_c_155_n N_A_586_94#_M1004_g 0.00409479f $X=4.675 $Y=2.105
+ $X2=0 $Y2=0
cc_168 N_A_162_48#_c_151_n N_A_586_94#_c_383_n 0.0016349f $X=4.565 $Y=1.095
+ $X2=0 $Y2=0
cc_169 N_A_162_48#_c_148_n N_A_586_94#_c_408_n 0.0142089f $X=3.36 $Y=0.34 $X2=0
+ $Y2=0
cc_170 N_A_162_48#_c_146_n N_A_586_94#_c_384_n 0.00331391f $X=2.645 $Y=1.095
+ $X2=0 $Y2=0
cc_171 N_A_162_48#_c_157_n N_A_586_94#_c_384_n 0.00488541f $X=2.3 $Y=1.095 $X2=0
+ $Y2=0
cc_172 N_A_162_48#_c_155_n N_A_586_94#_c_395_n 0.00414326f $X=4.675 $Y=2.105
+ $X2=0 $Y2=0
cc_173 N_A_162_48#_c_151_n N_A_586_94#_c_385_n 0.0156104f $X=4.565 $Y=1.095
+ $X2=0 $Y2=0
cc_174 N_A_162_48#_c_155_n N_A_586_94#_c_385_n 0.0185329f $X=4.675 $Y=2.105
+ $X2=0 $Y2=0
cc_175 N_A_162_48#_c_151_n N_A_586_94#_c_386_n 0.00303502f $X=4.565 $Y=1.095
+ $X2=0 $Y2=0
cc_176 N_A_162_48#_c_146_n N_A_586_94#_c_387_n 0.00545578f $X=2.645 $Y=1.095
+ $X2=0 $Y2=0
cc_177 N_A_162_48#_c_152_n N_A_586_94#_c_387_n 0.00975088f $X=3.53 $Y=1.095
+ $X2=0 $Y2=0
cc_178 N_A_162_48#_c_155_n N_B2_M1009_g 4.20847e-19 $X=4.675 $Y=2.105 $X2=0
+ $Y2=0
cc_179 N_A_162_48#_c_154_n N_B2_M1001_g 0.00307188f $X=4.69 $Y=1.01 $X2=0 $Y2=0
cc_180 N_A_162_48#_c_155_n N_B2_M1001_g 0.00184906f $X=4.675 $Y=2.105 $X2=0
+ $Y2=0
cc_181 N_A_162_48#_c_156_n N_B2_M1001_g 0.0132302f $X=5.6 $Y=0.515 $X2=0 $Y2=0
cc_182 N_A_162_48#_c_158_n N_B2_M1001_g 0.0029913f $X=4.69 $Y=1.095 $X2=0 $Y2=0
cc_183 N_A_162_48#_c_156_n N_B2_M1011_g 0.00337267f $X=5.6 $Y=0.515 $X2=0 $Y2=0
cc_184 N_A_162_48#_c_155_n B2 0.0145622f $X=4.675 $Y=2.105 $X2=0 $Y2=0
cc_185 N_A_162_48#_c_155_n N_B2_c_471_n 0.00779214f $X=4.675 $Y=2.105 $X2=0
+ $Y2=0
cc_186 N_A_162_48#_M1012_g N_VPWR_c_561_n 0.00742848f $X=0.95 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A_162_48#_M1016_g N_VPWR_c_562_n 0.00329146f $X=1.4 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A_162_48#_M1018_g N_VPWR_c_562_n 0.00329146f $X=1.85 $Y=2.4 $X2=0 $Y2=0
cc_189 N_A_162_48#_M1020_g N_VPWR_c_563_n 0.00940768f $X=2.3 $Y=2.4 $X2=0 $Y2=0
cc_190 N_A_162_48#_M1012_g N_VPWR_c_566_n 0.005209f $X=0.95 $Y=2.4 $X2=0 $Y2=0
cc_191 N_A_162_48#_M1016_g N_VPWR_c_566_n 0.005209f $X=1.4 $Y=2.4 $X2=0 $Y2=0
cc_192 N_A_162_48#_M1018_g N_VPWR_c_571_n 0.005209f $X=1.85 $Y=2.4 $X2=0 $Y2=0
cc_193 N_A_162_48#_M1020_g N_VPWR_c_571_n 0.005209f $X=2.3 $Y=2.4 $X2=0 $Y2=0
cc_194 N_A_162_48#_M1012_g N_VPWR_c_560_n 0.00987399f $X=0.95 $Y=2.4 $X2=0 $Y2=0
cc_195 N_A_162_48#_M1016_g N_VPWR_c_560_n 0.00982266f $X=1.4 $Y=2.4 $X2=0 $Y2=0
cc_196 N_A_162_48#_M1018_g N_VPWR_c_560_n 0.00982266f $X=1.85 $Y=2.4 $X2=0 $Y2=0
cc_197 N_A_162_48#_M1020_g N_VPWR_c_560_n 0.00982496f $X=2.3 $Y=2.4 $X2=0 $Y2=0
cc_198 N_A_162_48#_M1012_g N_X_c_651_n 0.0162518f $X=0.95 $Y=2.4 $X2=0 $Y2=0
cc_199 N_A_162_48#_c_159_n N_X_c_651_n 7.7481e-19 $X=2.3 $Y=1.465 $X2=0 $Y2=0
cc_200 N_A_162_48#_M1000_g N_X_c_647_n 0.0223647f $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A_162_48#_M1012_g N_X_c_647_n 0.00589889f $X=0.95 $Y=2.4 $X2=0 $Y2=0
cc_202 N_A_162_48#_M1007_g N_X_c_647_n 5.75161e-19 $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A_162_48#_c_230_p N_X_c_647_n 0.0370738f $X=2.215 $Y=1.465 $X2=0 $Y2=0
cc_204 N_A_162_48#_c_159_n N_X_c_647_n 0.0169446f $X=2.3 $Y=1.465 $X2=0 $Y2=0
cc_205 N_A_162_48#_M1000_g N_X_c_648_n 0.0128625f $X=0.885 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A_162_48#_M1007_g N_X_c_648_n 3.97481e-19 $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A_162_48#_M1012_g N_X_c_653_n 0.019068f $X=0.95 $Y=2.4 $X2=0 $Y2=0
cc_208 N_A_162_48#_M1016_g N_X_c_653_n 0.0143027f $X=1.4 $Y=2.4 $X2=0 $Y2=0
cc_209 N_A_162_48#_M1018_g N_X_c_653_n 6.97946e-19 $X=1.85 $Y=2.4 $X2=0 $Y2=0
cc_210 N_A_162_48#_M1007_g N_X_c_649_n 0.0124434f $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A_162_48#_M1010_g N_X_c_649_n 0.0120709f $X=1.745 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A_162_48#_c_230_p N_X_c_649_n 0.0657213f $X=2.215 $Y=1.465 $X2=0 $Y2=0
cc_213 N_A_162_48#_c_157_n N_X_c_649_n 0.00497192f $X=2.3 $Y=1.095 $X2=0 $Y2=0
cc_214 N_A_162_48#_c_159_n N_X_c_649_n 0.00536003f $X=2.3 $Y=1.465 $X2=0 $Y2=0
cc_215 N_A_162_48#_M1016_g N_X_c_654_n 0.012931f $X=1.4 $Y=2.4 $X2=0 $Y2=0
cc_216 N_A_162_48#_M1018_g N_X_c_654_n 0.0142852f $X=1.85 $Y=2.4 $X2=0 $Y2=0
cc_217 N_A_162_48#_M1020_g N_X_c_654_n 0.00441435f $X=2.3 $Y=2.4 $X2=0 $Y2=0
cc_218 N_A_162_48#_c_230_p N_X_c_654_n 0.0672186f $X=2.215 $Y=1.465 $X2=0 $Y2=0
cc_219 N_A_162_48#_c_157_n N_X_c_654_n 0.00201744f $X=2.3 $Y=1.095 $X2=0 $Y2=0
cc_220 N_A_162_48#_c_159_n N_X_c_654_n 0.00482403f $X=2.3 $Y=1.465 $X2=0 $Y2=0
cc_221 N_A_162_48#_M1007_g N_X_c_650_n 6.20738e-19 $X=1.315 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A_162_48#_M1010_g N_X_c_650_n 0.00866629f $X=1.745 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A_162_48#_M1021_g N_X_c_650_n 3.97481e-19 $X=2.175 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A_162_48#_M1016_g N_X_c_655_n 6.97946e-19 $X=1.4 $Y=2.4 $X2=0 $Y2=0
cc_225 N_A_162_48#_M1018_g N_X_c_655_n 0.0143027f $X=1.85 $Y=2.4 $X2=0 $Y2=0
cc_226 N_A_162_48#_M1020_g N_X_c_655_n 0.0125234f $X=2.3 $Y=2.4 $X2=0 $Y2=0
cc_227 N_A_162_48#_M1012_g N_X_c_656_n 0.00170136f $X=0.95 $Y=2.4 $X2=0 $Y2=0
cc_228 N_A_162_48#_M1016_g N_X_c_656_n 0.00134521f $X=1.4 $Y=2.4 $X2=0 $Y2=0
cc_229 N_A_162_48#_c_230_p N_X_c_656_n 0.0255674f $X=2.215 $Y=1.465 $X2=0 $Y2=0
cc_230 N_A_162_48#_c_159_n N_X_c_656_n 0.0023727f $X=2.3 $Y=1.465 $X2=0 $Y2=0
cc_231 N_A_162_48#_M1003_d N_A_820_392#_c_719_n 0.00165831f $X=4.54 $Y=1.96
+ $X2=0 $Y2=0
cc_232 N_A_162_48#_c_155_n N_A_820_392#_c_719_n 0.0118736f $X=4.675 $Y=2.105
+ $X2=0 $Y2=0
cc_233 N_A_162_48#_c_155_n N_A_820_392#_c_721_n 0.00659243f $X=4.675 $Y=2.105
+ $X2=0 $Y2=0
cc_234 N_A_162_48#_c_146_n N_VGND_M1021_d 0.00860096f $X=2.645 $Y=1.095 $X2=0
+ $Y2=0
cc_235 N_A_162_48#_c_147_n N_VGND_M1021_d 0.00604133f $X=2.73 $Y=1.01 $X2=0
+ $Y2=0
cc_236 N_A_162_48#_c_157_n N_VGND_M1021_d 0.0011083f $X=2.3 $Y=1.095 $X2=0 $Y2=0
cc_237 N_A_162_48#_c_150_n N_VGND_M1022_d 0.0129017f $X=3.445 $Y=1.01 $X2=0
+ $Y2=0
cc_238 N_A_162_48#_c_151_n N_VGND_M1022_d 0.0164421f $X=4.565 $Y=1.095 $X2=0
+ $Y2=0
cc_239 N_A_162_48#_c_152_n N_VGND_M1022_d 6.25458e-19 $X=3.53 $Y=1.095 $X2=0
+ $Y2=0
cc_240 N_A_162_48#_M1000_g N_VGND_c_780_n 0.00466772f $X=0.885 $Y=0.74 $X2=0
+ $Y2=0
cc_241 N_A_162_48#_M1000_g N_VGND_c_781_n 5.05592e-19 $X=0.885 $Y=0.74 $X2=0
+ $Y2=0
cc_242 N_A_162_48#_M1007_g N_VGND_c_781_n 0.00914496f $X=1.315 $Y=0.74 $X2=0
+ $Y2=0
cc_243 N_A_162_48#_M1010_g N_VGND_c_781_n 0.00183835f $X=1.745 $Y=0.74 $X2=0
+ $Y2=0
cc_244 N_A_162_48#_M1010_g N_VGND_c_782_n 5.20618e-19 $X=1.745 $Y=0.74 $X2=0
+ $Y2=0
cc_245 N_A_162_48#_M1021_g N_VGND_c_782_n 0.0117339f $X=2.175 $Y=0.74 $X2=0
+ $Y2=0
cc_246 N_A_162_48#_c_146_n N_VGND_c_782_n 0.00724091f $X=2.645 $Y=1.095 $X2=0
+ $Y2=0
cc_247 N_A_162_48#_c_147_n N_VGND_c_782_n 0.0310611f $X=2.73 $Y=1.01 $X2=0 $Y2=0
cc_248 N_A_162_48#_c_149_n N_VGND_c_782_n 0.0146659f $X=2.815 $Y=0.34 $X2=0
+ $Y2=0
cc_249 N_A_162_48#_c_157_n N_VGND_c_782_n 0.00887034f $X=2.3 $Y=1.095 $X2=0
+ $Y2=0
cc_250 N_A_162_48#_c_159_n N_VGND_c_782_n 5.02668e-19 $X=2.3 $Y=1.465 $X2=0
+ $Y2=0
cc_251 N_A_162_48#_c_148_n N_VGND_c_783_n 0.0158668f $X=3.36 $Y=0.34 $X2=0 $Y2=0
cc_252 N_A_162_48#_c_150_n N_VGND_c_783_n 0.0337298f $X=3.445 $Y=1.01 $X2=0
+ $Y2=0
cc_253 N_A_162_48#_c_151_n N_VGND_c_783_n 0.0507639f $X=4.565 $Y=1.095 $X2=0
+ $Y2=0
cc_254 N_A_162_48#_c_153_n N_VGND_c_783_n 0.0109137f $X=4.69 $Y=0.6 $X2=0 $Y2=0
cc_255 N_A_162_48#_M1000_g N_VGND_c_786_n 0.00434272f $X=0.885 $Y=0.74 $X2=0
+ $Y2=0
cc_256 N_A_162_48#_M1007_g N_VGND_c_786_n 0.00383152f $X=1.315 $Y=0.74 $X2=0
+ $Y2=0
cc_257 N_A_162_48#_M1010_g N_VGND_c_788_n 0.00434272f $X=1.745 $Y=0.74 $X2=0
+ $Y2=0
cc_258 N_A_162_48#_M1021_g N_VGND_c_788_n 0.00383152f $X=2.175 $Y=0.74 $X2=0
+ $Y2=0
cc_259 N_A_162_48#_c_153_n N_VGND_c_792_n 0.0111552f $X=4.69 $Y=0.6 $X2=0 $Y2=0
cc_260 N_A_162_48#_c_156_n N_VGND_c_792_n 0.0388592f $X=5.6 $Y=0.515 $X2=0 $Y2=0
cc_261 N_A_162_48#_c_148_n N_VGND_c_794_n 0.0472364f $X=3.36 $Y=0.34 $X2=0 $Y2=0
cc_262 N_A_162_48#_c_149_n N_VGND_c_794_n 0.0121867f $X=2.815 $Y=0.34 $X2=0
+ $Y2=0
cc_263 N_A_162_48#_M1000_g N_VGND_c_796_n 0.00825283f $X=0.885 $Y=0.74 $X2=0
+ $Y2=0
cc_264 N_A_162_48#_M1007_g N_VGND_c_796_n 0.0075754f $X=1.315 $Y=0.74 $X2=0
+ $Y2=0
cc_265 N_A_162_48#_M1010_g N_VGND_c_796_n 0.00820284f $X=1.745 $Y=0.74 $X2=0
+ $Y2=0
cc_266 N_A_162_48#_M1021_g N_VGND_c_796_n 0.0075754f $X=2.175 $Y=0.74 $X2=0
+ $Y2=0
cc_267 N_A_162_48#_c_148_n N_VGND_c_796_n 0.027092f $X=3.36 $Y=0.34 $X2=0 $Y2=0
cc_268 N_A_162_48#_c_149_n N_VGND_c_796_n 0.00660921f $X=2.815 $Y=0.34 $X2=0
+ $Y2=0
cc_269 N_A_162_48#_c_153_n N_VGND_c_796_n 0.00923333f $X=4.69 $Y=0.6 $X2=0 $Y2=0
cc_270 N_A_162_48#_c_156_n N_VGND_c_796_n 0.033121f $X=5.6 $Y=0.515 $X2=0 $Y2=0
cc_271 N_A_162_48#_c_156_n N_A_1009_74#_M1001_d 0.00332037f $X=5.6 $Y=0.515
+ $X2=-0.19 $Y2=-0.245
cc_272 N_A_162_48#_M1001_s N_A_1009_74#_c_875_n 0.00176801f $X=5.46 $Y=0.37
+ $X2=0 $Y2=0
cc_273 N_A_162_48#_c_154_n N_A_1009_74#_c_875_n 0.0191245f $X=4.69 $Y=1.01 $X2=0
+ $Y2=0
cc_274 N_A_162_48#_c_156_n N_A_1009_74#_c_875_n 0.0438027f $X=5.6 $Y=0.515 $X2=0
+ $Y2=0
cc_275 N_A_162_48#_c_158_n N_A_1009_74#_c_875_n 0.00683847f $X=4.69 $Y=1.095
+ $X2=0 $Y2=0
cc_276 N_A_162_48#_c_156_n N_A_1009_74#_c_876_n 0.010629f $X=5.6 $Y=0.515 $X2=0
+ $Y2=0
cc_277 N_A1_N_M1002_g N_A2_N_M1006_g 0.0519612f $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_278 N_A1_N_M1014_g N_A2_N_M1022_g 0.0234549f $X=2.855 $Y=0.79 $X2=0 $Y2=0
cc_279 N_A1_N_c_305_n N_A2_N_c_344_n 0.0519612f $X=2.765 $Y=1.515 $X2=0 $Y2=0
cc_280 N_A1_N_c_306_n N_A2_N_c_344_n 3.74559e-19 $X=2.765 $Y=1.515 $X2=0 $Y2=0
cc_281 N_A1_N_M1014_g N_A_586_94#_c_384_n 0.00872368f $X=2.855 $Y=0.79 $X2=0
+ $Y2=0
cc_282 N_A1_N_c_306_n N_A_586_94#_c_384_n 0.0320025f $X=2.765 $Y=1.515 $X2=0
+ $Y2=0
cc_283 N_A1_N_M1002_g N_A_586_94#_c_394_n 0.00234609f $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_284 N_A1_N_M1002_g N_A_586_94#_c_396_n 0.00135549f $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_285 N_A1_N_M1014_g N_A_586_94#_c_387_n 6.65078e-19 $X=2.855 $Y=0.79 $X2=0
+ $Y2=0
cc_286 N_A1_N_M1002_g N_VPWR_c_563_n 0.0221989f $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_287 N_A1_N_c_305_n N_VPWR_c_563_n 7.80375e-19 $X=2.765 $Y=1.515 $X2=0 $Y2=0
cc_288 N_A1_N_c_306_n N_VPWR_c_563_n 0.0169894f $X=2.765 $Y=1.515 $X2=0 $Y2=0
cc_289 N_A1_N_M1002_g N_VPWR_c_572_n 0.00460063f $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_290 N_A1_N_M1002_g N_VPWR_c_560_n 0.00908061f $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_291 N_A1_N_M1002_g N_X_c_654_n 6.13915e-19 $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_292 N_A1_N_M1002_g N_X_c_655_n 2.26923e-19 $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_293 N_A1_N_M1014_g N_VGND_c_782_n 0.00145351f $X=2.855 $Y=0.79 $X2=0 $Y2=0
cc_294 N_A1_N_M1014_g N_VGND_c_794_n 7.822e-19 $X=2.855 $Y=0.79 $X2=0 $Y2=0
cc_295 A2_N N_A_586_94#_M1017_g 0.00262375f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_296 N_A2_N_M1006_g N_A_586_94#_c_384_n 0.00694339f $X=3.23 $Y=2.4 $X2=0 $Y2=0
cc_297 A2_N N_A_586_94#_c_384_n 0.0310564f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_298 N_A2_N_c_344_n N_A_586_94#_c_384_n 0.00876725f $X=3.445 $Y=1.515 $X2=0
+ $Y2=0
cc_299 N_A2_N_M1006_g N_A_586_94#_c_394_n 0.016131f $X=3.23 $Y=2.4 $X2=0 $Y2=0
cc_300 N_A2_N_M1006_g N_A_586_94#_c_396_n 0.016288f $X=3.23 $Y=2.4 $X2=0 $Y2=0
cc_301 A2_N N_A_586_94#_c_396_n 0.0253713f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_302 N_A2_N_c_344_n N_A_586_94#_c_396_n 0.00133254f $X=3.445 $Y=1.515 $X2=0
+ $Y2=0
cc_303 N_A2_N_M1006_g N_A_586_94#_c_385_n 0.00218401f $X=3.23 $Y=2.4 $X2=0 $Y2=0
cc_304 A2_N N_A_586_94#_c_385_n 0.0243455f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_305 N_A2_N_c_344_n N_A_586_94#_c_385_n 2.11902e-19 $X=3.445 $Y=1.515 $X2=0
+ $Y2=0
cc_306 N_A2_N_M1006_g N_A_586_94#_c_386_n 0.00212665f $X=3.23 $Y=2.4 $X2=0 $Y2=0
cc_307 A2_N N_A_586_94#_c_386_n 0.00238956f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_308 N_A2_N_c_344_n N_A_586_94#_c_386_n 0.0131988f $X=3.445 $Y=1.515 $X2=0
+ $Y2=0
cc_309 N_A2_N_M1022_g N_A_586_94#_c_387_n 0.00532649f $X=3.285 $Y=0.79 $X2=0
+ $Y2=0
cc_310 N_A2_N_M1006_g N_VPWR_c_563_n 0.00303692f $X=3.23 $Y=2.4 $X2=0 $Y2=0
cc_311 N_A2_N_M1006_g N_VPWR_c_572_n 0.005209f $X=3.23 $Y=2.4 $X2=0 $Y2=0
cc_312 N_A2_N_M1006_g N_VPWR_c_560_n 0.00988003f $X=3.23 $Y=2.4 $X2=0 $Y2=0
cc_313 N_A2_N_M1022_g N_VGND_c_783_n 4.48089e-19 $X=3.285 $Y=0.79 $X2=0 $Y2=0
cc_314 N_A2_N_M1022_g N_VGND_c_794_n 7.82463e-19 $X=3.285 $Y=0.79 $X2=0 $Y2=0
cc_315 N_A_586_94#_c_382_n N_B2_M1009_g 0.0211214f $X=4.81 $Y=1.725 $X2=0 $Y2=0
cc_316 N_A_586_94#_c_382_n B2 4.93152e-19 $X=4.81 $Y=1.725 $X2=0 $Y2=0
cc_317 N_A_586_94#_c_394_n N_VPWR_c_563_n 0.0265385f $X=3.455 $Y=2.815 $X2=0
+ $Y2=0
cc_318 N_A_586_94#_c_396_n N_VPWR_c_563_n 0.0107238f $X=3.62 $Y=2.035 $X2=0
+ $Y2=0
cc_319 N_A_586_94#_M1004_g N_VPWR_c_564_n 3.82437e-19 $X=4.9 $Y=2.46 $X2=0 $Y2=0
cc_320 N_A_586_94#_M1003_g N_VPWR_c_572_n 0.00333896f $X=4.45 $Y=2.46 $X2=0
+ $Y2=0
cc_321 N_A_586_94#_M1004_g N_VPWR_c_572_n 0.00333896f $X=4.9 $Y=2.46 $X2=0 $Y2=0
cc_322 N_A_586_94#_c_394_n N_VPWR_c_572_n 0.014549f $X=3.455 $Y=2.815 $X2=0
+ $Y2=0
cc_323 N_A_586_94#_M1003_g N_VPWR_c_560_n 0.00427818f $X=4.45 $Y=2.46 $X2=0
+ $Y2=0
cc_324 N_A_586_94#_M1004_g N_VPWR_c_560_n 0.00422796f $X=4.9 $Y=2.46 $X2=0 $Y2=0
cc_325 N_A_586_94#_c_394_n N_VPWR_c_560_n 0.0119743f $X=3.455 $Y=2.815 $X2=0
+ $Y2=0
cc_326 N_A_586_94#_c_384_n A_586_368# 0.0014055f $X=3.105 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_327 N_A_586_94#_c_396_n A_586_368# 0.00419084f $X=3.62 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_328 N_A_586_94#_c_395_n N_A_820_392#_M1003_s 0.00299216f $X=3.855 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_329 N_A_586_94#_M1003_g N_A_820_392#_c_718_n 0.00971842f $X=4.45 $Y=2.46
+ $X2=0 $Y2=0
cc_330 N_A_586_94#_M1004_g N_A_820_392#_c_718_n 5.56591e-19 $X=4.9 $Y=2.46 $X2=0
+ $Y2=0
cc_331 N_A_586_94#_c_394_n N_A_820_392#_c_718_n 0.0265266f $X=3.455 $Y=2.815
+ $X2=0 $Y2=0
cc_332 N_A_586_94#_c_395_n N_A_820_392#_c_718_n 0.00813517f $X=3.855 $Y=2.035
+ $X2=0 $Y2=0
cc_333 N_A_586_94#_c_386_n N_A_820_392#_c_718_n 0.00552791f $X=3.985 $Y=1.635
+ $X2=0 $Y2=0
cc_334 N_A_586_94#_M1003_g N_A_820_392#_c_719_n 0.0115958f $X=4.45 $Y=2.46 $X2=0
+ $Y2=0
cc_335 N_A_586_94#_M1004_g N_A_820_392#_c_719_n 0.0132535f $X=4.9 $Y=2.46 $X2=0
+ $Y2=0
cc_336 N_A_586_94#_M1003_g N_A_820_392#_c_720_n 0.00291744f $X=4.45 $Y=2.46
+ $X2=0 $Y2=0
cc_337 N_A_586_94#_c_394_n N_A_820_392#_c_720_n 0.00343054f $X=3.455 $Y=2.815
+ $X2=0 $Y2=0
cc_338 N_A_586_94#_M1004_g N_A_820_392#_c_721_n 0.00353824f $X=4.9 $Y=2.46 $X2=0
+ $Y2=0
cc_339 N_A_586_94#_M1003_g N_A_820_392#_c_742_n 6.28799e-19 $X=4.45 $Y=2.46
+ $X2=0 $Y2=0
cc_340 N_A_586_94#_M1004_g N_A_820_392#_c_742_n 0.0105282f $X=4.9 $Y=2.46 $X2=0
+ $Y2=0
cc_341 N_A_586_94#_M1017_g N_VGND_c_783_n 0.016897f $X=4.435 $Y=0.74 $X2=0 $Y2=0
cc_342 N_A_586_94#_M1017_g N_VGND_c_792_n 0.00383152f $X=4.435 $Y=0.74 $X2=0
+ $Y2=0
cc_343 N_A_586_94#_M1017_g N_VGND_c_796_n 0.00762539f $X=4.435 $Y=0.74 $X2=0
+ $Y2=0
cc_344 N_B2_M1013_g N_B1_M1015_g 0.0195547f $X=5.8 $Y=2.46 $X2=0 $Y2=0
cc_345 N_B2_M1011_g N_B1_M1005_g 0.0181154f $X=5.815 $Y=0.69 $X2=0 $Y2=0
cc_346 B2 B1 0.0356352f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_347 N_B2_c_471_n B1 2.24997e-19 $X=5.815 $Y=1.425 $X2=0 $Y2=0
cc_348 B2 N_B1_c_520_n 0.00559665f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_349 N_B2_c_471_n N_B1_c_520_n 0.0195547f $X=5.815 $Y=1.425 $X2=0 $Y2=0
cc_350 N_B2_M1009_g N_VPWR_c_564_n 0.011752f $X=5.35 $Y=2.46 $X2=0 $Y2=0
cc_351 N_B2_M1013_g N_VPWR_c_564_n 0.002979f $X=5.8 $Y=2.46 $X2=0 $Y2=0
cc_352 N_B2_M1013_g N_VPWR_c_568_n 0.005209f $X=5.8 $Y=2.46 $X2=0 $Y2=0
cc_353 N_B2_M1009_g N_VPWR_c_572_n 0.00460063f $X=5.35 $Y=2.46 $X2=0 $Y2=0
cc_354 N_B2_M1009_g N_VPWR_c_560_n 0.00908665f $X=5.35 $Y=2.46 $X2=0 $Y2=0
cc_355 N_B2_M1013_g N_VPWR_c_560_n 0.00982376f $X=5.8 $Y=2.46 $X2=0 $Y2=0
cc_356 N_B2_M1009_g N_A_820_392#_c_719_n 0.00101073f $X=5.35 $Y=2.46 $X2=0 $Y2=0
cc_357 N_B2_M1009_g N_A_820_392#_c_722_n 0.01879f $X=5.35 $Y=2.46 $X2=0 $Y2=0
cc_358 N_B2_M1013_g N_A_820_392#_c_722_n 0.012931f $X=5.8 $Y=2.46 $X2=0 $Y2=0
cc_359 B2 N_A_820_392#_c_722_n 0.0358836f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_360 N_B2_c_471_n N_A_820_392#_c_722_n 4.03951e-19 $X=5.815 $Y=1.425 $X2=0
+ $Y2=0
cc_361 N_B2_M1009_g N_A_820_392#_c_723_n 6.74232e-19 $X=5.35 $Y=2.46 $X2=0 $Y2=0
cc_362 N_B2_M1013_g N_A_820_392#_c_723_n 0.0121322f $X=5.8 $Y=2.46 $X2=0 $Y2=0
cc_363 N_B2_M1013_g N_A_820_392#_c_727_n 0.00100213f $X=5.8 $Y=2.46 $X2=0 $Y2=0
cc_364 B2 N_A_820_392#_c_727_n 0.0230491f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_365 N_B2_M1001_g N_VGND_c_792_n 0.00291649f $X=5.385 $Y=0.69 $X2=0 $Y2=0
cc_366 N_B2_M1011_g N_VGND_c_792_n 0.00433162f $X=5.815 $Y=0.69 $X2=0 $Y2=0
cc_367 N_B2_M1001_g N_VGND_c_796_n 0.0036412f $X=5.385 $Y=0.69 $X2=0 $Y2=0
cc_368 N_B2_M1011_g N_VGND_c_796_n 0.00432528f $X=5.815 $Y=0.69 $X2=0 $Y2=0
cc_369 N_B2_M1001_g N_A_1009_74#_c_875_n 0.017183f $X=5.385 $Y=0.69 $X2=0 $Y2=0
cc_370 N_B2_M1011_g N_A_1009_74#_c_875_n 0.0144965f $X=5.815 $Y=0.69 $X2=0 $Y2=0
cc_371 B2 N_A_1009_74#_c_875_n 0.0434573f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_372 N_B2_c_471_n N_A_1009_74#_c_875_n 0.00460578f $X=5.815 $Y=1.425 $X2=0
+ $Y2=0
cc_373 B2 N_A_1009_74#_c_879_n 0.015544f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_374 N_B1_M1015_g N_VPWR_c_565_n 0.0027763f $X=6.25 $Y=2.46 $X2=0 $Y2=0
cc_375 N_B1_M1019_g N_VPWR_c_565_n 0.0027763f $X=6.7 $Y=2.46 $X2=0 $Y2=0
cc_376 N_B1_M1015_g N_VPWR_c_568_n 0.005209f $X=6.25 $Y=2.46 $X2=0 $Y2=0
cc_377 N_B1_M1019_g N_VPWR_c_573_n 0.005209f $X=6.7 $Y=2.46 $X2=0 $Y2=0
cc_378 N_B1_M1015_g N_VPWR_c_560_n 0.00982376f $X=6.25 $Y=2.46 $X2=0 $Y2=0
cc_379 N_B1_M1019_g N_VPWR_c_560_n 0.0098599f $X=6.7 $Y=2.46 $X2=0 $Y2=0
cc_380 N_B1_M1015_g N_A_820_392#_c_723_n 0.0119338f $X=6.25 $Y=2.46 $X2=0 $Y2=0
cc_381 N_B1_M1019_g N_A_820_392#_c_723_n 6.50516e-19 $X=6.7 $Y=2.46 $X2=0 $Y2=0
cc_382 N_B1_M1015_g N_A_820_392#_c_724_n 0.0174816f $X=6.25 $Y=2.46 $X2=0 $Y2=0
cc_383 N_B1_M1019_g N_A_820_392#_c_724_n 0.012931f $X=6.7 $Y=2.46 $X2=0 $Y2=0
cc_384 B1 N_A_820_392#_c_724_n 0.0312334f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_385 N_B1_c_520_n N_A_820_392#_c_724_n 4.05102e-19 $X=6.715 $Y=1.425 $X2=0
+ $Y2=0
cc_386 N_B1_M1019_g N_A_820_392#_c_725_n 0.00108119f $X=6.7 $Y=2.46 $X2=0 $Y2=0
cc_387 B1 N_A_820_392#_c_725_n 0.0285352f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_388 N_B1_M1015_g N_A_820_392#_c_726_n 6.50516e-19 $X=6.25 $Y=2.46 $X2=0 $Y2=0
cc_389 N_B1_M1019_g N_A_820_392#_c_726_n 0.0121004f $X=6.7 $Y=2.46 $X2=0 $Y2=0
cc_390 N_B1_M1015_g N_A_820_392#_c_727_n 0.00212471f $X=6.25 $Y=2.46 $X2=0 $Y2=0
cc_391 N_B1_M1005_g N_VGND_c_790_n 0.00502457f $X=6.245 $Y=0.69 $X2=0 $Y2=0
cc_392 N_B1_M1008_g N_VGND_c_790_n 0.00503476f $X=6.715 $Y=0.69 $X2=0 $Y2=0
cc_393 N_B1_M1005_g N_VGND_c_791_n 0.00226696f $X=6.245 $Y=0.69 $X2=0 $Y2=0
cc_394 N_B1_M1008_g N_VGND_c_791_n 0.00568798f $X=6.715 $Y=0.69 $X2=0 $Y2=0
cc_395 N_B1_M1005_g N_VGND_c_792_n 0.00434272f $X=6.245 $Y=0.69 $X2=0 $Y2=0
cc_396 N_B1_M1008_g N_VGND_c_795_n 0.00383152f $X=6.715 $Y=0.69 $X2=0 $Y2=0
cc_397 N_B1_M1005_g N_VGND_c_796_n 0.00821754f $X=6.245 $Y=0.69 $X2=0 $Y2=0
cc_398 N_B1_M1008_g N_VGND_c_796_n 0.00761163f $X=6.715 $Y=0.69 $X2=0 $Y2=0
cc_399 N_B1_M1005_g N_A_1009_74#_c_877_n 0.0180055f $X=6.245 $Y=0.69 $X2=0 $Y2=0
cc_400 N_B1_M1008_g N_A_1009_74#_c_877_n 0.0140902f $X=6.715 $Y=0.69 $X2=0 $Y2=0
cc_401 B1 N_A_1009_74#_c_877_n 0.0580465f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_402 N_B1_c_520_n N_A_1009_74#_c_877_n 0.00375093f $X=6.715 $Y=1.425 $X2=0
+ $Y2=0
cc_403 N_B1_M1008_g N_A_1009_74#_c_878_n 4.43891e-19 $X=6.715 $Y=0.69 $X2=0
+ $Y2=0
cc_404 N_VPWR_M1012_s N_X_c_647_n 0.00749944f $X=0.6 $Y=1.84 $X2=0 $Y2=0
cc_405 N_VPWR_c_561_n N_X_c_647_n 0.0180926f $X=0.725 $Y=2.305 $X2=0 $Y2=0
cc_406 N_VPWR_c_561_n N_X_c_653_n 0.0283501f $X=0.725 $Y=2.305 $X2=0 $Y2=0
cc_407 N_VPWR_c_562_n N_X_c_653_n 0.0283117f $X=1.625 $Y=2.305 $X2=0 $Y2=0
cc_408 N_VPWR_c_566_n N_X_c_653_n 0.0144623f $X=1.54 $Y=3.33 $X2=0 $Y2=0
cc_409 N_VPWR_c_560_n N_X_c_653_n 0.0118344f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_410 N_VPWR_M1016_s N_X_c_654_n 0.00165831f $X=1.49 $Y=1.84 $X2=0 $Y2=0
cc_411 N_VPWR_c_562_n N_X_c_654_n 0.0126919f $X=1.625 $Y=2.305 $X2=0 $Y2=0
cc_412 N_VPWR_c_562_n N_X_c_655_n 0.0283117f $X=1.625 $Y=2.305 $X2=0 $Y2=0
cc_413 N_VPWR_c_563_n N_X_c_655_n 0.0386643f $X=2.595 $Y=2.115 $X2=0 $Y2=0
cc_414 N_VPWR_c_571_n N_X_c_655_n 0.0144623f $X=2.41 $Y=3.33 $X2=0 $Y2=0
cc_415 N_VPWR_c_560_n N_X_c_655_n 0.0118344f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_416 N_VPWR_c_564_n N_A_820_392#_c_719_n 0.010126f $X=5.575 $Y=2.455 $X2=0
+ $Y2=0
cc_417 N_VPWR_c_572_n N_A_820_392#_c_719_n 0.0536089f $X=5.41 $Y=3.33 $X2=0
+ $Y2=0
cc_418 N_VPWR_c_560_n N_A_820_392#_c_719_n 0.0296408f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_419 N_VPWR_c_572_n N_A_820_392#_c_720_n 0.0235512f $X=5.41 $Y=3.33 $X2=0
+ $Y2=0
cc_420 N_VPWR_c_560_n N_A_820_392#_c_720_n 0.0126924f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_421 N_VPWR_M1009_d N_A_820_392#_c_722_n 0.00165831f $X=5.44 $Y=1.96 $X2=0
+ $Y2=0
cc_422 N_VPWR_c_564_n N_A_820_392#_c_722_n 0.0148589f $X=5.575 $Y=2.455 $X2=0
+ $Y2=0
cc_423 N_VPWR_c_564_n N_A_820_392#_c_723_n 0.0234083f $X=5.575 $Y=2.455 $X2=0
+ $Y2=0
cc_424 N_VPWR_c_565_n N_A_820_392#_c_723_n 0.0233699f $X=6.475 $Y=2.455 $X2=0
+ $Y2=0
cc_425 N_VPWR_c_568_n N_A_820_392#_c_723_n 0.0144623f $X=6.39 $Y=3.33 $X2=0
+ $Y2=0
cc_426 N_VPWR_c_560_n N_A_820_392#_c_723_n 0.0118344f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_427 N_VPWR_M1015_d N_A_820_392#_c_724_n 0.00165831f $X=6.34 $Y=1.96 $X2=0
+ $Y2=0
cc_428 N_VPWR_c_565_n N_A_820_392#_c_724_n 0.0126919f $X=6.475 $Y=2.455 $X2=0
+ $Y2=0
cc_429 N_VPWR_c_565_n N_A_820_392#_c_726_n 0.0233699f $X=6.475 $Y=2.455 $X2=0
+ $Y2=0
cc_430 N_VPWR_c_573_n N_A_820_392#_c_726_n 0.014549f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_431 N_VPWR_c_560_n N_A_820_392#_c_726_n 0.0119743f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_432 N_X_c_647_n N_VGND_M1000_d 0.00300749f $X=0.835 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_433 N_X_c_649_n N_VGND_M1007_d 0.00176461f $X=1.795 $Y=1.045 $X2=0 $Y2=0
cc_434 N_X_c_647_n N_VGND_c_780_n 0.0224079f $X=0.835 $Y=1.885 $X2=0 $Y2=0
cc_435 N_X_c_648_n N_VGND_c_780_n 0.0158413f $X=1.1 $Y=0.515 $X2=0 $Y2=0
cc_436 N_X_c_648_n N_VGND_c_781_n 0.0158413f $X=1.1 $Y=0.515 $X2=0 $Y2=0
cc_437 N_X_c_649_n N_VGND_c_781_n 0.0152916f $X=1.795 $Y=1.045 $X2=0 $Y2=0
cc_438 N_X_c_650_n N_VGND_c_781_n 0.0158413f $X=1.96 $Y=0.515 $X2=0 $Y2=0
cc_439 N_X_c_650_n N_VGND_c_782_n 0.0175587f $X=1.96 $Y=0.515 $X2=0 $Y2=0
cc_440 N_X_c_648_n N_VGND_c_786_n 0.0109942f $X=1.1 $Y=0.515 $X2=0 $Y2=0
cc_441 N_X_c_650_n N_VGND_c_788_n 0.0109942f $X=1.96 $Y=0.515 $X2=0 $Y2=0
cc_442 N_X_c_648_n N_VGND_c_796_n 0.00904371f $X=1.1 $Y=0.515 $X2=0 $Y2=0
cc_443 N_X_c_650_n N_VGND_c_796_n 0.00904371f $X=1.96 $Y=0.515 $X2=0 $Y2=0
cc_444 N_VGND_c_796_n N_A_1009_74#_c_875_n 0.00730683f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_445 N_VGND_c_790_n N_A_1009_74#_c_876_n 0.0152763f $X=6.48 $Y=0.55 $X2=0
+ $Y2=0
cc_446 N_VGND_c_792_n N_A_1009_74#_c_876_n 0.00749631f $X=6.495 $Y=0 $X2=0 $Y2=0
cc_447 N_VGND_c_796_n N_A_1009_74#_c_876_n 0.0062048f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_448 N_VGND_M1005_s N_A_1009_74#_c_877_n 0.00218982f $X=6.32 $Y=0.37 $X2=0
+ $Y2=0
cc_449 N_VGND_c_790_n N_A_1009_74#_c_877_n 0.019937f $X=6.48 $Y=0.55 $X2=0 $Y2=0
cc_450 N_VGND_c_790_n N_A_1009_74#_c_878_n 0.0153177f $X=6.48 $Y=0.55 $X2=0
+ $Y2=0
cc_451 N_VGND_c_795_n N_A_1009_74#_c_878_n 0.011066f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_452 N_VGND_c_796_n N_A_1009_74#_c_878_n 0.00915947f $X=6.96 $Y=0 $X2=0 $Y2=0

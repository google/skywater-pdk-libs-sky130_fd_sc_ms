* File: sky130_fd_sc_ms__mux2_1.spice
* Created: Fri Aug 28 17:39:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__mux2_1.pex.spice"
.subckt sky130_fd_sc_ms__mux2_1  VNB VPB S A1 A0 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A0	A0
* A1	A1
* S	S
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_S_M1006_g N_A_27_112#_M1006_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.123281 AS=0.15675 PD=0.98062 PS=1.67 NRD=13.632 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75003.5 A=0.0825 P=1.4 MULT=1
MM1008 A_226_74# N_S_M1008_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.165869 PD=0.98 PS=1.31938 NRD=10.536 NRS=11.34 M=1 R=4.93333 SA=75000.6
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1007 N_A_304_74#_M1007_d N_A1_M1007_g A_226_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.20165 AS=0.0888 PD=1.285 PS=0.98 NRD=21.072 NRS=10.536 M=1 R=4.93333
+ SA=75001 SB=75002.6 A=0.111 P=1.78 MULT=1
MM1002 A_443_74# N_A0_M1002_g N_A_304_74#_M1007_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2997 AS=0.20165 PD=1.55 PS=1.285 NRD=56.748 NRS=21.888 M=1 R=4.93333
+ SA=75001.7 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_27_112#_M1009_g A_443_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.20905 AS=0.2997 PD=1.305 PS=1.55 NRD=23.508 NRS=56.748 M=1 R=4.93333
+ SA=75002.7 SB=75000.9 A=0.111 P=1.78 MULT=1
MM1010 N_X_M1010_d N_A_304_74#_M1010_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.20905 PD=2.05 PS=1.305 NRD=0 NRS=22.692 M=1 R=4.93333
+ SA=75003.4 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_VPWR_M1003_d N_S_M1003_g N_A_27_112#_M1003_s VPB PSHORT L=0.18 W=0.84
+ AD=0.156587 AS=0.2352 PD=1.23717 PS=2.24 NRD=18.7544 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90003.4 A=0.1512 P=2.04 MULT=1
MM1011 A_226_368# N_S_M1011_g N_VPWR_M1003_d VPB PSHORT L=0.18 W=1 AD=0.3925
+ AS=0.186413 PD=1.785 PS=1.47283 NRD=66.4678 NRS=0 M=1 R=5.55556 SA=90000.6
+ SB=90002.9 A=0.18 P=2.36 MULT=1
MM1000 N_A_304_74#_M1000_d N_A0_M1000_g A_226_368# VPB PSHORT L=0.18 W=1 AD=0.18
+ AS=0.3925 PD=1.36 PS=1.785 NRD=0 NRS=66.4678 M=1 R=5.55556 SA=90001.6
+ SB=90001.9 A=0.18 P=2.36 MULT=1
MM1005 A_527_368# N_A1_M1005_g N_A_304_74#_M1000_d VPB PSHORT L=0.18 W=1
+ AD=0.195 AS=0.18 PD=1.39 PS=1.36 NRD=27.5603 NRS=16.7253 M=1 R=5.55556
+ SA=90002.1 SB=90001.4 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_A_27_112#_M1004_g A_527_368# VPB PSHORT L=0.18 W=1
+ AD=0.226226 AS=0.195 PD=1.4717 PS=1.39 NRD=22.9702 NRS=27.5603 M=1 R=5.55556
+ SA=90002.7 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1001 N_X_M1001_d N_A_304_74#_M1001_g N_VPWR_M1004_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.253374 PD=2.8 PS=1.6483 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__mux2_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__dlrbp_1.pex.spice
* Created: Fri Aug 28 17:27:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLRBP_1%D 3 7 9 12
r35 12 15 40.7727 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.615
+ $X2=0.59 $Y2=1.78
r36 12 14 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.615
+ $X2=0.59 $Y2=1.45
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.615 $X2=0.6 $Y2=1.615
r38 9 13 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.72 $Y=1.615 $X2=0.6
+ $Y2=1.615
r39 7 14 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.495 $Y=0.985
+ $X2=0.495 $Y2=1.45
r40 3 15 244.887 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=0.505 $Y=2.41
+ $X2=0.505 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_1%GATE 3 7 9 12
r38 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.615
+ $X2=1.14 $Y2=1.78
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.615
+ $X2=1.14 $Y2=1.45
r40 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=1.615 $X2=1.14 $Y2=1.615
r41 7 15 244.887 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=1.125 $Y=2.41
+ $X2=1.125 $Y2=1.78
r42 3 14 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.055 $Y=0.89
+ $X2=1.055 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_1%A_226_104# 1 2 7 11 15 17 19 20 21 25 26 27
+ 28 29 36 37 39 41 42 46 48 50 56
c148 41 0 6.32864e-20 $X=3.74 $Y=0.345
c149 21 0 2.87737e-19 $X=3.225 $Y=1.765
c150 20 0 5.71781e-20 $X=3.725 $Y=1.765
r151 49 56 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.71 $Y=1.585
+ $X2=1.71 $Y2=1.495
r152 48 51 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.675 $Y=1.585
+ $X2=1.675 $Y2=1.75
r153 48 50 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.675 $Y=1.585
+ $X2=1.675 $Y2=1.42
r154 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.585 $X2=1.71 $Y2=1.585
r155 46 50 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.56 $Y=1.28
+ $X2=1.56 $Y2=1.42
r156 42 62 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.74 $Y=0.345
+ $X2=3.74 $Y2=0.51
r157 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.74
+ $Y=0.345 $X2=3.74 $Y2=0.345
r158 39 54 18.4631 $w=1.68e-07 $l=2.83e-07 $layer=LI1_cond $X=2.905 $Y=0.382
+ $X2=2.905 $Y2=0.665
r159 39 41 33.8954 $w=2.53e-07 $l=7.5e-07 $layer=LI1_cond $X=2.99 $Y=0.382
+ $X2=3.74 $Y2=0.382
r160 38 45 6.07722 $w=1.7e-07 $l=2.49199e-07 $layer=LI1_cond $X=1.645 $Y=0.665
+ $X2=1.415 $Y2=0.625
r161 37 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.82 $Y=0.665
+ $X2=2.905 $Y2=0.665
r162 37 38 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=2.82 $Y=0.665
+ $X2=1.645 $Y2=0.665
r163 36 51 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.56 $Y=1.97
+ $X2=1.56 $Y2=1.75
r164 29 36 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.475 $Y=2.095
+ $X2=1.56 $Y2=1.97
r165 29 31 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.475 $Y=2.095
+ $X2=1.385 $Y2=2.095
r166 28 46 10.9702 $w=4.58e-07 $l=2.3e-07 $layer=LI1_cond $X=1.415 $Y=1.05
+ $X2=1.415 $Y2=1.28
r167 27 45 2.81353 $w=4.6e-07 $l=1.25e-07 $layer=LI1_cond $X=1.415 $Y=0.75
+ $X2=1.415 $Y2=0.625
r168 27 28 7.80051 $w=4.58e-07 $l=3e-07 $layer=LI1_cond $X=1.415 $Y=0.75
+ $X2=1.415 $Y2=1.05
r169 25 62 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.8 $Y=0.83 $X2=3.8
+ $Y2=0.51
r170 23 25 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=3.8 $Y=1.69 $X2=3.8
+ $Y2=0.83
r171 20 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.725 $Y=1.765
+ $X2=3.8 $Y2=1.69
r172 20 21 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.725 $Y=1.765
+ $X2=3.225 $Y2=1.765
r173 17 21 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.135 $Y=1.84
+ $X2=3.225 $Y2=1.765
r174 17 19 166.022 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=3.135 $Y=1.84
+ $X2=3.135 $Y2=2.46
r175 13 26 18.8402 $w=1.65e-07 $l=2.81425e-07 $layer=POLY_cond $X=2.205 $Y=1.66
+ $X2=2.115 $Y2=1.42
r176 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.205 $Y=1.66
+ $X2=2.205 $Y2=2.38
r177 9 26 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=2.19 $Y=1.42
+ $X2=2.115 $Y2=1.42
r178 9 11 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.19 $Y=1.42
+ $X2=2.19 $Y2=0.86
r179 8 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.875 $Y=1.495
+ $X2=1.71 $Y2=1.495
r180 7 26 6.66866 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.115 $Y=1.495
+ $X2=2.115 $Y2=1.42
r181 7 8 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.115 $Y=1.495
+ $X2=1.875 $Y2=1.495
r182 2 31 600 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=1.215
+ $Y=1.99 $X2=1.385 $Y2=2.135
r183 1 45 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=1.13
+ $Y=0.52 $X2=1.35 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_1%A_27_142# 1 2 9 15 16 17 18 24 25 26 28 29
+ 31 32 34 35 39
c92 34 0 1.36773e-19 $X=2.67 $Y=1.635
c93 28 0 2.09267e-19 $X=2.59 $Y=2.39
c94 17 0 1.91696e-19 $X=2.77 $Y=1.265
c95 9 0 1.32022e-19 $X=2.745 $Y=2.46
r96 35 40 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.635
+ $X2=2.67 $Y2=1.8
r97 35 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.635
+ $X2=2.67 $Y2=1.47
r98 34 37 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.67 $Y=1.635
+ $X2=2.67 $Y2=1.8
r99 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.635 $X2=2.67 $Y2=1.635
r100 31 32 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.27 $Y=2.135
+ $X2=0.27 $Y2=1.97
r101 29 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.18 $Y=1.28
+ $X2=0.18 $Y2=1.97
r102 28 37 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.59 $Y=2.39
+ $X2=2.59 $Y2=1.8
r103 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.505 $Y=2.475
+ $X2=2.59 $Y2=2.39
r104 25 26 134.396 $w=1.68e-07 $l=2.06e-06 $layer=LI1_cond $X=2.505 $Y=2.475
+ $X2=0.445 $Y2=2.475
r105 24 26 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=0.27 $Y=2.39
+ $X2=0.445 $Y2=2.475
r106 23 31 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=0.27 $Y=2.145
+ $X2=0.27 $Y2=2.135
r107 23 24 8.0671 $w=3.48e-07 $l=2.45e-07 $layer=LI1_cond $X=0.27 $Y=2.145
+ $X2=0.27 $Y2=2.39
r108 18 29 8.81775 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=0.27 $Y=1.105
+ $X2=0.27 $Y2=1.28
r109 18 20 4.18286 $w=3.5e-07 $l=1.2e-07 $layer=LI1_cond $X=0.27 $Y=1.105
+ $X2=0.27 $Y2=0.985
r110 17 39 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.76 $Y=1.265
+ $X2=2.76 $Y2=1.47
r111 16 17 63.4211 $w=1.7e-07 $l=1.5e-07 $layer=POLY_cond $X=2.77 $Y=1.115
+ $X2=2.77 $Y2=1.265
r112 15 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.78 $Y=0.72
+ $X2=2.78 $Y2=1.115
r113 9 40 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.745 $Y=2.46
+ $X2=2.745 $Y2=1.8
r114 2 31 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.99 $X2=0.28 $Y2=2.135
r115 1 20 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.71 $X2=0.28 $Y2=0.985
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_1%A_353_98# 1 2 9 12 15 16 17 19 21 22 23 26
+ 27 32 39 41 45 48
c123 45 0 1.54446e-19 $X=3.23 $Y=1.315
c124 41 0 1.6995e-19 $X=3.2 $Y=1.215
c125 17 0 7.89243e-20 $X=2.215 $Y=1.215
c126 15 0 1.32022e-19 $X=2.13 $Y=1.94
r127 45 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.23 $Y=1.315
+ $X2=3.23 $Y2=1.15
r128 44 46 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=3.2 $Y=1.315
+ $X2=3.2 $Y2=1.48
r129 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.23
+ $Y=1.315 $X2=3.23 $Y2=1.315
r130 41 44 2.95498 $w=3.88e-07 $l=1e-07 $layer=LI1_cond $X=3.2 $Y=1.215 $X2=3.2
+ $Y2=1.315
r131 37 39 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.94 $Y=2.055
+ $X2=3.09 $Y2=2.055
r132 35 36 6.60399 $w=3.51e-07 $l=1.9e-07 $layer=LI1_cond $X=1.94 $Y=1.11
+ $X2=2.13 $Y2=1.11
r133 30 32 6.1738 $w=2.78e-07 $l=1.5e-07 $layer=LI1_cond $X=1.98 $Y=2.08
+ $X2=2.13 $Y2=2.08
r134 27 50 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=3.85 $Y=2.215
+ $X2=3.69 $Y2=2.215
r135 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.85
+ $Y=2.215 $X2=3.85 $Y2=2.215
r136 24 26 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=3.85 $Y=2.905
+ $X2=3.85 $Y2=2.215
r137 22 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.685 $Y=2.99
+ $X2=3.85 $Y2=2.905
r138 22 23 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=3.685 $Y=2.99
+ $X2=3.025 $Y2=2.99
r139 21 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.09 $Y=1.97
+ $X2=3.09 $Y2=2.055
r140 21 46 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.09 $Y=1.97
+ $X2=3.09 $Y2=1.48
r141 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.94 $Y=2.905
+ $X2=3.025 $Y2=2.99
r142 18 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.94 $Y=2.14
+ $X2=2.94 $Y2=2.055
r143 18 19 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.94 $Y=2.14
+ $X2=2.94 $Y2=2.905
r144 17 36 6.20757 $w=3.51e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.215 $Y=1.215
+ $X2=2.13 $Y2=1.11
r145 16 41 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=3.005 $Y=1.215
+ $X2=3.2 $Y2=1.215
r146 16 17 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=3.005 $Y=1.215
+ $X2=2.215 $Y2=1.215
r147 15 32 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.13 $Y=1.94
+ $X2=2.13 $Y2=2.08
r148 14 36 4.99104 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.13 $Y=1.3 $X2=2.13
+ $Y2=1.11
r149 14 15 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.13 $Y=1.3 $X2=2.13
+ $Y2=1.94
r150 10 50 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.69 $Y=2.38
+ $X2=3.69 $Y2=2.215
r151 10 12 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=3.69 $Y=2.38
+ $X2=3.69 $Y2=2.75
r152 9 48 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.14 $Y=0.72
+ $X2=3.14 $Y2=1.15
r153 2 30 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=1.835
+ $Y=1.96 $X2=1.98 $Y2=2.12
r154 1 35 182 $w=1.7e-07 $l=6.76868e-07 $layer=licon1_NDIFF $count=1 $X=1.765
+ $Y=0.49 $X2=1.94 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_1%A_823_98# 1 2 7 9 14 18 22 24 28 34 37 39 40
+ 41 42 45 49 55 57 61 64 65 66 72 74
c156 66 0 4.3223e-20 $X=5.332 $Y=1.72
c157 57 0 7.12526e-20 $X=6.005 $Y=1.805
c158 42 0 1.06492e-20 $X=5.085 $Y=2.155
c159 7 0 6.32864e-20 $X=4.19 $Y=1.115
r160 74 75 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.17 $Y=1.425
+ $X2=6.17 $Y2=1.35
r161 65 68 4.34938 $w=4.93e-07 $l=1.8e-07 $layer=LI1_cond $X=5.332 $Y=1.805
+ $X2=5.332 $Y2=1.985
r162 65 66 7.55351 $w=4.93e-07 $l=8.5e-08 $layer=LI1_cond $X=5.332 $Y=1.805
+ $X2=5.332 $Y2=1.72
r163 64 66 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.17 $Y=1.13
+ $X2=5.17 $Y2=1.72
r164 62 77 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.17 $Y=1.515
+ $X2=6.17 $Y2=1.68
r165 62 74 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.17 $Y=1.515
+ $X2=6.17 $Y2=1.425
r166 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.17
+ $Y=1.515 $X2=6.17 $Y2=1.515
r167 59 61 7.26926 $w=3.23e-07 $l=2.05e-07 $layer=LI1_cond $X=6.167 $Y=1.72
+ $X2=6.167 $Y2=1.515
r168 58 65 7.09362 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=5.58 $Y=1.805
+ $X2=5.332 $Y2=1.805
r169 57 59 7.72402 $w=1.7e-07 $l=2.00035e-07 $layer=LI1_cond $X=6.005 $Y=1.805
+ $X2=6.167 $Y2=1.72
r170 57 58 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=6.005 $Y=1.805
+ $X2=5.58 $Y2=1.805
r171 55 70 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=5.415 $Y=2.815
+ $X2=5.415 $Y2=2.32
r172 47 64 10.8817 $w=4.53e-07 $l=2.27e-07 $layer=LI1_cond $X=5.027 $Y=0.903
+ $X2=5.027 $Y2=1.13
r173 47 49 10.1995 $w=4.53e-07 $l=3.88e-07 $layer=LI1_cond $X=5.027 $Y=0.903
+ $X2=5.027 $Y2=0.515
r174 45 73 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.39 $Y=2.155
+ $X2=4.39 $Y2=2.32
r175 45 72 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.39 $Y=2.155
+ $X2=4.39 $Y2=1.99
r176 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.39
+ $Y=2.155 $X2=4.39 $Y2=2.155
r177 42 70 5.31902 $w=4.93e-07 $l=1.65e-07 $layer=LI1_cond $X=5.332 $Y=2.155
+ $X2=5.332 $Y2=2.32
r178 42 68 4.10774 $w=4.93e-07 $l=1.7e-07 $layer=LI1_cond $X=5.332 $Y=2.155
+ $X2=5.332 $Y2=1.985
r179 42 44 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.085 $Y=2.155
+ $X2=4.39 $Y2=2.155
r180 40 41 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=7.117 $Y=1.89
+ $X2=7.117 $Y2=2.04
r181 35 37 56.4043 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=4.19 $Y=1.19
+ $X2=4.3 $Y2=1.19
r182 34 41 133.889 $w=1.8e-07 $l=5e-07 $layer=POLY_cond $X=7.15 $Y=2.54 $X2=7.15
+ $Y2=2.04
r183 30 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.07 $Y=1.5
+ $X2=7.07 $Y2=1.425
r184 30 40 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=7.07 $Y=1.5
+ $X2=7.07 $Y2=1.89
r185 26 39 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.07 $Y=1.35
+ $X2=7.07 $Y2=1.425
r186 26 28 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=7.07 $Y=1.35
+ $X2=7.07 $Y2=0.645
r187 25 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.335 $Y=1.425
+ $X2=6.17 $Y2=1.425
r188 24 39 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.995 $Y=1.425
+ $X2=7.07 $Y2=1.425
r189 24 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.995 $Y=1.425
+ $X2=6.335 $Y2=1.425
r190 22 77 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.14 $Y=2.4
+ $X2=6.14 $Y2=1.68
r191 18 75 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.08 $Y=0.74
+ $X2=6.08 $Y2=1.35
r192 14 73 167.145 $w=1.8e-07 $l=4.3e-07 $layer=POLY_cond $X=4.345 $Y=2.75
+ $X2=4.345 $Y2=2.32
r193 10 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.3 $Y=1.265
+ $X2=4.3 $Y2=1.19
r194 10 72 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=4.3 $Y=1.265
+ $X2=4.3 $Y2=1.99
r195 7 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.19 $Y=1.115
+ $X2=4.19 $Y2=1.19
r196 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.19 $Y=1.115 $X2=4.19
+ $Y2=0.83
r197 2 68 400 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=5.255
+ $Y=1.84 $X2=5.415 $Y2=1.985
r198 2 55 400 $w=1.7e-07 $l=1.05196e-06 $layer=licon1_PDIFF $count=1 $X=5.255
+ $Y=1.84 $X2=5.415 $Y2=2.815
r199 1 49 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.82
+ $Y=0.37 $X2=4.965 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_1%A_643_80# 1 2 9 13 15 16 17 24 25 26 28 29
+ 35
c88 29 0 4.70832e-20 $X=3.355 $Y=2.405
c89 26 0 1.43227e-19 $X=3.75 $Y=1.735
c90 9 0 7.12526e-20 $X=5.165 $Y=2.4
r91 35 38 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=4.75 $Y=1.515
+ $X2=4.75 $Y2=1.735
r92 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.75
+ $Y=1.515 $X2=4.75 $Y2=1.515
r93 31 33 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.43 $Y=1.735
+ $X2=3.665 $Y2=1.735
r94 28 29 8.46025 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.355 $Y=2.57
+ $X2=3.355 $Y2=2.405
r95 26 33 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.75 $Y=1.735
+ $X2=3.665 $Y2=1.735
r96 25 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.585 $Y=1.735
+ $X2=4.75 $Y2=1.735
r97 25 26 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=4.585 $Y=1.735
+ $X2=3.75 $Y2=1.735
r98 24 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.665 $Y=1.65
+ $X2=3.665 $Y2=1.735
r99 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.665 $Y=0.96
+ $X2=3.665 $Y2=1.65
r100 21 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=1.82
+ $X2=3.43 $Y2=1.735
r101 21 29 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.43 $Y=1.82
+ $X2=3.43 $Y2=2.405
r102 17 23 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.58 $Y=0.835
+ $X2=3.665 $Y2=0.96
r103 17 19 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=3.58 $Y=0.835
+ $X2=3.47 $Y2=0.835
r104 15 36 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=5.075 $Y=1.515
+ $X2=4.75 $Y2=1.515
r105 15 16 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.075 $Y=1.515
+ $X2=5.165 $Y2=1.515
r106 11 16 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=5.18 $Y=1.35
+ $X2=5.165 $Y2=1.515
r107 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.18 $Y=1.35
+ $X2=5.18 $Y2=0.74
r108 7 16 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=5.165 $Y=1.68
+ $X2=5.165 $Y2=1.515
r109 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.165 $Y=1.68
+ $X2=5.165 $Y2=2.4
r110 2 28 600 $w=1.7e-07 $l=6.78638e-07 $layer=licon1_PDIFF $count=1 $X=3.225
+ $Y=1.96 $X2=3.37 $Y2=2.57
r111 1 19 182 $w=1.7e-07 $l=5.88855e-07 $layer=licon1_NDIFF $count=1 $X=3.215
+ $Y=0.4 $X2=3.47 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_1%RESET_B 3 6 8 11 12 13
c38 13 0 2.2426e-19 $X=5.63 $Y=1.22
c39 6 0 1.06492e-20 $X=5.64 $Y=2.4
r40 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.63 $Y=1.385
+ $X2=5.63 $Y2=1.55
r41 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.63 $Y=1.385
+ $X2=5.63 $Y2=1.22
r42 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.63
+ $Y=1.385 $X2=5.63 $Y2=1.385
r43 8 12 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=5.52 $Y=1.365
+ $X2=5.63 $Y2=1.365
r44 6 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=5.64 $Y=2.4 $X2=5.64
+ $Y2=1.55
r45 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.57 $Y=0.74 $X2=5.57
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_1%A_1342_74# 1 2 9 13 16 19 23 24 27 30
c58 19 0 6.46507e-20 $X=6.925 $Y=2.265
r59 27 29 9.87261 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=6.855 $Y=0.625
+ $X2=6.855 $Y2=0.84
r60 24 33 40.8642 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=7.565 $Y=1.485
+ $X2=7.565 $Y2=1.65
r61 24 32 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=7.565 $Y=1.485
+ $X2=7.565 $Y2=1.32
r62 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.55
+ $Y=1.485 $X2=7.55 $Y2=1.485
r63 21 30 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=7.02 $Y=1.485 $X2=6.93
+ $Y2=1.485
r64 21 23 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=7.02 $Y=1.485
+ $X2=7.55 $Y2=1.485
r65 17 30 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=6.925 $Y=1.65
+ $X2=6.93 $Y2=1.485
r66 17 19 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=6.925 $Y=1.65
+ $X2=6.925 $Y2=2.265
r67 16 30 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=6.93 $Y=1.32
+ $X2=6.93 $Y2=1.485
r68 16 29 29.5758 $w=1.78e-07 $l=4.8e-07 $layer=LI1_cond $X=6.93 $Y=1.32
+ $X2=6.93 $Y2=0.84
r69 13 33 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=7.655 $Y=2.4
+ $X2=7.655 $Y2=1.65
r70 9 32 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.58 $Y=0.74 $X2=7.58
+ $Y2=1.32
r71 2 19 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=6.78
+ $Y=2.12 $X2=6.925 $Y2=2.265
r72 1 27 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=6.71
+ $Y=0.37 $X2=6.855 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_1%VPWR 1 2 3 4 5 20 24 28 32 34 36 44 49 54 61
+ 62 65 68 71 78 81
r89 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r90 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r91 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r92 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r93 62 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r94 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r95 59 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.54 $Y=3.33
+ $X2=7.375 $Y2=3.33
r96 59 61 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=7.54 $Y=3.33
+ $X2=7.92 $Y2=3.33
r97 58 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r98 58 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33 $X2=6
+ $Y2=3.33
r99 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r100 55 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.03 $Y=3.33
+ $X2=5.905 $Y2=3.33
r101 55 57 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=6.03 $Y=3.33
+ $X2=6.96 $Y2=3.33
r102 54 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.21 $Y=3.33
+ $X2=7.375 $Y2=3.33
r103 54 57 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=7.21 $Y=3.33
+ $X2=6.96 $Y2=3.33
r104 53 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r105 53 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r106 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r107 50 52 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.08 $Y=3.33
+ $X2=5.52 $Y2=3.33
r108 49 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.78 $Y=3.33
+ $X2=5.905 $Y2=3.33
r109 49 52 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.78 $Y=3.33
+ $X2=5.52 $Y2=3.33
r110 45 68 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.685 $Y=3.33
+ $X2=2.517 $Y2=3.33
r111 45 47 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=2.685 $Y=3.33
+ $X2=4.08 $Y2=3.33
r112 44 50 9.08255 $w=1.7e-07 $l=3.38e-07 $layer=LI1_cond $X=4.742 $Y=3.33
+ $X2=5.08 $Y2=3.33
r113 44 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r114 44 71 9.12564 $w=6.73e-07 $l=5.15e-07 $layer=LI1_cond $X=4.742 $Y=3.33
+ $X2=4.742 $Y2=2.815
r115 44 47 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.405 $Y=3.33
+ $X2=4.08 $Y2=3.33
r116 43 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r117 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r118 40 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r119 40 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r120 39 42 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r121 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r122 37 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r123 37 39 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=1.2 $Y2=3.33
r124 36 68 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=2.35 $Y=3.33
+ $X2=2.517 $Y2=3.33
r125 36 42 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.35 $Y=3.33
+ $X2=2.16 $Y2=3.33
r126 34 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r127 34 69 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r128 34 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r129 30 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.375 $Y=3.245
+ $X2=7.375 $Y2=3.33
r130 30 32 34.2241 $w=3.28e-07 $l=9.8e-07 $layer=LI1_cond $X=7.375 $Y=3.245
+ $X2=7.375 $Y2=2.265
r131 26 78 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.905 $Y=3.245
+ $X2=5.905 $Y2=3.33
r132 26 28 47.0197 $w=2.48e-07 $l=1.02e-06 $layer=LI1_cond $X=5.905 $Y=3.245
+ $X2=5.905 $Y2=2.225
r133 22 68 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.517 $Y=3.245
+ $X2=2.517 $Y2=3.33
r134 22 24 14.7926 $w=3.33e-07 $l=4.3e-07 $layer=LI1_cond $X=2.517 $Y=3.245
+ $X2=2.517 $Y2=2.815
r135 18 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r136 18 20 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.895
r137 5 32 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=7.24
+ $Y=2.12 $X2=7.375 $Y2=2.265
r138 4 28 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=5.73
+ $Y=1.84 $X2=5.865 $Y2=2.225
r139 3 71 300 $w=1.7e-07 $l=6.01997e-07 $layer=licon1_PDIFF $count=2 $X=4.435
+ $Y=2.54 $X2=4.915 $Y2=2.815
r140 2 24 600 $w=1.7e-07 $l=9.5871e-07 $layer=licon1_PDIFF $count=1 $X=2.295
+ $Y=1.96 $X2=2.515 $Y2=2.815
r141 1 20 600 $w=1.7e-07 $l=1.00902e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.99 $X2=0.815 $Y2=2.895
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_1%Q 1 2 9 15 19 20 21 22
c40 9 0 1.81037e-19 $X=6.295 $Y=0.515
r41 21 22 9.41594 $w=4.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.435 $Y=2.405
+ $X2=6.435 $Y2=2.775
r42 19 20 9.33757 $w=4.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.435 $Y=2.225
+ $X2=6.435 $Y2=2.06
r43 17 21 2.79933 $w=4.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.435 $Y=2.295
+ $X2=6.435 $Y2=2.405
r44 17 19 1.78139 $w=4.68e-07 $l=7e-08 $layer=LI1_cond $X=6.435 $Y=2.295
+ $X2=6.435 $Y2=2.225
r45 11 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.585 $Y=1.18
+ $X2=6.585 $Y2=1.095
r46 11 20 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=6.585 $Y=1.18
+ $X2=6.585 $Y2=2.06
r47 7 15 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.295 $Y=1.095
+ $X2=6.585 $Y2=1.095
r48 7 9 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=6.295 $Y=1.01
+ $X2=6.295 $Y2=0.515
r49 2 19 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=6.23
+ $Y=1.84 $X2=6.365 $Y2=2.225
r50 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.155
+ $Y=0.37 $X2=6.295 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_1%Q_N 1 2 9 14 15 16 17 28
r22 21 28 1.90404 $w=3.43e-07 $l=5.7e-08 $layer=LI1_cond $X=7.882 $Y=0.868
+ $X2=7.882 $Y2=0.925
r23 17 30 6.34154 $w=3.43e-07 $l=1.01e-07 $layer=LI1_cond $X=7.882 $Y=0.939
+ $X2=7.882 $Y2=1.04
r24 17 28 0.467658 $w=3.43e-07 $l=1.4e-08 $layer=LI1_cond $X=7.882 $Y=0.939
+ $X2=7.882 $Y2=0.925
r25 17 21 0.467658 $w=3.43e-07 $l=1.4e-08 $layer=LI1_cond $X=7.882 $Y=0.854
+ $X2=7.882 $Y2=0.868
r26 16 17 11.324 $w=3.43e-07 $l=3.39e-07 $layer=LI1_cond $X=7.882 $Y=0.515
+ $X2=7.882 $Y2=0.854
r27 15 30 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=7.97 $Y=1.82
+ $X2=7.97 $Y2=1.04
r28 14 15 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=7.885 $Y=1.985
+ $X2=7.885 $Y2=1.82
r29 7 14 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=7.885 $Y=1.99
+ $X2=7.885 $Y2=1.985
r30 7 9 27.9637 $w=3.38e-07 $l=8.25e-07 $layer=LI1_cond $X=7.885 $Y=1.99
+ $X2=7.885 $Y2=2.815
r31 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.745
+ $Y=1.84 $X2=7.88 $Y2=1.985
r32 2 9 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.745
+ $Y=1.84 $X2=7.88 $Y2=2.815
r33 1 16 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=7.655
+ $Y=0.37 $X2=7.875 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBP_1%VGND 1 2 3 4 5 18 24 28 32 37 38 39 41 46 54
+ 63 72 73 76 80 86 89
r94 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r95 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r96 80 83 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.485 $Y=0
+ $X2=2.485 $Y2=0.325
r97 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r98 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r99 73 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r100 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r101 70 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.53 $Y=0 $X2=7.365
+ $Y2=0
r102 70 72 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=7.53 $Y=0 $X2=7.92
+ $Y2=0
r103 69 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r104 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r105 66 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r106 65 68 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r107 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r108 63 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.2 $Y=0 $X2=7.365
+ $Y2=0
r109 63 68 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=7.2 $Y=0 $X2=6.96
+ $Y2=0
r110 62 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r111 62 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r112 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r113 59 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.57 $Y=0 $X2=4.405
+ $Y2=0
r114 59 61 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=4.57 $Y=0 $X2=5.52
+ $Y2=0
r115 55 80 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.65 $Y=0 $X2=2.485
+ $Y2=0
r116 55 57 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=2.65 $Y=0 $X2=4.08
+ $Y2=0
r117 54 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.24 $Y=0 $X2=4.405
+ $Y2=0
r118 54 57 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.24 $Y=0 $X2=4.08
+ $Y2=0
r119 53 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r120 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r121 50 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r122 50 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r123 49 52 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r124 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r125 47 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r126 47 49 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r127 46 80 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.32 $Y=0 $X2=2.485
+ $Y2=0
r128 46 52 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.32 $Y=0 $X2=2.16
+ $Y2=0
r129 44 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r130 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r131 41 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r132 41 43 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r133 39 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r134 39 81 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=2.64 $Y2=0
r135 39 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r136 37 61 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=5.62 $Y=0 $X2=5.52
+ $Y2=0
r137 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.62 $Y=0 $X2=5.785
+ $Y2=0
r138 36 65 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=5.95 $Y=0 $X2=6 $Y2=0
r139 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.95 $Y=0 $X2=5.785
+ $Y2=0
r140 32 34 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=7.365 $Y=0.495
+ $X2=7.365 $Y2=0.855
r141 30 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.365 $Y=0.085
+ $X2=7.365 $Y2=0
r142 30 32 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=7.365 $Y=0.085
+ $X2=7.365 $Y2=0.495
r143 26 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.785 $Y=0.085
+ $X2=5.785 $Y2=0
r144 26 28 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=5.785 $Y=0.085
+ $X2=5.785 $Y2=0.495
r145 22 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.405 $Y=0.085
+ $X2=4.405 $Y2=0
r146 22 24 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=4.405 $Y=0.085
+ $X2=4.405 $Y2=0.83
r147 18 20 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.79 $Y=0.665
+ $X2=0.79 $Y2=1.115
r148 16 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0
r149 16 18 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0.665
r150 5 34 182 $w=1.7e-07 $l=5.84744e-07 $layer=licon1_NDIFF $count=1 $X=7.145
+ $Y=0.37 $X2=7.365 $Y2=0.855
r151 5 32 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=7.145
+ $Y=0.37 $X2=7.365 $Y2=0.495
r152 4 28 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=5.645
+ $Y=0.37 $X2=5.785 $Y2=0.495
r153 3 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.265
+ $Y=0.62 $X2=4.405 $Y2=0.83
r154 2 83 182 $w=1.7e-07 $l=2.91033e-07 $layer=licon1_NDIFF $count=1 $X=2.265
+ $Y=0.49 $X2=2.485 $Y2=0.325
r155 1 20 182 $w=1.7e-07 $l=5.03115e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.71 $X2=0.79 $Y2=1.115
r156 1 18 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.71 $X2=0.79 $Y2=0.665
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfrtp_2 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
M1000 a_390_81# D a_343_483# VPB pshort w=640000u l=180000u
+  ad=5.4e+11p pd=5.28e+06u as=1.472e+11p ps=1.74e+06u
M1001 VPWR a_2495_392# Q VPB pshort w=1.12e+06u l=180000u
+  ad=2.9811e+12p pd=2.35e+07u as=3.024e+11p ps=2.78e+06u
M1002 a_1235_119# a_1037_119# a_390_81# VPB pshort w=420000u l=180000u
+  ad=2.394e+11p pd=2.82e+06u as=0p ps=0u
M1003 Q a_2495_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=2.0718e+12p ps=1.661e+07u
M1004 VGND RESET_B a_225_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.52e+11p ps=2.88e+06u
M1005 VPWR a_2082_446# a_2040_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1006 a_1383_349# a_1235_119# VPWR VPB pshort w=1e+06u l=180000u
+  ad=4.6755e+11p pd=3.07e+06u as=0p ps=0u
M1007 VGND RESET_B a_1432_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1008 a_547_81# SCE a_390_81# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.927e+11p ps=3.55e+06u
M1009 a_2078_74# a_837_119# a_1824_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=5.504e+11p ps=3.72e+06u
M1010 VGND a_2082_446# a_2078_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR SCE a_27_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1012 a_343_483# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1235_119# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_312_81# a_27_74# a_225_81# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1015 a_390_81# D a_312_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND CLK a_837_119# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.0225e+11p ps=2.04e+06u
M1017 a_1037_119# a_837_119# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.998e+11p pd=2.02e+06u as=0p ps=0u
M1018 a_2082_446# a_1824_74# a_2242_74# VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1019 a_2082_446# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1020 a_1824_74# a_837_119# a_1383_349# VPB pshort w=1e+06u l=180000u
+  ad=4.2595e+11p pd=3.6e+06u as=0p ps=0u
M1021 a_2040_508# a_1037_119# a_1824_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1432_119# a_1383_349# a_1354_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1023 a_390_81# RESET_B VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_1824_74# a_2082_446# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_1339_457# a_837_119# a_1235_119# VPB pshort w=420000u l=180000u
+  ad=9.24e+10p pd=1.28e+06u as=0p ps=0u
M1026 a_2242_74# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR CLK a_837_119# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1028 a_1824_74# a_1037_119# a_1383_349# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.627e+11p ps=2.19e+06u
M1029 a_2495_392# a_1824_74# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1030 VGND a_2495_392# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1235_119# a_837_119# a_390_81# VNB nlowvt w=420000u l=150000u
+  ad=1.869e+11p pd=1.73e+06u as=0p ps=0u
M1032 a_1354_119# a_1037_119# a_1235_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR a_1383_349# a_1339_457# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1037_119# a_837_119# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1035 a_225_81# SCD a_547_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND SCE a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1037 a_2495_392# a_1824_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1038 a_517_483# a_27_74# a_390_81# VPB pshort w=640000u l=180000u
+  ad=2.304e+11p pd=2e+06u as=0p ps=0u
M1039 VPWR SCD a_517_483# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1383_349# a_1235_119# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 Q a_2495_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_ms__a311o_1.pex.spice
* Created: Wed Sep  2 11:54:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A311O_1%A_89_270# 1 2 3 12 14 16 17 18 19 23 27 36
+ 42 43 44 48
c99 48 0 1.98395e-19 $X=0.735 $Y=1.515
c100 36 0 1.72877e-19 $X=2.405 $Y=1.005
c101 19 0 1.06923e-19 $X=3.245 $Y=1.53
c102 17 0 4.83091e-20 $X=2.24 $Y=1.195
r103 42 43 5.27442 $w=4.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.34 $Y=2.105
+ $X2=3.34 $Y2=1.94
r104 38 39 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.405 $Y=1.195
+ $X2=2.405 $Y2=1.53
r105 36 38 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.405 $Y=1.005
+ $X2=2.405 $Y2=1.195
r106 34 48 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.645 $Y=1.515
+ $X2=0.735 $Y2=1.515
r107 34 45 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=0.645 $Y=1.515
+ $X2=0.535 $Y2=1.515
r108 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.645
+ $Y=1.515 $X2=0.645 $Y2=1.515
r109 29 44 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.41 $Y=1.615
+ $X2=3.41 $Y2=1.53
r110 29 43 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.41 $Y=1.615
+ $X2=3.41 $Y2=1.94
r111 25 44 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.41 $Y=1.445
+ $X2=3.41 $Y2=1.53
r112 25 27 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=3.41 $Y=1.445
+ $X2=3.41 $Y2=1.105
r113 21 42 1.78139 $w=4.68e-07 $l=7e-08 $layer=LI1_cond $X=3.34 $Y=2.175
+ $X2=3.34 $Y2=2.105
r114 21 23 16.287 $w=4.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.34 $Y=2.175
+ $X2=3.34 $Y2=2.815
r115 20 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.57 $Y=1.53
+ $X2=2.405 $Y2=1.53
r116 19 44 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=1.53
+ $X2=3.41 $Y2=1.53
r117 19 20 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=3.245 $Y=1.53
+ $X2=2.57 $Y2=1.53
r118 18 33 11.4824 $w=3.4e-07 $l=4.20666e-07 $layer=LI1_cond $X=0.945 $Y=1.195
+ $X2=0.712 $Y2=1.515
r119 17 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=1.195
+ $X2=2.405 $Y2=1.195
r120 17 18 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=2.24 $Y=1.195
+ $X2=0.945 $Y2=1.195
r121 14 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.735 $Y=1.35
+ $X2=0.735 $Y2=1.515
r122 14 16 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.735 $Y=1.35
+ $X2=0.735 $Y2=0.87
r123 10 45 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.68
+ $X2=0.535 $Y2=1.515
r124 10 12 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.535 $Y=1.68
+ $X2=0.535 $Y2=2.4
r125 3 42 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.135
+ $Y=1.96 $X2=3.27 $Y2=2.105
r126 3 23 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.135
+ $Y=1.96 $X2=3.27 $Y2=2.815
r127 2 27 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=3.27
+ $Y=0.615 $X2=3.41 $Y2=1.105
r128 1 36 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=2.265
+ $Y=0.615 $X2=2.405 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_1%A3 3 7 9 12
c36 9 0 1.98395e-19 $X=1.2 $Y=1.665
c37 7 0 1.5978e-19 $X=1.245 $Y=0.92
r38 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=1.615
+ $X2=1.2 $Y2=1.78
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=1.615
+ $X2=1.2 $Y2=1.45
r40 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.2
+ $Y=1.615 $X2=1.2 $Y2=1.615
r41 7 14 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.245 $Y=0.92
+ $X2=1.245 $Y2=1.45
r42 3 15 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=1.215 $Y=2.46
+ $X2=1.215 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_1%A2 3 7 9 12
c34 12 0 1.72877e-19 $X=1.74 $Y=1.615
c35 7 0 1.69592e-19 $X=1.72 $Y=0.935
c36 3 0 4.60934e-20 $X=1.665 $Y=2.46
r37 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.74 $Y=1.615
+ $X2=1.74 $Y2=1.78
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.74 $Y=1.615
+ $X2=1.74 $Y2=1.45
r39 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.74
+ $Y=1.615 $X2=1.74 $Y2=1.615
r40 7 14 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=1.72 $Y=0.935
+ $X2=1.72 $Y2=1.45
r41 3 15 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=1.665 $Y=2.46
+ $X2=1.665 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_1%A1 4 5 7 10 11 15 16 19
c50 16 0 1.83039e-19 $X=2.17 $Y=0.34
c51 15 0 1.46334e-19 $X=2.17 $Y=0.34
c52 7 0 1.06923e-19 $X=2.205 $Y=2.46
r53 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=0.34
+ $X2=2.17 $Y2=0.505
r54 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.17
+ $Y=0.34 $X2=2.17 $Y2=0.34
r55 11 16 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.17 $Y=0.555
+ $X2=2.17 $Y2=0.34
r56 11 19 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.17 $Y=0.555
+ $X2=2.005 $Y2=0.555
r57 10 19 16.2845 $w=2.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.68 $Y=0.555
+ $X2=2.005 $Y2=0.555
r58 5 9 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.205 $Y=1.42 $X2=2.205
+ $Y2=1.33
r59 5 7 404.258 $w=1.8e-07 $l=1.04e-06 $layer=POLY_cond $X=2.205 $Y=1.42
+ $X2=2.205 $Y2=2.46
r60 4 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.19 $Y=0.935
+ $X2=2.19 $Y2=1.33
r61 4 18 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.19 $Y=0.935
+ $X2=2.19 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_1%B1 4 7 10 11 14
c41 10 0 1.12525e-19 $X=2.645 $Y=1.48
c42 4 0 4.83091e-20 $X=2.62 $Y=0.935
r43 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=0.34
+ $X2=2.71 $Y2=0.505
r44 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.71
+ $Y=0.34 $X2=2.71 $Y2=0.34
r45 11 15 9.04483 $w=2.9e-07 $l=2.15e-07 $layer=LI1_cond $X=2.7 $Y=0.555 $X2=2.7
+ $Y2=0.34
r46 9 10 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.645 $Y=1.33
+ $X2=2.645 $Y2=1.48
r47 7 10 380.935 $w=1.8e-07 $l=9.8e-07 $layer=POLY_cond $X=2.655 $Y=2.46
+ $X2=2.655 $Y2=1.48
r48 4 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.62 $Y=0.935
+ $X2=2.62 $Y2=1.33
r49 4 17 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.62 $Y=0.935
+ $X2=2.62 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_1%C1 3 8 11 13 14 17 18
r40 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=0.34 $X2=3.55 $Y2=0.34
r41 14 18 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=3.55 $Y=0.555
+ $X2=3.55 $Y2=0.34
r42 13 17 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=3.27 $Y=0.34
+ $X2=3.55 $Y2=0.34
r43 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.195 $Y=1.33
+ $X2=3.195 $Y2=1.405
r44 6 8 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.195 $Y=1.33
+ $X2=3.195 $Y2=0.935
r45 5 13 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.195 $Y=0.505
+ $X2=3.27 $Y2=0.34
r46 5 8 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.195 $Y=0.505
+ $X2=3.195 $Y2=0.935
r47 1 11 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.045 $Y=1.405
+ $X2=3.195 $Y2=1.405
r48 1 3 380.935 $w=1.8e-07 $l=9.8e-07 $layer=POLY_cond $X=3.045 $Y=1.48
+ $X2=3.045 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_1%X 1 2 9 11 17 18 19 26 35
r21 24 26 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=0.3 $Y=2.025 $X2=0.3
+ $Y2=2.035
r22 18 19 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.3 $Y=2.405 $X2=0.3
+ $Y2=2.775
r23 17 24 1.25122 $w=3.48e-07 $l=3.8e-08 $layer=LI1_cond $X=0.3 $Y=1.987 $X2=0.3
+ $Y2=2.025
r24 17 35 7.56653 $w=3.48e-07 $l=1.37e-07 $layer=LI1_cond $X=0.3 $Y=1.987
+ $X2=0.3 $Y2=1.85
r25 17 18 10.9647 $w=3.48e-07 $l=3.33e-07 $layer=LI1_cond $X=0.3 $Y=2.072
+ $X2=0.3 $Y2=2.405
r26 17 26 1.2183 $w=3.48e-07 $l=3.7e-08 $layer=LI1_cond $X=0.3 $Y=2.072 $X2=0.3
+ $Y2=2.035
r27 9 13 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.48 $Y=1.095 $X2=0.21
+ $Y2=1.095
r28 9 11 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=0.48 $Y=1.01
+ $X2=0.48 $Y2=0.645
r29 7 13 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.21 $Y=1.18 $X2=0.21
+ $Y2=1.095
r30 7 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.21 $Y=1.18 $X2=0.21
+ $Y2=1.85
r31 2 17 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.185
+ $Y=1.84 $X2=0.31 $Y2=2.015
r32 2 19 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.185
+ $Y=1.84 $X2=0.31 $Y2=2.815
r33 1 11 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.395
+ $Y=0.5 $X2=0.52 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_1%VPWR 1 2 11 17 20 21 22 32 33 36
r43 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r45 30 33 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r46 29 32 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r47 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 27 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 24 36 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=1.105 $Y=3.33
+ $X2=0.875 $Y2=3.33
r51 24 26 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=1.105 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 22 30 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 22 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 20 26 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.805 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 20 21 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.805 $Y=3.33
+ $X2=1.95 $Y2=3.33
r56 19 29 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 19 21 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.095 $Y=3.33
+ $X2=1.95 $Y2=3.33
r58 15 21 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.95 $Y=3.245
+ $X2=1.95 $Y2=3.33
r59 15 17 31.3941 $w=2.88e-07 $l=7.9e-07 $layer=LI1_cond $X=1.95 $Y=3.245
+ $X2=1.95 $Y2=2.455
r60 11 14 18.2012 $w=4.58e-07 $l=7e-07 $layer=LI1_cond $X=0.875 $Y=2.115
+ $X2=0.875 $Y2=2.815
r61 9 36 1.85547 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.875 $Y=3.245
+ $X2=0.875 $Y2=3.33
r62 9 14 11.1807 $w=4.58e-07 $l=4.3e-07 $layer=LI1_cond $X=0.875 $Y=3.245
+ $X2=0.875 $Y2=2.815
r63 2 17 300 $w=1.7e-07 $l=5.6723e-07 $layer=licon1_PDIFF $count=2 $X=1.755
+ $Y=1.96 $X2=1.91 $Y2=2.455
r64 1 14 400 $w=1.7e-07 $l=1.09287e-06 $layer=licon1_PDIFF $count=1 $X=0.625
+ $Y=1.84 $X2=0.875 $Y2=2.815
r65 1 11 400 $w=1.7e-07 $l=3.79967e-07 $layer=licon1_PDIFF $count=1 $X=0.625
+ $Y=1.84 $X2=0.875 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_1%A_261_392# 1 2 7 9 11 13 15
c41 13 0 1.58618e-19 $X=2.43 $Y=2.12
r42 13 20 2.68829 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.43 $Y=2.12 $X2=2.43
+ $Y2=2.03
r43 13 15 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.43 $Y=2.12
+ $X2=2.43 $Y2=2.815
r44 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.605 $Y=2.035
+ $X2=1.44 $Y2=2.035
r45 11 20 5.07788 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=2.265 $Y=2.035
+ $X2=2.43 $Y2=2.03
r46 11 12 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=2.265 $Y=2.035
+ $X2=1.605 $Y2=2.035
r47 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.44 $Y=2.12 $X2=1.44
+ $Y2=2.035
r48 7 9 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.44 $Y=2.12 $X2=1.44
+ $Y2=2.815
r49 2 20 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.295
+ $Y=1.96 $X2=2.43 $Y2=2.105
r50 2 15 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.295
+ $Y=1.96 $X2=2.43 $Y2=2.815
r51 1 18 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=1.305
+ $Y=1.96 $X2=1.44 $Y2=2.115
r52 1 9 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.305
+ $Y=1.96 $X2=1.44 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__A311O_1%VGND 1 2 9 12 14 15 18 24 30 31 34
r48 34 35 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r49 31 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r50 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r51 28 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.13
+ $Y2=0
r52 28 30 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.6
+ $Y2=0
r53 26 27 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 24 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.045 $Y=0 $X2=3.13
+ $Y2=0
r55 24 26 120.369 $w=1.68e-07 $l=1.845e-06 $layer=LI1_cond $X=3.045 $Y=0 $X2=1.2
+ $Y2=0
r56 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r57 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r58 18 35 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=3.12
+ $Y2=0
r59 18 27 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r60 14 21 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=0.785 $Y=0 $X2=0.72
+ $Y2=0
r61 14 15 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.785 $Y=0 $X2=0.95
+ $Y2=0
r62 13 26 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.2
+ $Y2=0
r63 13 15 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=0.95
+ $Y2=0
r64 12 17 15.8187 $w=3.2e-07 $l=4.12414e-07 $layer=LI1_cond $X=3.13 $Y=0.675
+ $X2=2.982 $Y2=1.02
r65 11 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=0.085
+ $X2=3.13 $Y2=0
r66 11 12 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.13 $Y=0.085
+ $X2=3.13 $Y2=0.675
r67 7 15 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.95 $Y=0.085 $X2=0.95
+ $Y2=0
r68 7 9 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=0.95 $Y=0.085 $X2=0.95
+ $Y2=0.775
r69 2 17 182 $w=1.7e-07 $l=5.03115e-07 $layer=licon1_NDIFF $count=1 $X=2.695
+ $Y=0.615 $X2=2.915 $Y2=1.02
r70 1 9 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.81
+ $Y=0.5 $X2=0.95 $Y2=0.775
.ends


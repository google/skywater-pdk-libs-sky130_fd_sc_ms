* File: sky130_fd_sc_ms__dlxbp_1.spice
* Created: Wed Sep  2 12:06:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dlxbp_1.pex.spice"
.subckt sky130_fd_sc_ms__dlxbp_1  VNB VPB D GATE VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_D_M1005_g N_A_27_413#_M1005_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.129591 AS=0.15675 PD=0.997674 PS=1.67 NRD=18 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1002 N_A_231_74#_M1002_d N_GATE_M1002_g N_VGND_M1005_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1019 N_VGND_M1019_d N_A_231_74#_M1019_g N_A_373_82#_M1019_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.224922 AS=0.2109 PD=1.57116 PS=2.05 NRD=40.368 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002 A=0.111 P=1.78 MULT=1
MM1012 A_589_80# N_A_27_413#_M1012_g N_VGND_M1019_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.194528 PD=0.88 PS=1.35884 NRD=12.18 NRS=21.552 M=1 R=4.26667
+ SA=75000.8 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1011 N_A_667_80#_M1011_d N_A_373_82#_M1011_g A_589_80# VNB NLOWVT L=0.15
+ W=0.64 AD=0.182823 AS=0.0768 PD=1.48528 PS=0.88 NRD=29.052 NRS=12.18 M=1
+ R=4.26667 SA=75001.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1003 A_815_124# N_A_231_74#_M1003_g N_A_667_80#_M1011_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.119977 PD=0.66 PS=0.974717 NRD=18.564 NRS=44.28 M=1
+ R=2.8 SA=75002 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_863_98#_M1020_g A_815_124# VNB NLOWVT L=0.15 W=0.42
+ AD=0.106521 AS=0.0504 PD=0.847241 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8
+ SA=75002.4 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1007 N_A_863_98#_M1007_d N_A_667_80#_M1007_g N_VGND_M1020_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.187679 PD=2.05 PS=1.49276 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_A_863_98#_M1015_g N_Q_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.137674 AS=0.2072 PD=1.25054 PS=2.04 NRD=5.664 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1018 N_A_1350_116#_M1018_d N_A_863_98#_M1018_g N_VGND_M1015_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.15675 AS=0.102326 PD=1.67 PS=0.929457 NRD=0 NRS=7.632 M=1
+ R=3.66667 SA=75000.7 SB=75000.2 A=0.0825 P=1.4 MULT=1
MM1008 N_Q_N_M1008_d N_A_1350_116#_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_VPWR_M1010_d N_D_M1010_g N_A_27_413#_M1010_s VPB PSHORT L=0.18 W=0.84
+ AD=0.2212 AS=0.231 PD=1.56 PS=2.23 NRD=48.856 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1013 N_A_231_74#_M1013_d N_GATE_M1013_g N_VPWR_M1010_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.2212 PD=2.24 PS=1.56 NRD=0 NRS=48.856 M=1 R=4.66667
+ SA=90000.8 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1000 N_VPWR_M1000_d N_A_231_74#_M1000_g N_A_373_82#_M1000_s VPB PSHORT L=0.18
+ W=0.84 AD=0.210023 AS=0.2352 PD=1.42891 PS=2.24 NRD=45.7237 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90001.8 A=0.1512 P=2.04 MULT=1
MM1001 A_589_392# N_A_27_413#_M1001_g N_VPWR_M1000_d VPB PSHORT L=0.18 W=1
+ AD=0.105 AS=0.250027 PD=1.21 PS=1.70109 NRD=9.8303 NRS=16.7253 M=1 R=5.55556
+ SA=90000.7 SB=90001.4 A=0.18 P=2.36 MULT=1
MM1016 N_A_667_80#_M1016_d N_A_231_74#_M1016_g A_589_392# VPB PSHORT L=0.18 W=1
+ AD=0.215845 AS=0.105 PD=1.90141 PS=1.21 NRD=0 NRS=9.8303 M=1 R=5.55556
+ SA=90001.1 SB=90001 A=0.18 P=2.36 MULT=1
MM1021 A_773_508# N_A_373_82#_M1021_g N_A_667_80#_M1016_d VPB PSHORT L=0.18
+ W=0.42 AD=0.09975 AS=0.0906549 PD=0.895 PS=0.798592 NRD=85.5965 NRS=75.4313
+ M=1 R=2.33333 SA=90001.5 SB=90001.6 A=0.0756 P=1.2 MULT=1
MM1006 N_VPWR_M1006_d N_A_863_98#_M1006_g A_773_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.109009 AS=0.09975 PD=0.902727 PS=0.895 NRD=46.886 NRS=85.5965 M=1
+ R=2.33333 SA=90002.2 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1004 N_A_863_98#_M1004_d N_A_667_80#_M1004_g N_VPWR_M1006_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.290691 PD=2.8 PS=2.40727 NRD=0 NRS=27.2451 M=1 R=6.22222
+ SA=90001.2 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1017 N_VPWR_M1017_d N_A_863_98#_M1017_g N_Q_M1017_s VPB PSHORT L=0.18 W=1.12
+ AD=0.196 AS=0.3136 PD=1.65143 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1014 N_A_1350_116#_M1014_d N_A_863_98#_M1014_g N_VPWR_M1017_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.231 AS=0.147 PD=2.23 PS=1.23857 NRD=0 NRS=11.7215 M=1
+ R=4.66667 SA=90000.7 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1009 N_Q_N_M1009_d N_A_1350_116#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.18
+ W=1.12 AD=0.308 AS=0.308 PD=2.79 PS=2.79 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX22_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_ms__dlxbp_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__a2bb2oi_4.pex.spice
* Created: Wed Sep  2 11:54:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A2BB2OI_4%A2_N 3 7 9 10 11 13 14 15 16 22
c50 7 0 3.35904e-19 $X=0.945 $Y=2.46
r51 29 30 43.6418 $w=4.97e-07 $l=4.5e-07 $layer=POLY_cond $X=0.495 $Y=1.477
+ $X2=0.945 $Y2=1.477
r52 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.29
+ $Y=1.605 $X2=0.29 $Y2=1.605
r53 20 29 15.0322 $w=4.97e-07 $l=1.55e-07 $layer=POLY_cond $X=0.34 $Y=1.477
+ $X2=0.495 $Y2=1.477
r54 20 26 4.84909 $w=4.97e-07 $l=5e-08 $layer=POLY_cond $X=0.34 $Y=1.477
+ $X2=0.29 $Y2=1.477
r55 20 22 91.1834 $w=4.3e-07 $l=7.05e-07 $layer=POLY_cond $X=0.34 $Y=1.29
+ $X2=0.34 $Y2=0.585
r56 16 27 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.605
r57 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=0.925
+ $X2=0.29 $Y2=1.295
r58 14 15 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=0.555
+ $X2=0.29 $Y2=0.925
r59 14 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.29
+ $Y=0.585 $X2=0.29 $Y2=0.585
r60 11 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.32 $Y=1.185
+ $X2=1.32 $Y2=0.74
r61 10 30 34.5746 $w=4.97e-07 $l=2.58107e-07 $layer=POLY_cond $X=1.035 $Y=1.26
+ $X2=0.945 $Y2=1.477
r62 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.245 $Y=1.26
+ $X2=1.32 $Y2=1.185
r63 9 10 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.245 $Y=1.26
+ $X2=1.035 $Y2=1.26
r64 5 30 26.715 $w=1.8e-07 $l=2.93e-07 $layer=POLY_cond $X=0.945 $Y=1.77
+ $X2=0.945 $Y2=1.477
r65 5 7 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=0.945 $Y=1.77 $X2=0.945
+ $Y2=2.46
r66 1 29 26.715 $w=1.8e-07 $l=2.93e-07 $layer=POLY_cond $X=0.495 $Y=1.77
+ $X2=0.495 $Y2=1.477
r67 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=0.495 $Y=1.77 $X2=0.495
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_4%A1_N 3 7 11 13 14 20
c47 20 0 6.19774e-20 $X=1.77 $Y=1.635
c48 7 0 3.63668e-19 $X=1.75 $Y=0.74
r49 20 22 14.8156 $w=2.44e-07 $l=7.5e-08 $layer=POLY_cond $X=1.77 $Y=1.635
+ $X2=1.845 $Y2=1.635
r50 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.77
+ $Y=1.635 $X2=1.77 $Y2=1.635
r51 18 20 3.95082 $w=2.44e-07 $l=2e-08 $layer=POLY_cond $X=1.75 $Y=1.635
+ $X2=1.77 $Y2=1.635
r52 14 21 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.16 $Y=1.635
+ $X2=1.77 $Y2=1.635
r53 13 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.68 $Y=1.635 $X2=1.77
+ $Y2=1.635
r54 9 22 9.95785 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.8
+ $X2=1.845 $Y2=1.635
r55 9 11 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.845 $Y=1.8
+ $X2=1.845 $Y2=2.46
r56 5 18 14.1583 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.47
+ $X2=1.75 $Y2=1.635
r57 5 7 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=1.75 $Y=1.47 $X2=1.75
+ $Y2=0.74
r58 1 18 70.1271 $w=2.44e-07 $l=4.29651e-07 $layer=POLY_cond $X=1.395 $Y=1.8
+ $X2=1.75 $Y2=1.635
r59 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.395 $Y=1.8 $X2=1.395
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_4%A_117_392# 1 2 7 9 11 12 14 17 19 21 24 26
+ 28 29 33 35 39 41 44 46 47 50 54 56 59 63 65 72
c140 54 0 6.19774e-20 $X=2.995 $Y=1.34
c141 33 0 1.69337e-19 $X=3.945 $Y=2.4
c142 26 0 1.39795e-19 $X=3.51 $Y=1.22
c143 19 0 1.39795e-19 $X=3.08 $Y=1.22
c144 12 0 1.44963e-19 $X=2.65 $Y=1.22
r145 71 72 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.51 $Y=1.385
+ $X2=3.585 $Y2=1.385
r146 70 71 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.495 $Y=1.385
+ $X2=3.51 $Y2=1.385
r147 67 68 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=3.045 $Y=1.385
+ $X2=3.08 $Y2=1.385
r148 64 65 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.65 $Y=1.385
+ $X2=2.575 $Y2=1.385
r149 62 67 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=2.74 $Y=1.385
+ $X2=3.045 $Y2=1.385
r150 62 64 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.74 $Y=1.385
+ $X2=2.65 $Y2=1.385
r151 61 63 8.7366 $w=4.18e-07 $l=1.65e-07 $layer=LI1_cond $X=2.74 $Y=1.34
+ $X2=2.575 $Y2=1.34
r152 61 62 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.74
+ $Y=1.385 $X2=2.74 $Y2=1.385
r153 57 70 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.42 $Y=1.385
+ $X2=3.495 $Y2=1.385
r154 57 68 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.42 $Y=1.385
+ $X2=3.08 $Y2=1.385
r155 56 57 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.42
+ $Y=1.385 $X2=3.42 $Y2=1.385
r156 54 61 6.99698 $w=4.18e-07 $l=2.55e-07 $layer=LI1_cond $X=2.995 $Y=1.34
+ $X2=2.74 $Y2=1.34
r157 54 56 11.6616 $w=4.18e-07 $l=4.25e-07 $layer=LI1_cond $X=2.995 $Y=1.34
+ $X2=3.42 $Y2=1.34
r158 53 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=1.215
+ $X2=1.535 $Y2=1.215
r159 53 63 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.62 $Y=1.215
+ $X2=2.575 $Y2=1.215
r160 48 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=1.13
+ $X2=1.535 $Y2=1.215
r161 48 50 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.535 $Y=1.13
+ $X2=1.535 $Y2=0.515
r162 46 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.45 $Y=1.215
+ $X2=1.535 $Y2=1.215
r163 46 47 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.45 $Y=1.215
+ $X2=0.885 $Y2=1.215
r164 42 47 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.76 $Y=1.3
+ $X2=0.885 $Y2=1.215
r165 42 44 37.1087 $w=2.48e-07 $l=8.05e-07 $layer=LI1_cond $X=0.76 $Y=1.3
+ $X2=0.76 $Y2=2.105
r166 37 39 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=4.395 $Y=1.55
+ $X2=4.395 $Y2=2.4
r167 36 41 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.035 $Y=1.475
+ $X2=3.945 $Y2=1.475
r168 35 37 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.305 $Y=1.475
+ $X2=4.395 $Y2=1.55
r169 35 36 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.305 $Y=1.475
+ $X2=4.035 $Y2=1.475
r170 31 41 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.945 $Y=1.55
+ $X2=3.945 $Y2=1.475
r171 31 33 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.945 $Y=1.55
+ $X2=3.945 $Y2=2.4
r172 29 41 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.855 $Y=1.475
+ $X2=3.945 $Y2=1.475
r173 29 72 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.855 $Y=1.475
+ $X2=3.585 $Y2=1.475
r174 26 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.51 $Y=1.22
+ $X2=3.51 $Y2=1.385
r175 26 28 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.51 $Y=1.22
+ $X2=3.51 $Y2=0.74
r176 22 70 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.495 $Y=1.55
+ $X2=3.495 $Y2=1.385
r177 22 24 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.495 $Y=1.55
+ $X2=3.495 $Y2=2.4
r178 19 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.08 $Y=1.22
+ $X2=3.08 $Y2=1.385
r179 19 21 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.08 $Y=1.22
+ $X2=3.08 $Y2=0.74
r180 15 67 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.045 $Y=1.55
+ $X2=3.045 $Y2=1.385
r181 15 17 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.045 $Y=1.55
+ $X2=3.045 $Y2=2.4
r182 12 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.65 $Y=1.22
+ $X2=2.65 $Y2=1.385
r183 12 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.65 $Y=1.22
+ $X2=2.65 $Y2=0.74
r184 11 65 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.295 $Y=1.295
+ $X2=2.575 $Y2=1.295
r185 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.22 $Y=1.22
+ $X2=2.295 $Y2=1.295
r186 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.22 $Y=1.22 $X2=2.22
+ $Y2=0.74
r187 2 44 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.96 $X2=0.72 $Y2=2.105
r188 1 50 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.395
+ $Y=0.37 $X2=1.535 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_4%B2 3 7 11 15 19 23 27 31 33 34 35 36 55
c86 36 0 1.69337e-19 $X=6 $Y=1.665
r87 54 55 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=6.195 $Y=1.515
+ $X2=6.2 $Y2=1.515
r88 52 54 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=5.94 $Y=1.515
+ $X2=6.195 $Y2=1.515
r89 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.94
+ $Y=1.515 $X2=5.94 $Y2=1.515
r90 50 52 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=5.77 $Y=1.515
+ $X2=5.94 $Y2=1.515
r91 49 50 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=5.745 $Y=1.515
+ $X2=5.77 $Y2=1.515
r92 48 49 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=5.34 $Y=1.515
+ $X2=5.745 $Y2=1.515
r93 47 48 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=5.295 $Y=1.515
+ $X2=5.34 $Y2=1.515
r94 45 47 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=4.92 $Y=1.515
+ $X2=5.295 $Y2=1.515
r95 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.92
+ $Y=1.515 $X2=4.92 $Y2=1.515
r96 43 45 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=4.91 $Y=1.515 $X2=4.92
+ $Y2=1.515
r97 41 43 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=4.845 $Y=1.515
+ $X2=4.91 $Y2=1.515
r98 36 53 1.60806 $w=4.28e-07 $l=6e-08 $layer=LI1_cond $X=6 $Y=1.565 $X2=5.94
+ $Y2=1.565
r99 35 53 11.2564 $w=4.28e-07 $l=4.2e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.94 $Y2=1.565
r100 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.52 $Y2=1.565
r101 34 46 3.21612 $w=4.28e-07 $l=1.2e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=4.92 $Y2=1.565
r102 33 46 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.92 $Y2=1.565
r103 29 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.2 $Y=1.35
+ $X2=6.2 $Y2=1.515
r104 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.2 $Y=1.35 $X2=6.2
+ $Y2=0.74
r105 25 54 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.195 $Y=1.68
+ $X2=6.195 $Y2=1.515
r106 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.195 $Y=1.68
+ $X2=6.195 $Y2=2.4
r107 21 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.77 $Y=1.35
+ $X2=5.77 $Y2=1.515
r108 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.77 $Y=1.35
+ $X2=5.77 $Y2=0.74
r109 17 49 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.745 $Y=1.68
+ $X2=5.745 $Y2=1.515
r110 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.745 $Y=1.68
+ $X2=5.745 $Y2=2.4
r111 13 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.34 $Y=1.35
+ $X2=5.34 $Y2=1.515
r112 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.34 $Y=1.35
+ $X2=5.34 $Y2=0.74
r113 9 47 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.295 $Y=1.68
+ $X2=5.295 $Y2=1.515
r114 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.295 $Y=1.68
+ $X2=5.295 $Y2=2.4
r115 5 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.91 $Y=1.35
+ $X2=4.91 $Y2=1.515
r116 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.91 $Y=1.35 $X2=4.91
+ $Y2=0.74
r117 1 41 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.845 $Y=1.68
+ $X2=4.845 $Y2=1.515
r118 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.845 $Y=1.68
+ $X2=4.845 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_4%B1 3 7 11 15 19 23 27 31 33 34 35 36 54
c83 3 0 2.04552e-19 $X=6.63 $Y=0.74
r84 52 54 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.92 $Y=1.515
+ $X2=7.995 $Y2=1.515
r85 50 52 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=7.545 $Y=1.515
+ $X2=7.92 $Y2=1.515
r86 49 50 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=7.49 $Y=1.515
+ $X2=7.545 $Y2=1.515
r87 48 49 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=7.095 $Y=1.515
+ $X2=7.49 $Y2=1.515
r88 47 48 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=7.06 $Y=1.515
+ $X2=7.095 $Y2=1.515
r89 45 47 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=6.9 $Y=1.515
+ $X2=7.06 $Y2=1.515
r90 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.9
+ $Y=1.515 $X2=6.9 $Y2=1.515
r91 43 45 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=6.645 $Y=1.515
+ $X2=6.9 $Y2=1.515
r92 41 43 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.63 $Y=1.515
+ $X2=6.645 $Y2=1.515
r93 35 36 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.92 $Y=1.565
+ $X2=8.4 $Y2=1.565
r94 35 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.92
+ $Y=1.515 $X2=7.92 $Y2=1.515
r95 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.92 $Y2=1.565
r96 33 34 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.44 $Y2=1.565
r97 33 46 1.60806 $w=4.28e-07 $l=6e-08 $layer=LI1_cond $X=6.96 $Y=1.565 $X2=6.9
+ $Y2=1.565
r98 29 54 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.995 $Y=1.68
+ $X2=7.995 $Y2=1.515
r99 29 31 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.995 $Y=1.68
+ $X2=7.995 $Y2=2.4
r100 25 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.92 $Y=1.35
+ $X2=7.92 $Y2=1.515
r101 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.92 $Y=1.35
+ $X2=7.92 $Y2=0.74
r102 21 50 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.545 $Y=1.68
+ $X2=7.545 $Y2=1.515
r103 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.545 $Y=1.68
+ $X2=7.545 $Y2=2.4
r104 17 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.49 $Y=1.35
+ $X2=7.49 $Y2=1.515
r105 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.49 $Y=1.35
+ $X2=7.49 $Y2=0.74
r106 13 48 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.095 $Y=1.68
+ $X2=7.095 $Y2=1.515
r107 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.095 $Y=1.68
+ $X2=7.095 $Y2=2.4
r108 9 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.06 $Y=1.35
+ $X2=7.06 $Y2=1.515
r109 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.06 $Y=1.35
+ $X2=7.06 $Y2=0.74
r110 5 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.645 $Y=1.68
+ $X2=6.645 $Y2=1.515
r111 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.645 $Y=1.68
+ $X2=6.645 $Y2=2.4
r112 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.63 $Y=1.35
+ $X2=6.63 $Y2=1.515
r113 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.63 $Y=1.35 $X2=6.63
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_4%A_29_392# 1 2 3 12 16 17 18 22 24 26
c45 18 0 1.47912e-19 $X=1.17 $Y=2.14
r46 24 31 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=2.14 $X2=2.07
+ $Y2=2.055
r47 24 26 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.07 $Y=2.14
+ $X2=2.07 $Y2=2.815
r48 23 29 3.40825 $w=1.7e-07 $l=9.21954e-08 $layer=LI1_cond $X=1.255 $Y=2.055
+ $X2=1.17 $Y2=2.04
r49 22 31 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=2.055
+ $X2=2.07 $Y2=2.055
r50 22 23 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.905 $Y=2.055
+ $X2=1.255 $Y2=2.055
r51 19 21 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.17 $Y=2.905 $X2=1.17
+ $Y2=2.815
r52 18 29 3.40825 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.17 $Y=2.14 $X2=1.17
+ $Y2=2.04
r53 18 21 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.17 $Y=2.14
+ $X2=1.17 $Y2=2.815
r54 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.085 $Y=2.99
+ $X2=1.17 $Y2=2.905
r55 16 17 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.085 $Y=2.99
+ $X2=0.435 $Y2=2.99
r56 12 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.27 $Y=2.105
+ $X2=0.27 $Y2=2.815
r57 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.27 $Y=2.905
+ $X2=0.435 $Y2=2.99
r58 10 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=2.905 $X2=0.27
+ $Y2=2.815
r59 3 31 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=1.96 $X2=2.07 $Y2=2.135
r60 3 26 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=1.96 $X2=2.07 $Y2=2.815
r61 2 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.96 $X2=1.17 $Y2=2.105
r62 2 21 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.96 $X2=1.17 $Y2=2.815
r63 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.96 $X2=0.27 $Y2=2.815
r64 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.96 $X2=0.27 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_4%VPWR 1 2 3 4 5 18 20 24 28 32 36 39 40 42
+ 43 44 46 54 67 68 71 74 77
c104 18 0 1.87992e-19 $X=1.62 $Y=2.475
r105 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r106 74 75 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r107 71 72 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r108 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r109 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r110 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r111 62 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r112 62 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r113 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r114 59 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.135 $Y=3.33
+ $X2=6.01 $Y2=3.33
r115 59 61 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.135 $Y=3.33
+ $X2=6.48 $Y2=3.33
r116 58 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r117 58 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r118 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r119 55 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.155 $Y=3.33
+ $X2=5.07 $Y2=3.33
r120 55 57 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.155 $Y=3.33
+ $X2=5.52 $Y2=3.33
r121 54 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.885 $Y=3.33
+ $X2=6.01 $Y2=3.33
r122 54 57 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.885 $Y=3.33
+ $X2=5.52 $Y2=3.33
r123 53 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r124 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r125 49 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r126 48 52 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r127 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r128 46 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.455 $Y=3.33
+ $X2=1.58 $Y2=3.33
r129 46 52 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.455 $Y=3.33
+ $X2=1.2 $Y2=3.33
r130 44 75 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=5.04 $Y2=3.33
r131 44 72 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=1.68 $Y2=3.33
r132 42 64 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.685 $Y=3.33
+ $X2=7.44 $Y2=3.33
r133 42 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.685 $Y=3.33
+ $X2=7.77 $Y2=3.33
r134 41 67 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=7.855 $Y=3.33
+ $X2=8.4 $Y2=3.33
r135 41 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.855 $Y=3.33
+ $X2=7.77 $Y2=3.33
r136 39 61 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.705 $Y=3.33
+ $X2=6.48 $Y2=3.33
r137 39 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.705 $Y=3.33
+ $X2=6.83 $Y2=3.33
r138 38 64 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=6.955 $Y=3.33
+ $X2=7.44 $Y2=3.33
r139 38 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.955 $Y=3.33
+ $X2=6.83 $Y2=3.33
r140 34 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.77 $Y=3.245
+ $X2=7.77 $Y2=3.33
r141 34 36 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=7.77 $Y=3.245
+ $X2=7.77 $Y2=2.455
r142 30 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.83 $Y=3.245
+ $X2=6.83 $Y2=3.33
r143 30 32 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=6.83 $Y=3.245
+ $X2=6.83 $Y2=2.455
r144 26 77 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.01 $Y=3.245
+ $X2=6.01 $Y2=3.33
r145 26 28 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=6.01 $Y=3.245
+ $X2=6.01 $Y2=2.455
r146 22 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.07 $Y=3.245
+ $X2=5.07 $Y2=3.33
r147 22 24 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=5.07 $Y=3.245
+ $X2=5.07 $Y2=2.455
r148 21 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.705 $Y=3.33
+ $X2=1.58 $Y2=3.33
r149 20 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.985 $Y=3.33
+ $X2=5.07 $Y2=3.33
r150 20 21 213.989 $w=1.68e-07 $l=3.28e-06 $layer=LI1_cond $X=4.985 $Y=3.33
+ $X2=1.705 $Y2=3.33
r151 16 71 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=3.245
+ $X2=1.58 $Y2=3.33
r152 16 18 35.4952 $w=2.48e-07 $l=7.7e-07 $layer=LI1_cond $X=1.58 $Y=3.245
+ $X2=1.58 $Y2=2.475
r153 5 36 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=7.635
+ $Y=1.84 $X2=7.77 $Y2=2.455
r154 4 32 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=6.735
+ $Y=1.84 $X2=6.87 $Y2=2.455
r155 3 28 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=5.835
+ $Y=1.84 $X2=5.97 $Y2=2.455
r156 2 24 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=4.935
+ $Y=1.84 $X2=5.07 $Y2=2.455
r157 1 18 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.96 $X2=1.62 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_4%A_539_368# 1 2 3 4 5 6 7 24 28 29 32 34 36
+ 39 40 44 46 50 52 56 58 60 62 64 68 70 72
c117 70 0 1.52151e-19 $X=6.42 $Y=1.985
r118 60 74 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.22 $Y=2.12 $X2=8.22
+ $Y2=2.035
r119 60 62 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=8.22 $Y=2.12
+ $X2=8.22 $Y2=2.815
r120 59 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.485 $Y=2.035
+ $X2=7.32 $Y2=2.035
r121 58 74 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.055 $Y=2.035
+ $X2=8.22 $Y2=2.035
r122 58 59 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.055 $Y=2.035
+ $X2=7.485 $Y2=2.035
r123 54 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.32 $Y=2.12
+ $X2=7.32 $Y2=2.035
r124 54 56 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=7.32 $Y=2.12
+ $X2=7.32 $Y2=2.815
r125 53 70 5.16603 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=6.505 $Y=2.035
+ $X2=6.42 $Y2=1.97
r126 52 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.155 $Y=2.035
+ $X2=7.32 $Y2=2.035
r127 52 53 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=7.155 $Y=2.035
+ $X2=6.505 $Y2=2.035
r128 48 70 1.34256 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.42 $Y=2.12
+ $X2=6.42 $Y2=1.97
r129 48 50 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=6.42 $Y=2.12
+ $X2=6.42 $Y2=2.4
r130 47 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.685 $Y=2.035
+ $X2=5.52 $Y2=2.035
r131 46 70 5.16603 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=6.335 $Y=2.035
+ $X2=6.42 $Y2=1.97
r132 46 47 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.335 $Y=2.035
+ $X2=5.685 $Y2=2.035
r133 42 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.52 $Y=2.12
+ $X2=5.52 $Y2=2.035
r134 42 44 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.52 $Y=2.12
+ $X2=5.52 $Y2=2.815
r135 41 66 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.785 $Y=2.035
+ $X2=4.62 $Y2=2.035
r136 40 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.355 $Y=2.035
+ $X2=5.52 $Y2=2.035
r137 40 41 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.355 $Y=2.035
+ $X2=4.785 $Y2=2.035
r138 37 39 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.62 $Y=2.905
+ $X2=4.62 $Y2=2.815
r139 36 66 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.62 $Y=2.12 $X2=4.62
+ $Y2=2.035
r140 36 39 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.62 $Y=2.12
+ $X2=4.62 $Y2=2.815
r141 35 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=2.99
+ $X2=3.72 $Y2=2.99
r142 34 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.455 $Y=2.99
+ $X2=4.62 $Y2=2.905
r143 34 35 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.455 $Y=2.99
+ $X2=3.885 $Y2=2.99
r144 30 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=2.905
+ $X2=3.72 $Y2=2.99
r145 30 32 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.72 $Y=2.905
+ $X2=3.72 $Y2=2.225
r146 28 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=2.99
+ $X2=3.72 $Y2=2.99
r147 28 29 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.555 $Y=2.99
+ $X2=2.985 $Y2=2.99
r148 24 27 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.82 $Y=1.985
+ $X2=2.82 $Y2=2.815
r149 22 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.82 $Y=2.905
+ $X2=2.985 $Y2=2.99
r150 22 27 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.82 $Y=2.905
+ $X2=2.82 $Y2=2.815
r151 7 74 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=8.085
+ $Y=1.84 $X2=8.22 $Y2=2.115
r152 7 62 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.085
+ $Y=1.84 $X2=8.22 $Y2=2.815
r153 6 72 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=7.185
+ $Y=1.84 $X2=7.32 $Y2=2.115
r154 6 56 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.185
+ $Y=1.84 $X2=7.32 $Y2=2.815
r155 5 70 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.285
+ $Y=1.84 $X2=6.42 $Y2=1.985
r156 5 50 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=6.285
+ $Y=1.84 $X2=6.42 $Y2=2.4
r157 4 68 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=5.385
+ $Y=1.84 $X2=5.52 $Y2=2.115
r158 4 44 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.385
+ $Y=1.84 $X2=5.52 $Y2=2.815
r159 3 66 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=4.485
+ $Y=1.84 $X2=4.62 $Y2=2.115
r160 3 39 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.485
+ $Y=1.84 $X2=4.62 $Y2=2.815
r161 2 32 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=3.585
+ $Y=1.84 $X2=3.72 $Y2=2.225
r162 1 27 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=2.695
+ $Y=1.84 $X2=2.82 $Y2=2.815
r163 1 24 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.695
+ $Y=1.84 $X2=2.82 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_4%Y 1 2 3 4 5 6 19 21 23 27 31 33 34 35 39
+ 43 45 50 52 55 56 57
c86 45 0 4.29123e-20 $X=5.985 $Y=0.95
c87 31 0 2.7959e-19 $X=3.295 $Y=0.515
c88 21 0 3.44467e-19 $X=2.435 $Y=0.515
c89 19 0 1.64164e-19 $X=2.395 $Y=0.79
r90 57 60 6.557 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=4.11 $Y=1.295
+ $X2=4.11 $Y2=1.13
r91 56 60 0.883768 $w=2.9e-07 $l=1.7e-07 $layer=LI1_cond $X=4.11 $Y=0.96
+ $X2=4.11 $Y2=1.13
r92 54 55 5.33064 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=0.95
+ $X2=4.96 $Y2=0.95
r93 51 57 16.8893 $w=2.88e-07 $l=4.25e-07 $layer=LI1_cond $X=4.11 $Y=1.72
+ $X2=4.11 $Y2=1.295
r94 51 52 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=1.72 $X2=4.11
+ $Y2=1.805
r95 43 54 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=5.14 $Y=0.95
+ $X2=5.125 $Y2=0.95
r96 43 45 27.0504 $w=3.58e-07 $l=8.45e-07 $layer=LI1_cond $X=5.14 $Y=0.95
+ $X2=5.985 $Y2=0.95
r97 42 56 5.74179 $w=2.55e-07 $l=1.45e-07 $layer=LI1_cond $X=4.255 $Y=0.96
+ $X2=4.11 $Y2=0.96
r98 42 55 23.8962 $w=3.38e-07 $l=7.05e-07 $layer=LI1_cond $X=4.255 $Y=0.96
+ $X2=4.96 $Y2=0.96
r99 37 52 3.98977 $w=2.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=4.17 $Y=1.89
+ $X2=4.11 $Y2=1.805
r100 37 39 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=4.17 $Y=1.89
+ $X2=4.17 $Y2=1.985
r101 36 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.38 $Y=0.875
+ $X2=3.295 $Y2=0.875
r102 35 56 5.74179 $w=2.55e-07 $l=1.8262e-07 $layer=LI1_cond $X=3.965 $Y=0.875
+ $X2=4.11 $Y2=0.96
r103 35 36 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.965 $Y=0.875
+ $X2=3.38 $Y2=0.875
r104 33 52 2.45049 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.965 $Y=1.805
+ $X2=4.11 $Y2=1.805
r105 33 34 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.965 $Y=1.805
+ $X2=3.355 $Y2=1.805
r106 29 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.295 $Y=0.79
+ $X2=3.295 $Y2=0.875
r107 29 31 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.295 $Y=0.79
+ $X2=3.295 $Y2=0.515
r108 25 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.27 $Y=1.89
+ $X2=3.355 $Y2=1.805
r109 25 27 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.27 $Y=1.89
+ $X2=3.27 $Y2=1.985
r110 24 48 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.52 $Y=0.875
+ $X2=2.395 $Y2=0.875
r111 23 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.21 $Y=0.875
+ $X2=3.295 $Y2=0.875
r112 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.21 $Y=0.875
+ $X2=2.52 $Y2=0.875
r113 19 48 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.395 $Y=0.79
+ $X2=2.395 $Y2=0.875
r114 19 21 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=2.395 $Y=0.79
+ $X2=2.395 $Y2=0.515
r115 6 39 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=4.035
+ $Y=1.84 $X2=4.17 $Y2=1.985
r116 5 27 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.135
+ $Y=1.84 $X2=3.27 $Y2=1.985
r117 4 45 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=5.845
+ $Y=0.37 $X2=5.985 $Y2=0.95
r118 3 54 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=4.985
+ $Y=0.37 $X2=5.125 $Y2=0.95
r119 2 50 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=3.155
+ $Y=0.37 $X2=3.295 $Y2=0.875
r120 2 31 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.155
+ $Y=0.37 $X2=3.295 $Y2=0.515
r121 1 48 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=2.295
+ $Y=0.37 $X2=2.435 $Y2=0.875
r122 1 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.295
+ $Y=0.37 $X2=2.435 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_4%VGND 1 2 3 4 5 6 21 25 29 31 35 39 43 46
+ 47 49 50 51 52 54 55 57 58 59 82 83 86
r111 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r112 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r113 80 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=8.4
+ $Y2=0
r114 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r115 77 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r116 76 77 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r117 74 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r118 73 76 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6.48
+ $Y2=0
r119 73 74 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r120 71 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.89 $Y=0 $X2=3.725
+ $Y2=0
r121 71 73 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.89 $Y=0 $X2=4.08
+ $Y2=0
r122 70 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r123 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r124 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r125 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r126 63 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r127 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r128 59 77 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=6.48 $Y2=0
r129 59 74 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.08 $Y2=0
r130 57 79 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=7.54 $Y=0 $X2=7.44
+ $Y2=0
r131 57 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.54 $Y=0 $X2=7.665
+ $Y2=0
r132 56 82 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.79 $Y=0 $X2=8.4
+ $Y2=0
r133 56 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.79 $Y=0 $X2=7.665
+ $Y2=0
r134 54 76 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=6.68 $Y=0 $X2=6.48
+ $Y2=0
r135 54 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.68 $Y=0 $X2=6.805
+ $Y2=0
r136 53 79 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.93 $Y=0 $X2=7.44
+ $Y2=0
r137 53 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.93 $Y=0 $X2=6.805
+ $Y2=0
r138 51 69 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=2.7 $Y=0 $X2=2.64
+ $Y2=0
r139 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.7 $Y=0 $X2=2.865
+ $Y2=0
r140 49 66 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.8 $Y=0 $X2=1.68
+ $Y2=0
r141 49 50 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.8 $Y=0 $X2=1.945
+ $Y2=0
r142 48 69 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.09 $Y=0 $X2=2.64
+ $Y2=0
r143 48 50 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=2.09 $Y=0 $X2=1.945
+ $Y2=0
r144 46 62 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.94 $Y=0 $X2=0.72
+ $Y2=0
r145 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.94 $Y=0 $X2=1.105
+ $Y2=0
r146 45 66 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.27 $Y=0 $X2=1.68
+ $Y2=0
r147 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.27 $Y=0 $X2=1.105
+ $Y2=0
r148 41 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.665 $Y=0.085
+ $X2=7.665 $Y2=0
r149 41 43 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=7.665 $Y=0.085
+ $X2=7.665 $Y2=0.675
r150 37 55 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.805 $Y=0.085
+ $X2=6.805 $Y2=0
r151 37 39 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=6.805 $Y=0.085
+ $X2=6.805 $Y2=0.675
r152 33 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.725 $Y=0.085
+ $X2=3.725 $Y2=0
r153 33 35 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.725 $Y=0.085
+ $X2=3.725 $Y2=0.525
r154 32 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.03 $Y=0 $X2=2.865
+ $Y2=0
r155 31 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.56 $Y=0 $X2=3.725
+ $Y2=0
r156 31 32 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.56 $Y=0 $X2=3.03
+ $Y2=0
r157 27 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=0.085
+ $X2=2.865 $Y2=0
r158 27 29 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=2.865 $Y=0.085
+ $X2=2.865 $Y2=0.525
r159 23 50 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.945 $Y=0.085
+ $X2=1.945 $Y2=0
r160 23 25 25.2345 $w=2.88e-07 $l=6.35e-07 $layer=LI1_cond $X=1.945 $Y=0.085
+ $X2=1.945 $Y2=0.72
r161 19 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.105 $Y=0.085
+ $X2=1.105 $Y2=0
r162 19 21 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=1.105 $Y=0.085
+ $X2=1.105 $Y2=0.525
r163 6 43 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=7.565
+ $Y=0.37 $X2=7.705 $Y2=0.675
r164 5 39 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=6.705
+ $Y=0.37 $X2=6.845 $Y2=0.675
r165 4 35 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.37 $X2=3.725 $Y2=0.525
r166 3 29 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=2.725
+ $Y=0.37 $X2=2.865 $Y2=0.525
r167 2 25 182 $w=1.7e-07 $l=4.22493e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.37 $X2=1.985 $Y2=0.72
r168 1 21 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.37 $X2=1.105 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_4%A_914_74# 1 2 3 4 5 16 22 26 27 30 32 36
+ 40
c54 26 0 1.52151e-19 $X=7.11 $Y=1.095
c55 22 0 1.6164e-19 $X=6.415 $Y=0.6
r56 34 36 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=8.135 $Y=1.01
+ $X2=8.135 $Y2=0.515
r57 33 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.36 $Y=1.095
+ $X2=7.235 $Y2=1.095
r58 32 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.97 $Y=1.095
+ $X2=8.135 $Y2=1.01
r59 32 33 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.97 $Y=1.095
+ $X2=7.36 $Y2=1.095
r60 28 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.235 $Y=1.01
+ $X2=7.235 $Y2=1.095
r61 28 30 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=7.235 $Y=1.01
+ $X2=7.235 $Y2=0.515
r62 26 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.11 $Y=1.095
+ $X2=7.235 $Y2=1.095
r63 26 27 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.11 $Y=1.095
+ $X2=6.5 $Y2=1.095
r64 23 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.415 $Y=1.01
+ $X2=6.5 $Y2=1.095
r65 23 25 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=6.415 $Y=1.01
+ $X2=6.415 $Y2=0.965
r66 22 39 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.415 $Y=0.6
+ $X2=6.415 $Y2=0.475
r67 22 25 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.415 $Y=0.6
+ $X2=6.415 $Y2=0.965
r68 18 21 39.644 $w=2.48e-07 $l=8.6e-07 $layer=LI1_cond $X=4.695 $Y=0.475
+ $X2=5.555 $Y2=0.475
r69 16 39 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.33 $Y=0.475
+ $X2=6.415 $Y2=0.475
r70 16 21 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=6.33 $Y=0.475
+ $X2=5.555 $Y2=0.475
r71 5 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.995
+ $Y=0.37 $X2=8.135 $Y2=0.515
r72 4 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.135
+ $Y=0.37 $X2=7.275 $Y2=0.515
r73 3 39 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.275
+ $Y=0.37 $X2=6.415 $Y2=0.515
r74 3 25 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=6.275
+ $Y=0.37 $X2=6.415 $Y2=0.965
r75 2 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.415
+ $Y=0.37 $X2=5.555 $Y2=0.515
r76 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.57
+ $Y=0.37 $X2=4.695 $Y2=0.515
.ends


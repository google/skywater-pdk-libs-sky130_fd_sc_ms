* File: sky130_fd_sc_ms__mux4_1.spice
* Created: Fri Aug 28 17:40:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__mux4_1.pex.spice"
.subckt sky130_fd_sc_ms__mux4_1  VNB VPB A0 A1 A2 S0 A3 S1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* S1	S1
* A3	A3
* S0	S0
* A2	A2
* A1	A1
* A0	A0
* VPB	VPB
* VNB	VNB
MM1021 N_VGND_M1021_d N_S0_M1021_g N_A_27_74#_M1021_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.192 AS=0.1824 PD=1.24 PS=1.85 NRD=34.68 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75004.9 A=0.096 P=1.58 MULT=1
MM1014 A_264_74# N_A0_M1014_g N_VGND_M1021_d VNB NLOWVT L=0.15 W=0.64 AD=0.0768
+ AS=0.192 PD=0.88 PS=1.24 NRD=12.18 NRS=25.308 M=1 R=4.26667 SA=75001
+ SB=75004.2 A=0.096 P=1.58 MULT=1
MM1015 N_A_342_74#_M1015_d N_A_27_74#_M1015_g A_264_74# VNB NLOWVT L=0.15 W=0.64
+ AD=0.1248 AS=0.0768 PD=1.03 PS=0.88 NRD=20.616 NRS=12.18 M=1 R=4.26667
+ SA=75001.3 SB=75003.8 A=0.096 P=1.58 MULT=1
MM1019 A_450_74# N_S0_M1019_g N_A_342_74#_M1015_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.24 AS=0.1248 PD=1.39 PS=1.03 NRD=60 NRS=0 M=1 R=4.26667 SA=75001.9
+ SB=75003.2 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1001_d N_A1_M1001_g A_450_74# VNB NLOWVT L=0.15 W=0.64 AD=0.1728
+ AS=0.24 PD=1.18 PS=1.39 NRD=24.372 NRS=60 M=1 R=4.26667 SA=75002.8 SB=75002.3
+ A=0.096 P=1.58 MULT=1
MM1023 A_768_74# N_A2_M1023_g N_VGND_M1001_d VNB NLOWVT L=0.15 W=0.64 AD=0.0768
+ AS=0.1728 PD=0.88 PS=1.18 NRD=12.18 NRS=24.372 M=1 R=4.26667 SA=75003.5
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1022 N_A_846_74#_M1022_d N_A_27_74#_M1022_g A_768_74# VNB NLOWVT L=0.15 W=0.64
+ AD=0.1648 AS=0.0768 PD=1.155 PS=0.88 NRD=21.552 NRS=12.18 M=1 R=4.26667
+ SA=75003.9 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1003 A_979_74# N_S0_M1003_g N_A_846_74#_M1022_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1648 PD=0.88 PS=1.155 NRD=12.18 NRS=22.488 M=1 R=4.26667
+ SA=75004.5 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1025 N_VGND_M1025_d N_A3_M1025_g A_979_74# VNB NLOWVT L=0.15 W=0.64 AD=0.1824
+ AS=0.0768 PD=1.85 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667 SA=75004.9 SB=75000.2
+ A=0.096 P=1.58 MULT=1
MM1004 N_A_1338_125#_M1004_d N_S1_M1004_g N_A_846_74#_M1004_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0928 AS=0.454475 PD=0.93 PS=3.19 NRD=0.936 NRS=46.872 M=1
+ R=4.26667 SA=75000.3 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1024 N_A_342_74#_M1024_d N_A_1396_99#_M1024_g N_A_1338_125#_M1004_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.0928 PD=1.85 PS=0.93 NRD=0 NRS=0.936 M=1
+ R=4.26667 SA=75000.8 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1011 N_VGND_M1011_d N_S1_M1011_g N_A_1396_99#_M1011_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.136255 AS=0.1824 PD=1.07594 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1017 N_X_M1017_d N_A_1338_125#_M1017_g N_VGND_M1011_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.157545 PD=2.05 PS=1.24406 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_VPWR_M1009_d N_S0_M1009_g N_A_27_74#_M1009_s VPB PSHORT L=0.18 W=1
+ AD=0.214312 AS=0.28 PD=1.54 PS=2.56 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90004.4 A=0.18 P=2.36 MULT=1
MM1020 A_258_341# N_A0_M1020_g N_VPWR_M1009_d VPB PSHORT L=0.18 W=1 AD=0.39
+ AS=0.214312 PD=1.78 PS=1.54 NRD=65.9753 NRS=16.0752 M=1 R=5.55556 SA=90000.7
+ SB=90004.2 A=0.18 P=2.36 MULT=1
MM1010 N_A_342_74#_M1010_d N_S0_M1010_g A_258_341# VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.39 PD=1.27 PS=1.78 NRD=0 NRS=65.9753 M=1 R=5.55556 SA=90001.7
+ SB=90003.2 A=0.18 P=2.36 MULT=1
MM1013 A_540_341# N_A_27_74#_M1013_g N_A_342_74#_M1010_d VPB PSHORT L=0.18 W=1
+ AD=0.165 AS=0.135 PD=1.33 PS=1.27 NRD=21.6503 NRS=0 M=1 R=5.55556 SA=90002.1
+ SB=90002.8 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g A_540_341# VPB PSHORT L=0.18 W=1 AD=0.2606
+ AS=0.165 PD=1.72 PS=1.33 NRD=40.4835 NRS=21.6503 M=1 R=5.55556 SA=90002.6
+ SB=90002.3 A=0.18 P=2.36 MULT=1
MM1002 A_766_341# N_A2_M1002_g N_VPWR_M1000_d VPB PSHORT L=0.18 W=1 AD=0.182625
+ AS=0.2606 PD=1.555 PS=1.72 NRD=25.1372 NRS=40.4835 M=1 R=5.55556 SA=90003.2
+ SB=90001.7 A=0.18 P=2.36 MULT=1
MM1008 N_A_846_74#_M1008_d N_S0_M1008_g A_766_341# VPB PSHORT L=0.18 W=1
+ AD=0.4125 AS=0.182625 PD=1.825 PS=1.555 NRD=0 NRS=25.1372 M=1 R=5.55556
+ SA=90003 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1005 A_1068_387# N_A_27_74#_M1005_g N_A_846_74#_M1008_d VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.4125 PD=1.24 PS=1.825 NRD=12.7853 NRS=0 M=1 R=5.55556 SA=90004
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_A3_M1012_g A_1068_387# VPB PSHORT L=0.18 W=1 AD=0.28
+ AS=0.12 PD=2.56 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556 SA=90004.4 SB=90000.2
+ A=0.18 P=2.36 MULT=1
MM1007 N_A_1338_125#_M1007_d N_S1_M1007_g N_A_342_74#_M1007_s VPB PSHORT L=0.18
+ W=1 AD=0.16 AS=0.28 PD=1.32 PS=2.56 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1006 N_A_846_74#_M1006_d N_A_1396_99#_M1006_g N_A_1338_125#_M1007_d VPB PSHORT
+ L=0.18 W=1 AD=0.33 AS=0.16 PD=2.66 PS=1.32 NRD=8.8453 NRS=0 M=1 R=5.55556
+ SA=90000.7 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1016 N_VPWR_M1016_d N_S1_M1016_g N_A_1396_99#_M1016_s VPB PSHORT L=0.18 W=1
+ AD=0.302241 AS=0.33 PD=1.63208 PS=2.66 NRD=65.995 NRS=8.8453 M=1 R=5.55556
+ SA=90000.2 SB=90001 A=0.18 P=2.36 MULT=1
MM1018 N_X_M1018_d N_A_1338_125#_M1018_g N_VPWR_M1016_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3304 AS=0.338509 PD=2.83 PS=1.82792 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.9
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX26_noxref VNB VPB NWDIODE A=19.0461 P=23.95
c_182 VPB 0 1.25754e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__mux4_1.pxi.spice"
*
.ends
*
*

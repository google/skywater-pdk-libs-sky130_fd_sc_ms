* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
M1000 a_225_82# C VPWR VPB pshort w=1e+06u l=180000u
+  ad=8.1e+11p pd=5.62e+06u as=1.854e+12p ps=1.212e+07u
M1001 VPWR D a_225_82# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_390_82# a_354_252# a_312_82# VNB nlowvt w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=1.776e+11p ps=1.96e+06u
M1003 X a_225_82# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=1.0454e+12p ps=7.35e+06u
M1004 a_312_82# a_27_74# a_225_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1005 a_354_252# B_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.478e+11p pd=2.27e+06u as=0p ps=0u
M1006 a_354_252# B_N VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1007 VGND a_225_82# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_225_82# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1009 VPWR a_225_82# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_498_82# C a_390_82# VNB nlowvt w=740000u l=150000u
+  ad=2.664e+11p pd=2.2e+06u as=0p ps=0u
M1011 VGND D a_498_82# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_354_252# a_225_82# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_225_82# a_27_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A_N a_27_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1015 VPWR A_N a_27_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
.ends

* File: sky130_fd_sc_ms__sdfxtp_1.pxi.spice
* Created: Fri Aug 28 18:14:25 2020
* 
x_PM_SKY130_FD_SC_MS__SDFXTP_1%A_35_74# N_A_35_74#_M1006_s N_A_35_74#_M1014_s
+ N_A_35_74#_M1020_g N_A_35_74#_M1027_g N_A_35_74#_c_234_n N_A_35_74#_c_227_n
+ N_A_35_74#_c_235_n N_A_35_74#_c_236_n N_A_35_74#_c_228_n N_A_35_74#_c_229_n
+ N_A_35_74#_c_230_n N_A_35_74#_c_231_n N_A_35_74#_c_232_n
+ PM_SKY130_FD_SC_MS__SDFXTP_1%A_35_74#
x_PM_SKY130_FD_SC_MS__SDFXTP_1%SCE N_SCE_c_321_n N_SCE_c_322_n N_SCE_c_323_n
+ N_SCE_c_332_n N_SCE_c_333_n N_SCE_M1006_g N_SCE_c_334_n N_SCE_M1014_g
+ N_SCE_c_335_n N_SCE_c_336_n N_SCE_M1012_g N_SCE_M1029_g N_SCE_c_337_n
+ N_SCE_c_325_n N_SCE_c_326_n N_SCE_c_327_n SCE N_SCE_c_328_n N_SCE_c_329_n
+ N_SCE_c_330_n PM_SKY130_FD_SC_MS__SDFXTP_1%SCE
x_PM_SKY130_FD_SC_MS__SDFXTP_1%D N_D_M1021_g N_D_M1025_g D N_D_c_409_n
+ N_D_c_410_n PM_SKY130_FD_SC_MS__SDFXTP_1%D
x_PM_SKY130_FD_SC_MS__SDFXTP_1%SCD N_SCD_M1002_g N_SCD_M1028_g N_SCD_c_448_n
+ N_SCD_c_453_n SCD N_SCD_c_450_n PM_SKY130_FD_SC_MS__SDFXTP_1%SCD
x_PM_SKY130_FD_SC_MS__SDFXTP_1%CLK N_CLK_c_493_n N_CLK_M1003_g N_CLK_M1004_g CLK
+ N_CLK_c_496_n PM_SKY130_FD_SC_MS__SDFXTP_1%CLK
x_PM_SKY130_FD_SC_MS__SDFXTP_1%A_828_74# N_A_828_74#_M1018_d N_A_828_74#_M1008_d
+ N_A_828_74#_M1015_g N_A_828_74#_c_536_n N_A_828_74#_M1030_g
+ N_A_828_74#_M1000_g N_A_828_74#_M1010_g N_A_828_74#_c_556_n
+ N_A_828_74#_c_537_n N_A_828_74#_c_538_n N_A_828_74#_c_539_n
+ N_A_828_74#_c_540_n N_A_828_74#_c_541_n N_A_828_74#_c_542_n
+ N_A_828_74#_c_543_n N_A_828_74#_c_544_n N_A_828_74#_c_614_p
+ N_A_828_74#_c_630_p N_A_828_74#_c_545_n N_A_828_74#_c_546_n
+ N_A_828_74#_c_547_n N_A_828_74#_c_558_n N_A_828_74#_c_548_n
+ N_A_828_74#_c_560_n N_A_828_74#_c_561_n N_A_828_74#_c_549_n
+ N_A_828_74#_c_715_p N_A_828_74#_c_550_n N_A_828_74#_c_551_n
+ N_A_828_74#_c_552_n N_A_828_74#_c_553_n PM_SKY130_FD_SC_MS__SDFXTP_1%A_828_74#
x_PM_SKY130_FD_SC_MS__SDFXTP_1%A_630_74# N_A_630_74#_M1003_d N_A_630_74#_M1004_d
+ N_A_630_74#_M1018_g N_A_630_74#_c_734_n N_A_630_74#_M1008_g
+ N_A_630_74#_c_736_n N_A_630_74#_M1007_g N_A_630_74#_c_753_n
+ N_A_630_74#_M1013_g N_A_630_74#_M1026_g N_A_630_74#_c_738_n
+ N_A_630_74#_c_739_n N_A_630_74#_c_740_n N_A_630_74#_c_741_n
+ N_A_630_74#_M1023_g N_A_630_74#_c_742_n N_A_630_74#_c_743_n
+ N_A_630_74#_c_744_n N_A_630_74#_c_757_n N_A_630_74#_c_745_n
+ N_A_630_74#_c_746_n N_A_630_74#_c_779_n N_A_630_74#_c_747_n
+ N_A_630_74#_c_748_n N_A_630_74#_c_759_n N_A_630_74#_c_760_n
+ N_A_630_74#_c_867_p N_A_630_74#_c_761_n N_A_630_74#_c_749_n
+ N_A_630_74#_c_762_n N_A_630_74#_c_763_n N_A_630_74#_c_750_n
+ N_A_630_74#_c_751_n N_A_630_74#_c_766_n PM_SKY130_FD_SC_MS__SDFXTP_1%A_630_74#
x_PM_SKY130_FD_SC_MS__SDFXTP_1%A_1239_74# N_A_1239_74#_M1011_d
+ N_A_1239_74#_M1016_d N_A_1239_74#_M1024_g N_A_1239_74#_c_952_n
+ N_A_1239_74#_M1019_g N_A_1239_74#_c_945_n N_A_1239_74#_c_946_n
+ N_A_1239_74#_c_947_n N_A_1239_74#_c_948_n N_A_1239_74#_c_955_n
+ N_A_1239_74#_c_949_n N_A_1239_74#_c_967_n N_A_1239_74#_c_950_n
+ N_A_1239_74#_c_951_n PM_SKY130_FD_SC_MS__SDFXTP_1%A_1239_74#
x_PM_SKY130_FD_SC_MS__SDFXTP_1%A_1018_100# N_A_1018_100#_M1007_d
+ N_A_1018_100#_M1015_d N_A_1018_100#_M1016_g N_A_1018_100#_M1011_g
+ N_A_1018_100#_c_1023_n N_A_1018_100#_c_1029_n N_A_1018_100#_c_1024_n
+ N_A_1018_100#_c_1025_n N_A_1018_100#_c_1031_n N_A_1018_100#_c_1032_n
+ N_A_1018_100#_c_1026_n N_A_1018_100#_c_1027_n
+ PM_SKY130_FD_SC_MS__SDFXTP_1%A_1018_100#
x_PM_SKY130_FD_SC_MS__SDFXTP_1%A_1736_74# N_A_1736_74#_M1009_d
+ N_A_1736_74#_M1031_d N_A_1736_74#_c_1112_n N_A_1736_74#_M1005_g
+ N_A_1736_74#_c_1122_n N_A_1736_74#_M1022_g N_A_1736_74#_c_1113_n
+ N_A_1736_74#_M1001_g N_A_1736_74#_M1017_g N_A_1736_74#_c_1125_n
+ N_A_1736_74#_c_1116_n N_A_1736_74#_c_1117_n N_A_1736_74#_c_1118_n
+ N_A_1736_74#_c_1119_n N_A_1736_74#_c_1120_n N_A_1736_74#_c_1126_n
+ N_A_1736_74#_c_1127_n N_A_1736_74#_c_1121_n
+ PM_SKY130_FD_SC_MS__SDFXTP_1%A_1736_74#
x_PM_SKY130_FD_SC_MS__SDFXTP_1%A_1520_74# N_A_1520_74#_M1000_d
+ N_A_1520_74#_M1026_d N_A_1520_74#_M1031_g N_A_1520_74#_M1009_g
+ N_A_1520_74#_c_1205_n N_A_1520_74#_c_1206_n N_A_1520_74#_c_1207_n
+ N_A_1520_74#_c_1199_n N_A_1520_74#_c_1208_n N_A_1520_74#_c_1200_n
+ N_A_1520_74#_c_1201_n N_A_1520_74#_c_1202_n N_A_1520_74#_c_1203_n
+ PM_SKY130_FD_SC_MS__SDFXTP_1%A_1520_74#
x_PM_SKY130_FD_SC_MS__SDFXTP_1%VPWR N_VPWR_M1014_d N_VPWR_M1002_d N_VPWR_M1008_s
+ N_VPWR_M1019_d N_VPWR_M1022_d N_VPWR_M1001_s N_VPWR_c_1288_n N_VPWR_c_1289_n
+ N_VPWR_c_1290_n N_VPWR_c_1291_n N_VPWR_c_1292_n N_VPWR_c_1293_n
+ N_VPWR_c_1294_n N_VPWR_c_1295_n N_VPWR_c_1296_n N_VPWR_c_1297_n
+ N_VPWR_c_1298_n N_VPWR_c_1299_n VPWR N_VPWR_c_1300_n N_VPWR_c_1301_n
+ N_VPWR_c_1302_n N_VPWR_c_1303_n N_VPWR_c_1287_n N_VPWR_c_1305_n
+ N_VPWR_c_1306_n N_VPWR_c_1307_n PM_SKY130_FD_SC_MS__SDFXTP_1%VPWR
x_PM_SKY130_FD_SC_MS__SDFXTP_1%A_301_74# N_A_301_74#_M1021_d N_A_301_74#_M1007_s
+ N_A_301_74#_M1025_d N_A_301_74#_M1015_s N_A_301_74#_c_1422_n
+ N_A_301_74#_c_1415_n N_A_301_74#_c_1407_n N_A_301_74#_c_1408_n
+ N_A_301_74#_c_1409_n N_A_301_74#_c_1410_n N_A_301_74#_c_1462_n
+ N_A_301_74#_c_1417_n N_A_301_74#_c_1411_n N_A_301_74#_c_1412_n
+ N_A_301_74#_c_1470_n N_A_301_74#_c_1413_n N_A_301_74#_c_1418_n
+ N_A_301_74#_c_1419_n N_A_301_74#_c_1420_n N_A_301_74#_c_1527_n
+ N_A_301_74#_c_1421_n N_A_301_74#_c_1414_n
+ PM_SKY130_FD_SC_MS__SDFXTP_1%A_301_74#
x_PM_SKY130_FD_SC_MS__SDFXTP_1%Q N_Q_M1017_d N_Q_M1001_d Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_MS__SDFXTP_1%Q
x_PM_SKY130_FD_SC_MS__SDFXTP_1%VGND N_VGND_M1006_d N_VGND_M1028_d N_VGND_M1018_s
+ N_VGND_M1024_d N_VGND_M1005_d N_VGND_M1017_s N_VGND_c_1556_n N_VGND_c_1557_n
+ N_VGND_c_1558_n N_VGND_c_1559_n N_VGND_c_1560_n N_VGND_c_1561_n
+ N_VGND_c_1562_n N_VGND_c_1563_n N_VGND_c_1564_n N_VGND_c_1565_n VGND
+ N_VGND_c_1566_n N_VGND_c_1567_n N_VGND_c_1568_n N_VGND_c_1569_n
+ N_VGND_c_1570_n N_VGND_c_1571_n N_VGND_c_1572_n N_VGND_c_1573_n
+ N_VGND_c_1574_n N_VGND_c_1575_n PM_SKY130_FD_SC_MS__SDFXTP_1%VGND
cc_1 VNB N_A_35_74#_M1020_g 0.0493688f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.58
cc_2 VNB N_A_35_74#_c_227_n 0.029403f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=1.525
cc_3 VNB N_A_35_74#_c_228_n 0.00230899f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.635
cc_4 VNB N_A_35_74#_c_229_n 0.0176748f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.635
cc_5 VNB N_A_35_74#_c_230_n 0.0207287f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=0.565
cc_6 VNB N_A_35_74#_c_231_n 0.0214782f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.69
cc_7 VNB N_A_35_74#_c_232_n 0.00801772f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=1.825
cc_8 VNB N_SCE_c_321_n 0.0229485f $X=-0.19 $Y=-0.245 $X2=0.245 $Y2=2.32
cc_9 VNB N_SCE_c_322_n 0.0112516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_SCE_c_323_n 0.010922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_SCE_M1006_g 0.0245768f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.58
cc_12 VNB N_SCE_c_325_n 0.031826f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.635
cc_13 VNB N_SCE_c_326_n 0.0175089f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=0.567
cc_14 VNB N_SCE_c_327_n 0.0303895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_SCE_c_328_n 0.0199759f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.69
cc_16 VNB N_SCE_c_329_n 0.00701215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_SCE_c_330_n 0.00651353f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.525
cc_18 VNB N_D_M1021_g 0.0517631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_D_c_409_n 0.0161794f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=2.64
cc_20 VNB N_D_c_410_n 0.00377665f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=2.64
cc_21 VNB N_SCD_M1028_g 0.0524176f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.525
cc_22 VNB N_SCD_c_448_n 0.00166739f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=2.14
cc_23 VNB SCD 0.00342799f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=2.64
cc_24 VNB N_SCD_c_450_n 0.0165724f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=2.14
cc_25 VNB N_CLK_c_493_n 0.0214812f $X=-0.19 $Y=-0.245 $X2=0.175 $Y2=0.37
cc_26 VNB N_CLK_M1004_g 0.00749619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB CLK 0.00809038f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.58
cc_28 VNB N_CLK_c_496_n 0.0531476f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=2.14
cc_29 VNB N_A_828_74#_c_536_n 0.0183603f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=2.14
cc_30 VNB N_A_828_74#_c_537_n 0.00996782f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=2.04
cc_31 VNB N_A_828_74#_c_538_n 0.0164465f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.635
cc_32 VNB N_A_828_74#_c_539_n 0.00365087f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.635
cc_33 VNB N_A_828_74#_c_540_n 0.00639393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_828_74#_c_541_n 0.0174224f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=0.567
cc_35 VNB N_A_828_74#_c_542_n 6.88452e-19 $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=0.565
cc_36 VNB N_A_828_74#_c_543_n 0.00279686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_828_74#_c_544_n 0.0394958f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.825
cc_38 VNB N_A_828_74#_c_545_n 0.00869027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_828_74#_c_546_n 0.00244258f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.69
cc_40 VNB N_A_828_74#_c_547_n 0.0175834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_828_74#_c_548_n 0.0242021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_828_74#_c_549_n 0.00123754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_828_74#_c_550_n 0.0066909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_828_74#_c_551_n 0.0342754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_828_74#_c_552_n 0.00190275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_828_74#_c_553_n 0.0197728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_630_74#_M1018_g 0.0264372f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.58
cc_48 VNB N_A_630_74#_c_734_n 0.0122933f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=2.14
cc_49 VNB N_A_630_74#_M1008_g 0.00193628f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.975
cc_50 VNB N_A_630_74#_c_736_n 0.0262728f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=0.785
cc_51 VNB N_A_630_74#_M1007_g 0.0464438f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=2.465
cc_52 VNB N_A_630_74#_c_738_n 0.0258932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_630_74#_c_739_n 0.0183966f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.825
cc_54 VNB N_A_630_74#_c_740_n 0.00994721f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.825
cc_55 VNB N_A_630_74#_c_741_n 0.0176984f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.69
cc_56 VNB N_A_630_74#_c_742_n 0.00995479f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.635
cc_57 VNB N_A_630_74#_c_743_n 0.00867977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_630_74#_c_744_n 0.00761442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_630_74#_c_745_n 0.00808997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_630_74#_c_746_n 2.58108e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_630_74#_c_747_n 5.94375e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_630_74#_c_748_n 0.0400274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_630_74#_c_749_n 0.00329671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_630_74#_c_750_n 6.18184e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_630_74#_c_751_n 0.0136293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1239_74#_c_945_n 0.0235398f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=2.14
cc_67 VNB N_A_1239_74#_c_946_n 0.0122231f $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=0.785
cc_68 VNB N_A_1239_74#_c_947_n 0.0304611f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=2.465
cc_69 VNB N_A_1239_74#_c_948_n 8.08094e-19 $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=2.04
cc_70 VNB N_A_1239_74#_c_949_n 0.00383613f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.635
cc_71 VNB N_A_1239_74#_c_950_n 0.00196184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1239_74#_c_951_n 0.0208314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1018_100#_M1011_g 0.0523031f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=2.64
cc_74 VNB N_A_1018_100#_c_1023_n 0.0157486f $X=-0.19 $Y=-0.245 $X2=0.17
+ $Y2=0.785
cc_75 VNB N_A_1018_100#_c_1024_n 0.0103148f $X=-0.19 $Y=-0.245 $X2=2.03
+ $Y2=1.955
cc_76 VNB N_A_1018_100#_c_1025_n 8.56573e-19 $X=-0.19 $Y=-0.245 $X2=2.03
+ $Y2=1.635
cc_77 VNB N_A_1018_100#_c_1026_n 0.00359804f $X=-0.19 $Y=-0.245 $X2=0.17
+ $Y2=0.567
cc_78 VNB N_A_1018_100#_c_1027_n 0.0154872f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.69
cc_79 VNB N_A_1736_74#_c_1112_n 0.017257f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.525
cc_80 VNB N_A_1736_74#_c_1113_n 0.0159888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1736_74#_M1001_g 6.91195e-19 $X=-0.19 $Y=-0.245 $X2=0.17 $Y2=0.785
cc_82 VNB N_A_1736_74#_M1017_g 0.0280762f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=2.465
cc_83 VNB N_A_1736_74#_c_1116_n 0.0532604f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.635
cc_84 VNB N_A_1736_74#_c_1117_n 0.0173802f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.635
cc_85 VNB N_A_1736_74#_c_1118_n 0.00485979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1736_74#_c_1119_n 0.00913282f $X=-0.19 $Y=-0.245 $X2=0.66
+ $Y2=1.825
cc_87 VNB N_A_1736_74#_c_1120_n 0.0269789f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.69
cc_88 VNB N_A_1736_74#_c_1121_n 0.0565155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1520_74#_M1009_g 0.0533763f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=2.64
cc_90 VNB N_A_1520_74#_c_1199_n 0.00359946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1520_74#_c_1200_n 0.00184614f $X=-0.19 $Y=-0.245 $X2=2.03
+ $Y2=1.635
cc_92 VNB N_A_1520_74#_c_1201_n 0.0108024f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.635
cc_93 VNB N_A_1520_74#_c_1202_n 0.0140958f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=0.565
cc_94 VNB N_A_1520_74#_c_1203_n 3.57783e-19 $X=-0.19 $Y=-0.245 $X2=0.17
+ $Y2=1.825
cc_95 VNB N_VPWR_c_1287_n 0.462217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_301_74#_c_1407_n 0.00243276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_301_74#_c_1408_n 0.0153861f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=2.04
cc_98 VNB N_A_301_74#_c_1409_n 0.00219671f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=2.04
cc_99 VNB N_A_301_74#_c_1410_n 0.00557658f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.635
cc_100 VNB N_A_301_74#_c_1411_n 0.00388435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_301_74#_c_1412_n 0.00224253f $X=-0.19 $Y=-0.245 $X2=0.32
+ $Y2=0.567
cc_102 VNB N_A_301_74#_c_1413_n 0.0117089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_301_74#_c_1414_n 0.00658719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB Q 0.054179f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.525
cc_105 VNB N_VGND_c_1556_n 0.00655155f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=2.465
cc_106 VNB N_VGND_c_1557_n 0.00807568f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.955
cc_107 VNB N_VGND_c_1558_n 0.00939245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1559_n 0.00822673f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=0.565
cc_109 VNB N_VGND_c_1560_n 0.0173663f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.825
cc_110 VNB N_VGND_c_1561_n 0.019401f $X=-0.19 $Y=-0.245 $X2=0.825 $Y2=1.825
cc_111 VNB N_VGND_c_1562_n 0.0513128f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.69
cc_112 VNB N_VGND_c_1563_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.525
cc_113 VNB N_VGND_c_1564_n 0.0209223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1565_n 0.00613324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1566_n 0.0181062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1567_n 0.057222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1568_n 0.0565515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1569_n 0.0194903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1570_n 0.0192125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1571_n 0.606411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1572_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1573_n 0.00477982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1574_n 0.0129835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1575_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VPB N_A_35_74#_M1027_g 0.0243628f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=2.64
cc_126 VPB N_A_35_74#_c_234_n 0.0136529f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=2.14
cc_127 VPB N_A_35_74#_c_235_n 0.0404316f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=2.465
cc_128 VPB N_A_35_74#_c_236_n 0.0225459f $X=-0.19 $Y=1.66 $X2=1.865 $Y2=2.04
cc_129 VPB N_A_35_74#_c_229_n 0.0214258f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.635
cc_130 VPB N_A_35_74#_c_231_n 0.0241408f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.69
cc_131 VPB N_A_35_74#_c_232_n 0.0227388f $X=-0.19 $Y=1.66 $X2=0.825 $Y2=1.825
cc_132 VPB N_SCE_c_321_n 0.0258923f $X=-0.19 $Y=1.66 $X2=0.245 $Y2=2.32
cc_133 VPB N_SCE_c_332_n 0.0191236f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_SCE_c_333_n 0.010921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_SCE_c_334_n 0.0216639f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=2.14
cc_136 VPB N_SCE_c_335_n 0.0226181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_SCE_c_336_n 0.0166285f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=2.14
cc_138 VPB N_SCE_c_337_n 0.00494854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_D_M1025_g 0.0448062f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.525
cc_140 VPB N_D_c_409_n 0.0117982f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=2.64
cc_141 VPB N_D_c_410_n 0.00352995f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=2.64
cc_142 VPB N_SCD_M1002_g 0.0268527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_SCD_c_448_n 0.0218151f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=2.14
cc_144 VPB N_SCD_c_453_n 0.0156983f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=2.64
cc_145 VPB SCD 0.00470416f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=2.64
cc_146 VPB N_CLK_M1004_g 0.027759f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_828_74#_M1015_g 0.0276023f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=0.58
cc_148 VPB N_A_828_74#_M1010_g 0.0368783f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=2.125
cc_149 VPB N_A_828_74#_c_556_n 0.0255241f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=2.465
cc_150 VPB N_A_828_74#_c_540_n 0.00308658f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_828_74#_c_558_n 9.29659e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_828_74#_c_548_n 0.0184465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_828_74#_c_560_n 0.0144773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_828_74#_c_561_n 0.0476956f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_630_74#_M1008_g 0.0303927f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.975
cc_156 VPB N_A_630_74#_c_753_n 0.0572036f $X=-0.19 $Y=1.66 $X2=1.865 $Y2=2.04
cc_157 VPB N_A_630_74#_M1013_g 0.0317305f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_630_74#_M1026_g 0.0283715f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=0.565
cc_159 VPB N_A_630_74#_c_743_n 0.0102901f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_630_74#_c_757_n 0.0136179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_630_74#_c_747_n 0.00321728f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_630_74#_c_759_n 0.00564588f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_A_630_74#_c_760_n 0.00752343f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_630_74#_c_761_n 0.00153764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_630_74#_c_762_n 0.0143045f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_630_74#_c_763_n 0.00776005f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_A_630_74#_c_750_n 0.00377631f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_630_74#_c_751_n 0.0335981f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_630_74#_c_766_n 0.015142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_A_1239_74#_c_952_n 0.00652147f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_A_1239_74#_M1019_g 0.0216857f $X=-0.19 $Y=1.66 $X2=1.985 $Y2=2.64
cc_172 VPB N_A_1239_74#_c_945_n 0.0352247f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=2.14
cc_173 VPB N_A_1239_74#_c_955_n 0.00332302f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.635
cc_174 VPB N_A_1239_74#_c_949_n 0.00458138f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.635
cc_175 VPB N_A_1018_100#_M1016_g 0.0283338f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=0.58
cc_176 VPB N_A_1018_100#_c_1029_n 0.00274525f $X=-0.19 $Y=1.66 $X2=1.865
+ $Y2=2.04
cc_177 VPB N_A_1018_100#_c_1024_n 0.0103824f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.955
cc_178 VPB N_A_1018_100#_c_1031_n 0.00697767f $X=-0.19 $Y=1.66 $X2=2.03
+ $Y2=1.635
cc_179 VPB N_A_1018_100#_c_1032_n 0.00256207f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_1018_100#_c_1026_n 0.0035137f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=0.567
cc_181 VPB N_A_1018_100#_c_1027_n 0.0335046f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.69
cc_182 VPB N_A_1736_74#_c_1122_n 0.0182928f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_1736_74#_c_1113_n 0.0318383f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_1736_74#_M1001_g 0.0308727f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=0.785
cc_185 VPB N_A_1736_74#_c_1125_n 0.0200252f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.955
cc_186 VPB N_A_1736_74#_c_1126_n 0.0151692f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_1736_74#_c_1127_n 0.00869523f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.69
cc_188 VPB N_A_1520_74#_M1031_g 0.0283477f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=0.58
cc_189 VPB N_A_1520_74#_c_1205_n 0.00467912f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.975
cc_190 VPB N_A_1520_74#_c_1206_n 0.0039298f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=0.785
cc_191 VPB N_A_1520_74#_c_1207_n 0.0222238f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=2.125
cc_192 VPB N_A_1520_74#_c_1208_n 0.00237715f $X=-0.19 $Y=1.66 $X2=0.825 $Y2=2.04
cc_193 VPB N_A_1520_74#_c_1200_n 0.00894446f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.635
cc_194 VPB N_A_1520_74#_c_1201_n 0.0316652f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.635
cc_195 VPB N_A_1520_74#_c_1203_n 0.00161002f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=1.825
cc_196 VPB N_VPWR_c_1288_n 0.00856778f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=2.465
cc_197 VPB N_VPWR_c_1289_n 0.00841791f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.955
cc_198 VPB N_VPWR_c_1290_n 0.0128761f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1291_n 0.00771885f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=0.565
cc_200 VPB N_VPWR_c_1292_n 0.00902245f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.825
cc_201 VPB N_VPWR_c_1293_n 0.0215292f $X=-0.19 $Y=1.66 $X2=0.825 $Y2=1.825
cc_202 VPB N_VPWR_c_1294_n 0.0215455f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1295_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1296_n 0.0486086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1297_n 0.00949348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1298_n 0.0204869f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1299_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1300_n 0.0214173f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1301_n 0.0560572f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1302_n 0.0586206f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1303_n 0.019908f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1287_n 0.131435f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1305_n 0.00959004f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1306_n 0.00631473f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1307_n 0.0108399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_301_74#_c_1415_n 0.0142211f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=2.125
cc_217 VPB N_A_301_74#_c_1410_n 0.0037373f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.635
cc_218 VPB N_A_301_74#_c_1417_n 0.00165322f $X=-0.19 $Y=1.66 $X2=0.17 $Y2=0.567
cc_219 VPB N_A_301_74#_c_1418_n 0.00168453f $X=-0.19 $Y=1.66 $X2=0.32 $Y2=1.825
cc_220 VPB N_A_301_74#_c_1419_n 0.0114349f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.69
cc_221 VPB N_A_301_74#_c_1420_n 0.00475731f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.635
cc_222 VPB N_A_301_74#_c_1421_n 0.00927489f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.69
cc_223 VPB Q 0.0540116f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.525
cc_224 N_A_35_74#_M1020_g N_SCE_c_321_n 0.00319777f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_225 N_A_35_74#_c_227_n N_SCE_c_321_n 0.0166247f $X=0.17 $Y=1.525 $X2=0 $Y2=0
cc_226 N_A_35_74#_c_231_n N_SCE_c_321_n 0.0181152f $X=0.66 $Y=1.69 $X2=0 $Y2=0
cc_227 N_A_35_74#_c_232_n N_SCE_c_321_n 0.0234495f $X=0.825 $Y=1.825 $X2=0 $Y2=0
cc_228 N_A_35_74#_c_232_n N_SCE_c_322_n 0.00797249f $X=0.825 $Y=1.825 $X2=0
+ $Y2=0
cc_229 N_A_35_74#_c_227_n N_SCE_c_323_n 0.00937938f $X=0.17 $Y=1.525 $X2=0 $Y2=0
cc_230 N_A_35_74#_c_230_n N_SCE_c_323_n 0.00519217f $X=0.32 $Y=0.565 $X2=0 $Y2=0
cc_231 N_A_35_74#_c_235_n N_SCE_c_332_n 0.0103233f $X=0.39 $Y=2.465 $X2=0 $Y2=0
cc_232 N_A_35_74#_c_231_n N_SCE_c_332_n 0.0181427f $X=0.66 $Y=1.69 $X2=0 $Y2=0
cc_233 N_A_35_74#_c_232_n N_SCE_c_332_n 0.00738429f $X=0.825 $Y=1.825 $X2=0
+ $Y2=0
cc_234 N_A_35_74#_c_235_n N_SCE_c_333_n 0.00764266f $X=0.39 $Y=2.465 $X2=0 $Y2=0
cc_235 N_A_35_74#_c_232_n N_SCE_c_333_n 0.00129587f $X=0.825 $Y=1.825 $X2=0
+ $Y2=0
cc_236 N_A_35_74#_M1020_g N_SCE_M1006_g 0.0154845f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_237 N_A_35_74#_c_227_n N_SCE_M1006_g 0.00558859f $X=0.17 $Y=1.525 $X2=0 $Y2=0
cc_238 N_A_35_74#_c_230_n N_SCE_M1006_g 8.85432e-19 $X=0.32 $Y=0.565 $X2=0 $Y2=0
cc_239 N_A_35_74#_c_235_n N_SCE_c_334_n 0.0110849f $X=0.39 $Y=2.465 $X2=0 $Y2=0
cc_240 N_A_35_74#_c_236_n N_SCE_c_335_n 0.0149882f $X=1.865 $Y=2.04 $X2=0 $Y2=0
cc_241 N_A_35_74#_c_231_n N_SCE_c_335_n 0.00723285f $X=0.66 $Y=1.69 $X2=0 $Y2=0
cc_242 N_A_35_74#_c_232_n N_SCE_c_335_n 0.00384547f $X=0.825 $Y=1.825 $X2=0
+ $Y2=0
cc_243 N_A_35_74#_c_235_n N_SCE_c_336_n 4.29561e-19 $X=0.39 $Y=2.465 $X2=0 $Y2=0
cc_244 N_A_35_74#_c_235_n N_SCE_c_337_n 0.00615422f $X=0.39 $Y=2.465 $X2=0 $Y2=0
cc_245 N_A_35_74#_c_232_n N_SCE_c_337_n 0.0101853f $X=0.825 $Y=1.825 $X2=0 $Y2=0
cc_246 N_A_35_74#_M1020_g N_SCE_c_325_n 0.0213749f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_247 N_A_35_74#_c_227_n N_SCE_c_325_n 0.00126186f $X=0.17 $Y=1.525 $X2=0 $Y2=0
cc_248 N_A_35_74#_c_231_n N_SCE_c_325_n 0.013832f $X=0.66 $Y=1.69 $X2=0 $Y2=0
cc_249 N_A_35_74#_c_232_n N_SCE_c_325_n 0.00102275f $X=0.825 $Y=1.825 $X2=0
+ $Y2=0
cc_250 N_A_35_74#_c_228_n N_SCE_c_326_n 0.0260915f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_251 N_A_35_74#_c_229_n N_SCE_c_326_n 0.00136357f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_252 N_A_35_74#_c_228_n N_SCE_c_327_n 3.10542e-19 $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_253 N_A_35_74#_c_229_n N_SCE_c_327_n 0.0152145f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_254 N_A_35_74#_M1020_g N_SCE_c_329_n 0.0152416f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_255 N_A_35_74#_c_227_n N_SCE_c_329_n 0.0256551f $X=0.17 $Y=1.525 $X2=0 $Y2=0
cc_256 N_A_35_74#_c_236_n N_SCE_c_329_n 0.0137806f $X=1.865 $Y=2.04 $X2=0 $Y2=0
cc_257 N_A_35_74#_c_231_n N_SCE_c_329_n 0.00570233f $X=0.66 $Y=1.69 $X2=0 $Y2=0
cc_258 N_A_35_74#_c_232_n N_SCE_c_329_n 0.0244961f $X=0.825 $Y=1.825 $X2=0 $Y2=0
cc_259 N_A_35_74#_M1020_g N_SCE_c_330_n 0.00958558f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_260 N_A_35_74#_M1020_g N_D_M1021_g 0.0647188f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_261 N_A_35_74#_M1027_g N_D_M1025_g 0.0164941f $X=1.985 $Y=2.64 $X2=0 $Y2=0
cc_262 N_A_35_74#_c_236_n N_D_M1025_g 0.0178488f $X=1.865 $Y=2.04 $X2=0 $Y2=0
cc_263 N_A_35_74#_c_228_n N_D_M1025_g 0.00111327f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_264 N_A_35_74#_c_229_n N_D_M1025_g 0.0196508f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_265 N_A_35_74#_c_231_n N_D_M1025_g 9.65951e-19 $X=0.66 $Y=1.69 $X2=0 $Y2=0
cc_266 N_A_35_74#_c_232_n N_D_M1025_g 0.00297182f $X=0.825 $Y=1.825 $X2=0 $Y2=0
cc_267 N_A_35_74#_M1020_g N_D_c_409_n 0.0142617f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_268 N_A_35_74#_c_236_n N_D_c_409_n 0.00371768f $X=1.865 $Y=2.04 $X2=0 $Y2=0
cc_269 N_A_35_74#_c_228_n N_D_c_409_n 3.9661e-19 $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_270 N_A_35_74#_c_229_n N_D_c_409_n 0.0198258f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_271 N_A_35_74#_c_231_n N_D_c_409_n 0.0021383f $X=0.66 $Y=1.69 $X2=0 $Y2=0
cc_272 N_A_35_74#_M1020_g N_D_c_410_n 0.00420444f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_273 N_A_35_74#_c_236_n N_D_c_410_n 0.0431554f $X=1.865 $Y=2.04 $X2=0 $Y2=0
cc_274 N_A_35_74#_c_228_n N_D_c_410_n 0.0208514f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_275 N_A_35_74#_c_229_n N_D_c_410_n 0.00109252f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_276 N_A_35_74#_c_231_n N_D_c_410_n 0.00527649f $X=0.66 $Y=1.69 $X2=0 $Y2=0
cc_277 N_A_35_74#_c_232_n N_D_c_410_n 0.0157949f $X=0.825 $Y=1.825 $X2=0 $Y2=0
cc_278 N_A_35_74#_M1027_g N_SCD_M1002_g 0.0333797f $X=1.985 $Y=2.64 $X2=0 $Y2=0
cc_279 N_A_35_74#_c_234_n N_SCD_c_448_n 0.0205499f $X=2.03 $Y=2.14 $X2=0 $Y2=0
cc_280 N_A_35_74#_c_236_n N_SCD_c_448_n 6.39715e-19 $X=1.865 $Y=2.04 $X2=0 $Y2=0
cc_281 N_A_35_74#_c_236_n SCD 0.0123499f $X=1.865 $Y=2.04 $X2=0 $Y2=0
cc_282 N_A_35_74#_c_228_n SCD 0.0307081f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_283 N_A_35_74#_c_229_n SCD 0.00192082f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_284 N_A_35_74#_c_228_n N_SCD_c_450_n 0.00168573f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_285 N_A_35_74#_c_229_n N_SCD_c_450_n 0.0205499f $X=2.03 $Y=1.635 $X2=0 $Y2=0
cc_286 N_A_35_74#_c_235_n N_VPWR_c_1288_n 0.0285143f $X=0.39 $Y=2.465 $X2=0
+ $Y2=0
cc_287 N_A_35_74#_c_232_n N_VPWR_c_1288_n 0.0263993f $X=0.825 $Y=1.825 $X2=0
+ $Y2=0
cc_288 N_A_35_74#_c_235_n N_VPWR_c_1294_n 0.0207959f $X=0.39 $Y=2.465 $X2=0
+ $Y2=0
cc_289 N_A_35_74#_M1027_g N_VPWR_c_1296_n 0.005209f $X=1.985 $Y=2.64 $X2=0 $Y2=0
cc_290 N_A_35_74#_M1027_g N_VPWR_c_1287_n 0.00537521f $X=1.985 $Y=2.64 $X2=0
+ $Y2=0
cc_291 N_A_35_74#_c_235_n N_VPWR_c_1287_n 0.0171449f $X=0.39 $Y=2.465 $X2=0
+ $Y2=0
cc_292 N_A_35_74#_M1020_g N_A_301_74#_c_1422_n 9.49989e-19 $X=1.04 $Y=0.58 $X2=0
+ $Y2=0
cc_293 N_A_35_74#_M1027_g N_A_301_74#_c_1415_n 0.010261f $X=1.985 $Y=2.64 $X2=0
+ $Y2=0
cc_294 N_A_35_74#_c_234_n N_A_301_74#_c_1415_n 8.35672e-19 $X=2.03 $Y=2.14 $X2=0
+ $Y2=0
cc_295 N_A_35_74#_c_236_n N_A_301_74#_c_1415_n 0.0209566f $X=1.865 $Y=2.04 $X2=0
+ $Y2=0
cc_296 N_A_35_74#_M1027_g N_A_301_74#_c_1420_n 0.0116864f $X=1.985 $Y=2.64 $X2=0
+ $Y2=0
cc_297 N_A_35_74#_c_234_n N_A_301_74#_c_1420_n 2.33387e-19 $X=2.03 $Y=2.14 $X2=0
+ $Y2=0
cc_298 N_A_35_74#_c_236_n N_A_301_74#_c_1420_n 0.0263677f $X=1.865 $Y=2.04 $X2=0
+ $Y2=0
cc_299 N_A_35_74#_M1020_g N_VGND_c_1556_n 0.00578925f $X=1.04 $Y=0.58 $X2=0
+ $Y2=0
cc_300 N_A_35_74#_c_230_n N_VGND_c_1556_n 0.0163081f $X=0.32 $Y=0.565 $X2=0
+ $Y2=0
cc_301 N_A_35_74#_M1020_g N_VGND_c_1562_n 0.00461464f $X=1.04 $Y=0.58 $X2=0
+ $Y2=0
cc_302 N_A_35_74#_c_230_n N_VGND_c_1566_n 0.0137679f $X=0.32 $Y=0.565 $X2=0
+ $Y2=0
cc_303 N_A_35_74#_M1020_g N_VGND_c_1571_n 0.0081824f $X=1.04 $Y=0.58 $X2=0 $Y2=0
cc_304 N_A_35_74#_c_230_n N_VGND_c_1571_n 0.0116365f $X=0.32 $Y=0.565 $X2=0
+ $Y2=0
cc_305 N_SCE_c_326_n N_D_M1021_g 0.0242708f $X=2.085 $Y=1.065 $X2=0 $Y2=0
cc_306 N_SCE_c_327_n N_D_M1021_g 0.00867602f $X=2.085 $Y=1.065 $X2=0 $Y2=0
cc_307 N_SCE_c_328_n N_D_M1021_g 0.0129182f $X=2.085 $Y=0.9 $X2=0 $Y2=0
cc_308 N_SCE_c_330_n N_D_M1021_g 0.00225056f $X=1.315 $Y=1.047 $X2=0 $Y2=0
cc_309 N_SCE_c_335_n N_D_M1025_g 0.0532994f $X=1.025 $Y=2.17 $X2=0 $Y2=0
cc_310 N_SCE_c_326_n N_D_c_409_n 0.00459016f $X=2.085 $Y=1.065 $X2=0 $Y2=0
cc_311 N_SCE_c_335_n N_D_c_410_n 5.5141e-19 $X=1.025 $Y=2.17 $X2=0 $Y2=0
cc_312 N_SCE_c_330_n N_D_c_410_n 0.0460537f $X=1.315 $Y=1.047 $X2=0 $Y2=0
cc_313 N_SCE_c_326_n N_SCD_M1028_g 7.27759e-19 $X=2.085 $Y=1.065 $X2=0 $Y2=0
cc_314 N_SCE_c_328_n N_SCD_M1028_g 0.053304f $X=2.085 $Y=0.9 $X2=0 $Y2=0
cc_315 N_SCE_c_334_n N_VPWR_c_1288_n 0.00351947f $X=0.615 $Y=2.245 $X2=0 $Y2=0
cc_316 N_SCE_c_335_n N_VPWR_c_1288_n 0.00323965f $X=1.025 $Y=2.17 $X2=0 $Y2=0
cc_317 N_SCE_c_336_n N_VPWR_c_1288_n 0.0173553f $X=1.115 $Y=2.245 $X2=0 $Y2=0
cc_318 N_SCE_c_334_n N_VPWR_c_1294_n 0.005209f $X=0.615 $Y=2.245 $X2=0 $Y2=0
cc_319 N_SCE_c_336_n N_VPWR_c_1296_n 0.00460063f $X=1.115 $Y=2.245 $X2=0 $Y2=0
cc_320 N_SCE_c_334_n N_VPWR_c_1287_n 0.0098615f $X=0.615 $Y=2.245 $X2=0 $Y2=0
cc_321 N_SCE_c_336_n N_VPWR_c_1287_n 0.00908371f $X=1.115 $Y=2.245 $X2=0 $Y2=0
cc_322 N_SCE_c_326_n N_A_301_74#_c_1422_n 0.0568015f $X=2.085 $Y=1.065 $X2=0
+ $Y2=0
cc_323 N_SCE_c_327_n N_A_301_74#_c_1422_n 0.00395514f $X=2.085 $Y=1.065 $X2=0
+ $Y2=0
cc_324 N_SCE_c_328_n N_A_301_74#_c_1422_n 0.018235f $X=2.085 $Y=0.9 $X2=0 $Y2=0
cc_325 N_SCE_c_326_n N_A_301_74#_c_1407_n 0.0182629f $X=2.085 $Y=1.065 $X2=0
+ $Y2=0
cc_326 N_SCE_c_327_n N_A_301_74#_c_1407_n 6.89219e-19 $X=2.085 $Y=1.065 $X2=0
+ $Y2=0
cc_327 N_SCE_c_328_n N_A_301_74#_c_1407_n 0.0034424f $X=2.085 $Y=0.9 $X2=0 $Y2=0
cc_328 N_SCE_c_326_n N_A_301_74#_c_1409_n 0.0139422f $X=2.085 $Y=1.065 $X2=0
+ $Y2=0
cc_329 N_SCE_c_327_n N_A_301_74#_c_1409_n 3.81179e-19 $X=2.085 $Y=1.065 $X2=0
+ $Y2=0
cc_330 N_SCE_c_336_n N_A_301_74#_c_1420_n 0.0018968f $X=1.115 $Y=2.245 $X2=0
+ $Y2=0
cc_331 N_SCE_M1006_g N_VGND_c_1556_n 0.0121355f $X=0.535 $Y=0.58 $X2=0 $Y2=0
cc_332 N_SCE_c_325_n N_VGND_c_1556_n 0.00320419f $X=0.59 $Y=1.12 $X2=0 $Y2=0
cc_333 N_SCE_c_329_n N_VGND_c_1556_n 0.0248464f $X=1.085 $Y=1.047 $X2=0 $Y2=0
cc_334 N_SCE_c_328_n N_VGND_c_1562_n 0.00298292f $X=2.085 $Y=0.9 $X2=0 $Y2=0
cc_335 N_SCE_M1006_g N_VGND_c_1566_n 0.00383152f $X=0.535 $Y=0.58 $X2=0 $Y2=0
cc_336 N_SCE_M1006_g N_VGND_c_1571_n 0.00761327f $X=0.535 $Y=0.58 $X2=0 $Y2=0
cc_337 N_SCE_c_328_n N_VGND_c_1571_n 0.00367497f $X=2.085 $Y=0.9 $X2=0 $Y2=0
cc_338 N_SCE_c_330_n N_VGND_c_1571_n 0.0087477f $X=1.315 $Y=1.047 $X2=0 $Y2=0
cc_339 N_D_M1025_g N_VPWR_c_1288_n 0.00249078f $X=1.535 $Y=2.64 $X2=0 $Y2=0
cc_340 N_D_M1025_g N_VPWR_c_1296_n 0.005209f $X=1.535 $Y=2.64 $X2=0 $Y2=0
cc_341 N_D_M1025_g N_VPWR_c_1287_n 0.00983291f $X=1.535 $Y=2.64 $X2=0 $Y2=0
cc_342 N_D_M1021_g N_A_301_74#_c_1422_n 0.0126349f $X=1.43 $Y=0.58 $X2=0 $Y2=0
cc_343 N_D_M1025_g N_A_301_74#_c_1420_n 0.0134434f $X=1.535 $Y=2.64 $X2=0 $Y2=0
cc_344 N_D_M1021_g N_VGND_c_1562_n 0.00439708f $X=1.43 $Y=0.58 $X2=0 $Y2=0
cc_345 N_D_M1021_g N_VGND_c_1571_n 0.0083885f $X=1.43 $Y=0.58 $X2=0 $Y2=0
cc_346 N_SCD_M1028_g N_CLK_c_493_n 0.0271743f $X=2.565 $Y=0.58 $X2=-0.19
+ $Y2=-0.245
cc_347 N_SCD_M1002_g N_CLK_M1004_g 0.0171374f $X=2.525 $Y=2.64 $X2=0 $Y2=0
cc_348 N_SCD_c_448_n N_CLK_M1004_g 0.00794241f $X=2.57 $Y=1.975 $X2=0 $Y2=0
cc_349 N_SCD_M1028_g N_CLK_c_496_n 0.00161101f $X=2.565 $Y=0.58 $X2=0 $Y2=0
cc_350 N_SCD_c_450_n N_CLK_c_496_n 0.00794241f $X=2.57 $Y=1.635 $X2=0 $Y2=0
cc_351 N_SCD_M1028_g N_A_630_74#_c_746_n 5.10107e-19 $X=2.565 $Y=0.58 $X2=0
+ $Y2=0
cc_352 N_SCD_M1002_g N_VPWR_c_1289_n 0.00651263f $X=2.525 $Y=2.64 $X2=0 $Y2=0
cc_353 N_SCD_M1002_g N_VPWR_c_1296_n 0.00553757f $X=2.525 $Y=2.64 $X2=0 $Y2=0
cc_354 N_SCD_M1002_g N_VPWR_c_1287_n 0.0056107f $X=2.525 $Y=2.64 $X2=0 $Y2=0
cc_355 N_SCD_M1028_g N_A_301_74#_c_1422_n 0.00976024f $X=2.565 $Y=0.58 $X2=0
+ $Y2=0
cc_356 N_SCD_M1002_g N_A_301_74#_c_1415_n 0.0149545f $X=2.525 $Y=2.64 $X2=0
+ $Y2=0
cc_357 N_SCD_c_453_n N_A_301_74#_c_1415_n 0.00103741f $X=2.57 $Y=2.14 $X2=0
+ $Y2=0
cc_358 SCD N_A_301_74#_c_1415_n 0.0259252f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_359 N_SCD_M1028_g N_A_301_74#_c_1407_n 0.0105397f $X=2.565 $Y=0.58 $X2=0
+ $Y2=0
cc_360 N_SCD_M1028_g N_A_301_74#_c_1408_n 0.005999f $X=2.565 $Y=0.58 $X2=0 $Y2=0
cc_361 SCD N_A_301_74#_c_1408_n 0.0116904f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_362 N_SCD_c_450_n N_A_301_74#_c_1408_n 6.61574e-19 $X=2.57 $Y=1.635 $X2=0
+ $Y2=0
cc_363 N_SCD_M1028_g N_A_301_74#_c_1409_n 0.00455678f $X=2.565 $Y=0.58 $X2=0
+ $Y2=0
cc_364 SCD N_A_301_74#_c_1409_n 0.0146897f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_365 N_SCD_c_450_n N_A_301_74#_c_1409_n 5.47548e-19 $X=2.57 $Y=1.635 $X2=0
+ $Y2=0
cc_366 N_SCD_M1002_g N_A_301_74#_c_1410_n 0.00337201f $X=2.525 $Y=2.64 $X2=0
+ $Y2=0
cc_367 N_SCD_M1028_g N_A_301_74#_c_1410_n 0.00333054f $X=2.565 $Y=0.58 $X2=0
+ $Y2=0
cc_368 SCD N_A_301_74#_c_1410_n 0.052777f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_369 N_SCD_c_450_n N_A_301_74#_c_1410_n 0.00233284f $X=2.57 $Y=1.635 $X2=0
+ $Y2=0
cc_370 N_SCD_M1002_g N_A_301_74#_c_1420_n 0.00229868f $X=2.525 $Y=2.64 $X2=0
+ $Y2=0
cc_371 N_SCD_M1028_g N_VGND_c_1557_n 0.00630066f $X=2.565 $Y=0.58 $X2=0 $Y2=0
cc_372 N_SCD_M1028_g N_VGND_c_1562_n 0.00352596f $X=2.565 $Y=0.58 $X2=0 $Y2=0
cc_373 N_SCD_M1028_g N_VGND_c_1571_n 0.00547145f $X=2.565 $Y=0.58 $X2=0 $Y2=0
cc_374 CLK N_A_630_74#_M1018_g 4.50002e-19 $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_375 N_CLK_c_496_n N_A_630_74#_M1018_g 0.00213289f $X=3.235 $Y=1.385 $X2=0
+ $Y2=0
cc_376 N_CLK_c_493_n N_A_630_74#_c_744_n 0.00521767f $X=3.075 $Y=1.22 $X2=0
+ $Y2=0
cc_377 N_CLK_M1004_g N_A_630_74#_c_757_n 0.00537037f $X=3.235 $Y=2.4 $X2=0 $Y2=0
cc_378 CLK N_A_630_74#_c_757_n 0.0223297f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_379 N_CLK_c_496_n N_A_630_74#_c_757_n 0.00544741f $X=3.235 $Y=1.385 $X2=0
+ $Y2=0
cc_380 CLK N_A_630_74#_c_745_n 0.0153326f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_381 N_CLK_c_496_n N_A_630_74#_c_745_n 7.56949e-19 $X=3.235 $Y=1.385 $X2=0
+ $Y2=0
cc_382 N_CLK_c_493_n N_A_630_74#_c_746_n 0.00395607f $X=3.075 $Y=1.22 $X2=0
+ $Y2=0
cc_383 CLK N_A_630_74#_c_746_n 0.0147852f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_384 N_CLK_c_496_n N_A_630_74#_c_746_n 0.00451028f $X=3.235 $Y=1.385 $X2=0
+ $Y2=0
cc_385 N_CLK_c_496_n N_A_630_74#_c_779_n 2.27554e-19 $X=3.235 $Y=1.385 $X2=0
+ $Y2=0
cc_386 N_CLK_M1004_g N_A_630_74#_c_747_n 0.00503406f $X=3.235 $Y=2.4 $X2=0 $Y2=0
cc_387 N_CLK_M1004_g N_A_630_74#_c_748_n 0.0024946f $X=3.235 $Y=2.4 $X2=0 $Y2=0
cc_388 CLK N_A_630_74#_c_748_n 0.00170318f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_389 N_CLK_c_496_n N_A_630_74#_c_748_n 0.015847f $X=3.235 $Y=1.385 $X2=0 $Y2=0
cc_390 CLK N_A_630_74#_c_749_n 0.0291649f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_391 N_CLK_c_496_n N_A_630_74#_c_749_n 2.12609e-19 $X=3.235 $Y=1.385 $X2=0
+ $Y2=0
cc_392 N_CLK_M1004_g N_VPWR_c_1289_n 0.0288306f $X=3.235 $Y=2.4 $X2=0 $Y2=0
cc_393 N_CLK_M1004_g N_VPWR_c_1290_n 0.00980791f $X=3.235 $Y=2.4 $X2=0 $Y2=0
cc_394 N_CLK_M1004_g N_VPWR_c_1300_n 0.00460063f $X=3.235 $Y=2.4 $X2=0 $Y2=0
cc_395 N_CLK_M1004_g N_VPWR_c_1287_n 0.00468499f $X=3.235 $Y=2.4 $X2=0 $Y2=0
cc_396 N_CLK_c_493_n N_A_301_74#_c_1407_n 0.00144764f $X=3.075 $Y=1.22 $X2=0
+ $Y2=0
cc_397 N_CLK_c_493_n N_A_301_74#_c_1408_n 0.00858861f $X=3.075 $Y=1.22 $X2=0
+ $Y2=0
cc_398 CLK N_A_301_74#_c_1408_n 0.00984264f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_399 N_CLK_c_496_n N_A_301_74#_c_1408_n 0.00291916f $X=3.235 $Y=1.385 $X2=0
+ $Y2=0
cc_400 CLK N_A_301_74#_c_1410_n 0.0189121f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_401 N_CLK_c_496_n N_A_301_74#_c_1410_n 0.0203085f $X=3.235 $Y=1.385 $X2=0
+ $Y2=0
cc_402 N_CLK_M1004_g N_A_301_74#_c_1462_n 0.0209338f $X=3.235 $Y=2.4 $X2=0 $Y2=0
cc_403 N_CLK_c_493_n N_VGND_c_1557_n 0.00319344f $X=3.075 $Y=1.22 $X2=0 $Y2=0
cc_404 N_CLK_c_493_n N_VGND_c_1558_n 0.00324671f $X=3.075 $Y=1.22 $X2=0 $Y2=0
cc_405 N_CLK_c_493_n N_VGND_c_1564_n 0.00434272f $X=3.075 $Y=1.22 $X2=0 $Y2=0
cc_406 N_CLK_c_493_n N_VGND_c_1571_n 0.00826076f $X=3.075 $Y=1.22 $X2=0 $Y2=0
cc_407 N_A_828_74#_c_537_n N_A_630_74#_M1018_g 0.0015901f $X=4.28 $Y=0.515 $X2=0
+ $Y2=0
cc_408 N_A_828_74#_c_539_n N_A_630_74#_M1018_g 0.00266901f $X=4.445 $Y=0.34
+ $X2=0 $Y2=0
cc_409 N_A_828_74#_c_537_n N_A_630_74#_c_734_n 0.00119028f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_410 N_A_828_74#_c_540_n N_A_630_74#_M1008_g 5.82776e-19 $X=5.14 $Y=2.05 $X2=0
+ $Y2=0
cc_411 N_A_828_74#_c_560_n N_A_630_74#_M1008_g 8.469e-19 $X=5.12 $Y=2.215 $X2=0
+ $Y2=0
cc_412 N_A_828_74#_c_561_n N_A_630_74#_M1008_g 0.00582615f $X=5.12 $Y=2.215
+ $X2=0 $Y2=0
cc_413 N_A_828_74#_c_560_n N_A_630_74#_c_736_n 0.00242763f $X=5.12 $Y=2.215
+ $X2=0 $Y2=0
cc_414 N_A_828_74#_c_536_n N_A_630_74#_M1007_g 0.0133683f $X=5.695 $Y=1.03 $X2=0
+ $Y2=0
cc_415 N_A_828_74#_c_537_n N_A_630_74#_M1007_g 0.00315776f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_416 N_A_828_74#_c_538_n N_A_630_74#_M1007_g 0.00881128f $X=5.055 $Y=0.34
+ $X2=0 $Y2=0
cc_417 N_A_828_74#_c_540_n N_A_630_74#_M1007_g 0.028068f $X=5.14 $Y=2.05 $X2=0
+ $Y2=0
cc_418 N_A_828_74#_c_549_n N_A_630_74#_M1007_g 0.00175971f $X=5.14 $Y=0.34 $X2=0
+ $Y2=0
cc_419 N_A_828_74#_c_540_n N_A_630_74#_c_753_n 0.0083267f $X=5.14 $Y=2.05 $X2=0
+ $Y2=0
cc_420 N_A_828_74#_c_543_n N_A_630_74#_c_753_n 2.41031e-19 $X=5.82 $Y=1.195
+ $X2=0 $Y2=0
cc_421 N_A_828_74#_c_544_n N_A_630_74#_c_753_n 0.0133536f $X=5.82 $Y=1.195 $X2=0
+ $Y2=0
cc_422 N_A_828_74#_c_561_n N_A_630_74#_c_753_n 0.00817017f $X=5.12 $Y=2.215
+ $X2=0 $Y2=0
cc_423 N_A_828_74#_c_561_n N_A_630_74#_M1013_g 0.0185677f $X=5.12 $Y=2.215 $X2=0
+ $Y2=0
cc_424 N_A_828_74#_c_556_n N_A_630_74#_M1026_g 0.0190696f $X=8.47 $Y=1.91 $X2=0
+ $Y2=0
cc_425 N_A_828_74#_c_558_n N_A_630_74#_M1026_g 5.48409e-19 $X=8.47 $Y=1.57 $X2=0
+ $Y2=0
cc_426 N_A_828_74#_c_547_n N_A_630_74#_c_738_n 0.0224602f $X=8.07 $Y=1.275 $X2=0
+ $Y2=0
cc_427 N_A_828_74#_c_558_n N_A_630_74#_c_738_n 0.00137931f $X=8.47 $Y=1.57 $X2=0
+ $Y2=0
cc_428 N_A_828_74#_c_548_n N_A_630_74#_c_738_n 0.0223365f $X=8.47 $Y=1.57 $X2=0
+ $Y2=0
cc_429 N_A_828_74#_c_550_n N_A_630_74#_c_738_n 0.00145063f $X=7.57 $Y=1.195
+ $X2=0 $Y2=0
cc_430 N_A_828_74#_c_547_n N_A_630_74#_c_739_n 0.00640549f $X=8.07 $Y=1.275
+ $X2=0 $Y2=0
cc_431 N_A_828_74#_c_548_n N_A_630_74#_c_739_n 0.00754759f $X=8.47 $Y=1.57 $X2=0
+ $Y2=0
cc_432 N_A_828_74#_c_551_n N_A_630_74#_c_740_n 0.0210721f $X=7.57 $Y=1.195 $X2=0
+ $Y2=0
cc_433 N_A_828_74#_c_552_n N_A_630_74#_c_740_n 0.00129449f $X=7.65 $Y=1.03 $X2=0
+ $Y2=0
cc_434 N_A_828_74#_c_553_n N_A_630_74#_c_740_n 4.15839e-19 $X=7.57 $Y=1.03 $X2=0
+ $Y2=0
cc_435 N_A_828_74#_c_545_n N_A_630_74#_c_741_n 0.0011964f $X=7.645 $Y=0.34 $X2=0
+ $Y2=0
cc_436 N_A_828_74#_c_552_n N_A_630_74#_c_741_n 0.00213389f $X=7.65 $Y=1.03 $X2=0
+ $Y2=0
cc_437 N_A_828_74#_c_553_n N_A_630_74#_c_741_n 0.00408693f $X=7.57 $Y=1.03 $X2=0
+ $Y2=0
cc_438 N_A_828_74#_c_537_n N_A_630_74#_c_742_n 0.00118383f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_439 N_A_828_74#_c_540_n N_A_630_74#_c_743_n 0.0110783f $X=5.14 $Y=2.05 $X2=0
+ $Y2=0
cc_440 N_A_828_74#_c_560_n N_A_630_74#_c_743_n 0.00121268f $X=5.12 $Y=2.215
+ $X2=0 $Y2=0
cc_441 N_A_828_74#_c_561_n N_A_630_74#_c_743_n 0.0222307f $X=5.12 $Y=2.215 $X2=0
+ $Y2=0
cc_442 N_A_828_74#_c_556_n N_A_630_74#_c_761_n 7.44721e-19 $X=8.47 $Y=1.91 $X2=0
+ $Y2=0
cc_443 N_A_828_74#_c_558_n N_A_630_74#_c_761_n 0.00361184f $X=8.47 $Y=1.57 $X2=0
+ $Y2=0
cc_444 N_A_828_74#_c_537_n N_A_630_74#_c_749_n 0.00648541f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_445 N_A_828_74#_c_547_n N_A_630_74#_c_750_n 0.00493576f $X=8.07 $Y=1.275
+ $X2=0 $Y2=0
cc_446 N_A_828_74#_c_558_n N_A_630_74#_c_750_n 0.0120505f $X=8.47 $Y=1.57 $X2=0
+ $Y2=0
cc_447 N_A_828_74#_c_548_n N_A_630_74#_c_750_n 0.0011416f $X=8.47 $Y=1.57 $X2=0
+ $Y2=0
cc_448 N_A_828_74#_c_550_n N_A_630_74#_c_750_n 0.0164206f $X=7.57 $Y=1.195 $X2=0
+ $Y2=0
cc_449 N_A_828_74#_c_551_n N_A_630_74#_c_750_n 3.83408e-19 $X=7.57 $Y=1.195
+ $X2=0 $Y2=0
cc_450 N_A_828_74#_c_547_n N_A_630_74#_c_751_n 0.00324689f $X=8.07 $Y=1.275
+ $X2=0 $Y2=0
cc_451 N_A_828_74#_c_558_n N_A_630_74#_c_751_n 2.22243e-19 $X=8.47 $Y=1.57 $X2=0
+ $Y2=0
cc_452 N_A_828_74#_c_548_n N_A_630_74#_c_751_n 0.00491918f $X=8.47 $Y=1.57 $X2=0
+ $Y2=0
cc_453 N_A_828_74#_c_550_n N_A_630_74#_c_751_n 0.00253213f $X=7.57 $Y=1.195
+ $X2=0 $Y2=0
cc_454 N_A_828_74#_c_551_n N_A_630_74#_c_751_n 0.00934794f $X=7.57 $Y=1.195
+ $X2=0 $Y2=0
cc_455 N_A_828_74#_c_561_n N_A_630_74#_c_766_n 0.00320751f $X=5.12 $Y=2.215
+ $X2=0 $Y2=0
cc_456 N_A_828_74#_c_545_n N_A_1239_74#_M1011_d 0.00181776f $X=7.645 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_457 N_A_828_74#_c_543_n N_A_1239_74#_c_946_n 0.0216554f $X=5.82 $Y=1.195
+ $X2=0 $Y2=0
cc_458 N_A_828_74#_c_544_n N_A_1239_74#_c_946_n 0.0011618f $X=5.82 $Y=1.195
+ $X2=0 $Y2=0
cc_459 N_A_828_74#_c_614_p N_A_1239_74#_c_946_n 0.0575793f $X=6.805 $Y=0.775
+ $X2=0 $Y2=0
cc_460 N_A_828_74#_c_545_n N_A_1239_74#_c_946_n 0.00392224f $X=7.645 $Y=0.34
+ $X2=0 $Y2=0
cc_461 N_A_828_74#_c_543_n N_A_1239_74#_c_947_n 4.15752e-19 $X=5.82 $Y=1.195
+ $X2=0 $Y2=0
cc_462 N_A_828_74#_c_544_n N_A_1239_74#_c_947_n 0.020933f $X=5.82 $Y=1.195 $X2=0
+ $Y2=0
cc_463 N_A_828_74#_c_614_p N_A_1239_74#_c_947_n 0.00422584f $X=6.805 $Y=0.775
+ $X2=0 $Y2=0
cc_464 N_A_828_74#_c_552_n N_A_1239_74#_c_948_n 0.00646115f $X=7.65 $Y=1.03
+ $X2=0 $Y2=0
cc_465 N_A_828_74#_c_553_n N_A_1239_74#_c_948_n 0.00125838f $X=7.57 $Y=1.03
+ $X2=0 $Y2=0
cc_466 N_A_828_74#_c_545_n N_A_1239_74#_c_967_n 0.0154872f $X=7.645 $Y=0.34
+ $X2=0 $Y2=0
cc_467 N_A_828_74#_c_553_n N_A_1239_74#_c_967_n 0.00414841f $X=7.57 $Y=1.03
+ $X2=0 $Y2=0
cc_468 N_A_828_74#_c_550_n N_A_1239_74#_c_950_n 0.0278269f $X=7.57 $Y=1.195
+ $X2=0 $Y2=0
cc_469 N_A_828_74#_c_551_n N_A_1239_74#_c_950_n 0.0025345f $X=7.57 $Y=1.195
+ $X2=0 $Y2=0
cc_470 N_A_828_74#_c_536_n N_A_1239_74#_c_951_n 0.0154821f $X=5.695 $Y=1.03
+ $X2=0 $Y2=0
cc_471 N_A_828_74#_c_541_n N_A_1239_74#_c_951_n 5.48134e-19 $X=5.735 $Y=0.34
+ $X2=0 $Y2=0
cc_472 N_A_828_74#_c_542_n N_A_1239_74#_c_951_n 0.00400832f $X=5.82 $Y=0.69
+ $X2=0 $Y2=0
cc_473 N_A_828_74#_c_543_n N_A_1239_74#_c_951_n 0.00382001f $X=5.82 $Y=1.195
+ $X2=0 $Y2=0
cc_474 N_A_828_74#_c_614_p N_A_1239_74#_c_951_n 0.0137143f $X=6.805 $Y=0.775
+ $X2=0 $Y2=0
cc_475 N_A_828_74#_c_630_p N_A_1239_74#_c_951_n 0.00299245f $X=6.89 $Y=0.69
+ $X2=0 $Y2=0
cc_476 N_A_828_74#_c_540_n N_A_1018_100#_M1007_d 0.0042575f $X=5.14 $Y=2.05
+ $X2=-0.19 $Y2=-0.245
cc_477 N_A_828_74#_c_545_n N_A_1018_100#_M1011_g 0.0118435f $X=7.645 $Y=0.34
+ $X2=0 $Y2=0
cc_478 N_A_828_74#_c_550_n N_A_1018_100#_M1011_g 2.84017e-19 $X=7.57 $Y=1.195
+ $X2=0 $Y2=0
cc_479 N_A_828_74#_c_551_n N_A_1018_100#_M1011_g 0.0171198f $X=7.57 $Y=1.195
+ $X2=0 $Y2=0
cc_480 N_A_828_74#_c_553_n N_A_1018_100#_M1011_g 0.0167881f $X=7.57 $Y=1.03
+ $X2=0 $Y2=0
cc_481 N_A_828_74#_c_536_n N_A_1018_100#_c_1023_n 0.00490388f $X=5.695 $Y=1.03
+ $X2=0 $Y2=0
cc_482 N_A_828_74#_c_540_n N_A_1018_100#_c_1023_n 0.0694974f $X=5.14 $Y=2.05
+ $X2=0 $Y2=0
cc_483 N_A_828_74#_c_541_n N_A_1018_100#_c_1023_n 0.012971f $X=5.735 $Y=0.34
+ $X2=0 $Y2=0
cc_484 N_A_828_74#_c_543_n N_A_1018_100#_c_1023_n 0.0344248f $X=5.82 $Y=1.195
+ $X2=0 $Y2=0
cc_485 N_A_828_74#_M1015_g N_A_1018_100#_c_1029_n 3.51291e-19 $X=5.435 $Y=2.75
+ $X2=0 $Y2=0
cc_486 N_A_828_74#_c_543_n N_A_1018_100#_c_1024_n 0.0198116f $X=5.82 $Y=1.195
+ $X2=0 $Y2=0
cc_487 N_A_828_74#_c_544_n N_A_1018_100#_c_1024_n 0.00346855f $X=5.82 $Y=1.195
+ $X2=0 $Y2=0
cc_488 N_A_828_74#_c_614_p N_A_1018_100#_c_1024_n 0.00499811f $X=6.805 $Y=0.775
+ $X2=0 $Y2=0
cc_489 N_A_828_74#_c_540_n N_A_1018_100#_c_1025_n 0.0142743f $X=5.14 $Y=2.05
+ $X2=0 $Y2=0
cc_490 N_A_828_74#_c_540_n N_A_1018_100#_c_1031_n 0.0252308f $X=5.14 $Y=2.05
+ $X2=0 $Y2=0
cc_491 N_A_828_74#_c_560_n N_A_1018_100#_c_1031_n 0.0249185f $X=5.12 $Y=2.215
+ $X2=0 $Y2=0
cc_492 N_A_828_74#_c_561_n N_A_1018_100#_c_1031_n 0.00798404f $X=5.12 $Y=2.215
+ $X2=0 $Y2=0
cc_493 N_A_828_74#_M1015_g N_A_1018_100#_c_1032_n 0.0139809f $X=5.435 $Y=2.75
+ $X2=0 $Y2=0
cc_494 N_A_828_74#_c_561_n N_A_1018_100#_c_1032_n 3.97086e-19 $X=5.12 $Y=2.215
+ $X2=0 $Y2=0
cc_495 N_A_828_74#_c_556_n N_A_1736_74#_c_1113_n 0.00580344f $X=8.47 $Y=1.91
+ $X2=0 $Y2=0
cc_496 N_A_828_74#_c_558_n N_A_1736_74#_c_1113_n 5.0811e-19 $X=8.47 $Y=1.57
+ $X2=0 $Y2=0
cc_497 N_A_828_74#_c_548_n N_A_1736_74#_c_1113_n 0.0347286f $X=8.47 $Y=1.57
+ $X2=0 $Y2=0
cc_498 N_A_828_74#_M1010_g N_A_1736_74#_c_1125_n 0.0421582f $X=8.365 $Y=2.75
+ $X2=0 $Y2=0
cc_499 N_A_828_74#_c_547_n N_A_1736_74#_c_1121_n 0.00109485f $X=8.07 $Y=1.275
+ $X2=0 $Y2=0
cc_500 N_A_828_74#_c_545_n N_A_1520_74#_M1000_d 0.00108545f $X=7.645 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_501 N_A_828_74#_c_552_n N_A_1520_74#_M1000_d 0.00741037f $X=7.65 $Y=1.03
+ $X2=-0.19 $Y2=-0.245
cc_502 N_A_828_74#_c_556_n N_A_1520_74#_c_1205_n 0.00199368f $X=8.47 $Y=1.91
+ $X2=0 $Y2=0
cc_503 N_A_828_74#_c_547_n N_A_1520_74#_c_1205_n 0.00224131f $X=8.07 $Y=1.275
+ $X2=0 $Y2=0
cc_504 N_A_828_74#_M1010_g N_A_1520_74#_c_1206_n 0.0146033f $X=8.365 $Y=2.75
+ $X2=0 $Y2=0
cc_505 N_A_828_74#_M1010_g N_A_1520_74#_c_1207_n 0.0185831f $X=8.365 $Y=2.75
+ $X2=0 $Y2=0
cc_506 N_A_828_74#_c_556_n N_A_1520_74#_c_1207_n 0.00401956f $X=8.47 $Y=1.91
+ $X2=0 $Y2=0
cc_507 N_A_828_74#_c_558_n N_A_1520_74#_c_1207_n 0.0192618f $X=8.47 $Y=1.57
+ $X2=0 $Y2=0
cc_508 N_A_828_74#_c_547_n N_A_1520_74#_c_1199_n 0.0187913f $X=8.07 $Y=1.275
+ $X2=0 $Y2=0
cc_509 N_A_828_74#_c_558_n N_A_1520_74#_c_1199_n 0.00802087f $X=8.47 $Y=1.57
+ $X2=0 $Y2=0
cc_510 N_A_828_74#_c_548_n N_A_1520_74#_c_1199_n 0.00129638f $X=8.47 $Y=1.57
+ $X2=0 $Y2=0
cc_511 N_A_828_74#_c_556_n N_A_1520_74#_c_1208_n 0.002823f $X=8.47 $Y=1.91 $X2=0
+ $Y2=0
cc_512 N_A_828_74#_c_558_n N_A_1520_74#_c_1208_n 0.0106323f $X=8.47 $Y=1.57
+ $X2=0 $Y2=0
cc_513 N_A_828_74#_c_547_n N_A_1520_74#_c_1202_n 0.0364823f $X=8.07 $Y=1.275
+ $X2=0 $Y2=0
cc_514 N_A_828_74#_c_548_n N_A_1520_74#_c_1202_n 0.00389197f $X=8.47 $Y=1.57
+ $X2=0 $Y2=0
cc_515 N_A_828_74#_c_552_n N_A_1520_74#_c_1202_n 0.0423843f $X=7.65 $Y=1.03
+ $X2=0 $Y2=0
cc_516 N_A_828_74#_c_558_n N_A_1520_74#_c_1203_n 0.0272725f $X=8.47 $Y=1.57
+ $X2=0 $Y2=0
cc_517 N_A_828_74#_c_548_n N_A_1520_74#_c_1203_n 0.00253041f $X=8.47 $Y=1.57
+ $X2=0 $Y2=0
cc_518 N_A_828_74#_M1010_g N_VPWR_c_1292_n 0.00211374f $X=8.365 $Y=2.75 $X2=0
+ $Y2=0
cc_519 N_A_828_74#_M1015_g N_VPWR_c_1301_n 0.00519794f $X=5.435 $Y=2.75 $X2=0
+ $Y2=0
cc_520 N_A_828_74#_M1010_g N_VPWR_c_1302_n 0.00553757f $X=8.365 $Y=2.75 $X2=0
+ $Y2=0
cc_521 N_A_828_74#_M1015_g N_VPWR_c_1287_n 0.00591991f $X=5.435 $Y=2.75 $X2=0
+ $Y2=0
cc_522 N_A_828_74#_M1010_g N_VPWR_c_1287_n 0.0109163f $X=8.365 $Y=2.75 $X2=0
+ $Y2=0
cc_523 N_A_828_74#_c_540_n N_A_301_74#_c_1417_n 0.00370176f $X=5.14 $Y=2.05
+ $X2=0 $Y2=0
cc_524 N_A_828_74#_c_560_n N_A_301_74#_c_1417_n 0.0167477f $X=5.12 $Y=2.215
+ $X2=0 $Y2=0
cc_525 N_A_828_74#_c_561_n N_A_301_74#_c_1417_n 2.0203e-19 $X=5.12 $Y=2.215
+ $X2=0 $Y2=0
cc_526 N_A_828_74#_c_537_n N_A_301_74#_c_1411_n 0.0022968f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_527 N_A_828_74#_c_540_n N_A_301_74#_c_1411_n 0.00887932f $X=5.14 $Y=2.05
+ $X2=0 $Y2=0
cc_528 N_A_828_74#_c_560_n N_A_301_74#_c_1411_n 0.0193726f $X=5.12 $Y=2.215
+ $X2=0 $Y2=0
cc_529 N_A_828_74#_c_537_n N_A_301_74#_c_1412_n 0.00879712f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_530 N_A_828_74#_M1008_d N_A_301_74#_c_1470_n 0.00263553f $X=4.515 $Y=1.84
+ $X2=0 $Y2=0
cc_531 N_A_828_74#_M1015_g N_A_301_74#_c_1470_n 0.0021205f $X=5.435 $Y=2.75
+ $X2=0 $Y2=0
cc_532 N_A_828_74#_c_537_n N_A_301_74#_c_1413_n 0.0147383f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_533 N_A_828_74#_c_540_n N_A_301_74#_c_1413_n 0.0273131f $X=5.14 $Y=2.05 $X2=0
+ $Y2=0
cc_534 N_A_828_74#_M1008_d N_A_301_74#_c_1418_n 0.00163615f $X=4.515 $Y=1.84
+ $X2=0 $Y2=0
cc_535 N_A_828_74#_M1008_d N_A_301_74#_c_1419_n 0.00284049f $X=4.515 $Y=1.84
+ $X2=0 $Y2=0
cc_536 N_A_828_74#_M1015_g N_A_301_74#_c_1419_n 0.00503824f $X=5.435 $Y=2.75
+ $X2=0 $Y2=0
cc_537 N_A_828_74#_c_560_n N_A_301_74#_c_1419_n 0.0227474f $X=5.12 $Y=2.215
+ $X2=0 $Y2=0
cc_538 N_A_828_74#_c_561_n N_A_301_74#_c_1419_n 0.00464433f $X=5.12 $Y=2.215
+ $X2=0 $Y2=0
cc_539 N_A_828_74#_M1008_d N_A_301_74#_c_1421_n 0.00503581f $X=4.515 $Y=1.84
+ $X2=0 $Y2=0
cc_540 N_A_828_74#_M1015_g N_A_301_74#_c_1421_n 0.00437377f $X=5.435 $Y=2.75
+ $X2=0 $Y2=0
cc_541 N_A_828_74#_c_560_n N_A_301_74#_c_1421_n 0.013477f $X=5.12 $Y=2.215 $X2=0
+ $Y2=0
cc_542 N_A_828_74#_c_537_n N_A_301_74#_c_1414_n 0.0276766f $X=4.28 $Y=0.515
+ $X2=0 $Y2=0
cc_543 N_A_828_74#_c_538_n N_A_301_74#_c_1414_n 0.0197906f $X=5.055 $Y=0.34
+ $X2=0 $Y2=0
cc_544 N_A_828_74#_c_540_n N_A_301_74#_c_1414_n 0.0124099f $X=5.14 $Y=2.05 $X2=0
+ $Y2=0
cc_545 N_A_828_74#_c_614_p N_VGND_M1024_d 0.0150959f $X=6.805 $Y=0.775 $X2=0
+ $Y2=0
cc_546 N_A_828_74#_c_630_p N_VGND_M1024_d 0.00439195f $X=6.89 $Y=0.69 $X2=0
+ $Y2=0
cc_547 N_A_828_74#_c_546_n N_VGND_M1024_d 6.26408e-19 $X=6.975 $Y=0.34 $X2=0
+ $Y2=0
cc_548 N_A_828_74#_c_539_n N_VGND_c_1558_n 0.0112234f $X=4.445 $Y=0.34 $X2=0
+ $Y2=0
cc_549 N_A_828_74#_c_541_n N_VGND_c_1559_n 0.00716007f $X=5.735 $Y=0.34 $X2=0
+ $Y2=0
cc_550 N_A_828_74#_c_542_n N_VGND_c_1559_n 0.00311855f $X=5.82 $Y=0.69 $X2=0
+ $Y2=0
cc_551 N_A_828_74#_c_614_p N_VGND_c_1559_n 0.0179784f $X=6.805 $Y=0.775 $X2=0
+ $Y2=0
cc_552 N_A_828_74#_c_630_p N_VGND_c_1559_n 0.00706899f $X=6.89 $Y=0.69 $X2=0
+ $Y2=0
cc_553 N_A_828_74#_c_546_n N_VGND_c_1559_n 0.0144033f $X=6.975 $Y=0.34 $X2=0
+ $Y2=0
cc_554 N_A_828_74#_c_536_n N_VGND_c_1567_n 7.26171e-19 $X=5.695 $Y=1.03 $X2=0
+ $Y2=0
cc_555 N_A_828_74#_c_538_n N_VGND_c_1567_n 0.0392369f $X=5.055 $Y=0.34 $X2=0
+ $Y2=0
cc_556 N_A_828_74#_c_539_n N_VGND_c_1567_n 0.0179217f $X=4.445 $Y=0.34 $X2=0
+ $Y2=0
cc_557 N_A_828_74#_c_541_n N_VGND_c_1567_n 0.0449818f $X=5.735 $Y=0.34 $X2=0
+ $Y2=0
cc_558 N_A_828_74#_c_614_p N_VGND_c_1567_n 0.00534483f $X=6.805 $Y=0.775 $X2=0
+ $Y2=0
cc_559 N_A_828_74#_c_549_n N_VGND_c_1567_n 0.0121867f $X=5.14 $Y=0.34 $X2=0
+ $Y2=0
cc_560 N_A_828_74#_c_715_p N_VGND_c_1567_n 0.00137281f $X=5.86 $Y=0.775 $X2=0
+ $Y2=0
cc_561 N_A_828_74#_c_614_p N_VGND_c_1568_n 0.00262318f $X=6.805 $Y=0.775 $X2=0
+ $Y2=0
cc_562 N_A_828_74#_c_545_n N_VGND_c_1568_n 0.0544154f $X=7.645 $Y=0.34 $X2=0
+ $Y2=0
cc_563 N_A_828_74#_c_546_n N_VGND_c_1568_n 0.0120795f $X=6.975 $Y=0.34 $X2=0
+ $Y2=0
cc_564 N_A_828_74#_c_553_n N_VGND_c_1568_n 0.00278271f $X=7.57 $Y=1.03 $X2=0
+ $Y2=0
cc_565 N_A_828_74#_c_538_n N_VGND_c_1571_n 0.0229266f $X=5.055 $Y=0.34 $X2=0
+ $Y2=0
cc_566 N_A_828_74#_c_539_n N_VGND_c_1571_n 0.00971942f $X=4.445 $Y=0.34 $X2=0
+ $Y2=0
cc_567 N_A_828_74#_c_541_n N_VGND_c_1571_n 0.025776f $X=5.735 $Y=0.34 $X2=0
+ $Y2=0
cc_568 N_A_828_74#_c_614_p N_VGND_c_1571_n 0.0165161f $X=6.805 $Y=0.775 $X2=0
+ $Y2=0
cc_569 N_A_828_74#_c_545_n N_VGND_c_1571_n 0.0304265f $X=7.645 $Y=0.34 $X2=0
+ $Y2=0
cc_570 N_A_828_74#_c_546_n N_VGND_c_1571_n 0.00658903f $X=6.975 $Y=0.34 $X2=0
+ $Y2=0
cc_571 N_A_828_74#_c_549_n N_VGND_c_1571_n 0.00660921f $X=5.14 $Y=0.34 $X2=0
+ $Y2=0
cc_572 N_A_828_74#_c_715_p N_VGND_c_1571_n 0.00232932f $X=5.86 $Y=0.775 $X2=0
+ $Y2=0
cc_573 N_A_828_74#_c_553_n N_VGND_c_1571_n 0.00358571f $X=7.57 $Y=1.03 $X2=0
+ $Y2=0
cc_574 N_A_828_74#_c_542_n A_1154_100# 0.00242668f $X=5.82 $Y=0.69 $X2=-0.19
+ $Y2=-0.245
cc_575 N_A_828_74#_c_543_n A_1154_100# 7.37711e-19 $X=5.82 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_576 N_A_828_74#_c_614_p A_1154_100# 0.00627545f $X=6.805 $Y=0.775 $X2=-0.19
+ $Y2=-0.245
cc_577 N_A_828_74#_c_715_p A_1154_100# 0.00184264f $X=5.86 $Y=0.775 $X2=-0.19
+ $Y2=-0.245
cc_578 N_A_630_74#_c_760_n N_A_1239_74#_M1016_d 0.0168685f $X=7.545 $Y=2.605
+ $X2=0 $Y2=0
cc_579 N_A_630_74#_M1013_g N_A_1239_74#_c_952_n 0.0434559f $X=5.935 $Y=2.75
+ $X2=0 $Y2=0
cc_580 N_A_630_74#_c_759_n N_A_1239_74#_c_952_n 0.00488263f $X=6.13 $Y=2.52
+ $X2=0 $Y2=0
cc_581 N_A_630_74#_c_760_n N_A_1239_74#_M1019_g 0.0184868f $X=7.545 $Y=2.605
+ $X2=0 $Y2=0
cc_582 N_A_630_74#_c_753_n N_A_1239_74#_c_945_n 0.0319501f $X=5.735 $Y=1.765
+ $X2=0 $Y2=0
cc_583 N_A_630_74#_M1013_g N_A_1239_74#_c_945_n 0.00473467f $X=5.935 $Y=2.75
+ $X2=0 $Y2=0
cc_584 N_A_630_74#_c_759_n N_A_1239_74#_c_945_n 0.00267751f $X=6.13 $Y=2.52
+ $X2=0 $Y2=0
cc_585 N_A_630_74#_c_763_n N_A_1239_74#_c_945_n 0.00821079f $X=6.13 $Y=2.035
+ $X2=0 $Y2=0
cc_586 N_A_630_74#_M1026_g N_A_1239_74#_c_955_n 9.98065e-19 $X=7.66 $Y=2.54
+ $X2=0 $Y2=0
cc_587 N_A_630_74#_c_760_n N_A_1239_74#_c_955_n 0.0234985f $X=7.545 $Y=2.605
+ $X2=0 $Y2=0
cc_588 N_A_630_74#_c_761_n N_A_1239_74#_c_955_n 0.0109032f $X=7.63 $Y=2.52 $X2=0
+ $Y2=0
cc_589 N_A_630_74#_M1026_g N_A_1239_74#_c_949_n 6.20776e-19 $X=7.66 $Y=2.54
+ $X2=0 $Y2=0
cc_590 N_A_630_74#_c_738_n N_A_1239_74#_c_949_n 0.00508347f $X=8.02 $Y=1.6 $X2=0
+ $Y2=0
cc_591 N_A_630_74#_c_761_n N_A_1239_74#_c_949_n 0.0103312f $X=7.63 $Y=2.52 $X2=0
+ $Y2=0
cc_592 N_A_630_74#_c_750_n N_A_1239_74#_c_949_n 0.021245f $X=7.735 $Y=1.765
+ $X2=0 $Y2=0
cc_593 N_A_630_74#_c_751_n N_A_1239_74#_c_949_n 0.00111668f $X=7.735 $Y=1.765
+ $X2=0 $Y2=0
cc_594 N_A_630_74#_M1026_g N_A_1018_100#_M1016_g 0.0218236f $X=7.66 $Y=2.54
+ $X2=0 $Y2=0
cc_595 N_A_630_74#_c_760_n N_A_1018_100#_M1016_g 0.0177366f $X=7.545 $Y=2.605
+ $X2=0 $Y2=0
cc_596 N_A_630_74#_M1007_g N_A_1018_100#_c_1023_n 0.002957f $X=5.015 $Y=0.71
+ $X2=0 $Y2=0
cc_597 N_A_630_74#_M1013_g N_A_1018_100#_c_1029_n 0.00792053f $X=5.935 $Y=2.75
+ $X2=0 $Y2=0
cc_598 N_A_630_74#_c_753_n N_A_1018_100#_c_1024_n 0.0139864f $X=5.735 $Y=1.765
+ $X2=0 $Y2=0
cc_599 N_A_630_74#_c_763_n N_A_1018_100#_c_1024_n 0.0354589f $X=6.13 $Y=2.035
+ $X2=0 $Y2=0
cc_600 N_A_630_74#_c_753_n N_A_1018_100#_c_1025_n 0.00440036f $X=5.735 $Y=1.765
+ $X2=0 $Y2=0
cc_601 N_A_630_74#_c_743_n N_A_1018_100#_c_1025_n 9.11089e-19 $X=5.015 $Y=1.555
+ $X2=0 $Y2=0
cc_602 N_A_630_74#_c_753_n N_A_1018_100#_c_1031_n 0.0127816f $X=5.735 $Y=1.765
+ $X2=0 $Y2=0
cc_603 N_A_630_74#_M1013_g N_A_1018_100#_c_1031_n 0.00134966f $X=5.935 $Y=2.75
+ $X2=0 $Y2=0
cc_604 N_A_630_74#_c_759_n N_A_1018_100#_c_1031_n 0.00618484f $X=6.13 $Y=2.52
+ $X2=0 $Y2=0
cc_605 N_A_630_74#_c_762_n N_A_1018_100#_c_1031_n 0.0029426f $X=5.9 $Y=2.035
+ $X2=0 $Y2=0
cc_606 N_A_630_74#_c_763_n N_A_1018_100#_c_1031_n 0.0254592f $X=6.13 $Y=2.035
+ $X2=0 $Y2=0
cc_607 N_A_630_74#_c_753_n N_A_1018_100#_c_1032_n 0.00284089f $X=5.735 $Y=1.765
+ $X2=0 $Y2=0
cc_608 N_A_630_74#_M1013_g N_A_1018_100#_c_1032_n 0.00451493f $X=5.935 $Y=2.75
+ $X2=0 $Y2=0
cc_609 N_A_630_74#_c_759_n N_A_1018_100#_c_1032_n 0.0115661f $X=6.13 $Y=2.52
+ $X2=0 $Y2=0
cc_610 N_A_630_74#_c_867_p N_A_1018_100#_c_1032_n 0.00730162f $X=6.215 $Y=2.605
+ $X2=0 $Y2=0
cc_611 N_A_630_74#_c_763_n N_A_1018_100#_c_1032_n 0.0114884f $X=6.13 $Y=2.035
+ $X2=0 $Y2=0
cc_612 N_A_630_74#_c_766_n N_A_1018_100#_c_1032_n 0.00278262f $X=5.9 $Y=2.2
+ $X2=0 $Y2=0
cc_613 N_A_630_74#_c_760_n N_A_1018_100#_c_1026_n 0.00819615f $X=7.545 $Y=2.605
+ $X2=0 $Y2=0
cc_614 N_A_630_74#_c_763_n N_A_1018_100#_c_1026_n 0.00240996f $X=6.13 $Y=2.035
+ $X2=0 $Y2=0
cc_615 N_A_630_74#_c_760_n N_A_1018_100#_c_1027_n 0.00105513f $X=7.545 $Y=2.605
+ $X2=0 $Y2=0
cc_616 N_A_630_74#_c_750_n N_A_1018_100#_c_1027_n 9.72318e-19 $X=7.735 $Y=1.765
+ $X2=0 $Y2=0
cc_617 N_A_630_74#_c_751_n N_A_1018_100#_c_1027_n 0.00907639f $X=7.735 $Y=1.765
+ $X2=0 $Y2=0
cc_618 N_A_630_74#_c_741_n N_A_1736_74#_c_1112_n 0.0202694f $X=8.365 $Y=1.015
+ $X2=0 $Y2=0
cc_619 N_A_630_74#_c_739_n N_A_1736_74#_c_1121_n 0.0202694f $X=8.29 $Y=1.09
+ $X2=0 $Y2=0
cc_620 N_A_630_74#_M1026_g N_A_1520_74#_c_1205_n 0.00293691f $X=7.66 $Y=2.54
+ $X2=0 $Y2=0
cc_621 N_A_630_74#_c_761_n N_A_1520_74#_c_1205_n 0.0239941f $X=7.63 $Y=2.52
+ $X2=0 $Y2=0
cc_622 N_A_630_74#_c_750_n N_A_1520_74#_c_1205_n 0.001265f $X=7.735 $Y=1.765
+ $X2=0 $Y2=0
cc_623 N_A_630_74#_c_751_n N_A_1520_74#_c_1205_n 0.00753796f $X=7.735 $Y=1.765
+ $X2=0 $Y2=0
cc_624 N_A_630_74#_M1026_g N_A_1520_74#_c_1206_n 0.0100066f $X=7.66 $Y=2.54
+ $X2=0 $Y2=0
cc_625 N_A_630_74#_c_760_n N_A_1520_74#_c_1206_n 0.0137305f $X=7.545 $Y=2.605
+ $X2=0 $Y2=0
cc_626 N_A_630_74#_c_761_n N_A_1520_74#_c_1206_n 0.00752589f $X=7.63 $Y=2.52
+ $X2=0 $Y2=0
cc_627 N_A_630_74#_c_738_n N_A_1520_74#_c_1199_n 0.00134724f $X=8.02 $Y=1.6
+ $X2=0 $Y2=0
cc_628 N_A_630_74#_c_739_n N_A_1520_74#_c_1202_n 0.00500602f $X=8.29 $Y=1.09
+ $X2=0 $Y2=0
cc_629 N_A_630_74#_c_740_n N_A_1520_74#_c_1202_n 0.00811832f $X=8.095 $Y=1.09
+ $X2=0 $Y2=0
cc_630 N_A_630_74#_c_741_n N_A_1520_74#_c_1202_n 0.0164162f $X=8.365 $Y=1.015
+ $X2=0 $Y2=0
cc_631 N_A_630_74#_c_757_n N_VPWR_M1008_s 0.00770541f $X=3.855 $Y=1.98 $X2=0
+ $Y2=0
cc_632 N_A_630_74#_c_760_n N_VPWR_M1019_d 0.00799866f $X=7.545 $Y=2.605 $X2=0
+ $Y2=0
cc_633 N_A_630_74#_M1008_g N_VPWR_c_1290_n 0.0169885f $X=4.425 $Y=2.4 $X2=0
+ $Y2=0
cc_634 N_A_630_74#_c_760_n N_VPWR_c_1291_n 0.0248918f $X=7.545 $Y=2.605 $X2=0
+ $Y2=0
cc_635 N_A_630_74#_M1008_g N_VPWR_c_1301_n 0.00460063f $X=4.425 $Y=2.4 $X2=0
+ $Y2=0
cc_636 N_A_630_74#_M1013_g N_VPWR_c_1301_n 0.005209f $X=5.935 $Y=2.75 $X2=0
+ $Y2=0
cc_637 N_A_630_74#_c_760_n N_VPWR_c_1301_n 0.00371686f $X=7.545 $Y=2.605 $X2=0
+ $Y2=0
cc_638 N_A_630_74#_c_867_p N_VPWR_c_1301_n 0.00259386f $X=6.215 $Y=2.605 $X2=0
+ $Y2=0
cc_639 N_A_630_74#_M1026_g N_VPWR_c_1302_n 0.00423418f $X=7.66 $Y=2.54 $X2=0
+ $Y2=0
cc_640 N_A_630_74#_c_760_n N_VPWR_c_1302_n 0.0141895f $X=7.545 $Y=2.605 $X2=0
+ $Y2=0
cc_641 N_A_630_74#_M1008_g N_VPWR_c_1287_n 0.00448128f $X=4.425 $Y=2.4 $X2=0
+ $Y2=0
cc_642 N_A_630_74#_M1013_g N_VPWR_c_1287_n 0.00983542f $X=5.935 $Y=2.75 $X2=0
+ $Y2=0
cc_643 N_A_630_74#_M1026_g N_VPWR_c_1287_n 0.00615705f $X=7.66 $Y=2.54 $X2=0
+ $Y2=0
cc_644 N_A_630_74#_c_760_n N_VPWR_c_1287_n 0.0325677f $X=7.545 $Y=2.605 $X2=0
+ $Y2=0
cc_645 N_A_630_74#_c_867_p N_VPWR_c_1287_n 0.00506366f $X=6.215 $Y=2.605 $X2=0
+ $Y2=0
cc_646 N_A_630_74#_c_746_n N_A_301_74#_c_1407_n 0.00504519f $X=3.455 $Y=0.875
+ $X2=0 $Y2=0
cc_647 N_A_630_74#_c_757_n N_A_301_74#_c_1410_n 0.0208559f $X=3.855 $Y=1.98
+ $X2=0 $Y2=0
cc_648 N_A_630_74#_c_757_n N_A_301_74#_c_1462_n 0.00209974f $X=3.855 $Y=1.98
+ $X2=0 $Y2=0
cc_649 N_A_630_74#_M1008_g N_A_301_74#_c_1417_n 0.0222436f $X=4.425 $Y=2.4 $X2=0
+ $Y2=0
cc_650 N_A_630_74#_c_743_n N_A_301_74#_c_1417_n 6.78967e-19 $X=5.015 $Y=1.555
+ $X2=0 $Y2=0
cc_651 N_A_630_74#_c_757_n N_A_301_74#_c_1417_n 0.0260964f $X=3.855 $Y=1.98
+ $X2=0 $Y2=0
cc_652 N_A_630_74#_c_747_n N_A_301_74#_c_1417_n 0.0128838f $X=3.955 $Y=1.465
+ $X2=0 $Y2=0
cc_653 N_A_630_74#_M1008_g N_A_301_74#_c_1411_n 0.00569613f $X=4.425 $Y=2.4
+ $X2=0 $Y2=0
cc_654 N_A_630_74#_c_736_n N_A_301_74#_c_1411_n 0.0165063f $X=4.94 $Y=1.555
+ $X2=0 $Y2=0
cc_655 N_A_630_74#_c_742_n N_A_301_74#_c_1411_n 0.00470969f $X=4.425 $Y=1.555
+ $X2=0 $Y2=0
cc_656 N_A_630_74#_c_734_n N_A_301_74#_c_1412_n 0.00679719f $X=4.335 $Y=1.555
+ $X2=0 $Y2=0
cc_657 N_A_630_74#_M1008_g N_A_301_74#_c_1412_n 4.2037e-19 $X=4.425 $Y=2.4 $X2=0
+ $Y2=0
cc_658 N_A_630_74#_c_742_n N_A_301_74#_c_1412_n 0.0010724f $X=4.425 $Y=1.555
+ $X2=0 $Y2=0
cc_659 N_A_630_74#_c_747_n N_A_301_74#_c_1412_n 0.0130528f $X=3.955 $Y=1.465
+ $X2=0 $Y2=0
cc_660 N_A_630_74#_M1018_g N_A_301_74#_c_1413_n 0.00628173f $X=4.065 $Y=0.74
+ $X2=0 $Y2=0
cc_661 N_A_630_74#_M1007_g N_A_301_74#_c_1413_n 0.0111103f $X=5.015 $Y=0.71
+ $X2=0 $Y2=0
cc_662 N_A_630_74#_c_779_n N_A_301_74#_c_1413_n 0.00527653f $X=3.955 $Y=1.4
+ $X2=0 $Y2=0
cc_663 N_A_630_74#_c_749_n N_A_301_74#_c_1413_n 0.00474003f $X=3.955 $Y=1.3
+ $X2=0 $Y2=0
cc_664 N_A_630_74#_M1008_g N_A_301_74#_c_1418_n 0.00568905f $X=4.425 $Y=2.4
+ $X2=0 $Y2=0
cc_665 N_A_630_74#_M1004_d N_A_301_74#_c_1421_n 0.00819631f $X=3.325 $Y=1.84
+ $X2=0 $Y2=0
cc_666 N_A_630_74#_M1008_g N_A_301_74#_c_1421_n 0.0231562f $X=4.425 $Y=2.4 $X2=0
+ $Y2=0
cc_667 N_A_630_74#_c_757_n N_A_301_74#_c_1421_n 0.0547723f $X=3.855 $Y=1.98
+ $X2=0 $Y2=0
cc_668 N_A_630_74#_c_748_n N_A_301_74#_c_1421_n 0.00494605f $X=3.955 $Y=1.465
+ $X2=0 $Y2=0
cc_669 N_A_630_74#_c_736_n N_A_301_74#_c_1414_n 0.00201345f $X=4.94 $Y=1.555
+ $X2=0 $Y2=0
cc_670 N_A_630_74#_M1007_g N_A_301_74#_c_1414_n 4.19896e-19 $X=5.015 $Y=0.71
+ $X2=0 $Y2=0
cc_671 N_A_630_74#_c_867_p A_1205_508# 0.00192409f $X=6.215 $Y=2.605 $X2=-0.19
+ $Y2=-0.245
cc_672 N_A_630_74#_c_745_n N_VGND_M1018_s 0.0074763f $X=3.855 $Y=0.875 $X2=0
+ $Y2=0
cc_673 N_A_630_74#_c_749_n N_VGND_M1018_s 0.00568518f $X=3.955 $Y=1.3 $X2=0
+ $Y2=0
cc_674 N_A_630_74#_c_744_n N_VGND_c_1557_n 0.0164209f $X=3.29 $Y=0.515 $X2=0
+ $Y2=0
cc_675 N_A_630_74#_M1018_g N_VGND_c_1558_n 0.00796029f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_676 N_A_630_74#_c_744_n N_VGND_c_1558_n 0.018203f $X=3.29 $Y=0.515 $X2=0
+ $Y2=0
cc_677 N_A_630_74#_c_745_n N_VGND_c_1558_n 0.0222318f $X=3.855 $Y=0.875 $X2=0
+ $Y2=0
cc_678 N_A_630_74#_c_748_n N_VGND_c_1558_n 4.14752e-19 $X=3.955 $Y=1.465 $X2=0
+ $Y2=0
cc_679 N_A_630_74#_c_741_n N_VGND_c_1560_n 0.00138935f $X=8.365 $Y=1.015 $X2=0
+ $Y2=0
cc_680 N_A_630_74#_c_744_n N_VGND_c_1564_n 0.0144497f $X=3.29 $Y=0.515 $X2=0
+ $Y2=0
cc_681 N_A_630_74#_M1018_g N_VGND_c_1567_n 0.00383152f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_682 N_A_630_74#_M1007_g N_VGND_c_1567_n 7.26171e-19 $X=5.015 $Y=0.71 $X2=0
+ $Y2=0
cc_683 N_A_630_74#_c_741_n N_VGND_c_1568_n 0.00466611f $X=8.365 $Y=1.015 $X2=0
+ $Y2=0
cc_684 N_A_630_74#_M1018_g N_VGND_c_1571_n 0.00728991f $X=4.065 $Y=0.74 $X2=0
+ $Y2=0
cc_685 N_A_630_74#_c_741_n N_VGND_c_1571_n 0.00505379f $X=8.365 $Y=1.015 $X2=0
+ $Y2=0
cc_686 N_A_630_74#_c_744_n N_VGND_c_1571_n 0.0119539f $X=3.29 $Y=0.515 $X2=0
+ $Y2=0
cc_687 N_A_630_74#_c_745_n N_VGND_c_1571_n 0.00989205f $X=3.855 $Y=0.875 $X2=0
+ $Y2=0
cc_688 N_A_1239_74#_c_945_n N_A_1018_100#_M1016_g 0.0305229f $X=6.335 $Y=2.315
+ $X2=0 $Y2=0
cc_689 N_A_1239_74#_c_955_n N_A_1018_100#_M1016_g 0.00748671f $X=7.195 $Y=2.265
+ $X2=0 $Y2=0
cc_690 N_A_1239_74#_c_949_n N_A_1018_100#_M1016_g 0.00431208f $X=7.195 $Y=2.1
+ $X2=0 $Y2=0
cc_691 N_A_1239_74#_c_945_n N_A_1018_100#_M1011_g 0.00521383f $X=6.335 $Y=2.315
+ $X2=0 $Y2=0
cc_692 N_A_1239_74#_c_946_n N_A_1018_100#_M1011_g 0.0192641f $X=7.145 $Y=1.195
+ $X2=0 $Y2=0
cc_693 N_A_1239_74#_c_947_n N_A_1018_100#_M1011_g 0.00662294f $X=6.36 $Y=1.195
+ $X2=0 $Y2=0
cc_694 N_A_1239_74#_c_948_n N_A_1018_100#_M1011_g 0.00782995f $X=7.23 $Y=1.03
+ $X2=0 $Y2=0
cc_695 N_A_1239_74#_c_949_n N_A_1018_100#_M1011_g 0.0115886f $X=7.195 $Y=2.1
+ $X2=0 $Y2=0
cc_696 N_A_1239_74#_c_967_n N_A_1018_100#_M1011_g 0.00298439f $X=7.31 $Y=0.685
+ $X2=0 $Y2=0
cc_697 N_A_1239_74#_c_950_n N_A_1018_100#_M1011_g 0.0027421f $X=7.23 $Y=1.195
+ $X2=0 $Y2=0
cc_698 N_A_1239_74#_c_951_n N_A_1018_100#_M1011_g 0.00857377f $X=6.36 $Y=1.03
+ $X2=0 $Y2=0
cc_699 N_A_1239_74#_M1019_g N_A_1018_100#_c_1029_n 0.00116915f $X=6.335 $Y=2.75
+ $X2=0 $Y2=0
cc_700 N_A_1239_74#_c_952_n N_A_1018_100#_c_1024_n 7.85116e-19 $X=6.335 $Y=2.405
+ $X2=0 $Y2=0
cc_701 N_A_1239_74#_c_945_n N_A_1018_100#_c_1024_n 0.0168872f $X=6.335 $Y=2.315
+ $X2=0 $Y2=0
cc_702 N_A_1239_74#_c_946_n N_A_1018_100#_c_1024_n 0.0337543f $X=7.145 $Y=1.195
+ $X2=0 $Y2=0
cc_703 N_A_1239_74#_c_947_n N_A_1018_100#_c_1024_n 0.00435089f $X=6.36 $Y=1.195
+ $X2=0 $Y2=0
cc_704 N_A_1239_74#_c_945_n N_A_1018_100#_c_1026_n 0.00151695f $X=6.335 $Y=2.315
+ $X2=0 $Y2=0
cc_705 N_A_1239_74#_c_946_n N_A_1018_100#_c_1026_n 0.0278385f $X=7.145 $Y=1.195
+ $X2=0 $Y2=0
cc_706 N_A_1239_74#_c_949_n N_A_1018_100#_c_1026_n 0.0288169f $X=7.195 $Y=2.1
+ $X2=0 $Y2=0
cc_707 N_A_1239_74#_c_945_n N_A_1018_100#_c_1027_n 0.0204867f $X=6.335 $Y=2.315
+ $X2=0 $Y2=0
cc_708 N_A_1239_74#_c_946_n N_A_1018_100#_c_1027_n 0.00369837f $X=7.145 $Y=1.195
+ $X2=0 $Y2=0
cc_709 N_A_1239_74#_c_955_n N_A_1018_100#_c_1027_n 0.00431986f $X=7.195 $Y=2.265
+ $X2=0 $Y2=0
cc_710 N_A_1239_74#_c_949_n N_A_1018_100#_c_1027_n 0.00879068f $X=7.195 $Y=2.1
+ $X2=0 $Y2=0
cc_711 N_A_1239_74#_M1019_g N_VPWR_c_1291_n 0.0041537f $X=6.335 $Y=2.75 $X2=0
+ $Y2=0
cc_712 N_A_1239_74#_M1019_g N_VPWR_c_1301_n 0.00392086f $X=6.335 $Y=2.75 $X2=0
+ $Y2=0
cc_713 N_A_1239_74#_M1019_g N_VPWR_c_1287_n 0.00496594f $X=6.335 $Y=2.75 $X2=0
+ $Y2=0
cc_714 N_A_1239_74#_c_951_n N_VGND_c_1559_n 0.00231554f $X=6.36 $Y=1.03 $X2=0
+ $Y2=0
cc_715 N_A_1239_74#_c_951_n N_VGND_c_1567_n 0.00378853f $X=6.36 $Y=1.03 $X2=0
+ $Y2=0
cc_716 N_A_1239_74#_c_951_n N_VGND_c_1571_n 0.00505379f $X=6.36 $Y=1.03 $X2=0
+ $Y2=0
cc_717 N_A_1018_100#_M1016_g N_VPWR_c_1291_n 0.00440778f $X=6.955 $Y=2.54 $X2=0
+ $Y2=0
cc_718 N_A_1018_100#_c_1029_n N_VPWR_c_1291_n 0.00189455f $X=5.71 $Y=2.75 $X2=0
+ $Y2=0
cc_719 N_A_1018_100#_c_1029_n N_VPWR_c_1301_n 0.0144416f $X=5.71 $Y=2.75 $X2=0
+ $Y2=0
cc_720 N_A_1018_100#_M1016_g N_VPWR_c_1302_n 0.00392086f $X=6.955 $Y=2.54 $X2=0
+ $Y2=0
cc_721 N_A_1018_100#_M1016_g N_VPWR_c_1287_n 0.00499039f $X=6.955 $Y=2.54 $X2=0
+ $Y2=0
cc_722 N_A_1018_100#_c_1029_n N_VPWR_c_1287_n 0.0119324f $X=5.71 $Y=2.75 $X2=0
+ $Y2=0
cc_723 N_A_1018_100#_c_1032_n N_VPWR_c_1287_n 0.00511545f $X=5.635 $Y=2.54 $X2=0
+ $Y2=0
cc_724 N_A_1018_100#_c_1029_n N_A_301_74#_c_1419_n 0.0120413f $X=5.71 $Y=2.75
+ $X2=0 $Y2=0
cc_725 N_A_1018_100#_M1011_g N_VGND_c_1559_n 0.00121379f $X=7.09 $Y=0.645 $X2=0
+ $Y2=0
cc_726 N_A_1018_100#_M1011_g N_VGND_c_1568_n 0.00278271f $X=7.09 $Y=0.645 $X2=0
+ $Y2=0
cc_727 N_A_1018_100#_M1011_g N_VGND_c_1571_n 0.00358571f $X=7.09 $Y=0.645 $X2=0
+ $Y2=0
cc_728 N_A_1736_74#_c_1122_n N_A_1520_74#_M1031_g 0.0110928f $X=8.785 $Y=2.465
+ $X2=0 $Y2=0
cc_729 N_A_1736_74#_c_1113_n N_A_1520_74#_M1031_g 0.0152056f $X=8.95 $Y=2.315
+ $X2=0 $Y2=0
cc_730 N_A_1736_74#_c_1126_n N_A_1520_74#_M1031_g 0.0256958f $X=9.755 $Y=2.265
+ $X2=0 $Y2=0
cc_731 N_A_1736_74#_c_1127_n N_A_1520_74#_M1031_g 0.00606936f $X=9.762 $Y=2.1
+ $X2=0 $Y2=0
cc_732 N_A_1736_74#_c_1112_n N_A_1520_74#_M1009_g 0.00620125f $X=8.755 $Y=1.015
+ $X2=0 $Y2=0
cc_733 N_A_1736_74#_c_1113_n N_A_1520_74#_M1009_g 0.00602362f $X=8.95 $Y=2.315
+ $X2=0 $Y2=0
cc_734 N_A_1736_74#_c_1116_n N_A_1520_74#_M1009_g 0.0167285f $X=10.45 $Y=1.485
+ $X2=0 $Y2=0
cc_735 N_A_1736_74#_c_1118_n N_A_1520_74#_M1009_g 0.0163877f $X=9.65 $Y=1.195
+ $X2=0 $Y2=0
cc_736 N_A_1736_74#_c_1119_n N_A_1520_74#_M1009_g 0.0201251f $X=9.815 $Y=0.645
+ $X2=0 $Y2=0
cc_737 N_A_1736_74#_c_1120_n N_A_1520_74#_M1009_g 0.0152668f $X=9.85 $Y=1.65
+ $X2=0 $Y2=0
cc_738 N_A_1736_74#_c_1121_n N_A_1520_74#_M1009_g 0.0223769f $X=8.95 $Y=1.187
+ $X2=0 $Y2=0
cc_739 N_A_1736_74#_c_1113_n N_A_1520_74#_c_1207_n 0.00258749f $X=8.95 $Y=2.315
+ $X2=0 $Y2=0
cc_740 N_A_1736_74#_c_1125_n N_A_1520_74#_c_1207_n 0.0170478f $X=8.95 $Y=2.39
+ $X2=0 $Y2=0
cc_741 N_A_1736_74#_c_1113_n N_A_1520_74#_c_1199_n 0.00673107f $X=8.95 $Y=2.315
+ $X2=0 $Y2=0
cc_742 N_A_1736_74#_c_1118_n N_A_1520_74#_c_1199_n 0.0158866f $X=9.65 $Y=1.195
+ $X2=0 $Y2=0
cc_743 N_A_1736_74#_c_1121_n N_A_1520_74#_c_1199_n 0.010589f $X=8.95 $Y=1.187
+ $X2=0 $Y2=0
cc_744 N_A_1736_74#_c_1113_n N_A_1520_74#_c_1208_n 0.00849239f $X=8.95 $Y=2.315
+ $X2=0 $Y2=0
cc_745 N_A_1736_74#_c_1113_n N_A_1520_74#_c_1200_n 0.0190414f $X=8.95 $Y=2.315
+ $X2=0 $Y2=0
cc_746 N_A_1736_74#_c_1118_n N_A_1520_74#_c_1200_n 0.0319279f $X=9.65 $Y=1.195
+ $X2=0 $Y2=0
cc_747 N_A_1736_74#_c_1120_n N_A_1520_74#_c_1200_n 0.00425106f $X=9.85 $Y=1.65
+ $X2=0 $Y2=0
cc_748 N_A_1736_74#_c_1127_n N_A_1520_74#_c_1200_n 0.0222566f $X=9.762 $Y=2.1
+ $X2=0 $Y2=0
cc_749 N_A_1736_74#_c_1121_n N_A_1520_74#_c_1200_n 0.00609519f $X=8.95 $Y=1.187
+ $X2=0 $Y2=0
cc_750 N_A_1736_74#_c_1113_n N_A_1520_74#_c_1201_n 0.018115f $X=8.95 $Y=2.315
+ $X2=0 $Y2=0
cc_751 N_A_1736_74#_c_1118_n N_A_1520_74#_c_1201_n 0.00507668f $X=9.65 $Y=1.195
+ $X2=0 $Y2=0
cc_752 N_A_1736_74#_c_1126_n N_A_1520_74#_c_1201_n 0.0026612f $X=9.755 $Y=2.265
+ $X2=0 $Y2=0
cc_753 N_A_1736_74#_c_1127_n N_A_1520_74#_c_1201_n 0.00722473f $X=9.762 $Y=2.1
+ $X2=0 $Y2=0
cc_754 N_A_1736_74#_c_1121_n N_A_1520_74#_c_1201_n 0.00259706f $X=8.95 $Y=1.187
+ $X2=0 $Y2=0
cc_755 N_A_1736_74#_c_1112_n N_A_1520_74#_c_1202_n 0.0132051f $X=8.755 $Y=1.015
+ $X2=0 $Y2=0
cc_756 N_A_1736_74#_c_1118_n N_A_1520_74#_c_1202_n 0.00982098f $X=9.65 $Y=1.195
+ $X2=0 $Y2=0
cc_757 N_A_1736_74#_c_1121_n N_A_1520_74#_c_1202_n 0.00873734f $X=8.95 $Y=1.187
+ $X2=0 $Y2=0
cc_758 N_A_1736_74#_c_1113_n N_A_1520_74#_c_1203_n 0.00274855f $X=8.95 $Y=2.315
+ $X2=0 $Y2=0
cc_759 N_A_1736_74#_c_1122_n N_VPWR_c_1292_n 0.0178456f $X=8.785 $Y=2.465 $X2=0
+ $Y2=0
cc_760 N_A_1736_74#_c_1125_n N_VPWR_c_1292_n 0.00578442f $X=8.95 $Y=2.39 $X2=0
+ $Y2=0
cc_761 N_A_1736_74#_c_1126_n N_VPWR_c_1292_n 0.0133266f $X=9.755 $Y=2.265 $X2=0
+ $Y2=0
cc_762 N_A_1736_74#_M1001_g N_VPWR_c_1293_n 0.00649215f $X=10.54 $Y=2.4 $X2=0
+ $Y2=0
cc_763 N_A_1736_74#_c_1116_n N_VPWR_c_1293_n 0.0053894f $X=10.45 $Y=1.485 $X2=0
+ $Y2=0
cc_764 N_A_1736_74#_c_1120_n N_VPWR_c_1293_n 0.00796601f $X=9.85 $Y=1.65 $X2=0
+ $Y2=0
cc_765 N_A_1736_74#_c_1127_n N_VPWR_c_1293_n 0.0794555f $X=9.762 $Y=2.1 $X2=0
+ $Y2=0
cc_766 N_A_1736_74#_c_1126_n N_VPWR_c_1298_n 0.0152183f $X=9.755 $Y=2.265 $X2=0
+ $Y2=0
cc_767 N_A_1736_74#_c_1122_n N_VPWR_c_1302_n 0.00460063f $X=8.785 $Y=2.465 $X2=0
+ $Y2=0
cc_768 N_A_1736_74#_M1001_g N_VPWR_c_1303_n 0.005209f $X=10.54 $Y=2.4 $X2=0
+ $Y2=0
cc_769 N_A_1736_74#_c_1122_n N_VPWR_c_1287_n 0.00908371f $X=8.785 $Y=2.465 $X2=0
+ $Y2=0
cc_770 N_A_1736_74#_M1001_g N_VPWR_c_1287_n 0.00991123f $X=10.54 $Y=2.4 $X2=0
+ $Y2=0
cc_771 N_A_1736_74#_c_1126_n N_VPWR_c_1287_n 0.0125283f $X=9.755 $Y=2.265 $X2=0
+ $Y2=0
cc_772 N_A_1736_74#_M1001_g Q 0.0239605f $X=10.54 $Y=2.4 $X2=0 $Y2=0
cc_773 N_A_1736_74#_M1017_g Q 0.0180582f $X=10.555 $Y=0.76 $X2=0 $Y2=0
cc_774 N_A_1736_74#_c_1117_n Q 0.0145147f $X=10.54 $Y=1.485 $X2=0 $Y2=0
cc_775 N_A_1736_74#_c_1120_n Q 0.0196039f $X=9.85 $Y=1.65 $X2=0 $Y2=0
cc_776 N_A_1736_74#_c_1127_n Q 0.00448272f $X=9.762 $Y=2.1 $X2=0 $Y2=0
cc_777 N_A_1736_74#_c_1112_n N_VGND_c_1560_n 0.0108466f $X=8.755 $Y=1.015 $X2=0
+ $Y2=0
cc_778 N_A_1736_74#_c_1118_n N_VGND_c_1560_n 0.0283129f $X=9.65 $Y=1.195 $X2=0
+ $Y2=0
cc_779 N_A_1736_74#_c_1119_n N_VGND_c_1560_n 0.018141f $X=9.815 $Y=0.645 $X2=0
+ $Y2=0
cc_780 N_A_1736_74#_c_1121_n N_VGND_c_1560_n 0.013912f $X=8.95 $Y=1.187 $X2=0
+ $Y2=0
cc_781 N_A_1736_74#_M1017_g N_VGND_c_1561_n 0.00650419f $X=10.555 $Y=0.76 $X2=0
+ $Y2=0
cc_782 N_A_1736_74#_c_1116_n N_VGND_c_1561_n 0.00630256f $X=10.45 $Y=1.485 $X2=0
+ $Y2=0
cc_783 N_A_1736_74#_c_1119_n N_VGND_c_1561_n 0.0503224f $X=9.815 $Y=0.645 $X2=0
+ $Y2=0
cc_784 N_A_1736_74#_c_1120_n N_VGND_c_1561_n 0.015294f $X=9.85 $Y=1.65 $X2=0
+ $Y2=0
cc_785 N_A_1736_74#_c_1112_n N_VGND_c_1568_n 0.00405273f $X=8.755 $Y=1.015 $X2=0
+ $Y2=0
cc_786 N_A_1736_74#_c_1119_n N_VGND_c_1569_n 0.0145639f $X=9.815 $Y=0.645 $X2=0
+ $Y2=0
cc_787 N_A_1736_74#_M1017_g N_VGND_c_1570_n 0.00532065f $X=10.555 $Y=0.76 $X2=0
+ $Y2=0
cc_788 N_A_1736_74#_c_1112_n N_VGND_c_1571_n 0.00424518f $X=8.755 $Y=1.015 $X2=0
+ $Y2=0
cc_789 N_A_1736_74#_M1017_g N_VGND_c_1571_n 0.00539454f $X=10.555 $Y=0.76 $X2=0
+ $Y2=0
cc_790 N_A_1736_74#_c_1119_n N_VGND_c_1571_n 0.0119984f $X=9.815 $Y=0.645 $X2=0
+ $Y2=0
cc_791 N_A_1520_74#_M1031_g N_VPWR_c_1292_n 0.00671754f $X=9.53 $Y=2.54 $X2=0
+ $Y2=0
cc_792 N_A_1520_74#_c_1207_n N_VPWR_c_1292_n 0.00254192f $X=8.725 $Y=2.33 $X2=0
+ $Y2=0
cc_793 N_A_1520_74#_M1031_g N_VPWR_c_1293_n 0.00450661f $X=9.53 $Y=2.54 $X2=0
+ $Y2=0
cc_794 N_A_1520_74#_M1031_g N_VPWR_c_1298_n 0.005209f $X=9.53 $Y=2.54 $X2=0
+ $Y2=0
cc_795 N_A_1520_74#_c_1206_n N_VPWR_c_1302_n 0.011066f $X=7.97 $Y=2.815 $X2=0
+ $Y2=0
cc_796 N_A_1520_74#_M1031_g N_VPWR_c_1287_n 0.00989015f $X=9.53 $Y=2.54 $X2=0
+ $Y2=0
cc_797 N_A_1520_74#_c_1206_n N_VPWR_c_1287_n 0.00915947f $X=7.97 $Y=2.815 $X2=0
+ $Y2=0
cc_798 N_A_1520_74#_M1009_g N_VGND_c_1560_n 0.00949323f $X=9.6 $Y=0.645 $X2=0
+ $Y2=0
cc_799 N_A_1520_74#_c_1202_n N_VGND_c_1560_n 0.017907f $X=8.15 $Y=0.71 $X2=0
+ $Y2=0
cc_800 N_A_1520_74#_M1009_g N_VGND_c_1561_n 0.00488821f $X=9.6 $Y=0.645 $X2=0
+ $Y2=0
cc_801 N_A_1520_74#_c_1202_n N_VGND_c_1568_n 0.00929885f $X=8.15 $Y=0.71 $X2=0
+ $Y2=0
cc_802 N_A_1520_74#_M1009_g N_VGND_c_1569_n 0.00434272f $X=9.6 $Y=0.645 $X2=0
+ $Y2=0
cc_803 N_A_1520_74#_M1009_g N_VGND_c_1571_n 0.00830058f $X=9.6 $Y=0.645 $X2=0
+ $Y2=0
cc_804 N_A_1520_74#_c_1202_n N_VGND_c_1571_n 0.0207933f $X=8.15 $Y=0.71 $X2=0
+ $Y2=0
cc_805 N_A_1520_74#_c_1202_n A_1688_100# 0.00353421f $X=8.15 $Y=0.71 $X2=-0.19
+ $Y2=-0.245
cc_806 N_VPWR_M1002_d N_A_301_74#_c_1415_n 0.00402448f $X=2.615 $Y=2.32 $X2=0
+ $Y2=0
cc_807 N_VPWR_c_1289_n N_A_301_74#_c_1415_n 0.0189203f $X=2.92 $Y=2.815 $X2=0
+ $Y2=0
cc_808 N_VPWR_c_1287_n N_A_301_74#_c_1415_n 0.0239379f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_809 N_VPWR_M1002_d N_A_301_74#_c_1410_n 0.0123482f $X=2.615 $Y=2.32 $X2=0
+ $Y2=0
cc_810 N_VPWR_M1002_d N_A_301_74#_c_1462_n 3.40545e-19 $X=2.615 $Y=2.32 $X2=0
+ $Y2=0
cc_811 N_VPWR_c_1289_n N_A_301_74#_c_1462_n 0.00276502f $X=2.92 $Y=2.815 $X2=0
+ $Y2=0
cc_812 N_VPWR_c_1287_n N_A_301_74#_c_1462_n 0.00504989f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_813 N_VPWR_M1008_s N_A_301_74#_c_1417_n 0.00963735f $X=3.875 $Y=1.84 $X2=0
+ $Y2=0
cc_814 N_VPWR_c_1290_n N_A_301_74#_c_1418_n 0.0109597f $X=4.11 $Y=2.815 $X2=0
+ $Y2=0
cc_815 N_VPWR_c_1301_n N_A_301_74#_c_1418_n 0.00750764f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_816 N_VPWR_c_1287_n N_A_301_74#_c_1418_n 0.00624857f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_817 N_VPWR_c_1301_n N_A_301_74#_c_1419_n 0.0277877f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_818 N_VPWR_c_1287_n N_A_301_74#_c_1419_n 0.023859f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_819 N_VPWR_c_1288_n N_A_301_74#_c_1420_n 0.0197668f $X=0.89 $Y=2.465 $X2=0
+ $Y2=0
cc_820 N_VPWR_c_1296_n N_A_301_74#_c_1420_n 0.0144468f $X=2.67 $Y=3.33 $X2=0
+ $Y2=0
cc_821 N_VPWR_c_1287_n N_A_301_74#_c_1420_n 0.0118283f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_822 N_VPWR_M1002_d N_A_301_74#_c_1527_n 0.00234998f $X=2.615 $Y=2.32 $X2=0
+ $Y2=0
cc_823 N_VPWR_c_1289_n N_A_301_74#_c_1527_n 0.0148861f $X=2.92 $Y=2.815 $X2=0
+ $Y2=0
cc_824 N_VPWR_c_1287_n N_A_301_74#_c_1527_n 6.0606e-19 $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_825 N_VPWR_M1008_s N_A_301_74#_c_1421_n 0.0130906f $X=3.875 $Y=1.84 $X2=0
+ $Y2=0
cc_826 N_VPWR_c_1290_n N_A_301_74#_c_1421_n 0.0371625f $X=4.11 $Y=2.815 $X2=0
+ $Y2=0
cc_827 N_VPWR_c_1287_n N_A_301_74#_c_1421_n 0.0267352f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_828 N_VPWR_c_1293_n Q 0.0396567f $X=10.315 $Y=1.985 $X2=0 $Y2=0
cc_829 N_VPWR_c_1303_n Q 0.0147721f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_830 N_VPWR_c_1287_n Q 0.0121589f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_831 N_VPWR_c_1293_n N_VGND_c_1561_n 0.00541092f $X=10.315 $Y=1.985 $X2=0
+ $Y2=0
cc_832 N_A_301_74#_c_1415_n A_415_464# 0.00498776f $X=2.91 $Y=2.395 $X2=-0.19
+ $Y2=-0.245
cc_833 N_A_301_74#_c_1422_n N_VGND_c_1557_n 0.0242843f $X=2.42 $Y=0.565 $X2=0
+ $Y2=0
cc_834 N_A_301_74#_c_1407_n N_VGND_c_1557_n 0.0039147f $X=2.505 $Y=1.13 $X2=0
+ $Y2=0
cc_835 N_A_301_74#_c_1408_n N_VGND_c_1557_n 0.0085837f $X=2.91 $Y=1.215 $X2=0
+ $Y2=0
cc_836 N_A_301_74#_c_1422_n N_VGND_c_1562_n 0.0341166f $X=2.42 $Y=0.565 $X2=0
+ $Y2=0
cc_837 N_A_301_74#_c_1422_n N_VGND_c_1571_n 0.0373562f $X=2.42 $Y=0.565 $X2=0
+ $Y2=0
cc_838 N_A_301_74#_c_1422_n A_450_74# 0.00622173f $X=2.42 $Y=0.565 $X2=-0.19
+ $Y2=-0.245
cc_839 N_A_301_74#_c_1407_n A_450_74# 6.84302e-19 $X=2.505 $Y=1.13 $X2=-0.19
+ $Y2=-0.245
cc_840 Q N_VGND_c_1561_n 0.0301457f $X=10.715 $Y=0.47 $X2=0 $Y2=0
cc_841 Q N_VGND_c_1570_n 0.0136693f $X=10.715 $Y=0.47 $X2=0 $Y2=0
cc_842 Q N_VGND_c_1571_n 0.0121248f $X=10.715 $Y=0.47 $X2=0 $Y2=0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or2_4 A B VGND VNB VPB VPWR X
X0 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X2 VPWR A a_496_388# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X3 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 X a_83_260# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 a_83_260# B a_496_388# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X6 VGND A a_83_260# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_83_260# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_496_388# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X9 X a_83_260# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X11 VPWR a_83_260# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X12 a_496_388# B a_83_260# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X13 VGND a_83_260# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

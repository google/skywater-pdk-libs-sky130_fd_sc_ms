* File: sky130_fd_sc_ms__a32o_2.pxi.spice
* Created: Fri Aug 28 17:07:59 2020
* 
x_PM_SKY130_FD_SC_MS__A32O_2%A_45_264# N_A_45_264#_M1011_d N_A_45_264#_M1001_d
+ N_A_45_264#_M1004_g N_A_45_264#_M1003_g N_A_45_264#_M1005_g
+ N_A_45_264#_M1009_g N_A_45_264#_c_79_n N_A_45_264#_c_91_p N_A_45_264#_c_125_p
+ N_A_45_264#_c_80_n N_A_45_264#_c_93_p N_A_45_264#_c_81_n N_A_45_264#_c_82_n
+ N_A_45_264#_c_94_p N_A_45_264#_c_83_n N_A_45_264#_c_84_n N_A_45_264#_c_130_p
+ N_A_45_264#_c_122_p N_A_45_264#_c_85_n PM_SKY130_FD_SC_MS__A32O_2%A_45_264#
x_PM_SKY130_FD_SC_MS__A32O_2%A3 N_A3_M1010_g N_A3_M1007_g A3 N_A3_c_192_n
+ N_A3_c_193_n PM_SKY130_FD_SC_MS__A32O_2%A3
x_PM_SKY130_FD_SC_MS__A32O_2%A2 N_A2_M1006_g N_A2_M1012_g A2 N_A2_c_228_n
+ N_A2_c_229_n PM_SKY130_FD_SC_MS__A32O_2%A2
x_PM_SKY130_FD_SC_MS__A32O_2%A1 N_A1_M1011_g N_A1_M1000_g A1 N_A1_c_263_n
+ N_A1_c_264_n PM_SKY130_FD_SC_MS__A32O_2%A1
x_PM_SKY130_FD_SC_MS__A32O_2%B1 N_B1_M1002_g N_B1_M1001_g B1 N_B1_c_303_n
+ PM_SKY130_FD_SC_MS__A32O_2%B1
x_PM_SKY130_FD_SC_MS__A32O_2%B2 N_B2_M1008_g N_B2_M1013_g B2 N_B2_c_339_n
+ N_B2_c_340_n PM_SKY130_FD_SC_MS__A32O_2%B2
x_PM_SKY130_FD_SC_MS__A32O_2%VPWR N_VPWR_M1004_s N_VPWR_M1005_s N_VPWR_M1012_d
+ N_VPWR_c_362_n N_VPWR_c_363_n N_VPWR_c_364_n N_VPWR_c_365_n VPWR
+ N_VPWR_c_366_n N_VPWR_c_367_n N_VPWR_c_368_n N_VPWR_c_361_n N_VPWR_c_370_n
+ N_VPWR_c_371_n PM_SKY130_FD_SC_MS__A32O_2%VPWR
x_PM_SKY130_FD_SC_MS__A32O_2%X N_X_M1003_s N_X_M1004_d N_X_c_416_n N_X_c_417_n X
+ N_X_c_418_n PM_SKY130_FD_SC_MS__A32O_2%X
x_PM_SKY130_FD_SC_MS__A32O_2%A_349_368# N_A_349_368#_M1010_d
+ N_A_349_368#_M1000_d N_A_349_368#_M1013_d N_A_349_368#_c_453_n
+ N_A_349_368#_c_454_n N_A_349_368#_c_462_n N_A_349_368#_c_447_n
+ N_A_349_368#_c_448_n N_A_349_368#_c_449_n N_A_349_368#_c_450_n
+ PM_SKY130_FD_SC_MS__A32O_2%A_349_368#
x_PM_SKY130_FD_SC_MS__A32O_2%VGND N_VGND_M1003_d N_VGND_M1009_d N_VGND_M1008_d
+ N_VGND_c_491_n N_VGND_c_492_n N_VGND_c_493_n N_VGND_c_494_n N_VGND_c_495_n
+ N_VGND_c_496_n VGND N_VGND_c_497_n N_VGND_c_498_n N_VGND_c_499_n
+ PM_SKY130_FD_SC_MS__A32O_2%VGND
cc_1 VNB N_A_45_264#_M1004_g 5.17164e-19 $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A_45_264#_M1003_g 0.0282752f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_3 VNB N_A_45_264#_M1005_g 4.93277e-19 $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_4 VNB N_A_45_264#_M1009_g 0.0244304f $X=-0.19 $Y=-0.245 $X2=1 $Y2=0.74
cc_5 VNB N_A_45_264#_c_79_n 3.74074e-19 $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=2.32
cc_6 VNB N_A_45_264#_c_80_n 0.00921004f $X=-0.19 $Y=-0.245 $X2=1.19 $Y2=1.95
cc_7 VNB N_A_45_264#_c_81_n 0.0335619f $X=-0.19 $Y=-0.245 $X2=2.775 $Y2=1.095
cc_8 VNB N_A_45_264#_c_82_n 8.19761e-19 $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=1.095
cc_9 VNB N_A_45_264#_c_83_n 0.00342903f $X=-0.19 $Y=-0.245 $X2=2.94 $Y2=0.515
cc_10 VNB N_A_45_264#_c_84_n 0.00395055f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.485
cc_11 VNB N_A_45_264#_c_85_n 0.0753176f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.485
cc_12 VNB N_A3_M1007_g 0.0265047f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.65
cc_13 VNB N_A3_c_192_n 0.0286464f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_14 VNB N_A3_c_193_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_15 VNB N_A2_M1006_g 0.0254275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A2_c_228_n 0.0270247f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_17 VNB N_A2_c_229_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_18 VNB N_A1_M1011_g 0.0278022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_263_n 0.0250761f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_20 VNB N_A1_c_264_n 0.00414591f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_21 VNB N_B1_M1002_g 0.0285948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB B1 0.0133269f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_23 VNB N_B1_c_303_n 0.0274234f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_24 VNB N_B2_M1008_g 0.0298505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B2_M1013_g 0.00188935f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.65
cc_26 VNB N_B2_c_339_n 0.0594419f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.65
cc_27 VNB N_B2_c_340_n 0.00521402f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_28 VNB N_VPWR_c_361_n 0.183584f $X=-0.19 $Y=-0.245 $X2=2.94 $Y2=0.515
cc_29 VNB N_X_c_416_n 0.00240426f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_30 VNB N_X_c_417_n 0.00136575f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_31 VNB N_X_c_418_n 0.00120578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_491_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_492_n 0.0482617f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_34 VNB N_VGND_c_493_n 0.0209012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_494_n 0.0099193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_495_n 0.0128247f $X=-0.19 $Y=-0.245 $X2=1 $Y2=0.74
cc_37 VNB N_VGND_c_496_n 0.040801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_497_n 0.0715204f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=2.405
cc_39 VNB N_VGND_c_498_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_499_n 0.292107f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.485
cc_41 VPB N_A_45_264#_M1004_g 0.0245552f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_42 VPB N_A_45_264#_M1005_g 0.0240549f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_43 VPB N_A_45_264#_c_79_n 0.00759572f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=2.32
cc_44 VPB N_A_45_264#_c_80_n 0.00344843f $X=-0.19 $Y=1.66 $X2=1.19 $Y2=1.95
cc_45 VPB N_A3_M1010_g 0.0223182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A3_c_192_n 0.00575519f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_47 VPB N_A3_c_193_n 0.00277039f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_48 VPB N_A2_M1012_g 0.0229979f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.65
cc_49 VPB N_A2_c_228_n 0.0056732f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_50 VPB N_A2_c_229_n 0.00208071f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_51 VPB N_A1_M1000_g 0.0217685f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.65
cc_52 VPB N_A1_c_263_n 0.00554211f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_53 VPB N_A1_c_264_n 0.00344296f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_54 VPB N_B1_M1001_g 0.0202329f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.65
cc_55 VPB B1 0.00555587f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_56 VPB N_B1_c_303_n 0.00545172f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_57 VPB N_B2_M1013_g 0.0274233f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.65
cc_58 VPB N_B2_c_340_n 0.00764817f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_59 VPB N_VPWR_c_362_n 0.0119967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_363_n 0.0215351f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_61 VPB N_VPWR_c_364_n 0.0145679f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_62 VPB N_VPWR_c_365_n 0.0176541f $X=-0.19 $Y=1.66 $X2=1 $Y2=0.74
cc_63 VPB N_VPWR_c_366_n 0.0206218f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=2.32
cc_64 VPB N_VPWR_c_367_n 0.0219379f $X=-0.19 $Y=1.66 $X2=1.19 $Y2=2.12
cc_65 VPB N_VPWR_c_368_n 0.0429452f $X=-0.19 $Y=1.66 $X2=2.94 $Y2=0.515
cc_66 VPB N_VPWR_c_361_n 0.0801501f $X=-0.19 $Y=1.66 $X2=2.94 $Y2=0.515
cc_67 VPB N_VPWR_c_370_n 0.00786036f $X=-0.19 $Y=1.66 $X2=0.39 $Y2=1.485
cc_68 VPB N_VPWR_c_371_n 0.00728331f $X=-0.19 $Y=1.66 $X2=1.19 $Y2=2.035
cc_69 VPB X 0.00218805f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_X_c_418_n 8.17269e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_349_368#_c_447_n 0.019349f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_72 VPB N_A_349_368#_c_448_n 0.00350307f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_73 VPB N_A_349_368#_c_449_n 0.0365874f $X=-0.19 $Y=1.66 $X2=1 $Y2=0.74
cc_74 VPB N_A_349_368#_c_450_n 0.00281339f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.65
cc_75 N_A_45_264#_M1005_g N_A3_M1010_g 0.0211388f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_76 N_A_45_264#_c_91_p N_A3_M1010_g 0.00177334f $X=1.105 $Y=2.405 $X2=0 $Y2=0
cc_77 N_A_45_264#_c_80_n N_A3_M1010_g 0.00366577f $X=1.19 $Y=1.95 $X2=0 $Y2=0
cc_78 N_A_45_264#_c_93_p N_A3_M1010_g 0.00364533f $X=1.19 $Y=2.32 $X2=0 $Y2=0
cc_79 N_A_45_264#_c_94_p N_A3_M1010_g 0.0170881f $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_80 N_A_45_264#_M1009_g N_A3_M1007_g 0.016139f $X=1 $Y=0.74 $X2=0 $Y2=0
cc_81 N_A_45_264#_c_80_n N_A3_M1007_g 0.00314558f $X=1.19 $Y=1.95 $X2=0 $Y2=0
cc_82 N_A_45_264#_c_81_n N_A3_M1007_g 0.0157478f $X=2.775 $Y=1.095 $X2=0 $Y2=0
cc_83 N_A_45_264#_c_80_n N_A3_c_192_n 0.00248328f $X=1.19 $Y=1.95 $X2=0 $Y2=0
cc_84 N_A_45_264#_c_81_n N_A3_c_192_n 0.00125621f $X=2.775 $Y=1.095 $X2=0 $Y2=0
cc_85 N_A_45_264#_c_94_p N_A3_c_192_n 5.45341e-19 $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_86 N_A_45_264#_c_85_n N_A3_c_192_n 0.0085561f $X=0.955 $Y=1.485 $X2=0 $Y2=0
cc_87 N_A_45_264#_c_80_n N_A3_c_193_n 0.0327294f $X=1.19 $Y=1.95 $X2=0 $Y2=0
cc_88 N_A_45_264#_c_81_n N_A3_c_193_n 0.0247243f $X=2.775 $Y=1.095 $X2=0 $Y2=0
cc_89 N_A_45_264#_c_94_p N_A3_c_193_n 0.0219071f $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_90 N_A_45_264#_c_81_n N_A2_M1006_g 0.0154058f $X=2.775 $Y=1.095 $X2=0 $Y2=0
cc_91 N_A_45_264#_c_94_p N_A2_M1012_g 0.0127017f $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_92 N_A_45_264#_c_81_n N_A2_c_228_n 0.00125903f $X=2.775 $Y=1.095 $X2=0 $Y2=0
cc_93 N_A_45_264#_c_94_p N_A2_c_228_n 7.08634e-19 $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_94 N_A_45_264#_c_81_n N_A2_c_229_n 0.0247243f $X=2.775 $Y=1.095 $X2=0 $Y2=0
cc_95 N_A_45_264#_c_94_p N_A2_c_229_n 0.0229716f $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_96 N_A_45_264#_c_81_n N_A1_M1011_g 0.0161075f $X=2.775 $Y=1.095 $X2=0 $Y2=0
cc_97 N_A_45_264#_c_83_n N_A1_M1011_g 0.00449149f $X=2.94 $Y=0.515 $X2=0 $Y2=0
cc_98 N_A_45_264#_c_94_p N_A1_M1000_g 0.012729f $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_99 N_A_45_264#_c_81_n N_A1_c_263_n 0.0013639f $X=2.775 $Y=1.095 $X2=0 $Y2=0
cc_100 N_A_45_264#_c_94_p N_A1_c_263_n 6.49771e-19 $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_101 N_A_45_264#_c_81_n N_A1_c_264_n 0.030842f $X=2.775 $Y=1.095 $X2=0 $Y2=0
cc_102 N_A_45_264#_c_94_p N_A1_c_264_n 0.027438f $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_103 N_A_45_264#_c_81_n N_B1_M1002_g 0.00292704f $X=2.775 $Y=1.095 $X2=0 $Y2=0
cc_104 N_A_45_264#_c_83_n N_B1_M1002_g 0.0044057f $X=2.94 $Y=0.515 $X2=0 $Y2=0
cc_105 N_A_45_264#_c_94_p N_B1_M1001_g 0.0141869f $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_106 N_A_45_264#_c_94_p B1 0.0148329f $X=3.375 $Y=2.035 $X2=0 $Y2=0
cc_107 N_A_45_264#_c_122_p B1 0.0258499f $X=3.54 $Y=2.065 $X2=0 $Y2=0
cc_108 N_A_45_264#_c_122_p N_B1_c_303_n 5.85255e-19 $X=3.54 $Y=2.065 $X2=0 $Y2=0
cc_109 N_A_45_264#_c_79_n N_VPWR_M1004_s 0.0205644f $X=0.31 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_110 N_A_45_264#_c_125_p N_VPWR_M1004_s 0.00920379f $X=0.395 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_111 N_A_45_264#_c_91_p N_VPWR_M1005_s 0.00463428f $X=1.105 $Y=2.405 $X2=0
+ $Y2=0
cc_112 N_A_45_264#_c_80_n N_VPWR_M1005_s 0.0032334f $X=1.19 $Y=1.95 $X2=0 $Y2=0
cc_113 N_A_45_264#_c_93_p N_VPWR_M1005_s 0.00528913f $X=1.19 $Y=2.32 $X2=0 $Y2=0
cc_114 N_A_45_264#_c_94_p N_VPWR_M1005_s 0.0123997f $X=3.375 $Y=2.035 $X2=0
+ $Y2=0
cc_115 N_A_45_264#_c_130_p N_VPWR_M1005_s 0.00295606f $X=1.19 $Y=2.035 $X2=0
+ $Y2=0
cc_116 N_A_45_264#_c_94_p N_VPWR_M1012_d 0.0151027f $X=3.375 $Y=2.035 $X2=0
+ $Y2=0
cc_117 N_A_45_264#_M1004_g N_VPWR_c_363_n 0.012355f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A_45_264#_M1005_g N_VPWR_c_363_n 0.00130014f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_119 N_A_45_264#_c_91_p N_VPWR_c_363_n 0.0021187f $X=1.105 $Y=2.405 $X2=0
+ $Y2=0
cc_120 N_A_45_264#_c_125_p N_VPWR_c_363_n 0.0116597f $X=0.395 $Y=2.405 $X2=0
+ $Y2=0
cc_121 N_A_45_264#_M1005_g N_VPWR_c_364_n 0.00602407f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_122 N_A_45_264#_c_91_p N_VPWR_c_364_n 0.0148723f $X=1.105 $Y=2.405 $X2=0
+ $Y2=0
cc_123 N_A_45_264#_c_94_p N_VPWR_c_364_n 0.00799152f $X=3.375 $Y=2.035 $X2=0
+ $Y2=0
cc_124 N_A_45_264#_M1004_g N_VPWR_c_366_n 0.00460063f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_125 N_A_45_264#_M1005_g N_VPWR_c_366_n 0.00553757f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_126 N_A_45_264#_M1004_g N_VPWR_c_361_n 0.0046086f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_127 N_A_45_264#_M1005_g N_VPWR_c_361_n 0.00560227f $X=0.955 $Y=2.4 $X2=0
+ $Y2=0
cc_128 N_A_45_264#_c_91_p N_VPWR_c_361_n 0.0210935f $X=1.105 $Y=2.405 $X2=0
+ $Y2=0
cc_129 N_A_45_264#_c_125_p N_VPWR_c_361_n 6.15054e-19 $X=0.395 $Y=2.405 $X2=0
+ $Y2=0
cc_130 N_A_45_264#_c_91_p N_X_M1004_d 0.00472722f $X=1.105 $Y=2.405 $X2=0 $Y2=0
cc_131 N_A_45_264#_M1003_g N_X_c_416_n 0.00868565f $X=0.56 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A_45_264#_M1009_g N_X_c_416_n 0.0107619f $X=1 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A_45_264#_M1003_g N_X_c_417_n 0.00332192f $X=0.56 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A_45_264#_M1009_g N_X_c_417_n 0.00221233f $X=1 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A_45_264#_c_82_n N_X_c_417_n 0.00969158f $X=1.275 $Y=1.095 $X2=0 $Y2=0
cc_136 N_A_45_264#_M1004_g X 0.0058762f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A_45_264#_M1005_g X 0.00589497f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_138 N_A_45_264#_c_79_n X 0.0133159f $X=0.31 $Y=2.32 $X2=0 $Y2=0
cc_139 N_A_45_264#_c_91_p X 0.0196168f $X=1.105 $Y=2.405 $X2=0 $Y2=0
cc_140 N_A_45_264#_c_93_p X 0.00219866f $X=1.19 $Y=2.32 $X2=0 $Y2=0
cc_141 N_A_45_264#_c_130_p X 0.0141516f $X=1.19 $Y=2.035 $X2=0 $Y2=0
cc_142 N_A_45_264#_c_85_n X 0.0012997f $X=0.955 $Y=1.485 $X2=0 $Y2=0
cc_143 N_A_45_264#_M1004_g N_X_c_418_n 9.76882e-19 $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A_45_264#_M1003_g N_X_c_418_n 0.00286404f $X=0.56 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A_45_264#_M1005_g N_X_c_418_n 0.00379794f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_146 N_A_45_264#_M1009_g N_X_c_418_n 0.00323488f $X=1 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A_45_264#_c_79_n N_X_c_418_n 0.0057604f $X=0.31 $Y=2.32 $X2=0 $Y2=0
cc_148 N_A_45_264#_c_80_n N_X_c_418_n 0.0564947f $X=1.19 $Y=1.95 $X2=0 $Y2=0
cc_149 N_A_45_264#_c_84_n N_X_c_418_n 0.0239356f $X=0.39 $Y=1.485 $X2=0 $Y2=0
cc_150 N_A_45_264#_c_85_n N_X_c_418_n 0.0175067f $X=0.955 $Y=1.485 $X2=0 $Y2=0
cc_151 N_A_45_264#_c_94_p N_A_349_368#_M1010_d 0.00761058f $X=3.375 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_152 N_A_45_264#_c_94_p N_A_349_368#_M1000_d 0.00761058f $X=3.375 $Y=2.035
+ $X2=0 $Y2=0
cc_153 N_A_45_264#_c_94_p N_A_349_368#_c_453_n 0.0504818f $X=3.375 $Y=2.035
+ $X2=0 $Y2=0
cc_154 N_A_45_264#_c_94_p N_A_349_368#_c_454_n 0.0171782f $X=3.375 $Y=2.035
+ $X2=0 $Y2=0
cc_155 N_A_45_264#_c_122_p N_A_349_368#_c_447_n 0.0225479f $X=3.54 $Y=2.065
+ $X2=0 $Y2=0
cc_156 N_A_45_264#_M1005_g N_A_349_368#_c_450_n 7.84453e-19 $X=0.955 $Y=2.4
+ $X2=0 $Y2=0
cc_157 N_A_45_264#_c_91_p N_A_349_368#_c_450_n 0.00700984f $X=1.105 $Y=2.405
+ $X2=0 $Y2=0
cc_158 N_A_45_264#_c_93_p N_A_349_368#_c_450_n 0.00110642f $X=1.19 $Y=2.32 $X2=0
+ $Y2=0
cc_159 N_A_45_264#_c_94_p N_A_349_368#_c_450_n 0.0169008f $X=3.375 $Y=2.035
+ $X2=0 $Y2=0
cc_160 N_A_45_264#_c_81_n N_VGND_M1009_d 0.00551645f $X=2.775 $Y=1.095 $X2=0
+ $Y2=0
cc_161 N_A_45_264#_c_82_n N_VGND_M1009_d 0.00421237f $X=1.275 $Y=1.095 $X2=0
+ $Y2=0
cc_162 N_A_45_264#_M1003_g N_VGND_c_492_n 0.019585f $X=0.56 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A_45_264#_c_84_n N_VGND_c_492_n 0.0176651f $X=0.39 $Y=1.485 $X2=0 $Y2=0
cc_164 N_A_45_264#_c_85_n N_VGND_c_492_n 0.0016984f $X=0.955 $Y=1.485 $X2=0
+ $Y2=0
cc_165 N_A_45_264#_M1003_g N_VGND_c_493_n 0.00439591f $X=0.56 $Y=0.74 $X2=0
+ $Y2=0
cc_166 N_A_45_264#_M1009_g N_VGND_c_493_n 0.00451103f $X=1 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A_45_264#_M1009_g N_VGND_c_494_n 0.00798291f $X=1 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A_45_264#_c_81_n N_VGND_c_494_n 0.0194082f $X=2.775 $Y=1.095 $X2=0
+ $Y2=0
cc_169 N_A_45_264#_c_82_n N_VGND_c_494_n 0.0080244f $X=1.275 $Y=1.095 $X2=0
+ $Y2=0
cc_170 N_A_45_264#_c_83_n N_VGND_c_497_n 0.0146357f $X=2.94 $Y=0.515 $X2=0 $Y2=0
cc_171 N_A_45_264#_M1003_g N_VGND_c_499_n 0.00842009f $X=0.56 $Y=0.74 $X2=0
+ $Y2=0
cc_172 N_A_45_264#_M1009_g N_VGND_c_499_n 0.00878376f $X=1 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A_45_264#_c_83_n N_VGND_c_499_n 0.0121141f $X=2.94 $Y=0.515 $X2=0 $Y2=0
cc_174 N_A_45_264#_c_81_n A_355_74# 0.0048076f $X=2.775 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_175 N_A_45_264#_c_81_n A_433_74# 0.0120044f $X=2.775 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_176 N_A3_M1007_g N_A2_M1006_g 0.0395125f $X=1.7 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A3_M1010_g N_A2_M1012_g 0.0307472f $X=1.655 $Y=2.34 $X2=0 $Y2=0
cc_178 N_A3_c_193_n N_A2_M1012_g 5.9728e-19 $X=1.61 $Y=1.515 $X2=0 $Y2=0
cc_179 N_A3_c_192_n N_A2_c_228_n 0.0395125f $X=1.61 $Y=1.515 $X2=0 $Y2=0
cc_180 N_A3_c_193_n N_A2_c_228_n 0.00121489f $X=1.61 $Y=1.515 $X2=0 $Y2=0
cc_181 N_A3_c_192_n N_A2_c_229_n 0.00121489f $X=1.61 $Y=1.515 $X2=0 $Y2=0
cc_182 N_A3_c_193_n N_A2_c_229_n 0.0248916f $X=1.61 $Y=1.515 $X2=0 $Y2=0
cc_183 N_A3_M1010_g N_VPWR_c_364_n 0.00500933f $X=1.655 $Y=2.34 $X2=0 $Y2=0
cc_184 N_A3_M1010_g N_VPWR_c_367_n 0.00567889f $X=1.655 $Y=2.34 $X2=0 $Y2=0
cc_185 N_A3_M1010_g N_VPWR_c_361_n 0.00610055f $X=1.655 $Y=2.34 $X2=0 $Y2=0
cc_186 N_A3_M1007_g N_X_c_416_n 8.11115e-19 $X=1.7 $Y=0.74 $X2=0 $Y2=0
cc_187 N_A3_M1010_g N_A_349_368#_c_450_n 0.0108652f $X=1.655 $Y=2.34 $X2=0 $Y2=0
cc_188 N_A3_M1007_g N_VGND_c_494_n 0.0168903f $X=1.7 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A3_M1007_g N_VGND_c_497_n 0.00461464f $X=1.7 $Y=0.74 $X2=0 $Y2=0
cc_190 N_A3_M1007_g N_VGND_c_499_n 0.00911119f $X=1.7 $Y=0.74 $X2=0 $Y2=0
cc_191 N_A2_M1006_g N_A1_M1011_g 0.0343511f $X=2.09 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A2_M1012_g N_A1_M1000_g 0.0255177f $X=2.105 $Y=2.34 $X2=0 $Y2=0
cc_193 N_A2_c_229_n N_A1_M1000_g 2.64892e-19 $X=2.18 $Y=1.515 $X2=0 $Y2=0
cc_194 N_A2_c_228_n N_A1_c_263_n 0.0174173f $X=2.18 $Y=1.515 $X2=0 $Y2=0
cc_195 N_A2_c_229_n N_A1_c_263_n 3.73693e-19 $X=2.18 $Y=1.515 $X2=0 $Y2=0
cc_196 N_A2_M1012_g N_A1_c_264_n 3.02506e-19 $X=2.105 $Y=2.34 $X2=0 $Y2=0
cc_197 N_A2_c_228_n N_A1_c_264_n 0.00203135f $X=2.18 $Y=1.515 $X2=0 $Y2=0
cc_198 N_A2_c_229_n N_A1_c_264_n 0.0334556f $X=2.18 $Y=1.515 $X2=0 $Y2=0
cc_199 N_A2_M1012_g N_VPWR_c_365_n 0.00597119f $X=2.105 $Y=2.34 $X2=0 $Y2=0
cc_200 N_A2_M1012_g N_VPWR_c_367_n 0.00567889f $X=2.105 $Y=2.34 $X2=0 $Y2=0
cc_201 N_A2_M1012_g N_VPWR_c_361_n 0.00610055f $X=2.105 $Y=2.34 $X2=0 $Y2=0
cc_202 N_A2_M1012_g N_A_349_368#_c_453_n 0.0136887f $X=2.105 $Y=2.34 $X2=0 $Y2=0
cc_203 N_A2_M1012_g N_A_349_368#_c_462_n 7.71282e-19 $X=2.105 $Y=2.34 $X2=0
+ $Y2=0
cc_204 N_A2_M1012_g N_A_349_368#_c_450_n 0.00826575f $X=2.105 $Y=2.34 $X2=0
+ $Y2=0
cc_205 N_A2_M1006_g N_VGND_c_497_n 0.00461464f $X=2.09 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A2_M1006_g N_VGND_c_499_n 0.0091028f $X=2.09 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A1_M1011_g N_B1_M1002_g 0.0261158f $X=2.66 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A1_M1000_g N_B1_M1001_g 0.0309981f $X=2.815 $Y=2.34 $X2=0 $Y2=0
cc_209 N_A1_c_264_n N_B1_M1001_g 3.67631e-19 $X=2.75 $Y=1.515 $X2=0 $Y2=0
cc_210 N_A1_M1000_g B1 4.03377e-19 $X=2.815 $Y=2.34 $X2=0 $Y2=0
cc_211 N_A1_c_263_n B1 0.00121024f $X=2.75 $Y=1.515 $X2=0 $Y2=0
cc_212 N_A1_c_264_n B1 0.0266982f $X=2.75 $Y=1.515 $X2=0 $Y2=0
cc_213 N_A1_c_263_n N_B1_c_303_n 0.017626f $X=2.75 $Y=1.515 $X2=0 $Y2=0
cc_214 N_A1_c_264_n N_B1_c_303_n 4.19879e-19 $X=2.75 $Y=1.515 $X2=0 $Y2=0
cc_215 N_A1_M1000_g N_VPWR_c_365_n 0.00384059f $X=2.815 $Y=2.34 $X2=0 $Y2=0
cc_216 N_A1_M1000_g N_VPWR_c_368_n 0.00508554f $X=2.815 $Y=2.34 $X2=0 $Y2=0
cc_217 N_A1_M1000_g N_VPWR_c_361_n 0.00508379f $X=2.815 $Y=2.34 $X2=0 $Y2=0
cc_218 N_A1_M1000_g N_A_349_368#_c_453_n 0.0136887f $X=2.815 $Y=2.34 $X2=0 $Y2=0
cc_219 N_A1_M1000_g N_A_349_368#_c_454_n 8.84614e-19 $X=2.815 $Y=2.34 $X2=0
+ $Y2=0
cc_220 N_A1_M1000_g N_A_349_368#_c_462_n 0.00817391f $X=2.815 $Y=2.34 $X2=0
+ $Y2=0
cc_221 N_A1_M1000_g N_A_349_368#_c_448_n 0.00208236f $X=2.815 $Y=2.34 $X2=0
+ $Y2=0
cc_222 N_A1_M1000_g N_A_349_368#_c_450_n 7.60873e-19 $X=2.815 $Y=2.34 $X2=0
+ $Y2=0
cc_223 N_A1_M1011_g N_VGND_c_497_n 0.00461464f $X=2.66 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A1_M1011_g N_VGND_c_499_n 0.00911823f $X=2.66 $Y=0.74 $X2=0 $Y2=0
cc_225 N_B1_M1002_g N_B2_M1008_g 0.0306717f $X=3.23 $Y=0.74 $X2=0 $Y2=0
cc_226 N_B1_M1001_g N_B2_M1013_g 0.0151152f $X=3.265 $Y=2.34 $X2=0 $Y2=0
cc_227 B1 N_B2_c_339_n 0.00401057f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_228 N_B1_c_303_n N_B2_c_339_n 0.0174186f $X=3.32 $Y=1.515 $X2=0 $Y2=0
cc_229 N_B1_M1002_g N_B2_c_340_n 2.13129e-19 $X=3.23 $Y=0.74 $X2=0 $Y2=0
cc_230 B1 N_B2_c_340_n 0.0354768f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_231 N_B1_c_303_n N_B2_c_340_n 2.22391e-19 $X=3.32 $Y=1.515 $X2=0 $Y2=0
cc_232 N_B1_M1001_g N_VPWR_c_368_n 8.89343e-19 $X=3.265 $Y=2.34 $X2=0 $Y2=0
cc_233 N_B1_M1001_g N_A_349_368#_c_454_n 0.00235686f $X=3.265 $Y=2.34 $X2=0
+ $Y2=0
cc_234 N_B1_M1001_g N_A_349_368#_c_462_n 0.00741339f $X=3.265 $Y=2.34 $X2=0
+ $Y2=0
cc_235 N_B1_M1001_g N_A_349_368#_c_447_n 0.0108527f $X=3.265 $Y=2.34 $X2=0 $Y2=0
cc_236 N_B1_M1001_g N_A_349_368#_c_448_n 0.00141162f $X=3.265 $Y=2.34 $X2=0
+ $Y2=0
cc_237 N_B1_M1001_g N_A_349_368#_c_449_n 4.89222e-19 $X=3.265 $Y=2.34 $X2=0
+ $Y2=0
cc_238 N_B1_M1002_g N_VGND_c_496_n 0.00407036f $X=3.23 $Y=0.74 $X2=0 $Y2=0
cc_239 N_B1_M1002_g N_VGND_c_497_n 0.00461464f $X=3.23 $Y=0.74 $X2=0 $Y2=0
cc_240 N_B1_M1002_g N_VGND_c_499_n 0.00911823f $X=3.23 $Y=0.74 $X2=0 $Y2=0
cc_241 N_B2_M1013_g N_VPWR_c_368_n 8.89343e-19 $X=3.815 $Y=2.34 $X2=0 $Y2=0
cc_242 N_B2_M1013_g N_A_349_368#_c_462_n 4.17027e-19 $X=3.815 $Y=2.34 $X2=0
+ $Y2=0
cc_243 N_B2_M1013_g N_A_349_368#_c_447_n 0.0128353f $X=3.815 $Y=2.34 $X2=0 $Y2=0
cc_244 N_B2_M1013_g N_A_349_368#_c_449_n 0.0193497f $X=3.815 $Y=2.34 $X2=0 $Y2=0
cc_245 N_B2_c_339_n N_A_349_368#_c_449_n 0.00152096f $X=4.05 $Y=1.465 $X2=0
+ $Y2=0
cc_246 N_B2_c_340_n N_A_349_368#_c_449_n 0.0257606f $X=4.05 $Y=1.465 $X2=0 $Y2=0
cc_247 N_B2_M1008_g N_VGND_c_496_n 0.0240799f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_248 N_B2_c_339_n N_VGND_c_496_n 0.00284946f $X=4.05 $Y=1.465 $X2=0 $Y2=0
cc_249 N_B2_c_340_n N_VGND_c_496_n 0.0254821f $X=4.05 $Y=1.465 $X2=0 $Y2=0
cc_250 N_B2_M1008_g N_VGND_c_497_n 0.00383152f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_251 N_B2_M1008_g N_VGND_c_499_n 0.00758792f $X=3.8 $Y=0.74 $X2=0 $Y2=0
cc_252 N_VPWR_M1012_d N_A_349_368#_c_453_n 0.0113265f $X=2.195 $Y=1.84 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_365_n N_A_349_368#_c_453_n 0.0307535f $X=2.46 $Y=2.715 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_365_n N_A_349_368#_c_462_n 0.0171892f $X=2.46 $Y=2.715 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_368_n N_A_349_368#_c_447_n 0.0667586f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_256 N_VPWR_c_361_n N_A_349_368#_c_447_n 0.0380121f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_365_n N_A_349_368#_c_448_n 0.0119783f $X=2.46 $Y=2.715 $X2=0
+ $Y2=0
cc_258 N_VPWR_c_368_n N_A_349_368#_c_448_n 0.0236566f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_361_n N_A_349_368#_c_448_n 0.0128296f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_260 N_VPWR_c_364_n N_A_349_368#_c_450_n 0.00717656f $X=1.305 $Y=2.825 $X2=0
+ $Y2=0
cc_261 N_VPWR_c_365_n N_A_349_368#_c_450_n 0.0148393f $X=2.46 $Y=2.715 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_367_n N_A_349_368#_c_450_n 0.00955252f $X=2.265 $Y=3.33 $X2=0
+ $Y2=0
cc_263 N_VPWR_c_361_n N_A_349_368#_c_450_n 0.0110607f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_264 N_X_c_416_n N_VGND_c_492_n 0.0322525f $X=0.78 $Y=0.495 $X2=0 $Y2=0
cc_265 N_X_c_416_n N_VGND_c_493_n 0.0153382f $X=0.78 $Y=0.495 $X2=0 $Y2=0
cc_266 N_X_c_416_n N_VGND_c_494_n 0.0294488f $X=0.78 $Y=0.495 $X2=0 $Y2=0
cc_267 N_X_c_416_n N_VGND_c_499_n 0.0117503f $X=0.78 $Y=0.495 $X2=0 $Y2=0

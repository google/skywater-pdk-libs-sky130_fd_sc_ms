* File: sky130_fd_sc_ms__clkinv_16.pex.spice
* Created: Fri Aug 28 17:19:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__CLKINV_16%A 3 7 11 15 19 23 27 31 35 39 43 47 51 55
+ 59 63 67 71 75 79 83 87 91 95 99 103 107 111 115 119 123 127 131 135 139 143
+ 147 151 155 159 161 227 231 237 243 249 255 261 267 273 277
c413 227 0 1.45923e-19 $X=10.75 $Y=1.485
c414 95 0 1.88851e-19 $X=5.645 $Y=0.61
c415 55 0 1.6166e-19 $X=3.215 $Y=0.61
r416 274 277 1.84782 $w=2.3e-07 $l=2.88e-06 $layer=MET1_cond $X=7.83 $Y=1.295
+ $X2=10.71 $Y2=1.295
r417 273 277 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=10.71
+ $Y=1.295 $X2=10.71 $Y2=1.295
r418 273 274 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.83
+ $Y=1.295 $X2=7.83 $Y2=1.295
r419 268 274 0.718597 $w=2.3e-07 $l=1.12e-06 $layer=MET1_cond $X=6.71 $Y=1.295
+ $X2=7.83 $Y2=1.295
r420 267 268 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.71 $Y=1.295
+ $X2=6.71 $Y2=1.295
r421 261 262 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.76 $Y=1.295
+ $X2=5.76 $Y2=1.295
r422 256 262 0.538948 $w=2.3e-07 $l=8.4e-07 $layer=MET1_cond $X=4.92 $Y=1.295
+ $X2=5.76 $Y2=1.295
r423 255 256 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.92 $Y=1.295
+ $X2=4.92 $Y2=1.295
r424 250 256 0.635188 $w=2.3e-07 $l=9.9e-07 $layer=MET1_cond $X=3.93 $Y=1.295
+ $X2=4.92 $Y2=1.295
r425 249 250 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.93 $Y=1.295
+ $X2=3.93 $Y2=1.295
r426 244 250 0.596692 $w=2.3e-07 $l=9.3e-07 $layer=MET1_cond $X=3 $Y=1.295
+ $X2=3.93 $Y2=1.295
r427 243 244 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3 $Y=1.295 $X2=3
+ $Y2=1.295
r428 238 244 0.622356 $w=2.3e-07 $l=9.7e-07 $layer=MET1_cond $X=2.03 $Y=1.295
+ $X2=3 $Y2=1.295
r429 237 238 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.03 $Y=1.295
+ $X2=2.03 $Y2=1.295
r430 232 238 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=1.13 $Y=1.295
+ $X2=2.03 $Y2=1.295
r431 231 232 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.13 $Y=1.295
+ $X2=1.13 $Y2=1.295
r432 227 229 35.5794 $w=3.59e-07 $l=2.65e-07 $layer=POLY_cond $X=10.75 $Y=1.5
+ $X2=11.015 $Y2=1.5
r433 225 227 24.8384 $w=3.59e-07 $l=1.85e-07 $layer=POLY_cond $X=10.565 $Y=1.5
+ $X2=10.75 $Y2=1.5
r434 224 225 60.4178 $w=3.59e-07 $l=4.5e-07 $layer=POLY_cond $X=10.115 $Y=1.5
+ $X2=10.565 $Y2=1.5
r435 223 224 60.4178 $w=3.59e-07 $l=4.5e-07 $layer=POLY_cond $X=9.665 $Y=1.5
+ $X2=10.115 $Y2=1.5
r436 222 223 60.4178 $w=3.59e-07 $l=4.5e-07 $layer=POLY_cond $X=9.215 $Y=1.5
+ $X2=9.665 $Y2=1.5
r437 221 222 60.4178 $w=3.59e-07 $l=4.5e-07 $layer=POLY_cond $X=8.765 $Y=1.5
+ $X2=9.215 $Y2=1.5
r438 220 221 60.4178 $w=3.59e-07 $l=4.5e-07 $layer=POLY_cond $X=8.315 $Y=1.5
+ $X2=8.765 $Y2=1.5
r439 219 220 60.4178 $w=3.59e-07 $l=4.5e-07 $layer=POLY_cond $X=7.865 $Y=1.5
+ $X2=8.315 $Y2=1.5
r440 218 273 0.683776 $w=3.388e-06 $l=1.9e-07 $layer=LI1_cond $X=9.22 $Y=1.485
+ $X2=9.22 $Y2=1.295
r441 218 227 29.056 $w=1.7e-07 $l=8.5e-07 $layer=licon1_POLY $count=5 $X=10.75
+ $Y=1.485 $X2=10.75 $Y2=1.485
r442 217 219 23.4958 $w=3.59e-07 $l=1.75e-07 $layer=POLY_cond $X=7.69 $Y=1.5
+ $X2=7.865 $Y2=1.5
r443 217 218 29.056 $w=1.7e-07 $l=8.5e-07 $layer=licon1_POLY $count=5 $X=7.69
+ $Y=1.485 $X2=7.69 $Y2=1.485
r444 215 217 36.922 $w=3.59e-07 $l=2.75e-07 $layer=POLY_cond $X=7.415 $Y=1.5
+ $X2=7.69 $Y2=1.5
r445 214 215 6.71309 $w=3.59e-07 $l=5e-08 $layer=POLY_cond $X=7.365 $Y=1.5
+ $X2=7.415 $Y2=1.5
r446 213 214 57.7326 $w=3.59e-07 $l=4.3e-07 $layer=POLY_cond $X=6.935 $Y=1.5
+ $X2=7.365 $Y2=1.5
r447 212 213 4.02785 $w=3.59e-07 $l=3e-08 $layer=POLY_cond $X=6.905 $Y=1.5
+ $X2=6.935 $Y2=1.5
r448 211 267 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=6.71 $Y=1.485
+ $X2=6.71 $Y2=1.295
r449 210 212 26.1811 $w=3.59e-07 $l=1.95e-07 $layer=POLY_cond $X=6.71 $Y=1.5
+ $X2=6.905 $Y2=1.5
r450 210 211 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.71
+ $Y=1.485 $X2=6.71 $Y2=1.485
r451 208 210 27.5237 $w=3.59e-07 $l=2.05e-07 $layer=POLY_cond $X=6.505 $Y=1.5
+ $X2=6.71 $Y2=1.5
r452 207 208 13.4262 $w=3.59e-07 $l=1e-07 $layer=POLY_cond $X=6.405 $Y=1.5
+ $X2=6.505 $Y2=1.5
r453 206 207 44.3064 $w=3.59e-07 $l=3.3e-07 $layer=POLY_cond $X=6.075 $Y=1.5
+ $X2=6.405 $Y2=1.5
r454 205 206 16.1114 $w=3.59e-07 $l=1.2e-07 $layer=POLY_cond $X=5.955 $Y=1.5
+ $X2=6.075 $Y2=1.5
r455 204 261 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=5.76 $Y=1.485
+ $X2=5.76 $Y2=1.295
r456 203 205 26.1811 $w=3.59e-07 $l=1.95e-07 $layer=POLY_cond $X=5.76 $Y=1.5
+ $X2=5.955 $Y2=1.5
r457 203 204 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.76
+ $Y=1.485 $X2=5.76 $Y2=1.485
r458 201 203 15.4401 $w=3.59e-07 $l=1.15e-07 $layer=POLY_cond $X=5.645 $Y=1.5
+ $X2=5.76 $Y2=1.5
r459 200 201 25.5097 $w=3.59e-07 $l=1.9e-07 $layer=POLY_cond $X=5.455 $Y=1.5
+ $X2=5.645 $Y2=1.5
r460 199 200 32.2228 $w=3.59e-07 $l=2.4e-07 $layer=POLY_cond $X=5.215 $Y=1.5
+ $X2=5.455 $Y2=1.5
r461 198 199 28.195 $w=3.59e-07 $l=2.1e-07 $layer=POLY_cond $X=5.005 $Y=1.5
+ $X2=5.215 $Y2=1.5
r462 197 255 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.92 $Y=1.485
+ $X2=4.92 $Y2=1.295
r463 196 198 11.4123 $w=3.59e-07 $l=8.5e-08 $layer=POLY_cond $X=4.92 $Y=1.5
+ $X2=5.005 $Y2=1.5
r464 196 197 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.92
+ $Y=1.485 $X2=4.92 $Y2=1.485
r465 194 196 36.922 $w=3.59e-07 $l=2.75e-07 $layer=POLY_cond $X=4.645 $Y=1.5
+ $X2=4.92 $Y2=1.5
r466 193 194 12.0836 $w=3.59e-07 $l=9e-08 $layer=POLY_cond $X=4.555 $Y=1.5
+ $X2=4.645 $Y2=1.5
r467 192 193 45.649 $w=3.59e-07 $l=3.4e-07 $layer=POLY_cond $X=4.215 $Y=1.5
+ $X2=4.555 $Y2=1.5
r468 191 192 14.7688 $w=3.59e-07 $l=1.1e-07 $layer=POLY_cond $X=4.105 $Y=1.5
+ $X2=4.215 $Y2=1.5
r469 190 249 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.93 $Y=1.485
+ $X2=3.93 $Y2=1.295
r470 189 191 23.4958 $w=3.59e-07 $l=1.75e-07 $layer=POLY_cond $X=3.93 $Y=1.5
+ $X2=4.105 $Y2=1.5
r471 189 190 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.93
+ $Y=1.485 $X2=3.93 $Y2=1.485
r472 187 189 36.922 $w=3.59e-07 $l=2.75e-07 $layer=POLY_cond $X=3.655 $Y=1.5
+ $X2=3.93 $Y2=1.5
r473 186 187 1.34262 $w=3.59e-07 $l=1e-08 $layer=POLY_cond $X=3.645 $Y=1.5
+ $X2=3.655 $Y2=1.5
r474 185 186 57.7326 $w=3.59e-07 $l=4.3e-07 $layer=POLY_cond $X=3.215 $Y=1.5
+ $X2=3.645 $Y2=1.5
r475 184 185 1.34262 $w=3.59e-07 $l=1e-08 $layer=POLY_cond $X=3.205 $Y=1.5
+ $X2=3.215 $Y2=1.5
r476 183 243 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3 $Y=1.485 $X2=3
+ $Y2=1.295
r477 182 184 27.5237 $w=3.59e-07 $l=2.05e-07 $layer=POLY_cond $X=3 $Y=1.5
+ $X2=3.205 $Y2=1.5
r478 182 183 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3
+ $Y=1.485 $X2=3 $Y2=1.485
r479 180 182 32.8941 $w=3.59e-07 $l=2.45e-07 $layer=POLY_cond $X=2.755 $Y=1.5
+ $X2=3 $Y2=1.5
r480 179 180 5.37047 $w=3.59e-07 $l=4e-08 $layer=POLY_cond $X=2.715 $Y=1.5
+ $X2=2.755 $Y2=1.5
r481 178 179 55.0474 $w=3.59e-07 $l=4.1e-07 $layer=POLY_cond $X=2.305 $Y=1.5
+ $X2=2.715 $Y2=1.5
r482 177 178 2.68524 $w=3.59e-07 $l=2e-08 $layer=POLY_cond $X=2.285 $Y=1.5
+ $X2=2.305 $Y2=1.5
r483 176 237 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.03 $Y=1.485
+ $X2=2.03 $Y2=1.295
r484 175 177 34.2368 $w=3.59e-07 $l=2.55e-07 $layer=POLY_cond $X=2.03 $Y=1.5
+ $X2=2.285 $Y2=1.5
r485 175 176 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.03
+ $Y=1.485 $X2=2.03 $Y2=1.485
r486 173 175 23.4958 $w=3.59e-07 $l=1.75e-07 $layer=POLY_cond $X=1.855 $Y=1.5
+ $X2=2.03 $Y2=1.5
r487 172 173 9.39833 $w=3.59e-07 $l=7e-08 $layer=POLY_cond $X=1.785 $Y=1.5
+ $X2=1.855 $Y2=1.5
r488 171 172 51.0195 $w=3.59e-07 $l=3.8e-07 $layer=POLY_cond $X=1.405 $Y=1.5
+ $X2=1.785 $Y2=1.5
r489 170 171 6.71309 $w=3.59e-07 $l=5e-08 $layer=POLY_cond $X=1.355 $Y=1.5
+ $X2=1.405 $Y2=1.5
r490 169 231 6.84263 $w=3.18e-07 $l=1.9e-07 $layer=LI1_cond $X=1.135 $Y=1.485
+ $X2=1.135 $Y2=1.295
r491 168 170 30.2089 $w=3.59e-07 $l=2.25e-07 $layer=POLY_cond $X=1.13 $Y=1.5
+ $X2=1.355 $Y2=1.5
r492 168 169 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.485 $X2=1.13 $Y2=1.485
r493 166 168 23.4958 $w=3.59e-07 $l=1.75e-07 $layer=POLY_cond $X=0.955 $Y=1.5
+ $X2=1.13 $Y2=1.5
r494 165 166 4.02785 $w=3.59e-07 $l=3e-08 $layer=POLY_cond $X=0.925 $Y=1.5
+ $X2=0.955 $Y2=1.5
r495 164 165 56.39 $w=3.59e-07 $l=4.2e-07 $layer=POLY_cond $X=0.505 $Y=1.5
+ $X2=0.925 $Y2=1.5
r496 163 164 1.34262 $w=3.59e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.5
+ $X2=0.505 $Y2=1.5
r497 161 268 0.481203 $w=2.3e-07 $l=7.5e-07 $layer=MET1_cond $X=5.96 $Y=1.295
+ $X2=6.71 $Y2=1.295
r498 161 262 0.128321 $w=2.3e-07 $l=2e-07 $layer=MET1_cond $X=5.96 $Y=1.295
+ $X2=5.76 $Y2=1.295
r499 157 229 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=11.015 $Y=1.68
+ $X2=11.015 $Y2=1.5
r500 157 159 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=11.015 $Y=1.68
+ $X2=11.015 $Y2=2.4
r501 153 225 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=10.565 $Y=1.68
+ $X2=10.565 $Y2=1.5
r502 153 155 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=10.565 $Y=1.68
+ $X2=10.565 $Y2=2.4
r503 149 224 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=10.115 $Y=1.68
+ $X2=10.115 $Y2=1.5
r504 149 151 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=10.115 $Y=1.68
+ $X2=10.115 $Y2=2.4
r505 145 223 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=9.665 $Y=1.68
+ $X2=9.665 $Y2=1.5
r506 145 147 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=9.665 $Y=1.68
+ $X2=9.665 $Y2=2.4
r507 141 222 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=9.215 $Y=1.68
+ $X2=9.215 $Y2=1.5
r508 141 143 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=9.215 $Y=1.68
+ $X2=9.215 $Y2=2.4
r509 137 221 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=8.765 $Y=1.68
+ $X2=8.765 $Y2=1.5
r510 137 139 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.765 $Y=1.68
+ $X2=8.765 $Y2=2.4
r511 133 220 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=8.315 $Y=1.68
+ $X2=8.315 $Y2=1.5
r512 133 135 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.315 $Y=1.68
+ $X2=8.315 $Y2=2.4
r513 129 219 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=7.865 $Y=1.68
+ $X2=7.865 $Y2=1.5
r514 129 131 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.865 $Y=1.68
+ $X2=7.865 $Y2=2.4
r515 125 215 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=7.415 $Y=1.68
+ $X2=7.415 $Y2=1.5
r516 125 127 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.415 $Y=1.68
+ $X2=7.415 $Y2=2.4
r517 121 214 23.2387 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.365 $Y=1.32
+ $X2=7.365 $Y2=1.5
r518 121 123 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=7.365 $Y=1.32
+ $X2=7.365 $Y2=0.61
r519 117 213 23.2387 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.935 $Y=1.32
+ $X2=6.935 $Y2=1.5
r520 117 119 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.935 $Y=1.32
+ $X2=6.935 $Y2=0.61
r521 113 212 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=6.905 $Y=1.68
+ $X2=6.905 $Y2=1.5
r522 113 115 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.905 $Y=1.68
+ $X2=6.905 $Y2=2.4
r523 109 208 23.2387 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.505 $Y=1.32
+ $X2=6.505 $Y2=1.5
r524 109 111 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.505 $Y=1.32
+ $X2=6.505 $Y2=0.61
r525 105 207 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=6.405 $Y=1.68
+ $X2=6.405 $Y2=1.5
r526 105 107 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.405 $Y=1.68
+ $X2=6.405 $Y2=2.4
r527 101 206 23.2387 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.075 $Y=1.32
+ $X2=6.075 $Y2=1.5
r528 101 103 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.075 $Y=1.32
+ $X2=6.075 $Y2=0.61
r529 97 205 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=5.955 $Y=1.68
+ $X2=5.955 $Y2=1.5
r530 97 99 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.955 $Y=1.68
+ $X2=5.955 $Y2=2.4
r531 93 201 23.2387 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=5.645 $Y=1.32
+ $X2=5.645 $Y2=1.5
r532 93 95 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.645 $Y=1.32
+ $X2=5.645 $Y2=0.61
r533 89 200 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=5.455 $Y=1.68
+ $X2=5.455 $Y2=1.5
r534 89 91 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.455 $Y=1.68
+ $X2=5.455 $Y2=2.4
r535 85 199 23.2387 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=5.215 $Y=1.32
+ $X2=5.215 $Y2=1.5
r536 85 87 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.215 $Y=1.32
+ $X2=5.215 $Y2=0.61
r537 81 198 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=5.005 $Y=1.68
+ $X2=5.005 $Y2=1.5
r538 81 83 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.005 $Y=1.68
+ $X2=5.005 $Y2=2.4
r539 77 194 23.2387 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=4.645 $Y=1.32
+ $X2=4.645 $Y2=1.5
r540 77 79 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.645 $Y=1.32
+ $X2=4.645 $Y2=0.61
r541 73 193 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=4.555 $Y=1.68
+ $X2=4.555 $Y2=1.5
r542 73 75 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.555 $Y=1.68
+ $X2=4.555 $Y2=2.4
r543 69 192 23.2387 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=4.215 $Y=1.32
+ $X2=4.215 $Y2=1.5
r544 69 71 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.215 $Y=1.32
+ $X2=4.215 $Y2=0.61
r545 65 191 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=4.105 $Y=1.68
+ $X2=4.105 $Y2=1.5
r546 65 67 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.105 $Y=1.68
+ $X2=4.105 $Y2=2.4
r547 61 186 23.2387 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.645 $Y=1.32
+ $X2=3.645 $Y2=1.5
r548 61 63 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.645 $Y=1.32
+ $X2=3.645 $Y2=0.61
r549 57 187 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=3.655 $Y=1.68
+ $X2=3.655 $Y2=1.5
r550 57 59 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.655 $Y=1.68
+ $X2=3.655 $Y2=2.4
r551 53 185 23.2387 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.215 $Y=1.32
+ $X2=3.215 $Y2=1.5
r552 53 55 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.215 $Y=1.32
+ $X2=3.215 $Y2=0.61
r553 49 184 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=3.205 $Y=1.68
+ $X2=3.205 $Y2=1.5
r554 49 51 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.205 $Y=1.68
+ $X2=3.205 $Y2=2.4
r555 45 180 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=2.755 $Y=1.68
+ $X2=2.755 $Y2=1.5
r556 45 47 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.755 $Y=1.68
+ $X2=2.755 $Y2=2.4
r557 41 179 23.2387 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.715 $Y=1.32
+ $X2=2.715 $Y2=1.5
r558 41 43 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.715 $Y=1.32
+ $X2=2.715 $Y2=0.61
r559 37 178 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=2.305 $Y=1.68
+ $X2=2.305 $Y2=1.5
r560 37 39 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.305 $Y=1.68
+ $X2=2.305 $Y2=2.4
r561 33 177 23.2387 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.285 $Y=1.32
+ $X2=2.285 $Y2=1.5
r562 33 35 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.285 $Y=1.32
+ $X2=2.285 $Y2=0.61
r563 29 173 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=1.855 $Y=1.68
+ $X2=1.855 $Y2=1.5
r564 29 31 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.855 $Y=1.68
+ $X2=1.855 $Y2=2.4
r565 25 172 23.2387 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.785 $Y=1.32
+ $X2=1.785 $Y2=1.5
r566 25 27 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.785 $Y=1.32
+ $X2=1.785 $Y2=0.61
r567 21 171 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=1.405 $Y=1.68
+ $X2=1.405 $Y2=1.5
r568 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.405 $Y=1.68
+ $X2=1.405 $Y2=2.4
r569 17 170 23.2387 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.355 $Y=1.32
+ $X2=1.355 $Y2=1.5
r570 17 19 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.355 $Y=1.32
+ $X2=1.355 $Y2=0.61
r571 13 166 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=0.955 $Y=1.68
+ $X2=0.955 $Y2=1.5
r572 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.955 $Y=1.68
+ $X2=0.955 $Y2=2.4
r573 9 165 23.2387 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.925 $Y=1.32
+ $X2=0.925 $Y2=1.5
r574 9 11 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.925 $Y=1.32
+ $X2=0.925 $Y2=0.61
r575 5 163 23.2387 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.495 $Y=1.32
+ $X2=0.495 $Y2=1.5
r576 5 7 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.495 $Y=1.32
+ $X2=0.495 $Y2=0.61
r577 1 164 18.9031 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=0.505 $Y=1.68
+ $X2=0.505 $Y2=1.5
r578 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.505 $Y=1.68
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__CLKINV_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 40 42
+ 48 54 60 66 72 78 84 90 94 98 104 110 114 116 121 122 124 125 127 128 130 131
+ 133 134 136 137 139 140 141 142 143 170 175 180 189 192 195 199
r232 198 199 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r233 195 196 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r234 192 193 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r235 189 190 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r236 186 187 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r237 184 199 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r238 184 196 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=10.32 $Y2=3.33
r239 183 184 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r240 181 195 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.505 $Y=3.33
+ $X2=10.34 $Y2=3.33
r241 181 183 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.505 $Y=3.33
+ $X2=10.8 $Y2=3.33
r242 180 198 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=11.075 $Y=3.33
+ $X2=11.297 $Y2=3.33
r243 180 183 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.075 $Y=3.33
+ $X2=10.8 $Y2=3.33
r244 179 196 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r245 179 193 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r246 178 179 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r247 176 192 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.605 $Y=3.33
+ $X2=9.44 $Y2=3.33
r248 176 178 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.605 $Y=3.33
+ $X2=9.84 $Y2=3.33
r249 175 195 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.175 $Y=3.33
+ $X2=10.34 $Y2=3.33
r250 175 178 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=10.175 $Y=3.33
+ $X2=9.84 $Y2=3.33
r251 174 193 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r252 174 190 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r253 173 174 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r254 171 189 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.625 $Y=3.33
+ $X2=8.5 $Y2=3.33
r255 171 173 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.625 $Y=3.33
+ $X2=8.88 $Y2=3.33
r256 170 192 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.275 $Y=3.33
+ $X2=9.44 $Y2=3.33
r257 170 173 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=9.275 $Y=3.33
+ $X2=8.88 $Y2=3.33
r258 169 190 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r259 168 169 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r260 166 169 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r261 165 166 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r262 162 163 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r263 160 163 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r264 159 160 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r265 157 160 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r266 156 157 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r267 154 157 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r268 153 154 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r269 151 154 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r270 150 151 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r271 148 151 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r272 148 187 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r273 147 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r274 145 186 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r275 145 147 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r276 143 166 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=6.48 $Y2=3.33
r277 143 163 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=5.52 $Y2=3.33
r278 141 168 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=7.475 $Y=3.33
+ $X2=7.44 $Y2=3.33
r279 141 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.475 $Y=3.33
+ $X2=7.64 $Y2=3.33
r280 139 165 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=6.51 $Y=3.33
+ $X2=6.48 $Y2=3.33
r281 139 140 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=6.51 $Y=3.33
+ $X2=6.652 $Y2=3.33
r282 138 168 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=6.795 $Y=3.33
+ $X2=7.44 $Y2=3.33
r283 138 140 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=6.795 $Y=3.33
+ $X2=6.652 $Y2=3.33
r284 136 162 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=5.595 $Y=3.33
+ $X2=5.52 $Y2=3.33
r285 136 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.595 $Y=3.33
+ $X2=5.72 $Y2=3.33
r286 135 165 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=6.48 $Y2=3.33
r287 135 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=5.72 $Y2=3.33
r288 133 159 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.695 $Y=3.33
+ $X2=4.56 $Y2=3.33
r289 133 134 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.695 $Y=3.33
+ $X2=4.78 $Y2=3.33
r290 132 162 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.865 $Y=3.33
+ $X2=5.52 $Y2=3.33
r291 132 134 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.865 $Y=3.33
+ $X2=4.78 $Y2=3.33
r292 130 156 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.795 $Y=3.33
+ $X2=3.6 $Y2=3.33
r293 130 131 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.795 $Y=3.33
+ $X2=3.88 $Y2=3.33
r294 129 159 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.965 $Y=3.33
+ $X2=4.56 $Y2=3.33
r295 129 131 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.965 $Y=3.33
+ $X2=3.88 $Y2=3.33
r296 127 153 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=2.64 $Y2=3.33
r297 127 128 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=2.98 $Y2=3.33
r298 126 156 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.065 $Y=3.33
+ $X2=3.6 $Y2=3.33
r299 126 128 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=3.33
+ $X2=2.98 $Y2=3.33
r300 124 150 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=1.68 $Y2=3.33
r301 124 125 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=2.08 $Y2=3.33
r302 123 153 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.165 $Y=3.33
+ $X2=2.64 $Y2=3.33
r303 123 125 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=3.33
+ $X2=2.08 $Y2=3.33
r304 121 147 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r305 121 122 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.14 $Y2=3.33
r306 120 150 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.68 $Y2=3.33
r307 120 122 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.14 $Y2=3.33
r308 116 119 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=11.24 $Y=1.985
+ $X2=11.24 $Y2=2.815
r309 114 198 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=11.24 $Y=3.245
+ $X2=11.297 $Y2=3.33
r310 114 119 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.24 $Y=3.245
+ $X2=11.24 $Y2=2.815
r311 110 113 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=10.34 $Y=1.985
+ $X2=10.34 $Y2=2.815
r312 108 195 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.34 $Y=3.245
+ $X2=10.34 $Y2=3.33
r313 108 113 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.34 $Y=3.245
+ $X2=10.34 $Y2=2.815
r314 104 107 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=9.44 $Y=1.985
+ $X2=9.44 $Y2=2.815
r315 102 192 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.44 $Y=3.245
+ $X2=9.44 $Y2=3.33
r316 102 107 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=9.44 $Y=3.245
+ $X2=9.44 $Y2=2.815
r317 98 101 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=8.5 $Y=1.985
+ $X2=8.5 $Y2=2.815
r318 96 189 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.5 $Y=3.245
+ $X2=8.5 $Y2=3.33
r319 96 101 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.5 $Y=3.245
+ $X2=8.5 $Y2=2.815
r320 95 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.805 $Y=3.33
+ $X2=7.64 $Y2=3.33
r321 94 189 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.375 $Y=3.33
+ $X2=8.5 $Y2=3.33
r322 94 95 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.375 $Y=3.33
+ $X2=7.805 $Y2=3.33
r323 90 93 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=7.64 $Y=1.985
+ $X2=7.64 $Y2=2.815
r324 88 142 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.64 $Y=3.245
+ $X2=7.64 $Y2=3.33
r325 88 93 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.64 $Y=3.245
+ $X2=7.64 $Y2=2.815
r326 84 87 33.5624 $w=2.83e-07 $l=8.3e-07 $layer=LI1_cond $X=6.652 $Y=1.985
+ $X2=6.652 $Y2=2.815
r327 82 140 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=6.652 $Y=3.245
+ $X2=6.652 $Y2=3.33
r328 82 87 17.3877 $w=2.83e-07 $l=4.3e-07 $layer=LI1_cond $X=6.652 $Y=3.245
+ $X2=6.652 $Y2=2.815
r329 78 81 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=5.72 $Y=1.985
+ $X2=5.72 $Y2=2.815
r330 76 137 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.72 $Y=3.245
+ $X2=5.72 $Y2=3.33
r331 76 81 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.72 $Y=3.245
+ $X2=5.72 $Y2=2.815
r332 72 75 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.78 $Y=1.985
+ $X2=4.78 $Y2=2.815
r333 70 134 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.78 $Y=3.245
+ $X2=4.78 $Y2=3.33
r334 70 75 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.78 $Y=3.245
+ $X2=4.78 $Y2=2.815
r335 66 69 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.88 $Y=1.985
+ $X2=3.88 $Y2=2.815
r336 64 131 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.88 $Y=3.245
+ $X2=3.88 $Y2=3.33
r337 64 69 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.88 $Y=3.245
+ $X2=3.88 $Y2=2.815
r338 60 63 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.98 $Y=1.985
+ $X2=2.98 $Y2=2.815
r339 58 128 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=3.245
+ $X2=2.98 $Y2=3.33
r340 58 63 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.98 $Y=3.245
+ $X2=2.98 $Y2=2.815
r341 54 57 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.08 $Y=1.985
+ $X2=2.08 $Y2=2.815
r342 52 125 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=3.245
+ $X2=2.08 $Y2=3.33
r343 52 57 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.08 $Y=3.245
+ $X2=2.08 $Y2=2.815
r344 48 51 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=1.14 $Y=1.985
+ $X2=1.14 $Y2=2.815
r345 46 122 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=3.33
r346 46 51 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=2.815
r347 42 45 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r348 40 186 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r349 40 45 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r350 13 119 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=11.105
+ $Y=1.84 $X2=11.24 $Y2=2.815
r351 13 116 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=11.105
+ $Y=1.84 $X2=11.24 $Y2=1.985
r352 12 113 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.205
+ $Y=1.84 $X2=10.34 $Y2=2.815
r353 12 110 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.205
+ $Y=1.84 $X2=10.34 $Y2=1.985
r354 11 107 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.305
+ $Y=1.84 $X2=9.44 $Y2=2.815
r355 11 104 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.305
+ $Y=1.84 $X2=9.44 $Y2=1.985
r356 10 101 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.405
+ $Y=1.84 $X2=8.54 $Y2=2.815
r357 10 98 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.405
+ $Y=1.84 $X2=8.54 $Y2=1.985
r358 9 93 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.505
+ $Y=1.84 $X2=7.64 $Y2=2.815
r359 9 90 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.505
+ $Y=1.84 $X2=7.64 $Y2=1.985
r360 8 87 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.495
+ $Y=1.84 $X2=6.63 $Y2=2.815
r361 8 84 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.495
+ $Y=1.84 $X2=6.63 $Y2=1.985
r362 7 81 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.545
+ $Y=1.84 $X2=5.68 $Y2=2.815
r363 7 78 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.545
+ $Y=1.84 $X2=5.68 $Y2=1.985
r364 6 75 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.645
+ $Y=1.84 $X2=4.78 $Y2=2.815
r365 6 72 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.645
+ $Y=1.84 $X2=4.78 $Y2=1.985
r366 5 69 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.745
+ $Y=1.84 $X2=3.88 $Y2=2.815
r367 5 66 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.745
+ $Y=1.84 $X2=3.88 $Y2=1.985
r368 4 63 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.845
+ $Y=1.84 $X2=2.98 $Y2=2.815
r369 4 60 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.845
+ $Y=1.84 $X2=2.98 $Y2=1.985
r370 3 57 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.945
+ $Y=1.84 $X2=2.08 $Y2=2.815
r371 3 54 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.945
+ $Y=1.84 $X2=2.08 $Y2=1.985
r372 2 51 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.815
r373 2 48 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=1.985
r374 1 45 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r375 1 42 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__CLKINV_16%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 17 18 19 20 63 71 77 81 85 86 89 94 95 97 101 106 111 114 115 120 123 124 125
+ 128 135 142 149 155 162 172 180 188 196 199 204 205 209 210
c322 210 0 1.6166e-19 $X=2.53 $Y=1.885
c323 86 0 1.88851e-19 $X=6.217 $Y=1.638
r324 209 212 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.035
+ $X2=2.53 $Y2=2.035
r325 209 210 3.61044 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=2.53 $Y=1.985
+ $X2=2.53 $Y2=1.885
r326 207 212 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=1.63 $Y=2.035
+ $X2=2.53 $Y2=2.035
r327 204 207 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.63 $Y=2.035
+ $X2=1.63 $Y2=2.035
r328 204 205 4.56265 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.63 $Y=1.985
+ $X2=1.63 $Y2=1.885
r329 196 201 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=10.79 $Y=1.985
+ $X2=10.79 $Y2=2.815
r330 196 199 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.79 $Y=2.035
+ $X2=10.79 $Y2=2.035
r331 191 199 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=9.89 $Y=2.035
+ $X2=10.79 $Y2=2.035
r332 188 193 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=9.89 $Y=1.985
+ $X2=9.89 $Y2=2.815
r333 188 191 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=2.035
+ $X2=9.89 $Y2=2.035
r334 183 191 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=8.99 $Y=2.035
+ $X2=9.89 $Y2=2.035
r335 180 185 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=8.99 $Y=1.985
+ $X2=8.99 $Y2=2.815
r336 180 183 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.99 $Y=2.035
+ $X2=8.99 $Y2=2.035
r337 175 183 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=8.09 $Y=2.035
+ $X2=8.99 $Y2=2.035
r338 172 177 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=8.09 $Y=1.985
+ $X2=8.09 $Y2=2.815
r339 172 175 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.09 $Y=2.035
+ $X2=8.09 $Y2=2.035
r340 167 175 0.596692 $w=2.3e-07 $l=9.3e-07 $layer=MET1_cond $X=7.16 $Y=2.035
+ $X2=8.09 $Y2=2.035
r341 165 169 39.0419 $w=2.43e-07 $l=8.3e-07 $layer=LI1_cond $X=7.167 $Y=1.985
+ $X2=7.167 $Y2=2.815
r342 165 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.16 $Y=2.035
+ $X2=7.16 $Y2=2.035
r343 162 165 64.6779 $w=2.43e-07 $l=1.375e-06 $layer=LI1_cond $X=7.167 $Y=0.61
+ $X2=7.167 $Y2=1.985
r344 157 167 0.628772 $w=2.3e-07 $l=9.8e-07 $layer=MET1_cond $X=6.18 $Y=2.035
+ $X2=7.16 $Y2=2.035
r345 155 159 30.366 $w=3.13e-07 $l=8.3e-07 $layer=LI1_cond $X=6.172 $Y=1.985
+ $X2=6.172 $Y2=2.815
r346 155 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.18 $Y=2.035
+ $X2=6.18 $Y2=2.035
r347 149 152 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=5.23 $Y=2.035
+ $X2=5.23 $Y2=2.815
r348 149 150 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.23 $Y=2.035
+ $X2=5.23 $Y2=2.035
r349 144 150 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=4.33 $Y=2.035
+ $X2=5.23 $Y2=2.035
r350 142 146 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.33 $Y=1.985
+ $X2=4.33 $Y2=2.815
r351 142 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.33 $Y=2.035
+ $X2=4.33 $Y2=2.035
r352 137 144 0.558196 $w=2.3e-07 $l=8.7e-07 $layer=MET1_cond $X=3.46 $Y=2.035
+ $X2=4.33 $Y2=2.035
r353 137 212 0.596692 $w=2.3e-07 $l=9.3e-07 $layer=MET1_cond $X=3.46 $Y=2.035
+ $X2=2.53 $Y2=2.035
r354 135 139 36.7895 $w=2.58e-07 $l=8.3e-07 $layer=LI1_cond $X=3.465 $Y=1.985
+ $X2=3.465 $Y2=2.815
r355 135 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.46 $Y=2.035
+ $X2=3.46 $Y2=2.035
r356 130 207 0.58386 $w=2.3e-07 $l=9.1e-07 $layer=MET1_cond $X=0.72 $Y=2.035
+ $X2=1.63 $Y2=2.035
r357 128 132 48.4498 $w=1.88e-07 $l=8.3e-07 $layer=LI1_cond $X=0.72 $Y=1.985
+ $X2=0.72 $Y2=2.815
r358 128 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=2.035
+ $X2=0.72 $Y2=2.035
r359 125 157 0.272682 $w=2.3e-07 $l=4.25e-07 $layer=MET1_cond $X=5.755 $Y=2.035
+ $X2=6.18 $Y2=2.035
r360 125 150 0.336842 $w=2.3e-07 $l=5.25e-07 $layer=MET1_cond $X=5.755 $Y=2.035
+ $X2=5.23 $Y2=2.035
r361 123 124 13.8636 $w=1.78e-07 $l=2.25e-07 $layer=LI1_cond $X=6.25 $Y=1.01
+ $X2=6.25 $Y2=0.785
r362 122 155 0.292684 $w=3.13e-07 $l=8e-09 $layer=LI1_cond $X=6.172 $Y=1.977
+ $X2=6.172 $Y2=1.985
r363 117 120 2.62582 $w=3.93e-07 $l=9e-08 $layer=LI1_cond $X=5.34 $Y=0.577
+ $X2=5.43 $Y2=0.577
r364 116 149 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=5.23 $Y=2.01
+ $X2=5.23 $Y2=2.035
r365 114 116 0.901327 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=5.245 $Y=1.985
+ $X2=5.245 $Y2=2.01
r366 114 115 7.55066 $w=3.58e-07 $l=1.35e-07 $layer=LI1_cond $X=5.245 $Y=1.985
+ $X2=5.245 $Y2=1.85
r367 111 142 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.33 $Y=1.9
+ $X2=4.33 $Y2=1.985
r368 110 111 2.2967 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=4.345 $Y=1.85
+ $X2=4.345 $Y2=1.9
r369 108 135 53.6329 $w=2.58e-07 $l=1.21e-06 $layer=LI1_cond $X=3.465 $Y=0.775
+ $X2=3.465 $Y2=1.985
r370 106 108 6.63702 $w=2.93e-07 $l=1.65e-07 $layer=LI1_cond $X=3.447 $Y=0.61
+ $X2=3.447 $Y2=0.775
r371 103 210 42.6404 $w=2.98e-07 $l=1.11e-06 $layer=LI1_cond $X=2.515 $Y=0.775
+ $X2=2.515 $Y2=1.885
r372 101 103 6.07341 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=2.507 $Y=0.61
+ $X2=2.507 $Y2=0.775
r373 99 205 55.6179 $w=2.28e-07 $l=1.11e-06 $layer=LI1_cond $X=1.58 $Y=0.775
+ $X2=1.58 $Y2=1.885
r374 97 99 7.49534 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.57 $Y=0.61
+ $X2=1.57 $Y2=0.775
r375 94 128 4.08612 $w=1.88e-07 $l=7e-08 $layer=LI1_cond $X=0.72 $Y=1.915
+ $X2=0.72 $Y2=1.985
r376 94 95 5.58789 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=0.72 $Y=1.915
+ $X2=0.72 $Y2=1.82
r377 93 95 64.3889 $w=1.78e-07 $l=1.045e-06 $layer=LI1_cond $X=0.715 $Y=0.775
+ $X2=0.715 $Y2=1.82
r378 87 124 6.23075 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=6.272 $Y=0.673
+ $X2=6.272 $Y2=0.785
r379 87 89 3.22684 $w=2.23e-07 $l=6.3e-08 $layer=LI1_cond $X=6.272 $Y=0.673
+ $X2=6.272 $Y2=0.61
r380 86 122 15.0393 $w=2.75e-07 $l=3.60799e-07 $layer=LI1_cond $X=6.217 $Y=1.638
+ $X2=6.172 $Y2=1.977
r381 85 123 6.57226 $w=2.43e-07 $l=1.22e-07 $layer=LI1_cond $X=6.217 $Y=1.132
+ $X2=6.217 $Y2=1.01
r382 85 86 23.8015 $w=2.43e-07 $l=5.06e-07 $layer=LI1_cond $X=6.217 $Y=1.132
+ $X2=6.217 $Y2=1.638
r383 83 117 5.70203 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=5.34 $Y=0.775
+ $X2=5.34 $Y2=0.577
r384 83 115 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=5.34 $Y=0.775
+ $X2=5.34 $Y2=1.85
r385 81 110 54.9627 $w=2.58e-07 $l=1.24e-06 $layer=LI1_cond $X=4.395 $Y=0.61
+ $X2=4.395 $Y2=1.85
r386 75 209 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=2.53 $Y=2.05
+ $X2=2.53 $Y2=1.985
r387 75 77 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=2.53 $Y=2.05
+ $X2=2.53 $Y2=2.815
r388 69 204 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=1.63 $Y=2.05
+ $X2=1.63 $Y2=1.985
r389 69 71 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=1.63 $Y=2.05
+ $X2=1.63 $Y2=2.815
r390 61 93 5.58789 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=0.71 $Y=0.68
+ $X2=0.71 $Y2=0.775
r391 61 63 4.08612 $w=1.88e-07 $l=7e-08 $layer=LI1_cond $X=0.71 $Y=0.68 $X2=0.71
+ $Y2=0.61
r392 20 201 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.655
+ $Y=1.84 $X2=10.79 $Y2=2.815
r393 20 196 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.655
+ $Y=1.84 $X2=10.79 $Y2=1.985
r394 19 193 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.755
+ $Y=1.84 $X2=9.89 $Y2=2.815
r395 19 188 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.755
+ $Y=1.84 $X2=9.89 $Y2=1.985
r396 18 185 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.855
+ $Y=1.84 $X2=8.99 $Y2=2.815
r397 18 180 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.855
+ $Y=1.84 $X2=8.99 $Y2=1.985
r398 17 177 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.955
+ $Y=1.84 $X2=8.09 $Y2=2.815
r399 17 172 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.955
+ $Y=1.84 $X2=8.09 $Y2=1.985
r400 16 169 400 $w=1.7e-07 $l=1.05428e-06 $layer=licon1_PDIFF $count=1 $X=6.995
+ $Y=1.84 $X2=7.16 $Y2=2.815
r401 16 165 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=6.995
+ $Y=1.84 $X2=7.16 $Y2=1.985
r402 15 159 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.045
+ $Y=1.84 $X2=6.18 $Y2=2.815
r403 15 155 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.045
+ $Y=1.84 $X2=6.18 $Y2=1.985
r404 14 152 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.095
+ $Y=1.84 $X2=5.23 $Y2=2.815
r405 14 114 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.095
+ $Y=1.84 $X2=5.23 $Y2=1.985
r406 13 146 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.195
+ $Y=1.84 $X2=4.33 $Y2=2.815
r407 13 142 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.195
+ $Y=1.84 $X2=4.33 $Y2=1.985
r408 12 139 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.295
+ $Y=1.84 $X2=3.43 $Y2=2.815
r409 12 135 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.295
+ $Y=1.84 $X2=3.43 $Y2=1.985
r410 11 209 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.395
+ $Y=1.84 $X2=2.53 $Y2=1.985
r411 11 77 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.395
+ $Y=1.84 $X2=2.53 $Y2=2.815
r412 10 204 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.84 $X2=1.63 $Y2=1.985
r413 10 71 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.84 $X2=1.63 $Y2=2.815
r414 9 132 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.815
r415 9 128 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=1.985
r416 8 162 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.01
+ $Y=0.4 $X2=7.15 $Y2=0.61
r417 7 89 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.15
+ $Y=0.4 $X2=6.29 $Y2=0.61
r418 6 120 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.29
+ $Y=0.4 $X2=5.43 $Y2=0.61
r419 5 81 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.29
+ $Y=0.4 $X2=4.43 $Y2=0.61
r420 4 106 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.29
+ $Y=0.4 $X2=3.43 $Y2=0.61
r421 3 101 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.36
+ $Y=0.4 $X2=2.5 $Y2=0.61
r422 2 97 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.43
+ $Y=0.4 $X2=1.57 $Y2=0.61
r423 1 63 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.4 $X2=0.71 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_MS__CLKINV_16%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46
+ 50 54 58 61 62 64 65 67 68 70 71 73 74 76 77 79 80 82 85 86 114 122 123 130
c146 30 0 1.45923e-19 $X=0.28 $Y=0.61
r147 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r148 129 132 4.06215 $w=7.93e-07 $l=2.7e-07 $layer=LI1_cond $X=7.65 $Y=0.312
+ $X2=7.92 $Y2=0.312
r149 129 130 11.4033 $w=7.93e-07 $l=1.65e-07 $layer=LI1_cond $X=7.65 $Y=0.312
+ $X2=7.485 $Y2=0.312
r150 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r151 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r152 120 123 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=11.28 $Y2=0
r153 119 122 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=9.84 $Y=0
+ $X2=11.28 $Y2=0
r154 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r155 117 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r156 117 133 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=7.92 $Y2=0
r157 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r158 114 132 5.4162 $w=7.93e-07 $l=3.6e-07 $layer=LI1_cond $X=8.28 $Y=0.312
+ $X2=7.92 $Y2=0.312
r159 114 116 16.2486 $w=7.93e-07 $l=1.08e-06 $layer=LI1_cond $X=8.28 $Y=0.312
+ $X2=9.36 $Y2=0.312
r160 113 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r161 112 130 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=7.44 $Y=0
+ $X2=7.485 $Y2=0
r162 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r163 109 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=7.44 $Y2=0
r164 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r165 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r166 103 106 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.52 $Y2=0
r167 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r168 100 103 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0
+ $X2=4.56 $Y2=0
r169 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r170 97 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r171 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r172 94 97 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r173 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r174 91 94 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r175 91 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r176 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r177 88 126 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r178 88 90 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r179 86 109 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=6.48 $Y2=0
r180 86 106 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=5.52 $Y2=0
r181 85 119 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=9.825 $Y=0
+ $X2=9.84 $Y2=0
r182 84 85 11.4033 $w=7.93e-07 $l=1.65e-07 $layer=LI1_cond $X=9.66 $Y=0.312
+ $X2=9.825 $Y2=0.312
r183 82 116 1.02306 $w=7.93e-07 $l=6.8e-08 $layer=LI1_cond $X=9.428 $Y=0.312
+ $X2=9.36 $Y2=0.312
r184 82 84 3.49044 $w=7.93e-07 $l=2.32e-07 $layer=LI1_cond $X=9.428 $Y=0.312
+ $X2=9.66 $Y2=0.312
r185 79 108 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.555 $Y=0
+ $X2=6.48 $Y2=0
r186 79 80 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=6.555 $Y=0 $X2=6.715
+ $Y2=0
r187 78 112 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=6.875 $Y=0
+ $X2=7.44 $Y2=0
r188 78 80 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=6.875 $Y=0 $X2=6.715
+ $Y2=0
r189 76 105 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.695 $Y=0
+ $X2=5.52 $Y2=0
r190 76 77 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=5.695 $Y=0
+ $X2=5.837 $Y2=0
r191 75 108 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=5.98 $Y=0 $X2=6.48
+ $Y2=0
r192 75 77 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=5.98 $Y=0 $X2=5.837
+ $Y2=0
r193 73 102 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.765 $Y=0
+ $X2=4.56 $Y2=0
r194 73 74 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=4.765 $Y=0 $X2=4.925
+ $Y2=0
r195 72 105 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=5.085 $Y=0
+ $X2=5.52 $Y2=0
r196 72 74 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=5.085 $Y=0 $X2=4.925
+ $Y2=0
r197 70 99 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.765 $Y=0 $X2=3.6
+ $Y2=0
r198 70 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.765 $Y=0 $X2=3.93
+ $Y2=0
r199 69 102 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=4.095 $Y=0
+ $X2=4.56 $Y2=0
r200 69 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.095 $Y=0 $X2=3.93
+ $Y2=0
r201 67 96 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.845 $Y=0
+ $X2=2.64 $Y2=0
r202 67 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.845 $Y=0 $X2=2.97
+ $Y2=0
r203 66 99 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=3.095 $Y=0 $X2=3.6
+ $Y2=0
r204 66 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.095 $Y=0 $X2=2.97
+ $Y2=0
r205 64 93 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.885 $Y=0
+ $X2=1.68 $Y2=0
r206 64 65 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.885 $Y=0 $X2=2.025
+ $Y2=0
r207 63 96 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.165 $Y=0
+ $X2=2.64 $Y2=0
r208 63 65 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.165 $Y=0 $X2=2.025
+ $Y2=0
r209 61 90 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0
+ $X2=0.72 $Y2=0
r210 61 62 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=0.975 $Y=0
+ $X2=1.117 $Y2=0
r211 60 93 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.68
+ $Y2=0
r212 60 62 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.117
+ $Y2=0
r213 56 80 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=6.715 $Y=0.085
+ $X2=6.715 $Y2=0
r214 56 58 18.9073 $w=3.18e-07 $l=5.25e-07 $layer=LI1_cond $X=6.715 $Y=0.085
+ $X2=6.715 $Y2=0.61
r215 52 77 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=5.837 $Y=0.085
+ $X2=5.837 $Y2=0
r216 52 54 21.2292 $w=2.83e-07 $l=5.25e-07 $layer=LI1_cond $X=5.837 $Y=0.085
+ $X2=5.837 $Y2=0.61
r217 48 74 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.925 $Y=0.085
+ $X2=4.925 $Y2=0
r218 48 50 18.9073 $w=3.18e-07 $l=5.25e-07 $layer=LI1_cond $X=4.925 $Y=0.085
+ $X2=4.925 $Y2=0.61
r219 44 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.93 $Y=0.085
+ $X2=3.93 $Y2=0
r220 44 46 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=3.93 $Y=0.085
+ $X2=3.93 $Y2=0.61
r221 40 68 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=0.085
+ $X2=2.97 $Y2=0
r222 40 42 24.2013 $w=2.48e-07 $l=5.25e-07 $layer=LI1_cond $X=2.97 $Y=0.085
+ $X2=2.97 $Y2=0.61
r223 36 65 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0
r224 36 38 21.6083 $w=2.78e-07 $l=5.25e-07 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0.61
r225 32 62 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.117 $Y=0.085
+ $X2=1.117 $Y2=0
r226 32 34 21.2292 $w=2.83e-07 $l=5.25e-07 $layer=LI1_cond $X=1.117 $Y=0.085
+ $X2=1.117 $Y2=0.61
r227 28 126 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r228 28 30 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.61
r229 9 129 60.6667 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=3
+ $X=7.44 $Y=0.4 $X2=7.65 $Y2=0.545
r230 9 84 60.6667 $w=1.7e-07 $l=2.29135e-06 $layer=licon1_NDIFF $count=3 $X=7.44
+ $Y=0.4 $X2=9.66 $Y2=0.545
r231 8 58 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.58
+ $Y=0.4 $X2=6.72 $Y2=0.61
r232 7 54 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.72
+ $Y=0.4 $X2=5.86 $Y2=0.61
r233 6 50 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=4.72
+ $Y=0.4 $X2=4.93 $Y2=0.61
r234 5 46 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=3.72
+ $Y=0.4 $X2=3.93 $Y2=0.61
r235 4 42 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.79
+ $Y=0.4 $X2=2.93 $Y2=0.61
r236 3 38 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.4 $X2=2 $Y2=0.61
r237 2 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1 $Y=0.4
+ $X2=1.14 $Y2=0.61
r238 1 30 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.4 $X2=0.28 $Y2=0.61
.ends


* File: sky130_fd_sc_ms__xnor2_4.pex.spice
* Created: Wed Sep  2 12:33:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__XNOR2_4%A 3 7 11 15 19 23 27 31 35 37 39 40 42 44 46
+ 52 54 55 58 61 67 77 90
c189 55 0 1.57454e-19 $X=1.345 $Y=1.665
c190 44 0 9.06279e-20 $X=6.815 $Y=1.725
c191 42 0 3.01101e-20 $X=6.55 $Y=0.74
c192 35 0 3.01101e-20 $X=5.96 $Y=0.74
c193 27 0 3.01105e-20 $X=5.53 $Y=0.74
c194 7 0 7.39126e-20 $X=0.495 $Y=0.69
r195 79 80 40.1667 $w=2.82e-07 $l=2.35e-07 $layer=POLY_cond $X=5.96 $Y=1.537
+ $X2=6.195 $Y2=1.537
r196 78 79 36.7482 $w=2.82e-07 $l=2.15e-07 $layer=POLY_cond $X=5.745 $Y=1.537
+ $X2=5.96 $Y2=1.537
r197 76 78 12.8191 $w=2.82e-07 $l=7.5e-08 $layer=POLY_cond $X=5.67 $Y=1.537
+ $X2=5.745 $Y2=1.537
r198 76 77 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.67
+ $Y=1.515 $X2=5.67 $Y2=1.515
r199 74 76 23.9291 $w=2.82e-07 $l=1.4e-07 $layer=POLY_cond $X=5.53 $Y=1.537
+ $X2=5.67 $Y2=1.537
r200 73 74 70.078 $w=2.82e-07 $l=4.1e-07 $layer=POLY_cond $X=5.12 $Y=1.537
+ $X2=5.53 $Y2=1.537
r201 72 77 18.4391 $w=4.23e-07 $l=6.8e-07 $layer=LI1_cond $X=4.99 $Y=1.562
+ $X2=5.67 $Y2=1.562
r202 71 73 22.2199 $w=2.82e-07 $l=1.3e-07 $layer=POLY_cond $X=4.99 $Y=1.537
+ $X2=5.12 $Y2=1.537
r203 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.99
+ $Y=1.515 $X2=4.99 $Y2=1.515
r204 69 71 8.5461 $w=2.82e-07 $l=5e-08 $layer=POLY_cond $X=4.94 $Y=1.537
+ $X2=4.99 $Y2=1.537
r205 67 68 5.96904 $w=3.23e-07 $l=4e-08 $layer=POLY_cond $X=0.955 $Y=1.485
+ $X2=0.995 $Y2=1.485
r206 64 65 1.49226 $w=3.23e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.485
+ $X2=0.505 $Y2=1.485
r207 58 90 3.96409 $w=4.58e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.55
+ $X2=1.085 $Y2=1.55
r208 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=1.665
+ $X2=1.2 $Y2=1.665
r209 55 57 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=1.665
+ $X2=1.2 $Y2=1.665
r210 54 61 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.415 $Y=1.665
+ $X2=4.56 $Y2=1.665
r211 54 55 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=4.415 $Y=1.665
+ $X2=1.345 $Y2=1.665
r212 52 72 11.66 $w=4.23e-07 $l=4.3e-07 $layer=LI1_cond $X=4.56 $Y=1.562
+ $X2=4.99 $Y2=1.562
r213 52 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=1.665
+ $X2=4.56 $Y2=1.665
r214 50 67 36.5604 $w=3.23e-07 $l=2.45e-07 $layer=POLY_cond $X=0.71 $Y=1.485
+ $X2=0.955 $Y2=1.485
r215 50 65 30.5913 $w=3.23e-07 $l=2.05e-07 $layer=POLY_cond $X=0.71 $Y=1.485
+ $X2=0.505 $Y2=1.485
r216 49 90 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=0.71 $Y=1.485
+ $X2=1.085 $Y2=1.485
r217 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.71
+ $Y=1.485 $X2=0.71 $Y2=1.485
r218 44 46 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=6.815 $Y=1.725
+ $X2=6.815 $Y2=2.4
r219 40 44 45.2943 $w=2.82e-07 $l=3.46475e-07 $layer=POLY_cond $X=6.55 $Y=1.537
+ $X2=6.815 $Y2=1.725
r220 40 80 60.6773 $w=2.82e-07 $l=3.55e-07 $layer=POLY_cond $X=6.55 $Y=1.537
+ $X2=6.195 $Y2=1.537
r221 40 42 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=6.55 $Y=1.425
+ $X2=6.55 $Y2=0.74
r222 37 80 13.2911 $w=1.8e-07 $l=1.88e-07 $layer=POLY_cond $X=6.195 $Y=1.725
+ $X2=6.195 $Y2=1.537
r223 37 39 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=6.195 $Y=1.725
+ $X2=6.195 $Y2=2.4
r224 33 79 17.5183 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=5.96 $Y=1.35
+ $X2=5.96 $Y2=1.537
r225 33 35 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.96 $Y=1.35
+ $X2=5.96 $Y2=0.74
r226 29 78 13.2911 $w=1.8e-07 $l=1.43e-07 $layer=POLY_cond $X=5.745 $Y=1.68
+ $X2=5.745 $Y2=1.537
r227 29 31 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.745 $Y=1.68
+ $X2=5.745 $Y2=2.4
r228 25 74 17.5183 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=5.53 $Y=1.35
+ $X2=5.53 $Y2=1.537
r229 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.53 $Y=1.35
+ $X2=5.53 $Y2=0.74
r230 21 73 13.2911 $w=1.8e-07 $l=1.43e-07 $layer=POLY_cond $X=5.12 $Y=1.68
+ $X2=5.12 $Y2=1.537
r231 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.12 $Y=1.68
+ $X2=5.12 $Y2=2.4
r232 17 69 17.5183 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=4.94 $Y=1.35
+ $X2=4.94 $Y2=1.537
r233 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.94 $Y=1.35
+ $X2=4.94 $Y2=0.74
r234 13 68 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.32
+ $X2=0.995 $Y2=1.485
r235 13 15 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.995 $Y=1.32
+ $X2=0.995 $Y2=0.69
r236 9 67 16.4327 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.65
+ $X2=0.955 $Y2=1.485
r237 9 11 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=0.955 $Y=1.65
+ $X2=0.955 $Y2=2.26
r238 5 64 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.32
+ $X2=0.495 $Y2=1.485
r239 5 7 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.495 $Y=1.32
+ $X2=0.495 $Y2=0.69
r240 1 65 16.4327 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.65
+ $X2=0.505 $Y2=1.485
r241 1 3 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=0.505 $Y=1.65
+ $X2=0.505 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR2_4%B 3 7 11 15 17 19 22 26 30 34 38 40 41 44 48
+ 50 53 54 55 56 57 58 60 61 62 63 64 65 87
c202 53 0 8.76351e-20 $X=2.07 $Y=1.68
c203 34 0 3.01101e-20 $X=8.035 $Y=0.74
c204 26 0 3.01105e-20 $X=7.605 $Y=0.74
c205 17 0 3.01105e-20 $X=6.98 $Y=1.185
c206 15 0 1.04341e-19 $X=1.925 $Y=0.69
r207 86 87 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.99
+ $Y=1.515 $X2=7.99 $Y2=1.515
r208 84 86 41.9462 $w=3.16e-07 $l=2.75e-07 $layer=POLY_cond $X=7.715 $Y=1.432
+ $X2=7.99 $Y2=1.432
r209 81 82 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.31
+ $Y=1.515 $X2=7.31 $Y2=1.515
r210 79 81 6.86392 $w=3.16e-07 $l=4.5e-08 $layer=POLY_cond $X=7.265 $Y=1.432
+ $X2=7.31 $Y2=1.432
r211 74 75 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=1.855 $Y=1.515
+ $X2=1.925 $Y2=1.515
r212 73 74 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.425 $Y=1.515
+ $X2=1.855 $Y2=1.515
r213 71 73 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.405 $Y=1.515
+ $X2=1.425 $Y2=1.515
r214 65 87 1.94388 $w=4.13e-07 $l=7e-08 $layer=LI1_cond $X=7.92 $Y=1.557
+ $X2=7.99 $Y2=1.557
r215 64 65 13.3295 $w=4.13e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.557
+ $X2=7.92 $Y2=1.557
r216 64 82 3.61006 $w=4.13e-07 $l=1.3e-07 $layer=LI1_cond $X=7.44 $Y=1.557
+ $X2=7.31 $Y2=1.557
r217 63 82 9.7194 $w=4.13e-07 $l=3.5e-07 $layer=LI1_cond $X=6.96 $Y=1.557
+ $X2=7.31 $Y2=1.557
r218 62 90 2.46632 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=6.45 $Y=1.557
+ $X2=6.535 $Y2=1.557
r219 62 63 11.3856 $w=4.13e-07 $l=4.1e-07 $layer=LI1_cond $X=6.55 $Y=1.557
+ $X2=6.96 $Y2=1.557
r220 62 90 0.416546 $w=4.13e-07 $l=1.5e-08 $layer=LI1_cond $X=6.55 $Y=1.557
+ $X2=6.535 $Y2=1.557
r221 61 75 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=1.99 $Y=1.515
+ $X2=1.925 $Y2=1.515
r222 60 61 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.99
+ $Y=1.515 $X2=1.99 $Y2=1.515
r223 57 62 6.03523 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=6.45 $Y=1.765
+ $X2=6.45 $Y2=1.557
r224 57 58 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.45 $Y=1.765
+ $X2=6.45 $Y2=1.945
r225 55 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.365 $Y=2.03
+ $X2=6.45 $Y2=1.945
r226 55 56 274.663 $w=1.68e-07 $l=4.21e-06 $layer=LI1_cond $X=6.365 $Y=2.03
+ $X2=2.155 $Y2=2.03
r227 54 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.07 $Y=1.945
+ $X2=2.155 $Y2=2.03
r228 53 60 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.07 $Y=1.68
+ $X2=2.07 $Y2=1.515
r229 53 54 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.07 $Y=1.68
+ $X2=2.07 $Y2=1.945
r230 46 50 18.8402 $w=1.65e-07 $l=7.98436e-08 $layer=POLY_cond $X=8.625 $Y=1.35
+ $X2=8.615 $Y2=1.425
r231 46 48 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.625 $Y=1.35
+ $X2=8.625 $Y2=0.74
r232 42 50 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=8.615 $Y=1.5
+ $X2=8.615 $Y2=1.425
r233 42 44 349.839 $w=1.8e-07 $l=9e-07 $layer=POLY_cond $X=8.615 $Y=1.5
+ $X2=8.615 $Y2=2.4
r234 41 89 27.0984 $w=3.16e-07 $l=9.34345e-08 $layer=POLY_cond $X=8.255 $Y=1.425
+ $X2=8.165 $Y2=1.432
r235 40 50 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.525 $Y=1.425
+ $X2=8.615 $Y2=1.425
r236 40 41 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=8.525 $Y=1.425
+ $X2=8.255 $Y2=1.425
r237 36 89 15.9236 $w=1.8e-07 $l=2.48e-07 $layer=POLY_cond $X=8.165 $Y=1.68
+ $X2=8.165 $Y2=1.432
r238 36 38 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.165 $Y=1.68
+ $X2=8.165 $Y2=2.4
r239 32 89 19.8291 $w=3.16e-07 $l=1.3e-07 $layer=POLY_cond $X=8.035 $Y=1.432
+ $X2=8.165 $Y2=1.432
r240 32 86 6.86392 $w=3.16e-07 $l=4.5e-08 $layer=POLY_cond $X=8.035 $Y=1.432
+ $X2=7.99 $Y2=1.432
r241 32 34 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.035 $Y=1.35
+ $X2=8.035 $Y2=0.74
r242 28 84 15.9236 $w=1.8e-07 $l=2.48e-07 $layer=POLY_cond $X=7.715 $Y=1.68
+ $X2=7.715 $Y2=1.432
r243 28 30 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.715 $Y=1.68
+ $X2=7.715 $Y2=2.4
r244 24 84 16.7785 $w=3.16e-07 $l=1.1e-07 $layer=POLY_cond $X=7.605 $Y=1.432
+ $X2=7.715 $Y2=1.432
r245 24 81 44.9968 $w=3.16e-07 $l=2.95e-07 $layer=POLY_cond $X=7.605 $Y=1.432
+ $X2=7.31 $Y2=1.432
r246 24 26 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.605 $Y=1.35
+ $X2=7.605 $Y2=0.74
r247 20 79 15.9236 $w=1.8e-07 $l=2.48e-07 $layer=POLY_cond $X=7.265 $Y=1.68
+ $X2=7.265 $Y2=1.432
r248 20 22 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.265 $Y=1.68
+ $X2=7.265 $Y2=2.4
r249 17 79 43.4715 $w=3.16e-07 $l=3.89384e-07 $layer=POLY_cond $X=6.98 $Y=1.185
+ $X2=7.265 $Y2=1.432
r250 17 19 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=6.98 $Y=1.185
+ $X2=6.98 $Y2=0.74
r251 13 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.35
+ $X2=1.925 $Y2=1.515
r252 13 15 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.925 $Y=1.35
+ $X2=1.925 $Y2=0.69
r253 9 74 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.68
+ $X2=1.855 $Y2=1.515
r254 9 11 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=1.855 $Y=1.68
+ $X2=1.855 $Y2=2.26
r255 5 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=1.515
r256 5 7 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=0.69
r257 1 71 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.68
+ $X2=1.405 $Y2=1.515
r258 1 3 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=1.405 $Y=1.68
+ $X2=1.405 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR2_4%A_119_368# 1 2 3 12 16 20 24 28 31 32 36 38
+ 39 41 42 45 47 48 50 51 54 57 60 62 63 66 70 80 83
c172 57 0 1.20688e-19 $X=3.92 $Y=1.515
c173 54 0 9.22535e-20 $X=2.48 $Y=1.35
r174 91 92 83.9334 $w=3.3e-07 $l=4.8e-07 $layer=POLY_cond $X=2.935 $Y=1.515
+ $X2=3.415 $Y2=1.515
r175 90 91 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.915 $Y=1.515
+ $X2=2.935 $Y2=1.515
r176 83 92 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.49 $Y=1.515
+ $X2=3.415 $Y2=1.515
r177 78 80 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.745 $Y=2.79
+ $X2=3.58 $Y2=2.79
r178 78 79 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.745
+ $Y=2.79 $X2=3.745 $Y2=2.79
r179 76 90 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.56 $Y=1.515
+ $X2=2.915 $Y2=1.515
r180 76 87 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.56 $Y=1.515
+ $X2=2.485 $Y2=1.515
r181 75 76 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.56
+ $Y=1.515 $X2=2.56 $Y2=1.515
r182 70 72 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.71 $Y=0.86
+ $X2=1.71 $Y2=1.095
r183 62 63 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.425
+ $Y=2.79 $X2=4.425 $Y2=2.79
r184 60 78 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.91 $Y=2.79
+ $X2=3.745 $Y2=2.79
r185 60 62 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=3.91 $Y=2.79
+ $X2=4.425 $Y2=2.79
r186 58 83 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.92 $Y=1.515
+ $X2=3.49 $Y2=1.515
r187 57 58 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.92
+ $Y=1.515 $X2=3.92 $Y2=1.515
r188 55 75 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.565 $Y=1.515
+ $X2=2.48 $Y2=1.515
r189 55 57 47.32 $w=3.28e-07 $l=1.355e-06 $layer=LI1_cond $X=2.565 $Y=1.515
+ $X2=3.92 $Y2=1.515
r190 54 75 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.48 $Y=1.35
+ $X2=2.48 $Y2=1.515
r191 53 54 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.48 $Y=1.18
+ $X2=2.48 $Y2=1.35
r192 52 72 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=1.095
+ $X2=1.71 $Y2=1.095
r193 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.395 $Y=1.095
+ $X2=2.48 $Y2=1.18
r194 51 52 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.395 $Y=1.095
+ $X2=1.875 $Y2=1.095
r195 50 80 116.455 $w=1.68e-07 $l=1.785e-06 $layer=LI1_cond $X=1.795 $Y=2.71
+ $X2=3.58 $Y2=2.71
r196 48 50 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.63 $Y=2.625
+ $X2=1.795 $Y2=2.71
r197 47 68 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=2.12 $X2=1.63
+ $Y2=2.035
r198 47 48 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=1.63 $Y=2.12
+ $X2=1.63 $Y2=2.625
r199 46 66 4.70058 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=0.895 $Y=2.035
+ $X2=0.73 $Y2=1.97
r200 45 68 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=2.035
+ $X2=1.63 $Y2=2.035
r201 45 46 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.465 $Y=2.035
+ $X2=0.895 $Y2=2.035
r202 41 79 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=3.935 $Y=2.79
+ $X2=3.745 $Y2=2.79
r203 41 42 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.935 $Y=2.79
+ $X2=4.01 $Y2=2.79
r204 40 63 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.085 $Y=2.79
+ $X2=4.425 $Y2=2.79
r205 40 42 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.085 $Y=2.79
+ $X2=4.01 $Y2=2.79
r206 38 58 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.935 $Y=1.515
+ $X2=3.92 $Y2=1.515
r207 38 39 6.91837 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.935 $Y=1.515
+ $X2=4.01 $Y2=1.515
r208 34 36 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.44 $Y=1.35
+ $X2=4.44 $Y2=0.74
r209 33 39 6.91837 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.085 $Y=1.425
+ $X2=4.01 $Y2=1.515
r210 32 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.365 $Y=1.425
+ $X2=4.44 $Y2=1.35
r211 32 33 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.365 $Y=1.425
+ $X2=4.085 $Y2=1.425
r212 31 42 16.9349 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.01 $Y=2.625
+ $X2=4.01 $Y2=2.79
r213 30 39 18.1359 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.01 $Y=1.68
+ $X2=4.01 $Y2=1.515
r214 30 31 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=4.01 $Y=1.68
+ $X2=4.01 $Y2=2.625
r215 26 39 18.1359 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.01 $Y=1.35
+ $X2=4.01 $Y2=1.515
r216 26 28 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.01 $Y=1.35
+ $X2=4.01 $Y2=0.74
r217 22 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.415 $Y=1.35
+ $X2=3.415 $Y2=1.515
r218 22 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.415 $Y=1.35
+ $X2=3.415 $Y2=0.74
r219 18 91 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.935 $Y=1.68
+ $X2=2.935 $Y2=1.515
r220 18 20 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.935 $Y=1.68
+ $X2=2.935 $Y2=2.4
r221 14 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=1.35
+ $X2=2.915 $Y2=1.515
r222 14 16 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.915 $Y=1.35
+ $X2=2.915 $Y2=0.74
r223 10 87 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.485 $Y=1.68
+ $X2=2.485 $Y2=1.515
r224 10 12 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.485 $Y=1.68
+ $X2=2.485 $Y2=2.4
r225 3 68 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.84 $X2=1.63 $Y2=2.115
r226 2 66 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=1.985
r227 1 70 182 $w=1.7e-07 $l=5.85662e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.71 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR2_4%VPWR 1 2 3 4 5 6 19 21 25 27 30 31 33 36 39
+ 45 56 65 66 72 79 86
r111 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r112 86 89 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=6.505 $Y=3.05
+ $X2=6.505 $Y2=3.33
r113 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r114 79 82 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=3.245 $Y=3.05
+ $X2=3.245 $Y2=3.33
r115 76 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r116 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r117 72 75 9.49071 $w=3.38e-07 $l=2.8e-07 $layer=LI1_cond $X=2.17 $Y=3.05
+ $X2=2.17 $Y2=3.33
r118 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r119 65 66 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r120 63 66 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.88 $Y2=3.33
r121 63 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r122 62 65 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=8.88 $Y2=3.33
r123 62 63 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r124 60 89 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.67 $Y=3.33
+ $X2=6.505 $Y2=3.33
r125 60 62 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.67 $Y=3.33
+ $X2=6.96 $Y2=3.33
r126 59 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r127 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r128 56 89 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.34 $Y=3.33
+ $X2=6.505 $Y2=3.33
r129 56 58 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.34 $Y=3.33 $X2=6
+ $Y2=3.33
r130 55 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r131 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r132 52 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r133 51 54 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r134 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r135 49 82 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.41 $Y=3.33
+ $X2=3.245 $Y2=3.33
r136 49 51 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.41 $Y=3.33
+ $X2=3.6 $Y2=3.33
r137 48 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r138 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r139 45 75 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2 $Y=3.33 $X2=2.17
+ $Y2=3.33
r140 45 47 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2 $Y=3.33 $X2=1.68
+ $Y2=3.33
r141 44 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r142 44 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r143 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r144 41 69 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r145 41 43 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r146 39 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r147 39 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=3.6 $Y2=3.33
r148 37 58 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=5.6 $Y=3.33 $X2=6
+ $Y2=3.33
r149 36 54 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.265 $Y=3.33
+ $X2=5.04 $Y2=3.33
r150 36 37 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=5.432 $Y=3.33
+ $X2=5.6 $Y2=3.33
r151 33 36 9.63236 $w=3.33e-07 $l=2.8e-07 $layer=LI1_cond $X=5.432 $Y=3.05
+ $X2=5.432 $Y2=3.33
r152 30 43 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.72 $Y2=3.33
r153 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.18 $Y2=3.33
r154 29 47 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.68 $Y2=3.33
r155 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.18 $Y2=3.33
r156 28 75 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.34 $Y=3.33
+ $X2=2.17 $Y2=3.33
r157 27 82 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=3.33
+ $X2=3.245 $Y2=3.33
r158 27 28 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=3.08 $Y=3.33
+ $X2=2.34 $Y2=3.33
r159 23 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r160 23 25 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.495
r161 19 69 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r162 19 21 58.0831 $w=2.48e-07 $l=1.26e-06 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=1.985
r163 6 86 600 $w=1.7e-07 $l=1.31541e-06 $layer=licon1_PDIFF $count=1 $X=6.285
+ $Y=1.84 $X2=6.505 $Y2=3.05
r164 5 33 600 $w=1.7e-07 $l=1.31541e-06 $layer=licon1_PDIFF $count=1 $X=5.21
+ $Y=1.84 $X2=5.43 $Y2=3.05
r165 4 79 600 $w=1.7e-07 $l=1.31541e-06 $layer=licon1_PDIFF $count=1 $X=3.025
+ $Y=1.84 $X2=3.245 $Y2=3.05
r166 3 72 600 $w=1.7e-07 $l=1.31771e-06 $layer=licon1_PDIFF $count=1 $X=1.945
+ $Y=1.84 $X2=2.17 $Y2=3.05
r167 2 25 600 $w=1.7e-07 $l=7.1934e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.495
r168 1 21 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR2_4%Y 1 2 3 4 5 16 22 24 25 28 30 32 37 38 41 42
+ 45
r127 42 45 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.49 $Y=2.02 $X2=7.49
+ $Y2=2.105
r128 42 45 0.244458 $w=3.28e-07 $l=7e-09 $layer=LI1_cond $X=7.49 $Y=2.112
+ $X2=7.49 $Y2=2.105
r129 39 42 6.04159 $w=3.28e-07 $l=1.73e-07 $layer=LI1_cond $X=7.49 $Y=2.285
+ $X2=7.49 $Y2=2.112
r130 37 41 3.70735 $w=2.5e-07 $l=9.44722e-08 $layer=LI1_cond $X=8.41 $Y=1.935
+ $X2=8.39 $Y2=2.02
r131 36 37 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=8.41 $Y=1.18
+ $X2=8.41 $Y2=1.935
r132 33 42 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.655 $Y=2.02
+ $X2=7.49 $Y2=2.02
r133 32 41 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.225 $Y=2.02
+ $X2=8.39 $Y2=2.02
r134 32 33 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.225 $Y=2.02
+ $X2=7.655 $Y2=2.02
r135 31 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.39 $Y=1.095
+ $X2=4.225 $Y2=1.095
r136 30 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.325 $Y=1.095
+ $X2=8.41 $Y2=1.18
r137 30 31 256.722 $w=1.68e-07 $l=3.935e-06 $layer=LI1_cond $X=8.325 $Y=1.095
+ $X2=4.39 $Y2=1.095
r138 26 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.225 $Y=1.01
+ $X2=4.225 $Y2=1.095
r139 26 28 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.225 $Y=1.01
+ $X2=4.225 $Y2=0.86
r140 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.06 $Y=1.095
+ $X2=4.225 $Y2=1.095
r141 24 25 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.06 $Y=1.095
+ $X2=3.365 $Y2=1.095
r142 20 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.2 $Y=1.01
+ $X2=3.365 $Y2=1.095
r143 20 22 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.2 $Y=1.01 $X2=3.2
+ $Y2=0.86
r144 16 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.325 $Y=2.37
+ $X2=7.49 $Y2=2.285
r145 16 18 301.086 $w=1.68e-07 $l=4.615e-06 $layer=LI1_cond $X=7.325 $Y=2.37
+ $X2=2.71 $Y2=2.37
r146 5 41 300 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_PDIFF $count=2 $X=8.255
+ $Y=1.84 $X2=8.39 $Y2=2.1
r147 4 42 300 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_PDIFF $count=2 $X=7.355
+ $Y=1.84 $X2=7.49 $Y2=2.1
r148 3 18 600 $w=1.7e-07 $l=5.93675e-07 $layer=licon1_PDIFF $count=1 $X=2.575
+ $Y=1.84 $X2=2.71 $Y2=2.37
r149 2 28 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=4.085
+ $Y=0.37 $X2=4.225 $Y2=0.86
r150 1 22 182 $w=1.7e-07 $l=5.85662e-07 $layer=licon1_NDIFF $count=1 $X=2.99
+ $Y=0.37 $X2=3.2 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR2_4%A_950_368# 1 2 3 4 5 18 20 24 26 30 34 41 42
+ 43 49
c66 20 0 9.06279e-20 $X=7.855 $Y=2.99
r67 46 47 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=7 $Y=2.8 $X2=7
+ $Y2=2.99
r68 43 46 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=7 $Y=2.71 $X2=7
+ $Y2=2.8
r69 40 42 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=5.97 $Y=2.802
+ $X2=6.135 $Y2=2.802
r70 40 41 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=5.97 $Y=2.802
+ $X2=5.805 $Y2=2.802
r71 34 37 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.935 $Y=2.71
+ $X2=4.935 $Y2=2.8
r72 30 33 32.9599 $w=2.48e-07 $l=7.15e-07 $layer=LI1_cond $X=8.88 $Y=2.1
+ $X2=8.88 $Y2=2.815
r73 28 33 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=8.88 $Y=2.905 $X2=8.88
+ $Y2=2.815
r74 27 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.025 $Y=2.99
+ $X2=7.94 $Y2=2.99
r75 26 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.755 $Y=2.99
+ $X2=8.88 $Y2=2.905
r76 26 27 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=8.755 $Y=2.99
+ $X2=8.025 $Y2=2.99
r77 22 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.94 $Y=2.905
+ $X2=7.94 $Y2=2.99
r78 22 24 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=7.94 $Y=2.905
+ $X2=7.94 $Y2=2.44
r79 21 47 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.125 $Y=2.99 $X2=7
+ $Y2=2.99
r80 20 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.855 $Y=2.99
+ $X2=7.94 $Y2=2.99
r81 20 21 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.855 $Y=2.99
+ $X2=7.125 $Y2=2.99
r82 18 43 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.875 $Y=2.71 $X2=7
+ $Y2=2.71
r83 18 42 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=6.875 $Y=2.71
+ $X2=6.135 $Y2=2.71
r84 17 34 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.06 $Y=2.71
+ $X2=4.935 $Y2=2.71
r85 17 41 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=5.06 $Y=2.71
+ $X2=5.805 $Y2=2.71
r86 5 33 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.705
+ $Y=1.84 $X2=8.84 $Y2=2.815
r87 5 30 400 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_PDIFF $count=1 $X=8.705
+ $Y=1.84 $X2=8.84 $Y2=2.1
r88 4 24 300 $w=1.7e-07 $l=6.64078e-07 $layer=licon1_PDIFF $count=2 $X=7.805
+ $Y=1.84 $X2=7.94 $Y2=2.44
r89 3 46 600 $w=1.7e-07 $l=1.02528e-06 $layer=licon1_PDIFF $count=1 $X=6.905
+ $Y=1.84 $X2=7.04 $Y2=2.8
r90 2 40 600 $w=1.7e-07 $l=1.02528e-06 $layer=licon1_PDIFF $count=1 $X=5.835
+ $Y=1.84 $X2=5.97 $Y2=2.8
r91 1 37 600 $w=1.7e-07 $l=1.02995e-06 $layer=licon1_PDIFF $count=1 $X=4.75
+ $Y=1.84 $X2=4.895 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR2_4%A_27_74# 1 2 3 12 14 15 16 17 20
c40 16 0 7.39126e-20 $X=1.21 $Y=0.6
c41 14 0 1.04341e-19 $X=1.045 $Y=1.065
r42 18 23 3.97509 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.475
+ $X2=1.21 $Y2=0.475
r43 18 20 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=1.375 $Y=0.475
+ $X2=2.14 $Y2=0.475
r44 16 23 3.01144 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=1.21 $Y=0.6 $X2=1.21
+ $Y2=0.475
r45 16 17 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.21 $Y=0.6 $X2=1.21
+ $Y2=0.98
r46 14 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.045 $Y=1.065
+ $X2=1.21 $Y2=0.98
r47 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.045 $Y=1.065
+ $X2=0.365 $Y2=1.065
r48 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.98
+ $X2=0.365 $Y2=1.065
r49 10 12 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=0.24 $Y=0.98
+ $X2=0.24 $Y2=0.515
r50 3 20 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2 $Y=0.37
+ $X2=2.14 $Y2=0.515
r51 2 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.37 $X2=1.21 $Y2=0.515
r52 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR2_4%VGND 1 2 3 4 5 18 22 26 30 34 37 38 40 41 43
+ 44 45 47 65 71 72 75 78
r117 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r118 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r119 72 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r120 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r121 69 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.495 $Y=0 $X2=8.33
+ $Y2=0
r122 69 71 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=8.495 $Y=0
+ $X2=8.88 $Y2=0
r123 68 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r124 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r125 65 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.165 $Y=0 $X2=8.33
+ $Y2=0
r126 65 67 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=8.165 $Y=0 $X2=7.92
+ $Y2=0
r127 64 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r128 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r129 61 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r130 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r131 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r132 57 58 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r133 55 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r134 54 57 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=5.04
+ $Y2=0
r135 54 55 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.2 $Y=0
+ $X2=1.2 $Y2=0
r136 52 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r137 52 54 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r138 50 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r139 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r140 47 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r141 47 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r142 45 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r143 45 55 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=1.2
+ $Y2=0
r144 43 63 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=7.11 $Y=0 $X2=6.96
+ $Y2=0
r145 43 44 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=7.11 $Y=0 $X2=7.292
+ $Y2=0
r146 42 67 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=7.475 $Y=0
+ $X2=7.92 $Y2=0
r147 42 44 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=7.475 $Y=0
+ $X2=7.292 $Y2=0
r148 40 60 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=6.09 $Y=0 $X2=6 $Y2=0
r149 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.09 $Y=0 $X2=6.255
+ $Y2=0
r150 39 63 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=6.42 $Y=0 $X2=6.96
+ $Y2=0
r151 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.42 $Y=0 $X2=6.255
+ $Y2=0
r152 37 57 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=5.07 $Y=0 $X2=5.04
+ $Y2=0
r153 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.07 $Y=0 $X2=5.235
+ $Y2=0
r154 36 60 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.4 $Y=0 $X2=6 $Y2=0
r155 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.4 $Y=0 $X2=5.235
+ $Y2=0
r156 32 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.33 $Y=0.085
+ $X2=8.33 $Y2=0
r157 32 34 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=8.33 $Y=0.085
+ $X2=8.33 $Y2=0.335
r158 28 44 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=7.292 $Y=0.085
+ $X2=7.292 $Y2=0
r159 28 30 7.89345 $w=3.63e-07 $l=2.5e-07 $layer=LI1_cond $X=7.292 $Y=0.085
+ $X2=7.292 $Y2=0.335
r160 24 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.255 $Y=0.085
+ $X2=6.255 $Y2=0
r161 24 26 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=6.255 $Y=0.085
+ $X2=6.255 $Y2=0.335
r162 20 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.235 $Y=0.085
+ $X2=5.235 $Y2=0
r163 20 22 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=5.235 $Y=0.085
+ $X2=5.235 $Y2=0.335
r164 16 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r165 16 18 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.58
r166 5 34 182 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_NDIFF $count=1 $X=8.11
+ $Y=0.37 $X2=8.33 $Y2=0.335
r167 4 30 182 $w=1.7e-07 $l=2.51893e-07 $layer=licon1_NDIFF $count=1 $X=7.055
+ $Y=0.37 $X2=7.29 $Y2=0.335
r168 3 26 182 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_NDIFF $count=1 $X=6.035
+ $Y=0.37 $X2=6.255 $Y2=0.335
r169 2 22 182 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_NDIFF $count=1 $X=5.015
+ $Y=0.37 $X2=5.235 $Y2=0.335
r170 1 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR2_4%A_511_74# 1 2 3 4 5 6 7 24 26 27 30 32 37 38
+ 39 40 42 44 46 48 53 58 63
c121 44 0 3.01105e-20 $X=8.675 $Y=0.755
c122 42 0 6.02202e-20 $X=7.655 $Y=0.755
c123 40 0 6.0221e-20 $X=6.6 $Y=0.755
c124 38 0 3.01101e-20 $X=5.58 $Y=0.755
r125 63 65 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=8.84 $Y=0.515
+ $X2=8.84 $Y2=0.755
r126 58 60 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=7.82 $Y=0.595
+ $X2=7.82 $Y2=0.755
r127 53 55 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=6.765 $Y=0.595
+ $X2=6.765 $Y2=0.755
r128 48 50 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=5.745 $Y=0.595
+ $X2=5.745 $Y2=0.755
r129 45 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.985 $Y=0.755
+ $X2=7.82 $Y2=0.755
r130 44 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.675 $Y=0.755
+ $X2=8.84 $Y2=0.755
r131 44 45 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.675 $Y=0.755
+ $X2=7.985 $Y2=0.755
r132 43 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.93 $Y=0.755
+ $X2=6.765 $Y2=0.755
r133 42 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.655 $Y=0.755
+ $X2=7.82 $Y2=0.755
r134 42 43 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=7.655 $Y=0.755
+ $X2=6.93 $Y2=0.755
r135 41 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.91 $Y=0.755
+ $X2=5.745 $Y2=0.755
r136 40 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.6 $Y=0.755
+ $X2=6.765 $Y2=0.755
r137 40 41 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.6 $Y=0.755
+ $X2=5.91 $Y2=0.755
r138 38 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.58 $Y=0.755
+ $X2=5.745 $Y2=0.755
r139 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.58 $Y=0.755
+ $X2=4.89 $Y2=0.755
r140 35 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.725 $Y=0.67
+ $X2=4.89 $Y2=0.755
r141 35 37 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=4.725 $Y=0.67
+ $X2=4.725 $Y2=0.595
r142 34 37 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.725 $Y=0.425
+ $X2=4.725 $Y2=0.595
r143 33 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.865 $Y=0.34
+ $X2=3.7 $Y2=0.34
r144 32 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.56 $Y=0.34
+ $X2=4.725 $Y2=0.425
r145 32 33 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.56 $Y=0.34
+ $X2=3.865 $Y2=0.34
r146 28 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.425 $X2=3.7
+ $Y2=0.34
r147 28 30 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.7 $Y=0.425
+ $X2=3.7 $Y2=0.595
r148 26 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.535 $Y=0.34
+ $X2=3.7 $Y2=0.34
r149 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.535 $Y=0.34
+ $X2=2.865 $Y2=0.34
r150 22 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.7 $Y=0.425
+ $X2=2.865 $Y2=0.34
r151 22 24 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.7 $Y=0.425
+ $X2=2.7 $Y2=0.595
r152 7 63 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.7
+ $Y=0.37 $X2=8.84 $Y2=0.515
r153 6 58 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=7.68
+ $Y=0.37 $X2=7.82 $Y2=0.595
r154 5 53 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=6.625
+ $Y=0.37 $X2=6.765 $Y2=0.595
r155 4 48 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=5.605
+ $Y=0.37 $X2=5.745 $Y2=0.595
r156 3 37 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=4.515
+ $Y=0.37 $X2=4.725 $Y2=0.595
r157 2 30 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=3.49
+ $Y=0.37 $X2=3.7 $Y2=0.595
r158 1 24 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=2.555
+ $Y=0.37 $X2=2.7 $Y2=0.595
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and4_4 A B C D VGND VNB VPB VPWR X
X0 a_119_392# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X1 VPWR A a_119_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X2 a_463_119# C a_32_119# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 VPWR a_119_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X4 a_463_119# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 a_32_119# C a_463_119# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 VGND a_119_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VPWR C a_119_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X8 VPWR D a_119_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X9 X a_119_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 X a_119_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_32_119# B a_119_119# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X12 a_119_392# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X13 VGND a_119_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 X a_119_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 a_119_392# C VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X16 X a_119_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X17 a_119_119# A a_119_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X18 a_119_392# D VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X19 VGND D a_463_119# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X20 VPWR a_119_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X21 a_119_119# B a_32_119# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X22 VPWR B a_119_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X23 a_119_392# A a_119_119# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_ms__mux2i_1 A0 A1 S VGND VNB VPB VPWR Y
*.PININFO A0:I A1:I S:I VGND:I VNB:I VPB:I VPWR:I Y:O
MMNA00 Y A0 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA01 smdNA0 Sb VNB nfet_01v8_lvt m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA10 Y A1 VNB nfet_01v8_lvt m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMNA11 sndNA1 S VNB nfet_01v8_lvt m=1 w=0.74 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 Sb S VNB nfet_01v8_lvt m=1 w=0.55 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA00 VPWR S VPB pfet_01v8 m=1 w=1.12 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMPA01 sndPS A0 VPB pfet_01v8 m=1 w=1.12 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA10 VPWR Sb VPB pfet_01v8 m=1 w=1.12 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMPA11 sndPSb A1 VPB pfet_01v8 m=1 w=1.12 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 Sb S VPB pfet_01v8 m=1 w=0.84 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_ms__mux2i_1

* NGSPICE file created from sky130_fd_sc_ms__xnor3_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__xnor3_2 A B C VGND VNB VPB VPWR X
M1000 a_335_373# B a_83_247# VPB pshort w=840000u l=180000u
+  ad=5.572e+11p pd=4.77e+06u as=7.096e+11p ps=5.58e+06u
M1001 a_83_247# a_397_21# a_329_81# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=5.174e+11p ps=4.63e+06u
M1002 a_83_247# a_397_21# a_335_373# VNB nlowvt w=640000u l=150000u
+  ad=5.925e+11p pd=4.86e+06u as=4.512e+11p ps=3.97e+06u
M1003 a_335_373# B a_27_373# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=3.886e+11p ps=3.85e+06u
M1004 a_27_373# a_397_21# a_329_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=4.22e+11p ps=4.25e+06u
M1005 a_1057_74# a_1027_48# a_335_373# VPB pshort w=840000u l=180000u
+  ad=4.0245e+11p pd=2.81e+06u as=0p ps=0u
M1006 X a_1057_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.5438e+12p ps=1.187e+07u
M1007 a_329_81# C a_1057_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_1057_74# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_1057_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=1.54235e+12p ps=1.041e+07u
M1010 a_83_247# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_373# a_397_21# a_335_373# VPB pshort w=640000u l=180000u
+  ad=4.656e+11p pd=4.42e+06u as=0p ps=0u
M1012 VGND a_83_247# a_27_373# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND C a_1027_48# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1014 a_329_81# B a_27_373# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_83_247# a_27_373# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND B a_397_21# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1017 VGND a_1057_74# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_329_81# B a_83_247# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_335_373# C a_1057_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.24e+11p ps=1.98e+06u
M1020 VPWR C a_1027_48# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.76e+11p ps=1.83e+06u
M1021 VPWR B a_397_21# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.08e+11p ps=2.79e+06u
M1022 a_83_247# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1057_74# a_1027_48# a_329_81# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


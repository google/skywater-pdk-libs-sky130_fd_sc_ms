* File: sky130_fd_sc_ms__or2_2.spice
* Created: Fri Aug 28 18:06:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__or2_2.pex.spice"
.subckt sky130_fd_sc_ms__or2_2  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1003 N_A_27_368#_M1003_d N_B_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1792 PD=0.92 PS=1.84 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1005 N_VGND_M1005_d N_A_M1005_g N_A_27_368#_M1003_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.118354 AS=0.0896 PD=1.01565 PS=0.92 NRD=14.052 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1005_d N_A_27_368#_M1001_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.136846 AS=0.1036 PD=1.17435 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_A_27_368#_M1006_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2479 AS=0.1036 PD=2.15 PS=1.02 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75001.4
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1004 A_117_368# N_B_M1004_g N_A_27_368#_M1004_s VPB PSHORT L=0.18 W=1 AD=0.105
+ AS=0.27 PD=1.21 PS=2.54 NRD=9.8303 NRS=0 M=1 R=5.55556 SA=90000.2 SB=90001.6
+ A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g A_117_368# VPB PSHORT L=0.18 W=1 AD=0.18566
+ AS=0.105 PD=1.39623 PS=1.21 NRD=17.7103 NRS=9.8303 M=1 R=5.55556 SA=90000.6
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1002 N_X_M1002_d N_A_27_368#_M1002_g N_VPWR_M1000_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1624 AS=0.20794 PD=1.41 PS=1.56377 NRD=0.8668 NRS=0 M=1 R=6.22222
+ SA=90001 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1007 N_X_M1002_d N_A_27_368#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1624 AS=0.3136 PD=1.41 PS=2.8 NRD=0.8668 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.1708 P=9.28
*
.include "sky130_fd_sc_ms__or2_2.pxi.spice"
*
.ends
*
*

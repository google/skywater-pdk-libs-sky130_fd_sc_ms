* File: sky130_fd_sc_ms__nor3_4.spice
* Created: Fri Aug 28 17:48:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nor3_4.pex.spice"
.subckt sky130_fd_sc_ms__nor3_4  VNB VPB A B C VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_M1004_g N_Y_M1004_s VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.1073 PD=2.05 PS=1.03 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2 SB=75002.9
+ A=0.111 P=1.78 MULT=1
MM1016 N_VGND_M1016_d N_A_M1016_g N_Y_M1004_s VNB NLOWVT L=0.15 W=0.74 AD=0.1517
+ AS=0.1073 PD=1.15 PS=1.03 NRD=9.72 NRS=1.62 M=1 R=4.93333 SA=75000.6
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1006 N_Y_M1006_d N_B_M1006_g N_VGND_M1016_d VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.1517 PD=1.02 PS=1.15 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.2 SB=75001.9
+ A=0.111 P=1.78 MULT=1
MM1013 N_Y_M1006_d N_B_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.6 SB=75001.5
+ A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_C_M1002_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.2 SB=75000.9
+ A=0.111 P=1.78 MULT=1
MM1007 N_Y_M1002_d N_C_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.40425 PD=1.02 PS=2.58 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.6 SB=75000.5
+ A=0.111 P=1.78 MULT=1
MM1008 N_A_27_368#_M1008_d N_A_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.308 AS=0.1512 PD=2.79 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90005.9 A=0.2016 P=2.6 MULT=1
MM1009 N_A_27_368#_M1009_d N_A_M1009_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90005.5 A=0.2016 P=2.6 MULT=1
MM1003 N_A_27_368#_M1009_d N_B_M1003_g N_A_298_368#_M1003_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2545 PD=1.39 PS=1.665 NRD=0 NRS=14.0658 M=1 R=6.22222
+ SA=90001.1 SB=90005 A=0.2016 P=2.6 MULT=1
MM1000 N_Y_M1000_d N_C_M1000_g N_A_298_368#_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.24465 AS=0.2545 PD=1.61 PS=1.665 NRD=13.1793 NRS=13.1793 M=1 R=6.22222
+ SA=90001.7 SB=90004.4 A=0.2016 P=2.6 MULT=1
MM1001 N_Y_M1000_d N_C_M1001_g N_A_298_368#_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.24465 AS=0.2576 PD=1.61 PS=1.67 NRD=13.1793 NRS=14.0658 M=1 R=6.22222
+ SA=90002.3 SB=90003.8 A=0.2016 P=2.6 MULT=1
MM1015 N_Y_M1015_d N_C_M1015_g N_A_298_368#_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.24465 AS=0.2576 PD=1.61 PS=1.67 NRD=13.1793 NRS=14.0658 M=1 R=6.22222
+ SA=90002.9 SB=90003.2 A=0.2016 P=2.6 MULT=1
MM1017 N_Y_M1015_d N_C_M1017_g N_A_298_368#_M1017_s VPB PSHORT L=0.18 W=1.12
+ AD=0.24465 AS=0.2576 PD=1.61 PS=1.67 NRD=13.1793 NRS=14.0658 M=1 R=6.22222
+ SA=90003.5 SB=90002.6 A=0.2016 P=2.6 MULT=1
MM1005 N_A_27_368#_M1005_d N_B_M1005_g N_A_298_368#_M1017_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2576 PD=1.39 PS=1.67 NRD=0 NRS=14.0658 M=1 R=6.22222
+ SA=90004.1 SB=90002 A=0.2016 P=2.6 MULT=1
MM1010 N_A_27_368#_M1005_d N_B_M1010_g N_A_298_368#_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90004.6 SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1011 N_A_27_368#_M1011_d N_B_M1011_g N_A_298_368#_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90005
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1012 N_A_27_368#_M1011_d N_A_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90005.5
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1014 N_A_27_368#_M1014_d N_A_M1014_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3024 AS=0.1512 PD=2.78 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90005.9
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX18_noxref VNB VPB NWDIODE A=13.3495 P=18.06
c_105 VPB 0 3.61225e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__nor3_4.pxi.spice"
*
.ends
*
*

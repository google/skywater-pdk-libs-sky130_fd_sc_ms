* File: sky130_fd_sc_ms__xor2_4.pex.spice
* Created: Wed Sep  2 12:34:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__XOR2_4%A 3 7 11 15 19 23 27 31 35 39 41 45 49 52 53
+ 55 57 58 60 63 66 67 68 70 71 72 73 74 75 76 81 88 96 97
c226 88 0 1.58295e-19 $X=1.05 $Y=1.585
c227 68 0 1.24044e-19 $X=3.04 $Y=1.105
c228 60 0 4.48662e-20 $X=0.945 $Y=1.585
c229 53 0 1.31802e-19 $X=6.345 $Y=1.485
c230 41 0 1.05217e-19 $X=6.255 $Y=1.485
c231 27 0 9.66338e-20 $X=5.315 $Y=2.4
c232 19 0 9.06279e-20 $X=4.725 $Y=2.4
c233 7 0 1.34713e-19 $X=0.725 $Y=0.86
r234 95 96 17.8155 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.765 $Y=1.515
+ $X2=5.855 $Y2=1.515
r235 93 95 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=5.45 $Y=1.515
+ $X2=5.765 $Y2=1.515
r236 93 94 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.45
+ $Y=1.515 $X2=5.45 $Y2=1.515
r237 91 93 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=5.335 $Y=1.515
+ $X2=5.45 $Y2=1.515
r238 90 91 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=5.315 $Y=1.515
+ $X2=5.335 $Y2=1.515
r239 85 86 27.2977 $w=3.09e-07 $l=1.75e-07 $layer=POLY_cond $X=0.55 $Y=1.585
+ $X2=0.725 $Y2=1.585
r240 84 94 9.21954 $w=4.23e-07 $l=3.4e-07 $layer=LI1_cond $X=5.11 $Y=1.562
+ $X2=5.45 $Y2=1.562
r241 83 84 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.11
+ $Y=1.515 $X2=5.11 $Y2=1.515
r242 81 90 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.225 $Y=1.515
+ $X2=5.315 $Y2=1.515
r243 81 83 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=5.225 $Y=1.515
+ $X2=5.11 $Y2=1.515
r244 76 94 1.89814 $w=4.23e-07 $l=7e-08 $layer=LI1_cond $X=5.52 $Y=1.562
+ $X2=5.45 $Y2=1.562
r245 75 84 1.89814 $w=4.23e-07 $l=7e-08 $layer=LI1_cond $X=5.04 $Y=1.562
+ $X2=5.11 $Y2=1.562
r246 74 75 13.0158 $w=4.23e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.562
+ $X2=5.04 $Y2=1.562
r247 74 97 4.60977 $w=4.23e-07 $l=1.7e-07 $layer=LI1_cond $X=4.56 $Y=1.562
+ $X2=4.39 $Y2=1.562
r248 73 97 9.38859 $w=4.25e-07 $l=3.1e-07 $layer=LI1_cond $X=4.08 $Y=1.562
+ $X2=4.39 $Y2=1.562
r249 71 72 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=1.275 $Y=0.675
+ $X2=1.445 $Y2=0.675
r250 70 73 8.18076 $w=3.43e-07 $l=3.18842e-07 $layer=LI1_cond $X=3.85 $Y=1.35
+ $X2=4.08 $Y2=1.562
r251 69 70 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.85 $Y=1.19
+ $X2=3.85 $Y2=1.35
r252 67 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.765 $Y=1.105
+ $X2=3.85 $Y2=1.19
r253 67 68 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.765 $Y=1.105
+ $X2=3.04 $Y2=1.105
r254 66 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.955 $Y=1.02
+ $X2=3.04 $Y2=1.105
r255 65 66 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.955 $Y=0.77
+ $X2=2.955 $Y2=1.02
r256 63 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.87 $Y=0.685
+ $X2=2.955 $Y2=0.77
r257 63 72 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=2.87 $Y=0.685
+ $X2=1.445 $Y2=0.685
r258 61 88 16.3786 $w=3.09e-07 $l=1.05e-07 $layer=POLY_cond $X=0.945 $Y=1.585
+ $X2=1.05 $Y2=1.585
r259 61 86 34.3172 $w=3.09e-07 $l=2.2e-07 $layer=POLY_cond $X=0.945 $Y=1.585
+ $X2=0.725 $Y2=1.585
r260 60 61 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.945
+ $Y=1.585 $X2=0.945 $Y2=1.585
r261 58 60 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=0.685 $Y=1.585
+ $X2=0.945 $Y2=1.585
r262 57 71 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.685 $Y=0.665
+ $X2=1.275 $Y2=0.665
r263 55 58 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.6 $Y=1.42
+ $X2=0.685 $Y2=1.585
r264 54 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.6 $Y=0.75
+ $X2=0.685 $Y2=0.665
r265 54 55 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.6 $Y=0.75 $X2=0.6
+ $Y2=1.42
r266 51 83 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=4.82 $Y=1.515
+ $X2=5.11 $Y2=1.515
r267 51 52 3.90195 $w=3.3e-07 $l=1.08e-07 $layer=POLY_cond $X=4.82 $Y=1.515
+ $X2=4.712 $Y2=1.515
r268 47 53 30.0832 $w=1.65e-07 $l=1.39911e-07 $layer=POLY_cond $X=6.355 $Y=1.35
+ $X2=6.345 $Y2=1.485
r269 47 49 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.355 $Y=1.35
+ $X2=6.355 $Y2=0.74
r270 43 53 30.0832 $w=1.65e-07 $l=1.35e-07 $layer=POLY_cond $X=6.345 $Y=1.62
+ $X2=6.345 $Y2=1.485
r271 43 45 303.194 $w=1.8e-07 $l=7.8e-07 $layer=POLY_cond $X=6.345 $Y=1.62
+ $X2=6.345 $Y2=2.4
r272 41 53 1.40033 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=6.255 $Y=1.485
+ $X2=6.345 $Y2=1.485
r273 41 96 88.8695 $w=2.7e-07 $l=4e-07 $layer=POLY_cond $X=6.255 $Y=1.485
+ $X2=5.855 $Y2=1.485
r274 37 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.765 $Y=1.35
+ $X2=5.765 $Y2=1.515
r275 37 39 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.765 $Y=1.35
+ $X2=5.765 $Y2=0.74
r276 33 95 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.765 $Y=1.68
+ $X2=5.765 $Y2=1.515
r277 33 35 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.765 $Y=1.68
+ $X2=5.765 $Y2=2.4
r278 29 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.335 $Y=1.35
+ $X2=5.335 $Y2=1.515
r279 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.335 $Y=1.35
+ $X2=5.335 $Y2=0.74
r280 25 90 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.315 $Y=1.68
+ $X2=5.315 $Y2=1.515
r281 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.315 $Y=1.68
+ $X2=5.315 $Y2=2.4
r282 21 52 34.7346 $w=1.65e-07 $l=1.80748e-07 $layer=POLY_cond $X=4.745 $Y=1.35
+ $X2=4.712 $Y2=1.515
r283 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.745 $Y=1.35
+ $X2=4.745 $Y2=0.74
r284 17 52 34.7346 $w=1.65e-07 $l=1.71377e-07 $layer=POLY_cond $X=4.725 $Y=1.68
+ $X2=4.712 $Y2=1.515
r285 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.725 $Y=1.68
+ $X2=4.725 $Y2=2.4
r286 13 88 16.3786 $w=3.09e-07 $l=2.11069e-07 $layer=POLY_cond $X=1.155 $Y=1.42
+ $X2=1.05 $Y2=1.585
r287 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.155 $Y=1.42
+ $X2=1.155 $Y2=0.86
r288 9 88 15.404 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.05 $Y=1.75
+ $X2=1.05 $Y2=1.585
r289 9 11 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=1.05 $Y=1.75
+ $X2=1.05 $Y2=2.46
r290 5 86 19.6649 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.725 $Y=1.42
+ $X2=0.725 $Y2=1.585
r291 5 7 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.725 $Y=1.42
+ $X2=0.725 $Y2=0.86
r292 1 85 15.404 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.55 $Y=1.75
+ $X2=0.55 $Y2=1.585
r293 1 3 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=0.55 $Y=1.75 $X2=0.55
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__XOR2_4%B 1 3 6 8 10 13 15 17 22 23 24 28 31 35 39 43
+ 45 47 52 53 55 56 57 59 60 61 65 66 67 68 69 90 94
c199 59 0 9.66338e-20 $X=5.89 $Y=1.78
c200 17 0 1.47912e-19 $X=6.795 $Y=2.4
c201 15 0 1.60229e-19 $X=6.795 $Y=1.275
c202 13 0 1.24044e-19 $X=2.285 $Y=0.86
c203 6 0 1.87977e-19 $X=1.745 $Y=0.86
r204 92 94 0.670025 $w=4.28e-07 $l=2.5e-08 $layer=LI1_cond $X=5.975 $Y=1.565
+ $X2=6 $Y2=1.565
r205 89 90 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8
+ $Y=1.515 $X2=8 $Y2=1.515
r206 84 86 51.6429 $w=3.5e-07 $l=3.75e-07 $layer=POLY_cond $X=7.32 $Y=1.432
+ $X2=7.695 $Y2=1.432
r207 84 85 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.32
+ $Y=1.515 $X2=7.32 $Y2=1.515
r208 82 84 10.3286 $w=3.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.245 $Y=1.432
+ $X2=7.32 $Y2=1.432
r209 81 82 4.13143 $w=3.5e-07 $l=3e-08 $layer=POLY_cond $X=7.215 $Y=1.432
+ $X2=7.245 $Y2=1.432
r210 76 77 32.8941 $w=3.59e-07 $l=2.45e-07 $layer=POLY_cond $X=1.5 $Y=1.685
+ $X2=1.745 $Y2=1.685
r211 69 90 2.14408 $w=4.28e-07 $l=8e-08 $layer=LI1_cond $X=7.92 $Y=1.565 $X2=8
+ $Y2=1.565
r212 68 69 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.92 $Y2=1.565
r213 68 85 3.21612 $w=4.28e-07 $l=1.2e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.32 $Y2=1.565
r214 67 85 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.32 $Y2=1.565
r215 66 67 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.96 $Y2=1.565
r216 65 92 2.44569 $w=4.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.89 $Y=1.565
+ $X2=5.975 $Y2=1.565
r217 65 66 12.0604 $w=4.28e-07 $l=4.5e-07 $layer=LI1_cond $X=6.03 $Y=1.565
+ $X2=6.48 $Y2=1.565
r218 65 94 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=6.03 $Y=1.565 $X2=6
+ $Y2=1.565
r219 61 63 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.57 $Y=1.935
+ $X2=3.57 $Y2=2.03
r220 59 65 6.18617 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=5.89 $Y=1.78
+ $X2=5.89 $Y2=1.565
r221 59 60 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.89 $Y=1.78
+ $X2=5.89 $Y2=1.945
r222 58 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.655 $Y=2.03
+ $X2=3.57 $Y2=2.03
r223 57 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.805 $Y=2.03
+ $X2=5.89 $Y2=1.945
r224 57 58 140.267 $w=1.68e-07 $l=2.15e-06 $layer=LI1_cond $X=5.805 $Y=2.03
+ $X2=3.655 $Y2=2.03
r225 55 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.485 $Y=1.935
+ $X2=3.57 $Y2=1.935
r226 55 56 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=3.485 $Y=1.935
+ $X2=2.36 $Y2=1.935
r227 53 80 12.0836 $w=3.59e-07 $l=9e-08 $layer=POLY_cond $X=2.195 $Y=1.685
+ $X2=2.285 $Y2=1.685
r228 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.195
+ $Y=1.635 $X2=2.195 $Y2=1.635
r229 50 56 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.195 $Y=1.85
+ $X2=2.36 $Y2=1.935
r230 50 52 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.195 $Y=1.85
+ $X2=2.195 $Y2=1.635
r231 45 89 19.9686 $w=3.5e-07 $l=1.45e-07 $layer=POLY_cond $X=8.145 $Y=1.432
+ $X2=8 $Y2=1.432
r232 45 47 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.145 $Y=1.35
+ $X2=8.145 $Y2=0.74
r233 41 45 18.307 $w=1.8e-07 $l=2.48e-07 $layer=POLY_cond $X=8.145 $Y=1.68
+ $X2=8.145 $Y2=1.432
r234 41 43 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.145 $Y=1.68
+ $X2=8.145 $Y2=2.4
r235 37 89 39.2486 $w=3.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.715 $Y=1.432
+ $X2=8 $Y2=1.432
r236 37 86 2.75429 $w=3.5e-07 $l=2e-08 $layer=POLY_cond $X=7.715 $Y=1.432
+ $X2=7.695 $Y2=1.432
r237 37 39 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.715 $Y=1.35
+ $X2=7.715 $Y2=0.74
r238 33 86 18.307 $w=1.8e-07 $l=2.48e-07 $layer=POLY_cond $X=7.695 $Y=1.68
+ $X2=7.695 $Y2=1.432
r239 33 35 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.695 $Y=1.68
+ $X2=7.695 $Y2=2.4
r240 29 82 18.307 $w=1.8e-07 $l=2.48e-07 $layer=POLY_cond $X=7.245 $Y=1.68
+ $X2=7.245 $Y2=1.432
r241 29 31 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.245 $Y=1.68
+ $X2=7.245 $Y2=2.4
r242 26 81 22.6286 $w=1.5e-07 $l=2.47e-07 $layer=POLY_cond $X=7.215 $Y=1.185
+ $X2=7.215 $Y2=1.432
r243 26 28 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=7.215 $Y=1.185
+ $X2=7.215 $Y2=0.74
r244 25 28 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=7.215 $Y=0.295
+ $X2=7.215 $Y2=0.74
r245 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.14 $Y=0.22
+ $X2=7.215 $Y2=0.295
r246 23 24 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=7.14 $Y=0.22
+ $X2=6.86 $Y2=0.22
r247 22 49 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=6.785 $Y=0.74
+ $X2=6.785 $Y2=1.185
r248 19 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.785 $Y=0.295
+ $X2=6.86 $Y2=0.22
r249 19 22 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=6.785 $Y=0.295
+ $X2=6.785 $Y2=0.74
r250 15 49 36.5962 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.795 $Y=1.275
+ $X2=6.795 $Y2=1.185
r251 15 17 437.298 $w=1.8e-07 $l=1.125e-06 $layer=POLY_cond $X=6.795 $Y=1.275
+ $X2=6.795 $Y2=2.4
r252 11 80 23.2387 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=2.285 $Y=1.47
+ $X2=2.285 $Y2=1.685
r253 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.285 $Y=1.47
+ $X2=2.285 $Y2=0.86
r254 8 53 32.8941 $w=3.59e-07 $l=2.45e-07 $layer=POLY_cond $X=1.95 $Y=1.685
+ $X2=2.195 $Y2=1.685
r255 8 77 27.5237 $w=3.59e-07 $l=2.05e-07 $layer=POLY_cond $X=1.95 $Y=1.685
+ $X2=1.745 $Y2=1.685
r256 8 10 164.683 $w=1.8e-07 $l=6.15e-07 $layer=POLY_cond $X=1.95 $Y=1.845
+ $X2=1.95 $Y2=2.46
r257 4 77 23.2387 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.745 $Y=1.47
+ $X2=1.745 $Y2=1.685
r258 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.745 $Y=1.47
+ $X2=1.745 $Y2=0.86
r259 1 76 18.9031 $w=1.8e-07 $l=2.15e-07 $layer=POLY_cond $X=1.5 $Y=1.9 $X2=1.5
+ $Y2=1.685
r260 1 3 149.956 $w=1.8e-07 $l=5.6e-07 $layer=POLY_cond $X=1.5 $Y=1.9 $X2=1.5
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__XOR2_4%A_160_98# 1 2 3 10 12 15 19 21 23 26 28 29 32
+ 34 38 40 45 46 51 57 58
c130 57 0 2.77823e-19 $X=1.105 $Y=1.085
r131 61 62 73.277 $w=2.96e-07 $l=4.5e-07 $layer=POLY_cond $X=2.925 $Y=1.515
+ $X2=3.375 $Y2=1.515
r132 60 61 8.14189 $w=2.96e-07 $l=5e-08 $layer=POLY_cond $X=2.875 $Y=1.515
+ $X2=2.925 $Y2=1.515
r133 55 57 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.94 $Y=1.085
+ $X2=1.105 $Y2=1.085
r134 52 64 26.0541 $w=2.96e-07 $l=1.6e-07 $layer=POLY_cond $X=3.43 $Y=1.515
+ $X2=3.59 $Y2=1.515
r135 52 62 8.95608 $w=2.96e-07 $l=5.5e-08 $layer=POLY_cond $X=3.43 $Y=1.515
+ $X2=3.375 $Y2=1.515
r136 51 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.43
+ $Y=1.515 $X2=3.43 $Y2=1.515
r137 49 60 20.3547 $w=2.96e-07 $l=1.25e-07 $layer=POLY_cond $X=2.75 $Y=1.515
+ $X2=2.875 $Y2=1.515
r138 48 51 24.4894 $w=3.18e-07 $l=6.8e-07 $layer=LI1_cond $X=2.75 $Y=1.52
+ $X2=3.43 $Y2=1.52
r139 48 49 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.75
+ $Y=1.515 $X2=2.75 $Y2=1.515
r140 46 48 1.80069 $w=3.18e-07 $l=5e-08 $layer=LI1_cond $X=2.7 $Y=1.52 $X2=2.75
+ $Y2=1.52
r141 45 46 7.68211 $w=3.2e-07 $l=1.9799e-07 $layer=LI1_cond $X=2.615 $Y=1.36
+ $X2=2.7 $Y2=1.52
r142 44 45 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.615 $Y=1.19
+ $X2=2.615 $Y2=1.36
r143 41 58 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.81 $Y=1.065
+ $X2=1.685 $Y2=1.065
r144 41 43 9.45003 $w=2.48e-07 $l=2.05e-07 $layer=LI1_cond $X=1.81 $Y=1.065
+ $X2=2.015 $Y2=1.065
r145 40 44 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.53 $Y=1.065
+ $X2=2.615 $Y2=1.19
r146 40 43 23.7403 $w=2.48e-07 $l=5.15e-07 $layer=LI1_cond $X=2.53 $Y=1.065
+ $X2=2.015 $Y2=1.065
r147 36 58 1.34256 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.685 $Y=1.19
+ $X2=1.685 $Y2=1.065
r148 36 38 42.1794 $w=2.48e-07 $l=9.15e-07 $layer=LI1_cond $X=1.685 $Y=1.19
+ $X2=1.685 $Y2=2.105
r149 34 58 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.56 $Y=1.065
+ $X2=1.685 $Y2=1.065
r150 34 57 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=1.56 $Y=1.065
+ $X2=1.105 $Y2=1.065
r151 30 32 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.275 $Y=1.68
+ $X2=4.275 $Y2=2.4
r152 28 30 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.185 $Y=1.605
+ $X2=4.275 $Y2=1.68
r153 28 29 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.185 $Y=1.605
+ $X2=3.915 $Y2=1.605
r154 24 29 26.359 $w=2.96e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.825 $Y=1.68
+ $X2=3.915 $Y2=1.605
r155 24 64 38.2669 $w=2.96e-07 $l=3.06594e-07 $layer=POLY_cond $X=3.825 $Y=1.68
+ $X2=3.59 $Y2=1.515
r156 24 26 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.825 $Y=1.68
+ $X2=3.825 $Y2=2.4
r157 21 64 18.6531 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.59 $Y=1.35
+ $X2=3.59 $Y2=1.515
r158 21 23 157.453 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=3.59 $Y=1.35
+ $X2=3.59 $Y2=0.86
r159 17 62 14.4094 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.375 $Y=1.68
+ $X2=3.375 $Y2=1.515
r160 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.375 $Y=1.68
+ $X2=3.375 $Y2=2.4
r161 13 61 14.4094 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.925 $Y=1.68
+ $X2=2.925 $Y2=1.515
r162 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.925 $Y=1.68
+ $X2=2.925 $Y2=2.4
r163 10 60 18.6531 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.875 $Y=1.35
+ $X2=2.875 $Y2=1.515
r164 10 12 157.453 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=2.875 $Y=1.35
+ $X2=2.875 $Y2=0.86
r165 3 38 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.59
+ $Y=1.96 $X2=1.725 $Y2=2.105
r166 2 43 182 $w=1.7e-07 $l=6.2494e-07 $layer=licon1_NDIFF $count=1 $X=1.82
+ $Y=0.49 $X2=2.015 $Y2=1.025
r167 1 55 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=0.8
+ $Y=0.49 $X2=0.94 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_MS__XOR2_4%A_36_392# 1 2 3 12 16 17 21 24 25 28
c43 17 0 1.58295e-19 $X=0.49 $Y=2.005
r44 26 28 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=2.175 $Y=2.905
+ $X2=2.175 $Y2=2.355
r45 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.01 $Y=2.99
+ $X2=2.175 $Y2=2.905
r46 24 25 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.01 $Y=2.99
+ $X2=1.36 $Y2=2.99
r47 21 23 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=1.235 $Y=2.105
+ $X2=1.235 $Y2=2.815
r48 19 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.235 $Y=2.905
+ $X2=1.36 $Y2=2.99
r49 19 23 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.235 $Y=2.905
+ $X2=1.235 $Y2=2.815
r50 18 21 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=1.235 $Y=2.09
+ $X2=1.235 $Y2=2.105
r51 16 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.11 $Y=2.005
+ $X2=1.235 $Y2=2.09
r52 16 17 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.11 $Y=2.005
+ $X2=0.49 $Y2=2.005
r53 12 14 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.325 $Y=2.105
+ $X2=0.325 $Y2=2.815
r54 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.325 $Y=2.09
+ $X2=0.49 $Y2=2.005
r55 10 12 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.325 $Y=2.09
+ $X2=0.325 $Y2=2.105
r56 3 28 300 $w=1.7e-07 $l=4.57548e-07 $layer=licon1_PDIFF $count=2 $X=2.04
+ $Y=1.96 $X2=2.175 $Y2=2.355
r57 2 23 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.14
+ $Y=1.96 $X2=1.275 $Y2=2.815
r58 2 21 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.14
+ $Y=1.96 $X2=1.275 $Y2=2.105
r59 1 14 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.18
+ $Y=1.96 $X2=0.325 $Y2=2.815
r60 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.18
+ $Y=1.96 $X2=0.325 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_MS__XOR2_4%VPWR 1 2 3 4 5 20 24 28 30 32 40 45 50 57 58
+ 61 64 71 78 81
r117 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r118 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r119 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r120 71 74 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=6.055 $Y=3.05
+ $X2=6.055 $Y2=3.33
r121 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r122 64 67 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=5.02 $Y=3.05
+ $X2=5.02 $Y2=3.33
r123 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r124 58 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r125 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r126 55 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.005 $Y=3.33
+ $X2=7.92 $Y2=3.33
r127 55 57 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=8.005 $Y=3.33
+ $X2=8.4 $Y2=3.33
r128 54 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r129 54 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r130 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r131 51 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.105 $Y=3.33
+ $X2=6.98 $Y2=3.33
r132 51 53 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.105 $Y=3.33
+ $X2=7.44 $Y2=3.33
r133 50 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.835 $Y=3.33
+ $X2=7.92 $Y2=3.33
r134 50 53 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=7.835 $Y=3.33
+ $X2=7.44 $Y2=3.33
r135 49 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r136 49 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r137 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r138 46 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.22 $Y=3.33
+ $X2=6.055 $Y2=3.33
r139 46 48 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.22 $Y=3.33
+ $X2=6.48 $Y2=3.33
r140 45 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.855 $Y=3.33
+ $X2=6.98 $Y2=3.33
r141 45 48 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.855 $Y=3.33
+ $X2=6.48 $Y2=3.33
r142 44 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r143 44 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r144 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r145 41 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.185 $Y=3.33
+ $X2=5.02 $Y2=3.33
r146 41 43 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.185 $Y=3.33
+ $X2=5.52 $Y2=3.33
r147 40 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.89 $Y=3.33
+ $X2=6.055 $Y2=3.33
r148 40 43 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.89 $Y=3.33
+ $X2=5.52 $Y2=3.33
r149 39 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r150 38 39 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r151 36 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r152 35 38 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=4.56 $Y2=3.33
r153 35 36 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r154 33 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.94 $Y=3.33
+ $X2=0.815 $Y2=3.33
r155 33 35 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.94 $Y=3.33
+ $X2=1.2 $Y2=3.33
r156 32 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=5.02 $Y2=3.33
r157 32 38 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=4.56 $Y2=3.33
r158 30 39 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r159 30 36 0.869652 $w=4.9e-07 $l=3.12e-06 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=1.2 $Y2=3.33
r160 26 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.92 $Y=3.245
+ $X2=7.92 $Y2=3.33
r161 26 28 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=7.92 $Y=3.245
+ $X2=7.92 $Y2=2.805
r162 22 78 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.98 $Y=3.245
+ $X2=6.98 $Y2=3.33
r163 22 24 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=6.98 $Y=3.245
+ $X2=6.98 $Y2=2.805
r164 18 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r165 18 20 37.8001 $w=2.48e-07 $l=8.2e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.425
r166 5 28 600 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=7.785
+ $Y=1.84 $X2=7.92 $Y2=2.805
r167 4 24 600 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=6.885
+ $Y=1.84 $X2=7.02 $Y2=2.805
r168 3 71 600 $w=1.7e-07 $l=1.30618e-06 $layer=licon1_PDIFF $count=1 $X=5.855
+ $Y=1.84 $X2=6.055 $Y2=3.05
r169 2 64 600 $w=1.7e-07 $l=1.30849e-06 $layer=licon1_PDIFF $count=1 $X=4.815
+ $Y=1.84 $X2=5.02 $Y2=3.05
r170 1 20 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=0.64
+ $Y=1.96 $X2=0.775 $Y2=2.425
.ends

.subckt PM_SKY130_FD_SC_MS__XOR2_4%A_514_368# 1 2 3 4 5 6 7 24 26 27 30 32 36 38
+ 39 40 44 48 49 57 58 64 66
c110 39 0 1.47912e-19 $X=6.57 $Y=2.625
c111 32 0 9.06279e-20 $X=4.415 $Y=2.99
r112 56 58 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=5.54 $Y=2.802
+ $X2=5.705 $Y2=2.802
r113 56 57 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=5.54 $Y=2.802
+ $X2=5.375 $Y2=2.802
r114 52 53 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=4.54 $Y=2.8
+ $X2=4.54 $Y2=2.99
r115 49 52 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.54 $Y=2.71 $X2=4.54
+ $Y2=2.8
r116 45 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.635 $Y=2.375
+ $X2=7.47 $Y2=2.375
r117 44 66 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.205 $Y=2.375
+ $X2=8.37 $Y2=2.375
r118 44 45 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.205 $Y=2.375
+ $X2=7.635 $Y2=2.375
r119 41 60 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.655 $Y=2.375
+ $X2=6.57 $Y2=2.375
r120 40 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.305 $Y=2.375
+ $X2=7.47 $Y2=2.375
r121 40 41 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=7.305 $Y=2.375
+ $X2=6.655 $Y2=2.375
r122 39 62 3.40825 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=6.57 $Y=2.625
+ $X2=6.57 $Y2=2.802
r123 38 60 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.57 $Y=2.46
+ $X2=6.57 $Y2=2.375
r124 38 39 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.57 $Y=2.46
+ $X2=6.57 $Y2=2.625
r125 36 62 3.40825 $w=1.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=6.485 $Y=2.71
+ $X2=6.57 $Y2=2.802
r126 36 58 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=6.485 $Y=2.71
+ $X2=5.705 $Y2=2.71
r127 35 49 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.665 $Y=2.71
+ $X2=4.54 $Y2=2.71
r128 35 57 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.665 $Y=2.71
+ $X2=5.375 $Y2=2.71
r129 33 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=2.99
+ $X2=3.6 $Y2=2.99
r130 32 53 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.415 $Y=2.99
+ $X2=4.54 $Y2=2.99
r131 32 33 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.415 $Y=2.99
+ $X2=3.685 $Y2=2.99
r132 28 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=2.905 $X2=3.6
+ $Y2=2.99
r133 28 30 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.6 $Y=2.905
+ $X2=3.6 $Y2=2.8
r134 26 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=2.99
+ $X2=3.6 $Y2=2.99
r135 26 27 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.515 $Y=2.99
+ $X2=2.785 $Y2=2.99
r136 22 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.66 $Y=2.905
+ $X2=2.785 $Y2=2.99
r137 22 24 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=2.66 $Y=2.905
+ $X2=2.66 $Y2=2.355
r138 7 66 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=8.235
+ $Y=1.84 $X2=8.37 $Y2=2.455
r139 6 64 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=7.335
+ $Y=1.84 $X2=7.47 $Y2=2.455
r140 5 62 600 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.435
+ $Y=1.84 $X2=6.57 $Y2=2.815
r141 5 60 600 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=1 $X=6.435
+ $Y=1.84 $X2=6.57 $Y2=2.455
r142 4 56 600 $w=1.7e-07 $l=1.02528e-06 $layer=licon1_PDIFF $count=1 $X=5.405
+ $Y=1.84 $X2=5.54 $Y2=2.8
r143 3 52 600 $w=1.7e-07 $l=1.02528e-06 $layer=licon1_PDIFF $count=1 $X=4.365
+ $Y=1.84 $X2=4.5 $Y2=2.8
r144 2 30 600 $w=1.7e-07 $l=1.02528e-06 $layer=licon1_PDIFF $count=1 $X=3.465
+ $Y=1.84 $X2=3.6 $Y2=2.8
r145 1 24 300 $w=1.7e-07 $l=5.76346e-07 $layer=licon1_PDIFF $count=2 $X=2.57
+ $Y=1.84 $X2=2.7 $Y2=2.355
.ends

.subckt PM_SKY130_FD_SC_MS__XOR2_4%X 1 2 3 4 5 18 21 22 24 25 27 28 29 32 34 38
+ 40 43 45 50 54 55 56 60 63
c164 29 0 1.05217e-19 $X=6.315 $Y=2.035
c165 24 0 2.92031e-19 $X=6.835 $Y=1.095
r166 59 60 9.22412 $w=4.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.05 $Y=2.51
+ $X2=3.885 $Y2=2.51
r167 56 63 8.42674 $w=4.48e-07 $l=1.35e-07 $layer=LI1_cond $X=4.08 $Y=2.51
+ $X2=4.215 $Y2=2.51
r168 56 59 0.797386 $w=4.48e-07 $l=3e-08 $layer=LI1_cond $X=4.08 $Y=2.51
+ $X2=4.05 $Y2=2.51
r169 50 52 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.375 $Y=0.66
+ $X2=3.375 $Y2=0.765
r170 45 47 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.15 $Y=2.275
+ $X2=3.15 $Y2=2.37
r171 42 43 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=8.42 $Y=1.18
+ $X2=8.42 $Y2=1.95
r172 41 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.015 $Y=1.095
+ $X2=7.93 $Y2=1.095
r173 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.335 $Y=1.095
+ $X2=8.42 $Y2=1.18
r174 40 41 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.335 $Y=1.095
+ $X2=8.015 $Y2=1.095
r175 36 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.93 $Y=1.01
+ $X2=7.93 $Y2=1.095
r176 36 38 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.93 $Y=1.01
+ $X2=7.93 $Y2=0.805
r177 35 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.165 $Y=1.095
+ $X2=7 $Y2=1.095
r178 34 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.845 $Y=1.095
+ $X2=7.93 $Y2=1.095
r179 34 35 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.845 $Y=1.095
+ $X2=7.165 $Y2=1.095
r180 30 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7 $Y=1.01 $X2=7
+ $Y2=1.095
r181 30 32 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=7 $Y=1.01 $X2=7
+ $Y2=0.76
r182 28 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.335 $Y=2.035
+ $X2=8.42 $Y2=1.95
r183 28 29 131.786 $w=1.68e-07 $l=2.02e-06 $layer=LI1_cond $X=8.335 $Y=2.035
+ $X2=6.315 $Y2=2.035
r184 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.23 $Y=2.12
+ $X2=6.315 $Y2=2.035
r185 26 27 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.23 $Y=2.12
+ $X2=6.23 $Y2=2.285
r186 24 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.835 $Y=1.095
+ $X2=7 $Y2=1.095
r187 24 25 167.016 $w=1.68e-07 $l=2.56e-06 $layer=LI1_cond $X=6.835 $Y=1.095
+ $X2=4.275 $Y2=1.095
r188 22 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.145 $Y=2.37
+ $X2=6.23 $Y2=2.285
r189 22 63 125.914 $w=1.68e-07 $l=1.93e-06 $layer=LI1_cond $X=6.145 $Y=2.37
+ $X2=4.215 $Y2=2.37
r190 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.19 $Y=1.01
+ $X2=4.275 $Y2=1.095
r191 20 21 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.19 $Y=0.85
+ $X2=4.19 $Y2=1.01
r192 19 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.54 $Y=0.765
+ $X2=3.375 $Y2=0.765
r193 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.105 $Y=0.765
+ $X2=4.19 $Y2=0.85
r194 18 19 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=4.105 $Y=0.765
+ $X2=3.54 $Y2=0.765
r195 17 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.315 $Y=2.37
+ $X2=3.15 $Y2=2.37
r196 17 60 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.315 $Y=2.37
+ $X2=3.885 $Y2=2.37
r197 5 59 600 $w=1.7e-07 $l=7.34405e-07 $layer=licon1_PDIFF $count=1 $X=3.915
+ $Y=1.84 $X2=4.05 $Y2=2.51
r198 4 45 300 $w=1.7e-07 $l=4.97946e-07 $layer=licon1_PDIFF $count=2 $X=3.015
+ $Y=1.84 $X2=3.15 $Y2=2.275
r199 3 38 182 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_NDIFF $count=1 $X=7.79
+ $Y=0.37 $X2=7.93 $Y2=0.805
r200 2 32 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=6.86
+ $Y=0.37 $X2=7 $Y2=0.76
r201 1 50 182 $w=1.7e-07 $l=5.02867e-07 $layer=licon1_NDIFF $count=1 $X=2.95
+ $Y=0.49 $X2=3.375 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_MS__XOR2_4%VGND 1 2 3 4 5 6 19 21 25 29 33 37 39 40 47
+ 48 49 55 63 67 77 78 84 87 90
r122 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r123 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r124 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r125 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r126 77 78 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r127 75 78 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r128 75 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r129 74 77 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r130 74 75 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r131 72 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.225 $Y=0 $X2=6.06
+ $Y2=0
r132 72 74 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.225 $Y=0
+ $X2=6.48 $Y2=0
r133 71 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r134 71 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r135 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r136 68 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.205 $Y=0 $X2=5.04
+ $Y2=0
r137 68 70 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.205 $Y=0
+ $X2=5.52 $Y2=0
r138 67 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.895 $Y=0 $X2=6.06
+ $Y2=0
r139 67 70 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.895 $Y=0
+ $X2=5.52 $Y2=0
r140 66 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r141 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r142 63 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.875 $Y=0 $X2=5.04
+ $Y2=0
r143 63 65 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.875 $Y=0
+ $X2=4.56 $Y2=0
r144 62 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r145 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r146 59 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.58
+ $Y2=0
r147 59 61 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=3.6
+ $Y2=0
r148 58 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r149 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r150 55 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=0 $X2=2.58
+ $Y2=0
r151 55 57 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.415 $Y=0
+ $X2=2.16 $Y2=0
r152 54 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r153 54 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r154 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r155 51 81 4.03846 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r156 51 53 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=1.2
+ $Y2=0
r157 49 66 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.56 $Y2=0
r158 49 62 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.32 $Y=0 $X2=3.6
+ $Y2=0
r159 47 61 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.72 $Y=0 $X2=3.6
+ $Y2=0
r160 47 48 10.0494 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=3.72 $Y=0 $X2=3.927
+ $Y2=0
r161 46 65 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=4.135 $Y=0
+ $X2=4.56 $Y2=0
r162 46 48 10.0494 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=4.135 $Y=0
+ $X2=3.927 $Y2=0
r163 42 57 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=1.615 $Y=0
+ $X2=2.16 $Y2=0
r164 40 53 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.2
+ $Y2=0
r165 39 44 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.45
+ $Y2=0.325
r166 39 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.615
+ $Y2=0
r167 39 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.285
+ $Y2=0
r168 35 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.06 $Y=0.085
+ $X2=6.06 $Y2=0
r169 35 37 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=6.06 $Y=0.085
+ $X2=6.06 $Y2=0.335
r170 31 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.04 $Y=0.085
+ $X2=5.04 $Y2=0
r171 31 33 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=5.04 $Y=0.085
+ $X2=5.04 $Y2=0.335
r172 27 48 1.57254 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.927 $Y=0.085
+ $X2=3.927 $Y2=0
r173 27 29 7.22012 $w=4.13e-07 $l=2.6e-07 $layer=LI1_cond $X=3.927 $Y=0.085
+ $X2=3.927 $Y2=0.345
r174 23 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=0.085
+ $X2=2.58 $Y2=0
r175 23 25 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.58 $Y=0.085
+ $X2=2.58 $Y2=0.335
r176 19 81 3.10471 $w=2.5e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.22 $Y=0.085
+ $X2=0.172 $Y2=0
r177 19 21 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=0.22 $Y=0.085
+ $X2=0.22 $Y2=0.635
r178 6 37 182 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_NDIFF $count=1 $X=5.84
+ $Y=0.37 $X2=6.06 $Y2=0.335
r179 5 33 182 $w=1.7e-07 $l=2.36854e-07 $layer=licon1_NDIFF $count=1 $X=4.82
+ $Y=0.37 $X2=5.04 $Y2=0.335
r180 4 29 182 $w=1.7e-07 $l=3.245e-07 $layer=licon1_NDIFF $count=1 $X=3.665
+ $Y=0.49 $X2=3.925 $Y2=0.345
r181 3 25 182 $w=1.7e-07 $l=2.87228e-07 $layer=licon1_NDIFF $count=1 $X=2.36
+ $Y=0.49 $X2=2.58 $Y2=0.335
r182 2 44 182 $w=1.7e-07 $l=2.91033e-07 $layer=licon1_NDIFF $count=1 $X=1.23
+ $Y=0.49 $X2=1.45 $Y2=0.325
r183 1 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.49 $X2=0.26 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_MS__XOR2_4%A_877_74# 1 2 3 4 5 20 23 24 25 28 30 34 37
+ 40 41 44
r77 39 41 9.45624 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=5.55 $Y=0.595
+ $X2=5.715 $Y2=0.595
r78 39 40 9.45624 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=5.55 $Y=0.595
+ $X2=5.385 $Y2=0.595
r79 32 34 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=8.36 $Y=0.425
+ $X2=8.36 $Y2=0.675
r80 31 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.665 $Y=0.34
+ $X2=7.5 $Y2=0.34
r81 30 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.195 $Y=0.34
+ $X2=8.36 $Y2=0.425
r82 30 31 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=8.195 $Y=0.34
+ $X2=7.665 $Y2=0.34
r83 26 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.5 $Y=0.425 $X2=7.5
+ $Y2=0.34
r84 26 28 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=7.5 $Y=0.425 $X2=7.5
+ $Y2=0.675
r85 24 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.335 $Y=0.34
+ $X2=7.5 $Y2=0.34
r86 24 25 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.335 $Y=0.34
+ $X2=6.655 $Y2=0.34
r87 23 43 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.53 $Y=0.67 $X2=6.53
+ $Y2=0.755
r88 22 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.53 $Y=0.425
+ $X2=6.655 $Y2=0.34
r89 22 23 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=6.53 $Y=0.425
+ $X2=6.53 $Y2=0.67
r90 20 43 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.405 $Y=0.755
+ $X2=6.53 $Y2=0.755
r91 20 41 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.405 $Y=0.755
+ $X2=5.715 $Y2=0.755
r92 19 37 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.695 $Y=0.755
+ $X2=4.57 $Y2=0.755
r93 19 40 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.695 $Y=0.755
+ $X2=5.385 $Y2=0.755
r94 5 34 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=8.22
+ $Y=0.37 $X2=8.36 $Y2=0.675
r95 4 28 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=7.29
+ $Y=0.37 $X2=7.5 $Y2=0.675
r96 3 43 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=6.43
+ $Y=0.37 $X2=6.57 $Y2=0.675
r97 2 39 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=5.41
+ $Y=0.37 $X2=5.55 $Y2=0.675
r98 1 37 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=4.385
+ $Y=0.37 $X2=4.53 $Y2=0.675
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 a_225_392# B1 a_230_79# VNB nlowvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=1.344e+11p ps=1.7e+06u
M1001 VGND A2 a_52_123# VNB nlowvt w=640000u l=150000u
+  ad=4.426e+11p pd=4.38e+06u as=3.52e+11p ps=3.66e+06u
M1002 X a_225_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=8.412e+11p ps=5.86e+06u
M1003 a_230_79# B2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_135_392# B1 a_225_392# VPB pshort w=1e+06u l=180000u
+  ad=6.3e+11p pd=5.26e+06u as=3e+11p ps=2.6e+06u
M1005 a_135_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_225_392# B2 a_135_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_52_123# A1 a_225_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_225_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1009 VPWR A1 a_135_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_ms__and2_1.spice
* Created: Wed Sep  2 11:56:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__and2_1.pex.spice"
.subckt sky130_fd_sc_ms__and2_1  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1004 A_143_136# N_A_M1004_g N_A_56_136#_M1004_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1376 AS=0.1824 PD=1.14 PS=1.85 NRD=30 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1003 N_VGND_M1003_d N_B_M1003_g A_143_136# VNB NLOWVT L=0.15 W=0.64
+ AD=0.144093 AS=0.1376 PD=1.08522 PS=1.14 NRD=14.988 NRS=30 M=1 R=4.26667
+ SA=75000.7 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1005 N_X_M1005_d N_A_56_136#_M1005_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.166607 PD=2.05 PS=1.25478 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_56_136#_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1344 AS=0.2394 PD=1.16 PS=2.25 NRD=10.5395 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90001.2 A=0.1512 P=2.04 MULT=1
MM1001 N_VPWR_M1001_d N_B_M1001_g N_A_56_136#_M1000_d VPB PSHORT L=0.18 W=0.84
+ AD=0.1578 AS=0.1344 PD=1.26429 PS=1.16 NRD=18.7544 NRS=0 M=1 R=4.66667
+ SA=90000.7 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1002 N_X_M1002_d N_A_56_136#_M1002_g N_VPWR_M1001_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.2104 PD=2.8 PS=1.68571 NRD=0 NRS=0 M=1 R=6.22222 SA=90001
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1708 P=9.28
*
.include "sky130_fd_sc_ms__and2_1.pxi.spice"
*
.ends
*
*

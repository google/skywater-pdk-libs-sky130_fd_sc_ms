* File: sky130_fd_sc_ms__mux4_4.pxi.spice
* Created: Wed Sep  2 12:12:34 2020
* 
x_PM_SKY130_FD_SC_MS__MUX4_4%A1 N_A1_M1003_g N_A1_M1025_g N_A1_M1033_g
+ N_A1_M1004_g A1 A1 N_A1_c_312_n PM_SKY130_FD_SC_MS__MUX4_4%A1
x_PM_SKY130_FD_SC_MS__MUX4_4%A0 N_A0_M1007_g N_A0_M1022_g N_A0_M1023_g
+ N_A0_M1011_g A0 A0 A0 N_A0_c_355_n N_A0_c_356_n PM_SKY130_FD_SC_MS__MUX4_4%A0
x_PM_SKY130_FD_SC_MS__MUX4_4%A_758_306# N_A_758_306#_M1016_s
+ N_A_758_306#_M1013_s N_A_758_306#_M1045_g N_A_758_306#_M1039_g
+ N_A_758_306#_M1049_g N_A_758_306#_M1043_g N_A_758_306#_c_414_n
+ N_A_758_306#_c_415_n N_A_758_306#_M1002_g N_A_758_306#_M1046_g
+ N_A_758_306#_c_416_n N_A_758_306#_M1006_g N_A_758_306#_M1050_g
+ N_A_758_306#_c_417_n N_A_758_306#_c_429_n N_A_758_306#_c_418_n
+ N_A_758_306#_c_524_p N_A_758_306#_c_419_n N_A_758_306#_c_420_n
+ N_A_758_306#_c_421_n N_A_758_306#_c_422_n N_A_758_306#_c_423_n
+ PM_SKY130_FD_SC_MS__MUX4_4%A_758_306#
x_PM_SKY130_FD_SC_MS__MUX4_4%S0 N_S0_M1000_g N_S0_M1009_g N_S0_c_548_n
+ N_S0_c_549_n N_S0_M1042_g N_S0_M1047_g N_S0_c_552_n N_S0_M1016_g N_S0_c_554_n
+ N_S0_M1013_g N_S0_c_556_n N_S0_M1012_g N_S0_M1001_g N_S0_M1041_g N_S0_M1008_g
+ N_S0_c_559_n N_S0_c_560_n N_S0_c_561_n N_S0_c_562_n N_S0_c_563_n N_S0_c_564_n
+ S0 S0 S0 N_S0_c_566_n PM_SKY130_FD_SC_MS__MUX4_4%S0
x_PM_SKY130_FD_SC_MS__MUX4_4%A2 N_A2_M1036_g N_A2_M1021_g N_A2_M1038_g
+ N_A2_M1040_g A2 A2 N_A2_c_724_n PM_SKY130_FD_SC_MS__MUX4_4%A2
x_PM_SKY130_FD_SC_MS__MUX4_4%A3 N_A3_M1018_g N_A3_M1005_g N_A3_c_779_n
+ N_A3_M1031_g N_A3_M1024_g N_A3_c_780_n N_A3_c_781_n A3 A3 N_A3_c_783_n
+ PM_SKY130_FD_SC_MS__MUX4_4%A3
x_PM_SKY130_FD_SC_MS__MUX4_4%S1 N_S1_M1017_g N_S1_M1032_g N_S1_M1019_g
+ N_S1_M1037_g N_S1_c_837_n N_S1_c_838_n N_S1_M1014_g N_S1_M1044_g N_S1_c_840_n
+ N_S1_c_841_n N_S1_c_842_n S1 N_S1_c_843_n N_S1_c_844_n S1 N_S1_c_845_n
+ N_S1_c_846_n PM_SKY130_FD_SC_MS__MUX4_4%S1
x_PM_SKY130_FD_SC_MS__MUX4_4%A_2489_347# N_A_2489_347#_M1014_s
+ N_A_2489_347#_M1044_s N_A_2489_347#_c_955_n N_A_2489_347#_M1028_g
+ N_A_2489_347#_M1015_g N_A_2489_347#_c_956_n N_A_2489_347#_M1029_g
+ N_A_2489_347#_M1048_g N_A_2489_347#_c_957_n N_A_2489_347#_c_958_n
+ N_A_2489_347#_c_951_n N_A_2489_347#_c_952_n N_A_2489_347#_c_953_n
+ N_A_2489_347#_c_962_n N_A_2489_347#_c_954_n
+ PM_SKY130_FD_SC_MS__MUX4_4%A_2489_347#
x_PM_SKY130_FD_SC_MS__MUX4_4%A_2199_74# N_A_2199_74#_M1017_s
+ N_A_2199_74#_M1019_s N_A_2199_74#_M1048_d N_A_2199_74#_M1032_d
+ N_A_2199_74#_M1037_d N_A_2199_74#_M1029_s N_A_2199_74#_M1010_g
+ N_A_2199_74#_M1020_g N_A_2199_74#_M1026_g N_A_2199_74#_M1027_g
+ N_A_2199_74#_M1030_g N_A_2199_74#_M1035_g N_A_2199_74#_M1034_g
+ N_A_2199_74#_M1051_g N_A_2199_74#_c_1042_n N_A_2199_74#_c_1071_n
+ N_A_2199_74#_c_1060_n N_A_2199_74#_c_1061_n N_A_2199_74#_c_1096_n
+ N_A_2199_74#_c_1043_n N_A_2199_74#_c_1077_n N_A_2199_74#_c_1044_n
+ N_A_2199_74#_c_1062_n N_A_2199_74#_c_1063_n N_A_2199_74#_c_1045_n
+ N_A_2199_74#_c_1046_n N_A_2199_74#_c_1047_n N_A_2199_74#_c_1048_n
+ N_A_2199_74#_c_1049_n N_A_2199_74#_c_1050_n N_A_2199_74#_c_1088_n
+ N_A_2199_74#_c_1051_n N_A_2199_74#_c_1052_n N_A_2199_74#_c_1053_n
+ N_A_2199_74#_c_1054_n PM_SKY130_FD_SC_MS__MUX4_4%A_2199_74#
x_PM_SKY130_FD_SC_MS__MUX4_4%VPWR N_VPWR_M1003_s N_VPWR_M1004_s N_VPWR_M1011_d
+ N_VPWR_M1013_d N_VPWR_M1036_s N_VPWR_M1038_s N_VPWR_M1024_s N_VPWR_M1044_d
+ N_VPWR_M1026_s N_VPWR_M1034_s N_VPWR_c_1241_n N_VPWR_c_1242_n N_VPWR_c_1243_n
+ N_VPWR_c_1244_n N_VPWR_c_1245_n N_VPWR_c_1246_n N_VPWR_c_1247_n
+ N_VPWR_c_1248_n N_VPWR_c_1249_n N_VPWR_c_1250_n N_VPWR_c_1251_n
+ N_VPWR_c_1252_n N_VPWR_c_1253_n N_VPWR_c_1254_n N_VPWR_c_1255_n
+ N_VPWR_c_1256_n N_VPWR_c_1257_n N_VPWR_c_1258_n VPWR N_VPWR_c_1259_n
+ N_VPWR_c_1260_n N_VPWR_c_1261_n N_VPWR_c_1262_n N_VPWR_c_1263_n
+ N_VPWR_c_1264_n N_VPWR_c_1265_n N_VPWR_c_1266_n N_VPWR_c_1267_n
+ N_VPWR_c_1240_n PM_SKY130_FD_SC_MS__MUX4_4%VPWR
x_PM_SKY130_FD_SC_MS__MUX4_4%A_119_392# N_A_119_392#_M1003_d
+ N_A_119_392#_M1045_d N_A_119_392#_c_1422_n N_A_119_392#_c_1423_n
+ N_A_119_392#_c_1424_n N_A_119_392#_c_1425_n N_A_119_392#_c_1420_n
+ N_A_119_392#_c_1421_n N_A_119_392#_c_1428_n
+ PM_SKY130_FD_SC_MS__MUX4_4%A_119_392#
x_PM_SKY130_FD_SC_MS__MUX4_4%A_299_392# N_A_299_392#_M1007_s
+ N_A_299_392#_M1000_s N_A_299_392#_c_1483_n N_A_299_392#_c_1484_n
+ N_A_299_392#_c_1485_n N_A_299_392#_c_1491_n
+ PM_SKY130_FD_SC_MS__MUX4_4%A_299_392#
x_PM_SKY130_FD_SC_MS__MUX4_4%A_509_392# N_A_509_392#_M1009_d
+ N_A_509_392#_M1047_d N_A_509_392#_M1043_s N_A_509_392#_M1015_s
+ N_A_509_392#_M1000_d N_A_509_392#_M1042_d N_A_509_392#_M1049_s
+ N_A_509_392#_M1032_s N_A_509_392#_c_1524_n N_A_509_392#_c_1512_n
+ N_A_509_392#_c_1525_n N_A_509_392#_c_1513_n N_A_509_392#_c_1514_n
+ N_A_509_392#_c_1526_n N_A_509_392#_c_1515_n N_A_509_392#_c_1527_n
+ N_A_509_392#_c_1516_n N_A_509_392#_c_1517_n N_A_509_392#_c_1599_n
+ N_A_509_392#_c_1528_n N_A_509_392#_c_1518_n N_A_509_392#_c_1529_n
+ N_A_509_392#_c_1519_n N_A_509_392#_c_1520_n N_A_509_392#_c_1521_n
+ N_A_509_392#_c_1604_n N_A_509_392#_c_1530_n N_A_509_392#_c_1531_n
+ N_A_509_392#_c_1532_n N_A_509_392#_c_1533_n N_A_509_392#_c_1522_n
+ N_A_509_392#_c_1523_n PM_SKY130_FD_SC_MS__MUX4_4%A_509_392#
x_PM_SKY130_FD_SC_MS__MUX4_4%A_1191_121# N_A_1191_121#_M1002_s
+ N_A_1191_121#_M1006_s N_A_1191_121#_M1041_s N_A_1191_121#_M1017_d
+ N_A_1191_121#_M1046_s N_A_1191_121#_M1050_s N_A_1191_121#_M1008_s
+ N_A_1191_121#_M1028_d N_A_1191_121#_c_1699_n N_A_1191_121#_c_1700_n
+ N_A_1191_121#_c_1709_n N_A_1191_121#_c_1710_n N_A_1191_121#_c_1727_n
+ N_A_1191_121#_c_1711_n N_A_1191_121#_c_1701_n N_A_1191_121#_c_1746_n
+ N_A_1191_121#_c_1702_n N_A_1191_121#_c_1834_p N_A_1191_121#_c_1703_n
+ N_A_1191_121#_c_1713_n N_A_1191_121#_c_1704_n N_A_1191_121#_c_1715_n
+ N_A_1191_121#_c_1705_n N_A_1191_121#_c_1706_n N_A_1191_121#_c_1716_n
+ N_A_1191_121#_c_1717_n N_A_1191_121#_c_1787_n N_A_1191_121#_c_1707_n
+ N_A_1191_121#_c_1718_n N_A_1191_121#_c_1708_n N_A_1191_121#_c_1719_n
+ PM_SKY130_FD_SC_MS__MUX4_4%A_1191_121#
x_PM_SKY130_FD_SC_MS__MUX4_4%A_1288_377# N_A_1288_377#_M1046_d
+ N_A_1288_377#_M1005_d N_A_1288_377#_c_1875_n N_A_1288_377#_c_1871_n
+ N_A_1288_377#_c_1872_n N_A_1288_377#_c_1873_n N_A_1288_377#_c_1886_n
+ N_A_1288_377#_c_1874_n PM_SKY130_FD_SC_MS__MUX4_4%A_1288_377#
x_PM_SKY130_FD_SC_MS__MUX4_4%A_1468_377# N_A_1468_377#_M1001_d
+ N_A_1468_377#_M1036_d N_A_1468_377#_c_1926_n N_A_1468_377#_c_1928_n
+ PM_SKY130_FD_SC_MS__MUX4_4%A_1468_377#
x_PM_SKY130_FD_SC_MS__MUX4_4%X N_X_M1020_d N_X_M1035_d N_X_M1010_d N_X_M1030_d
+ N_X_c_1954_n N_X_c_1947_n N_X_c_1955_n N_X_c_1956_n N_X_c_1948_n N_X_c_1949_n
+ N_X_c_1957_n N_X_c_1950_n N_X_c_1958_n N_X_c_1951_n N_X_c_1959_n N_X_c_1952_n
+ X X PM_SKY130_FD_SC_MS__MUX4_4%X
x_PM_SKY130_FD_SC_MS__MUX4_4%VGND N_VGND_M1025_d N_VGND_M1033_d N_VGND_M1023_s
+ N_VGND_M1016_d N_VGND_M1021_s N_VGND_M1040_s N_VGND_M1031_s N_VGND_M1014_d
+ N_VGND_M1027_s N_VGND_M1051_s N_VGND_c_2030_n N_VGND_c_2031_n N_VGND_c_2032_n
+ N_VGND_c_2033_n N_VGND_c_2034_n N_VGND_c_2072_n N_VGND_c_2035_n
+ N_VGND_c_2036_n N_VGND_c_2037_n N_VGND_c_2038_n N_VGND_c_2039_n
+ N_VGND_c_2040_n N_VGND_c_2041_n N_VGND_c_2042_n N_VGND_c_2043_n
+ N_VGND_c_2044_n N_VGND_c_2045_n N_VGND_c_2046_n N_VGND_c_2047_n
+ N_VGND_c_2048_n N_VGND_c_2049_n VGND N_VGND_c_2050_n N_VGND_c_2051_n
+ N_VGND_c_2052_n N_VGND_c_2053_n N_VGND_c_2054_n N_VGND_c_2055_n
+ N_VGND_c_2056_n N_VGND_c_2057_n N_VGND_c_2058_n
+ PM_SKY130_FD_SC_MS__MUX4_4%VGND
x_PM_SKY130_FD_SC_MS__MUX4_4%A_114_126# N_A_114_126#_M1025_s
+ N_A_114_126#_M1009_s N_A_114_126#_c_2232_n N_A_114_126#_c_2233_n
+ N_A_114_126#_c_2234_n N_A_114_126#_c_2235_n N_A_114_126#_c_2236_n
+ N_A_114_126#_c_2247_n N_A_114_126#_c_2237_n
+ PM_SKY130_FD_SC_MS__MUX4_4%A_114_126#
x_PM_SKY130_FD_SC_MS__MUX4_4%A_299_126# N_A_299_126#_M1022_d
+ N_A_299_126#_M1039_d N_A_299_126#_c_2282_n N_A_299_126#_c_2283_n
+ N_A_299_126#_c_2284_n N_A_299_126#_c_2285_n N_A_299_126#_c_2286_n
+ PM_SKY130_FD_SC_MS__MUX4_4%A_299_126#
x_PM_SKY130_FD_SC_MS__MUX4_4%A_1278_121# N_A_1278_121#_M1002_d
+ N_A_1278_121#_M1021_d N_A_1278_121#_c_2324_n N_A_1278_121#_c_2325_n
+ N_A_1278_121#_c_2326_n N_A_1278_121#_c_2327_n N_A_1278_121#_c_2328_n
+ N_A_1278_121#_c_2329_n N_A_1278_121#_c_2330_n
+ PM_SKY130_FD_SC_MS__MUX4_4%A_1278_121#
x_PM_SKY130_FD_SC_MS__MUX4_4%A_1450_121# N_A_1450_121#_M1012_d
+ N_A_1450_121#_M1018_d N_A_1450_121#_c_2377_n N_A_1450_121#_c_2378_n
+ N_A_1450_121#_c_2379_n N_A_1450_121#_c_2380_n N_A_1450_121#_c_2381_n
+ PM_SKY130_FD_SC_MS__MUX4_4%A_1450_121#
cc_1 VNB N_A1_M1025_g 0.0253008f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.95
cc_2 VNB N_A1_M1033_g 0.0200691f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.95
cc_3 VNB A1 0.00939308f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_A1_c_312_n 0.0369025f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.615
cc_5 VNB N_A0_M1022_g 0.0215995f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.95
cc_6 VNB N_A0_M1023_g 0.0253354f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.95
cc_7 VNB A0 0.00608988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A0_c_355_n 0.0211887f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.615
cc_9 VNB N_A0_c_356_n 0.0196575f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.615
cc_10 VNB N_A_758_306#_M1039_g 0.0170312f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.78
cc_11 VNB N_A_758_306#_M1043_g 0.020382f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.615
cc_12 VNB N_A_758_306#_c_414_n 0.0246973f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.615
cc_13 VNB N_A_758_306#_c_415_n 0.0194199f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.615
cc_14 VNB N_A_758_306#_c_416_n 0.014905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_758_306#_c_417_n 0.0143874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_758_306#_c_418_n 0.00207742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_758_306#_c_419_n 0.0298973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_758_306#_c_420_n 0.00188816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_758_306#_c_421_n 0.0218401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_758_306#_c_422_n 0.0150421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_758_306#_c_423_n 0.0478629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_S0_M1000_g 0.0121349f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_23 VNB N_S0_M1009_g 0.0240024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_S0_c_548_n 0.0191625f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.45
cc_25 VNB N_S0_c_549_n 0.012611f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.95
cc_26 VNB N_S0_M1042_g 0.0108562f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.78
cc_27 VNB N_S0_M1047_g 0.0228453f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_28 VNB N_S0_c_552_n 0.124248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_S0_M1016_g 0.0129586f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.615
cc_30 VNB N_S0_c_554_n 0.0085432f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.615
cc_31 VNB N_S0_M1013_g 0.0245856f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.615
cc_32 VNB N_S0_c_556_n 0.210692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_S0_M1012_g 0.015698f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_34 VNB N_S0_M1041_g 0.0199871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_S0_c_559_n 0.0674609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_S0_c_560_n 0.0143755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_S0_c_561_n 0.0116324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_S0_c_562_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_S0_c_563_n 0.00732516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_S0_c_564_n 0.0258376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB S0 0.00433756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_S0_c_566_n 0.0272342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A2_M1036_g 0.00379398f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_44 VNB N_A2_M1021_g 0.0272771f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.95
cc_45 VNB N_A2_M1038_g 0.00342908f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.95
cc_46 VNB N_A2_M1040_g 0.0232221f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.46
cc_47 VNB A2 0.00398279f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_48 VNB N_A2_c_724_n 0.0521622f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.615
cc_49 VNB N_A3_M1018_g 0.0343392f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_50 VNB N_A3_c_779_n 0.0173391f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.45
cc_51 VNB N_A3_c_780_n 0.0127568f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_52 VNB N_A3_c_781_n 0.0149455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB A3 0.00455884f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.615
cc_54 VNB N_A3_c_783_n 0.0315199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_S1_M1017_g 0.0250832f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.46
cc_56 VNB N_S1_M1032_g 0.00889551f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.95
cc_57 VNB N_S1_M1019_g 0.0246191f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.95
cc_58 VNB N_S1_M1037_g 0.00825093f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.46
cc_59 VNB N_S1_c_837_n 0.0298116f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_60 VNB N_S1_c_838_n 0.0209511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_S1_M1044_g 0.0079111f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.615
cc_62 VNB N_S1_c_840_n 0.055013f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.615
cc_63 VNB N_S1_c_841_n 0.0131301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_S1_c_842_n 0.026117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_S1_c_843_n 0.0348594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_S1_c_844_n 0.0364686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_S1_c_845_n 0.00294663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_S1_c_846_n 0.00253735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_2489_347#_M1015_g 0.0350434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_2489_347#_M1048_g 0.0395546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_2489_347#_c_951_n 0.00698854f $X=-0.19 $Y=-0.245 $X2=0.24
+ $Y2=1.615
cc_72 VNB N_A_2489_347#_c_952_n 7.73014e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_2489_347#_c_953_n 0.0268228f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_74 VNB N_A_2489_347#_c_954_n 0.00368999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_2199_74#_M1010_g 0.0016648f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.615
cc_76 VNB N_A_2199_74#_M1020_g 0.0242761f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.615
cc_77 VNB N_A_2199_74#_M1026_g 0.00160182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_2199_74#_M1027_g 0.0203684f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_79 VNB N_A_2199_74#_M1030_g 0.0016013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_2199_74#_M1035_g 0.0209263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_2199_74#_M1034_g 0.00169679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_2199_74#_M1051_g 0.0232593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_2199_74#_c_1042_n 0.00856582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_2199_74#_c_1043_n 0.00365532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_2199_74#_c_1044_n 0.0026202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_2199_74#_c_1045_n 0.00589658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_2199_74#_c_1046_n 0.0160232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_2199_74#_c_1047_n 0.00273158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_2199_74#_c_1048_n 0.00150988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_2199_74#_c_1049_n 0.012286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_2199_74#_c_1050_n 0.00378272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_2199_74#_c_1051_n 9.79592e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_2199_74#_c_1052_n 0.00151123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_2199_74#_c_1053_n 0.00325932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_2199_74#_c_1054_n 0.0925308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VPWR_c_1240_n 0.701046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_119_392#_c_1420_n 0.00638497f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.46
cc_98 VNB N_A_119_392#_c_1421_n 0.00221343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_509_392#_c_1512_n 0.00921432f $X=-0.19 $Y=-0.245 $X2=0.925
+ $Y2=1.615
cc_100 VNB N_A_509_392#_c_1513_n 0.00340257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_509_392#_c_1514_n 0.016329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_509_392#_c_1515_n 0.00636936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_509_392#_c_1516_n 0.00281722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_509_392#_c_1517_n 5.89755e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_509_392#_c_1518_n 0.0108906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_509_392#_c_1519_n 2.82947e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_509_392#_c_1520_n 0.00167754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_509_392#_c_1521_n 0.00269263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_509_392#_c_1522_n 0.00133979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_509_392#_c_1523_n 0.00187902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_1191_121#_c_1699_n 0.00217675f $X=-0.19 $Y=-0.245 $X2=0.725
+ $Y2=1.615
cc_112 VNB N_A_1191_121#_c_1700_n 0.00619748f $X=-0.19 $Y=-0.245 $X2=0.925
+ $Y2=1.615
cc_113 VNB N_A_1191_121#_c_1701_n 0.00140514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_1191_121#_c_1702_n 0.00347953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_1191_121#_c_1703_n 0.00196259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_1191_121#_c_1704_n 0.0279051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_1191_121#_c_1705_n 0.0034847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_1191_121#_c_1706_n 0.00905591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_1191_121#_c_1707_n 0.00101203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_1191_121#_c_1708_n 0.00157069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_X_c_1947_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.615
cc_122 VNB N_X_c_1948_n 0.00275044f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.615
cc_123 VNB N_X_c_1949_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.615
cc_124 VNB N_X_c_1950_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_X_c_1951_n 0.0087474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_X_c_1952_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB X 0.0265224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2030_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2031_n 0.0122963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2032_n 0.0415587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2033_n 0.00303884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2034_n 0.00401119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2035_n 0.0109437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2036_n 0.0136696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2037_n 0.00420208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2038_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2039_n 0.0109995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2040_n 0.00852643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2041_n 0.00420208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2042_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2043_n 0.0257769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2044_n 0.0134389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2045_n 0.0670697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2046_n 0.0163794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2047_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2048_n 0.0967389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2049_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2050_n 0.0391102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2051_n 0.0737216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2052_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2053_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2054_n 0.0063135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2055_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2056_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2057_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2058_n 0.831397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_A_114_126#_c_2232_n 0.00135554f $X=-0.19 $Y=-0.245 $X2=0.925
+ $Y2=1.45
cc_158 VNB N_A_114_126#_c_2233_n 0.0218796f $X=-0.19 $Y=-0.245 $X2=0.925
+ $Y2=0.95
cc_159 VNB N_A_114_126#_c_2234_n 0.00488309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_A_114_126#_c_2235_n 0.00331078f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.46
cc_161 VNB N_A_114_126#_c_2236_n 9.57738e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VNB N_A_114_126#_c_2237_n 0.00821615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_A_299_126#_c_2282_n 0.00949813f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=0.95
cc_164 VNB N_A_299_126#_c_2283_n 0.01887f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.45
cc_165 VNB N_A_299_126#_c_2284_n 0.00111857f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=1.78
cc_166 VNB N_A_299_126#_c_2285_n 0.00202937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_A_299_126#_c_2286_n 0.00574177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_A_1278_121#_c_2324_n 0.00265586f $X=-0.19 $Y=-0.245 $X2=0.925
+ $Y2=1.45
cc_169 VNB N_A_1278_121#_c_2325_n 0.0291012f $X=-0.19 $Y=-0.245 $X2=0.925
+ $Y2=0.95
cc_170 VNB N_A_1278_121#_c_2326_n 0.00341436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_A_1278_121#_c_2327_n 0.00206083f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.46
cc_172 VNB N_A_1278_121#_c_2328_n 0.00409716f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=2.46
cc_173 VNB N_A_1278_121#_c_2329_n 0.00151359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_174 VNB N_A_1278_121#_c_2330_n 0.00204804f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_175 VNB N_A_1450_121#_c_2377_n 0.00529172f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=0.95
cc_176 VNB N_A_1450_121#_c_2378_n 0.027156f $X=-0.19 $Y=-0.245 $X2=0.925
+ $Y2=1.45
cc_177 VNB N_A_1450_121#_c_2379_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.955
+ $Y2=1.78
cc_178 VNB N_A_1450_121#_c_2380_n 0.00187699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_179 VNB N_A_1450_121#_c_2381_n 0.00310731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_180 VPB N_A1_M1003_g 0.028312f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_181 VPB N_A1_M1004_g 0.0228738f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.46
cc_182 VPB A1 0.00572761f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_183 VPB N_A1_c_312_n 0.024504f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.615
cc_184 VPB N_A0_M1007_g 0.0215995f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_185 VPB N_A0_M1011_g 0.024574f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.46
cc_186 VPB A0 0.00431663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A0_c_355_n 0.0153453f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.615
cc_188 VPB N_A0_c_356_n 0.0167624f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.615
cc_189 VPB N_A_758_306#_M1045_g 0.0266838f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.45
cc_190 VPB N_A_758_306#_M1049_g 0.0321359f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_191 VPB N_A_758_306#_c_414_n 0.00418894f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.615
cc_192 VPB N_A_758_306#_M1046_g 0.0272367f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_193 VPB N_A_758_306#_M1050_g 0.021132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_758_306#_c_429_n 0.0156426f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_758_306#_c_418_n 5.65058e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_758_306#_c_419_n 0.012178f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_758_306#_c_420_n 5.97595e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_758_306#_c_422_n 0.00808002f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_758_306#_c_423_n 0.0123391f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_S0_M1000_g 0.0312412f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_201 VPB N_S0_M1042_g 0.0281133f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.78
cc_202 VPB N_S0_M1013_g 0.030717f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.615
cc_203 VPB N_S0_M1001_g 0.0196637f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_S0_M1008_g 0.0252259f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_S0_c_564_n 0.019332f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB S0 0.00850506f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_S0_c_566_n 0.00815027f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A2_M1036_g 0.0352421f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.46
cc_209 VPB N_A2_M1038_g 0.0307768f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.95
cc_210 VPB A2 0.00397864f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_211 VPB N_A3_M1005_g 0.0249148f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.95
cc_212 VPB N_A3_M1024_g 0.0246493f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.46
cc_213 VPB A3 0.00245853f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.615
cc_214 VPB N_A3_c_783_n 0.0168597f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_S1_M1032_g 0.0342236f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.95
cc_216 VPB N_S1_M1037_g 0.0294378f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.46
cc_217 VPB N_S1_M1044_g 0.0271421f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.615
cc_218 VPB N_S1_c_845_n 0.00376745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_2489_347#_c_955_n 0.016749f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.95
cc_220 VPB N_A_2489_347#_c_956_n 0.0223856f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.46
cc_221 VPB N_A_2489_347#_c_957_n 0.0219737f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.615
cc_222 VPB N_A_2489_347#_c_958_n 0.0223372f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.615
cc_223 VPB N_A_2489_347#_c_951_n 0.00106366f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_224 VPB N_A_2489_347#_c_952_n 0.00189656f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_A_2489_347#_c_953_n 0.048189f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_226 VPB N_A_2489_347#_c_962_n 0.00441519f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_2199_74#_M1010_g 0.0235202f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.615
cc_228 VPB N_A_2199_74#_M1026_g 0.0226708f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_2199_74#_M1030_g 0.0226671f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_2199_74#_M1034_g 0.0240888f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_2199_74#_c_1042_n 0.00977476f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_2199_74#_c_1060_n 0.00187959f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_2199_74#_c_1061_n 0.00223315f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_2199_74#_c_1062_n 0.00258185f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_2199_74#_c_1063_n 0.0135475f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1241_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1242_n 0.0513874f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_238 VPB N_VPWR_c_1243_n 0.00554449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1244_n 0.0117927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1245_n 0.0223252f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1246_n 0.00830185f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1247_n 0.00977897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1248_n 0.0081889f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1249_n 0.0131478f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1250_n 0.0438927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1251_n 0.0141519f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1252_n 0.0195396f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1253_n 0.0196689f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1254_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1255_n 0.092707f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1256_n 0.00614127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1257_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1258_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1259_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1260_n 0.0194914f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1261_n 0.0753721f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1262_n 0.0634408f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1263_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1264_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1265_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1266_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1267_n 0.0141887f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1240_n 0.177152f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_A_119_392#_c_1422_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.95
cc_265 VPB N_A_119_392#_c_1423_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.45
cc_266 VPB N_A_119_392#_c_1424_n 0.00738029f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.95
cc_267 VPB N_A_119_392#_c_1425_n 0.00502504f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.46
cc_268 VPB N_A_119_392#_c_1420_n 0.0102103f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.46
cc_269 VPB N_A_119_392#_c_1421_n 0.00118275f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_A_119_392#_c_1428_n 0.00292075f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_A_299_392#_c_1483_n 0.00834688f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.45
cc_272 VPB N_A_299_392#_c_1484_n 0.00265468f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.78
cc_273 VPB N_A_299_392#_c_1485_n 0.00275605f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_A_509_392#_c_1524_n 0.00210043f $X=-0.19 $Y=1.66 $X2=0.725
+ $Y2=1.615
cc_275 VPB N_A_509_392#_c_1525_n 0.00265247f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_A_509_392#_c_1526_n 0.00675638f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_A_509_392#_c_1527_n 0.00712058f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_A_509_392#_c_1528_n 0.00668636f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_A_509_392#_c_1529_n 0.0021475f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_A_509_392#_c_1530_n 0.0328248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_A_509_392#_c_1531_n 0.00237732f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_A_509_392#_c_1532_n 0.00344159f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_283 VPB N_A_509_392#_c_1533_n 7.8154e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_284 VPB N_A_509_392#_c_1522_n 0.00269527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 VPB N_A_509_392#_c_1523_n 0.00248628f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_286 VPB N_A_1191_121#_c_1709_n 0.00343247f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_287 VPB N_A_1191_121#_c_1710_n 0.0100835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_288 VPB N_A_1191_121#_c_1711_n 0.00321228f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_289 VPB N_A_1191_121#_c_1702_n 0.00331537f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_290 VPB N_A_1191_121#_c_1713_n 0.0391801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_291 VPB N_A_1191_121#_c_1704_n 0.00685901f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_292 VPB N_A_1191_121#_c_1715_n 0.0175193f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_293 VPB N_A_1191_121#_c_1716_n 0.0177838f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_294 VPB N_A_1191_121#_c_1717_n 0.00348146f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_295 VPB N_A_1191_121#_c_1718_n 2.03678e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_296 VPB N_A_1191_121#_c_1719_n 0.00961975f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_297 VPB N_A_1288_377#_c_1871_n 0.0191209f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.95
cc_298 VPB N_A_1288_377#_c_1872_n 0.00484594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_299 VPB N_A_1288_377#_c_1873_n 0.00754673f $X=-0.19 $Y=1.66 $X2=0.955
+ $Y2=1.78
cc_300 VPB N_A_1288_377#_c_1874_n 0.00793561f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_301 VPB N_A_1468_377#_c_1926_n 0.00582192f $X=-0.19 $Y=1.66 $X2=0.925
+ $Y2=1.45
cc_302 VPB N_X_c_1954_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.46
cc_303 VPB N_X_c_1955_n 0.00249468f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.615
cc_304 VPB N_X_c_1956_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.615
cc_305 VPB N_X_c_1957_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_306 VPB N_X_c_1958_n 0.0100349f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_307 VPB N_X_c_1959_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_308 VPB X 0.00728633f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_309 N_A1_M1004_g N_A0_M1007_g 0.0225081f $X=0.955 $Y=2.46 $X2=0 $Y2=0
cc_310 N_A1_M1033_g N_A0_M1022_g 0.0115976f $X=0.925 $Y=0.95 $X2=0 $Y2=0
cc_311 N_A1_c_312_n N_A0_M1022_g 9.69146e-19 $X=0.955 $Y=1.615 $X2=0 $Y2=0
cc_312 A1 A0 0.0247408f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_313 N_A1_c_312_n A0 0.00388406f $X=0.955 $Y=1.615 $X2=0 $Y2=0
cc_314 A1 N_A0_c_355_n 2.15092e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_315 N_A1_c_312_n N_A0_c_355_n 0.0225081f $X=0.955 $Y=1.615 $X2=0 $Y2=0
cc_316 N_A1_M1003_g N_VPWR_c_1242_n 0.0052517f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_317 A1 N_VPWR_c_1242_n 0.0205478f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_318 N_A1_c_312_n N_VPWR_c_1242_n 0.00335457f $X=0.955 $Y=1.615 $X2=0 $Y2=0
cc_319 N_A1_M1004_g N_VPWR_c_1243_n 0.002979f $X=0.955 $Y=2.46 $X2=0 $Y2=0
cc_320 N_A1_M1003_g N_VPWR_c_1259_n 0.005209f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_321 N_A1_M1004_g N_VPWR_c_1259_n 0.005209f $X=0.955 $Y=2.46 $X2=0 $Y2=0
cc_322 N_A1_M1003_g N_VPWR_c_1240_n 0.00986008f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_323 N_A1_M1004_g N_VPWR_c_1240_n 0.00982376f $X=0.955 $Y=2.46 $X2=0 $Y2=0
cc_324 N_A1_M1003_g N_A_119_392#_c_1422_n 0.00292762f $X=0.505 $Y=2.46 $X2=0
+ $Y2=0
cc_325 N_A1_M1004_g N_A_119_392#_c_1422_n 0.0014691f $X=0.955 $Y=2.46 $X2=0
+ $Y2=0
cc_326 A1 N_A_119_392#_c_1422_n 0.0271639f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_327 N_A1_c_312_n N_A_119_392#_c_1422_n 0.00215577f $X=0.955 $Y=1.615 $X2=0
+ $Y2=0
cc_328 N_A1_M1003_g N_A_119_392#_c_1423_n 0.011014f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_329 N_A1_M1004_g N_A_119_392#_c_1423_n 0.0116888f $X=0.955 $Y=2.46 $X2=0
+ $Y2=0
cc_330 N_A1_M1004_g N_A_119_392#_c_1424_n 0.017339f $X=0.955 $Y=2.46 $X2=0 $Y2=0
cc_331 A1 N_VGND_c_2031_n 0.0206322f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_332 N_A1_c_312_n N_VGND_c_2031_n 0.00337787f $X=0.955 $Y=1.615 $X2=0 $Y2=0
cc_333 N_A1_M1025_g N_VGND_c_2032_n 0.00290289f $X=0.495 $Y=0.95 $X2=0 $Y2=0
cc_334 N_A1_M1025_g N_VGND_c_2033_n 0.0145041f $X=0.495 $Y=0.95 $X2=0 $Y2=0
cc_335 N_A1_M1033_g N_VGND_c_2033_n 0.0154359f $X=0.925 $Y=0.95 $X2=0 $Y2=0
cc_336 A1 N_VGND_c_2033_n 0.0398625f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_337 N_A1_c_312_n N_VGND_c_2033_n 0.0055439f $X=0.955 $Y=1.615 $X2=0 $Y2=0
cc_338 N_A1_M1025_g N_VGND_c_2050_n 0.00354577f $X=0.495 $Y=0.95 $X2=0 $Y2=0
cc_339 N_A1_M1033_g N_VGND_c_2050_n 2.33667e-19 $X=0.925 $Y=0.95 $X2=0 $Y2=0
cc_340 N_A1_M1025_g N_VGND_c_2058_n 0.00391696f $X=0.495 $Y=0.95 $X2=0 $Y2=0
cc_341 N_A1_M1025_g N_A_114_126#_c_2232_n 0.00626483f $X=0.495 $Y=0.95 $X2=0
+ $Y2=0
cc_342 N_A1_M1033_g N_A_114_126#_c_2232_n 0.00727484f $X=0.925 $Y=0.95 $X2=0
+ $Y2=0
cc_343 N_A1_M1033_g N_A_114_126#_c_2233_n 0.00455657f $X=0.925 $Y=0.95 $X2=0
+ $Y2=0
cc_344 A0 N_S0_M1000_g 8.62325e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_345 N_A0_c_356_n N_S0_M1000_g 0.006695f $X=2.19 $Y=1.635 $X2=0 $Y2=0
cc_346 N_A0_M1007_g N_VPWR_c_1243_n 0.011811f $X=1.405 $Y=2.46 $X2=0 $Y2=0
cc_347 N_A0_M1011_g N_VPWR_c_1243_n 6.96611e-19 $X=1.905 $Y=2.46 $X2=0 $Y2=0
cc_348 N_A0_M1011_g N_VPWR_c_1244_n 0.00501904f $X=1.905 $Y=2.46 $X2=0 $Y2=0
cc_349 N_A0_M1007_g N_VPWR_c_1260_n 0.00460063f $X=1.405 $Y=2.46 $X2=0 $Y2=0
cc_350 N_A0_M1011_g N_VPWR_c_1260_n 0.005209f $X=1.905 $Y=2.46 $X2=0 $Y2=0
cc_351 N_A0_M1007_g N_VPWR_c_1240_n 0.00909043f $X=1.405 $Y=2.46 $X2=0 $Y2=0
cc_352 N_A0_M1011_g N_VPWR_c_1240_n 0.00541032f $X=1.905 $Y=2.46 $X2=0 $Y2=0
cc_353 N_A0_M1007_g N_A_119_392#_c_1423_n 9.63162e-19 $X=1.405 $Y=2.46 $X2=0
+ $Y2=0
cc_354 N_A0_M1007_g N_A_119_392#_c_1424_n 0.0165315f $X=1.405 $Y=2.46 $X2=0
+ $Y2=0
cc_355 N_A0_M1011_g N_A_119_392#_c_1424_n 0.0140119f $X=1.905 $Y=2.46 $X2=0
+ $Y2=0
cc_356 A0 N_A_119_392#_c_1424_n 0.0850177f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_357 N_A0_c_355_n N_A_119_392#_c_1424_n 0.00329647f $X=1.995 $Y=1.635 $X2=0
+ $Y2=0
cc_358 N_A0_c_356_n N_A_119_392#_c_1424_n 0.00792612f $X=2.19 $Y=1.635 $X2=0
+ $Y2=0
cc_359 N_A0_M1011_g N_A_119_392#_c_1425_n 0.0040545f $X=1.905 $Y=2.46 $X2=0
+ $Y2=0
cc_360 A0 N_A_119_392#_c_1425_n 0.00227977f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_361 A0 N_A_119_392#_c_1421_n 0.0151563f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_362 N_A0_c_356_n N_A_119_392#_c_1421_n 7.73608e-19 $X=2.19 $Y=1.635 $X2=0
+ $Y2=0
cc_363 N_A0_M1011_g N_A_299_392#_c_1483_n 0.0119395f $X=1.905 $Y=2.46 $X2=0
+ $Y2=0
cc_364 N_A0_M1011_g N_A_299_392#_c_1485_n 0.0129627f $X=1.905 $Y=2.46 $X2=0
+ $Y2=0
cc_365 N_A0_M1023_g N_A_509_392#_c_1518_n 0.00280676f $X=1.85 $Y=0.95 $X2=0
+ $Y2=0
cc_366 N_A0_M1022_g N_VGND_c_2034_n 0.00308767f $X=1.42 $Y=0.95 $X2=0 $Y2=0
cc_367 A0 N_VGND_c_2034_n 0.0228477f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_368 N_A0_c_355_n N_VGND_c_2034_n 8.05101e-19 $X=1.995 $Y=1.635 $X2=0 $Y2=0
cc_369 N_A0_M1022_g N_VGND_c_2072_n 0.00569723f $X=1.42 $Y=0.95 $X2=0 $Y2=0
cc_370 N_A0_M1023_g N_VGND_c_2072_n 5.68292e-19 $X=1.85 $Y=0.95 $X2=0 $Y2=0
cc_371 N_A0_M1023_g N_VGND_c_2050_n 0.00258164f $X=1.85 $Y=0.95 $X2=0 $Y2=0
cc_372 N_A0_M1023_g N_VGND_c_2058_n 0.00360493f $X=1.85 $Y=0.95 $X2=0 $Y2=0
cc_373 N_A0_M1022_g N_A_114_126#_c_2232_n 6.3983e-19 $X=1.42 $Y=0.95 $X2=0 $Y2=0
cc_374 N_A0_M1022_g N_A_114_126#_c_2233_n 0.00692429f $X=1.42 $Y=0.95 $X2=0
+ $Y2=0
cc_375 N_A0_M1022_g N_A_114_126#_c_2235_n 0.0029318f $X=1.42 $Y=0.95 $X2=0 $Y2=0
cc_376 N_A0_M1023_g N_A_114_126#_c_2235_n 0.0067325f $X=1.85 $Y=0.95 $X2=0 $Y2=0
cc_377 N_A0_M1022_g N_A_114_126#_c_2236_n 0.00180292f $X=1.42 $Y=0.95 $X2=0
+ $Y2=0
cc_378 N_A0_M1023_g N_A_114_126#_c_2236_n 0.0117504f $X=1.85 $Y=0.95 $X2=0 $Y2=0
cc_379 N_A0_M1023_g N_A_299_126#_c_2282_n 0.0106426f $X=1.85 $Y=0.95 $X2=0 $Y2=0
cc_380 A0 N_A_299_126#_c_2282_n 0.0412064f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_381 N_A0_c_355_n N_A_299_126#_c_2282_n 0.0098964f $X=1.995 $Y=1.635 $X2=0
+ $Y2=0
cc_382 N_A0_M1022_g N_A_299_126#_c_2285_n 5.84569e-19 $X=1.42 $Y=0.95 $X2=0
+ $Y2=0
cc_383 N_A0_M1023_g N_A_299_126#_c_2285_n 0.00900763f $X=1.85 $Y=0.95 $X2=0
+ $Y2=0
cc_384 A0 N_A_299_126#_c_2285_n 0.0196736f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_385 N_A0_c_355_n N_A_299_126#_c_2285_n 0.00228163f $X=1.995 $Y=1.635 $X2=0
+ $Y2=0
cc_386 N_A0_M1023_g N_A_299_126#_c_2286_n 0.00320159f $X=1.85 $Y=0.95 $X2=0
+ $Y2=0
cc_387 N_A_758_306#_c_414_n N_S0_M1042_g 0.0286939f $X=4.42 $Y=1.547 $X2=0 $Y2=0
cc_388 N_A_758_306#_M1039_g N_S0_M1047_g 0.0126979f $X=3.905 $Y=0.915 $X2=0
+ $Y2=0
cc_389 N_A_758_306#_M1039_g N_S0_c_552_n 0.00882199f $X=3.905 $Y=0.915 $X2=0
+ $Y2=0
cc_390 N_A_758_306#_M1043_g N_S0_c_552_n 0.00903828f $X=4.335 $Y=0.915 $X2=0
+ $Y2=0
cc_391 N_A_758_306#_c_417_n N_S0_c_552_n 0.00506365f $X=5.11 $Y=0.515 $X2=0
+ $Y2=0
cc_392 N_A_758_306#_c_417_n N_S0_M1016_g 0.0111534f $X=5.11 $Y=0.515 $X2=0 $Y2=0
cc_393 N_A_758_306#_c_429_n N_S0_M1013_g 0.00798142f $X=5.115 $Y=1.985 $X2=0
+ $Y2=0
cc_394 N_A_758_306#_c_418_n N_S0_M1013_g 8.06287e-19 $X=6.365 $Y=1.53 $X2=0
+ $Y2=0
cc_395 N_A_758_306#_c_419_n N_S0_M1013_g 0.0205612f $X=4.875 $Y=1.515 $X2=0
+ $Y2=0
cc_396 N_A_758_306#_c_420_n N_S0_M1013_g 0.0045242f $X=5.2 $Y=1.515 $X2=0 $Y2=0
cc_397 N_A_758_306#_c_421_n N_S0_M1013_g 0.0175612f $X=6.035 $Y=1.53 $X2=0 $Y2=0
cc_398 N_A_758_306#_c_423_n N_S0_M1013_g 0.00464349f $X=6.8 $Y=1.53 $X2=0 $Y2=0
cc_399 N_A_758_306#_c_415_n N_S0_c_556_n 0.00980793f $X=6.315 $Y=1.365 $X2=0
+ $Y2=0
cc_400 N_A_758_306#_c_416_n N_S0_c_556_n 0.00844637f $X=6.745 $Y=1.365 $X2=0
+ $Y2=0
cc_401 N_A_758_306#_c_416_n N_S0_M1012_g 0.0106844f $X=6.745 $Y=1.365 $X2=0
+ $Y2=0
cc_402 N_A_758_306#_c_423_n N_S0_M1012_g 0.011768f $X=6.8 $Y=1.53 $X2=0 $Y2=0
cc_403 N_A_758_306#_M1050_g N_S0_M1001_g 0.0160374f $X=6.8 $Y=2.385 $X2=0 $Y2=0
cc_404 N_A_758_306#_c_414_n N_S0_c_561_n 0.0126979f $X=4.42 $Y=1.547 $X2=0 $Y2=0
cc_405 N_A_758_306#_c_423_n N_S0_c_566_n 0.0160374f $X=6.8 $Y=1.53 $X2=0 $Y2=0
cc_406 N_A_758_306#_M1046_g N_VPWR_c_1245_n 0.00578993f $X=6.35 $Y=2.385 $X2=0
+ $Y2=0
cc_407 N_A_758_306#_c_429_n N_VPWR_c_1245_n 0.0408989f $X=5.115 $Y=1.985 $X2=0
+ $Y2=0
cc_408 N_A_758_306#_c_421_n N_VPWR_c_1245_n 0.0170561f $X=6.035 $Y=1.53 $X2=0
+ $Y2=0
cc_409 N_A_758_306#_M1045_g N_VPWR_c_1261_n 0.00333896f $X=3.88 $Y=2.46 $X2=0
+ $Y2=0
cc_410 N_A_758_306#_M1049_g N_VPWR_c_1261_n 0.00333882f $X=4.33 $Y=2.46 $X2=0
+ $Y2=0
cc_411 N_A_758_306#_c_429_n N_VPWR_c_1261_n 0.011066f $X=5.115 $Y=1.985 $X2=0
+ $Y2=0
cc_412 N_A_758_306#_M1046_g N_VPWR_c_1262_n 0.005403f $X=6.35 $Y=2.385 $X2=0
+ $Y2=0
cc_413 N_A_758_306#_M1050_g N_VPWR_c_1262_n 9.98368e-19 $X=6.8 $Y=2.385 $X2=0
+ $Y2=0
cc_414 N_A_758_306#_M1045_g N_VPWR_c_1240_n 0.00423029f $X=3.88 $Y=2.46 $X2=0
+ $Y2=0
cc_415 N_A_758_306#_M1049_g N_VPWR_c_1240_n 0.00427817f $X=4.33 $Y=2.46 $X2=0
+ $Y2=0
cc_416 N_A_758_306#_M1046_g N_VPWR_c_1240_n 0.0052212f $X=6.35 $Y=2.385 $X2=0
+ $Y2=0
cc_417 N_A_758_306#_c_429_n N_VPWR_c_1240_n 0.00915947f $X=5.115 $Y=1.985 $X2=0
+ $Y2=0
cc_418 N_A_758_306#_M1045_g N_A_119_392#_c_1420_n 0.0104102f $X=3.88 $Y=2.46
+ $X2=0 $Y2=0
cc_419 N_A_758_306#_M1049_g N_A_119_392#_c_1420_n 7.62301e-19 $X=4.33 $Y=2.46
+ $X2=0 $Y2=0
cc_420 N_A_758_306#_c_414_n N_A_119_392#_c_1420_n 0.0126969f $X=4.42 $Y=1.547
+ $X2=0 $Y2=0
cc_421 N_A_758_306#_M1045_g N_A_119_392#_c_1428_n 0.00453984f $X=3.88 $Y=2.46
+ $X2=0 $Y2=0
cc_422 N_A_758_306#_M1049_g N_A_119_392#_c_1428_n 0.00170793f $X=4.33 $Y=2.46
+ $X2=0 $Y2=0
cc_423 N_A_758_306#_M1045_g N_A_509_392#_c_1525_n 0.0132856f $X=3.88 $Y=2.46
+ $X2=0 $Y2=0
cc_424 N_A_758_306#_M1049_g N_A_509_392#_c_1525_n 6.80759e-19 $X=4.33 $Y=2.46
+ $X2=0 $Y2=0
cc_425 N_A_758_306#_M1039_g N_A_509_392#_c_1513_n 0.00203728f $X=3.905 $Y=0.915
+ $X2=0 $Y2=0
cc_426 N_A_758_306#_M1039_g N_A_509_392#_c_1514_n 0.00330666f $X=3.905 $Y=0.915
+ $X2=0 $Y2=0
cc_427 N_A_758_306#_M1043_g N_A_509_392#_c_1514_n 0.00283033f $X=4.335 $Y=0.915
+ $X2=0 $Y2=0
cc_428 N_A_758_306#_c_417_n N_A_509_392#_c_1514_n 0.00526842f $X=5.11 $Y=0.515
+ $X2=0 $Y2=0
cc_429 N_A_758_306#_M1045_g N_A_509_392#_c_1526_n 0.0116345f $X=3.88 $Y=2.46
+ $X2=0 $Y2=0
cc_430 N_A_758_306#_M1049_g N_A_509_392#_c_1526_n 0.0138856f $X=4.33 $Y=2.46
+ $X2=0 $Y2=0
cc_431 N_A_758_306#_c_429_n N_A_509_392#_c_1526_n 0.00526103f $X=5.115 $Y=1.985
+ $X2=0 $Y2=0
cc_432 N_A_758_306#_M1039_g N_A_509_392#_c_1515_n 7.22399e-19 $X=3.905 $Y=0.915
+ $X2=0 $Y2=0
cc_433 N_A_758_306#_M1043_g N_A_509_392#_c_1515_n 0.0098936f $X=4.335 $Y=0.915
+ $X2=0 $Y2=0
cc_434 N_A_758_306#_c_417_n N_A_509_392#_c_1515_n 0.0499741f $X=5.11 $Y=0.515
+ $X2=0 $Y2=0
cc_435 N_A_758_306#_M1049_g N_A_509_392#_c_1527_n 0.0114399f $X=4.33 $Y=2.46
+ $X2=0 $Y2=0
cc_436 N_A_758_306#_M1045_g N_A_509_392#_c_1529_n 0.0020162f $X=3.88 $Y=2.46
+ $X2=0 $Y2=0
cc_437 N_A_758_306#_M1043_g N_A_509_392#_c_1520_n 0.00183387f $X=4.335 $Y=0.915
+ $X2=0 $Y2=0
cc_438 N_A_758_306#_c_422_n N_A_509_392#_c_1520_n 0.00666801f $X=4.71 $Y=1.515
+ $X2=0 $Y2=0
cc_439 N_A_758_306#_M1013_s N_A_509_392#_c_1530_n 0.00365135f $X=4.97 $Y=1.84
+ $X2=0 $Y2=0
cc_440 N_A_758_306#_M1046_g N_A_509_392#_c_1530_n 0.00681486f $X=6.35 $Y=2.385
+ $X2=0 $Y2=0
cc_441 N_A_758_306#_M1050_g N_A_509_392#_c_1530_n 0.00681486f $X=6.8 $Y=2.385
+ $X2=0 $Y2=0
cc_442 N_A_758_306#_c_429_n N_A_509_392#_c_1530_n 0.0238995f $X=5.115 $Y=1.985
+ $X2=0 $Y2=0
cc_443 N_A_758_306#_c_418_n N_A_509_392#_c_1530_n 0.00395434f $X=6.365 $Y=1.53
+ $X2=0 $Y2=0
cc_444 N_A_758_306#_c_419_n N_A_509_392#_c_1530_n 0.00523275f $X=4.875 $Y=1.515
+ $X2=0 $Y2=0
cc_445 N_A_758_306#_c_420_n N_A_509_392#_c_1530_n 0.0100335f $X=5.2 $Y=1.515
+ $X2=0 $Y2=0
cc_446 N_A_758_306#_c_421_n N_A_509_392#_c_1530_n 0.0143559f $X=6.035 $Y=1.53
+ $X2=0 $Y2=0
cc_447 N_A_758_306#_c_429_n N_A_509_392#_c_1531_n 6.54704e-19 $X=5.115 $Y=1.985
+ $X2=0 $Y2=0
cc_448 N_A_758_306#_M1049_g N_A_509_392#_c_1532_n 0.0029499f $X=4.33 $Y=2.46
+ $X2=0 $Y2=0
cc_449 N_A_758_306#_c_429_n N_A_509_392#_c_1532_n 0.0626517f $X=5.115 $Y=1.985
+ $X2=0 $Y2=0
cc_450 N_A_758_306#_c_422_n N_A_509_392#_c_1532_n 0.00572494f $X=4.71 $Y=1.515
+ $X2=0 $Y2=0
cc_451 N_A_758_306#_M1045_g N_A_509_392#_c_1523_n 8.05383e-19 $X=3.88 $Y=2.46
+ $X2=0 $Y2=0
cc_452 N_A_758_306#_M1049_g N_A_509_392#_c_1523_n 0.00736331f $X=4.33 $Y=2.46
+ $X2=0 $Y2=0
cc_453 N_A_758_306#_M1043_g N_A_509_392#_c_1523_n 0.00492997f $X=4.335 $Y=0.915
+ $X2=0 $Y2=0
cc_454 N_A_758_306#_c_414_n N_A_509_392#_c_1523_n 0.0098422f $X=4.42 $Y=1.547
+ $X2=0 $Y2=0
cc_455 N_A_758_306#_c_417_n N_A_509_392#_c_1523_n 0.00515416f $X=5.11 $Y=0.515
+ $X2=0 $Y2=0
cc_456 N_A_758_306#_c_429_n N_A_509_392#_c_1523_n 0.00809031f $X=5.115 $Y=1.985
+ $X2=0 $Y2=0
cc_457 N_A_758_306#_c_419_n N_A_509_392#_c_1523_n 4.37509e-19 $X=4.875 $Y=1.515
+ $X2=0 $Y2=0
cc_458 N_A_758_306#_c_420_n N_A_509_392#_c_1523_n 0.0248912f $X=5.2 $Y=1.515
+ $X2=0 $Y2=0
cc_459 N_A_758_306#_c_422_n N_A_509_392#_c_1523_n 0.0126905f $X=4.71 $Y=1.515
+ $X2=0 $Y2=0
cc_460 N_A_758_306#_c_421_n N_A_1191_121#_c_1699_n 0.0208194f $X=6.035 $Y=1.53
+ $X2=0 $Y2=0
cc_461 N_A_758_306#_c_423_n N_A_1191_121#_c_1699_n 0.00347152f $X=6.8 $Y=1.53
+ $X2=0 $Y2=0
cc_462 N_A_758_306#_c_415_n N_A_1191_121#_c_1700_n 4.43891e-19 $X=6.315 $Y=1.365
+ $X2=0 $Y2=0
cc_463 N_A_758_306#_c_418_n N_A_1191_121#_c_1709_n 0.013784f $X=6.365 $Y=1.53
+ $X2=0 $Y2=0
cc_464 N_A_758_306#_c_421_n N_A_1191_121#_c_1709_n 0.00116029f $X=6.035 $Y=1.53
+ $X2=0 $Y2=0
cc_465 N_A_758_306#_c_423_n N_A_1191_121#_c_1709_n 0.00407674f $X=6.8 $Y=1.53
+ $X2=0 $Y2=0
cc_466 N_A_758_306#_M1046_g N_A_1191_121#_c_1710_n 0.00107927f $X=6.35 $Y=2.385
+ $X2=0 $Y2=0
cc_467 N_A_758_306#_c_415_n N_A_1191_121#_c_1727_n 0.0119972f $X=6.315 $Y=1.365
+ $X2=0 $Y2=0
cc_468 N_A_758_306#_c_416_n N_A_1191_121#_c_1727_n 0.0115176f $X=6.745 $Y=1.365
+ $X2=0 $Y2=0
cc_469 N_A_758_306#_c_418_n N_A_1191_121#_c_1727_n 0.0317383f $X=6.365 $Y=1.53
+ $X2=0 $Y2=0
cc_470 N_A_758_306#_c_423_n N_A_1191_121#_c_1727_n 0.00243905f $X=6.8 $Y=1.53
+ $X2=0 $Y2=0
cc_471 N_A_758_306#_M1046_g N_A_1191_121#_c_1711_n 0.0114106f $X=6.35 $Y=2.385
+ $X2=0 $Y2=0
cc_472 N_A_758_306#_M1050_g N_A_1191_121#_c_1711_n 0.0136866f $X=6.8 $Y=2.385
+ $X2=0 $Y2=0
cc_473 N_A_758_306#_c_418_n N_A_1191_121#_c_1711_n 0.0336884f $X=6.365 $Y=1.53
+ $X2=0 $Y2=0
cc_474 N_A_758_306#_c_423_n N_A_1191_121#_c_1711_n 0.00337308f $X=6.8 $Y=1.53
+ $X2=0 $Y2=0
cc_475 N_A_758_306#_c_416_n N_A_1191_121#_c_1702_n 0.00221303f $X=6.745 $Y=1.365
+ $X2=0 $Y2=0
cc_476 N_A_758_306#_c_524_p N_A_1191_121#_c_1702_n 0.0206343f $X=6.54 $Y=1.53
+ $X2=0 $Y2=0
cc_477 N_A_758_306#_c_423_n N_A_1191_121#_c_1702_n 0.00715517f $X=6.8 $Y=1.53
+ $X2=0 $Y2=0
cc_478 N_A_758_306#_c_416_n N_A_1191_121#_c_1707_n 4.93723e-19 $X=6.745 $Y=1.365
+ $X2=0 $Y2=0
cc_479 N_A_758_306#_c_423_n N_A_1191_121#_c_1707_n 5.44986e-19 $X=6.8 $Y=1.53
+ $X2=0 $Y2=0
cc_480 N_A_758_306#_M1046_g N_A_1288_377#_c_1875_n 0.00975814f $X=6.35 $Y=2.385
+ $X2=0 $Y2=0
cc_481 N_A_758_306#_M1050_g N_A_1288_377#_c_1875_n 0.0105237f $X=6.8 $Y=2.385
+ $X2=0 $Y2=0
cc_482 N_A_758_306#_M1050_g N_A_1288_377#_c_1871_n 0.0116285f $X=6.8 $Y=2.385
+ $X2=0 $Y2=0
cc_483 N_A_758_306#_M1046_g N_A_1288_377#_c_1872_n 0.00700898f $X=6.35 $Y=2.385
+ $X2=0 $Y2=0
cc_484 N_A_758_306#_M1050_g N_A_1288_377#_c_1872_n 0.00204203f $X=6.8 $Y=2.385
+ $X2=0 $Y2=0
cc_485 N_A_758_306#_c_415_n N_VGND_c_2036_n 0.00251838f $X=6.315 $Y=1.365 $X2=0
+ $Y2=0
cc_486 N_A_758_306#_c_417_n N_VGND_c_2036_n 0.0300842f $X=5.11 $Y=0.515 $X2=0
+ $Y2=0
cc_487 N_A_758_306#_c_421_n N_VGND_c_2036_n 0.0217489f $X=6.035 $Y=1.53 $X2=0
+ $Y2=0
cc_488 N_A_758_306#_c_417_n N_VGND_c_2051_n 0.0112807f $X=5.11 $Y=0.515 $X2=0
+ $Y2=0
cc_489 N_A_758_306#_c_415_n N_VGND_c_2058_n 7.88433e-19 $X=6.315 $Y=1.365 $X2=0
+ $Y2=0
cc_490 N_A_758_306#_c_417_n N_VGND_c_2058_n 0.0083297f $X=5.11 $Y=0.515 $X2=0
+ $Y2=0
cc_491 N_A_758_306#_M1039_g N_A_299_126#_c_2283_n 0.0108159f $X=3.905 $Y=0.915
+ $X2=0 $Y2=0
cc_492 N_A_758_306#_M1043_g N_A_299_126#_c_2283_n 0.00124776f $X=4.335 $Y=0.915
+ $X2=0 $Y2=0
cc_493 N_A_758_306#_c_414_n N_A_299_126#_c_2283_n 0.0103808f $X=4.42 $Y=1.547
+ $X2=0 $Y2=0
cc_494 N_A_758_306#_M1039_g N_A_299_126#_c_2284_n 0.00848904f $X=3.905 $Y=0.915
+ $X2=0 $Y2=0
cc_495 N_A_758_306#_c_415_n N_A_1278_121#_c_2324_n 0.00749799f $X=6.315 $Y=1.365
+ $X2=0 $Y2=0
cc_496 N_A_758_306#_c_416_n N_A_1278_121#_c_2324_n 0.00699059f $X=6.745 $Y=1.365
+ $X2=0 $Y2=0
cc_497 N_A_758_306#_c_416_n N_A_1278_121#_c_2325_n 0.00163034f $X=6.745 $Y=1.365
+ $X2=0 $Y2=0
cc_498 N_S0_c_564_n N_A2_M1036_g 0.00720075f $X=8.155 $Y=1.56 $X2=0 $Y2=0
cc_499 N_S0_c_556_n N_A2_M1021_g 0.016973f $X=8.155 $Y=0.18 $X2=0 $Y2=0
cc_500 N_S0_c_559_n A2 0.00102397f $X=8.23 $Y=1.395 $X2=0 $Y2=0
cc_501 N_S0_c_564_n A2 2.4966e-19 $X=8.155 $Y=1.56 $X2=0 $Y2=0
cc_502 S0 A2 0.0225759f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_503 N_S0_c_559_n N_A2_c_724_n 0.00720075f $X=8.23 $Y=1.395 $X2=0 $Y2=0
cc_504 S0 N_A2_c_724_n 0.00383373f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_505 N_S0_M1000_g N_VPWR_c_1244_n 0.00124669f $X=2.93 $Y=2.46 $X2=0 $Y2=0
cc_506 N_S0_M1013_g N_VPWR_c_1245_n 0.023878f $X=5.34 $Y=2.4 $X2=0 $Y2=0
cc_507 N_S0_M1000_g N_VPWR_c_1261_n 0.00335128f $X=2.93 $Y=2.46 $X2=0 $Y2=0
cc_508 N_S0_M1042_g N_VPWR_c_1261_n 0.00333921f $X=3.405 $Y=2.46 $X2=0 $Y2=0
cc_509 N_S0_M1013_g N_VPWR_c_1261_n 0.00460063f $X=5.34 $Y=2.4 $X2=0 $Y2=0
cc_510 N_S0_M1001_g N_VPWR_c_1262_n 9.79923e-19 $X=7.25 $Y=2.385 $X2=0 $Y2=0
cc_511 N_S0_M1008_g N_VPWR_c_1262_n 9.79923e-19 $X=7.7 $Y=2.385 $X2=0 $Y2=0
cc_512 N_S0_M1000_g N_VPWR_c_1240_n 0.0042716f $X=2.93 $Y=2.46 $X2=0 $Y2=0
cc_513 N_S0_M1042_g N_VPWR_c_1240_n 0.00423281f $X=3.405 $Y=2.46 $X2=0 $Y2=0
cc_514 N_S0_M1013_g N_VPWR_c_1240_n 0.00913687f $X=5.34 $Y=2.4 $X2=0 $Y2=0
cc_515 N_S0_M1000_g N_A_119_392#_c_1424_n 0.00397786f $X=2.93 $Y=2.46 $X2=0
+ $Y2=0
cc_516 N_S0_M1000_g N_A_119_392#_c_1425_n 0.00637317f $X=2.93 $Y=2.46 $X2=0
+ $Y2=0
cc_517 N_S0_M1000_g N_A_119_392#_c_1420_n 0.0141195f $X=2.93 $Y=2.46 $X2=0 $Y2=0
cc_518 N_S0_M1042_g N_A_119_392#_c_1420_n 0.0172461f $X=3.405 $Y=2.46 $X2=0
+ $Y2=0
cc_519 N_S0_c_560_n N_A_119_392#_c_1420_n 0.00150122f $X=2.957 $Y=1.46 $X2=0
+ $Y2=0
cc_520 N_S0_c_561_n N_A_119_392#_c_1420_n 0.00150122f $X=3.432 $Y=1.46 $X2=0
+ $Y2=0
cc_521 N_S0_M1000_g N_A_299_392#_c_1483_n 0.0134217f $X=2.93 $Y=2.46 $X2=0 $Y2=0
cc_522 N_S0_M1000_g N_A_299_392#_c_1484_n 0.0111107f $X=2.93 $Y=2.46 $X2=0 $Y2=0
cc_523 N_S0_M1042_g N_A_299_392#_c_1484_n 2.22854e-19 $X=3.405 $Y=2.46 $X2=0
+ $Y2=0
cc_524 N_S0_M1000_g N_A_299_392#_c_1491_n 0.00180857f $X=2.93 $Y=2.46 $X2=0
+ $Y2=0
cc_525 N_S0_M1000_g N_A_509_392#_c_1524_n 0.00957763f $X=2.93 $Y=2.46 $X2=0
+ $Y2=0
cc_526 N_S0_M1042_g N_A_509_392#_c_1524_n 0.0134135f $X=3.405 $Y=2.46 $X2=0
+ $Y2=0
cc_527 N_S0_M1009_g N_A_509_392#_c_1512_n 0.0125911f $X=3 $Y=0.915 $X2=0 $Y2=0
cc_528 N_S0_c_548_n N_A_509_392#_c_1512_n 0.0034051f $X=3.4 $Y=0.18 $X2=0 $Y2=0
cc_529 N_S0_M1047_g N_A_509_392#_c_1512_n 0.0165579f $X=3.475 $Y=0.915 $X2=0
+ $Y2=0
cc_530 N_S0_M1000_g N_A_509_392#_c_1525_n 6.74956e-19 $X=2.93 $Y=2.46 $X2=0
+ $Y2=0
cc_531 N_S0_M1042_g N_A_509_392#_c_1525_n 0.0112244f $X=3.405 $Y=2.46 $X2=0
+ $Y2=0
cc_532 N_S0_M1047_g N_A_509_392#_c_1513_n 0.00505756f $X=3.475 $Y=0.915 $X2=0
+ $Y2=0
cc_533 N_S0_c_552_n N_A_509_392#_c_1514_n 0.01748f $X=5.25 $Y=0.18 $X2=0 $Y2=0
cc_534 N_S0_M1016_g N_A_509_392#_c_1514_n 0.00174103f $X=5.325 $Y=0.74 $X2=0
+ $Y2=0
cc_535 N_S0_M1013_g N_A_509_392#_c_1526_n 0.00288376f $X=5.34 $Y=2.4 $X2=0 $Y2=0
cc_536 N_S0_M1000_g N_A_509_392#_c_1528_n 0.00771733f $X=2.93 $Y=2.46 $X2=0
+ $Y2=0
cc_537 N_S0_M1042_g N_A_509_392#_c_1528_n 5.35884e-19 $X=3.405 $Y=2.46 $X2=0
+ $Y2=0
cc_538 N_S0_M1009_g N_A_509_392#_c_1518_n 0.009152f $X=3 $Y=0.915 $X2=0 $Y2=0
cc_539 N_S0_M1042_g N_A_509_392#_c_1529_n 0.0014927f $X=3.405 $Y=2.46 $X2=0
+ $Y2=0
cc_540 N_S0_c_552_n N_A_509_392#_c_1519_n 0.00470837f $X=5.25 $Y=0.18 $X2=0
+ $Y2=0
cc_541 N_S0_M1013_g N_A_509_392#_c_1530_n 0.0080131f $X=5.34 $Y=2.4 $X2=0 $Y2=0
cc_542 S0 N_A_509_392#_c_1530_n 0.00940257f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_543 N_S0_M1016_g N_A_1191_121#_c_1699_n 0.00179375f $X=5.325 $Y=0.74 $X2=0
+ $Y2=0
cc_544 N_S0_c_554_n N_A_1191_121#_c_1699_n 2.94405e-19 $X=5.34 $Y=1.275 $X2=0
+ $Y2=0
cc_545 N_S0_M1016_g N_A_1191_121#_c_1700_n 8.46248e-19 $X=5.325 $Y=0.74 $X2=0
+ $Y2=0
cc_546 N_S0_c_556_n N_A_1191_121#_c_1700_n 0.00494503f $X=8.155 $Y=0.18 $X2=0
+ $Y2=0
cc_547 N_S0_M1013_g N_A_1191_121#_c_1710_n 0.00148983f $X=5.34 $Y=2.4 $X2=0
+ $Y2=0
cc_548 N_S0_M1012_g N_A_1191_121#_c_1701_n 6.552e-19 $X=7.175 $Y=0.925 $X2=0
+ $Y2=0
cc_549 N_S0_M1012_g N_A_1191_121#_c_1746_n 0.00407014f $X=7.175 $Y=0.925 $X2=0
+ $Y2=0
cc_550 N_S0_M1041_g N_A_1191_121#_c_1746_n 4.70674e-19 $X=7.605 $Y=0.925 $X2=0
+ $Y2=0
cc_551 N_S0_M1012_g N_A_1191_121#_c_1702_n 0.00313646f $X=7.175 $Y=0.925 $X2=0
+ $Y2=0
cc_552 N_S0_M1041_g N_A_1191_121#_c_1702_n 6.31438e-19 $X=7.605 $Y=0.925 $X2=0
+ $Y2=0
cc_553 S0 N_A_1191_121#_c_1702_n 0.0267198f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_554 N_S0_c_566_n N_A_1191_121#_c_1702_n 0.00937479f $X=7.79 $Y=1.56 $X2=0
+ $Y2=0
cc_555 N_S0_M1012_g N_A_1191_121#_c_1703_n 0.0103465f $X=7.175 $Y=0.925 $X2=0
+ $Y2=0
cc_556 N_S0_M1041_g N_A_1191_121#_c_1703_n 0.00968335f $X=7.605 $Y=0.925 $X2=0
+ $Y2=0
cc_557 N_S0_M1001_g N_A_1191_121#_c_1713_n 0.0183488f $X=7.25 $Y=2.385 $X2=0
+ $Y2=0
cc_558 N_S0_M1008_g N_A_1191_121#_c_1713_n 0.00964311f $X=7.7 $Y=2.385 $X2=0
+ $Y2=0
cc_559 N_S0_c_564_n N_A_1191_121#_c_1713_n 0.0030281f $X=8.155 $Y=1.56 $X2=0
+ $Y2=0
cc_560 S0 N_A_1191_121#_c_1713_n 0.0791022f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_561 N_S0_c_566_n N_A_1191_121#_c_1713_n 5.47363e-19 $X=7.79 $Y=1.56 $X2=0
+ $Y2=0
cc_562 N_S0_M1012_g N_A_1191_121#_c_1707_n 0.00265737f $X=7.175 $Y=0.925 $X2=0
+ $Y2=0
cc_563 N_S0_M1001_g N_A_1191_121#_c_1718_n 6.21494e-19 $X=7.25 $Y=2.385 $X2=0
+ $Y2=0
cc_564 N_S0_M1041_g N_A_1191_121#_c_1708_n 5.15987e-19 $X=7.605 $Y=0.925 $X2=0
+ $Y2=0
cc_565 N_S0_c_559_n N_A_1191_121#_c_1708_n 0.00476489f $X=8.23 $Y=1.395 $X2=0
+ $Y2=0
cc_566 N_S0_M1001_g N_A_1288_377#_c_1875_n 9.10491e-19 $X=7.25 $Y=2.385 $X2=0
+ $Y2=0
cc_567 N_S0_M1001_g N_A_1288_377#_c_1871_n 0.01414f $X=7.25 $Y=2.385 $X2=0 $Y2=0
cc_568 N_S0_M1008_g N_A_1288_377#_c_1871_n 0.0117384f $X=7.7 $Y=2.385 $X2=0
+ $Y2=0
cc_569 N_S0_M1008_g N_A_1288_377#_c_1874_n 0.0086845f $X=7.7 $Y=2.385 $X2=0
+ $Y2=0
cc_570 N_S0_M1008_g N_A_1468_377#_c_1926_n 0.0128978f $X=7.7 $Y=2.385 $X2=0
+ $Y2=0
cc_571 N_S0_M1001_g N_A_1468_377#_c_1928_n 0.00678324f $X=7.25 $Y=2.385 $X2=0
+ $Y2=0
cc_572 N_S0_M1008_g N_A_1468_377#_c_1928_n 0.0118885f $X=7.7 $Y=2.385 $X2=0
+ $Y2=0
cc_573 N_S0_c_549_n N_VGND_c_2035_n 0.00227104f $X=3.075 $Y=0.18 $X2=0 $Y2=0
cc_574 N_S0_M1016_g N_VGND_c_2036_n 0.0147983f $X=5.325 $Y=0.74 $X2=0 $Y2=0
cc_575 N_S0_c_554_n N_VGND_c_2036_n 9.78193e-19 $X=5.34 $Y=1.275 $X2=0 $Y2=0
cc_576 N_S0_c_556_n N_VGND_c_2036_n 0.0187754f $X=8.155 $Y=0.18 $X2=0 $Y2=0
cc_577 N_S0_c_563_n N_VGND_c_2036_n 0.00460513f $X=5.325 $Y=0.18 $X2=0 $Y2=0
cc_578 N_S0_c_556_n N_VGND_c_2044_n 0.00443934f $X=8.155 $Y=0.18 $X2=0 $Y2=0
cc_579 N_S0_c_559_n N_VGND_c_2044_n 6.29386e-19 $X=8.23 $Y=1.395 $X2=0 $Y2=0
cc_580 N_S0_c_556_n N_VGND_c_2045_n 0.0604235f $X=8.155 $Y=0.18 $X2=0 $Y2=0
cc_581 N_S0_c_549_n N_VGND_c_2051_n 0.0586296f $X=3.075 $Y=0.18 $X2=0 $Y2=0
cc_582 N_S0_c_548_n N_VGND_c_2058_n 0.00777952f $X=3.4 $Y=0.18 $X2=0 $Y2=0
cc_583 N_S0_c_549_n N_VGND_c_2058_n 0.00604517f $X=3.075 $Y=0.18 $X2=0 $Y2=0
cc_584 N_S0_c_552_n N_VGND_c_2058_n 0.0489771f $X=5.25 $Y=0.18 $X2=0 $Y2=0
cc_585 N_S0_c_556_n N_VGND_c_2058_n 0.0737993f $X=8.155 $Y=0.18 $X2=0 $Y2=0
cc_586 N_S0_c_562_n N_VGND_c_2058_n 0.00370846f $X=3.475 $Y=0.18 $X2=0 $Y2=0
cc_587 N_S0_c_563_n N_VGND_c_2058_n 0.00749832f $X=5.325 $Y=0.18 $X2=0 $Y2=0
cc_588 N_S0_M1009_g N_A_114_126#_c_2247_n 0.0155442f $X=3 $Y=0.915 $X2=0 $Y2=0
cc_589 N_S0_c_561_n N_A_114_126#_c_2247_n 3.36668e-19 $X=3.432 $Y=1.46 $X2=0
+ $Y2=0
cc_590 N_S0_M1009_g N_A_114_126#_c_2237_n 0.00991756f $X=3 $Y=0.915 $X2=0 $Y2=0
cc_591 N_S0_c_560_n N_A_114_126#_c_2237_n 3.2644e-19 $X=2.957 $Y=1.46 $X2=0
+ $Y2=0
cc_592 N_S0_M1009_g N_A_299_126#_c_2283_n 0.00490473f $X=3 $Y=0.915 $X2=0 $Y2=0
cc_593 N_S0_M1047_g N_A_299_126#_c_2283_n 0.00850432f $X=3.475 $Y=0.915 $X2=0
+ $Y2=0
cc_594 N_S0_c_560_n N_A_299_126#_c_2283_n 0.00997967f $X=2.957 $Y=1.46 $X2=0
+ $Y2=0
cc_595 N_S0_c_561_n N_A_299_126#_c_2283_n 0.00925259f $X=3.432 $Y=1.46 $X2=0
+ $Y2=0
cc_596 N_S0_M1047_g N_A_299_126#_c_2284_n 9.78227e-19 $X=3.475 $Y=0.915 $X2=0
+ $Y2=0
cc_597 N_S0_M1009_g N_A_299_126#_c_2286_n 0.00440371f $X=3 $Y=0.915 $X2=0 $Y2=0
cc_598 N_S0_c_560_n N_A_299_126#_c_2286_n 6.41487e-19 $X=2.957 $Y=1.46 $X2=0
+ $Y2=0
cc_599 N_S0_M1012_g N_A_1278_121#_c_2324_n 6.67018e-19 $X=7.175 $Y=0.925 $X2=0
+ $Y2=0
cc_600 N_S0_c_556_n N_A_1278_121#_c_2325_n 0.0264241f $X=8.155 $Y=0.18 $X2=0
+ $Y2=0
cc_601 N_S0_M1012_g N_A_1278_121#_c_2325_n 0.00115636f $X=7.175 $Y=0.925 $X2=0
+ $Y2=0
cc_602 N_S0_M1041_g N_A_1278_121#_c_2325_n 0.00115673f $X=7.605 $Y=0.925 $X2=0
+ $Y2=0
cc_603 N_S0_c_559_n N_A_1278_121#_c_2325_n 0.00580058f $X=8.23 $Y=1.395 $X2=0
+ $Y2=0
cc_604 N_S0_c_556_n N_A_1278_121#_c_2326_n 0.00727301f $X=8.155 $Y=0.18 $X2=0
+ $Y2=0
cc_605 N_S0_M1041_g N_A_1278_121#_c_2327_n 5.73967e-19 $X=7.605 $Y=0.925 $X2=0
+ $Y2=0
cc_606 N_S0_c_559_n N_A_1278_121#_c_2327_n 0.0068488f $X=8.23 $Y=1.395 $X2=0
+ $Y2=0
cc_607 N_S0_c_559_n N_A_1278_121#_c_2329_n 0.00783294f $X=8.23 $Y=1.395 $X2=0
+ $Y2=0
cc_608 N_S0_M1041_g N_A_1450_121#_c_2377_n 0.00950725f $X=7.605 $Y=0.925 $X2=0
+ $Y2=0
cc_609 N_S0_c_559_n N_A_1450_121#_c_2377_n 0.0012418f $X=8.23 $Y=1.395 $X2=0
+ $Y2=0
cc_610 S0 N_A_1450_121#_c_2377_n 0.0446554f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_611 N_S0_c_566_n N_A_1450_121#_c_2377_n 0.00699396f $X=7.79 $Y=1.56 $X2=0
+ $Y2=0
cc_612 N_S0_c_559_n N_A_1450_121#_c_2378_n 0.0010042f $X=8.23 $Y=1.395 $X2=0
+ $Y2=0
cc_613 S0 N_A_1450_121#_c_2378_n 0.00925546f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_614 N_S0_M1041_g N_A_1450_121#_c_2380_n 0.00485385f $X=7.605 $Y=0.925 $X2=0
+ $Y2=0
cc_615 N_S0_c_559_n N_A_1450_121#_c_2380_n 5.67881e-19 $X=8.23 $Y=1.395 $X2=0
+ $Y2=0
cc_616 S0 N_A_1450_121#_c_2380_n 0.0196697f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_617 N_S0_c_566_n N_A_1450_121#_c_2380_n 0.00276176f $X=7.79 $Y=1.56 $X2=0
+ $Y2=0
cc_618 N_S0_M1041_g N_A_1450_121#_c_2381_n 7.7137e-19 $X=7.605 $Y=0.925 $X2=0
+ $Y2=0
cc_619 N_S0_c_559_n N_A_1450_121#_c_2381_n 0.0153513f $X=8.23 $Y=1.395 $X2=0
+ $Y2=0
cc_620 S0 N_A_1450_121#_c_2381_n 0.0129022f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_621 N_A2_M1040_g N_A3_M1018_g 0.0219085f $X=9.385 $Y=0.69 $X2=0 $Y2=0
cc_622 A2 N_A3_M1018_g 0.00454402f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_623 N_A2_M1038_g N_A3_M1005_g 0.0356084f $X=9.245 $Y=2.46 $X2=0 $Y2=0
cc_624 N_A2_M1038_g A3 6.45648e-19 $X=9.245 $Y=2.46 $X2=0 $Y2=0
cc_625 A2 A3 0.0235668f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_626 N_A2_c_724_n A3 6.12354e-19 $X=9.385 $Y=1.425 $X2=0 $Y2=0
cc_627 N_A2_M1038_g N_A3_c_783_n 0.00506598f $X=9.245 $Y=2.46 $X2=0 $Y2=0
cc_628 A2 N_A3_c_783_n 0.00144227f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_629 N_A2_c_724_n N_A3_c_783_n 0.0219085f $X=9.385 $Y=1.425 $X2=0 $Y2=0
cc_630 N_A2_M1038_g N_VPWR_c_1251_n 0.00367331f $X=9.245 $Y=2.46 $X2=0 $Y2=0
cc_631 N_A2_M1036_g N_VPWR_c_1252_n 0.00377953f $X=8.795 $Y=2.46 $X2=0 $Y2=0
cc_632 N_A2_M1038_g N_VPWR_c_1252_n 0.00377953f $X=9.245 $Y=2.46 $X2=0 $Y2=0
cc_633 N_A2_M1036_g N_VPWR_c_1267_n 0.00531893f $X=8.795 $Y=2.46 $X2=0 $Y2=0
cc_634 N_A2_M1036_g N_VPWR_c_1240_n 0.0047145f $X=8.795 $Y=2.46 $X2=0 $Y2=0
cc_635 N_A2_M1038_g N_VPWR_c_1240_n 0.00467891f $X=9.245 $Y=2.46 $X2=0 $Y2=0
cc_636 A2 N_A_509_392#_c_1530_n 0.00557945f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_637 N_A2_M1036_g N_A_1191_121#_c_1713_n 0.0156191f $X=8.795 $Y=2.46 $X2=0
+ $Y2=0
cc_638 N_A2_M1038_g N_A_1191_121#_c_1713_n 0.0142026f $X=9.245 $Y=2.46 $X2=0
+ $Y2=0
cc_639 A2 N_A_1191_121#_c_1713_n 0.0504049f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_640 N_A2_c_724_n N_A_1191_121#_c_1713_n 9.6499e-19 $X=9.385 $Y=1.425 $X2=0
+ $Y2=0
cc_641 N_A2_M1036_g N_A_1288_377#_c_1873_n 0.0143319f $X=8.795 $Y=2.46 $X2=0
+ $Y2=0
cc_642 N_A2_M1038_g N_A_1288_377#_c_1873_n 0.0156433f $X=9.245 $Y=2.46 $X2=0
+ $Y2=0
cc_643 N_A2_M1038_g N_A_1288_377#_c_1886_n 0.00149905f $X=9.245 $Y=2.46 $X2=0
+ $Y2=0
cc_644 N_A2_M1036_g N_A_1288_377#_c_1874_n 0.00447523f $X=8.795 $Y=2.46 $X2=0
+ $Y2=0
cc_645 N_A2_M1036_g N_A_1468_377#_c_1926_n 0.0117087f $X=8.795 $Y=2.46 $X2=0
+ $Y2=0
cc_646 N_A2_M1038_g N_A_1468_377#_c_1926_n 0.00474014f $X=9.245 $Y=2.46 $X2=0
+ $Y2=0
cc_647 N_A2_M1021_g N_VGND_c_2037_n 4.68597e-19 $X=8.955 $Y=0.69 $X2=0 $Y2=0
cc_648 N_A2_M1040_g N_VGND_c_2037_n 0.00822569f $X=9.385 $Y=0.69 $X2=0 $Y2=0
cc_649 N_A2_M1021_g N_VGND_c_2044_n 0.00240369f $X=8.955 $Y=0.69 $X2=0 $Y2=0
cc_650 N_A2_M1021_g N_VGND_c_2046_n 0.00316493f $X=8.955 $Y=0.69 $X2=0 $Y2=0
cc_651 N_A2_M1040_g N_VGND_c_2046_n 0.00383152f $X=9.385 $Y=0.69 $X2=0 $Y2=0
cc_652 N_A2_M1021_g N_VGND_c_2058_n 0.00394055f $X=8.955 $Y=0.69 $X2=0 $Y2=0
cc_653 N_A2_M1040_g N_VGND_c_2058_n 0.0075754f $X=9.385 $Y=0.69 $X2=0 $Y2=0
cc_654 N_A2_M1021_g N_A_1278_121#_c_2325_n 5.24269e-19 $X=8.955 $Y=0.69 $X2=0
+ $Y2=0
cc_655 N_A2_M1021_g N_A_1278_121#_c_2327_n 0.00226665f $X=8.955 $Y=0.69 $X2=0
+ $Y2=0
cc_656 N_A2_M1021_g N_A_1278_121#_c_2328_n 0.00981813f $X=8.955 $Y=0.69 $X2=0
+ $Y2=0
cc_657 N_A2_M1021_g N_A_1278_121#_c_2330_n 0.00953282f $X=8.955 $Y=0.69 $X2=0
+ $Y2=0
cc_658 N_A2_M1021_g N_A_1450_121#_c_2378_n 0.0115689f $X=8.955 $Y=0.69 $X2=0
+ $Y2=0
cc_659 N_A2_M1040_g N_A_1450_121#_c_2378_n 0.0142932f $X=9.385 $Y=0.69 $X2=0
+ $Y2=0
cc_660 A2 N_A_1450_121#_c_2378_n 0.054183f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_661 N_A2_c_724_n N_A_1450_121#_c_2378_n 0.00815787f $X=9.385 $Y=1.425 $X2=0
+ $Y2=0
cc_662 N_A2_M1040_g N_A_1450_121#_c_2379_n 9.61031e-19 $X=9.385 $Y=0.69 $X2=0
+ $Y2=0
cc_663 N_A2_M1021_g N_A_1450_121#_c_2381_n 0.00262376f $X=8.955 $Y=0.69 $X2=0
+ $Y2=0
cc_664 N_A3_M1024_g N_VPWR_c_1246_n 0.00481605f $X=10.325 $Y=2.46 $X2=0 $Y2=0
cc_665 N_A3_M1005_g N_VPWR_c_1251_n 0.00338518f $X=9.875 $Y=2.46 $X2=0 $Y2=0
cc_666 N_A3_M1005_g N_VPWR_c_1253_n 0.00373263f $X=9.875 $Y=2.46 $X2=0 $Y2=0
cc_667 N_A3_M1024_g N_VPWR_c_1253_n 0.00519767f $X=10.325 $Y=2.46 $X2=0 $Y2=0
cc_668 N_A3_M1005_g N_VPWR_c_1240_n 0.00461573f $X=9.875 $Y=2.46 $X2=0 $Y2=0
cc_669 N_A3_M1024_g N_VPWR_c_1240_n 0.0098373f $X=10.325 $Y=2.46 $X2=0 $Y2=0
cc_670 A3 N_A_509_392#_c_1530_n 0.00519452f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_671 N_A3_M1005_g N_A_1191_121#_c_1713_n 0.0141877f $X=9.875 $Y=2.46 $X2=0
+ $Y2=0
cc_672 N_A3_M1024_g N_A_1191_121#_c_1713_n 0.018194f $X=10.325 $Y=2.46 $X2=0
+ $Y2=0
cc_673 A3 N_A_1191_121#_c_1713_n 0.0472952f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_674 N_A3_c_783_n N_A_1191_121#_c_1713_n 0.00320407f $X=10.325 $Y=1.61 $X2=0
+ $Y2=0
cc_675 N_A3_c_779_n N_A_1191_121#_c_1704_n 0.00188304f $X=10.245 $Y=1.085 $X2=0
+ $Y2=0
cc_676 N_A3_c_781_n N_A_1191_121#_c_1704_n 0.0108756f $X=10.335 $Y=1.16 $X2=0
+ $Y2=0
cc_677 A3 N_A_1191_121#_c_1704_n 0.0196213f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_678 N_A3_c_783_n N_A_1191_121#_c_1704_n 0.00714223f $X=10.325 $Y=1.61 $X2=0
+ $Y2=0
cc_679 N_A3_M1024_g N_A_1191_121#_c_1715_n 0.00516999f $X=10.325 $Y=2.46 $X2=0
+ $Y2=0
cc_680 N_A3_c_779_n N_A_1191_121#_c_1705_n 6.63977e-19 $X=10.245 $Y=1.085 $X2=0
+ $Y2=0
cc_681 N_A3_M1005_g N_A_1288_377#_c_1873_n 0.0163434f $X=9.875 $Y=2.46 $X2=0
+ $Y2=0
cc_682 N_A3_M1024_g N_A_1288_377#_c_1873_n 0.00492236f $X=10.325 $Y=2.46 $X2=0
+ $Y2=0
cc_683 N_A3_M1005_g N_A_1288_377#_c_1886_n 0.00778425f $X=9.875 $Y=2.46 $X2=0
+ $Y2=0
cc_684 N_A3_M1024_g N_A_1288_377#_c_1886_n 0.00463641f $X=10.325 $Y=2.46 $X2=0
+ $Y2=0
cc_685 N_A3_M1005_g N_A_1468_377#_c_1926_n 7.36526e-19 $X=9.875 $Y=2.46 $X2=0
+ $Y2=0
cc_686 N_A3_M1018_g N_VGND_c_2037_n 0.00160688f $X=9.815 $Y=0.69 $X2=0 $Y2=0
cc_687 N_A3_M1018_g N_VGND_c_2038_n 0.00434272f $X=9.815 $Y=0.69 $X2=0 $Y2=0
cc_688 N_A3_c_779_n N_VGND_c_2038_n 0.00383152f $X=10.245 $Y=1.085 $X2=0 $Y2=0
cc_689 N_A3_M1018_g N_VGND_c_2039_n 5.59381e-19 $X=9.815 $Y=0.69 $X2=0 $Y2=0
cc_690 N_A3_c_779_n N_VGND_c_2039_n 0.0129152f $X=10.245 $Y=1.085 $X2=0 $Y2=0
cc_691 N_A3_c_781_n N_VGND_c_2039_n 0.00323003f $X=10.335 $Y=1.16 $X2=0 $Y2=0
cc_692 A3 N_VGND_c_2039_n 0.00601406f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_693 N_A3_M1018_g N_VGND_c_2058_n 0.00820382f $X=9.815 $Y=0.69 $X2=0 $Y2=0
cc_694 N_A3_c_779_n N_VGND_c_2058_n 0.0075754f $X=10.245 $Y=1.085 $X2=0 $Y2=0
cc_695 N_A3_M1018_g N_A_1450_121#_c_2378_n 0.0135496f $X=9.815 $Y=0.69 $X2=0
+ $Y2=0
cc_696 N_A3_c_779_n N_A_1450_121#_c_2378_n 0.00109283f $X=10.245 $Y=1.085 $X2=0
+ $Y2=0
cc_697 A3 N_A_1450_121#_c_2378_n 0.0177215f $X=10.235 $Y=1.58 $X2=0 $Y2=0
cc_698 N_A3_c_783_n N_A_1450_121#_c_2378_n 0.00305517f $X=10.325 $Y=1.61 $X2=0
+ $Y2=0
cc_699 N_A3_M1018_g N_A_1450_121#_c_2379_n 0.00754481f $X=9.815 $Y=0.69 $X2=0
+ $Y2=0
cc_700 N_S1_M1019_g N_A_2489_347#_M1015_g 0.00828914f $X=11.945 $Y=0.69 $X2=0
+ $Y2=0
cc_701 N_S1_c_842_n N_A_2489_347#_M1015_g 0.00441765f $X=13.54 $Y=1.215 $X2=0
+ $Y2=0
cc_702 N_S1_c_843_n N_A_2489_347#_M1015_g 0.0182158f $X=12.315 $Y=1.36 $X2=0
+ $Y2=0
cc_703 N_S1_c_846_n N_A_2489_347#_M1015_g 0.0109898f $X=12.835 $Y=1.455 $X2=0
+ $Y2=0
cc_704 N_S1_c_842_n N_A_2489_347#_M1048_g 0.01631f $X=13.54 $Y=1.215 $X2=0 $Y2=0
cc_705 N_S1_c_844_n N_A_2489_347#_M1048_g 0.0145818f $X=13.87 $Y=1.385 $X2=0
+ $Y2=0
cc_706 N_S1_c_846_n N_A_2489_347#_M1048_g 9.7513e-19 $X=12.835 $Y=1.455 $X2=0
+ $Y2=0
cc_707 N_S1_c_842_n N_A_2489_347#_c_957_n 0.0333171f $X=13.54 $Y=1.215 $X2=0
+ $Y2=0
cc_708 N_S1_c_844_n N_A_2489_347#_c_957_n 0.00250238f $X=13.87 $Y=1.385 $X2=0
+ $Y2=0
cc_709 N_S1_M1044_g N_A_2489_347#_c_958_n 0.00154565f $X=14.3 $Y=2.4 $X2=0 $Y2=0
cc_710 N_S1_c_837_n N_A_2489_347#_c_951_n 0.0209844f $X=14.21 $Y=1.37 $X2=0
+ $Y2=0
cc_711 N_S1_c_838_n N_A_2489_347#_c_951_n 0.00537771f $X=14.285 $Y=1.22 $X2=0
+ $Y2=0
cc_712 N_S1_M1044_g N_A_2489_347#_c_951_n 0.00634256f $X=14.3 $Y=2.4 $X2=0 $Y2=0
cc_713 N_S1_c_842_n N_A_2489_347#_c_951_n 0.0307762f $X=13.54 $Y=1.215 $X2=0
+ $Y2=0
cc_714 N_S1_c_844_n N_A_2489_347#_c_951_n 2.10237e-19 $X=13.87 $Y=1.385 $X2=0
+ $Y2=0
cc_715 N_S1_c_842_n N_A_2489_347#_c_952_n 0.0293493f $X=13.54 $Y=1.215 $X2=0
+ $Y2=0
cc_716 N_S1_c_844_n N_A_2489_347#_c_952_n 3.06382e-19 $X=13.87 $Y=1.385 $X2=0
+ $Y2=0
cc_717 N_S1_c_846_n N_A_2489_347#_c_952_n 0.0246532f $X=12.835 $Y=1.455 $X2=0
+ $Y2=0
cc_718 N_S1_M1037_g N_A_2489_347#_c_953_n 0.0267476f $X=12.035 $Y=2.46 $X2=0
+ $Y2=0
cc_719 N_S1_c_842_n N_A_2489_347#_c_953_n 0.00280142f $X=13.54 $Y=1.215 $X2=0
+ $Y2=0
cc_720 N_S1_c_843_n N_A_2489_347#_c_953_n 0.00228017f $X=12.315 $Y=1.36 $X2=0
+ $Y2=0
cc_721 N_S1_c_844_n N_A_2489_347#_c_953_n 0.00530331f $X=13.87 $Y=1.385 $X2=0
+ $Y2=0
cc_722 N_S1_c_845_n N_A_2489_347#_c_953_n 0.00977718f $X=12.665 $Y=1.455 $X2=0
+ $Y2=0
cc_723 N_S1_c_846_n N_A_2489_347#_c_953_n 0.0161033f $X=12.835 $Y=1.455 $X2=0
+ $Y2=0
cc_724 N_S1_c_837_n N_A_2489_347#_c_962_n 0.00681687f $X=14.21 $Y=1.37 $X2=0
+ $Y2=0
cc_725 N_S1_M1044_g N_A_2489_347#_c_962_n 0.00520612f $X=14.3 $Y=2.4 $X2=0 $Y2=0
cc_726 N_S1_c_837_n N_A_2489_347#_c_954_n 0.00474764f $X=14.21 $Y=1.37 $X2=0
+ $Y2=0
cc_727 N_S1_M1044_g N_A_2199_74#_M1010_g 0.00956567f $X=14.3 $Y=2.4 $X2=0 $Y2=0
cc_728 N_S1_c_838_n N_A_2199_74#_M1020_g 0.00759404f $X=14.285 $Y=1.22 $X2=0
+ $Y2=0
cc_729 N_S1_c_841_n N_A_2199_74#_M1020_g 0.00421747f $X=14.3 $Y=1.37 $X2=0 $Y2=0
cc_730 N_S1_M1017_g N_A_2199_74#_c_1042_n 0.00631046f $X=11.355 $Y=0.69 $X2=0
+ $Y2=0
cc_731 N_S1_M1032_g N_A_2199_74#_c_1042_n 0.0239305f $X=11.535 $Y=2.46 $X2=0
+ $Y2=0
cc_732 N_S1_M1037_g N_A_2199_74#_c_1042_n 9.25587e-19 $X=12.035 $Y=2.46 $X2=0
+ $Y2=0
cc_733 N_S1_c_840_n N_A_2199_74#_c_1042_n 0.0182011f $X=12.125 $Y=1.36 $X2=0
+ $Y2=0
cc_734 N_S1_M1032_g N_A_2199_74#_c_1071_n 0.00976504f $X=11.535 $Y=2.46 $X2=0
+ $Y2=0
cc_735 N_S1_M1037_g N_A_2199_74#_c_1071_n 0.014515f $X=12.035 $Y=2.46 $X2=0
+ $Y2=0
cc_736 N_S1_M1032_g N_A_2199_74#_c_1060_n 8.63924e-19 $X=11.535 $Y=2.46 $X2=0
+ $Y2=0
cc_737 N_S1_c_843_n N_A_2199_74#_c_1061_n 0.00151635f $X=12.315 $Y=1.36 $X2=0
+ $Y2=0
cc_738 N_S1_c_845_n N_A_2199_74#_c_1061_n 0.0293853f $X=12.665 $Y=1.455 $X2=0
+ $Y2=0
cc_739 N_S1_c_843_n N_A_2199_74#_c_1043_n 5.84221e-19 $X=12.315 $Y=1.36 $X2=0
+ $Y2=0
cc_740 N_S1_c_845_n N_A_2199_74#_c_1077_n 0.0170653f $X=12.665 $Y=1.455 $X2=0
+ $Y2=0
cc_741 N_S1_c_838_n N_A_2199_74#_c_1045_n 0.00475331f $X=14.285 $Y=1.22 $X2=0
+ $Y2=0
cc_742 N_S1_c_842_n N_A_2199_74#_c_1045_n 0.0274492f $X=13.54 $Y=1.215 $X2=0
+ $Y2=0
cc_743 N_S1_c_844_n N_A_2199_74#_c_1045_n 8.35195e-19 $X=13.87 $Y=1.385 $X2=0
+ $Y2=0
cc_744 N_S1_c_838_n N_A_2199_74#_c_1046_n 0.0160644f $X=14.285 $Y=1.22 $X2=0
+ $Y2=0
cc_745 N_S1_c_838_n N_A_2199_74#_c_1047_n 0.00694011f $X=14.285 $Y=1.22 $X2=0
+ $Y2=0
cc_746 N_S1_c_841_n N_A_2199_74#_c_1047_n 0.00251423f $X=14.3 $Y=1.37 $X2=0
+ $Y2=0
cc_747 N_S1_M1044_g N_A_2199_74#_c_1048_n 0.00285462f $X=14.3 $Y=2.4 $X2=0 $Y2=0
cc_748 N_S1_c_841_n N_A_2199_74#_c_1048_n 0.00746893f $X=14.3 $Y=1.37 $X2=0
+ $Y2=0
cc_749 N_S1_M1017_g N_A_2199_74#_c_1050_n 0.0123838f $X=11.355 $Y=0.69 $X2=0
+ $Y2=0
cc_750 N_S1_M1019_g N_A_2199_74#_c_1050_n 4.89925e-19 $X=11.945 $Y=0.69 $X2=0
+ $Y2=0
cc_751 N_S1_M1019_g N_A_2199_74#_c_1088_n 0.00816632f $X=11.945 $Y=0.69 $X2=0
+ $Y2=0
cc_752 N_S1_c_840_n N_A_2199_74#_c_1088_n 0.00448553f $X=12.125 $Y=1.36 $X2=0
+ $Y2=0
cc_753 N_S1_M1017_g N_A_2199_74#_c_1051_n 8.90513e-19 $X=11.355 $Y=0.69 $X2=0
+ $Y2=0
cc_754 N_S1_M1019_g N_A_2199_74#_c_1051_n 0.00988861f $X=11.945 $Y=0.69 $X2=0
+ $Y2=0
cc_755 N_S1_c_841_n N_A_2199_74#_c_1054_n 0.00956567f $X=14.3 $Y=1.37 $X2=0
+ $Y2=0
cc_756 N_S1_M1044_g N_VPWR_c_1247_n 0.0198695f $X=14.3 $Y=2.4 $X2=0 $Y2=0
cc_757 N_S1_M1032_g N_VPWR_c_1255_n 0.00333926f $X=11.535 $Y=2.46 $X2=0 $Y2=0
cc_758 N_S1_M1037_g N_VPWR_c_1255_n 0.00333926f $X=12.035 $Y=2.46 $X2=0 $Y2=0
cc_759 N_S1_M1044_g N_VPWR_c_1255_n 0.0050621f $X=14.3 $Y=2.4 $X2=0 $Y2=0
cc_760 N_S1_M1032_g N_VPWR_c_1240_n 0.00428309f $X=11.535 $Y=2.46 $X2=0 $Y2=0
cc_761 N_S1_M1037_g N_VPWR_c_1240_n 0.00423742f $X=12.035 $Y=2.46 $X2=0 $Y2=0
cc_762 N_S1_M1044_g N_VPWR_c_1240_n 0.0100401f $X=14.3 $Y=2.4 $X2=0 $Y2=0
cc_763 N_S1_M1019_g N_A_509_392#_c_1516_n 0.00609692f $X=11.945 $Y=0.69 $X2=0
+ $Y2=0
cc_764 N_S1_c_840_n N_A_509_392#_c_1516_n 0.0100701f $X=12.125 $Y=1.36 $X2=0
+ $Y2=0
cc_765 N_S1_c_845_n N_A_509_392#_c_1516_n 0.0135925f $X=12.665 $Y=1.455 $X2=0
+ $Y2=0
cc_766 N_S1_M1017_g N_A_509_392#_c_1517_n 6.78751e-19 $X=11.355 $Y=0.69 $X2=0
+ $Y2=0
cc_767 N_S1_M1019_g N_A_509_392#_c_1517_n 0.00528673f $X=11.945 $Y=0.69 $X2=0
+ $Y2=0
cc_768 N_S1_c_845_n N_A_509_392#_c_1599_n 0.00877217f $X=12.665 $Y=1.455 $X2=0
+ $Y2=0
cc_769 N_S1_c_846_n N_A_509_392#_c_1599_n 0.0128809f $X=12.835 $Y=1.455 $X2=0
+ $Y2=0
cc_770 N_S1_M1019_g N_A_509_392#_c_1521_n 0.00323735f $X=11.945 $Y=0.69 $X2=0
+ $Y2=0
cc_771 N_S1_c_843_n N_A_509_392#_c_1521_n 0.00385917f $X=12.315 $Y=1.36 $X2=0
+ $Y2=0
cc_772 N_S1_c_845_n N_A_509_392#_c_1521_n 0.0137977f $X=12.665 $Y=1.455 $X2=0
+ $Y2=0
cc_773 N_S1_c_842_n N_A_509_392#_c_1604_n 0.0196914f $X=13.54 $Y=1.215 $X2=0
+ $Y2=0
cc_774 N_S1_M1032_g N_A_509_392#_c_1530_n 0.00751613f $X=11.535 $Y=2.46 $X2=0
+ $Y2=0
cc_775 N_S1_M1032_g N_A_509_392#_c_1533_n 0.00170083f $X=11.535 $Y=2.46 $X2=0
+ $Y2=0
cc_776 N_S1_M1017_g N_A_509_392#_c_1522_n 3.16363e-19 $X=11.355 $Y=0.69 $X2=0
+ $Y2=0
cc_777 N_S1_M1032_g N_A_509_392#_c_1522_n 0.00437332f $X=11.535 $Y=2.46 $X2=0
+ $Y2=0
cc_778 N_S1_M1019_g N_A_509_392#_c_1522_n 0.00546568f $X=11.945 $Y=0.69 $X2=0
+ $Y2=0
cc_779 N_S1_M1037_g N_A_509_392#_c_1522_n 0.017577f $X=12.035 $Y=2.46 $X2=0
+ $Y2=0
cc_780 N_S1_c_840_n N_A_509_392#_c_1522_n 0.0281339f $X=12.125 $Y=1.36 $X2=0
+ $Y2=0
cc_781 N_S1_c_845_n N_A_509_392#_c_1522_n 0.0403568f $X=12.665 $Y=1.455 $X2=0
+ $Y2=0
cc_782 N_S1_M1017_g N_A_1191_121#_c_1704_n 0.00687329f $X=11.355 $Y=0.69 $X2=0
+ $Y2=0
cc_783 N_S1_c_840_n N_A_1191_121#_c_1704_n 0.00219734f $X=12.125 $Y=1.36 $X2=0
+ $Y2=0
cc_784 N_S1_M1032_g N_A_1191_121#_c_1715_n 0.00447947f $X=11.535 $Y=2.46 $X2=0
+ $Y2=0
cc_785 N_S1_M1017_g N_A_1191_121#_c_1706_n 0.0115258f $X=11.355 $Y=0.69 $X2=0
+ $Y2=0
cc_786 N_S1_M1019_g N_A_1191_121#_c_1706_n 0.00147484f $X=11.945 $Y=0.69 $X2=0
+ $Y2=0
cc_787 N_S1_M1032_g N_A_1191_121#_c_1716_n 0.0123831f $X=11.535 $Y=2.46 $X2=0
+ $Y2=0
cc_788 N_S1_M1037_g N_A_1191_121#_c_1716_n 0.0106408f $X=12.035 $Y=2.46 $X2=0
+ $Y2=0
cc_789 N_S1_M1032_g N_A_1191_121#_c_1719_n 2.22328e-19 $X=11.535 $Y=2.46 $X2=0
+ $Y2=0
cc_790 N_S1_M1044_g N_X_c_1954_n 2.62384e-19 $X=14.3 $Y=2.4 $X2=0 $Y2=0
cc_791 N_S1_c_838_n N_VGND_c_2040_n 0.00177323f $X=14.285 $Y=1.22 $X2=0 $Y2=0
cc_792 N_S1_M1017_g N_VGND_c_2048_n 0.00278271f $X=11.355 $Y=0.69 $X2=0 $Y2=0
cc_793 N_S1_M1019_g N_VGND_c_2048_n 0.00311652f $X=11.945 $Y=0.69 $X2=0 $Y2=0
cc_794 N_S1_c_838_n N_VGND_c_2048_n 0.00278271f $X=14.285 $Y=1.22 $X2=0 $Y2=0
cc_795 N_S1_M1017_g N_VGND_c_2058_n 0.00359811f $X=11.355 $Y=0.69 $X2=0 $Y2=0
cc_796 N_S1_M1019_g N_VGND_c_2058_n 0.00396569f $X=11.945 $Y=0.69 $X2=0 $Y2=0
cc_797 N_S1_c_838_n N_VGND_c_2058_n 0.00360685f $X=14.285 $Y=1.22 $X2=0 $Y2=0
cc_798 N_A_2489_347#_c_955_n N_A_2199_74#_c_1071_n 0.00233756f $X=12.535
+ $Y=1.885 $X2=0 $Y2=0
cc_799 N_A_2489_347#_c_955_n N_A_2199_74#_c_1061_n 0.00316619f $X=12.535
+ $Y=1.885 $X2=0 $Y2=0
cc_800 N_A_2489_347#_c_956_n N_A_2199_74#_c_1061_n 5.1526e-19 $X=13.035 $Y=1.885
+ $X2=0 $Y2=0
cc_801 N_A_2489_347#_c_955_n N_A_2199_74#_c_1096_n 0.00657868f $X=12.535
+ $Y=1.885 $X2=0 $Y2=0
cc_802 N_A_2489_347#_c_956_n N_A_2199_74#_c_1096_n 2.72638e-19 $X=13.035
+ $Y=1.885 $X2=0 $Y2=0
cc_803 N_A_2489_347#_c_955_n N_A_2199_74#_c_1077_n 0.0115135f $X=12.535 $Y=1.885
+ $X2=0 $Y2=0
cc_804 N_A_2489_347#_c_956_n N_A_2199_74#_c_1077_n 0.0163264f $X=13.035 $Y=1.885
+ $X2=0 $Y2=0
cc_805 N_A_2489_347#_c_952_n N_A_2199_74#_c_1077_n 0.00954425f $X=13.165
+ $Y=1.635 $X2=0 $Y2=0
cc_806 N_A_2489_347#_c_953_n N_A_2199_74#_c_1077_n 0.00408375f $X=13.165
+ $Y=1.635 $X2=0 $Y2=0
cc_807 N_A_2489_347#_M1015_g N_A_2199_74#_c_1044_n 0.0116317f $X=12.795 $Y=0.69
+ $X2=0 $Y2=0
cc_808 N_A_2489_347#_M1048_g N_A_2199_74#_c_1044_n 0.0137009f $X=13.225 $Y=0.69
+ $X2=0 $Y2=0
cc_809 N_A_2489_347#_c_957_n N_A_2199_74#_c_1062_n 0.0120254f $X=13.875 $Y=1.805
+ $X2=0 $Y2=0
cc_810 N_A_2489_347#_c_958_n N_A_2199_74#_c_1062_n 0.00830695f $X=14.04 $Y=1.985
+ $X2=0 $Y2=0
cc_811 N_A_2489_347#_c_952_n N_A_2199_74#_c_1062_n 0.0146444f $X=13.165 $Y=1.635
+ $X2=0 $Y2=0
cc_812 N_A_2489_347#_c_953_n N_A_2199_74#_c_1062_n 0.00130939f $X=13.165
+ $Y=1.635 $X2=0 $Y2=0
cc_813 N_A_2489_347#_c_956_n N_A_2199_74#_c_1063_n 4.81024e-19 $X=13.035
+ $Y=1.885 $X2=0 $Y2=0
cc_814 N_A_2489_347#_c_958_n N_A_2199_74#_c_1063_n 0.0345589f $X=14.04 $Y=1.985
+ $X2=0 $Y2=0
cc_815 N_A_2489_347#_c_954_n N_A_2199_74#_c_1045_n 0.0244318f $X=14.07 $Y=0.775
+ $X2=0 $Y2=0
cc_816 N_A_2489_347#_M1014_s N_A_2199_74#_c_1046_n 0.00273752f $X=13.925 $Y=0.37
+ $X2=0 $Y2=0
cc_817 N_A_2489_347#_c_954_n N_A_2199_74#_c_1046_n 0.0184007f $X=14.07 $Y=0.775
+ $X2=0 $Y2=0
cc_818 N_A_2489_347#_c_951_n N_A_2199_74#_c_1047_n 0.0135902f $X=14.12 $Y=1.72
+ $X2=0 $Y2=0
cc_819 N_A_2489_347#_c_951_n N_A_2199_74#_c_1048_n 0.0255059f $X=14.12 $Y=1.72
+ $X2=0 $Y2=0
cc_820 N_A_2489_347#_M1015_g N_A_2199_74#_c_1051_n 0.00280783f $X=12.795 $Y=0.69
+ $X2=0 $Y2=0
cc_821 N_A_2489_347#_c_958_n N_VPWR_c_1247_n 0.0416899f $X=14.04 $Y=1.985 $X2=0
+ $Y2=0
cc_822 N_A_2489_347#_c_962_n N_VPWR_c_1247_n 0.00352479f $X=14.04 $Y=1.805 $X2=0
+ $Y2=0
cc_823 N_A_2489_347#_c_955_n N_VPWR_c_1255_n 0.00333926f $X=12.535 $Y=1.885
+ $X2=0 $Y2=0
cc_824 N_A_2489_347#_c_956_n N_VPWR_c_1255_n 0.00517089f $X=13.035 $Y=1.885
+ $X2=0 $Y2=0
cc_825 N_A_2489_347#_c_958_n N_VPWR_c_1255_n 0.0146357f $X=14.04 $Y=1.985 $X2=0
+ $Y2=0
cc_826 N_A_2489_347#_c_955_n N_VPWR_c_1240_n 0.00423742f $X=12.535 $Y=1.885
+ $X2=0 $Y2=0
cc_827 N_A_2489_347#_c_956_n N_VPWR_c_1240_n 0.00984196f $X=13.035 $Y=1.885
+ $X2=0 $Y2=0
cc_828 N_A_2489_347#_c_958_n N_VPWR_c_1240_n 0.0121141f $X=14.04 $Y=1.985 $X2=0
+ $Y2=0
cc_829 N_A_2489_347#_M1015_g N_A_509_392#_c_1599_n 0.010582f $X=12.795 $Y=0.69
+ $X2=0 $Y2=0
cc_830 N_A_2489_347#_M1015_g N_A_509_392#_c_1521_n 0.00360839f $X=12.795 $Y=0.69
+ $X2=0 $Y2=0
cc_831 N_A_2489_347#_M1015_g N_A_509_392#_c_1604_n 0.00828563f $X=12.795 $Y=0.69
+ $X2=0 $Y2=0
cc_832 N_A_2489_347#_M1048_g N_A_509_392#_c_1604_n 0.00453241f $X=13.225 $Y=0.69
+ $X2=0 $Y2=0
cc_833 N_A_2489_347#_c_953_n N_A_509_392#_c_1522_n 9.1605e-19 $X=13.165 $Y=1.635
+ $X2=0 $Y2=0
cc_834 N_A_2489_347#_c_955_n N_A_1191_121#_c_1716_n 0.0121668f $X=12.535
+ $Y=1.885 $X2=0 $Y2=0
cc_835 N_A_2489_347#_c_956_n N_A_1191_121#_c_1716_n 0.00710719f $X=13.035
+ $Y=1.885 $X2=0 $Y2=0
cc_836 N_A_2489_347#_c_956_n N_A_1191_121#_c_1787_n 0.00632425f $X=13.035
+ $Y=1.885 $X2=0 $Y2=0
cc_837 N_A_2489_347#_c_962_n N_X_c_1956_n 6.16393e-19 $X=14.04 $Y=1.805 $X2=0
+ $Y2=0
cc_838 N_A_2489_347#_M1015_g N_VGND_c_2048_n 0.00278271f $X=12.795 $Y=0.69 $X2=0
+ $Y2=0
cc_839 N_A_2489_347#_M1048_g N_VGND_c_2048_n 0.00278271f $X=13.225 $Y=0.69 $X2=0
+ $Y2=0
cc_840 N_A_2489_347#_M1015_g N_VGND_c_2058_n 0.0035536f $X=12.795 $Y=0.69 $X2=0
+ $Y2=0
cc_841 N_A_2489_347#_M1048_g N_VGND_c_2058_n 0.00358427f $X=13.225 $Y=0.69 $X2=0
+ $Y2=0
cc_842 N_A_2199_74#_M1010_g N_VPWR_c_1247_n 0.00382644f $X=14.815 $Y=2.4 $X2=0
+ $Y2=0
cc_843 N_A_2199_74#_c_1048_n N_VPWR_c_1247_n 0.0145005f $X=14.545 $Y=1.465 $X2=0
+ $Y2=0
cc_844 N_A_2199_74#_c_1049_n N_VPWR_c_1247_n 0.0129622f $X=16.125 $Y=1.465 $X2=0
+ $Y2=0
cc_845 N_A_2199_74#_M1026_g N_VPWR_c_1248_n 0.00366558f $X=15.265 $Y=2.4 $X2=0
+ $Y2=0
cc_846 N_A_2199_74#_M1030_g N_VPWR_c_1248_n 0.00250919f $X=15.765 $Y=2.4 $X2=0
+ $Y2=0
cc_847 N_A_2199_74#_M1034_g N_VPWR_c_1250_n 0.00643907f $X=16.215 $Y=2.4 $X2=0
+ $Y2=0
cc_848 N_A_2199_74#_c_1063_n N_VPWR_c_1255_n 0.0146357f $X=13.31 $Y=2.485 $X2=0
+ $Y2=0
cc_849 N_A_2199_74#_M1010_g N_VPWR_c_1257_n 0.005209f $X=14.815 $Y=2.4 $X2=0
+ $Y2=0
cc_850 N_A_2199_74#_M1026_g N_VPWR_c_1257_n 0.005209f $X=15.265 $Y=2.4 $X2=0
+ $Y2=0
cc_851 N_A_2199_74#_M1030_g N_VPWR_c_1263_n 0.005209f $X=15.765 $Y=2.4 $X2=0
+ $Y2=0
cc_852 N_A_2199_74#_M1034_g N_VPWR_c_1263_n 0.005209f $X=16.215 $Y=2.4 $X2=0
+ $Y2=0
cc_853 N_A_2199_74#_M1010_g N_VPWR_c_1240_n 0.00982289f $X=14.815 $Y=2.4 $X2=0
+ $Y2=0
cc_854 N_A_2199_74#_M1026_g N_VPWR_c_1240_n 0.00982754f $X=15.265 $Y=2.4 $X2=0
+ $Y2=0
cc_855 N_A_2199_74#_M1030_g N_VPWR_c_1240_n 0.00982082f $X=15.765 $Y=2.4 $X2=0
+ $Y2=0
cc_856 N_A_2199_74#_M1034_g N_VPWR_c_1240_n 0.00985583f $X=16.215 $Y=2.4 $X2=0
+ $Y2=0
cc_857 N_A_2199_74#_c_1063_n N_VPWR_c_1240_n 0.0121141f $X=13.31 $Y=2.485 $X2=0
+ $Y2=0
cc_858 N_A_2199_74#_c_1044_n N_A_509_392#_M1015_s 0.00176461f $X=13.345 $Y=0.34
+ $X2=0 $Y2=0
cc_859 N_A_2199_74#_c_1071_n N_A_509_392#_M1032_s 0.00420664f $X=12.145 $Y=2.65
+ $X2=0 $Y2=0
cc_860 N_A_2199_74#_M1019_s N_A_509_392#_c_1516_n 0.00394438f $X=12.02 $Y=0.37
+ $X2=0 $Y2=0
cc_861 N_A_2199_74#_c_1043_n N_A_509_392#_c_1516_n 0.00829606f $X=12.493
+ $Y=0.437 $X2=0 $Y2=0
cc_862 N_A_2199_74#_c_1088_n N_A_509_392#_c_1516_n 0.00937046f $X=11.985 $Y=0.51
+ $X2=0 $Y2=0
cc_863 N_A_2199_74#_c_1050_n N_A_509_392#_c_1517_n 0.0117142f $X=11.265 $Y=0.68
+ $X2=0 $Y2=0
cc_864 N_A_2199_74#_c_1088_n N_A_509_392#_c_1517_n 0.0216666f $X=11.985 $Y=0.51
+ $X2=0 $Y2=0
cc_865 N_A_2199_74#_M1019_s N_A_509_392#_c_1599_n 0.00500868f $X=12.02 $Y=0.37
+ $X2=0 $Y2=0
cc_866 N_A_2199_74#_c_1044_n N_A_509_392#_c_1599_n 0.00445011f $X=13.345 $Y=0.34
+ $X2=0 $Y2=0
cc_867 N_A_2199_74#_c_1052_n N_A_509_392#_c_1599_n 0.0125748f $X=12.675 $Y=0.437
+ $X2=0 $Y2=0
cc_868 N_A_2199_74#_M1019_s N_A_509_392#_c_1521_n 0.00692408f $X=12.02 $Y=0.37
+ $X2=0 $Y2=0
cc_869 N_A_2199_74#_c_1043_n N_A_509_392#_c_1521_n 0.0131573f $X=12.493 $Y=0.437
+ $X2=0 $Y2=0
cc_870 N_A_2199_74#_c_1044_n N_A_509_392#_c_1604_n 0.0142275f $X=13.345 $Y=0.34
+ $X2=0 $Y2=0
cc_871 N_A_2199_74#_c_1042_n N_A_509_392#_c_1530_n 0.0390311f $X=11.31 $Y=2.105
+ $X2=0 $Y2=0
cc_872 N_A_2199_74#_c_1071_n N_A_509_392#_c_1530_n 0.00380869f $X=12.145 $Y=2.65
+ $X2=0 $Y2=0
cc_873 N_A_2199_74#_c_1042_n N_A_509_392#_c_1533_n 0.00230511f $X=11.31 $Y=2.105
+ $X2=0 $Y2=0
cc_874 N_A_2199_74#_c_1071_n N_A_509_392#_c_1533_n 0.0021623f $X=12.145 $Y=2.65
+ $X2=0 $Y2=0
cc_875 N_A_2199_74#_c_1061_n N_A_509_392#_c_1533_n 0.00133571f $X=12.31 $Y=2.23
+ $X2=0 $Y2=0
cc_876 N_A_2199_74#_c_1042_n N_A_509_392#_c_1522_n 0.0847402f $X=11.31 $Y=2.105
+ $X2=0 $Y2=0
cc_877 N_A_2199_74#_c_1071_n N_A_509_392#_c_1522_n 0.0182199f $X=12.145 $Y=2.65
+ $X2=0 $Y2=0
cc_878 N_A_2199_74#_c_1061_n N_A_509_392#_c_1522_n 0.0108722f $X=12.31 $Y=2.23
+ $X2=0 $Y2=0
cc_879 N_A_2199_74#_c_1088_n N_A_1191_121#_M1017_d 0.00871026f $X=11.985 $Y=0.51
+ $X2=0 $Y2=0
cc_880 N_A_2199_74#_c_1077_n N_A_1191_121#_M1028_d 0.00535325f $X=13.145
+ $Y=2.145 $X2=0 $Y2=0
cc_881 N_A_2199_74#_c_1042_n N_A_1191_121#_c_1704_n 0.0539165f $X=11.31 $Y=2.105
+ $X2=0 $Y2=0
cc_882 N_A_2199_74#_c_1050_n N_A_1191_121#_c_1704_n 0.0344938f $X=11.265 $Y=0.68
+ $X2=0 $Y2=0
cc_883 N_A_2199_74#_c_1042_n N_A_1191_121#_c_1715_n 0.0355988f $X=11.31 $Y=2.105
+ $X2=0 $Y2=0
cc_884 N_A_2199_74#_c_1060_n N_A_1191_121#_c_1715_n 0.0143581f $X=11.475 $Y=2.65
+ $X2=0 $Y2=0
cc_885 N_A_2199_74#_M1017_s N_A_1191_121#_c_1706_n 0.00441657f $X=10.995 $Y=0.37
+ $X2=0 $Y2=0
cc_886 N_A_2199_74#_c_1050_n N_A_1191_121#_c_1706_n 0.0231725f $X=11.265 $Y=0.68
+ $X2=0 $Y2=0
cc_887 N_A_2199_74#_c_1088_n N_A_1191_121#_c_1706_n 0.0222818f $X=11.985 $Y=0.51
+ $X2=0 $Y2=0
cc_888 N_A_2199_74#_c_1051_n N_A_1191_121#_c_1706_n 0.012401f $X=12.155 $Y=0.51
+ $X2=0 $Y2=0
cc_889 N_A_2199_74#_M1032_d N_A_1191_121#_c_1716_n 0.00266942f $X=11.165 $Y=1.96
+ $X2=0 $Y2=0
cc_890 N_A_2199_74#_M1037_d N_A_1191_121#_c_1716_n 0.00218982f $X=12.125 $Y=1.96
+ $X2=0 $Y2=0
cc_891 N_A_2199_74#_c_1071_n N_A_1191_121#_c_1716_n 0.0528479f $X=12.145 $Y=2.65
+ $X2=0 $Y2=0
cc_892 N_A_2199_74#_c_1060_n N_A_1191_121#_c_1716_n 0.0205753f $X=11.475 $Y=2.65
+ $X2=0 $Y2=0
cc_893 N_A_2199_74#_c_1077_n N_A_1191_121#_c_1716_n 0.00318644f $X=13.145
+ $Y=2.145 $X2=0 $Y2=0
cc_894 N_A_2199_74#_c_1063_n N_A_1191_121#_c_1716_n 0.0039531f $X=13.31 $Y=2.485
+ $X2=0 $Y2=0
cc_895 N_A_2199_74#_c_1077_n N_A_1191_121#_c_1787_n 0.0189154f $X=13.145
+ $Y=2.145 $X2=0 $Y2=0
cc_896 N_A_2199_74#_c_1042_n N_A_1191_121#_c_1719_n 0.0129149f $X=11.31 $Y=2.105
+ $X2=0 $Y2=0
cc_897 N_A_2199_74#_M1010_g N_X_c_1954_n 0.0124852f $X=14.815 $Y=2.4 $X2=0 $Y2=0
cc_898 N_A_2199_74#_M1026_g N_X_c_1954_n 0.0145605f $X=15.265 $Y=2.4 $X2=0 $Y2=0
cc_899 N_A_2199_74#_M1030_g N_X_c_1954_n 6.79538e-19 $X=15.765 $Y=2.4 $X2=0
+ $Y2=0
cc_900 N_A_2199_74#_M1020_g N_X_c_1947_n 0.00760419f $X=15.015 $Y=0.74 $X2=0
+ $Y2=0
cc_901 N_A_2199_74#_M1027_g N_X_c_1947_n 3.97481e-19 $X=15.445 $Y=0.74 $X2=0
+ $Y2=0
cc_902 N_A_2199_74#_M1026_g N_X_c_1955_n 0.0132272f $X=15.265 $Y=2.4 $X2=0 $Y2=0
cc_903 N_A_2199_74#_M1030_g N_X_c_1955_n 0.0132272f $X=15.765 $Y=2.4 $X2=0 $Y2=0
cc_904 N_A_2199_74#_c_1049_n N_X_c_1955_n 0.045409f $X=16.125 $Y=1.465 $X2=0
+ $Y2=0
cc_905 N_A_2199_74#_c_1054_n N_X_c_1955_n 0.00369047f $X=16.215 $Y=1.465 $X2=0
+ $Y2=0
cc_906 N_A_2199_74#_M1010_g N_X_c_1956_n 0.00301176f $X=14.815 $Y=2.4 $X2=0
+ $Y2=0
cc_907 N_A_2199_74#_M1026_g N_X_c_1956_n 0.00135419f $X=15.265 $Y=2.4 $X2=0
+ $Y2=0
cc_908 N_A_2199_74#_c_1049_n N_X_c_1956_n 0.0275631f $X=16.125 $Y=1.465 $X2=0
+ $Y2=0
cc_909 N_A_2199_74#_c_1054_n N_X_c_1956_n 0.00245159f $X=16.215 $Y=1.465 $X2=0
+ $Y2=0
cc_910 N_A_2199_74#_M1027_g N_X_c_1948_n 0.0124899f $X=15.445 $Y=0.74 $X2=0
+ $Y2=0
cc_911 N_A_2199_74#_M1035_g N_X_c_1948_n 0.01115f $X=15.875 $Y=0.74 $X2=0 $Y2=0
cc_912 N_A_2199_74#_c_1049_n N_X_c_1948_n 0.0447482f $X=16.125 $Y=1.465 $X2=0
+ $Y2=0
cc_913 N_A_2199_74#_c_1054_n N_X_c_1948_n 0.00263605f $X=16.215 $Y=1.465 $X2=0
+ $Y2=0
cc_914 N_A_2199_74#_M1020_g N_X_c_1949_n 0.00245337f $X=15.015 $Y=0.74 $X2=0
+ $Y2=0
cc_915 N_A_2199_74#_c_1049_n N_X_c_1949_n 0.0209731f $X=16.125 $Y=1.465 $X2=0
+ $Y2=0
cc_916 N_A_2199_74#_c_1054_n N_X_c_1949_n 0.00272398f $X=16.215 $Y=1.465 $X2=0
+ $Y2=0
cc_917 N_A_2199_74#_M1026_g N_X_c_1957_n 6.46654e-19 $X=15.265 $Y=2.4 $X2=0
+ $Y2=0
cc_918 N_A_2199_74#_M1030_g N_X_c_1957_n 0.0139698f $X=15.765 $Y=2.4 $X2=0 $Y2=0
cc_919 N_A_2199_74#_M1034_g N_X_c_1957_n 0.0184131f $X=16.215 $Y=2.4 $X2=0 $Y2=0
cc_920 N_A_2199_74#_M1027_g N_X_c_1950_n 6.20738e-19 $X=15.445 $Y=0.74 $X2=0
+ $Y2=0
cc_921 N_A_2199_74#_M1035_g N_X_c_1950_n 0.00866629f $X=15.875 $Y=0.74 $X2=0
+ $Y2=0
cc_922 N_A_2199_74#_M1051_g N_X_c_1950_n 3.97481e-19 $X=16.305 $Y=0.74 $X2=0
+ $Y2=0
cc_923 N_A_2199_74#_M1034_g N_X_c_1958_n 0.0159354f $X=16.215 $Y=2.4 $X2=0 $Y2=0
cc_924 N_A_2199_74#_c_1049_n N_X_c_1958_n 0.0038938f $X=16.125 $Y=1.465 $X2=0
+ $Y2=0
cc_925 N_A_2199_74#_c_1054_n N_X_c_1958_n 0.00234636f $X=16.215 $Y=1.465 $X2=0
+ $Y2=0
cc_926 N_A_2199_74#_M1051_g N_X_c_1951_n 0.0158737f $X=16.305 $Y=0.74 $X2=0
+ $Y2=0
cc_927 N_A_2199_74#_c_1049_n N_X_c_1951_n 0.0025934f $X=16.125 $Y=1.465 $X2=0
+ $Y2=0
cc_928 N_A_2199_74#_M1030_g N_X_c_1959_n 0.00135419f $X=15.765 $Y=2.4 $X2=0
+ $Y2=0
cc_929 N_A_2199_74#_M1034_g N_X_c_1959_n 0.00135419f $X=16.215 $Y=2.4 $X2=0
+ $Y2=0
cc_930 N_A_2199_74#_c_1049_n N_X_c_1959_n 0.0275631f $X=16.125 $Y=1.465 $X2=0
+ $Y2=0
cc_931 N_A_2199_74#_c_1054_n N_X_c_1959_n 0.00245159f $X=16.215 $Y=1.465 $X2=0
+ $Y2=0
cc_932 N_A_2199_74#_M1035_g N_X_c_1952_n 9.7541e-19 $X=15.875 $Y=0.74 $X2=0
+ $Y2=0
cc_933 N_A_2199_74#_c_1049_n N_X_c_1952_n 0.0209731f $X=16.125 $Y=1.465 $X2=0
+ $Y2=0
cc_934 N_A_2199_74#_c_1054_n N_X_c_1952_n 0.00272398f $X=16.215 $Y=1.465 $X2=0
+ $Y2=0
cc_935 N_A_2199_74#_M1034_g X 0.00632079f $X=16.215 $Y=2.4 $X2=0 $Y2=0
cc_936 N_A_2199_74#_M1051_g X 0.0169854f $X=16.305 $Y=0.74 $X2=0 $Y2=0
cc_937 N_A_2199_74#_c_1049_n X 0.0209823f $X=16.125 $Y=1.465 $X2=0 $Y2=0
cc_938 N_A_2199_74#_c_1046_n N_VGND_M1014_d 5.37942e-19 $X=14.375 $Y=0.34 $X2=0
+ $Y2=0
cc_939 N_A_2199_74#_c_1047_n N_VGND_M1014_d 0.00934994f $X=14.46 $Y=1.3 $X2=0
+ $Y2=0
cc_940 N_A_2199_74#_M1020_g N_VGND_c_2040_n 0.00262092f $X=15.015 $Y=0.74 $X2=0
+ $Y2=0
cc_941 N_A_2199_74#_c_1046_n N_VGND_c_2040_n 0.014187f $X=14.375 $Y=0.34 $X2=0
+ $Y2=0
cc_942 N_A_2199_74#_c_1047_n N_VGND_c_2040_n 0.0512232f $X=14.46 $Y=1.3 $X2=0
+ $Y2=0
cc_943 N_A_2199_74#_c_1049_n N_VGND_c_2040_n 0.0148609f $X=16.125 $Y=1.465 $X2=0
+ $Y2=0
cc_944 N_A_2199_74#_c_1054_n N_VGND_c_2040_n 8.18019e-19 $X=16.215 $Y=1.465
+ $X2=0 $Y2=0
cc_945 N_A_2199_74#_M1020_g N_VGND_c_2041_n 5.05592e-19 $X=15.015 $Y=0.74 $X2=0
+ $Y2=0
cc_946 N_A_2199_74#_M1027_g N_VGND_c_2041_n 0.00914496f $X=15.445 $Y=0.74 $X2=0
+ $Y2=0
cc_947 N_A_2199_74#_M1035_g N_VGND_c_2041_n 0.00183835f $X=15.875 $Y=0.74 $X2=0
+ $Y2=0
cc_948 N_A_2199_74#_M1035_g N_VGND_c_2043_n 5.04273e-19 $X=15.875 $Y=0.74 $X2=0
+ $Y2=0
cc_949 N_A_2199_74#_M1051_g N_VGND_c_2043_n 0.0112604f $X=16.305 $Y=0.74 $X2=0
+ $Y2=0
cc_950 N_A_2199_74#_c_1046_n N_VGND_c_2048_n 0.0567846f $X=14.375 $Y=0.34 $X2=0
+ $Y2=0
cc_951 N_A_2199_74#_c_1088_n N_VGND_c_2048_n 0.00265664f $X=11.985 $Y=0.51 $X2=0
+ $Y2=0
cc_952 N_A_2199_74#_c_1051_n N_VGND_c_2048_n 0.089252f $X=12.155 $Y=0.51 $X2=0
+ $Y2=0
cc_953 N_A_2199_74#_c_1053_n N_VGND_c_2048_n 0.0237213f $X=13.51 $Y=0.34 $X2=0
+ $Y2=0
cc_954 N_A_2199_74#_M1020_g N_VGND_c_2052_n 0.00434272f $X=15.015 $Y=0.74 $X2=0
+ $Y2=0
cc_955 N_A_2199_74#_M1027_g N_VGND_c_2052_n 0.00383152f $X=15.445 $Y=0.74 $X2=0
+ $Y2=0
cc_956 N_A_2199_74#_M1035_g N_VGND_c_2053_n 0.00434272f $X=15.875 $Y=0.74 $X2=0
+ $Y2=0
cc_957 N_A_2199_74#_M1051_g N_VGND_c_2053_n 0.00383152f $X=16.305 $Y=0.74 $X2=0
+ $Y2=0
cc_958 N_A_2199_74#_M1020_g N_VGND_c_2058_n 0.00822542f $X=15.015 $Y=0.74 $X2=0
+ $Y2=0
cc_959 N_A_2199_74#_M1027_g N_VGND_c_2058_n 0.0075754f $X=15.445 $Y=0.74 $X2=0
+ $Y2=0
cc_960 N_A_2199_74#_M1035_g N_VGND_c_2058_n 0.00820284f $X=15.875 $Y=0.74 $X2=0
+ $Y2=0
cc_961 N_A_2199_74#_M1051_g N_VGND_c_2058_n 0.0075754f $X=16.305 $Y=0.74 $X2=0
+ $Y2=0
cc_962 N_A_2199_74#_c_1046_n N_VGND_c_2058_n 0.032237f $X=14.375 $Y=0.34 $X2=0
+ $Y2=0
cc_963 N_A_2199_74#_c_1088_n N_VGND_c_2058_n 0.00514655f $X=11.985 $Y=0.51 $X2=0
+ $Y2=0
cc_964 N_A_2199_74#_c_1051_n N_VGND_c_2058_n 0.0500945f $X=12.155 $Y=0.51 $X2=0
+ $Y2=0
cc_965 N_A_2199_74#_c_1053_n N_VGND_c_2058_n 0.0128418f $X=13.51 $Y=0.34 $X2=0
+ $Y2=0
cc_966 N_VPWR_c_1242_n N_A_119_392#_c_1422_n 0.00726648f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_967 N_VPWR_c_1242_n N_A_119_392#_c_1423_n 0.0283172f $X=0.28 $Y=2.115 $X2=0
+ $Y2=0
cc_968 N_VPWR_c_1243_n N_A_119_392#_c_1423_n 0.0227494f $X=1.18 $Y=2.475 $X2=0
+ $Y2=0
cc_969 N_VPWR_c_1259_n N_A_119_392#_c_1423_n 0.0144623f $X=1.095 $Y=3.33 $X2=0
+ $Y2=0
cc_970 N_VPWR_c_1240_n N_A_119_392#_c_1423_n 0.0118344f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_971 N_VPWR_M1004_s N_A_119_392#_c_1424_n 0.00332066f $X=1.045 $Y=1.96 $X2=0
+ $Y2=0
cc_972 N_VPWR_M1011_d N_A_119_392#_c_1424_n 0.00512823f $X=1.995 $Y=1.96 $X2=0
+ $Y2=0
cc_973 N_VPWR_c_1243_n N_A_119_392#_c_1424_n 0.0148589f $X=1.18 $Y=2.475 $X2=0
+ $Y2=0
cc_974 N_VPWR_M1011_d N_A_299_392#_c_1483_n 0.00538852f $X=1.995 $Y=1.96 $X2=0
+ $Y2=0
cc_975 N_VPWR_c_1244_n N_A_299_392#_c_1483_n 0.0193313f $X=2.13 $Y=2.815 $X2=0
+ $Y2=0
cc_976 N_VPWR_c_1240_n N_A_299_392#_c_1483_n 0.0153384f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_977 N_VPWR_c_1243_n N_A_299_392#_c_1485_n 0.0187702f $X=1.18 $Y=2.475 $X2=0
+ $Y2=0
cc_978 N_VPWR_c_1244_n N_A_299_392#_c_1485_n 0.011548f $X=2.13 $Y=2.815 $X2=0
+ $Y2=0
cc_979 N_VPWR_c_1260_n N_A_299_392#_c_1485_n 0.0145333f $X=2.045 $Y=3.33 $X2=0
+ $Y2=0
cc_980 N_VPWR_c_1240_n N_A_299_392#_c_1485_n 0.0119681f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_981 N_VPWR_c_1261_n N_A_509_392#_c_1524_n 0.0395821f $X=5.4 $Y=3.33 $X2=0
+ $Y2=0
cc_982 N_VPWR_c_1240_n N_A_509_392#_c_1524_n 0.0221587f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_983 N_VPWR_c_1261_n N_A_509_392#_c_1526_n 0.0594111f $X=5.4 $Y=3.33 $X2=0
+ $Y2=0
cc_984 N_VPWR_c_1240_n N_A_509_392#_c_1526_n 0.0327651f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_985 N_VPWR_c_1244_n N_A_509_392#_c_1528_n 0.0280957f $X=2.13 $Y=2.815 $X2=0
+ $Y2=0
cc_986 N_VPWR_c_1261_n N_A_509_392#_c_1528_n 0.0229864f $X=5.4 $Y=3.33 $X2=0
+ $Y2=0
cc_987 N_VPWR_c_1240_n N_A_509_392#_c_1528_n 0.0127058f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_988 N_VPWR_c_1261_n N_A_509_392#_c_1529_n 0.0235336f $X=5.4 $Y=3.33 $X2=0
+ $Y2=0
cc_989 N_VPWR_c_1240_n N_A_509_392#_c_1529_n 0.0126695f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_990 N_VPWR_c_1245_n N_A_509_392#_c_1530_n 0.0309855f $X=5.565 $Y=1.985 $X2=0
+ $Y2=0
cc_991 N_VPWR_c_1246_n N_A_509_392#_c_1530_n 0.00142931f $X=10.55 $Y=2.45 $X2=0
+ $Y2=0
cc_992 N_VPWR_c_1245_n N_A_1191_121#_c_1709_n 0.010962f $X=5.565 $Y=1.985 $X2=0
+ $Y2=0
cc_993 N_VPWR_c_1245_n N_A_1191_121#_c_1710_n 0.0565306f $X=5.565 $Y=1.985 $X2=0
+ $Y2=0
cc_994 N_VPWR_c_1262_n N_A_1191_121#_c_1710_n 0.00849124f $X=8.32 $Y=3.33 $X2=0
+ $Y2=0
cc_995 N_VPWR_c_1240_n N_A_1191_121#_c_1710_n 0.00873398f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_996 N_VPWR_M1036_s N_A_1191_121#_c_1713_n 0.00485901f $X=8.34 $Y=1.96 $X2=0
+ $Y2=0
cc_997 N_VPWR_M1038_s N_A_1191_121#_c_1713_n 0.00690064f $X=9.335 $Y=1.96 $X2=0
+ $Y2=0
cc_998 N_VPWR_M1024_s N_A_1191_121#_c_1713_n 0.00490197f $X=10.415 $Y=1.96 $X2=0
+ $Y2=0
cc_999 N_VPWR_c_1246_n N_A_1191_121#_c_1713_n 0.0118417f $X=10.55 $Y=2.45 $X2=0
+ $Y2=0
cc_1000 N_VPWR_c_1246_n N_A_1191_121#_c_1715_n 0.0458206f $X=10.55 $Y=2.45 $X2=0
+ $Y2=0
cc_1001 N_VPWR_c_1255_n N_A_1191_121#_c_1716_n 0.129486f $X=14.375 $Y=3.33 $X2=0
+ $Y2=0
cc_1002 N_VPWR_c_1240_n N_A_1191_121#_c_1716_n 0.0730129f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1003 N_VPWR_c_1246_n N_A_1191_121#_c_1717_n 0.0142846f $X=10.55 $Y=2.45 $X2=0
+ $Y2=0
cc_1004 N_VPWR_c_1255_n N_A_1191_121#_c_1717_n 0.0121867f $X=14.375 $Y=3.33
+ $X2=0 $Y2=0
cc_1005 N_VPWR_c_1240_n N_A_1191_121#_c_1717_n 0.00660921f $X=16.56 $Y=3.33
+ $X2=0 $Y2=0
cc_1006 N_VPWR_c_1262_n N_A_1288_377#_c_1871_n 0.0798496f $X=8.32 $Y=3.33 $X2=0
+ $Y2=0
cc_1007 N_VPWR_c_1240_n N_A_1288_377#_c_1871_n 0.0466173f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1008 N_VPWR_c_1262_n N_A_1288_377#_c_1872_n 0.0236566f $X=8.32 $Y=3.33 $X2=0
+ $Y2=0
cc_1009 N_VPWR_c_1240_n N_A_1288_377#_c_1872_n 0.0128296f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1010 N_VPWR_M1036_s N_A_1288_377#_c_1873_n 0.00801174f $X=8.34 $Y=1.96 $X2=0
+ $Y2=0
cc_1011 N_VPWR_M1038_s N_A_1288_377#_c_1873_n 0.0100362f $X=9.335 $Y=1.96 $X2=0
+ $Y2=0
cc_1012 N_VPWR_c_1246_n N_A_1288_377#_c_1873_n 0.0130478f $X=10.55 $Y=2.45 $X2=0
+ $Y2=0
cc_1013 N_VPWR_c_1251_n N_A_1288_377#_c_1873_n 0.0259142f $X=9.56 $Y=3.05 $X2=0
+ $Y2=0
cc_1014 N_VPWR_c_1252_n N_A_1288_377#_c_1873_n 0.0138438f $X=9.39 $Y=3.33 $X2=0
+ $Y2=0
cc_1015 N_VPWR_c_1253_n N_A_1288_377#_c_1873_n 0.0184002f $X=10.465 $Y=3.33
+ $X2=0 $Y2=0
cc_1016 N_VPWR_c_1262_n N_A_1288_377#_c_1873_n 0.00389376f $X=8.32 $Y=3.33 $X2=0
+ $Y2=0
cc_1017 N_VPWR_c_1267_n N_A_1288_377#_c_1873_n 0.024193f $X=8.485 $Y=3.05 $X2=0
+ $Y2=0
cc_1018 N_VPWR_c_1240_n N_A_1288_377#_c_1873_n 0.0475996f $X=16.56 $Y=3.33 $X2=0
+ $Y2=0
cc_1019 N_VPWR_c_1262_n N_A_1288_377#_c_1874_n 0.0116773f $X=8.32 $Y=3.33 $X2=0
+ $Y2=0
cc_1020 N_VPWR_c_1267_n N_A_1288_377#_c_1874_n 0.00872135f $X=8.485 $Y=3.05
+ $X2=0 $Y2=0
cc_1021 N_VPWR_c_1240_n N_A_1288_377#_c_1874_n 0.00646299f $X=16.56 $Y=3.33
+ $X2=0 $Y2=0
cc_1022 N_VPWR_M1036_s N_A_1468_377#_c_1926_n 0.00799039f $X=8.34 $Y=1.96 $X2=0
+ $Y2=0
cc_1023 N_VPWR_c_1247_n N_X_c_1954_n 0.0386506f $X=14.54 $Y=1.985 $X2=0 $Y2=0
cc_1024 N_VPWR_c_1248_n N_X_c_1954_n 0.0283501f $X=15.49 $Y=2.305 $X2=0 $Y2=0
cc_1025 N_VPWR_c_1257_n N_X_c_1954_n 0.0144623f $X=15.405 $Y=3.33 $X2=0 $Y2=0
cc_1026 N_VPWR_c_1240_n N_X_c_1954_n 0.0118344f $X=16.56 $Y=3.33 $X2=0 $Y2=0
cc_1027 N_VPWR_M1026_s N_X_c_1955_n 0.00218982f $X=15.355 $Y=1.84 $X2=0 $Y2=0
cc_1028 N_VPWR_c_1248_n N_X_c_1955_n 0.0167599f $X=15.49 $Y=2.305 $X2=0 $Y2=0
cc_1029 N_VPWR_c_1247_n N_X_c_1956_n 0.00711241f $X=14.54 $Y=1.985 $X2=0 $Y2=0
cc_1030 N_VPWR_c_1248_n N_X_c_1957_n 0.0322767f $X=15.49 $Y=2.305 $X2=0 $Y2=0
cc_1031 N_VPWR_c_1250_n N_X_c_1957_n 0.0323093f $X=16.49 $Y=2.305 $X2=0 $Y2=0
cc_1032 N_VPWR_c_1263_n N_X_c_1957_n 0.0144623f $X=16.325 $Y=3.33 $X2=0 $Y2=0
cc_1033 N_VPWR_c_1240_n N_X_c_1957_n 0.0118344f $X=16.56 $Y=3.33 $X2=0 $Y2=0
cc_1034 N_VPWR_M1034_s N_X_c_1958_n 0.00405359f $X=16.305 $Y=1.84 $X2=0 $Y2=0
cc_1035 N_VPWR_c_1250_n N_X_c_1958_n 0.0256273f $X=16.49 $Y=2.305 $X2=0 $Y2=0
cc_1036 N_VPWR_c_1242_n N_VGND_c_2031_n 3.21545e-19 $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_1037 N_A_119_392#_c_1424_n N_A_299_392#_M1007_s 0.0040648f $X=2.525 $Y=2.055
+ $X2=-0.19 $Y2=-0.245
cc_1038 N_A_119_392#_c_1424_n N_A_299_392#_c_1483_n 0.0587095f $X=2.525 $Y=2.055
+ $X2=0 $Y2=0
cc_1039 N_A_119_392#_c_1420_n N_A_299_392#_c_1483_n 0.00771619f $X=4.02 $Y=1.685
+ $X2=0 $Y2=0
cc_1040 N_A_119_392#_c_1424_n N_A_299_392#_c_1484_n 0.00915284f $X=2.525
+ $Y=2.055 $X2=0 $Y2=0
cc_1041 N_A_119_392#_c_1425_n N_A_299_392#_c_1484_n 0.00144817f $X=2.61 $Y=1.97
+ $X2=0 $Y2=0
cc_1042 N_A_119_392#_c_1420_n N_A_299_392#_c_1484_n 0.0256916f $X=4.02 $Y=1.685
+ $X2=0 $Y2=0
cc_1043 N_A_119_392#_c_1424_n N_A_299_392#_c_1485_n 0.01898f $X=2.525 $Y=2.055
+ $X2=0 $Y2=0
cc_1044 N_A_119_392#_c_1424_n N_A_509_392#_M1000_d 0.00487638f $X=2.525 $Y=2.055
+ $X2=0 $Y2=0
cc_1045 N_A_119_392#_c_1420_n N_A_509_392#_c_1525_n 0.0274296f $X=4.02 $Y=1.685
+ $X2=0 $Y2=0
cc_1046 N_A_119_392#_c_1428_n N_A_509_392#_c_1525_n 0.0262918f $X=4.105 $Y=2.105
+ $X2=0 $Y2=0
cc_1047 N_A_119_392#_M1045_d N_A_509_392#_c_1526_n 0.00165831f $X=3.97 $Y=1.96
+ $X2=0 $Y2=0
cc_1048 N_A_119_392#_c_1428_n N_A_509_392#_c_1526_n 0.0118736f $X=4.105 $Y=2.105
+ $X2=0 $Y2=0
cc_1049 N_A_119_392#_c_1428_n N_A_509_392#_c_1531_n 0.00151178f $X=4.105
+ $Y=2.105 $X2=0 $Y2=0
cc_1050 N_A_119_392#_c_1420_n N_A_509_392#_c_1523_n 0.0124745f $X=4.02 $Y=1.685
+ $X2=0 $Y2=0
cc_1051 N_A_119_392#_c_1428_n N_A_509_392#_c_1523_n 0.0402194f $X=4.105 $Y=2.105
+ $X2=0 $Y2=0
cc_1052 N_A_119_392#_c_1424_n N_A_299_126#_c_2282_n 0.00489672f $X=2.525
+ $Y=2.055 $X2=0 $Y2=0
cc_1053 N_A_119_392#_c_1420_n N_A_299_126#_c_2283_n 0.109901f $X=4.02 $Y=1.685
+ $X2=0 $Y2=0
cc_1054 N_A_119_392#_c_1421_n N_A_299_126#_c_2286_n 0.0145619f $X=2.695 $Y=1.685
+ $X2=0 $Y2=0
cc_1055 N_A_299_392#_c_1483_n N_A_509_392#_M1000_d 0.00680698f $X=2.99 $Y=2.395
+ $X2=0 $Y2=0
cc_1056 N_A_299_392#_M1000_s N_A_509_392#_c_1524_n 0.00192406f $X=3.02 $Y=1.96
+ $X2=0 $Y2=0
cc_1057 N_A_299_392#_c_1483_n N_A_509_392#_c_1524_n 0.00357384f $X=2.99 $Y=2.395
+ $X2=0 $Y2=0
cc_1058 N_A_299_392#_c_1491_n N_A_509_392#_c_1524_n 0.0146592f $X=3.145 $Y=2.395
+ $X2=0 $Y2=0
cc_1059 N_A_299_392#_c_1484_n N_A_509_392#_c_1525_n 0.0134237f $X=3.155 $Y=2.105
+ $X2=0 $Y2=0
cc_1060 N_A_299_392#_c_1483_n N_A_509_392#_c_1528_n 0.0210687f $X=2.99 $Y=2.395
+ $X2=0 $Y2=0
cc_1061 N_A_509_392#_c_1517_n N_A_1191_121#_M1017_d 0.00270563f $X=11.975
+ $Y=1.02 $X2=0 $Y2=0
cc_1062 N_A_509_392#_c_1530_n N_A_1191_121#_M1046_s 0.00182568f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1063 N_A_509_392#_c_1530_n N_A_1191_121#_M1050_s 0.00182568f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1064 N_A_509_392#_c_1530_n N_A_1191_121#_c_1709_n 0.00759437f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1065 N_A_509_392#_c_1530_n N_A_1191_121#_c_1710_n 0.0184402f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1066 N_A_509_392#_c_1530_n N_A_1191_121#_c_1711_n 0.0297173f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1067 N_A_509_392#_c_1530_n N_A_1191_121#_c_1713_n 0.181476f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1068 N_A_509_392#_M1032_s N_A_1191_121#_c_1716_n 0.00219516f $X=11.625
+ $Y=1.96 $X2=0 $Y2=0
cc_1069 N_A_509_392#_c_1530_n N_A_1191_121#_c_1718_n 0.0244822f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1070 N_A_509_392#_c_1530_n N_A_1191_121#_c_1719_n 0.0312882f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1071 N_A_509_392#_c_1530_n N_A_1288_377#_M1046_d 0.00200058f $X=11.615
+ $Y=2.035 $X2=-0.19 $Y2=-0.245
cc_1072 N_A_509_392#_c_1530_n N_A_1288_377#_c_1875_n 0.00903825f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1073 N_A_509_392#_c_1530_n N_A_1288_377#_c_1873_n 0.00617016f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1074 N_A_509_392#_c_1530_n N_A_1288_377#_c_1886_n 0.0027522f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1075 N_A_509_392#_c_1530_n N_A_1468_377#_c_1926_n 0.0115744f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1076 N_A_509_392#_c_1530_n N_A_1468_377#_c_1928_n 0.00266675f $X=11.615
+ $Y=2.035 $X2=0 $Y2=0
cc_1077 N_A_509_392#_c_1518_n N_VGND_c_2035_n 0.0131469f $X=2.705 $Y=0.34 $X2=0
+ $Y2=0
cc_1078 N_A_509_392#_c_1514_n N_VGND_c_2036_n 0.00284916f $X=4.375 $Y=0.34 $X2=0
+ $Y2=0
cc_1079 N_A_509_392#_c_1512_n N_VGND_c_2051_n 0.0464419f $X=3.605 $Y=0.34 $X2=0
+ $Y2=0
cc_1080 N_A_509_392#_c_1514_n N_VGND_c_2051_n 0.0617583f $X=4.375 $Y=0.34 $X2=0
+ $Y2=0
cc_1081 N_A_509_392#_c_1518_n N_VGND_c_2051_n 0.0224527f $X=2.705 $Y=0.34 $X2=0
+ $Y2=0
cc_1082 N_A_509_392#_c_1519_n N_VGND_c_2051_n 0.0115893f $X=3.69 $Y=0.34 $X2=0
+ $Y2=0
cc_1083 N_A_509_392#_c_1512_n N_VGND_c_2058_n 0.0246622f $X=3.605 $Y=0.34 $X2=0
+ $Y2=0
cc_1084 N_A_509_392#_c_1514_n N_VGND_c_2058_n 0.0318225f $X=4.375 $Y=0.34 $X2=0
+ $Y2=0
cc_1085 N_A_509_392#_c_1518_n N_VGND_c_2058_n 0.0125544f $X=2.705 $Y=0.34 $X2=0
+ $Y2=0
cc_1086 N_A_509_392#_c_1519_n N_VGND_c_2058_n 0.00583135f $X=3.69 $Y=0.34 $X2=0
+ $Y2=0
cc_1087 N_A_509_392#_c_1512_n N_A_114_126#_c_2247_n 0.0211399f $X=3.605 $Y=0.34
+ $X2=0 $Y2=0
cc_1088 N_A_509_392#_M1009_d N_A_114_126#_c_2237_n 0.00868512f $X=2.56 $Y=0.31
+ $X2=0 $Y2=0
cc_1089 N_A_509_392#_c_1512_n N_A_114_126#_c_2237_n 0.00360515f $X=3.605 $Y=0.34
+ $X2=0 $Y2=0
cc_1090 N_A_509_392#_c_1518_n N_A_114_126#_c_2237_n 0.0246598f $X=2.705 $Y=0.34
+ $X2=0 $Y2=0
cc_1091 N_A_509_392#_c_1513_n N_A_299_126#_c_2283_n 0.0138021f $X=3.69 $Y=0.87
+ $X2=0 $Y2=0
cc_1092 N_A_509_392#_c_1523_n N_A_299_126#_c_2283_n 0.0136127f $X=4.547 $Y=1.92
+ $X2=0 $Y2=0
cc_1093 N_A_509_392#_c_1514_n N_A_299_126#_c_2284_n 0.0168109f $X=4.375 $Y=0.34
+ $X2=0 $Y2=0
cc_1094 N_A_509_392#_c_1515_n N_A_299_126#_c_2284_n 0.026002f $X=4.55 $Y=0.755
+ $X2=0 $Y2=0
cc_1095 N_A_509_392#_M1009_d N_A_299_126#_c_2286_n 0.00330374f $X=2.56 $Y=0.31
+ $X2=0 $Y2=0
cc_1096 N_A_1191_121#_c_1711_n N_A_1288_377#_M1046_d 7.35179e-19 $X=6.94 $Y=1.95
+ $X2=-0.19 $Y2=-0.245
cc_1097 N_A_1191_121#_c_1713_n N_A_1288_377#_M1005_d 0.00165831f $X=10.715
+ $Y=2.03 $X2=0 $Y2=0
cc_1098 N_A_1191_121#_c_1710_n N_A_1288_377#_c_1875_n 0.0237048f $X=6.125
+ $Y=2.74 $X2=0 $Y2=0
cc_1099 N_A_1191_121#_c_1711_n N_A_1288_377#_c_1875_n 0.016716f $X=6.94 $Y=1.95
+ $X2=0 $Y2=0
cc_1100 N_A_1191_121#_c_1834_p N_A_1288_377#_c_1871_n 0.0131021f $X=7.025
+ $Y=2.57 $X2=0 $Y2=0
cc_1101 N_A_1191_121#_c_1713_n N_A_1288_377#_c_1873_n 0.0152652f $X=10.715
+ $Y=2.03 $X2=0 $Y2=0
cc_1102 N_A_1191_121#_c_1713_n N_A_1288_377#_c_1886_n 0.0153278f $X=10.715
+ $Y=2.03 $X2=0 $Y2=0
cc_1103 N_A_1191_121#_M1008_s N_A_1288_377#_c_1874_n 0.00523318f $X=7.79
+ $Y=1.885 $X2=0 $Y2=0
cc_1104 N_A_1191_121#_c_1713_n N_A_1468_377#_M1001_d 0.00312854f $X=10.715
+ $Y=2.03 $X2=-0.19 $Y2=-0.245
cc_1105 N_A_1191_121#_c_1713_n N_A_1468_377#_M1036_d 0.00166235f $X=10.715
+ $Y=2.03 $X2=0 $Y2=0
cc_1106 N_A_1191_121#_M1008_s N_A_1468_377#_c_1926_n 0.00610428f $X=7.79
+ $Y=1.885 $X2=0 $Y2=0
cc_1107 N_A_1191_121#_c_1713_n N_A_1468_377#_c_1926_n 0.0857646f $X=10.715
+ $Y=2.03 $X2=0 $Y2=0
cc_1108 N_A_1191_121#_c_1713_n N_A_1468_377#_c_1928_n 0.0149109f $X=10.715
+ $Y=2.03 $X2=0 $Y2=0
cc_1109 N_A_1191_121#_c_1699_n N_VGND_c_2036_n 0.0075116f $X=6.06 $Y=1.025 $X2=0
+ $Y2=0
cc_1110 N_A_1191_121#_c_1700_n N_VGND_c_2036_n 0.0290212f $X=6.1 $Y=0.75 $X2=0
+ $Y2=0
cc_1111 N_A_1191_121#_c_1704_n N_VGND_c_2039_n 0.0460466f $X=10.8 $Y=1.945 $X2=0
+ $Y2=0
cc_1112 N_A_1191_121#_c_1705_n N_VGND_c_2039_n 0.0146661f $X=10.885 $Y=0.34
+ $X2=0 $Y2=0
cc_1113 N_A_1191_121#_c_1700_n N_VGND_c_2045_n 0.00553716f $X=6.1 $Y=0.75 $X2=0
+ $Y2=0
cc_1114 N_A_1191_121#_c_1705_n N_VGND_c_2048_n 0.0121867f $X=10.885 $Y=0.34
+ $X2=0 $Y2=0
cc_1115 N_A_1191_121#_c_1706_n N_VGND_c_2048_n 0.0591438f $X=11.65 $Y=0.34 $X2=0
+ $Y2=0
cc_1116 N_A_1191_121#_M1017_d N_VGND_c_2058_n 0.00246676f $X=11.43 $Y=0.37 $X2=0
+ $Y2=0
cc_1117 N_A_1191_121#_c_1700_n N_VGND_c_2058_n 0.00678664f $X=6.1 $Y=0.75 $X2=0
+ $Y2=0
cc_1118 N_A_1191_121#_c_1705_n N_VGND_c_2058_n 0.00660921f $X=10.885 $Y=0.34
+ $X2=0 $Y2=0
cc_1119 N_A_1191_121#_c_1706_n N_VGND_c_2058_n 0.0342794f $X=11.65 $Y=0.34 $X2=0
+ $Y2=0
cc_1120 N_A_1191_121#_c_1727_n N_A_1278_121#_M1002_d 0.00330483f $X=6.875
+ $Y=1.11 $X2=-0.19 $Y2=-0.245
cc_1121 N_A_1191_121#_c_1700_n N_A_1278_121#_c_2324_n 0.0104051f $X=6.1 $Y=0.75
+ $X2=0 $Y2=0
cc_1122 N_A_1191_121#_c_1727_n N_A_1278_121#_c_2324_n 0.0169041f $X=6.875
+ $Y=1.11 $X2=0 $Y2=0
cc_1123 N_A_1191_121#_c_1701_n N_A_1278_121#_c_2324_n 0.00652315f $X=7 $Y=0.765
+ $X2=0 $Y2=0
cc_1124 N_A_1191_121#_c_1727_n N_A_1278_121#_c_2325_n 0.00425327f $X=6.875
+ $Y=1.11 $X2=0 $Y2=0
cc_1125 N_A_1191_121#_c_1701_n N_A_1278_121#_c_2325_n 0.0196444f $X=7 $Y=0.765
+ $X2=0 $Y2=0
cc_1126 N_A_1191_121#_c_1703_n N_A_1278_121#_c_2325_n 0.0422737f $X=7.735
+ $Y=0.68 $X2=0 $Y2=0
cc_1127 N_A_1191_121#_c_1708_n N_A_1278_121#_c_2325_n 0.0185406f $X=7.86 $Y=0.68
+ $X2=0 $Y2=0
cc_1128 N_A_1191_121#_c_1708_n N_A_1278_121#_c_2329_n 0.0125333f $X=7.86 $Y=0.68
+ $X2=0 $Y2=0
cc_1129 N_A_1191_121#_c_1703_n N_A_1450_121#_M1012_d 0.00168086f $X=7.735
+ $Y=0.68 $X2=-0.19 $Y2=-0.245
cc_1130 N_A_1191_121#_M1041_s N_A_1450_121#_c_2377_n 0.00486971f $X=7.68
+ $Y=0.605 $X2=0 $Y2=0
cc_1131 N_A_1191_121#_c_1703_n N_A_1450_121#_c_2377_n 0.00498063f $X=7.735
+ $Y=0.68 $X2=0 $Y2=0
cc_1132 N_A_1191_121#_c_1708_n N_A_1450_121#_c_2377_n 0.0189683f $X=7.86 $Y=0.68
+ $X2=0 $Y2=0
cc_1133 N_A_1191_121#_c_1704_n N_A_1450_121#_c_2378_n 0.00207966f $X=10.8
+ $Y=1.945 $X2=0 $Y2=0
cc_1134 N_A_1191_121#_c_1703_n N_A_1450_121#_c_2380_n 0.0144331f $X=7.735
+ $Y=0.68 $X2=0 $Y2=0
cc_1135 N_A_1191_121#_c_1707_n N_A_1450_121#_c_2380_n 0.00998734f $X=7 $Y=1.145
+ $X2=0 $Y2=0
cc_1136 N_A_1191_121#_c_1708_n N_A_1450_121#_c_2381_n 3.61824e-19 $X=7.86
+ $Y=0.68 $X2=0 $Y2=0
cc_1137 N_A_1288_377#_c_1873_n N_A_1468_377#_M1036_d 0.00402069f $X=9.935
+ $Y=2.71 $X2=0 $Y2=0
cc_1138 N_A_1288_377#_c_1871_n N_A_1468_377#_c_1926_n 0.0106263f $X=7.98 $Y=2.99
+ $X2=0 $Y2=0
cc_1139 N_A_1288_377#_c_1873_n N_A_1468_377#_c_1926_n 0.0601271f $X=9.935
+ $Y=2.71 $X2=0 $Y2=0
cc_1140 N_A_1288_377#_c_1874_n N_A_1468_377#_c_1926_n 0.0129848f $X=8.065
+ $Y=2.71 $X2=0 $Y2=0
cc_1141 N_A_1288_377#_c_1871_n N_A_1468_377#_c_1928_n 0.0199555f $X=7.98 $Y=2.99
+ $X2=0 $Y2=0
cc_1142 N_A_1288_377#_c_1874_n N_A_1468_377#_c_1928_n 0.00476684f $X=8.065
+ $Y=2.71 $X2=0 $Y2=0
cc_1143 N_X_c_1948_n N_VGND_M1027_s 0.00176461f $X=15.925 $Y=1.045 $X2=0 $Y2=0
cc_1144 N_X_c_1951_n N_VGND_M1051_s 0.00338075f $X=16.445 $Y=1.045 $X2=0 $Y2=0
cc_1145 N_X_c_1947_n N_VGND_c_2040_n 0.0216048f $X=15.23 $Y=0.515 $X2=0 $Y2=0
cc_1146 N_X_c_1949_n N_VGND_c_2040_n 0.00752767f $X=15.315 $Y=1.045 $X2=0 $Y2=0
cc_1147 N_X_c_1947_n N_VGND_c_2041_n 0.0158413f $X=15.23 $Y=0.515 $X2=0 $Y2=0
cc_1148 N_X_c_1948_n N_VGND_c_2041_n 0.0152916f $X=15.925 $Y=1.045 $X2=0 $Y2=0
cc_1149 N_X_c_1950_n N_VGND_c_2041_n 0.0158413f $X=16.09 $Y=0.515 $X2=0 $Y2=0
cc_1150 N_X_c_1950_n N_VGND_c_2043_n 0.0164981f $X=16.09 $Y=0.515 $X2=0 $Y2=0
cc_1151 N_X_c_1951_n N_VGND_c_2043_n 0.023173f $X=16.445 $Y=1.045 $X2=0 $Y2=0
cc_1152 N_X_c_1947_n N_VGND_c_2052_n 0.0109942f $X=15.23 $Y=0.515 $X2=0 $Y2=0
cc_1153 N_X_c_1950_n N_VGND_c_2053_n 0.0109942f $X=16.09 $Y=0.515 $X2=0 $Y2=0
cc_1154 N_X_c_1947_n N_VGND_c_2058_n 0.00904371f $X=15.23 $Y=0.515 $X2=0 $Y2=0
cc_1155 N_X_c_1950_n N_VGND_c_2058_n 0.00904371f $X=16.09 $Y=0.515 $X2=0 $Y2=0
cc_1156 N_VGND_c_2033_n N_A_114_126#_M1025_s 0.00178571f $X=1.045 $Y=1.155
+ $X2=-0.19 $Y2=-0.245
cc_1157 N_VGND_c_2032_n N_A_114_126#_c_2232_n 0.0201555f $X=0.28 $Y=0.775 $X2=0
+ $Y2=0
cc_1158 N_VGND_c_2033_n N_A_114_126#_c_2232_n 0.0173292f $X=1.045 $Y=1.155 $X2=0
+ $Y2=0
cc_1159 N_VGND_c_2033_n N_A_114_126#_c_2233_n 0.00448545f $X=1.045 $Y=1.155
+ $X2=0 $Y2=0
cc_1160 N_VGND_c_2072_n N_A_114_126#_c_2233_n 0.022569f $X=1.17 $Y=0.805 $X2=0
+ $Y2=0
cc_1161 N_VGND_c_2035_n N_A_114_126#_c_2233_n 0.0154808f $X=2.145 $Y=0.365 $X2=0
+ $Y2=0
cc_1162 N_VGND_c_2050_n N_A_114_126#_c_2233_n 0.0550594f $X=1.98 $Y=0 $X2=0
+ $Y2=0
cc_1163 N_VGND_c_2058_n N_A_114_126#_c_2233_n 0.0350536f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1164 N_VGND_c_2032_n N_A_114_126#_c_2234_n 0.0162425f $X=0.28 $Y=0.775 $X2=0
+ $Y2=0
cc_1165 N_VGND_c_2050_n N_A_114_126#_c_2234_n 0.0207641f $X=1.98 $Y=0 $X2=0
+ $Y2=0
cc_1166 N_VGND_c_2058_n N_A_114_126#_c_2234_n 0.0126529f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1167 N_VGND_M1023_s N_A_114_126#_c_2236_n 0.0111424f $X=1.925 $Y=0.63 $X2=0
+ $Y2=0
cc_1168 N_VGND_c_2072_n N_A_114_126#_c_2236_n 0.0105495f $X=1.17 $Y=0.805 $X2=0
+ $Y2=0
cc_1169 N_VGND_c_2035_n N_A_114_126#_c_2236_n 0.0127545f $X=2.145 $Y=0.365 $X2=0
+ $Y2=0
cc_1170 N_VGND_c_2050_n N_A_114_126#_c_2236_n 0.00298933f $X=1.98 $Y=0 $X2=0
+ $Y2=0
cc_1171 N_VGND_c_2058_n N_A_114_126#_c_2236_n 0.00562944f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1172 N_VGND_M1023_s N_A_114_126#_c_2237_n 0.00425076f $X=1.925 $Y=0.63 $X2=0
+ $Y2=0
cc_1173 N_VGND_c_2035_n N_A_114_126#_c_2237_n 0.00511893f $X=2.145 $Y=0.365
+ $X2=0 $Y2=0
cc_1174 N_VGND_c_2058_n N_A_114_126#_c_2237_n 0.00983818f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1175 N_VGND_M1023_s N_A_299_126#_c_2282_n 0.00470132f $X=1.925 $Y=0.63 $X2=0
+ $Y2=0
cc_1176 N_VGND_c_2034_n N_A_299_126#_c_2285_n 0.0104027f $X=1.207 $Y=1.03 $X2=0
+ $Y2=0
cc_1177 N_VGND_c_2036_n N_A_1278_121#_c_2324_n 0.00470266f $X=5.54 $Y=0.515
+ $X2=0 $Y2=0
cc_1178 N_VGND_c_2044_n N_A_1278_121#_c_2325_n 0.0137091f $X=8.66 $Y=0 $X2=0
+ $Y2=0
cc_1179 N_VGND_c_2045_n N_A_1278_121#_c_2325_n 0.105357f $X=8.495 $Y=0 $X2=0
+ $Y2=0
cc_1180 N_VGND_c_2058_n N_A_1278_121#_c_2325_n 0.054907f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1181 N_VGND_c_2036_n N_A_1278_121#_c_2326_n 0.00581676f $X=5.54 $Y=0.515
+ $X2=0 $Y2=0
cc_1182 N_VGND_c_2045_n N_A_1278_121#_c_2326_n 0.0222946f $X=8.495 $Y=0 $X2=0
+ $Y2=0
cc_1183 N_VGND_c_2058_n N_A_1278_121#_c_2326_n 0.0112784f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1184 N_VGND_M1021_s N_A_1278_121#_c_2328_n 0.00797645f $X=8.515 $Y=0.18 $X2=0
+ $Y2=0
cc_1185 N_VGND_c_2044_n N_A_1278_121#_c_2328_n 0.0245264f $X=8.66 $Y=0 $X2=0
+ $Y2=0
cc_1186 N_VGND_c_2045_n N_A_1278_121#_c_2328_n 0.0034901f $X=8.495 $Y=0 $X2=0
+ $Y2=0
cc_1187 N_VGND_c_2046_n N_A_1278_121#_c_2328_n 0.0029521f $X=9.435 $Y=0 $X2=0
+ $Y2=0
cc_1188 N_VGND_c_2058_n N_A_1278_121#_c_2328_n 0.0115245f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1189 N_VGND_c_2037_n N_A_1278_121#_c_2330_n 0.0144673f $X=9.6 $Y=0.55 $X2=0
+ $Y2=0
cc_1190 N_VGND_c_2044_n N_A_1278_121#_c_2330_n 0.00282013f $X=8.66 $Y=0 $X2=0
+ $Y2=0
cc_1191 N_VGND_c_2046_n N_A_1278_121#_c_2330_n 0.0105866f $X=9.435 $Y=0 $X2=0
+ $Y2=0
cc_1192 N_VGND_c_2058_n N_A_1278_121#_c_2330_n 0.00888607f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1193 N_VGND_M1021_s N_A_1450_121#_c_2378_n 0.00419342f $X=8.515 $Y=0.18 $X2=0
+ $Y2=0
cc_1194 N_VGND_M1040_s N_A_1450_121#_c_2378_n 0.00176461f $X=9.46 $Y=0.37 $X2=0
+ $Y2=0
cc_1195 N_VGND_c_2037_n N_A_1450_121#_c_2378_n 0.0153337f $X=9.6 $Y=0.55 $X2=0
+ $Y2=0
cc_1196 N_VGND_c_2039_n N_A_1450_121#_c_2378_n 0.00464574f $X=10.46 $Y=0.515
+ $X2=0 $Y2=0
cc_1197 N_VGND_c_2037_n N_A_1450_121#_c_2379_n 0.0144673f $X=9.6 $Y=0.55 $X2=0
+ $Y2=0
cc_1198 N_VGND_c_2038_n N_A_1450_121#_c_2379_n 0.0109942f $X=10.295 $Y=0 $X2=0
+ $Y2=0
cc_1199 N_VGND_c_2039_n N_A_1450_121#_c_2379_n 0.0203066f $X=10.46 $Y=0.515
+ $X2=0 $Y2=0
cc_1200 N_VGND_c_2058_n N_A_1450_121#_c_2379_n 0.00904371f $X=16.56 $Y=0 $X2=0
+ $Y2=0
cc_1201 N_A_114_126#_c_2236_n N_A_299_126#_M1022_d 0.00316283f $X=2.14 $Y=0.875
+ $X2=-0.19 $Y2=-0.245
cc_1202 N_A_114_126#_c_2236_n N_A_299_126#_c_2282_n 0.0170749f $X=2.14 $Y=0.875
+ $X2=0 $Y2=0
cc_1203 N_A_114_126#_c_2237_n N_A_299_126#_c_2282_n 0.0289644f $X=3.05 $Y=0.842
+ $X2=0 $Y2=0
cc_1204 N_A_114_126#_c_2247_n N_A_299_126#_c_2283_n 0.0223181f $X=3.215 $Y=0.84
+ $X2=0 $Y2=0
cc_1205 N_A_114_126#_c_2237_n N_A_299_126#_c_2283_n 0.0155869f $X=3.05 $Y=0.842
+ $X2=0 $Y2=0
cc_1206 N_A_114_126#_c_2233_n N_A_299_126#_c_2285_n 8.50133e-19 $X=1.575
+ $Y=0.372 $X2=0 $Y2=0
cc_1207 N_A_114_126#_c_2236_n N_A_299_126#_c_2285_n 0.0138528f $X=2.14 $Y=0.875
+ $X2=0 $Y2=0
cc_1208 N_A_114_126#_c_2237_n N_A_299_126#_c_2286_n 0.0129027f $X=3.05 $Y=0.842
+ $X2=0 $Y2=0
cc_1209 N_A_1278_121#_c_2325_n N_A_1450_121#_c_2377_n 0.00484741f $X=8.155
+ $Y=0.34 $X2=0 $Y2=0
cc_1210 N_A_1278_121#_M1021_d N_A_1450_121#_c_2378_n 0.00176461f $X=9.03 $Y=0.37
+ $X2=0 $Y2=0
cc_1211 N_A_1278_121#_c_2328_n N_A_1450_121#_c_2378_n 0.0451131f $X=9.005
+ $Y=0.665 $X2=0 $Y2=0
cc_1212 N_A_1278_121#_c_2330_n N_A_1450_121#_c_2378_n 0.0146914f $X=9.17 $Y=0.55
+ $X2=0 $Y2=0
cc_1213 N_A_1278_121#_c_2329_n N_A_1450_121#_c_2381_n 0.0133492f $X=8.325
+ $Y=0.665 $X2=0 $Y2=0

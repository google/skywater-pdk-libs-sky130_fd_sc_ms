* File: sky130_fd_sc_ms__a31o_2.pxi.spice
* Created: Wed Sep  2 11:55:08 2020
* 
x_PM_SKY130_FD_SC_MS__A31O_2%A_97_296# N_A_97_296#_M1011_d N_A_97_296#_M1010_d
+ N_A_97_296#_M1002_g N_A_97_296#_M1007_g N_A_97_296#_M1008_g
+ N_A_97_296#_M1003_g N_A_97_296#_c_65_n N_A_97_296#_c_79_p N_A_97_296#_c_153_p
+ N_A_97_296#_c_71_n N_A_97_296#_c_102_p N_A_97_296#_c_66_n N_A_97_296#_c_72_n
+ N_A_97_296#_c_67_n N_A_97_296#_c_68_n PM_SKY130_FD_SC_MS__A31O_2%A_97_296#
x_PM_SKY130_FD_SC_MS__A31O_2%A3 N_A3_M1004_g N_A3_M1001_g A3 N_A3_c_173_n
+ N_A3_c_174_n PM_SKY130_FD_SC_MS__A31O_2%A3
x_PM_SKY130_FD_SC_MS__A31O_2%A2 N_A2_M1006_g N_A2_M1005_g A2 N_A2_c_208_n
+ N_A2_c_209_n N_A2_c_210_n PM_SKY130_FD_SC_MS__A31O_2%A2
x_PM_SKY130_FD_SC_MS__A31O_2%A1 N_A1_M1011_g N_A1_M1009_g A1 N_A1_c_241_n
+ N_A1_c_242_n PM_SKY130_FD_SC_MS__A31O_2%A1
x_PM_SKY130_FD_SC_MS__A31O_2%B1 N_B1_c_274_n N_B1_M1000_g N_B1_M1010_g B1
+ N_B1_c_277_n PM_SKY130_FD_SC_MS__A31O_2%B1
x_PM_SKY130_FD_SC_MS__A31O_2%VPWR N_VPWR_M1002_s N_VPWR_M1003_s N_VPWR_M1005_d
+ N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_302_n VPWR
+ N_VPWR_c_303_n N_VPWR_c_304_n N_VPWR_c_305_n N_VPWR_c_298_n N_VPWR_c_307_n
+ N_VPWR_c_308_n PM_SKY130_FD_SC_MS__A31O_2%VPWR
x_PM_SKY130_FD_SC_MS__A31O_2%X N_X_M1007_s N_X_M1002_d N_X_c_348_n N_X_c_349_n X
+ X X X N_X_c_350_n PM_SKY130_FD_SC_MS__A31O_2%X
x_PM_SKY130_FD_SC_MS__A31O_2%A_365_368# N_A_365_368#_M1004_d
+ N_A_365_368#_M1009_d N_A_365_368#_c_383_n N_A_365_368#_c_379_n
+ N_A_365_368#_c_380_n PM_SKY130_FD_SC_MS__A31O_2%A_365_368#
x_PM_SKY130_FD_SC_MS__A31O_2%VGND N_VGND_M1007_d N_VGND_M1008_d N_VGND_M1000_d
+ N_VGND_c_405_n N_VGND_c_406_n N_VGND_c_407_n N_VGND_c_408_n VGND
+ N_VGND_c_409_n N_VGND_c_410_n N_VGND_c_411_n N_VGND_c_412_n
+ PM_SKY130_FD_SC_MS__A31O_2%VGND
cc_1 VNB N_A_97_296#_M1002_g 0.00231818f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.4
cc_2 VNB N_A_97_296#_M1007_g 0.0260123f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_3 VNB N_A_97_296#_M1008_g 0.0235682f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_4 VNB N_A_97_296#_M1003_g 0.00180134f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=2.4
cc_5 VNB N_A_97_296#_c_65_n 0.00317249f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=1.3
cc_6 VNB N_A_97_296#_c_66_n 0.00335352f $X=-0.19 $Y=-0.245 $X2=3.015 $Y2=0.495
cc_7 VNB N_A_97_296#_c_67_n 0.00590395f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=1.465
cc_8 VNB N_A_97_296#_c_68_n 0.0665637f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.465
cc_9 VNB N_A3_M1004_g 0.00668438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB A3 0.00334701f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.4
cc_11 VNB N_A3_c_173_n 0.0332288f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.3
cc_12 VNB N_A3_c_174_n 0.0188039f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_13 VNB N_A2_M1005_g 0.00691403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_208_n 0.0279589f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.3
cc_15 VNB N_A2_c_209_n 0.00752993f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_16 VNB N_A2_c_210_n 0.0183498f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_17 VNB N_A1_M1009_g 0.00711974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB A1 0.0109964f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.4
cc_19 VNB N_A1_c_241_n 0.0280958f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.3
cc_20 VNB N_A1_c_242_n 0.0198831f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_21 VNB N_B1_c_274_n 0.0220404f $X=-0.19 $Y=-0.245 $X2=2.815 $Y2=0.37
cc_22 VNB N_B1_M1010_g 0.00957504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB B1 0.00926001f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.4
cc_24 VNB N_B1_c_277_n 0.0579546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_298_n 0.163682f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=1.465
cc_26 VNB N_X_c_348_n 0.00229096f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.4
cc_27 VNB N_X_c_349_n 0.00306343f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_28 VNB N_X_c_350_n 0.00113823f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=1.89
cc_29 VNB N_VGND_c_405_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_406_n 0.0550278f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_31 VNB N_VGND_c_407_n 0.0131437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_408_n 0.0344105f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_33 VNB N_VGND_c_409_n 0.0172472f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=2.4
cc_34 VNB N_VGND_c_410_n 0.0489588f $X=-0.19 $Y=-0.245 $X2=2.85 $Y2=0.925
cc_35 VNB N_VGND_c_411_n 0.0187802f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=1.985
cc_36 VNB N_VGND_c_412_n 0.228974f $X=-0.19 $Y=-0.245 $X2=3.015 $Y2=0.925
cc_37 VPB N_A_97_296#_M1002_g 0.0273997f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=2.4
cc_38 VPB N_A_97_296#_M1003_g 0.0254398f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=2.4
cc_39 VPB N_A_97_296#_c_71_n 0.0376948f $X=-0.19 $Y=1.66 $X2=3.385 $Y2=1.805
cc_40 VPB N_A_97_296#_c_72_n 0.040239f $X=-0.19 $Y=1.66 $X2=3.555 $Y2=1.985
cc_41 VPB N_A_97_296#_c_67_n 0.00232704f $X=-0.19 $Y=1.66 $X2=1.12 $Y2=1.465
cc_42 VPB N_A3_M1004_g 0.0234322f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A2_M1005_g 0.0229569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A1_M1009_g 0.023553f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_B1_M1010_g 0.028768f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_299_n 0.012885f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_300_n 0.0637942f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_48 VPB N_VPWR_c_301_n 0.0130389f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_302_n 0.0199866f $X=-0.19 $Y=1.66 $X2=1.22 $Y2=1.3
cc_50 VPB N_VPWR_c_303_n 0.0181766f $X=-0.19 $Y=1.66 $X2=1.305 $Y2=1.805
cc_51 VPB N_VPWR_c_304_n 0.0209833f $X=-0.19 $Y=1.66 $X2=3.555 $Y2=1.89
cc_52 VPB N_VPWR_c_305_n 0.034947f $X=-0.19 $Y=1.66 $X2=1.12 $Y2=1.465
cc_53 VPB N_VPWR_c_298_n 0.0797034f $X=-0.19 $Y=1.66 $X2=1.12 $Y2=1.465
cc_54 VPB N_VPWR_c_307_n 0.0100751f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.465
cc_55 VPB N_VPWR_c_308_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB X 0.0038778f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB X 0.00233713f $X=-0.19 $Y=1.66 $X2=1.22 $Y2=1.3
cc_58 VPB N_X_c_350_n 8.38119e-19 $X=-0.19 $Y=1.66 $X2=3.555 $Y2=1.89
cc_59 VPB N_A_365_368#_c_379_n 0.0028233f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_365_368#_c_380_n 0.00331839f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_61 N_A_97_296#_M1003_g N_A3_M1004_g 0.0134217f $X=1.025 $Y=2.4 $X2=0 $Y2=0
cc_62 N_A_97_296#_c_71_n N_A3_M1004_g 0.0171914f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_63 N_A_97_296#_c_67_n N_A3_M1004_g 0.00332609f $X=1.12 $Y=1.465 $X2=0 $Y2=0
cc_64 N_A_97_296#_c_68_n N_A3_M1004_g 0.00243134f $X=1.025 $Y=1.465 $X2=0 $Y2=0
cc_65 N_A_97_296#_c_65_n A3 0.00757247f $X=1.22 $Y=1.3 $X2=0 $Y2=0
cc_66 N_A_97_296#_c_79_p A3 0.0228656f $X=2.85 $Y=0.925 $X2=0 $Y2=0
cc_67 N_A_97_296#_c_71_n A3 0.024317f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_68 N_A_97_296#_c_67_n A3 0.0164597f $X=1.12 $Y=1.465 $X2=0 $Y2=0
cc_69 N_A_97_296#_c_68_n A3 3.04404e-19 $X=1.025 $Y=1.465 $X2=0 $Y2=0
cc_70 N_A_97_296#_M1008_g N_A3_c_173_n 0.00147268f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_71 N_A_97_296#_c_65_n N_A3_c_173_n 6.42308e-19 $X=1.22 $Y=1.3 $X2=0 $Y2=0
cc_72 N_A_97_296#_c_79_p N_A3_c_173_n 0.00100851f $X=2.85 $Y=0.925 $X2=0 $Y2=0
cc_73 N_A_97_296#_c_71_n N_A3_c_173_n 0.00104059f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_74 N_A_97_296#_c_67_n N_A3_c_173_n 0.00153381f $X=1.12 $Y=1.465 $X2=0 $Y2=0
cc_75 N_A_97_296#_c_68_n N_A3_c_173_n 0.0133463f $X=1.025 $Y=1.465 $X2=0 $Y2=0
cc_76 N_A_97_296#_M1008_g N_A3_c_174_n 0.00877705f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_77 N_A_97_296#_c_65_n N_A3_c_174_n 0.00315986f $X=1.22 $Y=1.3 $X2=0 $Y2=0
cc_78 N_A_97_296#_c_79_p N_A3_c_174_n 0.0126481f $X=2.85 $Y=0.925 $X2=0 $Y2=0
cc_79 N_A_97_296#_c_71_n N_A2_M1005_g 0.0124988f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_80 N_A_97_296#_c_79_p N_A2_c_208_n 0.00101866f $X=2.85 $Y=0.925 $X2=0 $Y2=0
cc_81 N_A_97_296#_c_71_n N_A2_c_208_n 0.00336308f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_82 N_A_97_296#_c_79_p N_A2_c_209_n 0.0250213f $X=2.85 $Y=0.925 $X2=0 $Y2=0
cc_83 N_A_97_296#_c_71_n N_A2_c_209_n 0.0283471f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_84 N_A_97_296#_c_79_p N_A2_c_210_n 0.0122562f $X=2.85 $Y=0.925 $X2=0 $Y2=0
cc_85 N_A_97_296#_c_71_n N_A1_M1009_g 0.0127848f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_86 N_A_97_296#_c_72_n N_A1_M1009_g 8.56666e-19 $X=3.555 $Y=1.985 $X2=0 $Y2=0
cc_87 N_A_97_296#_c_79_p A1 0.012294f $X=2.85 $Y=0.925 $X2=0 $Y2=0
cc_88 N_A_97_296#_c_71_n A1 0.0435494f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_89 N_A_97_296#_c_102_p A1 0.0277108f $X=3.015 $Y=0.84 $X2=0 $Y2=0
cc_90 N_A_97_296#_c_71_n N_A1_c_241_n 0.00363888f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_91 N_A_97_296#_c_102_p N_A1_c_241_n 9.57669e-19 $X=3.015 $Y=0.84 $X2=0 $Y2=0
cc_92 N_A_97_296#_c_79_p N_A1_c_242_n 0.012933f $X=2.85 $Y=0.925 $X2=0 $Y2=0
cc_93 N_A_97_296#_c_66_n N_A1_c_242_n 0.00348158f $X=3.015 $Y=0.495 $X2=0 $Y2=0
cc_94 N_A_97_296#_c_66_n N_B1_c_274_n 0.00298143f $X=3.015 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_95 N_A_97_296#_c_71_n N_B1_M1010_g 0.0217728f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_96 N_A_97_296#_c_72_n N_B1_M1010_g 0.0131289f $X=3.555 $Y=1.985 $X2=0 $Y2=0
cc_97 N_A_97_296#_c_71_n B1 0.0272055f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_98 N_A_97_296#_c_71_n N_B1_c_277_n 0.00245357f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_99 N_A_97_296#_c_71_n N_VPWR_M1003_s 0.00342895f $X=3.385 $Y=1.805 $X2=0
+ $Y2=0
cc_100 N_A_97_296#_c_67_n N_VPWR_M1003_s 0.00177236f $X=1.12 $Y=1.465 $X2=0
+ $Y2=0
cc_101 N_A_97_296#_c_71_n N_VPWR_M1005_d 0.00395823f $X=3.385 $Y=1.805 $X2=0
+ $Y2=0
cc_102 N_A_97_296#_M1002_g N_VPWR_c_300_n 0.00516118f $X=0.575 $Y=2.4 $X2=0
+ $Y2=0
cc_103 N_A_97_296#_M1002_g N_VPWR_c_301_n 6.03e-19 $X=0.575 $Y=2.4 $X2=0 $Y2=0
cc_104 N_A_97_296#_M1003_g N_VPWR_c_301_n 0.0213519f $X=1.025 $Y=2.4 $X2=0 $Y2=0
cc_105 N_A_97_296#_c_71_n N_VPWR_c_301_n 0.022988f $X=3.385 $Y=1.805 $X2=0 $Y2=0
cc_106 N_A_97_296#_c_67_n N_VPWR_c_301_n 0.0132323f $X=1.12 $Y=1.465 $X2=0 $Y2=0
cc_107 N_A_97_296#_c_68_n N_VPWR_c_301_n 5.99168e-19 $X=1.025 $Y=1.465 $X2=0
+ $Y2=0
cc_108 N_A_97_296#_M1002_g N_VPWR_c_303_n 0.0048691f $X=0.575 $Y=2.4 $X2=0 $Y2=0
cc_109 N_A_97_296#_M1003_g N_VPWR_c_303_n 0.00475445f $X=1.025 $Y=2.4 $X2=0
+ $Y2=0
cc_110 N_A_97_296#_c_72_n N_VPWR_c_305_n 0.0100594f $X=3.555 $Y=1.985 $X2=0
+ $Y2=0
cc_111 N_A_97_296#_M1002_g N_VPWR_c_298_n 0.00876167f $X=0.575 $Y=2.4 $X2=0
+ $Y2=0
cc_112 N_A_97_296#_M1003_g N_VPWR_c_298_n 0.00938661f $X=1.025 $Y=2.4 $X2=0
+ $Y2=0
cc_113 N_A_97_296#_c_72_n N_VPWR_c_298_n 0.0115169f $X=3.555 $Y=1.985 $X2=0
+ $Y2=0
cc_114 N_A_97_296#_M1007_g N_X_c_348_n 0.0078359f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_115 N_A_97_296#_M1008_g N_X_c_348_n 5.92016e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A_97_296#_M1007_g N_X_c_349_n 0.00164237f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_117 N_A_97_296#_c_65_n N_X_c_349_n 0.00392342f $X=1.22 $Y=1.3 $X2=0 $Y2=0
cc_118 N_A_97_296#_c_68_n N_X_c_349_n 0.00199986f $X=1.025 $Y=1.465 $X2=0 $Y2=0
cc_119 N_A_97_296#_M1002_g X 0.0028171f $X=0.575 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A_97_296#_M1003_g X 5.63769e-19 $X=1.025 $Y=2.4 $X2=0 $Y2=0
cc_121 N_A_97_296#_c_67_n X 0.00141813f $X=1.12 $Y=1.465 $X2=0 $Y2=0
cc_122 N_A_97_296#_c_68_n X 0.00266746f $X=1.025 $Y=1.465 $X2=0 $Y2=0
cc_123 N_A_97_296#_M1002_g X 0.0150828f $X=0.575 $Y=2.4 $X2=0 $Y2=0
cc_124 N_A_97_296#_M1002_g N_X_c_350_n 0.00982755f $X=0.575 $Y=2.4 $X2=0 $Y2=0
cc_125 N_A_97_296#_M1007_g N_X_c_350_n 0.00856132f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A_97_296#_M1008_g N_X_c_350_n 9.64425e-19 $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A_97_296#_M1003_g N_X_c_350_n 0.00109596f $X=1.025 $Y=2.4 $X2=0 $Y2=0
cc_128 N_A_97_296#_c_65_n N_X_c_350_n 0.00544148f $X=1.22 $Y=1.3 $X2=0 $Y2=0
cc_129 N_A_97_296#_c_67_n N_X_c_350_n 0.0304594f $X=1.12 $Y=1.465 $X2=0 $Y2=0
cc_130 N_A_97_296#_c_68_n N_X_c_350_n 0.0243631f $X=1.025 $Y=1.465 $X2=0 $Y2=0
cc_131 N_A_97_296#_c_71_n N_A_365_368#_M1004_d 0.00165831f $X=3.385 $Y=1.805
+ $X2=-0.19 $Y2=-0.245
cc_132 N_A_97_296#_c_71_n N_A_365_368#_M1009_d 0.00218982f $X=3.385 $Y=1.805
+ $X2=0 $Y2=0
cc_133 N_A_97_296#_c_71_n N_A_365_368#_c_383_n 0.0453975f $X=3.385 $Y=1.805
+ $X2=0 $Y2=0
cc_134 N_A_97_296#_M1003_g N_A_365_368#_c_379_n 2.1828e-19 $X=1.025 $Y=2.4 $X2=0
+ $Y2=0
cc_135 N_A_97_296#_c_71_n N_A_365_368#_c_379_n 0.0171782f $X=3.385 $Y=1.805
+ $X2=0 $Y2=0
cc_136 N_A_97_296#_c_71_n N_A_365_368#_c_380_n 0.019003f $X=3.385 $Y=1.805 $X2=0
+ $Y2=0
cc_137 N_A_97_296#_c_72_n N_A_365_368#_c_380_n 0.0245379f $X=3.555 $Y=1.985
+ $X2=0 $Y2=0
cc_138 N_A_97_296#_c_65_n N_VGND_M1008_d 0.00324595f $X=1.22 $Y=1.3 $X2=0 $Y2=0
cc_139 N_A_97_296#_c_79_p N_VGND_M1008_d 0.0156289f $X=2.85 $Y=0.925 $X2=0 $Y2=0
cc_140 N_A_97_296#_c_153_p N_VGND_M1008_d 0.00542593f $X=1.305 $Y=0.925 $X2=0
+ $Y2=0
cc_141 N_A_97_296#_M1007_g N_VGND_c_406_n 0.0184209f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_142 N_A_97_296#_c_66_n N_VGND_c_408_n 0.0183215f $X=3.015 $Y=0.495 $X2=0
+ $Y2=0
cc_143 N_A_97_296#_M1007_g N_VGND_c_409_n 0.00434272f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_144 N_A_97_296#_M1008_g N_VGND_c_409_n 0.004307f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A_97_296#_c_66_n N_VGND_c_410_n 0.0146038f $X=3.015 $Y=0.495 $X2=0
+ $Y2=0
cc_146 N_A_97_296#_M1007_g N_VGND_c_411_n 4.01823e-19 $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_147 N_A_97_296#_M1008_g N_VGND_c_411_n 0.00736755f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_148 N_A_97_296#_c_79_p N_VGND_c_411_n 0.021742f $X=2.85 $Y=0.925 $X2=0 $Y2=0
cc_149 N_A_97_296#_c_153_p N_VGND_c_411_n 0.0111679f $X=1.305 $Y=0.925 $X2=0
+ $Y2=0
cc_150 N_A_97_296#_c_68_n N_VGND_c_411_n 7.08609e-19 $X=1.025 $Y=1.465 $X2=0
+ $Y2=0
cc_151 N_A_97_296#_M1007_g N_VGND_c_412_n 0.00823934f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_152 N_A_97_296#_M1008_g N_VGND_c_412_n 0.00847524f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_153 N_A_97_296#_c_79_p N_VGND_c_412_n 0.0372445f $X=2.85 $Y=0.925 $X2=0 $Y2=0
cc_154 N_A_97_296#_c_153_p N_VGND_c_412_n 7.38843e-19 $X=1.305 $Y=0.925 $X2=0
+ $Y2=0
cc_155 N_A_97_296#_c_66_n N_VGND_c_412_n 0.0121018f $X=3.015 $Y=0.495 $X2=0
+ $Y2=0
cc_156 N_A_97_296#_c_79_p A_371_74# 0.00734082f $X=2.85 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_157 N_A_97_296#_c_79_p A_449_74# 0.0147367f $X=2.85 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_158 N_A3_M1004_g N_A2_M1005_g 0.0339866f $X=1.735 $Y=2.34 $X2=0 $Y2=0
cc_159 N_A3_c_173_n N_A2_c_208_n 0.0359536f $X=1.69 $Y=1.385 $X2=0 $Y2=0
cc_160 A3 N_A2_c_209_n 0.0271823f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_161 N_A3_c_174_n N_A2_c_209_n 0.00224187f $X=1.69 $Y=1.22 $X2=0 $Y2=0
cc_162 A3 N_A2_c_210_n 4.24429e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_163 N_A3_c_174_n N_A2_c_210_n 0.0359536f $X=1.69 $Y=1.22 $X2=0 $Y2=0
cc_164 N_A3_M1004_g N_VPWR_c_301_n 0.00716894f $X=1.735 $Y=2.34 $X2=0 $Y2=0
cc_165 N_A3_M1004_g N_VPWR_c_304_n 0.00567889f $X=1.735 $Y=2.34 $X2=0 $Y2=0
cc_166 N_A3_M1004_g N_VPWR_c_298_n 0.00610055f $X=1.735 $Y=2.34 $X2=0 $Y2=0
cc_167 N_A3_M1004_g N_A_365_368#_c_379_n 0.0118817f $X=1.735 $Y=2.34 $X2=0 $Y2=0
cc_168 N_A3_c_174_n N_VGND_c_410_n 0.00384553f $X=1.69 $Y=1.22 $X2=0 $Y2=0
cc_169 N_A3_c_174_n N_VGND_c_411_n 0.0103313f $X=1.69 $Y=1.22 $X2=0 $Y2=0
cc_170 N_A3_c_174_n N_VGND_c_412_n 0.00383677f $X=1.69 $Y=1.22 $X2=0 $Y2=0
cc_171 N_A2_M1005_g N_A1_M1009_g 0.0325142f $X=2.185 $Y=2.34 $X2=0 $Y2=0
cc_172 N_A2_c_208_n A1 4.18553e-19 $X=2.26 $Y=1.385 $X2=0 $Y2=0
cc_173 N_A2_c_209_n A1 0.0224075f $X=2.26 $Y=1.385 $X2=0 $Y2=0
cc_174 N_A2_c_208_n N_A1_c_241_n 0.0181621f $X=2.26 $Y=1.385 $X2=0 $Y2=0
cc_175 N_A2_c_209_n N_A1_c_241_n 4.20673e-19 $X=2.26 $Y=1.385 $X2=0 $Y2=0
cc_176 N_A2_c_210_n N_A1_c_242_n 0.0301845f $X=2.26 $Y=1.22 $X2=0 $Y2=0
cc_177 N_A2_M1005_g N_VPWR_c_302_n 0.00796671f $X=2.185 $Y=2.34 $X2=0 $Y2=0
cc_178 N_A2_M1005_g N_VPWR_c_304_n 0.00567889f $X=2.185 $Y=2.34 $X2=0 $Y2=0
cc_179 N_A2_M1005_g N_VPWR_c_298_n 0.00610055f $X=2.185 $Y=2.34 $X2=0 $Y2=0
cc_180 N_A2_M1005_g N_A_365_368#_c_383_n 0.0138062f $X=2.185 $Y=2.34 $X2=0 $Y2=0
cc_181 N_A2_M1005_g N_A_365_368#_c_379_n 0.0127267f $X=2.185 $Y=2.34 $X2=0 $Y2=0
cc_182 N_A2_M1005_g N_A_365_368#_c_380_n 8.38761e-19 $X=2.185 $Y=2.34 $X2=0
+ $Y2=0
cc_183 N_A2_c_210_n N_VGND_c_410_n 0.00461464f $X=2.26 $Y=1.22 $X2=0 $Y2=0
cc_184 N_A2_c_210_n N_VGND_c_411_n 0.00178416f $X=2.26 $Y=1.22 $X2=0 $Y2=0
cc_185 N_A2_c_210_n N_VGND_c_412_n 0.00465551f $X=2.26 $Y=1.22 $X2=0 $Y2=0
cc_186 A1 N_B1_c_274_n 0.00355487f $X=3.035 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_187 N_A1_c_242_n N_B1_c_274_n 0.0234037f $X=2.83 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_188 N_A1_M1009_g N_B1_M1010_g 0.0276124f $X=2.825 $Y=2.34 $X2=0 $Y2=0
cc_189 A1 B1 0.0290828f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_190 N_A1_c_241_n B1 2.16754e-19 $X=2.83 $Y=1.385 $X2=0 $Y2=0
cc_191 N_A1_c_241_n N_B1_c_277_n 0.0182029f $X=2.83 $Y=1.385 $X2=0 $Y2=0
cc_192 N_A1_M1009_g N_VPWR_c_302_n 0.00640175f $X=2.825 $Y=2.34 $X2=0 $Y2=0
cc_193 N_A1_M1009_g N_VPWR_c_305_n 0.00567889f $X=2.825 $Y=2.34 $X2=0 $Y2=0
cc_194 N_A1_M1009_g N_VPWR_c_298_n 0.00610055f $X=2.825 $Y=2.34 $X2=0 $Y2=0
cc_195 N_A1_M1009_g N_A_365_368#_c_383_n 0.0138062f $X=2.825 $Y=2.34 $X2=0 $Y2=0
cc_196 N_A1_M1009_g N_A_365_368#_c_379_n 8.47283e-19 $X=2.825 $Y=2.34 $X2=0
+ $Y2=0
cc_197 N_A1_M1009_g N_A_365_368#_c_380_n 0.0123814f $X=2.825 $Y=2.34 $X2=0 $Y2=0
cc_198 N_A1_c_242_n N_VGND_c_408_n 7.29208e-19 $X=2.83 $Y=1.22 $X2=0 $Y2=0
cc_199 N_A1_c_242_n N_VGND_c_410_n 0.00461464f $X=2.83 $Y=1.22 $X2=0 $Y2=0
cc_200 N_A1_c_242_n N_VGND_c_412_n 0.00467093f $X=2.83 $Y=1.22 $X2=0 $Y2=0
cc_201 N_B1_M1010_g N_VPWR_c_305_n 0.00567889f $X=3.325 $Y=2.34 $X2=0 $Y2=0
cc_202 N_B1_M1010_g N_VPWR_c_298_n 0.00610055f $X=3.325 $Y=2.34 $X2=0 $Y2=0
cc_203 N_B1_M1010_g N_A_365_368#_c_380_n 8.87887e-19 $X=3.325 $Y=2.34 $X2=0
+ $Y2=0
cc_204 N_B1_c_274_n N_VGND_c_408_n 0.0134916f $X=3.31 $Y=1.22 $X2=0 $Y2=0
cc_205 B1 N_VGND_c_408_n 0.0232669f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_206 N_B1_c_277_n N_VGND_c_408_n 0.00190792f $X=3.57 $Y=1.385 $X2=0 $Y2=0
cc_207 N_B1_c_274_n N_VGND_c_410_n 0.00383152f $X=3.31 $Y=1.22 $X2=0 $Y2=0
cc_208 N_B1_c_274_n N_VGND_c_412_n 0.00758792f $X=3.31 $Y=1.22 $X2=0 $Y2=0
cc_209 N_VPWR_c_300_n X 0.0446957f $X=0.35 $Y=1.985 $X2=0 $Y2=0
cc_210 N_VPWR_c_301_n X 0.0379525f $X=1.255 $Y=2.145 $X2=0 $Y2=0
cc_211 N_VPWR_c_303_n X 0.01379f $X=1.09 $Y=3.33 $X2=0 $Y2=0
cc_212 N_VPWR_c_298_n X 0.0112756f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_213 N_VPWR_M1005_d N_A_365_368#_c_383_n 0.00869539f $X=2.275 $Y=1.84 $X2=0
+ $Y2=0
cc_214 N_VPWR_c_302_n N_A_365_368#_c_383_n 0.0266042f $X=2.515 $Y=2.565 $X2=0
+ $Y2=0
cc_215 N_VPWR_c_301_n N_A_365_368#_c_379_n 0.0244519f $X=1.255 $Y=2.145 $X2=0
+ $Y2=0
cc_216 N_VPWR_c_302_n N_A_365_368#_c_379_n 0.0288221f $X=2.515 $Y=2.565 $X2=0
+ $Y2=0
cc_217 N_VPWR_c_304_n N_A_365_368#_c_379_n 0.00968502f $X=2.35 $Y=3.33 $X2=0
+ $Y2=0
cc_218 N_VPWR_c_298_n N_A_365_368#_c_379_n 0.0111457f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_219 N_VPWR_c_302_n N_A_365_368#_c_380_n 0.015552f $X=2.515 $Y=2.565 $X2=0
+ $Y2=0
cc_220 N_VPWR_c_305_n N_A_365_368#_c_380_n 0.00975961f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_221 N_VPWR_c_298_n N_A_365_368#_c_380_n 0.0111753f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_222 N_X_c_348_n N_VGND_c_406_n 0.0300058f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_223 N_X_c_348_n N_VGND_c_409_n 0.0121098f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_224 N_X_c_348_n N_VGND_c_411_n 0.0112219f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_225 N_X_c_348_n N_VGND_c_412_n 0.00996704f $X=0.78 $Y=0.515 $X2=0 $Y2=0

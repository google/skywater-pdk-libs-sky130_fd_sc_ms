* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__xor3_2 A B C VGND VNB VPB VPWR X
X0 X a_1198_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 a_416_113# a_440_315# a_83_289# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X2 a_83_289# B a_416_113# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 a_1162_379# C VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X4 a_27_134# a_83_289# VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X5 a_440_315# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 VGND a_1198_424# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_416_113# a_1162_379# a_1198_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X8 a_1162_379# C VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X9 a_416_113# a_440_315# a_27_134# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X10 a_83_289# B a_375_419# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X11 VGND A a_83_289# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X12 a_27_134# B a_416_113# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X13 X a_1198_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 VPWR a_1198_424# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 a_375_419# a_440_315# a_83_289# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X16 a_27_134# a_83_289# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X17 a_1198_424# C a_416_113# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X18 a_440_315# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X19 a_27_134# B a_375_419# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X20 a_375_419# a_440_315# a_27_134# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X21 a_1198_424# C a_375_419# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X22 VPWR A a_83_289# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X23 a_375_419# a_1162_379# a_1198_424# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends

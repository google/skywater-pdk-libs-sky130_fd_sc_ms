* File: sky130_fd_sc_ms__dfrbp_1.pex.spice
* Created: Wed Sep  2 12:02:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DFRBP_1%D 3 7 10 11 12 13 19 22 23
r33 22 24 45.79 $w=4.05e-07 $l=1.65e-07 $layer=POLY_cond $X=0.422 $Y=1.165
+ $X2=0.422 $Y2=1
r34 22 23 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.165 $X2=0.385 $Y2=1.165
r35 19 20 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.845 $X2=0.385 $Y2=1.845
r36 17 22 5.08091 $w=4.05e-07 $l=3.7e-08 $layer=POLY_cond $X=0.422 $Y=1.202
+ $X2=0.422 $Y2=1.165
r37 17 19 88.298 $w=4.05e-07 $l=6.43e-07 $layer=POLY_cond $X=0.422 $Y=1.202
+ $X2=0.422 $Y2=1.845
r38 13 20 5.5434 $w=3.93e-07 $l=1.9e-07 $layer=LI1_cond $X=0.322 $Y=2.035
+ $X2=0.322 $Y2=1.845
r39 12 20 5.25164 $w=3.93e-07 $l=1.8e-07 $layer=LI1_cond $X=0.322 $Y=1.665
+ $X2=0.322 $Y2=1.845
r40 11 12 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=0.322 $Y=1.295
+ $X2=0.322 $Y2=1.665
r41 11 23 3.79285 $w=3.93e-07 $l=1.3e-07 $layer=LI1_cond $X=0.322 $Y=1.295
+ $X2=0.322 $Y2=1.165
r42 9 19 41.6085 $w=4.05e-07 $l=3.03e-07 $layer=POLY_cond $X=0.422 $Y=2.148
+ $X2=0.422 $Y2=1.845
r43 9 10 41.5847 $w=4.05e-07 $l=2.02e-07 $layer=POLY_cond $X=0.422 $Y=2.148
+ $X2=0.422 $Y2=2.35
r44 7 24 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.55 $Y=0.6 $X2=0.55
+ $Y2=1
r45 3 10 155.484 $w=1.8e-07 $l=4e-07 $layer=POLY_cond $X=0.505 $Y=2.75 $X2=0.505
+ $Y2=2.35
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_1%CLK 3 7 8 11 13
c46 8 0 1.864e-19 $X=2.16 $Y=1.665
c47 3 0 1.39129e-19 $X=1.965 $Y=2.495
r48 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.95 $Y=1.61
+ $X2=1.95 $Y2=1.775
r49 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.95 $Y=1.61
+ $X2=1.95 $Y2=1.445
r50 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.95
+ $Y=1.61 $X2=1.95 $Y2=1.61
r51 8 12 5.48608 $w=4.67e-07 $l=2.1e-07 $layer=LI1_cond $X=2.16 $Y=1.545
+ $X2=1.95 $Y2=1.545
r52 7 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.995 $Y=0.965
+ $X2=1.995 $Y2=1.445
r53 3 14 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.965 $Y=2.495
+ $X2=1.965 $Y2=1.775
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_1%A_501_387# 1 2 9 11 14 15 17 18 20 21 22 25
+ 29 31 36 37 40 41 42 44 45 46 49 51 52 54 55 57 62 66
c204 66 0 2.21368e-19 $X=3.415 $Y=1.76
c205 62 0 1.864e-19 $X=2.975 $Y=1.907
c206 57 0 1.65606e-19 $X=2.852 $Y=0.34
c207 51 0 1.08581e-19 $X=6.735 $Y=1.865
c208 46 0 1.02425e-19 $X=6.255 $Y=1.065
c209 42 0 1.61434e-19 $X=4.52 $Y=0.665
c210 9 0 1.76128e-19 $X=3.455 $Y=2.525
r211 65 69 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.415 $Y=1.85
+ $X2=3.415 $Y2=2.015
r212 65 66 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.415 $Y=1.85
+ $X2=3.415 $Y2=1.76
r213 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.415
+ $Y=1.85 $X2=3.415 $Y2=1.85
r214 62 64 11.1833 $w=4.8e-07 $l=4.4e-07 $layer=LI1_cond $X=2.975 $Y=1.907
+ $X2=3.415 $Y2=1.907
r215 60 61 4.526 $w=5.23e-07 $l=8.5e-08 $layer=LI1_cond $X=2.852 $Y=0.72
+ $X2=2.852 $Y2=0.805
r216 57 60 8.65733 $w=5.23e-07 $l=3.8e-07 $layer=LI1_cond $X=2.852 $Y=0.34
+ $X2=2.852 $Y2=0.72
r217 55 76 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.205 $Y=2.03
+ $X2=7.205 $Y2=2.195
r218 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.205
+ $Y=2.03 $X2=7.205 $Y2=2.03
r219 52 54 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=6.82 $Y=2.03
+ $X2=7.205 $Y2=2.03
r220 51 52 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.735 $Y=1.865
+ $X2=6.82 $Y2=2.03
r221 50 51 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.735 $Y=1.23
+ $X2=6.735 $Y2=1.865
r222 49 72 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=6.645 $Y=1.065
+ $X2=6.645 $Y2=1.16
r223 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.645
+ $Y=1.065 $X2=6.645 $Y2=1.065
r224 46 48 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=6.255 $Y=1.065
+ $X2=6.645 $Y2=1.065
r225 45 50 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.65 $Y=1.065
+ $X2=6.735 $Y2=1.23
r226 45 48 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=6.65 $Y=1.065
+ $X2=6.645 $Y2=1.065
r227 44 46 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.17 $Y=0.9
+ $X2=6.255 $Y2=1.065
r228 43 44 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=6.17 $Y=0.75
+ $X2=6.17 $Y2=0.9
r229 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.085 $Y=0.665
+ $X2=6.17 $Y2=0.75
r230 41 42 102.102 $w=1.68e-07 $l=1.565e-06 $layer=LI1_cond $X=6.085 $Y=0.665
+ $X2=4.52 $Y2=0.665
r231 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.435 $Y=0.58
+ $X2=4.52 $Y2=0.665
r232 39 40 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.435 $Y=0.425
+ $X2=4.435 $Y2=0.58
r233 38 57 7.46409 $w=1.7e-07 $l=2.63e-07 $layer=LI1_cond $X=3.115 $Y=0.34
+ $X2=2.852 $Y2=0.34
r234 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.35 $Y=0.34
+ $X2=4.435 $Y2=0.425
r235 37 38 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=4.35 $Y=0.34
+ $X2=3.115 $Y2=0.34
r236 36 62 3.8908 $w=2.8e-07 $l=3.32e-07 $layer=LI1_cond $X=2.975 $Y=1.575
+ $X2=2.975 $Y2=1.907
r237 36 61 31.6922 $w=2.78e-07 $l=7.7e-07 $layer=LI1_cond $X=2.975 $Y=1.575
+ $X2=2.975 $Y2=0.805
r238 31 62 6.50234 $w=4.8e-07 $l=2.6163e-07 $layer=LI1_cond $X=2.79 $Y=2.092
+ $X2=2.975 $Y2=1.907
r239 31 33 5.85988 $w=2.93e-07 $l=1.5e-07 $layer=LI1_cond $X=2.79 $Y=2.092
+ $X2=2.64 $Y2=2.092
r240 27 29 56.4043 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=3.975 $Y=1.17
+ $X2=4.085 $Y2=1.17
r241 25 76 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=7.25 $Y=2.565
+ $X2=7.25 $Y2=2.195
r242 21 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.48 $Y=1.16
+ $X2=6.645 $Y2=1.16
r243 21 22 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=6.48 $Y=1.16
+ $X2=6.12 $Y2=1.16
r244 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.045 $Y=1.085
+ $X2=6.12 $Y2=1.16
r245 18 20 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.045 $Y=1.085
+ $X2=6.045 $Y2=0.69
r246 15 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.085 $Y=1.095
+ $X2=4.085 $Y2=1.17
r247 15 17 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.085 $Y=1.095
+ $X2=4.085 $Y2=0.805
r248 13 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.975 $Y=1.245
+ $X2=3.975 $Y2=1.17
r249 13 14 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=3.975 $Y=1.245
+ $X2=3.975 $Y2=1.685
r250 12 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.58 $Y=1.76
+ $X2=3.415 $Y2=1.76
r251 11 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.9 $Y=1.76
+ $X2=3.975 $Y2=1.685
r252 11 12 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.9 $Y=1.76
+ $X2=3.58 $Y2=1.76
r253 9 69 198.242 $w=1.8e-07 $l=5.1e-07 $layer=POLY_cond $X=3.455 $Y=2.525
+ $X2=3.455 $Y2=2.015
r254 2 33 600 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=2.505
+ $Y=1.935 $X2=2.64 $Y2=2.1
r255 1 60 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=2.59
+ $Y=0.595 $X2=2.755 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_1%A_841_401# 1 2 9 13 16 17 22 23 25 26 27 28
+ 29 30 33
c110 26 0 5.58686e-20 $X=4.63 $Y=1.005
c111 17 0 1.85606e-19 $X=4.417 $Y=2.155
c112 13 0 3.41044e-19 $X=4.475 $Y=0.805
r113 33 35 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=6.355 $Y=1.88
+ $X2=6.355 $Y2=2.59
r114 31 33 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=6.355 $Y=1.57
+ $X2=6.355 $Y2=1.88
r115 29 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.23 $Y=1.485
+ $X2=6.355 $Y2=1.57
r116 29 30 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.23 $Y=1.485
+ $X2=5.915 $Y2=1.485
r117 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.83 $Y=1.4
+ $X2=5.915 $Y2=1.485
r118 27 38 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.83 $Y=1.09
+ $X2=5.83 $Y2=1.005
r119 27 28 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.83 $Y=1.09
+ $X2=5.83 $Y2=1.4
r120 25 38 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.745 $Y=1.005
+ $X2=5.83 $Y2=1.005
r121 25 26 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=5.745 $Y=1.005
+ $X2=4.63 $Y2=1.005
r122 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.465
+ $Y=1.65 $X2=4.465 $Y2=1.65
r123 20 26 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=4.49 $Y=1.09
+ $X2=4.63 $Y2=1.005
r124 20 22 23.0489 $w=2.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.49 $Y=1.09
+ $X2=4.49 $Y2=1.65
r125 19 23 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.465 $Y=1.485
+ $X2=4.465 $Y2=1.65
r126 16 23 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=4.465 $Y=2.005
+ $X2=4.465 $Y2=1.65
r127 16 17 38.0674 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=4.417 $Y=2.005
+ $X2=4.417 $Y2=2.155
r128 13 19 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.475 $Y=0.805
+ $X2=4.475 $Y2=1.485
r129 9 17 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=4.295 $Y=2.525
+ $X2=4.295 $Y2=2.155
r130 2 35 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=6.18
+ $Y=1.735 $X2=6.315 $Y2=2.59
r131 2 33 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.18
+ $Y=1.735 $X2=6.315 $Y2=1.88
r132 1 38 182 $w=1.7e-07 $l=7.36834e-07 $layer=licon1_NDIFF $count=1 $X=5.53
+ $Y=0.37 $X2=5.75 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_1%RESET_B 4 6 9 11 12 16 18 21 25 29 32 34 35
+ 36 37 38 43 46 49 50 53 54 57 61 62
c211 54 0 1.26008e-19 $X=1.165 $Y=1.295
c212 43 0 6.85463e-20 $X=7.92 $Y=2.035
c213 36 0 1.31208e-20 $X=1.345 $Y=2.035
c214 11 0 4.00428e-20 $X=4.79 $Y=0.18
r215 61 64 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.135 $Y=2
+ $X2=8.135 $Y2=2.165
r216 61 63 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.135 $Y=2
+ $X2=8.135 $Y2=1.835
r217 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.135
+ $Y=2 $X2=8.135 $Y2=2
r218 57 59 41.4566 $w=4.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.097 $Y=1.975
+ $X2=1.097 $Y2=2.14
r219 57 58 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.165
+ $Y=1.975 $X2=1.165 $Y2=1.975
r220 54 58 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.165 $Y=1.295
+ $X2=1.165 $Y2=1.975
r221 53 55 47.3569 $w=4.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.097 $Y=1.295
+ $X2=1.097 $Y2=1.13
r222 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.165
+ $Y=1.295 $X2=1.165 $Y2=1.295
r223 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.395
+ $Y=1.99 $X2=5.395 $Y2=1.99
r224 46 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.035
+ $X2=1.2 $Y2=2.035
r225 44 62 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=7.92 $Y=2
+ $X2=8.135 $Y2=2
r226 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r227 40 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=2.035
+ $X2=5.52 $Y2=2.035
r228 38 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=2.035
+ $X2=5.52 $Y2=2.035
r229 37 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r230 37 38 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=5.665 $Y2=2.035
r231 36 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=2.035
+ $X2=1.2 $Y2=2.035
r232 35 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=2.035
+ $X2=5.52 $Y2=2.035
r233 35 36 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=5.375 $Y=2.035
+ $X2=1.345 $Y2=2.035
r234 33 49 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=5.02 $Y=1.99
+ $X2=5.395 $Y2=1.99
r235 33 34 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.02 $Y=1.99 $X2=4.93
+ $Y2=1.99
r236 31 32 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=4.89 $Y=1.09 $X2=4.89
+ $Y2=1.24
r237 29 64 155.484 $w=1.8e-07 $l=4e-07 $layer=POLY_cond $X=8.18 $Y=2.565
+ $X2=8.18 $Y2=2.165
r238 25 63 643.521 $w=1.5e-07 $l=1.255e-06 $layer=POLY_cond $X=8.045 $Y=0.58
+ $X2=8.045 $Y2=1.835
r239 19 34 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=4.93 $Y=2.155
+ $X2=4.93 $Y2=1.99
r240 19 21 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=4.93 $Y=2.155
+ $X2=4.93 $Y2=2.525
r241 18 34 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=4.915 $Y=1.825
+ $X2=4.93 $Y2=1.99
r242 18 32 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=4.915 $Y=1.825
+ $X2=4.915 $Y2=1.24
r243 16 31 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.865 $Y=0.805
+ $X2=4.865 $Y2=1.09
r244 13 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.865 $Y=0.255
+ $X2=4.865 $Y2=0.805
r245 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.79 $Y=0.18
+ $X2=4.865 $Y2=0.255
r246 11 12 1935.69 $w=1.5e-07 $l=3.775e-06 $layer=POLY_cond $X=4.79 $Y=0.18
+ $X2=1.015 $Y2=0.18
r247 9 59 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=0.955 $Y=2.75
+ $X2=0.955 $Y2=2.14
r248 6 57 8.0134 $w=4.65e-07 $l=6.7e-08 $layer=POLY_cond $X=1.097 $Y=1.908
+ $X2=1.097 $Y2=1.975
r249 5 53 8.0134 $w=4.65e-07 $l=6.7e-08 $layer=POLY_cond $X=1.097 $Y=1.362
+ $X2=1.097 $Y2=1.295
r250 5 6 65.3032 $w=4.65e-07 $l=5.46e-07 $layer=POLY_cond $X=1.097 $Y=1.362
+ $X2=1.097 $Y2=1.908
r251 4 55 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.94 $Y=0.6 $X2=0.94
+ $Y2=1.13
r252 1 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.94 $Y=0.255
+ $X2=1.015 $Y2=0.18
r253 1 4 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=0.94 $Y=0.255
+ $X2=0.94 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_1%A_709_463# 1 2 3 12 14 16 18 24 25 28 32 35
+ 36 37 40 41
c127 37 0 1.55214e-19 $X=4.975 $Y=1.45
c128 35 0 7.39987e-20 $X=4.01 $Y=2.585
c129 32 0 1.09016e-19 $X=4.095 $Y=0.812
c130 24 0 2.17414e-19 $X=4.095 $Y=2.415
c131 14 0 2.11006e-19 $X=6 $Y=1.54
r132 41 43 7.32792 $w=3.08e-07 $l=1.85e-07 $layer=LI1_cond $X=4.975 $Y=2.515
+ $X2=5.16 $Y2=2.515
r133 40 46 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.395 $Y=1.45
+ $X2=5.395 $Y2=1.54
r134 40 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.395 $Y=1.45
+ $X2=5.395 $Y2=1.285
r135 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.395
+ $Y=1.45 $X2=5.395 $Y2=1.45
r136 37 39 20.6613 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=4.975 $Y=1.45
+ $X2=5.395 $Y2=1.45
r137 34 36 8.81087 $w=3.38e-07 $l=1.75e-07 $layer=LI1_cond $X=4.095 $Y=2.585
+ $X2=4.27 $Y2=2.585
r138 34 35 4.09336 $w=3.38e-07 $l=8.5e-08 $layer=LI1_cond $X=4.095 $Y=2.585
+ $X2=4.01 $Y2=2.585
r139 30 32 5.96091 $w=4.33e-07 $l=2.25e-07 $layer=LI1_cond $X=3.87 $Y=0.812
+ $X2=4.095 $Y2=0.812
r140 28 41 4.21588 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.975 $Y=2.35
+ $X2=4.975 $Y2=2.515
r141 27 37 2.94836 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.975 $Y=1.615
+ $X2=4.975 $Y2=1.45
r142 27 28 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=4.975 $Y=1.615
+ $X2=4.975 $Y2=2.35
r143 25 41 5.79756 $w=3.08e-07 $l=9.21954e-08 $layer=LI1_cond $X=4.89 $Y=2.5
+ $X2=4.975 $Y2=2.515
r144 25 36 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.89 $Y=2.5
+ $X2=4.27 $Y2=2.5
r145 24 34 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.095 $Y=2.415
+ $X2=4.095 $Y2=2.585
r146 23 32 6.29128 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=4.095 $Y=1.03
+ $X2=4.095 $Y2=0.812
r147 23 24 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=4.095 $Y=1.03
+ $X2=4.095 $Y2=2.415
r148 21 35 16.5351 $w=2.28e-07 $l=3.3e-07 $layer=LI1_cond $X=3.68 $Y=2.64
+ $X2=4.01 $Y2=2.64
r149 16 18 166.022 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=6.09 $Y=1.615
+ $X2=6.09 $Y2=2.235
r150 15 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.56 $Y=1.54
+ $X2=5.395 $Y2=1.54
r151 14 16 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6 $Y=1.54
+ $X2=6.09 $Y2=1.615
r152 14 15 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=6 $Y=1.54 $X2=5.56
+ $Y2=1.54
r153 12 45 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=5.455 $Y=0.69
+ $X2=5.455 $Y2=1.285
r154 3 43 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=5.02
+ $Y=2.315 $X2=5.16 $Y2=2.515
r155 2 21 600 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_PDIFF $count=1 $X=3.545
+ $Y=2.315 $X2=3.68 $Y2=2.61
r156 1 30 182 $w=1.7e-07 $l=3.02283e-07 $layer=licon1_NDIFF $count=1 $X=3.66
+ $Y=0.595 $X2=3.87 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_1%A_307_387# 1 2 9 11 13 15 17 18 19 20 21 24
+ 28 30 35 36 37 40 42 43 45 46 49 51 58
c189 51 0 1.65606e-19 $X=1.735 $Y=0.715
c190 49 0 3.57624e-20 $X=2.555 $Y=1.44
c191 42 0 1.19314e-19 $X=2.95 $Y=2.2
c192 24 0 1.58258e-20 $X=3.585 $Y=0.805
c193 20 0 4.1286e-20 $X=3.51 $Y=1.4
c194 17 0 7.39987e-20 $X=2.935 $Y=3.075
r195 62 66 51.2207 $w=3.67e-07 $l=3.9e-07 $layer=POLY_cond $X=2.56 $Y=1.55
+ $X2=2.95 $Y2=1.55
r196 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.56
+ $Y=1.61 $X2=2.56 $Y2=1.61
r197 53 54 7.09776 $w=4.48e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=1.055
+ $X2=1.695 $Y2=1.14
r198 51 53 9.03704 $w=4.48e-07 $l=3.4e-07 $layer=LI1_cond $X=1.695 $Y=0.715
+ $X2=1.695 $Y2=1.055
r199 49 61 9.5639 $w=2.2e-07 $l=1.7e-07 $layer=LI1_cond $X=2.555 $Y=1.44
+ $X2=2.555 $Y2=1.61
r200 48 49 15.7151 $w=2.18e-07 $l=3e-07 $layer=LI1_cond $X=2.555 $Y=1.14
+ $X2=2.555 $Y2=1.44
r201 47 53 6.50032 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=1.92 $Y=1.055
+ $X2=1.695 $Y2=1.055
r202 46 48 9.16439 $w=1.48e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.445 $Y=1.055
+ $X2=2.555 $Y2=1.14
r203 46 47 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.445 $Y=1.055
+ $X2=1.92 $Y2=1.055
r204 45 58 4.10192 $w=2.93e-07 $l=1.05e-07 $layer=LI1_cond $X=1.555 $Y=2.092
+ $X2=1.66 $Y2=2.092
r205 45 54 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.555 $Y=1.945
+ $X2=1.555 $Y2=1.14
r206 38 40 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=7.095 $Y=1.475
+ $X2=7.095 $Y2=0.58
r207 36 38 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.02 $Y=1.55
+ $X2=7.095 $Y2=1.475
r208 36 37 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=7.02 $Y=1.55
+ $X2=6.63 $Y2=1.55
r209 33 35 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=6.54 $Y=3.075
+ $X2=6.54 $Y2=2.235
r210 32 37 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.54 $Y=1.625
+ $X2=6.63 $Y2=1.55
r211 32 35 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=6.54 $Y=1.625
+ $X2=6.54 $Y2=2.235
r212 31 43 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.995 $Y=3.15
+ $X2=3.905 $Y2=3.15
r213 30 33 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.45 $Y=3.15
+ $X2=6.54 $Y2=3.075
r214 30 31 1258.84 $w=1.5e-07 $l=2.455e-06 $layer=POLY_cond $X=6.45 $Y=3.15
+ $X2=3.995 $Y2=3.15
r215 26 43 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.905 $Y=3.075
+ $X2=3.905 $Y2=3.15
r216 26 28 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=3.905 $Y=3.075
+ $X2=3.905 $Y2=2.525
r217 22 24 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=3.585 $Y=1.325
+ $X2=3.585 $Y2=0.805
r218 21 66 37.0402 $w=3.67e-07 $l=2.12132e-07 $layer=POLY_cond $X=3.1 $Y=1.4
+ $X2=2.95 $Y2=1.55
r219 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.51 $Y=1.4
+ $X2=3.585 $Y2=1.325
r220 20 21 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.51 $Y=1.4 $X2=3.1
+ $Y2=1.4
r221 18 43 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.815 $Y=3.15
+ $X2=3.905 $Y2=3.15
r222 18 19 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=3.815 $Y=3.15
+ $X2=3.01 $Y2=3.15
r223 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.935 $Y=3.075
+ $X2=3.01 $Y2=3.15
r224 17 42 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=2.935 $Y=3.075
+ $X2=2.935 $Y2=2.2
r225 15 42 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.95 $Y=2.11 $X2=2.95
+ $Y2=2.2
r226 14 66 19.4219 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=2.95 $Y=1.775
+ $X2=2.95 $Y2=1.55
r227 14 15 130.218 $w=1.8e-07 $l=3.35e-07 $layer=POLY_cond $X=2.95 $Y=1.775
+ $X2=2.95 $Y2=2.11
r228 11 62 5.91008 $w=3.67e-07 $l=4.5e-08 $layer=POLY_cond $X=2.515 $Y=1.55
+ $X2=2.56 $Y2=1.55
r229 11 63 13.1335 $w=3.67e-07 $l=1e-07 $layer=POLY_cond $X=2.515 $Y=1.55
+ $X2=2.415 $Y2=1.55
r230 11 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.515 $Y=1.41
+ $X2=2.515 $Y2=0.965
r231 7 63 19.4219 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=2.415 $Y=1.775
+ $X2=2.415 $Y2=1.55
r232 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.415 $Y=1.775
+ $X2=2.415 $Y2=2.495
r233 2 58 600 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=1 $X=1.535
+ $Y=1.935 $X2=1.66 $Y2=2.1
r234 1 51 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.59
+ $Y=0.59 $X2=1.735 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_1%A_1482_48# 1 2 7 9 12 14 17 20 23 24 37 39
+ 43
c93 37 0 6.85463e-20 $X=8.885 $Y=1.85
c94 14 0 1.98491e-19 $X=8.485 $Y=0.985
r95 35 37 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.555 $Y=1.85
+ $X2=8.885 $Y2=1.85
r96 28 43 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.595 $Y=1.065
+ $X2=7.67 $Y2=1.065
r97 28 40 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=7.595 $Y=1.065
+ $X2=7.485 $Y2=1.065
r98 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.595
+ $Y=1.065 $X2=7.595 $Y2=1.065
r99 24 27 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.595 $Y=0.985
+ $X2=7.595 $Y2=1.065
r100 23 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.885 $Y=1.765
+ $X2=8.885 $Y2=1.85
r101 22 39 2.90768 $w=3.27e-07 $l=1.95944e-07 $layer=LI1_cond $X=8.885 $Y=1.07
+ $X2=8.727 $Y2=0.985
r102 22 23 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=8.885 $Y=1.07
+ $X2=8.885 $Y2=1.765
r103 18 39 2.90768 $w=3.27e-07 $l=8.5e-08 $layer=LI1_cond $X=8.727 $Y=0.9
+ $X2=8.727 $Y2=0.985
r104 18 20 7.89165 $w=4.83e-07 $l=3.2e-07 $layer=LI1_cond $X=8.727 $Y=0.9
+ $X2=8.727 $Y2=0.58
r105 17 31 4.37637 $w=3.93e-07 $l=1.5e-07 $layer=LI1_cond $X=8.555 $Y=2.532
+ $X2=8.405 $Y2=2.532
r106 16 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.555 $Y=1.935
+ $X2=8.555 $Y2=1.85
r107 16 17 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=8.555 $Y=1.935
+ $X2=8.555 $Y2=2.335
r108 15 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.76 $Y=0.985
+ $X2=7.595 $Y2=0.985
r109 14 39 3.78066 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=8.485 $Y=0.985
+ $X2=8.727 $Y2=0.985
r110 14 15 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=8.485 $Y=0.985
+ $X2=7.76 $Y2=0.985
r111 10 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.67 $Y=1.23
+ $X2=7.67 $Y2=1.065
r112 10 12 518.927 $w=1.8e-07 $l=1.335e-06 $layer=POLY_cond $X=7.67 $Y=1.23
+ $X2=7.67 $Y2=2.565
r113 7 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.485 $Y=0.9
+ $X2=7.485 $Y2=1.065
r114 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.485 $Y=0.9
+ $X2=7.485 $Y2=0.58
r115 2 31 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=8.27
+ $Y=2.355 $X2=8.405 $Y2=2.565
r116 1 20 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.51
+ $Y=0.37 $X2=8.65 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_1%A_1224_74# 1 2 9 13 15 16 19 23 25 26 29 33
+ 37 38 42 47 48 49 51 52 54 56
c159 51 0 1.03385e-19 $X=7.58 $Y=2.365
c160 29 0 1.88583e-19 $X=10.5 $Y=2.54
c161 16 0 1.98491e-19 $X=8.72 $Y=1.43
r162 57 64 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=8.495 $Y=1.43
+ $X2=8.63 $Y2=1.43
r163 57 61 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=8.495 $Y=1.43
+ $X2=8.435 $Y2=1.43
r164 56 59 3.07318 $w=2.98e-07 $l=8e-08 $layer=LI1_cond $X=8.48 $Y=1.43 $X2=8.48
+ $Y2=1.51
r165 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.495
+ $Y=1.43 $X2=8.495 $Y2=1.43
r166 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.665 $Y=1.51
+ $X2=7.58 $Y2=1.51
r167 52 59 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=8.33 $Y=1.51 $X2=8.48
+ $Y2=1.51
r168 52 53 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=8.33 $Y=1.51
+ $X2=7.665 $Y2=1.51
r169 50 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.58 $Y=1.595
+ $X2=7.58 $Y2=1.51
r170 50 51 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=7.58 $Y=1.595
+ $X2=7.58 $Y2=2.365
r171 48 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.495 $Y=1.51
+ $X2=7.58 $Y2=1.51
r172 48 49 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.495 $Y=1.51
+ $X2=7.16 $Y2=1.51
r173 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.075 $Y=1.425
+ $X2=7.16 $Y2=1.51
r174 46 47 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=7.075 $Y=0.73
+ $X2=7.075 $Y2=1.425
r175 42 51 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.495 $Y=2.53
+ $X2=7.58 $Y2=2.365
r176 42 44 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=7.495 $Y=2.53
+ $X2=6.89 $Y2=2.53
r177 38 46 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.99 $Y=0.565
+ $X2=7.075 $Y2=0.73
r178 38 40 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.99 $Y=0.565
+ $X2=6.695 $Y2=0.565
r179 35 36 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=9.145 $Y=1.43
+ $X2=9.44 $Y2=1.43
r180 31 37 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=10.515
+ $Y=1.265 $X2=10.5 $Y2=1.43
r181 31 33 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=10.515 $Y=1.265
+ $X2=10.515 $Y2=0.645
r182 27 37 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=10.5 $Y=1.595
+ $X2=10.5 $Y2=1.43
r183 27 29 367.331 $w=1.8e-07 $l=9.45e-07 $layer=POLY_cond $X=10.5 $Y=1.595
+ $X2=10.5 $Y2=2.54
r184 26 36 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.515 $Y=1.43
+ $X2=9.44 $Y2=1.43
r185 25 37 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=10.41 $Y=1.43
+ $X2=10.5 $Y2=1.43
r186 25 26 156.501 $w=3.3e-07 $l=8.95e-07 $layer=POLY_cond $X=10.41 $Y=1.43
+ $X2=9.515 $Y2=1.43
r187 21 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.44 $Y=1.265
+ $X2=9.44 $Y2=1.43
r188 21 23 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=9.44 $Y=1.265
+ $X2=9.44 $Y2=0.74
r189 17 35 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.145 $Y=1.595
+ $X2=9.145 $Y2=1.43
r190 17 19 312.911 $w=1.8e-07 $l=8.05e-07 $layer=POLY_cond $X=9.145 $Y=1.595
+ $X2=9.145 $Y2=2.4
r191 16 64 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.72 $Y=1.43 $X2=8.63
+ $Y2=1.43
r192 15 35 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.055 $Y=1.43
+ $X2=9.145 $Y2=1.43
r193 15 16 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=9.055 $Y=1.43
+ $X2=8.72 $Y2=1.43
r194 11 64 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.63 $Y=1.595
+ $X2=8.63 $Y2=1.43
r195 11 13 377.048 $w=1.8e-07 $l=9.7e-07 $layer=POLY_cond $X=8.63 $Y=1.595
+ $X2=8.63 $Y2=2.565
r196 7 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.435 $Y=1.265
+ $X2=8.435 $Y2=1.43
r197 7 9 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=8.435 $Y=1.265
+ $X2=8.435 $Y2=0.58
r198 2 44 600 $w=1.7e-07 $l=9.15819e-07 $layer=licon1_PDIFF $count=1 $X=6.63
+ $Y=1.735 $X2=6.89 $Y2=2.53
r199 1 40 182 $w=1.7e-07 $l=6.65395e-07 $layer=licon1_NDIFF $count=1 $X=6.12
+ $Y=0.37 $X2=6.695 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_1%A_2026_424# 1 2 9 13 17 21 25 26 28
r52 26 31 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.965 $Y=1.465
+ $X2=10.965 $Y2=1.63
r53 26 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.965 $Y=1.465
+ $X2=10.965 $Y2=1.3
r54 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.965
+ $Y=1.465 $X2=10.965 $Y2=1.465
r55 23 28 0.364692 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=10.44 $Y=1.465
+ $X2=10.315 $Y2=1.465
r56 23 25 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=10.44 $Y=1.465
+ $X2=10.965 $Y2=1.465
r57 19 28 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=10.315 $Y=1.63
+ $X2=10.315 $Y2=1.465
r58 19 21 29.5025 $w=2.48e-07 $l=6.4e-07 $layer=LI1_cond $X=10.315 $Y=1.63
+ $X2=10.315 $Y2=2.27
r59 15 28 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=10.315 $Y=1.3
+ $X2=10.315 $Y2=1.465
r60 15 17 30.4245 $w=2.48e-07 $l=6.6e-07 $layer=LI1_cond $X=10.315 $Y=1.3
+ $X2=10.315 $Y2=0.64
r61 13 30 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.015 $Y=0.74
+ $X2=11.015 $Y2=1.3
r62 9 31 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=11.015 $Y=2.4
+ $X2=11.015 $Y2=1.63
r63 2 21 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=10.13
+ $Y=2.12 $X2=10.275 $Y2=2.27
r64 1 17 182 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_NDIFF $count=1 $X=10.155
+ $Y=0.37 $X2=10.3 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_1%VPWR 1 2 3 4 5 6 7 8 25 27 31 35 39 43 49 51
+ 55 59 63 65 70 75 83 88 93 103 104 110 113 116 119 122 125 128
r146 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r147 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r148 123 126 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r149 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r150 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r151 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r152 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r153 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r154 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r155 104 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r156 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r157 101 128 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=10.905 $Y=3.33
+ $X2=10.757 $Y2=3.33
r158 101 103 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=10.905 $Y=3.33
+ $X2=11.28 $Y2=3.33
r159 100 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r160 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r161 97 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r162 97 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r163 96 99 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r164 96 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r165 94 125 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=9.025 $Y=3.33
+ $X2=8.917 $Y2=3.33
r166 94 96 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.025 $Y=3.33
+ $X2=9.36 $Y2=3.33
r167 93 128 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=10.61 $Y=3.33
+ $X2=10.757 $Y2=3.33
r168 93 99 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=10.61 $Y=3.33
+ $X2=10.32 $Y2=3.33
r169 92 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r170 92 120 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6 $Y2=3.33
r171 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r172 89 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.03 $Y=3.33
+ $X2=5.905 $Y2=3.33
r173 89 91 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=6.03 $Y=3.33
+ $X2=7.44 $Y2=3.33
r174 88 122 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=7.835 $Y=3.33
+ $X2=7.947 $Y2=3.33
r175 88 91 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=7.835 $Y=3.33
+ $X2=7.44 $Y2=3.33
r176 87 117 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r177 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r178 84 116 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=4.785 $Y=3.33
+ $X2=4.612 $Y2=3.33
r179 84 86 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=4.785 $Y=3.33
+ $X2=5.52 $Y2=3.33
r180 83 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.78 $Y=3.33
+ $X2=5.905 $Y2=3.33
r181 83 86 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.78 $Y=3.33
+ $X2=5.52 $Y2=3.33
r182 82 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r183 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r184 79 82 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r185 79 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r186 78 81 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r187 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r188 76 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=3.33
+ $X2=2.19 $Y2=3.33
r189 76 78 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.355 $Y=3.33
+ $X2=2.64 $Y2=3.33
r190 75 116 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=4.44 $Y=3.33
+ $X2=4.612 $Y2=3.33
r191 75 81 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.44 $Y=3.33
+ $X2=4.08 $Y2=3.33
r192 74 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r193 74 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r194 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r195 71 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.18 $Y2=3.33
r196 71 73 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r197 70 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=2.19 $Y2=3.33
r198 70 73 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=1.68 $Y2=3.33
r199 69 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r200 69 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r201 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r202 66 107 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r203 66 68 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r204 65 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.18 $Y2=3.33
r205 65 68 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r206 63 120 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=6 $Y2=3.33
r207 63 87 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=5.52 $Y2=3.33
r208 59 62 16.2123 $w=2.93e-07 $l=4.15e-07 $layer=LI1_cond $X=10.757 $Y=1.985
+ $X2=10.757 $Y2=2.4
r209 57 128 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=10.757 $Y=3.245
+ $X2=10.757 $Y2=3.33
r210 57 62 33.0107 $w=2.93e-07 $l=8.45e-07 $layer=LI1_cond $X=10.757 $Y=3.245
+ $X2=10.757 $Y2=2.4
r211 53 125 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=8.917 $Y=3.245
+ $X2=8.917 $Y2=3.33
r212 53 55 52.262 $w=2.13e-07 $l=9.75e-07 $layer=LI1_cond $X=8.917 $Y=3.245
+ $X2=8.917 $Y2=2.27
r213 52 122 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=8.06 $Y=3.33
+ $X2=7.947 $Y2=3.33
r214 51 125 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=8.81 $Y=3.33
+ $X2=8.917 $Y2=3.33
r215 51 52 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=8.81 $Y=3.33
+ $X2=8.06 $Y2=3.33
r216 47 122 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=7.947 $Y=3.245
+ $X2=7.947 $Y2=3.33
r217 47 49 34.8294 $w=2.23e-07 $l=6.8e-07 $layer=LI1_cond $X=7.947 $Y=3.245
+ $X2=7.947 $Y2=2.565
r218 43 46 31.5769 $w=2.48e-07 $l=6.85e-07 $layer=LI1_cond $X=5.905 $Y=1.905
+ $X2=5.905 $Y2=2.59
r219 41 119 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.905 $Y=3.245
+ $X2=5.905 $Y2=3.33
r220 41 46 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=5.905 $Y=3.245
+ $X2=5.905 $Y2=2.59
r221 37 116 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=4.612 $Y=3.245
+ $X2=4.612 $Y2=3.33
r222 37 39 13.5287 $w=3.43e-07 $l=4.05e-07 $layer=LI1_cond $X=4.612 $Y=3.245
+ $X2=4.612 $Y2=2.84
r223 33 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=3.33
r224 33 35 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=2.835
r225 29 110 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r226 29 31 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.835
r227 25 107 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r228 25 27 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.75
r229 8 62 300 $w=1.7e-07 $l=3.54965e-07 $layer=licon1_PDIFF $count=2 $X=10.59
+ $Y=2.12 $X2=10.76 $Y2=2.4
r230 8 59 600 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_PDIFF $count=1 $X=10.59
+ $Y=2.12 $X2=10.79 $Y2=1.985
r231 7 55 300 $w=1.7e-07 $l=2.38747e-07 $layer=licon1_PDIFF $count=2 $X=8.72
+ $Y=2.355 $X2=8.92 $Y2=2.27
r232 6 49 600 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=2.355 $X2=7.92 $Y2=2.565
r233 5 46 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.72
+ $Y=1.735 $X2=5.865 $Y2=2.59
r234 5 43 400 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=5.72
+ $Y=1.735 $X2=5.865 $Y2=1.905
r235 4 39 600 $w=1.7e-07 $l=6.27495e-07 $layer=licon1_PDIFF $count=1 $X=4.385
+ $Y=2.315 $X2=4.61 $Y2=2.84
r236 3 35 600 $w=1.7e-07 $l=9.65142e-07 $layer=licon1_PDIFF $count=1 $X=2.055
+ $Y=1.935 $X2=2.19 $Y2=2.835
r237 2 31 600 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=2.54 $X2=1.18 $Y2=2.835
r238 1 27 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.28 $Y2=2.75
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_1%A_38_78# 1 2 3 4 13 17 20 21 25 27 30 32 36
+ 38 43
c117 38 0 1.19314e-19 $X=3.205 $Y=2.495
r118 38 40 1.47581 $w=2.48e-07 $l=3e-08 $layer=LI1_cond $X=3.205 $Y=2.495
+ $X2=3.205 $Y2=2.525
r119 37 38 11.0685 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=3.205 $Y=2.27
+ $X2=3.205 $Y2=2.495
r120 32 34 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.335 $Y=0.6
+ $X2=0.335 $Y2=0.745
r121 29 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.755 $Y=1.37
+ $X2=3.755 $Y2=1.285
r122 29 30 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=3.755 $Y=1.37
+ $X2=3.755 $Y2=2.185
r123 28 37 2.94836 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.345 $Y=2.27
+ $X2=3.205 $Y2=2.27
r124 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.67 $Y=2.27
+ $X2=3.755 $Y2=2.185
r125 27 28 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.67 $Y=2.27
+ $X2=3.345 $Y2=2.27
r126 23 43 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.41 $Y=1.285
+ $X2=3.755 $Y2=1.285
r127 23 25 17.9781 $w=2.48e-07 $l=3.9e-07 $layer=LI1_cond $X=3.41 $Y=1.2
+ $X2=3.41 $Y2=0.81
r128 22 36 2.36881 $w=1.7e-07 $l=3.37268e-07 $layer=LI1_cond $X=0.89 $Y=2.495
+ $X2=0.565 $Y2=2.52
r129 21 38 2.94836 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.065 $Y=2.495
+ $X2=3.205 $Y2=2.495
r130 21 22 141.898 $w=1.68e-07 $l=2.175e-06 $layer=LI1_cond $X=3.065 $Y=2.495
+ $X2=0.89 $Y2=2.495
r131 20 36 4.06715 $w=2.25e-07 $l=2.5923e-07 $layer=LI1_cond $X=0.775 $Y=2.41
+ $X2=0.565 $Y2=2.52
r132 19 20 103.08 $w=1.68e-07 $l=1.58e-06 $layer=LI1_cond $X=0.775 $Y=0.83
+ $X2=0.775 $Y2=2.41
r133 15 36 4.06715 $w=2.25e-07 $l=1.85203e-07 $layer=LI1_cond $X=0.705 $Y=2.625
+ $X2=0.565 $Y2=2.52
r134 15 17 5.14483 $w=2.78e-07 $l=1.25e-07 $layer=LI1_cond $X=0.705 $Y=2.625
+ $X2=0.705 $Y2=2.75
r135 14 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.5 $Y=0.745
+ $X2=0.335 $Y2=0.745
r136 13 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.69 $Y=0.745
+ $X2=0.775 $Y2=0.83
r137 13 14 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.69 $Y=0.745
+ $X2=0.5 $Y2=0.745
r138 4 40 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=3.085
+ $Y=2.315 $X2=3.23 $Y2=2.525
r139 3 17 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=2.54 $X2=0.73 $Y2=2.75
r140 2 25 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=3.225
+ $Y=0.595 $X2=3.37 $Y2=0.81
r141 1 32 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.19
+ $Y=0.39 $X2=0.335 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_1%Q_N 1 2 9 11 12 13 26
c24 12 0 1.88583e-19 $X=9.84 $Y=2.405
r25 26 27 5.27602 $w=6.88e-07 $l=1.75e-07 $layer=LI1_cond $X=9.605 $Y=1.985
+ $X2=9.605 $Y2=1.81
r26 13 23 0.693379 $w=6.88e-07 $l=4e-08 $layer=LI1_cond $X=9.605 $Y=2.775
+ $X2=9.605 $Y2=2.815
r27 12 13 6.41375 $w=6.88e-07 $l=3.7e-07 $layer=LI1_cond $X=9.605 $Y=2.405
+ $X2=9.605 $Y2=2.775
r28 12 17 4.33362 $w=6.88e-07 $l=2.5e-07 $layer=LI1_cond $X=9.605 $Y=2.405
+ $X2=9.605 $Y2=2.155
r29 11 17 2.08014 $w=6.88e-07 $l=1.2e-07 $layer=LI1_cond $X=9.605 $Y=2.035
+ $X2=9.605 $Y2=2.155
r30 11 26 0.866723 $w=6.88e-07 $l=5e-08 $layer=LI1_cond $X=9.605 $Y=2.035
+ $X2=9.605 $Y2=1.985
r31 9 27 38.267 $w=3.88e-07 $l=1.295e-06 $layer=LI1_cond $X=9.755 $Y=0.515
+ $X2=9.755 $Y2=1.81
r32 2 26 200 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=3 $X=9.235
+ $Y=1.84 $X2=9.37 $Y2=1.985
r33 2 23 200 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=3 $X=9.235
+ $Y=1.84 $X2=9.37 $Y2=2.815
r34 1 9 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=9.515
+ $Y=0.37 $X2=9.725 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_1%Q 1 2 9 10 11 24 27 35
r24 33 35 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=11.35 $Y=1.13
+ $X2=11.35 $Y2=1.82
r25 25 27 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=11.255 $Y=2
+ $X2=11.255 $Y2=2.035
r26 17 24 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=11.25 $Y=0.945
+ $X2=11.25 $Y2=0.925
r27 11 25 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=11.255 $Y=1.975
+ $X2=11.255 $Y2=2
r28 11 35 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=11.255 $Y=1.975
+ $X2=11.255 $Y2=1.82
r29 11 30 24.1693 $w=3.58e-07 $l=7.55e-07 $layer=LI1_cond $X=11.255 $Y=2.06
+ $X2=11.255 $Y2=2.815
r30 11 27 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=11.255 $Y=2.06
+ $X2=11.255 $Y2=2.035
r31 10 33 8.16504 $w=3.68e-07 $l=1.53e-07 $layer=LI1_cond $X=11.25 $Y=0.977
+ $X2=11.25 $Y2=1.13
r32 10 17 0.996707 $w=3.68e-07 $l=3.2e-08 $layer=LI1_cond $X=11.25 $Y=0.977
+ $X2=11.25 $Y2=0.945
r33 10 24 1.02785 $w=3.68e-07 $l=3.3e-08 $layer=LI1_cond $X=11.25 $Y=0.892
+ $X2=11.25 $Y2=0.925
r34 9 10 11.7425 $w=3.68e-07 $l=3.77e-07 $layer=LI1_cond $X=11.25 $Y=0.515
+ $X2=11.25 $Y2=0.892
r35 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=11.105
+ $Y=1.84 $X2=11.24 $Y2=1.985
r36 2 30 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=11.105
+ $Y=1.84 $X2=11.24 $Y2=2.815
r37 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.09
+ $Y=0.37 $X2=11.23 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFRBP_1%VGND 1 2 3 4 5 6 21 23 27 31 35 39 43 45 50
+ 55 63 68 75 76 79 82 86 92 95 98
c115 76 0 1.90308e-19 $X=11.28 $Y=0
r116 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r117 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r118 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r119 86 89 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=5.16 $Y=0 $X2=5.16
+ $Y2=0.325
r120 86 87 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r121 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r122 80 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r123 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r124 76 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r125 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r126 73 98 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.895 $Y=0
+ $X2=10.77 $Y2=0
r127 73 75 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.895 $Y=0
+ $X2=11.28 $Y2=0
r128 72 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r129 72 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.36 $Y2=0
r130 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r131 69 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.39 $Y=0 $X2=9.265
+ $Y2=0
r132 69 71 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=9.39 $Y=0 $X2=10.32
+ $Y2=0
r133 68 98 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.645 $Y=0
+ $X2=10.77 $Y2=0
r134 68 71 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=10.645 $Y=0
+ $X2=10.32 $Y2=0
r135 67 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r136 67 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=7.92
+ $Y2=0
r137 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r138 64 92 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=7.995 $Y=0 $X2=7.765
+ $Y2=0
r139 64 66 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=7.995 $Y=0 $X2=8.88
+ $Y2=0
r140 63 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.14 $Y=0 $X2=9.265
+ $Y2=0
r141 63 66 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=9.14 $Y=0 $X2=8.88
+ $Y2=0
r142 62 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r143 61 62 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r144 59 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r145 58 61 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=7.44
+ $Y2=0
r146 58 59 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r147 56 86 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.325 $Y=0 $X2=5.16
+ $Y2=0
r148 56 58 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.325 $Y=0
+ $X2=5.52 $Y2=0
r149 55 92 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=7.535 $Y=0 $X2=7.765
+ $Y2=0
r150 55 61 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=7.535 $Y=0 $X2=7.44
+ $Y2=0
r151 54 87 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=5.04
+ $Y2=0
r152 54 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r153 53 54 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r154 51 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.42 $Y=0 $X2=2.255
+ $Y2=0
r155 51 53 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.42 $Y=0 $X2=2.64
+ $Y2=0
r156 50 86 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.995 $Y=0 $X2=5.16
+ $Y2=0
r157 50 53 153.642 $w=1.68e-07 $l=2.355e-06 $layer=LI1_cond $X=4.995 $Y=0
+ $X2=2.64 $Y2=0
r158 48 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r159 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r160 45 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=1.155
+ $Y2=0
r161 45 47 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=0.72
+ $Y2=0
r162 43 62 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=7.44 $Y2=0
r163 43 59 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=5.52 $Y2=0
r164 39 41 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=10.77 $Y=0.515
+ $X2=10.77 $Y2=0.965
r165 37 98 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.77 $Y=0.085
+ $X2=10.77 $Y2=0
r166 37 39 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.77 $Y=0.085
+ $X2=10.77 $Y2=0.515
r167 33 95 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.265 $Y=0.085
+ $X2=9.265 $Y2=0
r168 33 35 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.265 $Y=0.085
+ $X2=9.265 $Y2=0.515
r169 29 92 1.85547 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.765 $Y=0.085
+ $X2=7.765 $Y2=0
r170 29 31 12.2208 $w=4.58e-07 $l=4.7e-07 $layer=LI1_cond $X=7.765 $Y=0.085
+ $X2=7.765 $Y2=0.555
r171 25 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.255 $Y=0.085
+ $X2=2.255 $Y2=0
r172 25 27 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=2.255 $Y=0.085
+ $X2=2.255 $Y2=0.715
r173 24 79 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.155
+ $Y2=0
r174 23 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.09 $Y=0 $X2=2.255
+ $Y2=0
r175 23 24 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.09 $Y=0 $X2=1.28
+ $Y2=0
r176 19 79 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0
r177 19 21 23.7403 $w=2.48e-07 $l=5.15e-07 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0.6
r178 6 41 182 $w=1.7e-07 $l=6.87768e-07 $layer=licon1_NDIFF $count=1 $X=10.59
+ $Y=0.37 $X2=10.79 $Y2=0.965
r179 6 39 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=10.59
+ $Y=0.37 $X2=10.79 $Y2=0.515
r180 5 35 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=9.08
+ $Y=0.37 $X2=9.225 $Y2=0.515
r181 4 31 182 $w=1.7e-07 $l=2.82754e-07 $layer=licon1_NDIFF $count=1 $X=7.56
+ $Y=0.37 $X2=7.765 $Y2=0.555
r182 3 89 182 $w=1.7e-07 $l=3.63731e-07 $layer=licon1_NDIFF $count=1 $X=4.94
+ $Y=0.595 $X2=5.16 $Y2=0.325
r183 2 27 182 $w=1.7e-07 $l=2.37539e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.595 $X2=2.255 $Y2=0.715
r184 1 21 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.39 $X2=1.195 $Y2=0.6
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__o21ba_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__o21ba_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.175000 1.450000 4.675000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.552000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.845000 1.450000 6.115000 1.780000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.180000 0.835000 1.550000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  1.026600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.550000 1.315000 1.820000 ;
        RECT 1.085000 1.820000 2.345000 2.220000 ;
        RECT 1.145000 0.350000 1.340000 0.950000 ;
        RECT 1.145000 0.950000 2.210000 1.120000 ;
        RECT 1.145000 1.120000 1.315000 1.550000 ;
        RECT 1.960000 0.350000 2.210000 0.950000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.240000 0.085000 ;
        RECT 0.645000  0.085000 0.975000 1.010000 ;
        RECT 1.530000  0.085000 1.780000 0.780000 ;
        RECT 2.390000  0.085000 2.640000 1.120000 ;
        RECT 4.500000  0.085000 4.750000 0.940000 ;
        RECT 5.360000  0.085000 5.610000 0.940000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 6.240000 3.415000 ;
        RECT 0.615000 2.730000 0.995000 3.245000 ;
        RECT 1.565000 2.730000 1.895000 3.245000 ;
        RECT 2.465000 2.730000 3.205000 3.245000 ;
        RECT 3.945000 2.470000 4.275000 3.245000 ;
        RECT 5.875000 1.950000 6.125000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.350000 0.475000 1.010000 ;
      RECT 0.085000 1.010000 0.255000 1.820000 ;
      RECT 0.085000 1.820000 0.445000 2.390000 ;
      RECT 0.085000 2.390000 3.320000 2.560000 ;
      RECT 0.085000 2.560000 0.445000 2.980000 ;
      RECT 1.485000 1.290000 3.830000 1.460000 ;
      RECT 1.485000 1.460000 2.980000 1.620000 ;
      RECT 2.810000 0.255000 3.830000 0.425000 ;
      RECT 2.810000 0.425000 2.980000 1.290000 ;
      RECT 3.150000 0.595000 3.320000 0.950000 ;
      RECT 3.150000 0.950000 4.330000 1.110000 ;
      RECT 3.150000 1.110000 6.125000 1.120000 ;
      RECT 3.150000 1.630000 3.490000 1.960000 ;
      RECT 3.150000 1.960000 3.320000 2.390000 ;
      RECT 3.490000 2.130000 5.145000 2.300000 ;
      RECT 3.490000 2.300000 3.740000 2.980000 ;
      RECT 3.500000 0.425000 3.830000 0.780000 ;
      RECT 3.660000 1.460000 3.830000 1.950000 ;
      RECT 3.660000 1.950000 5.145000 2.130000 ;
      RECT 4.000000 0.605000 4.330000 0.950000 ;
      RECT 4.000000 1.120000 6.125000 1.280000 ;
      RECT 4.445000 2.470000 4.775000 2.905000 ;
      RECT 4.445000 2.905000 5.675000 3.075000 ;
      RECT 4.930000 0.605000 5.180000 1.110000 ;
      RECT 4.975000 2.300000 5.145000 2.735000 ;
      RECT 5.345000 1.950000 5.675000 2.905000 ;
      RECT 5.790000 0.605000 6.125000 1.110000 ;
  END
END sky130_fd_sc_ms__o21ba_4

* File: sky130_fd_sc_ms__a41o_1.spice
* Created: Fri Aug 28 17:09:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a41o_1.pex.spice"
.subckt sky130_fd_sc_ms__a41o_1  VNB VPB B1 A1 A2 A3 A4 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_83_244#_M1005_g N_X_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.7104 PD=1.16 PS=3.4 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.9
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1008 N_A_83_244#_M1008_d N_B1_M1008_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.5
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1003 A_449_74# N_A1_M1003_g N_A_83_244#_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1184 AS=0.1036 PD=1.06 PS=1.02 NRD=17.016 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1000 A_543_74# N_A2_M1000_g A_449_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.1184 PD=1.16 PS=1.06 NRD=25.128 NRS=17.016 M=1 R=4.93333 SA=75002.4
+ SB=75001.4 A=0.111 P=1.78 MULT=1
MM1006 A_657_74# N_A3_M1006_g A_543_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.1554 PD=1.16 PS=1.16 NRD=25.128 NRS=25.128 M=1 R=4.93333 SA=75002.9
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A4_M1009_g A_657_74# VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=25.128 M=1 R=4.93333 SA=75003.5 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1001 N_VPWR_M1001_d N_A_83_244#_M1001_g N_X_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.3136 PD=2.8 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1010 N_A_357_392#_M1010_d N_B1_M1010_g N_A_83_244#_M1010_s VPB PSHORT L=0.18
+ W=1 AD=0.16 AS=0.28 PD=1.32 PS=2.56 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90002.3 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1011_d N_A1_M1011_g N_A_357_392#_M1010_d VPB PSHORT L=0.18 W=1
+ AD=0.2 AS=0.16 PD=1.4 PS=1.32 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90000.7
+ SB=90001.8 A=0.18 P=2.36 MULT=1
MM1002 N_A_357_392#_M1002_d N_A2_M1002_g N_VPWR_M1011_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.2 PD=1.27 PS=1.4 NRD=0 NRS=14.7553 M=1 R=5.55556 SA=90001.3
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_A3_M1004_g N_A_357_392#_M1002_d VPB PSHORT L=0.18 W=1
+ AD=0.195 AS=0.135 PD=1.39 PS=1.27 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90001.7
+ SB=90000.8 A=0.18 P=2.36 MULT=1
MM1007 N_A_357_392#_M1007_d N_A4_M1007_g N_VPWR_M1004_d VPB PSHORT L=0.18 W=1
+ AD=0.28 AS=0.195 PD=2.56 PS=1.39 NRD=0 NRS=12.7853 M=1 R=5.55556 SA=90002.3
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__a41o_1.pxi.spice"
*
.ends
*
*

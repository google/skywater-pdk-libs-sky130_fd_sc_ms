* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor2b_2 A B_N VGND VNB VPB VPWR Y
M1000 a_228_368# a_27_392# Y VPB pshort w=1.12e+06u l=180000u
+  ad=9.24e+11p pd=8.37e+06u as=3.024e+11p ps=2.78e+06u
M1001 VPWR A a_228_368# VPB pshort w=1.12e+06u l=180000u
+  ad=5.824e+11p pd=5.34e+06u as=0p ps=0u
M1002 a_228_368# A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y a_27_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.884e+11p pd=4.28e+06u as=7.744e+11p ps=6.56e+06u
M1004 VPWR B_N a_27_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.75e+11p ps=2.55e+06u
M1005 VGND B_N a_27_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1006 VGND a_27_392# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_27_392# a_228_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

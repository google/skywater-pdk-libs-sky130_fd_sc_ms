* File: sky130_fd_sc_ms__dlrbn_1.spice
* Created: Wed Sep  2 12:04:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dlrbn_1.pex.spice"
.subckt sky130_fd_sc_ms__dlrbn_1  VNB VPB D GATE_N RESET_B VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_D_M1008_g N_A_27_424#_M1008_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.129591 AS=0.15675 PD=0.997674 PS=1.67 NRD=18 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1003 N_A_231_74#_M1003_d N_GATE_N_M1003_g N_VGND_M1008_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1015_d N_A_231_74#_M1015_g N_A_373_74#_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.215887 AS=0.2109 PD=1.42638 PS=2.05 NRD=30.804 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002 A=0.111 P=1.78 MULT=1
MM1001 A_608_74# N_A_27_424#_M1001_g N_VGND_M1015_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.186713 PD=0.88 PS=1.23362 NRD=12.18 NRS=22.488 M=1 R=4.26667
+ SA=75000.9 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1002 N_A_686_74#_M1002_d N_A_231_74#_M1002_g A_608_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.231547 AS=0.0768 PD=1.52755 PS=0.88 NRD=28.116 NRS=12.18 M=1
+ R=4.26667 SA=75001.3 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1014 A_841_118# N_A_373_74#_M1014_g N_A_686_74#_M1002_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.151953 PD=0.66 PS=1.00245 NRD=18.564 NRS=57.132 M=1
+ R=2.8 SA=75002.1 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_A_889_92#_M1023_g A_841_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1533 AS=0.0504 PD=1.57 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8 SA=75002.5
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1017 A_1133_74# N_A_686_74#_M1017_g N_A_889_92#_M1017_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_RESET_B_M1005_g A_1133_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1443 AS=0.0888 PD=1.13 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75000.6
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1018 N_Q_M1018_d N_A_889_92#_M1018_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1443 PD=2.05 PS=1.13 NRD=0 NRS=17.832 M=1 R=4.93333 SA=75001.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A_889_92#_M1010_g N_A_1437_112#_M1010_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.109083 AS=0.1925 PD=0.942248 PS=1.8 NRD=19.08 NRS=0 M=1
+ R=3.66667 SA=75000.3 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1020 N_Q_N_M1020_d N_A_1437_112#_M1020_g N_VGND_M1010_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.146767 PD=2.05 PS=1.26775 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1012 N_VPWR_M1012_d N_D_M1012_g N_A_27_424#_M1012_s VPB PSHORT L=0.18 W=0.84
+ AD=0.2436 AS=0.2352 PD=1.42 PS=2.24 NRD=0 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.9 A=0.1512 P=2.04 MULT=1
MM1007 N_A_231_74#_M1007_d N_GATE_N_M1007_g N_VPWR_M1012_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.2436 PD=2.24 PS=1.42 NRD=0 NRS=71.511 M=1 R=4.66667
+ SA=90000.9 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1022 N_VPWR_M1022_d N_A_231_74#_M1022_g N_A_373_74#_M1022_s VPB PSHORT L=0.18
+ W=0.84 AD=0.217898 AS=0.3704 PD=1.47 PS=2.85 NRD=47.9301 NRS=19.9167 M=1
+ R=4.66667 SA=90000.3 SB=90002.2 A=0.1512 P=2.04 MULT=1
MM1019 A_614_392# N_A_27_424#_M1019_g N_VPWR_M1022_d VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.259402 PD=1.24 PS=1.75 NRD=12.7853 NRS=16.7253 M=1 R=5.55556
+ SA=90000.8 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1006 N_A_686_74#_M1006_d N_A_373_74#_M1006_g A_614_392# VPB PSHORT L=0.18 W=1
+ AD=0.219366 AS=0.12 PD=1.90845 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556
+ SA=90001.2 SB=90001.3 A=0.18 P=2.36 MULT=1
MM1004 A_805_508# N_A_231_74#_M1004_g N_A_686_74#_M1006_d VPB PSHORT L=0.18
+ W=0.42 AD=0.10605 AS=0.0921338 PD=0.925 PS=0.801549 NRD=92.6294 NRS=39.8531
+ M=1 R=2.33333 SA=90001.6 SB=90002.2 A=0.0756 P=1.2 MULT=1
MM1011 N_VPWR_M1011_d N_A_889_92#_M1011_g A_805_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.124377 AS=0.10605 PD=1.08818 PS=0.925 NRD=0 NRS=92.6294 M=1 R=2.33333
+ SA=90002.3 SB=90001.5 A=0.0756 P=1.2 MULT=1
MM1013 N_A_889_92#_M1013_d N_A_686_74#_M1013_g N_VPWR_M1011_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1568 AS=0.331673 PD=1.4 PS=2.90182 NRD=0.8668 NRS=6.1464 M=1
+ R=6.22222 SA=90001 SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1000 N_VPWR_M1000_d N_RESET_B_M1000_g N_A_889_92#_M1013_d VPB PSHORT L=0.18
+ W=1.12 AD=0.196 AS=0.1568 PD=1.47 PS=1.4 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90001.5 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1016 N_Q_M1016_d N_A_889_92#_M1016_g N_VPWR_M1000_d VPB PSHORT L=0.18 W=1.12
+ AD=0.308 AS=0.196 PD=2.79 PS=1.47 NRD=1.7533 NRS=4.3931 M=1 R=6.22222 SA=90002
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1021 N_VPWR_M1021_d N_A_889_92#_M1021_g N_A_1437_112#_M1021_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1608 AS=0.2184 PD=1.26857 PS=2.2 NRD=37.5088 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1009 N_Q_N_M1009_d N_A_1437_112#_M1009_g N_VPWR_M1021_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.2144 PD=2.8 PS=1.69143 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX24_noxref VNB VPB NWDIODE A=17.3933 P=22.02
c_80 VNB 0 5.58535e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__dlrbn_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__or2_2.pxi.spice
* Created: Wed Sep  2 12:27:37 2020
* 
x_PM_SKY130_FD_SC_MS__OR2_2%B N_B_M1004_g N_B_c_52_n N_B_M1003_g B N_B_c_54_n
+ PM_SKY130_FD_SC_MS__OR2_2%B
x_PM_SKY130_FD_SC_MS__OR2_2%A N_A_M1000_g N_A_M1005_g A A N_A_c_78_n N_A_c_79_n
+ PM_SKY130_FD_SC_MS__OR2_2%A
x_PM_SKY130_FD_SC_MS__OR2_2%A_27_368# N_A_27_368#_M1003_d N_A_27_368#_M1004_s
+ N_A_27_368#_M1002_g N_A_27_368#_M1001_g N_A_27_368#_M1006_g
+ N_A_27_368#_M1007_g N_A_27_368#_c_135_n N_A_27_368#_c_136_n
+ N_A_27_368#_c_145_n N_A_27_368#_c_126_n N_A_27_368#_c_127_n
+ N_A_27_368#_c_128_n N_A_27_368#_c_129_n N_A_27_368#_c_138_n
+ N_A_27_368#_c_130_n N_A_27_368#_c_140_n N_A_27_368#_c_174_p
+ N_A_27_368#_c_131_n N_A_27_368#_c_132_n PM_SKY130_FD_SC_MS__OR2_2%A_27_368#
x_PM_SKY130_FD_SC_MS__OR2_2%VPWR N_VPWR_M1000_d N_VPWR_M1007_s N_VPWR_c_225_n
+ N_VPWR_c_226_n N_VPWR_c_227_n VPWR N_VPWR_c_228_n N_VPWR_c_229_n
+ N_VPWR_c_230_n N_VPWR_c_224_n PM_SKY130_FD_SC_MS__OR2_2%VPWR
x_PM_SKY130_FD_SC_MS__OR2_2%X N_X_M1001_s N_X_M1002_d X X X X X
+ PM_SKY130_FD_SC_MS__OR2_2%X
x_PM_SKY130_FD_SC_MS__OR2_2%VGND N_VGND_M1003_s N_VGND_M1005_d N_VGND_M1006_d
+ N_VGND_c_280_n N_VGND_c_281_n N_VGND_c_282_n N_VGND_c_283_n N_VGND_c_284_n
+ VGND N_VGND_c_285_n N_VGND_c_286_n N_VGND_c_287_n N_VGND_c_288_n
+ PM_SKY130_FD_SC_MS__OR2_2%VGND
cc_1 VNB N_B_M1004_g 0.00908107f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.34
cc_2 VNB N_B_c_52_n 0.0205953f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.22
cc_3 VNB B 0.00785817f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_B_c_54_n 0.0586058f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.385
cc_5 VNB N_A_M1005_g 0.0238971f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.79
cc_6 VNB N_A_c_78_n 0.0238743f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.385
cc_7 VNB N_A_c_79_n 0.00542652f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.385
cc_8 VNB N_A_27_368#_M1002_g 0.00135811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_368#_M1001_g 0.0218443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_368#_M1006_g 0.0260244f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_11 VNB N_A_27_368#_M1007_g 0.00171063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_368#_c_126_n 0.00241395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_368#_c_127_n 0.00412876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_368#_c_128_n 0.00278905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_368#_c_129_n 0.00349145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_368#_c_130_n 0.00121168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_368#_c_131_n 0.00841735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_368#_c_132_n 0.0821122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_224_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB X 0.00356546f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.79
cc_21 VNB N_VGND_c_280_n 0.0120573f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_22 VNB N_VGND_c_281_n 0.0358796f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_23 VNB N_VGND_c_282_n 0.00647256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_283_n 0.0117383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_284_n 0.0441433f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_26 VNB N_VGND_c_285_n 0.0175968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_286_n 0.0168532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_287_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_288_n 0.164475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VPB N_B_M1004_g 0.0300626f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.34
cc_31 VPB N_A_M1000_g 0.019689f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.34
cc_32 VPB N_A_c_78_n 0.00592259f $X=-0.19 $Y=1.66 $X2=0.49 $Y2=1.385
cc_33 VPB N_A_c_79_n 0.00277411f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.385
cc_34 VPB N_A_27_368#_M1002_g 0.0236768f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_A_27_368#_M1007_g 0.0249238f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_A_27_368#_c_135_n 0.0214518f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_A_27_368#_c_136_n 0.017341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_A_27_368#_c_129_n 0.00111195f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_A_27_368#_c_138_n 0.00748573f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A_27_368#_c_130_n 0.0246694f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_A_27_368#_c_140_n 0.0071123f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_225_n 0.0102729f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_226_n 0.0119967f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_44 VPB N_VPWR_c_227_n 0.0208602f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_228_n 0.033055f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_46 VPB N_VPWR_c_229_n 0.0183953f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_230_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_224_n 0.0598866f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB X 0.00209756f $X=-0.19 $Y=1.66 $X2=0.49 $Y2=0.79
cc_50 VPB X 5.28466e-19 $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_51 N_B_M1004_g N_A_M1000_g 0.0495275f $X=0.495 $Y=2.34 $X2=0 $Y2=0
cc_52 N_B_c_52_n N_A_M1005_g 0.00980177f $X=0.49 $Y=1.22 $X2=0 $Y2=0
cc_53 B N_A_M1005_g 7.98305e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_54 N_B_c_54_n N_A_M1005_g 0.00662485f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_55 N_B_c_54_n N_A_c_78_n 0.0495275f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_56 B N_A_c_79_n 0.0161951f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_57 N_B_c_54_n N_A_c_79_n 0.0107812f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_58 N_B_M1004_g N_A_27_368#_c_135_n 0.00765481f $X=0.495 $Y=2.34 $X2=0 $Y2=0
cc_59 B N_A_27_368#_c_135_n 0.0196739f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_60 N_B_c_54_n N_A_27_368#_c_135_n 0.00223706f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_61 N_B_M1004_g N_A_27_368#_c_136_n 0.00768334f $X=0.495 $Y=2.34 $X2=0 $Y2=0
cc_62 N_B_M1004_g N_A_27_368#_c_145_n 0.0138299f $X=0.495 $Y=2.34 $X2=0 $Y2=0
cc_63 N_B_c_52_n N_A_27_368#_c_128_n 0.00218762f $X=0.49 $Y=1.22 $X2=0 $Y2=0
cc_64 N_B_M1004_g N_A_27_368#_c_140_n 4.64231e-19 $X=0.495 $Y=2.34 $X2=0 $Y2=0
cc_65 N_B_M1004_g N_VPWR_c_228_n 0.00567889f $X=0.495 $Y=2.34 $X2=0 $Y2=0
cc_66 N_B_M1004_g N_VPWR_c_224_n 0.00610055f $X=0.495 $Y=2.34 $X2=0 $Y2=0
cc_67 N_B_c_52_n N_VGND_c_281_n 0.0148675f $X=0.49 $Y=1.22 $X2=0 $Y2=0
cc_68 B N_VGND_c_281_n 0.0246129f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_69 N_B_c_54_n N_VGND_c_281_n 0.00198461f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_70 N_B_c_52_n N_VGND_c_285_n 0.00421418f $X=0.49 $Y=1.22 $X2=0 $Y2=0
cc_71 N_B_c_52_n N_VGND_c_288_n 0.00432128f $X=0.49 $Y=1.22 $X2=0 $Y2=0
cc_72 N_A_M1000_g N_A_27_368#_M1002_g 0.0352119f $X=0.885 $Y=2.34 $X2=0 $Y2=0
cc_73 N_A_c_79_n N_A_27_368#_M1002_g 0.00138818f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_74 N_A_M1005_g N_A_27_368#_M1001_g 0.0224491f $X=0.92 $Y=0.79 $X2=0 $Y2=0
cc_75 N_A_M1000_g N_A_27_368#_c_135_n 0.0010561f $X=0.885 $Y=2.34 $X2=0 $Y2=0
cc_76 N_A_c_79_n N_A_27_368#_c_135_n 0.013208f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_77 N_A_M1000_g N_A_27_368#_c_136_n 0.0013909f $X=0.885 $Y=2.34 $X2=0 $Y2=0
cc_78 N_A_M1000_g N_A_27_368#_c_145_n 0.0132832f $X=0.885 $Y=2.34 $X2=0 $Y2=0
cc_79 N_A_c_78_n N_A_27_368#_c_145_n 0.00200733f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_80 N_A_c_79_n N_A_27_368#_c_145_n 0.0224983f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_81 N_A_M1005_g N_A_27_368#_c_126_n 0.00781094f $X=0.92 $Y=0.79 $X2=0 $Y2=0
cc_82 N_A_M1005_g N_A_27_368#_c_127_n 0.0113358f $X=0.92 $Y=0.79 $X2=0 $Y2=0
cc_83 N_A_c_78_n N_A_27_368#_c_127_n 0.00338829f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_84 N_A_c_79_n N_A_27_368#_c_127_n 0.0134037f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_85 N_A_M1005_g N_A_27_368#_c_128_n 0.00137818f $X=0.92 $Y=0.79 $X2=0 $Y2=0
cc_86 N_A_c_78_n N_A_27_368#_c_128_n 3.91013e-19 $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_87 N_A_c_79_n N_A_27_368#_c_128_n 0.0229711f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_88 N_A_M1000_g N_A_27_368#_c_129_n 0.00470061f $X=0.885 $Y=2.34 $X2=0 $Y2=0
cc_89 N_A_M1005_g N_A_27_368#_c_129_n 0.00340254f $X=0.92 $Y=0.79 $X2=0 $Y2=0
cc_90 N_A_c_78_n N_A_27_368#_c_129_n 0.00204642f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_91 N_A_c_79_n N_A_27_368#_c_129_n 0.0625705f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_92 N_A_M1005_g N_A_27_368#_c_132_n 0.00157274f $X=0.92 $Y=0.79 $X2=0 $Y2=0
cc_93 N_A_c_78_n N_A_27_368#_c_132_n 0.0204574f $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_94 N_A_c_79_n N_A_27_368#_c_132_n 2.84616e-19 $X=0.96 $Y=1.515 $X2=0 $Y2=0
cc_95 N_A_c_79_n A_117_368# 0.00106497f $X=0.96 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_96 N_A_c_79_n N_VPWR_M1000_d 0.00288519f $X=0.96 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_97 N_A_M1000_g N_VPWR_c_225_n 0.00605343f $X=0.885 $Y=2.34 $X2=0 $Y2=0
cc_98 N_A_M1000_g N_VPWR_c_228_n 0.0059286f $X=0.885 $Y=2.34 $X2=0 $Y2=0
cc_99 N_A_M1000_g N_VPWR_c_224_n 0.00610055f $X=0.885 $Y=2.34 $X2=0 $Y2=0
cc_100 N_A_M1005_g N_VGND_c_281_n 5.06989e-19 $X=0.92 $Y=0.79 $X2=0 $Y2=0
cc_101 N_A_M1005_g N_VGND_c_282_n 0.00365474f $X=0.92 $Y=0.79 $X2=0 $Y2=0
cc_102 N_A_M1005_g N_VGND_c_285_n 0.00485498f $X=0.92 $Y=0.79 $X2=0 $Y2=0
cc_103 N_A_M1005_g N_VGND_c_288_n 0.00514438f $X=0.92 $Y=0.79 $X2=0 $Y2=0
cc_104 N_A_27_368#_c_145_n A_117_368# 0.00295057f $X=1.215 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_105 N_A_27_368#_c_145_n N_VPWR_M1000_d 0.00678223f $X=1.215 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_106 N_A_27_368#_c_129_n N_VPWR_M1000_d 0.00472713f $X=1.3 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_107 N_A_27_368#_c_174_p N_VPWR_M1000_d 6.76789e-19 $X=1.3 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_108 N_A_27_368#_c_138_n N_VPWR_M1007_s 0.00479283f $X=2.125 $Y=2.405 $X2=0
+ $Y2=0
cc_109 N_A_27_368#_c_130_n N_VPWR_M1007_s 0.00841337f $X=2.21 $Y=2.32 $X2=0
+ $Y2=0
cc_110 N_A_27_368#_M1002_g N_VPWR_c_225_n 0.0119276f $X=1.425 $Y=2.4 $X2=0 $Y2=0
cc_111 N_A_27_368#_M1007_g N_VPWR_c_225_n 0.00127857f $X=1.895 $Y=2.4 $X2=0
+ $Y2=0
cc_112 N_A_27_368#_c_136_n N_VPWR_c_225_n 0.00576986f $X=0.27 $Y=2.695 $X2=0
+ $Y2=0
cc_113 N_A_27_368#_c_145_n N_VPWR_c_225_n 0.0142094f $X=1.215 $Y=2.405 $X2=0
+ $Y2=0
cc_114 N_A_27_368#_c_174_p N_VPWR_c_225_n 0.0078538f $X=1.3 $Y=2.405 $X2=0 $Y2=0
cc_115 N_A_27_368#_M1002_g N_VPWR_c_227_n 0.00127857f $X=1.425 $Y=2.4 $X2=0
+ $Y2=0
cc_116 N_A_27_368#_M1007_g N_VPWR_c_227_n 0.0120007f $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_117 N_A_27_368#_c_138_n N_VPWR_c_227_n 0.0227017f $X=2.125 $Y=2.405 $X2=0
+ $Y2=0
cc_118 N_A_27_368#_c_136_n N_VPWR_c_228_n 0.00975961f $X=0.27 $Y=2.695 $X2=0
+ $Y2=0
cc_119 N_A_27_368#_M1002_g N_VPWR_c_229_n 0.00460063f $X=1.425 $Y=2.4 $X2=0
+ $Y2=0
cc_120 N_A_27_368#_M1007_g N_VPWR_c_229_n 0.00460063f $X=1.895 $Y=2.4 $X2=0
+ $Y2=0
cc_121 N_A_27_368#_M1002_g N_VPWR_c_224_n 0.00461026f $X=1.425 $Y=2.4 $X2=0
+ $Y2=0
cc_122 N_A_27_368#_M1007_g N_VPWR_c_224_n 0.00461061f $X=1.895 $Y=2.4 $X2=0
+ $Y2=0
cc_123 N_A_27_368#_c_136_n N_VPWR_c_224_n 0.0111753f $X=0.27 $Y=2.695 $X2=0
+ $Y2=0
cc_124 N_A_27_368#_c_145_n N_VPWR_c_224_n 0.0202141f $X=1.215 $Y=2.405 $X2=0
+ $Y2=0
cc_125 N_A_27_368#_c_138_n N_VPWR_c_224_n 0.0192277f $X=2.125 $Y=2.405 $X2=0
+ $Y2=0
cc_126 N_A_27_368#_c_174_p N_VPWR_c_224_n 0.00118003f $X=1.3 $Y=2.405 $X2=0
+ $Y2=0
cc_127 N_A_27_368#_c_138_n N_X_M1002_d 0.00533145f $X=2.125 $Y=2.405 $X2=0 $Y2=0
cc_128 N_A_27_368#_M1002_g X 0.00162375f $X=1.425 $Y=2.4 $X2=0 $Y2=0
cc_129 N_A_27_368#_M1001_g X 0.00175981f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A_27_368#_M1006_g X 0.0173853f $X=1.855 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A_27_368#_M1007_g X 0.00206483f $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_132 N_A_27_368#_c_127_n X 0.0099082f $X=1.215 $Y=1.095 $X2=0 $Y2=0
cc_133 N_A_27_368#_c_129_n X 0.0575862f $X=1.3 $Y=2.32 $X2=0 $Y2=0
cc_134 N_A_27_368#_c_130_n X 0.00920493f $X=2.21 $Y=2.32 $X2=0 $Y2=0
cc_135 N_A_27_368#_c_131_n X 0.0241749f $X=2.13 $Y=1.465 $X2=0 $Y2=0
cc_136 N_A_27_368#_c_132_n X 0.0212739f $X=2.13 $Y=1.465 $X2=0 $Y2=0
cc_137 N_A_27_368#_M1007_g X 0.00687034f $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_138 N_A_27_368#_c_138_n X 0.0163632f $X=2.125 $Y=2.405 $X2=0 $Y2=0
cc_139 N_A_27_368#_c_130_n X 0.0159954f $X=2.21 $Y=2.32 $X2=0 $Y2=0
cc_140 N_A_27_368#_c_127_n N_VGND_M1005_d 0.00267951f $X=1.215 $Y=1.095 $X2=0
+ $Y2=0
cc_141 N_A_27_368#_c_126_n N_VGND_c_281_n 0.0204407f $X=0.705 $Y=0.615 $X2=0
+ $Y2=0
cc_142 N_A_27_368#_M1001_g N_VGND_c_282_n 0.0111891f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_143 N_A_27_368#_M1006_g N_VGND_c_282_n 5.12656e-19 $X=1.855 $Y=0.74 $X2=0
+ $Y2=0
cc_144 N_A_27_368#_c_126_n N_VGND_c_282_n 0.0139492f $X=0.705 $Y=0.615 $X2=0
+ $Y2=0
cc_145 N_A_27_368#_c_127_n N_VGND_c_282_n 0.0208721f $X=1.215 $Y=1.095 $X2=0
+ $Y2=0
cc_146 N_A_27_368#_M1006_g N_VGND_c_284_n 0.0185053f $X=1.855 $Y=0.74 $X2=0
+ $Y2=0
cc_147 N_A_27_368#_c_131_n N_VGND_c_284_n 0.0281178f $X=2.13 $Y=1.465 $X2=0
+ $Y2=0
cc_148 N_A_27_368#_c_132_n N_VGND_c_284_n 0.00255514f $X=2.13 $Y=1.465 $X2=0
+ $Y2=0
cc_149 N_A_27_368#_c_126_n N_VGND_c_285_n 0.0078096f $X=0.705 $Y=0.615 $X2=0
+ $Y2=0
cc_150 N_A_27_368#_M1001_g N_VGND_c_286_n 0.00383152f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_151 N_A_27_368#_M1006_g N_VGND_c_286_n 0.00445602f $X=1.855 $Y=0.74 $X2=0
+ $Y2=0
cc_152 N_A_27_368#_M1001_g N_VGND_c_288_n 0.0075754f $X=1.425 $Y=0.74 $X2=0
+ $Y2=0
cc_153 N_A_27_368#_M1006_g N_VGND_c_288_n 0.00860452f $X=1.855 $Y=0.74 $X2=0
+ $Y2=0
cc_154 N_A_27_368#_c_126_n N_VGND_c_288_n 0.0085649f $X=0.705 $Y=0.615 $X2=0
+ $Y2=0
cc_155 X N_VGND_c_282_n 0.0177481f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_156 X N_VGND_c_284_n 0.0287813f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_157 X N_VGND_c_286_n 0.0105779f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_158 X N_VGND_c_288_n 0.00872261f $X=1.595 $Y=0.47 $X2=0 $Y2=0

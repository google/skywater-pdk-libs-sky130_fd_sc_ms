* File: sky130_fd_sc_ms__nor4b_1.pxi.spice
* Created: Wed Sep  2 12:16:57 2020
* 
x_PM_SKY130_FD_SC_MS__NOR4B_1%D_N N_D_N_M1008_g N_D_N_M1004_g D_N N_D_N_c_64_n
+ PM_SKY130_FD_SC_MS__NOR4B_1%D_N
x_PM_SKY130_FD_SC_MS__NOR4B_1%A N_A_M1006_g N_A_M1009_g A N_A_c_99_n N_A_c_100_n
+ PM_SKY130_FD_SC_MS__NOR4B_1%A
x_PM_SKY130_FD_SC_MS__NOR4B_1%B N_B_M1001_g N_B_M1003_g B N_B_c_136_n
+ N_B_c_137_n PM_SKY130_FD_SC_MS__NOR4B_1%B
x_PM_SKY130_FD_SC_MS__NOR4B_1%C N_C_M1007_g N_C_M1000_g C N_C_c_174_n
+ N_C_c_175_n PM_SKY130_FD_SC_MS__NOR4B_1%C
x_PM_SKY130_FD_SC_MS__NOR4B_1%A_57_368# N_A_57_368#_M1004_s N_A_57_368#_M1008_s
+ N_A_57_368#_M1002_g N_A_57_368#_M1005_g N_A_57_368#_c_224_n
+ N_A_57_368#_c_218_n N_A_57_368#_c_213_n N_A_57_368#_c_219_n
+ N_A_57_368#_c_214_n N_A_57_368#_c_221_n N_A_57_368#_c_215_n
+ N_A_57_368#_c_216_n PM_SKY130_FD_SC_MS__NOR4B_1%A_57_368#
x_PM_SKY130_FD_SC_MS__NOR4B_1%VPWR N_VPWR_M1008_d N_VPWR_c_290_n N_VPWR_c_291_n
+ N_VPWR_c_292_n VPWR N_VPWR_c_293_n N_VPWR_c_289_n
+ PM_SKY130_FD_SC_MS__NOR4B_1%VPWR
x_PM_SKY130_FD_SC_MS__NOR4B_1%Y N_Y_M1009_d N_Y_M1000_d N_Y_M1005_d N_Y_c_319_n
+ N_Y_c_320_n N_Y_c_321_n N_Y_c_322_n N_Y_c_323_n N_Y_c_324_n Y Y Y N_Y_c_325_n
+ PM_SKY130_FD_SC_MS__NOR4B_1%Y
x_PM_SKY130_FD_SC_MS__NOR4B_1%VGND N_VGND_M1004_d N_VGND_M1003_d N_VGND_M1002_d
+ N_VGND_c_380_n N_VGND_c_381_n N_VGND_c_382_n N_VGND_c_383_n N_VGND_c_384_n
+ N_VGND_c_385_n N_VGND_c_386_n N_VGND_c_387_n VGND N_VGND_c_388_n
+ N_VGND_c_389_n PM_SKY130_FD_SC_MS__NOR4B_1%VGND
cc_1 VNB N_D_N_M1008_g 0.0134167f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.26
cc_2 VNB N_D_N_M1004_g 0.0280622f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.645
cc_3 VNB D_N 0.00776204f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_D_N_c_64_n 0.0354648f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.275
cc_5 VNB N_A_M1009_g 0.0259031f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.645
cc_6 VNB N_A_c_99_n 0.0265536f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.275
cc_7 VNB N_A_c_100_n 0.00355186f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.275
cc_8 VNB N_B_M1003_g 0.0258898f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.645
cc_9 VNB N_B_c_136_n 0.0262325f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.275
cc_10 VNB N_B_c_137_n 0.00165719f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.275
cc_11 VNB N_C_M1000_g 0.0258908f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.645
cc_12 VNB N_C_c_174_n 0.0242452f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.275
cc_13 VNB N_C_c_175_n 0.00381276f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.275
cc_14 VNB N_A_57_368#_M1002_g 0.0264924f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_15 VNB N_A_57_368#_c_213_n 0.0401545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_57_368#_c_214_n 0.0356004f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_57_368#_c_215_n 0.00512013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_57_368#_c_216_n 0.0273053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_289_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_319_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.275
cc_21 VNB N_Y_c_320_n 0.00823886f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.11
cc_22 VNB N_Y_c_321_n 0.0090164f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.44
cc_23 VNB N_Y_c_322_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.275
cc_24 VNB N_Y_c_323_n 0.0181248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_324_n 0.00775352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_325_n 0.0230123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_380_n 0.0134539f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.275
cc_28 VNB N_VGND_c_381_n 0.00907103f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.275
cc_29 VNB N_VGND_c_382_n 0.0158851f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.275
cc_30 VNB N_VGND_c_383_n 0.0313058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_384_n 0.0232674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_385_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_386_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_387_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_388_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_389_n 0.211126f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VPB N_D_N_M1008_g 0.0288699f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.26
cc_38 VPB N_A_M1006_g 0.0233108f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.26
cc_39 VPB N_A_c_99_n 0.00565213f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.275
cc_40 VPB N_A_c_100_n 0.00248627f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.275
cc_41 VPB N_B_M1001_g 0.0216209f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.26
cc_42 VPB N_B_c_136_n 0.00559488f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.275
cc_43 VPB N_B_c_137_n 0.00268169f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.275
cc_44 VPB N_C_M1007_g 0.0232209f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.26
cc_45 VPB N_C_c_174_n 0.00547464f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.275
cc_46 VPB N_C_c_175_n 0.00299982f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.275
cc_47 VPB N_A_57_368#_M1005_g 0.0269122f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.275
cc_48 VPB N_A_57_368#_c_218_n 0.00141324f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_57_368#_c_219_n 0.0218206f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_57_368#_c_214_n 0.00813055f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A_57_368#_c_221_n 0.032593f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_57_368#_c_215_n 4.03371e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_57_368#_c_216_n 0.00763791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_290_n 0.0169528f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=0.645
cc_55 VPB N_VPWR_c_291_n 0.0265205f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_56 VPB N_VPWR_c_292_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_293_n 0.0689598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_289_n 0.101036f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB Y 0.048721f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_Y_c_325_n 0.00902776f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 N_D_N_M1008_g N_A_M1006_g 0.0244596f $X=0.655 $Y=2.26 $X2=0 $Y2=0
cc_62 N_D_N_M1004_g N_A_M1009_g 0.0184418f $X=0.67 $Y=0.645 $X2=0 $Y2=0
cc_63 D_N N_A_M1009_g 0.00400388f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_64 N_D_N_c_64_n N_A_M1009_g 0.00644195f $X=0.61 $Y=1.275 $X2=0 $Y2=0
cc_65 N_D_N_M1008_g N_A_c_99_n 0.0135411f $X=0.655 $Y=2.26 $X2=0 $Y2=0
cc_66 D_N N_A_c_99_n 5.07587e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_67 N_D_N_c_64_n N_A_c_99_n 0.00563717f $X=0.61 $Y=1.275 $X2=0 $Y2=0
cc_68 N_D_N_M1008_g N_A_c_100_n 0.00385965f $X=0.655 $Y=2.26 $X2=0 $Y2=0
cc_69 D_N N_A_c_100_n 0.00714274f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_70 N_D_N_M1008_g N_A_57_368#_c_224_n 0.0158258f $X=0.655 $Y=2.26 $X2=0 $Y2=0
cc_71 D_N N_A_57_368#_c_224_n 0.00581508f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_72 N_D_N_M1004_g N_A_57_368#_c_213_n 0.0111596f $X=0.67 $Y=0.645 $X2=0 $Y2=0
cc_73 D_N N_A_57_368#_c_213_n 0.0144068f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_74 N_D_N_c_64_n N_A_57_368#_c_213_n 0.00359014f $X=0.61 $Y=1.275 $X2=0 $Y2=0
cc_75 N_D_N_M1008_g N_A_57_368#_c_219_n 0.00488975f $X=0.655 $Y=2.26 $X2=0 $Y2=0
cc_76 D_N N_A_57_368#_c_219_n 0.00677334f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_77 N_D_N_c_64_n N_A_57_368#_c_219_n 0.00245637f $X=0.61 $Y=1.275 $X2=0 $Y2=0
cc_78 N_D_N_M1008_g N_A_57_368#_c_214_n 0.0116522f $X=0.655 $Y=2.26 $X2=0 $Y2=0
cc_79 N_D_N_M1004_g N_A_57_368#_c_214_n 0.0049454f $X=0.67 $Y=0.645 $X2=0 $Y2=0
cc_80 D_N N_A_57_368#_c_214_n 0.0249903f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_81 N_D_N_c_64_n N_A_57_368#_c_214_n 0.00231223f $X=0.61 $Y=1.275 $X2=0 $Y2=0
cc_82 N_D_N_M1008_g N_A_57_368#_c_221_n 0.0134806f $X=0.655 $Y=2.26 $X2=0 $Y2=0
cc_83 N_D_N_M1008_g N_VPWR_c_290_n 0.00693742f $X=0.655 $Y=2.26 $X2=0 $Y2=0
cc_84 N_D_N_M1008_g N_VPWR_c_291_n 0.00465228f $X=0.655 $Y=2.26 $X2=0 $Y2=0
cc_85 N_D_N_M1008_g N_VPWR_c_289_n 0.00555093f $X=0.655 $Y=2.26 $X2=0 $Y2=0
cc_86 N_D_N_M1004_g N_Y_c_319_n 4.34666e-19 $X=0.67 $Y=0.645 $X2=0 $Y2=0
cc_87 N_D_N_M1004_g N_Y_c_321_n 4.50506e-19 $X=0.67 $Y=0.645 $X2=0 $Y2=0
cc_88 D_N N_Y_c_321_n 0.00269803f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_89 N_D_N_M1004_g N_VGND_c_380_n 0.00693523f $X=0.67 $Y=0.645 $X2=0 $Y2=0
cc_90 D_N N_VGND_c_380_n 0.00212308f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_91 N_D_N_M1004_g N_VGND_c_384_n 0.00433162f $X=0.67 $Y=0.645 $X2=0 $Y2=0
cc_92 N_D_N_M1004_g N_VGND_c_389_n 0.00821785f $X=0.67 $Y=0.645 $X2=0 $Y2=0
cc_93 N_A_M1006_g N_B_M1001_g 0.0789063f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_94 N_A_M1009_g N_B_M1003_g 0.019972f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_95 N_A_c_99_n N_B_c_136_n 0.0201104f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_96 N_A_c_100_n N_B_c_136_n 0.00114936f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_97 N_A_M1006_g N_B_c_137_n 5.64277e-19 $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_98 N_A_c_99_n N_B_c_137_n 0.00114936f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_99 N_A_c_100_n N_B_c_137_n 0.0276387f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_100 N_A_M1006_g N_A_57_368#_c_224_n 0.0165696f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_101 N_A_c_99_n N_A_57_368#_c_224_n 7.08634e-19 $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_102 N_A_c_100_n N_A_57_368#_c_224_n 0.0229716f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_103 N_A_M1006_g N_A_57_368#_c_219_n 0.00136424f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_104 N_A_M1006_g N_VPWR_c_290_n 0.0185439f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_105 N_A_M1006_g N_VPWR_c_293_n 0.00460063f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A_M1006_g N_VPWR_c_289_n 0.00908371f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_107 N_A_M1009_g N_Y_c_319_n 0.00863911f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_108 N_A_M1009_g N_Y_c_321_n 0.00453747f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_109 N_A_c_100_n N_Y_c_321_n 0.00196319f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_110 N_A_M1009_g N_VGND_c_380_n 0.00545144f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_111 N_A_c_99_n N_VGND_c_380_n 8.85031e-19 $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_112 N_A_c_100_n N_VGND_c_380_n 0.00542787f $X=1.15 $Y=1.515 $X2=0 $Y2=0
cc_113 N_A_M1009_g N_VGND_c_386_n 0.00434272f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_114 N_A_M1009_g N_VGND_c_389_n 0.0082141f $X=1.24 $Y=0.74 $X2=0 $Y2=0
cc_115 N_B_M1001_g N_C_M1007_g 0.0611181f $X=1.645 $Y=2.4 $X2=0 $Y2=0
cc_116 N_B_c_137_n N_C_M1007_g 3.56938e-19 $X=1.69 $Y=1.515 $X2=0 $Y2=0
cc_117 N_B_M1003_g N_C_M1000_g 0.0252177f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_118 N_B_c_136_n N_C_c_174_n 0.0206935f $X=1.69 $Y=1.515 $X2=0 $Y2=0
cc_119 N_B_c_137_n N_C_c_174_n 3.99347e-19 $X=1.69 $Y=1.515 $X2=0 $Y2=0
cc_120 N_B_M1001_g N_C_c_175_n 2.87335e-19 $X=1.645 $Y=2.4 $X2=0 $Y2=0
cc_121 N_B_c_136_n N_C_c_175_n 0.00188716f $X=1.69 $Y=1.515 $X2=0 $Y2=0
cc_122 N_B_c_137_n N_C_c_175_n 0.0318721f $X=1.69 $Y=1.515 $X2=0 $Y2=0
cc_123 N_B_M1001_g N_A_57_368#_c_224_n 0.0172246f $X=1.645 $Y=2.4 $X2=0 $Y2=0
cc_124 N_B_c_136_n N_A_57_368#_c_224_n 5.44636e-19 $X=1.69 $Y=1.515 $X2=0 $Y2=0
cc_125 N_B_c_137_n N_A_57_368#_c_224_n 0.0219071f $X=1.69 $Y=1.515 $X2=0 $Y2=0
cc_126 N_B_M1001_g N_VPWR_c_290_n 0.00385865f $X=1.645 $Y=2.4 $X2=0 $Y2=0
cc_127 N_B_M1001_g N_VPWR_c_293_n 0.00553757f $X=1.645 $Y=2.4 $X2=0 $Y2=0
cc_128 N_B_M1001_g N_VPWR_c_289_n 0.0109022f $X=1.645 $Y=2.4 $X2=0 $Y2=0
cc_129 N_B_M1003_g N_Y_c_319_n 0.00969128f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_130 N_B_M1003_g N_Y_c_320_n 0.0118338f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_131 N_B_c_136_n N_Y_c_320_n 7.68393e-19 $X=1.69 $Y=1.515 $X2=0 $Y2=0
cc_132 N_B_c_137_n N_Y_c_320_n 0.0175347f $X=1.69 $Y=1.515 $X2=0 $Y2=0
cc_133 N_B_M1003_g N_Y_c_321_n 0.0015571f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_134 N_B_c_136_n N_Y_c_321_n 5.42338e-19 $X=1.69 $Y=1.515 $X2=0 $Y2=0
cc_135 N_B_c_137_n N_Y_c_321_n 0.00799991f $X=1.69 $Y=1.515 $X2=0 $Y2=0
cc_136 N_B_M1003_g N_Y_c_322_n 8.70047e-19 $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_137 N_B_M1003_g N_VGND_c_381_n 0.00491516f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_138 N_B_M1003_g N_VGND_c_386_n 0.00434272f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_139 N_B_M1003_g N_VGND_c_389_n 0.00821482f $X=1.67 $Y=0.74 $X2=0 $Y2=0
cc_140 N_C_M1000_g N_A_57_368#_M1002_g 0.0199815f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_141 N_C_M1007_g N_A_57_368#_M1005_g 0.0461884f $X=2.155 $Y=2.4 $X2=0 $Y2=0
cc_142 N_C_c_175_n N_A_57_368#_M1005_g 3.24695e-19 $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_143 N_C_M1007_g N_A_57_368#_c_224_n 0.0180436f $X=2.155 $Y=2.4 $X2=0 $Y2=0
cc_144 N_C_c_174_n N_A_57_368#_c_224_n 7.02991e-19 $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_145 N_C_c_175_n N_A_57_368#_c_224_n 0.0238723f $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_146 N_C_M1007_g N_A_57_368#_c_218_n 0.00333705f $X=2.155 $Y=2.4 $X2=0 $Y2=0
cc_147 N_C_c_175_n N_A_57_368#_c_218_n 0.0079642f $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_148 N_C_c_174_n N_A_57_368#_c_215_n 0.00187066f $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_149 N_C_c_175_n N_A_57_368#_c_215_n 0.0264357f $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_150 N_C_c_174_n N_A_57_368#_c_216_n 0.02065f $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_151 N_C_c_175_n N_A_57_368#_c_216_n 3.77186e-19 $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_152 N_C_M1007_g N_VPWR_c_293_n 0.00553757f $X=2.155 $Y=2.4 $X2=0 $Y2=0
cc_153 N_C_M1007_g N_VPWR_c_289_n 0.0109155f $X=2.155 $Y=2.4 $X2=0 $Y2=0
cc_154 N_C_M1000_g N_Y_c_319_n 8.64794e-19 $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_155 N_C_M1000_g N_Y_c_320_n 0.0118338f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_156 N_C_c_174_n N_Y_c_320_n 7.65086e-19 $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_157 N_C_c_175_n N_Y_c_320_n 0.0191575f $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_158 N_C_M1000_g N_Y_c_322_n 0.00980887f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_159 N_C_M1000_g N_Y_c_324_n 0.0015571f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_160 N_C_c_174_n N_Y_c_324_n 5.46117e-19 $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_161 N_C_c_175_n N_Y_c_324_n 0.00799991f $X=2.23 $Y=1.515 $X2=0 $Y2=0
cc_162 N_C_M1000_g N_VGND_c_381_n 0.0061968f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_163 N_C_M1000_g N_VGND_c_388_n 0.00434272f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_164 N_C_M1000_g N_VGND_c_389_n 0.00821706f $X=2.25 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A_57_368#_c_224_n N_VPWR_M1008_d 0.0117084f $X=2.565 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_166 N_A_57_368#_c_224_n N_VPWR_c_290_n 0.0218557f $X=2.565 $Y=2.035 $X2=0
+ $Y2=0
cc_167 N_A_57_368#_c_221_n N_VPWR_c_290_n 0.0251858f $X=0.35 $Y=2.035 $X2=0
+ $Y2=0
cc_168 N_A_57_368#_c_221_n N_VPWR_c_291_n 0.00991858f $X=0.35 $Y=2.035 $X2=0
+ $Y2=0
cc_169 N_A_57_368#_M1005_g N_VPWR_c_293_n 0.00553757f $X=2.725 $Y=2.4 $X2=0
+ $Y2=0
cc_170 N_A_57_368#_M1005_g N_VPWR_c_289_n 0.0109501f $X=2.725 $Y=2.4 $X2=0 $Y2=0
cc_171 N_A_57_368#_c_221_n N_VPWR_c_289_n 0.0148286f $X=0.35 $Y=2.035 $X2=0
+ $Y2=0
cc_172 N_A_57_368#_c_224_n A_263_368# 0.0096152f $X=2.565 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_173 N_A_57_368#_c_224_n A_347_368# 0.0146552f $X=2.565 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_174 N_A_57_368#_c_224_n A_449_368# 0.0180737f $X=2.565 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_175 N_A_57_368#_c_218_n A_449_368# 0.00142693f $X=2.65 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_176 N_A_57_368#_M1002_g N_Y_c_322_n 0.01371f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A_57_368#_M1002_g N_Y_c_323_n 0.0129008f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A_57_368#_c_215_n N_Y_c_323_n 0.0224209f $X=2.77 $Y=1.515 $X2=0 $Y2=0
cc_179 N_A_57_368#_c_216_n N_Y_c_323_n 0.00427209f $X=2.77 $Y=1.515 $X2=0 $Y2=0
cc_180 N_A_57_368#_M1002_g N_Y_c_324_n 0.00155819f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_181 N_A_57_368#_c_215_n N_Y_c_324_n 0.00553408f $X=2.77 $Y=1.515 $X2=0 $Y2=0
cc_182 N_A_57_368#_M1005_g Y 0.0419957f $X=2.725 $Y=2.4 $X2=0 $Y2=0
cc_183 N_A_57_368#_c_224_n Y 0.0140855f $X=2.565 $Y=2.035 $X2=0 $Y2=0
cc_184 N_A_57_368#_c_218_n Y 0.0074344f $X=2.65 $Y=1.95 $X2=0 $Y2=0
cc_185 N_A_57_368#_c_215_n Y 0.00239484f $X=2.77 $Y=1.515 $X2=0 $Y2=0
cc_186 N_A_57_368#_c_216_n Y 6.75574e-19 $X=2.77 $Y=1.515 $X2=0 $Y2=0
cc_187 N_A_57_368#_M1002_g N_Y_c_325_n 0.00477786f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_188 N_A_57_368#_M1005_g N_Y_c_325_n 0.00321217f $X=2.725 $Y=2.4 $X2=0 $Y2=0
cc_189 N_A_57_368#_c_218_n N_Y_c_325_n 0.00676433f $X=2.65 $Y=1.95 $X2=0 $Y2=0
cc_190 N_A_57_368#_c_215_n N_Y_c_325_n 0.0249903f $X=2.77 $Y=1.515 $X2=0 $Y2=0
cc_191 N_A_57_368#_c_216_n N_Y_c_325_n 0.00231223f $X=2.77 $Y=1.515 $X2=0 $Y2=0
cc_192 N_A_57_368#_c_213_n N_VGND_c_380_n 0.0252474f $X=0.455 $Y=0.645 $X2=0
+ $Y2=0
cc_193 N_A_57_368#_M1002_g N_VGND_c_383_n 0.0141934f $X=2.68 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A_57_368#_c_213_n N_VGND_c_384_n 0.0225742f $X=0.455 $Y=0.645 $X2=0
+ $Y2=0
cc_195 N_A_57_368#_M1002_g N_VGND_c_388_n 0.00434272f $X=2.68 $Y=0.74 $X2=0
+ $Y2=0
cc_196 N_A_57_368#_M1002_g N_VGND_c_389_n 0.00824301f $X=2.68 $Y=0.74 $X2=0
+ $Y2=0
cc_197 N_A_57_368#_c_213_n N_VGND_c_389_n 0.0187953f $X=0.455 $Y=0.645 $X2=0
+ $Y2=0
cc_198 N_VPWR_c_293_n Y 0.0164205f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_199 N_VPWR_c_289_n Y 0.0135915f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_200 N_Y_c_320_n N_VGND_M1003_d 0.00374272f $X=2.3 $Y=1.095 $X2=0 $Y2=0
cc_201 N_Y_c_323_n N_VGND_M1002_d 0.00411309f $X=3.105 $Y=1.095 $X2=0 $Y2=0
cc_202 N_Y_c_319_n N_VGND_c_380_n 0.0229287f $X=1.455 $Y=0.515 $X2=0 $Y2=0
cc_203 N_Y_c_319_n N_VGND_c_381_n 0.0191765f $X=1.455 $Y=0.515 $X2=0 $Y2=0
cc_204 N_Y_c_320_n N_VGND_c_381_n 0.0257093f $X=2.3 $Y=1.095 $X2=0 $Y2=0
cc_205 N_Y_c_322_n N_VGND_c_381_n 0.0183215f $X=2.465 $Y=0.515 $X2=0 $Y2=0
cc_206 N_Y_c_322_n N_VGND_c_383_n 0.0191765f $X=2.465 $Y=0.515 $X2=0 $Y2=0
cc_207 N_Y_c_323_n N_VGND_c_383_n 0.0260326f $X=3.105 $Y=1.095 $X2=0 $Y2=0
cc_208 N_Y_c_319_n N_VGND_c_386_n 0.0144922f $X=1.455 $Y=0.515 $X2=0 $Y2=0
cc_209 N_Y_c_322_n N_VGND_c_388_n 0.0144922f $X=2.465 $Y=0.515 $X2=0 $Y2=0
cc_210 N_Y_c_319_n N_VGND_c_389_n 0.0118826f $X=1.455 $Y=0.515 $X2=0 $Y2=0
cc_211 N_Y_c_322_n N_VGND_c_389_n 0.0118826f $X=2.465 $Y=0.515 $X2=0 $Y2=0

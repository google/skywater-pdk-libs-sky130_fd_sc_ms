* File: sky130_fd_sc_ms__and4b_2.pex.spice
* Created: Fri Aug 28 17:14:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__AND4B_2%A_N 3 7 9 13 16
c30 7 0 6.09845e-20 $X=0.495 $Y=0.835
r31 15 16 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.465
+ $X2=0.505 $Y2=1.465
r32 12 15 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.29 $Y=1.465
+ $X2=0.495 $Y2=1.465
r33 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.465 $X2=0.29 $Y2=1.465
r34 9 13 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.29 $Y=1.665 $X2=0.29
+ $Y2=1.465
r35 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.465
r36 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=0.835
r37 1 16 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=1.465
r38 1 3 244.887 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_2%A_186_48# 1 2 3 12 16 20 24 29 30 31 32 36
+ 40 43 45 50
c109 31 0 1.93659e-19 $X=1.78 $Y=1.045
r110 49 50 9.69969 $w=3.23e-07 $l=6.5e-08 $layer=POLY_cond $X=1.435 $Y=1.465
+ $X2=1.5 $Y2=1.465
r111 48 49 57.452 $w=3.23e-07 $l=3.85e-07 $layer=POLY_cond $X=1.05 $Y=1.465
+ $X2=1.435 $Y2=1.465
r112 47 48 6.71517 $w=3.23e-07 $l=4.5e-08 $layer=POLY_cond $X=1.005 $Y=1.465
+ $X2=1.05 $Y2=1.465
r113 44 50 8.95356 $w=3.23e-07 $l=6e-08 $layer=POLY_cond $X=1.56 $Y=1.465
+ $X2=1.5 $Y2=1.465
r114 43 46 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.587 $Y=1.465
+ $X2=1.587 $Y2=1.63
r115 43 45 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=1.587 $Y=1.465
+ $X2=1.587 $Y2=1.3
r116 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.56
+ $Y=1.465 $X2=1.56 $Y2=1.465
r117 38 40 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.905 $Y=0.96
+ $X2=3.905 $Y2=0.515
r118 34 36 50.938 $w=2.48e-07 $l=1.105e-06 $layer=LI1_cond $X=2.355 $Y=2.075
+ $X2=3.46 $Y2=2.075
r119 32 34 26.5062 $w=2.48e-07 $l=5.75e-07 $layer=LI1_cond $X=1.78 $Y=2.075
+ $X2=2.355 $Y2=2.075
r120 30 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.74 $Y=1.045
+ $X2=3.905 $Y2=0.96
r121 30 31 127.872 $w=1.68e-07 $l=1.96e-06 $layer=LI1_cond $X=3.74 $Y=1.045
+ $X2=1.78 $Y2=1.045
r122 29 32 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.695 $Y=1.95
+ $X2=1.78 $Y2=2.075
r123 29 46 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.695 $Y=1.95
+ $X2=1.695 $Y2=1.63
r124 26 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.695 $Y=1.13
+ $X2=1.78 $Y2=1.045
r125 26 45 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.695 $Y=1.13
+ $X2=1.695 $Y2=1.3
r126 22 50 16.4327 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.5 $Y=1.63
+ $X2=1.5 $Y2=1.465
r127 22 24 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.5 $Y=1.63 $X2=1.5
+ $Y2=2.4
r128 18 49 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.435 $Y=1.3
+ $X2=1.435 $Y2=1.465
r129 18 20 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.435 $Y=1.3
+ $X2=1.435 $Y2=0.74
r130 14 48 16.4327 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.05 $Y=1.63
+ $X2=1.05 $Y2=1.465
r131 14 16 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.05 $Y=1.63
+ $X2=1.05 $Y2=2.4
r132 10 47 20.7134 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.3
+ $X2=1.005 $Y2=1.465
r133 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.005 $Y=1.3
+ $X2=1.005 $Y2=0.74
r134 3 36 600 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_PDIFF $count=1 $X=3.305
+ $Y=1.84 $X2=3.46 $Y2=2.035
r135 2 34 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=2.21
+ $Y=1.84 $X2=2.355 $Y2=2.035
r136 1 40 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.765
+ $Y=0.37 $X2=3.905 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_2%D 3 7 9 12 13
c36 3 0 2.8843e-19 $X=2.12 $Y=2.34
r37 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.515
+ $X2=2.13 $Y2=1.68
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.515
+ $X2=2.13 $Y2=1.35
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.515 $X2=2.13 $Y2=1.515
r40 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.13 $Y=1.665
+ $X2=2.13 $Y2=1.515
r41 7 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.22 $Y=0.74 $X2=2.22
+ $Y2=1.35
r42 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.12 $Y=2.34 $X2=2.12
+ $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_2%C 3 7 9 12 13
c34 13 0 1.1138e-19 $X=2.67 $Y=1.515
r35 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.515
+ $X2=2.67 $Y2=1.68
r36 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.67 $Y=1.515
+ $X2=2.67 $Y2=1.35
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.515 $X2=2.67 $Y2=1.515
r38 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.67 $Y=1.665
+ $X2=2.67 $Y2=1.515
r39 7 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.61 $Y=0.74 $X2=2.61
+ $Y2=1.35
r40 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.595 $Y=2.34
+ $X2=2.595 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_2%B 3 7 9 12 13
r35 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.24 $Y=1.515
+ $X2=3.24 $Y2=1.68
r36 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.24 $Y=1.515
+ $X2=3.24 $Y2=1.35
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.24
+ $Y=1.515 $X2=3.24 $Y2=1.515
r38 9 13 4.32166 $w=3.98e-07 $l=1.5e-07 $layer=LI1_cond $X=3.205 $Y=1.665
+ $X2=3.205 $Y2=1.515
r39 7 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.215 $Y=2.34
+ $X2=3.215 $Y2=1.68
r40 3 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.15 $Y=0.74 $X2=3.15
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_2%A_27_112# 1 2 9 13 17 19 20 22 23 26 28 32
+ 34
r86 32 38 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.78 $Y=1.515
+ $X2=3.78 $Y2=1.68
r87 32 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.78 $Y=1.515
+ $X2=3.78 $Y2=1.35
r88 31 34 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=3.78 $Y=1.515 $X2=3.9
+ $Y2=1.515
r89 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.78
+ $Y=1.515 $X2=3.78 $Y2=1.515
r90 28 29 6.8562 $w=6.05e-07 $l=3.4e-07 $layer=LI1_cond $X=0.455 $Y=2.115
+ $X2=0.455 $Y2=2.455
r91 25 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.9 $Y=1.68 $X2=3.9
+ $Y2=1.515
r92 25 26 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.9 $Y=1.68 $X2=3.9
+ $Y2=2.37
r93 24 29 8.37032 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=0.795 $Y=2.455
+ $X2=0.455 $Y2=2.455
r94 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.815 $Y=2.455
+ $X2=3.9 $Y2=2.37
r95 23 24 197.027 $w=1.68e-07 $l=3.02e-06 $layer=LI1_cond $X=3.815 $Y=2.455
+ $X2=0.795 $Y2=2.455
r96 22 28 10.3924 $w=6.05e-07 $l=3.27261e-07 $layer=LI1_cond $X=0.71 $Y=1.95
+ $X2=0.455 $Y2=2.115
r97 21 22 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.71 $Y=1.13
+ $X2=0.71 $Y2=1.95
r98 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.625 $Y=1.045
+ $X2=0.71 $Y2=1.13
r99 19 20 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.625 $Y=1.045
+ $X2=0.445 $Y2=1.045
r100 15 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.96
+ $X2=0.445 $Y2=1.045
r101 15 17 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=0.28 $Y=0.96
+ $X2=0.28 $Y2=0.835
r102 13 38 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.705 $Y=2.34
+ $X2=3.705 $Y2=1.68
r103 9 37 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.69 $Y=0.74
+ $X2=3.69 $Y2=1.35
r104 2 28 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r105 1 17 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.28 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_2%VPWR 1 2 3 4 17 19 23 27 29 31 34 35 36 42
+ 47 50 54
r54 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r55 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 48 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 45 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r59 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r60 42 53 4.96106 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.85 $Y=3.33
+ $X2=4.085 $Y2=3.33
r61 42 44 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.85 $Y=3.33 $X2=3.6
+ $Y2=3.33
r62 41 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r63 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r64 38 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=3.33
+ $X2=1.81 $Y2=3.33
r65 38 40 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.975 $Y=3.33
+ $X2=2.64 $Y2=3.33
r66 36 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r67 36 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r68 34 40 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.74 $Y=3.33 $X2=2.64
+ $Y2=3.33
r69 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.74 $Y=3.33
+ $X2=2.905 $Y2=3.33
r70 33 44 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.07 $Y=3.33 $X2=3.6
+ $Y2=3.33
r71 33 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.07 $Y=3.33
+ $X2=2.905 $Y2=3.33
r72 29 53 3.01886 $w=3.55e-07 $l=1.1025e-07 $layer=LI1_cond $X=4.027 $Y=3.245
+ $X2=4.085 $Y2=3.33
r73 29 31 14.2838 $w=3.53e-07 $l=4.4e-07 $layer=LI1_cond $X=4.027 $Y=3.245
+ $X2=4.027 $Y2=2.805
r74 25 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.905 $Y=3.245
+ $X2=2.905 $Y2=3.33
r75 25 27 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=2.905 $Y=3.245
+ $X2=2.905 $Y2=2.805
r76 21 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.81 $Y=3.245
+ $X2=1.81 $Y2=3.33
r77 21 23 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=1.81 $Y=3.245
+ $X2=1.81 $Y2=2.805
r78 20 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r79 19 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.645 $Y=3.33
+ $X2=1.81 $Y2=3.33
r80 19 20 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.645 $Y=3.33
+ $X2=0.98 $Y2=3.33
r81 15 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r82 15 17 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.805
r83 4 31 600 $w=1.7e-07 $l=1.07386e-06 $layer=licon1_PDIFF $count=1 $X=3.795
+ $Y=1.84 $X2=4.025 $Y2=2.805
r84 3 27 600 $w=1.7e-07 $l=1.06936e-06 $layer=licon1_PDIFF $count=1 $X=2.685
+ $Y=1.84 $X2=2.905 $Y2=2.805
r85 2 23 600 $w=1.7e-07 $l=1.06936e-06 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=1.84 $X2=1.81 $Y2=2.805
r86 1 17 600 $w=1.7e-07 $l=1.06936e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.815 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_2%X 1 2 9 12 13 14
c37 14 0 1.7705e-19 $X=1.2 $Y=2.035
c38 13 0 6.09845e-20 $X=1.22 $Y=1.13
r39 14 16 1.81965 $w=3.78e-07 $l=6e-08 $layer=LI1_cond $X=1.2 $Y=2.01 $X2=1.14
+ $Y2=2.01
r40 12 16 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.14 $Y=1.82 $X2=1.14
+ $Y2=2.01
r41 12 13 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.14 $Y=1.82 $X2=1.14
+ $Y2=1.13
r42 7 13 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.22 $Y=0.965
+ $X2=1.22 $Y2=1.13
r43 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.22 $Y=0.965 $X2=1.22
+ $Y2=0.515
r44 2 14 600 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=1.14
+ $Y=1.84 $X2=1.275 $Y2=2.01
r45 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.08
+ $Y=0.37 $X2=1.22 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__AND4B_2%VGND 1 2 9 13 15 17 22 29 30 33 36
r44 36 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r45 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r46 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r47 27 36 12.6759 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=2.165 $Y=0 $X2=1.86
+ $Y2=0
r48 27 29 124.936 $w=1.68e-07 $l=1.915e-06 $layer=LI1_cond $X=2.165 $Y=0
+ $X2=4.08 $Y2=0
r49 26 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r50 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r51 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r52 23 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.75
+ $Y2=0
r53 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r54 22 36 12.6759 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=1.555 $Y=0 $X2=1.86
+ $Y2=0
r55 22 25 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.555 $Y=0 $X2=1.2
+ $Y2=0
r56 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r57 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r58 17 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.75
+ $Y2=0
r59 17 19 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.24
+ $Y2=0
r60 15 30 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r61 15 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r62 15 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r63 11 36 2.55884 $w=6.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.86 $Y=0.085
+ $X2=1.86 $Y2=0
r64 11 13 10.5882 $w=6.08e-07 $l=5.4e-07 $layer=LI1_cond $X=1.86 $Y=0.085
+ $X2=1.86 $Y2=0.625
r65 7 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r66 7 9 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=0.75 $Y=0.085 $X2=0.75
+ $Y2=0.625
r67 2 13 91 $w=1.7e-07 $l=6.09303e-07 $layer=licon1_NDIFF $count=2 $X=1.51
+ $Y=0.37 $X2=2.005 $Y2=0.625
r68 1 9 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=0.57 $Y=0.56
+ $X2=0.79 $Y2=0.625
.ends


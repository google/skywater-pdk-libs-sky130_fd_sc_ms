* File: sky130_fd_sc_ms__a211o_4.pxi.spice
* Created: Wed Sep  2 11:50:12 2020
* 
x_PM_SKY130_FD_SC_MS__A211O_4%A_105_280# N_A_105_280#_M1005_d
+ N_A_105_280#_M1021_d N_A_105_280#_M1002_d N_A_105_280#_M1009_d
+ N_A_105_280#_M1006_g N_A_105_280#_c_125_n N_A_105_280#_c_126_n
+ N_A_105_280#_M1011_g N_A_105_280#_M1001_g N_A_105_280#_M1015_g
+ N_A_105_280#_c_130_n N_A_105_280#_M1007_g N_A_105_280#_M1016_g
+ N_A_105_280#_c_132_n N_A_105_280#_M1008_g N_A_105_280#_c_133_n
+ N_A_105_280#_M1019_g N_A_105_280#_c_134_n N_A_105_280#_c_135_n
+ N_A_105_280#_c_136_n N_A_105_280#_c_137_n N_A_105_280#_c_149_n
+ N_A_105_280#_c_151_p N_A_105_280#_c_138_n N_A_105_280#_c_179_p
+ N_A_105_280#_c_139_n N_A_105_280#_c_140_n N_A_105_280#_c_141_n
+ N_A_105_280#_c_142_n N_A_105_280#_c_143_n
+ PM_SKY130_FD_SC_MS__A211O_4%A_105_280#
x_PM_SKY130_FD_SC_MS__A211O_4%B1 N_B1_M1010_g N_B1_M1005_g N_B1_M1018_g
+ N_B1_M1013_g N_B1_c_307_n N_B1_c_301_n N_B1_c_302_n B1 B1 N_B1_c_304_n
+ PM_SKY130_FD_SC_MS__A211O_4%B1
x_PM_SKY130_FD_SC_MS__A211O_4%C1 N_C1_M1020_g N_C1_M1009_g N_C1_M1012_g
+ N_C1_c_402_n N_C1_M1021_g C1 N_C1_c_404_n PM_SKY130_FD_SC_MS__A211O_4%C1
x_PM_SKY130_FD_SC_MS__A211O_4%A1 N_A1_M1003_g N_A1_M1002_g N_A1_M1022_g
+ N_A1_M1017_g A1 A1 A1 N_A1_c_460_n PM_SKY130_FD_SC_MS__A211O_4%A1
x_PM_SKY130_FD_SC_MS__A211O_4%A2 N_A2_M1004_g N_A2_c_509_n N_A2_c_510_n
+ N_A2_M1000_g N_A2_c_512_n N_A2_c_513_n N_A2_M1014_g N_A2_M1023_g A2
+ N_A2_c_517_n PM_SKY130_FD_SC_MS__A211O_4%A2
x_PM_SKY130_FD_SC_MS__A211O_4%VPWR N_VPWR_M1006_s N_VPWR_M1011_s N_VPWR_M1016_s
+ N_VPWR_M1004_s N_VPWR_M1022_d N_VPWR_c_573_n N_VPWR_c_574_n N_VPWR_c_575_n
+ N_VPWR_c_576_n N_VPWR_c_577_n N_VPWR_c_578_n N_VPWR_c_579_n N_VPWR_c_580_n
+ N_VPWR_c_581_n N_VPWR_c_582_n VPWR N_VPWR_c_583_n N_VPWR_c_584_n
+ N_VPWR_c_572_n N_VPWR_c_586_n N_VPWR_c_587_n N_VPWR_c_588_n
+ PM_SKY130_FD_SC_MS__A211O_4%VPWR
x_PM_SKY130_FD_SC_MS__A211O_4%X N_X_M1001_d N_X_M1008_d N_X_M1006_d N_X_M1015_d
+ N_X_c_665_n N_X_c_671_n N_X_c_666_n N_X_c_667_n N_X_c_672_n N_X_c_668_n
+ N_X_c_673_n N_X_c_695_n N_X_c_698_n N_X_c_699_n X X N_X_c_702_n N_X_c_669_n
+ PM_SKY130_FD_SC_MS__A211O_4%X
x_PM_SKY130_FD_SC_MS__A211O_4%A_517_392# N_A_517_392#_M1010_s
+ N_A_517_392#_M1018_s N_A_517_392#_M1003_s N_A_517_392#_M1014_d
+ N_A_517_392#_c_746_n N_A_517_392#_c_748_n N_A_517_392#_c_759_n
+ N_A_517_392#_c_736_n N_A_517_392#_c_768_n N_A_517_392#_c_737_n
+ N_A_517_392#_c_738_n N_A_517_392#_c_739_n N_A_517_392#_c_740_n
+ N_A_517_392#_c_741_n N_A_517_392#_c_762_n N_A_517_392#_c_742_n
+ PM_SKY130_FD_SC_MS__A211O_4%A_517_392#
x_PM_SKY130_FD_SC_MS__A211O_4%A_605_392# N_A_605_392#_M1010_d
+ N_A_605_392#_M1012_s N_A_605_392#_c_809_n
+ PM_SKY130_FD_SC_MS__A211O_4%A_605_392#
x_PM_SKY130_FD_SC_MS__A211O_4%VGND N_VGND_M1001_s N_VGND_M1007_s N_VGND_M1019_s
+ N_VGND_M1020_s N_VGND_M1013_s N_VGND_M1023_s N_VGND_c_823_n N_VGND_c_824_n
+ N_VGND_c_825_n N_VGND_c_826_n N_VGND_c_827_n N_VGND_c_828_n N_VGND_c_829_n
+ N_VGND_c_830_n N_VGND_c_831_n N_VGND_c_832_n N_VGND_c_833_n N_VGND_c_834_n
+ VGND N_VGND_c_835_n N_VGND_c_836_n N_VGND_c_837_n N_VGND_c_838_n
+ N_VGND_c_839_n N_VGND_c_840_n N_VGND_c_841_n N_VGND_c_842_n
+ PM_SKY130_FD_SC_MS__A211O_4%VGND
x_PM_SKY130_FD_SC_MS__A211O_4%A_1064_123# N_A_1064_123#_M1000_d
+ N_A_1064_123#_M1017_s N_A_1064_123#_c_927_n N_A_1064_123#_c_924_n
+ N_A_1064_123#_c_925_n PM_SKY130_FD_SC_MS__A211O_4%A_1064_123#
cc_1 VNB N_A_105_280#_M1006_g 0.00871317f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.4
cc_2 VNB N_A_105_280#_c_125_n 0.0144728f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.475
cc_3 VNB N_A_105_280#_c_126_n 0.0203032f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.475
cc_4 VNB N_A_105_280#_M1011_g 0.0057674f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.4
cc_5 VNB N_A_105_280#_M1001_g 0.0325584f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=0.74
cc_6 VNB N_A_105_280#_M1015_g 0.00579577f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=2.4
cc_7 VNB N_A_105_280#_c_130_n 0.0155441f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.22
cc_8 VNB N_A_105_280#_M1016_g 0.00734244f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=2.4
cc_9 VNB N_A_105_280#_c_132_n 0.0157624f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=1.22
cc_10 VNB N_A_105_280#_c_133_n 0.0176521f $X=-0.19 $Y=-0.245 $X2=2.49 $Y2=1.22
cc_11 VNB N_A_105_280#_c_134_n 0.0104143f $X=-0.19 $Y=-0.245 $X2=2.445 $Y2=1.34
cc_12 VNB N_A_105_280#_c_135_n 0.0815917f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=1.385
cc_13 VNB N_A_105_280#_c_136_n 0.00244339f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=2.06
cc_14 VNB N_A_105_280#_c_137_n 0.00983787f $X=-0.19 $Y=-0.245 $X2=3.04 $Y2=1.215
cc_15 VNB N_A_105_280#_c_138_n 0.00241387f $X=-0.19 $Y=-0.245 $X2=3.195
+ $Y2=0.615
cc_16 VNB N_A_105_280#_c_139_n 0.0138404f $X=-0.19 $Y=-0.245 $X2=5.725 $Y2=1.195
cc_17 VNB N_A_105_280#_c_140_n 0.00306752f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=1.34
cc_18 VNB N_A_105_280#_c_141_n 0.0042379f $X=-0.19 $Y=-0.245 $X2=3.195 $Y2=0.965
cc_19 VNB N_A_105_280#_c_142_n 0.00283233f $X=-0.19 $Y=-0.245 $X2=4.14 $Y2=0.895
cc_20 VNB N_A_105_280#_c_143_n 0.00225819f $X=-0.19 $Y=-0.245 $X2=5.89 $Y2=1.105
cc_21 VNB N_B1_M1005_g 0.0301204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B1_M1013_g 0.0248495f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.4
cc_23 VNB N_B1_c_301_n 0.00156376f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.4
cc_24 VNB N_B1_c_302_n 0.0205075f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.4
cc_25 VNB B1 0.00539681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B1_c_304_n 0.0156366f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=0.74
cc_27 VNB N_C1_M1020_g 0.0210426f $X=-0.19 $Y=-0.245 $X2=5.75 $Y2=0.615
cc_28 VNB N_C1_M1009_g 0.00209214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_C1_M1012_g 0.00180727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_C1_c_402_n 0.0176663f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.55
cc_31 VNB C1 0.00323687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_C1_c_404_n 0.0410167f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=0.74
cc_33 VNB N_A1_M1002_g 0.019291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A1_M1017_g 0.0193558f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.4
cc_35 VNB A1 0.00339878f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.55
cc_36 VNB N_A1_c_460_n 0.0271394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A2_M1004_g 0.0113836f $X=-0.19 $Y=-0.245 $X2=5.75 $Y2=0.615
cc_38 VNB N_A2_c_509_n 0.0266867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A2_c_510_n 0.0102885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A2_M1000_g 0.0116349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A2_c_512_n 0.0902248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A2_c_513_n 0.00930251f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.55
cc_43 VNB N_A2_M1014_g 0.0156508f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.4
cc_44 VNB N_A2_M1023_g 0.0375929f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.4
cc_45 VNB A2 0.0135013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A2_c_517_n 0.047283f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=0.74
cc_47 VNB N_VPWR_c_572_n 0.302998f $X=-0.19 $Y=-0.245 $X2=5.725 $Y2=1.195
cc_48 VNB N_X_c_665_n 0.00104623f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.4
cc_49 VNB N_X_c_666_n 0.00375064f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.4
cc_50 VNB N_X_c_667_n 0.0134757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_X_c_668_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.55
cc_52 VNB N_X_c_669_n 0.00209458f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=1.215
cc_53 VNB N_VGND_c_823_n 0.0358565f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=2.4
cc_54 VNB N_VGND_c_824_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.4
cc_55 VNB N_VGND_c_825_n 0.00250542f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.55
cc_56 VNB N_VGND_c_826_n 0.00634533f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.22
cc_57 VNB N_VGND_c_827_n 0.0100309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_828_n 0.0131973f $X=-0.19 $Y=-0.245 $X2=2.49 $Y2=1.22
cc_59 VNB N_VGND_c_829_n 0.0495565f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=1.34
cc_60 VNB N_VGND_c_830_n 0.0282373f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=1.385
cc_61 VNB N_VGND_c_831_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_832_n 0.0112126f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=1.55
cc_63 VNB N_VGND_c_833_n 0.0487363f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=2.06
cc_64 VNB N_VGND_c_834_n 0.00528596f $X=-0.19 $Y=-0.245 $X2=3.04 $Y2=1.215
cc_65 VNB N_VGND_c_835_n 0.0154855f $X=-0.19 $Y=-0.245 $X2=3.16 $Y2=0.615
cc_66 VNB N_VGND_c_836_n 0.0171837f $X=-0.19 $Y=-0.245 $X2=5.725 $Y2=1.195
cc_67 VNB N_VGND_c_837_n 0.0187793f $X=-0.19 $Y=-0.245 $X2=3.16 $Y2=1.215
cc_68 VNB N_VGND_c_838_n 0.422175f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.4
cc_69 VNB N_VGND_c_839_n 0.00601765f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.385
cc_70 VNB N_VGND_c_840_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=1.385
cc_71 VNB N_VGND_c_841_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_842_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1064_123#_c_924_n 0.00186167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1064_123#_c_925_n 0.00326506f $X=-0.19 $Y=-0.245 $X2=0.615
+ $Y2=1.55
cc_75 VPB N_A_105_280#_M1006_g 0.0274058f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=2.4
cc_76 VPB N_A_105_280#_M1011_g 0.0207573f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=2.4
cc_77 VPB N_A_105_280#_M1015_g 0.0213712f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=2.4
cc_78 VPB N_A_105_280#_M1016_g 0.024897f $X=-0.19 $Y=1.66 $X2=1.965 $Y2=2.4
cc_79 VPB N_A_105_280#_c_136_n 0.00764956f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=2.06
cc_80 VPB N_A_105_280#_c_149_n 0.00649353f $X=-0.19 $Y=1.66 $X2=2.615 $Y2=2.145
cc_81 VPB N_B1_M1010_g 0.0252088f $X=-0.19 $Y=1.66 $X2=5.75 $Y2=0.615
cc_82 VPB N_B1_M1018_g 0.021555f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_B1_c_307_n 0.0117614f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.475
cc_84 VPB N_B1_c_301_n 0.00229946f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=2.4
cc_85 VPB N_B1_c_302_n 0.015449f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=2.4
cc_86 VPB B1 0.00562661f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_B1_c_304_n 0.0120404f $X=-0.19 $Y=1.66 $X2=1.63 $Y2=0.74
cc_88 VPB N_C1_M1009_g 0.0280304f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_C1_M1012_g 0.027204f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A1_M1003_g 0.0253114f $X=-0.19 $Y=1.66 $X2=5.75 $Y2=0.615
cc_91 VPB N_A1_M1022_g 0.0219597f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB A1 0.00962019f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=1.55
cc_93 VPB N_A1_c_460_n 0.015998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A2_M1004_g 0.0336081f $X=-0.19 $Y=1.66 $X2=5.75 $Y2=0.615
cc_95 VPB N_A2_M1014_g 0.040877f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=2.4
cc_96 VPB N_VPWR_c_573_n 0.0141609f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_574_n 0.0646892f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.475
cc_98 VPB N_VPWR_c_575_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_576_n 0.0049754f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_577_n 0.0206041f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=2.4
cc_101 VPB N_VPWR_c_578_n 0.0102648f $X=-0.19 $Y=1.66 $X2=1.63 $Y2=0.74
cc_102 VPB N_VPWR_c_579_n 0.00609297f $X=-0.19 $Y=1.66 $X2=2.06 $Y2=1.22
cc_103 VPB N_VPWR_c_580_n 0.00329801f $X=-0.19 $Y=1.66 $X2=2.49 $Y2=0.74
cc_104 VPB N_VPWR_c_581_n 0.0160978f $X=-0.19 $Y=1.66 $X2=2.13 $Y2=1.34
cc_105 VPB N_VPWR_c_582_n 0.00601644f $X=-0.19 $Y=1.66 $X2=2.13 $Y2=1.385
cc_106 VPB N_VPWR_c_583_n 0.0680039f $X=-0.19 $Y=1.66 $X2=2.53 $Y2=1.55
cc_107 VPB N_VPWR_c_584_n 0.0233618f $X=-0.19 $Y=1.66 $X2=3.28 $Y2=0.955
cc_108 VPB N_VPWR_c_572_n 0.0989674f $X=-0.19 $Y=1.66 $X2=5.725 $Y2=1.195
cc_109 VPB N_VPWR_c_586_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_587_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_588_n 0.0125785f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_X_c_665_n 5.61158e-19 $X=-0.19 $Y=1.66 $X2=0.615 $Y2=2.4
cc_113 VPB N_X_c_671_n 0.00202354f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.475
cc_114 VPB N_X_c_672_n 0.00737223f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.4
cc_115 VPB N_X_c_673_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.63 $Y2=1.22
cc_116 VPB N_A_517_392#_c_736_n 0.00231289f $X=-0.19 $Y=1.66 $X2=1.065 $Y2=1.55
cc_117 VPB N_A_517_392#_c_737_n 0.00237722f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=0.74
cc_118 VPB N_A_517_392#_c_738_n 0.00603908f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=1.55
cc_119 VPB N_A_517_392#_c_739_n 0.0127915f $X=-0.19 $Y=1.66 $X2=1.515 $Y2=2.4
cc_120 VPB N_A_517_392#_c_740_n 0.0352797f $X=-0.19 $Y=1.66 $X2=1.63 $Y2=1.22
cc_121 VPB N_A_517_392#_c_741_n 0.0045725f $X=-0.19 $Y=1.66 $X2=1.63 $Y2=0.74
cc_122 VPB N_A_517_392#_c_742_n 0.00204906f $X=-0.19 $Y=1.66 $X2=2.49 $Y2=0.74
cc_123 VPB N_A_605_392#_c_809_n 0.00760109f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 N_A_105_280#_c_136_n N_B1_M1010_g 0.00609624f $X=2.53 $Y=2.06 $X2=0 $Y2=0
cc_125 N_A_105_280#_c_151_p N_B1_M1010_g 0.013555f $X=3.66 $Y=2.145 $X2=0 $Y2=0
cc_126 N_A_105_280#_c_133_n N_B1_M1005_g 0.0217726f $X=2.49 $Y=1.22 $X2=0 $Y2=0
cc_127 N_A_105_280#_c_135_n N_B1_M1005_g 0.00124571f $X=2.13 $Y=1.385 $X2=0
+ $Y2=0
cc_128 N_A_105_280#_c_137_n N_B1_M1005_g 0.0127351f $X=3.04 $Y=1.215 $X2=0 $Y2=0
cc_129 N_A_105_280#_c_138_n N_B1_M1005_g 0.00433283f $X=3.195 $Y=0.615 $X2=0
+ $Y2=0
cc_130 N_A_105_280#_c_140_n N_B1_M1005_g 0.00427034f $X=2.53 $Y=1.34 $X2=0 $Y2=0
cc_131 N_A_105_280#_c_141_n N_B1_M1005_g 0.006532f $X=3.195 $Y=0.965 $X2=0 $Y2=0
cc_132 N_A_105_280#_c_151_p N_B1_M1018_g 2.56637e-19 $X=3.66 $Y=2.145 $X2=0
+ $Y2=0
cc_133 N_A_105_280#_c_139_n N_B1_M1013_g 0.0147131f $X=5.725 $Y=1.195 $X2=0
+ $Y2=0
cc_134 N_A_105_280#_c_142_n N_B1_M1013_g 0.00104272f $X=4.14 $Y=0.895 $X2=0
+ $Y2=0
cc_135 N_A_105_280#_c_151_p N_B1_c_307_n 0.0456792f $X=3.66 $Y=2.145 $X2=0 $Y2=0
cc_136 N_A_105_280#_c_141_n N_B1_c_307_n 0.00784836f $X=3.195 $Y=0.965 $X2=0
+ $Y2=0
cc_137 N_A_105_280#_c_136_n N_B1_c_301_n 0.0258245f $X=2.53 $Y=2.06 $X2=0 $Y2=0
cc_138 N_A_105_280#_c_137_n N_B1_c_301_n 0.0190372f $X=3.04 $Y=1.215 $X2=0 $Y2=0
cc_139 N_A_105_280#_c_151_p N_B1_c_301_n 0.020039f $X=3.66 $Y=2.145 $X2=0 $Y2=0
cc_140 N_A_105_280#_c_140_n N_B1_c_301_n 0.00670748f $X=2.53 $Y=1.34 $X2=0 $Y2=0
cc_141 N_A_105_280#_c_141_n N_B1_c_301_n 0.00536516f $X=3.195 $Y=0.965 $X2=0
+ $Y2=0
cc_142 N_A_105_280#_M1016_g N_B1_c_302_n 0.00236036f $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_143 N_A_105_280#_c_135_n N_B1_c_302_n 0.00156693f $X=2.13 $Y=1.385 $X2=0
+ $Y2=0
cc_144 N_A_105_280#_c_136_n N_B1_c_302_n 0.00278353f $X=2.53 $Y=2.06 $X2=0 $Y2=0
cc_145 N_A_105_280#_c_137_n N_B1_c_302_n 0.00124647f $X=3.04 $Y=1.215 $X2=0
+ $Y2=0
cc_146 N_A_105_280#_c_151_p N_B1_c_302_n 9.33085e-19 $X=3.66 $Y=2.145 $X2=0
+ $Y2=0
cc_147 N_A_105_280#_c_140_n N_B1_c_302_n 7.62508e-19 $X=2.53 $Y=1.34 $X2=0 $Y2=0
cc_148 N_A_105_280#_c_141_n N_B1_c_302_n 3.87822e-19 $X=3.195 $Y=0.965 $X2=0
+ $Y2=0
cc_149 N_A_105_280#_c_139_n B1 0.0185247f $X=5.725 $Y=1.195 $X2=0 $Y2=0
cc_150 N_A_105_280#_c_142_n B1 0.023578f $X=4.14 $Y=0.895 $X2=0 $Y2=0
cc_151 N_A_105_280#_c_139_n N_B1_c_304_n 8.23223e-19 $X=5.725 $Y=1.195 $X2=0
+ $Y2=0
cc_152 N_A_105_280#_c_142_n N_B1_c_304_n 4.58199e-19 $X=4.14 $Y=0.895 $X2=0
+ $Y2=0
cc_153 N_A_105_280#_c_179_p N_C1_M1020_g 0.0158149f $X=3.96 $Y=0.955 $X2=0 $Y2=0
cc_154 N_A_105_280#_c_141_n N_C1_M1020_g 0.00318964f $X=3.195 $Y=0.965 $X2=0
+ $Y2=0
cc_155 N_A_105_280#_c_142_n N_C1_M1020_g 0.00147283f $X=4.14 $Y=0.895 $X2=0
+ $Y2=0
cc_156 N_A_105_280#_c_151_p N_C1_M1009_g 0.0099235f $X=3.66 $Y=2.145 $X2=0 $Y2=0
cc_157 N_A_105_280#_c_151_p N_C1_M1012_g 0.00335283f $X=3.66 $Y=2.145 $X2=0
+ $Y2=0
cc_158 N_A_105_280#_c_179_p N_C1_c_402_n 0.0164949f $X=3.96 $Y=0.955 $X2=0 $Y2=0
cc_159 N_A_105_280#_c_142_n N_C1_c_402_n 0.0122258f $X=4.14 $Y=0.895 $X2=0 $Y2=0
cc_160 N_A_105_280#_c_179_p C1 0.0230486f $X=3.96 $Y=0.955 $X2=0 $Y2=0
cc_161 N_A_105_280#_c_141_n C1 0.00690772f $X=3.195 $Y=0.965 $X2=0 $Y2=0
cc_162 N_A_105_280#_c_142_n C1 0.00525028f $X=4.14 $Y=0.895 $X2=0 $Y2=0
cc_163 N_A_105_280#_c_179_p N_C1_c_404_n 9.07417e-19 $X=3.96 $Y=0.955 $X2=0
+ $Y2=0
cc_164 N_A_105_280#_c_139_n N_A1_M1002_g 0.00877195f $X=5.725 $Y=1.195 $X2=0
+ $Y2=0
cc_165 N_A_105_280#_c_143_n N_A1_M1002_g 0.00357018f $X=5.89 $Y=1.105 $X2=0
+ $Y2=0
cc_166 N_A_105_280#_c_143_n N_A1_M1017_g 0.00370955f $X=5.89 $Y=1.105 $X2=0
+ $Y2=0
cc_167 N_A_105_280#_c_139_n A1 0.0599227f $X=5.725 $Y=1.195 $X2=0 $Y2=0
cc_168 N_A_105_280#_c_143_n A1 0.0254529f $X=5.89 $Y=1.105 $X2=0 $Y2=0
cc_169 N_A_105_280#_c_139_n N_A1_c_460_n 0.00184523f $X=5.725 $Y=1.195 $X2=0
+ $Y2=0
cc_170 N_A_105_280#_c_143_n N_A1_c_460_n 0.00246465f $X=5.89 $Y=1.105 $X2=0
+ $Y2=0
cc_171 N_A_105_280#_c_139_n N_A2_c_510_n 0.0146651f $X=5.725 $Y=1.195 $X2=0
+ $Y2=0
cc_172 N_A_105_280#_c_139_n N_A2_M1000_g 0.013753f $X=5.725 $Y=1.195 $X2=0 $Y2=0
cc_173 N_A_105_280#_c_143_n N_A2_M1000_g 5.447e-19 $X=5.89 $Y=1.105 $X2=0 $Y2=0
cc_174 N_A_105_280#_c_139_n A2 0.0108974f $X=5.725 $Y=1.195 $X2=0 $Y2=0
cc_175 N_A_105_280#_c_139_n N_A2_c_517_n 5.5067e-19 $X=5.725 $Y=1.195 $X2=0
+ $Y2=0
cc_176 N_A_105_280#_M1006_g N_VPWR_c_574_n 0.00517359f $X=0.615 $Y=2.4 $X2=0
+ $Y2=0
cc_177 N_A_105_280#_M1006_g N_VPWR_c_575_n 0.005209f $X=0.615 $Y=2.4 $X2=0 $Y2=0
cc_178 N_A_105_280#_M1011_g N_VPWR_c_575_n 0.00460063f $X=1.065 $Y=2.4 $X2=0
+ $Y2=0
cc_179 N_A_105_280#_M1006_g N_VPWR_c_576_n 6.56346e-19 $X=0.615 $Y=2.4 $X2=0
+ $Y2=0
cc_180 N_A_105_280#_M1011_g N_VPWR_c_576_n 0.0170371f $X=1.065 $Y=2.4 $X2=0
+ $Y2=0
cc_181 N_A_105_280#_M1015_g N_VPWR_c_576_n 0.00383761f $X=1.515 $Y=2.4 $X2=0
+ $Y2=0
cc_182 N_A_105_280#_M1015_g N_VPWR_c_577_n 0.005209f $X=1.515 $Y=2.4 $X2=0 $Y2=0
cc_183 N_A_105_280#_M1016_g N_VPWR_c_577_n 0.005209f $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_184 N_A_105_280#_M1016_g N_VPWR_c_578_n 0.00628342f $X=1.965 $Y=2.4 $X2=0
+ $Y2=0
cc_185 N_A_105_280#_c_134_n N_VPWR_c_578_n 0.010202f $X=2.445 $Y=1.34 $X2=0
+ $Y2=0
cc_186 N_A_105_280#_c_135_n N_VPWR_c_578_n 0.00412269f $X=2.13 $Y=1.385 $X2=0
+ $Y2=0
cc_187 N_A_105_280#_c_136_n N_VPWR_c_578_n 0.0177406f $X=2.53 $Y=2.06 $X2=0
+ $Y2=0
cc_188 N_A_105_280#_c_149_n N_VPWR_c_578_n 0.0141315f $X=2.615 $Y=2.145 $X2=0
+ $Y2=0
cc_189 N_A_105_280#_M1006_g N_VPWR_c_572_n 0.00986333f $X=0.615 $Y=2.4 $X2=0
+ $Y2=0
cc_190 N_A_105_280#_M1011_g N_VPWR_c_572_n 0.00908554f $X=1.065 $Y=2.4 $X2=0
+ $Y2=0
cc_191 N_A_105_280#_M1015_g N_VPWR_c_572_n 0.00982266f $X=1.515 $Y=2.4 $X2=0
+ $Y2=0
cc_192 N_A_105_280#_M1016_g N_VPWR_c_572_n 0.00987399f $X=1.965 $Y=2.4 $X2=0
+ $Y2=0
cc_193 N_A_105_280#_M1006_g N_X_c_665_n 0.00867221f $X=0.615 $Y=2.4 $X2=0 $Y2=0
cc_194 N_A_105_280#_c_125_n N_X_c_665_n 0.01145f $X=0.975 $Y=1.475 $X2=0 $Y2=0
cc_195 N_A_105_280#_c_126_n N_X_c_665_n 0.00596361f $X=0.705 $Y=1.475 $X2=0
+ $Y2=0
cc_196 N_A_105_280#_M1011_g N_X_c_665_n 0.0043762f $X=1.065 $Y=2.4 $X2=0 $Y2=0
cc_197 N_A_105_280#_M1006_g N_X_c_671_n 0.0145309f $X=0.615 $Y=2.4 $X2=0 $Y2=0
cc_198 N_A_105_280#_M1011_g N_X_c_671_n 3.68116e-19 $X=1.065 $Y=2.4 $X2=0 $Y2=0
cc_199 N_A_105_280#_c_125_n N_X_c_666_n 0.00172879f $X=0.975 $Y=1.475 $X2=0
+ $Y2=0
cc_200 N_A_105_280#_M1001_g N_X_c_666_n 0.0135219f $X=1.2 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A_105_280#_c_135_n N_X_c_666_n 0.00873843f $X=2.13 $Y=1.385 $X2=0 $Y2=0
cc_202 N_A_105_280#_c_125_n N_X_c_667_n 0.00405513f $X=0.975 $Y=1.475 $X2=0
+ $Y2=0
cc_203 N_A_105_280#_c_126_n N_X_c_667_n 0.00100704f $X=0.705 $Y=1.475 $X2=0
+ $Y2=0
cc_204 N_A_105_280#_M1011_g N_X_c_672_n 0.0163535f $X=1.065 $Y=2.4 $X2=0 $Y2=0
cc_205 N_A_105_280#_M1015_g N_X_c_672_n 0.0158893f $X=1.515 $Y=2.4 $X2=0 $Y2=0
cc_206 N_A_105_280#_M1016_g N_X_c_672_n 0.00584392f $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_207 N_A_105_280#_c_135_n N_X_c_672_n 0.00516336f $X=2.13 $Y=1.385 $X2=0 $Y2=0
cc_208 N_A_105_280#_c_136_n N_X_c_672_n 0.00331571f $X=2.53 $Y=2.06 $X2=0 $Y2=0
cc_209 N_A_105_280#_M1001_g N_X_c_668_n 3.92313e-19 $X=1.2 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A_105_280#_c_130_n N_X_c_668_n 3.92313e-19 $X=1.63 $Y=1.22 $X2=0 $Y2=0
cc_211 N_A_105_280#_M1011_g N_X_c_673_n 8.30987e-19 $X=1.065 $Y=2.4 $X2=0 $Y2=0
cc_212 N_A_105_280#_M1015_g N_X_c_673_n 0.0154511f $X=1.515 $Y=2.4 $X2=0 $Y2=0
cc_213 N_A_105_280#_M1016_g N_X_c_673_n 0.014728f $X=1.965 $Y=2.4 $X2=0 $Y2=0
cc_214 N_A_105_280#_c_132_n N_X_c_695_n 0.00952589f $X=2.06 $Y=1.22 $X2=0 $Y2=0
cc_215 N_A_105_280#_c_134_n N_X_c_695_n 0.0137302f $X=2.445 $Y=1.34 $X2=0 $Y2=0
cc_216 N_A_105_280#_c_135_n N_X_c_695_n 0.00375306f $X=2.13 $Y=1.385 $X2=0 $Y2=0
cc_217 N_A_105_280#_M1006_g N_X_c_698_n 0.00705655f $X=0.615 $Y=2.4 $X2=0 $Y2=0
cc_218 N_A_105_280#_c_134_n N_X_c_699_n 0.0150761f $X=2.445 $Y=1.34 $X2=0 $Y2=0
cc_219 N_A_105_280#_c_135_n N_X_c_699_n 6.02637e-19 $X=2.13 $Y=1.385 $X2=0 $Y2=0
cc_220 N_A_105_280#_c_130_n X 0.00785688f $X=1.63 $Y=1.22 $X2=0 $Y2=0
cc_221 N_A_105_280#_c_134_n N_X_c_702_n 0.0143588f $X=2.445 $Y=1.34 $X2=0 $Y2=0
cc_222 N_A_105_280#_c_135_n N_X_c_702_n 0.0185963f $X=2.13 $Y=1.385 $X2=0 $Y2=0
cc_223 N_A_105_280#_M1001_g N_X_c_669_n 0.00371782f $X=1.2 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A_105_280#_c_130_n N_X_c_669_n 0.00610015f $X=1.63 $Y=1.22 $X2=0 $Y2=0
cc_225 N_A_105_280#_c_132_n N_X_c_669_n 0.00449938f $X=2.06 $Y=1.22 $X2=0 $Y2=0
cc_226 N_A_105_280#_c_134_n N_X_c_669_n 0.00966603f $X=2.445 $Y=1.34 $X2=0 $Y2=0
cc_227 N_A_105_280#_c_135_n N_X_c_669_n 8.70522e-19 $X=2.13 $Y=1.385 $X2=0 $Y2=0
cc_228 N_A_105_280#_c_136_n N_A_517_392#_M1010_s 0.00135002f $X=2.53 $Y=2.06
+ $X2=-0.19 $Y2=-0.245
cc_229 N_A_105_280#_c_149_n N_A_517_392#_M1010_s 6.03208e-19 $X=2.615 $Y=2.145
+ $X2=-0.19 $Y2=-0.245
cc_230 N_A_105_280#_c_151_p N_A_517_392#_M1010_s 0.00848742f $X=3.66 $Y=2.145
+ $X2=-0.19 $Y2=-0.245
cc_231 N_A_105_280#_M1009_d N_A_517_392#_c_746_n 0.00329004f $X=3.525 $Y=1.96
+ $X2=0 $Y2=0
cc_232 N_A_105_280#_c_151_p N_A_517_392#_c_746_n 0.0506264f $X=3.66 $Y=2.145
+ $X2=0 $Y2=0
cc_233 N_A_105_280#_c_151_p N_A_517_392#_c_748_n 0.0023583f $X=3.66 $Y=2.145
+ $X2=0 $Y2=0
cc_234 N_A_105_280#_c_149_n N_A_517_392#_c_741_n 0.00604908f $X=2.615 $Y=2.145
+ $X2=0 $Y2=0
cc_235 N_A_105_280#_c_151_p N_A_517_392#_c_741_n 0.0154635f $X=3.66 $Y=2.145
+ $X2=0 $Y2=0
cc_236 N_A_105_280#_c_151_p N_A_605_392#_M1010_d 0.00433523f $X=3.66 $Y=2.145
+ $X2=-0.19 $Y2=-0.245
cc_237 N_A_105_280#_M1009_d N_A_605_392#_c_809_n 0.00168223f $X=3.525 $Y=1.96
+ $X2=0 $Y2=0
cc_238 N_A_105_280#_c_179_p N_VGND_M1020_s 0.0044804f $X=3.96 $Y=0.955 $X2=0
+ $Y2=0
cc_239 N_A_105_280#_c_139_n N_VGND_M1013_s 0.0149463f $X=5.725 $Y=1.195 $X2=0
+ $Y2=0
cc_240 N_A_105_280#_c_125_n N_VGND_c_823_n 0.00151981f $X=0.975 $Y=1.475 $X2=0
+ $Y2=0
cc_241 N_A_105_280#_M1001_g N_VGND_c_823_n 0.0138061f $X=1.2 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A_105_280#_c_130_n N_VGND_c_823_n 4.56715e-19 $X=1.63 $Y=1.22 $X2=0
+ $Y2=0
cc_243 N_A_105_280#_M1001_g N_VGND_c_824_n 0.00383152f $X=1.2 $Y=0.74 $X2=0
+ $Y2=0
cc_244 N_A_105_280#_c_130_n N_VGND_c_824_n 0.00383152f $X=1.63 $Y=1.22 $X2=0
+ $Y2=0
cc_245 N_A_105_280#_M1001_g N_VGND_c_825_n 4.05984e-19 $X=1.2 $Y=0.74 $X2=0
+ $Y2=0
cc_246 N_A_105_280#_c_130_n N_VGND_c_825_n 0.00706531f $X=1.63 $Y=1.22 $X2=0
+ $Y2=0
cc_247 N_A_105_280#_c_132_n N_VGND_c_825_n 0.00843621f $X=2.06 $Y=1.22 $X2=0
+ $Y2=0
cc_248 N_A_105_280#_c_133_n N_VGND_c_825_n 9.20677e-19 $X=2.49 $Y=1.22 $X2=0
+ $Y2=0
cc_249 N_A_105_280#_c_132_n N_VGND_c_826_n 9.69054e-19 $X=2.06 $Y=1.22 $X2=0
+ $Y2=0
cc_250 N_A_105_280#_c_133_n N_VGND_c_826_n 0.0126826f $X=2.49 $Y=1.22 $X2=0
+ $Y2=0
cc_251 N_A_105_280#_c_137_n N_VGND_c_826_n 0.0197087f $X=3.04 $Y=1.215 $X2=0
+ $Y2=0
cc_252 N_A_105_280#_c_138_n N_VGND_c_826_n 0.0189796f $X=3.195 $Y=0.615 $X2=0
+ $Y2=0
cc_253 N_A_105_280#_c_140_n N_VGND_c_826_n 0.00433174f $X=2.53 $Y=1.34 $X2=0
+ $Y2=0
cc_254 N_A_105_280#_c_138_n N_VGND_c_827_n 0.00968381f $X=3.195 $Y=0.615 $X2=0
+ $Y2=0
cc_255 N_A_105_280#_c_179_p N_VGND_c_827_n 0.0201731f $X=3.96 $Y=0.955 $X2=0
+ $Y2=0
cc_256 N_A_105_280#_c_139_n N_VGND_c_828_n 0.0218816f $X=5.725 $Y=1.195 $X2=0
+ $Y2=0
cc_257 N_A_105_280#_c_142_n N_VGND_c_828_n 0.0131078f $X=4.14 $Y=0.895 $X2=0
+ $Y2=0
cc_258 N_A_105_280#_c_132_n N_VGND_c_835_n 0.00383152f $X=2.06 $Y=1.22 $X2=0
+ $Y2=0
cc_259 N_A_105_280#_c_133_n N_VGND_c_835_n 0.00383152f $X=2.49 $Y=1.22 $X2=0
+ $Y2=0
cc_260 N_A_105_280#_c_138_n N_VGND_c_836_n 0.00751838f $X=3.195 $Y=0.615 $X2=0
+ $Y2=0
cc_261 N_A_105_280#_c_142_n N_VGND_c_837_n 0.0053849f $X=4.14 $Y=0.895 $X2=0
+ $Y2=0
cc_262 N_A_105_280#_M1001_g N_VGND_c_838_n 0.0075754f $X=1.2 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A_105_280#_c_130_n N_VGND_c_838_n 0.00373265f $X=1.63 $Y=1.22 $X2=0
+ $Y2=0
cc_264 N_A_105_280#_c_132_n N_VGND_c_838_n 0.00373475f $X=2.06 $Y=1.22 $X2=0
+ $Y2=0
cc_265 N_A_105_280#_c_133_n N_VGND_c_838_n 0.0075754f $X=2.49 $Y=1.22 $X2=0
+ $Y2=0
cc_266 N_A_105_280#_c_138_n N_VGND_c_838_n 0.00822849f $X=3.195 $Y=0.615 $X2=0
+ $Y2=0
cc_267 N_A_105_280#_c_142_n N_VGND_c_838_n 0.00883028f $X=4.14 $Y=0.895 $X2=0
+ $Y2=0
cc_268 N_A_105_280#_c_139_n N_A_1064_123#_M1000_d 0.00216063f $X=5.725 $Y=1.195
+ $X2=-0.19 $Y2=-0.245
cc_269 N_A_105_280#_M1002_d N_A_1064_123#_c_927_n 0.00407798f $X=5.75 $Y=0.615
+ $X2=0 $Y2=0
cc_270 N_A_105_280#_c_139_n N_A_1064_123#_c_927_n 0.0157791f $X=5.725 $Y=1.195
+ $X2=0 $Y2=0
cc_271 N_A_105_280#_c_143_n N_A_1064_123#_c_927_n 0.015847f $X=5.89 $Y=1.105
+ $X2=0 $Y2=0
cc_272 N_A_105_280#_c_143_n N_A_1064_123#_c_925_n 0.0100053f $X=5.89 $Y=1.105
+ $X2=0 $Y2=0
cc_273 N_B1_M1005_g N_C1_M1020_g 0.0217088f $X=2.98 $Y=0.79 $X2=0 $Y2=0
cc_274 N_B1_M1010_g N_C1_M1009_g 0.0401733f $X=2.935 $Y=2.46 $X2=0 $Y2=0
cc_275 N_B1_c_307_n N_C1_M1009_g 0.0146739f $X=3.965 $Y=1.805 $X2=0 $Y2=0
cc_276 N_B1_c_301_n N_C1_M1009_g 7.90363e-19 $X=2.94 $Y=1.635 $X2=0 $Y2=0
cc_277 N_B1_c_302_n N_C1_M1009_g 0.0100167f $X=2.94 $Y=1.635 $X2=0 $Y2=0
cc_278 B1 N_C1_M1009_g 4.51928e-19 $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_279 N_B1_M1018_g N_C1_M1012_g 0.0393625f $X=4.36 $Y=2.46 $X2=0 $Y2=0
cc_280 N_B1_c_307_n N_C1_M1012_g 0.0159438f $X=3.965 $Y=1.805 $X2=0 $Y2=0
cc_281 B1 N_C1_M1012_g 0.00774604f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_282 N_B1_M1013_g N_C1_c_402_n 0.0226577f $X=4.375 $Y=0.935 $X2=0 $Y2=0
cc_283 N_B1_M1005_g C1 9.1033e-19 $X=2.98 $Y=0.79 $X2=0 $Y2=0
cc_284 N_B1_M1013_g C1 7.59958e-19 $X=4.375 $Y=0.935 $X2=0 $Y2=0
cc_285 N_B1_c_307_n C1 0.0245545f $X=3.965 $Y=1.805 $X2=0 $Y2=0
cc_286 N_B1_c_301_n C1 0.00339543f $X=2.94 $Y=1.635 $X2=0 $Y2=0
cc_287 N_B1_c_302_n C1 2.43307e-19 $X=2.94 $Y=1.635 $X2=0 $Y2=0
cc_288 B1 C1 0.00586513f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_289 N_B1_c_307_n N_C1_c_404_n 0.00263852f $X=3.965 $Y=1.805 $X2=0 $Y2=0
cc_290 N_B1_c_301_n N_C1_c_404_n 8.77101e-19 $X=2.94 $Y=1.635 $X2=0 $Y2=0
cc_291 N_B1_c_302_n N_C1_c_404_n 0.00920115f $X=2.94 $Y=1.635 $X2=0 $Y2=0
cc_292 B1 N_C1_c_404_n 0.00626662f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_293 N_B1_c_304_n N_C1_c_404_n 0.0213772f $X=4.35 $Y=1.635 $X2=0 $Y2=0
cc_294 B1 A1 0.0139741f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_295 N_B1_M1018_g N_A2_M1004_g 0.0131521f $X=4.36 $Y=2.46 $X2=0 $Y2=0
cc_296 B1 N_A2_M1004_g 0.00237142f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_297 N_B1_M1013_g N_A2_c_510_n 0.00796009f $X=4.375 $Y=0.935 $X2=0 $Y2=0
cc_298 B1 N_A2_c_510_n 0.00126353f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_299 N_B1_c_304_n N_A2_c_510_n 0.0199049f $X=4.35 $Y=1.635 $X2=0 $Y2=0
cc_300 N_B1_M1013_g N_A2_M1000_g 0.00842148f $X=4.375 $Y=0.935 $X2=0 $Y2=0
cc_301 N_B1_M1013_g A2 3.51473e-19 $X=4.375 $Y=0.935 $X2=0 $Y2=0
cc_302 N_B1_M1013_g N_A2_c_517_n 3.35183e-19 $X=4.375 $Y=0.935 $X2=0 $Y2=0
cc_303 N_B1_M1010_g N_VPWR_c_578_n 0.012055f $X=2.935 $Y=2.46 $X2=0 $Y2=0
cc_304 N_B1_M1018_g N_VPWR_c_579_n 5.90973e-19 $X=4.36 $Y=2.46 $X2=0 $Y2=0
cc_305 N_B1_M1010_g N_VPWR_c_583_n 0.00403327f $X=2.935 $Y=2.46 $X2=0 $Y2=0
cc_306 N_B1_M1018_g N_VPWR_c_583_n 0.00397082f $X=4.36 $Y=2.46 $X2=0 $Y2=0
cc_307 N_B1_M1010_g N_VPWR_c_572_n 0.00526422f $X=2.935 $Y=2.46 $X2=0 $Y2=0
cc_308 N_B1_M1018_g N_VPWR_c_572_n 0.00515236f $X=4.36 $Y=2.46 $X2=0 $Y2=0
cc_309 N_B1_M1010_g N_A_517_392#_c_746_n 0.0109404f $X=2.935 $Y=2.46 $X2=0 $Y2=0
cc_310 N_B1_M1018_g N_A_517_392#_c_746_n 0.0115538f $X=4.36 $Y=2.46 $X2=0 $Y2=0
cc_311 N_B1_c_307_n N_A_517_392#_c_746_n 0.00385591f $X=3.965 $Y=1.805 $X2=0
+ $Y2=0
cc_312 B1 N_A_517_392#_c_746_n 0.0169253f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_313 N_B1_c_304_n N_A_517_392#_c_746_n 2.275e-19 $X=4.35 $Y=1.635 $X2=0 $Y2=0
cc_314 N_B1_M1018_g N_A_517_392#_c_748_n 0.00309198f $X=4.36 $Y=2.46 $X2=0 $Y2=0
cc_315 B1 N_A_517_392#_c_748_n 0.0113294f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_316 N_B1_c_304_n N_A_517_392#_c_748_n 2.64051e-19 $X=4.35 $Y=1.635 $X2=0
+ $Y2=0
cc_317 N_B1_M1018_g N_A_517_392#_c_759_n 0.00322616f $X=4.36 $Y=2.46 $X2=0 $Y2=0
cc_318 N_B1_M1018_g N_A_517_392#_c_736_n 2.46921e-19 $X=4.36 $Y=2.46 $X2=0 $Y2=0
cc_319 N_B1_M1010_g N_A_517_392#_c_741_n 0.00614276f $X=2.935 $Y=2.46 $X2=0
+ $Y2=0
cc_320 N_B1_M1018_g N_A_517_392#_c_762_n 0.0011968f $X=4.36 $Y=2.46 $X2=0 $Y2=0
cc_321 B1 N_A_605_392#_M1012_s 0.00481243f $X=3.995 $Y=1.95 $X2=0 $Y2=0
cc_322 N_B1_M1010_g N_A_605_392#_c_809_n 9.52217e-19 $X=2.935 $Y=2.46 $X2=0
+ $Y2=0
cc_323 N_B1_M1018_g N_A_605_392#_c_809_n 0.00398994f $X=4.36 $Y=2.46 $X2=0 $Y2=0
cc_324 N_B1_M1005_g N_VGND_c_826_n 0.00435179f $X=2.98 $Y=0.79 $X2=0 $Y2=0
cc_325 N_B1_M1005_g N_VGND_c_827_n 4.1551e-19 $X=2.98 $Y=0.79 $X2=0 $Y2=0
cc_326 N_B1_M1013_g N_VGND_c_828_n 0.00879011f $X=4.375 $Y=0.935 $X2=0 $Y2=0
cc_327 N_B1_M1005_g N_VGND_c_836_n 0.00494504f $X=2.98 $Y=0.79 $X2=0 $Y2=0
cc_328 N_B1_M1013_g N_VGND_c_837_n 0.00349617f $X=4.375 $Y=0.935 $X2=0 $Y2=0
cc_329 N_B1_M1005_g N_VGND_c_838_n 0.00514438f $X=2.98 $Y=0.79 $X2=0 $Y2=0
cc_330 N_B1_M1013_g N_VGND_c_838_n 0.00396651f $X=4.375 $Y=0.935 $X2=0 $Y2=0
cc_331 N_C1_M1009_g N_VPWR_c_583_n 0.00348345f $X=3.435 $Y=2.46 $X2=0 $Y2=0
cc_332 N_C1_M1012_g N_VPWR_c_583_n 0.00348345f $X=3.885 $Y=2.46 $X2=0 $Y2=0
cc_333 N_C1_M1009_g N_VPWR_c_572_n 0.00428872f $X=3.435 $Y=2.46 $X2=0 $Y2=0
cc_334 N_C1_M1012_g N_VPWR_c_572_n 0.00428649f $X=3.885 $Y=2.46 $X2=0 $Y2=0
cc_335 N_C1_M1009_g N_A_517_392#_c_746_n 0.0118984f $X=3.435 $Y=2.46 $X2=0 $Y2=0
cc_336 N_C1_M1012_g N_A_517_392#_c_746_n 0.0134613f $X=3.885 $Y=2.46 $X2=0 $Y2=0
cc_337 N_C1_M1012_g N_A_517_392#_c_748_n 2.6828e-19 $X=3.885 $Y=2.46 $X2=0 $Y2=0
cc_338 N_C1_M1012_g N_A_517_392#_c_759_n 7.98669e-19 $X=3.885 $Y=2.46 $X2=0
+ $Y2=0
cc_339 N_C1_M1009_g N_A_517_392#_c_741_n 6.24855e-19 $X=3.435 $Y=2.46 $X2=0
+ $Y2=0
cc_340 N_C1_M1009_g N_A_605_392#_c_809_n 0.0115554f $X=3.435 $Y=2.46 $X2=0 $Y2=0
cc_341 N_C1_M1012_g N_A_605_392#_c_809_n 0.0115809f $X=3.885 $Y=2.46 $X2=0 $Y2=0
cc_342 N_C1_M1020_g N_VGND_c_827_n 0.00758501f $X=3.41 $Y=0.79 $X2=0 $Y2=0
cc_343 N_C1_c_402_n N_VGND_c_827_n 0.00282961f $X=3.9 $Y=1.29 $X2=0 $Y2=0
cc_344 N_C1_c_402_n N_VGND_c_828_n 0.00179111f $X=3.9 $Y=1.29 $X2=0 $Y2=0
cc_345 N_C1_M1020_g N_VGND_c_836_n 0.00421418f $X=3.41 $Y=0.79 $X2=0 $Y2=0
cc_346 N_C1_c_402_n N_VGND_c_837_n 0.00452791f $X=3.9 $Y=1.29 $X2=0 $Y2=0
cc_347 N_C1_M1020_g N_VGND_c_838_n 0.00432128f $X=3.41 $Y=0.79 $X2=0 $Y2=0
cc_348 N_C1_c_402_n N_VGND_c_838_n 0.00493565f $X=3.9 $Y=1.29 $X2=0 $Y2=0
cc_349 A1 N_A2_M1004_g 0.00539784f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_350 N_A1_c_460_n N_A2_M1004_g 0.0156388f $X=6.105 $Y=1.615 $X2=0 $Y2=0
cc_351 A1 N_A2_c_509_n 0.013926f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_352 N_A1_c_460_n N_A2_c_509_n 0.00197579f $X=6.105 $Y=1.615 $X2=0 $Y2=0
cc_353 N_A1_M1002_g N_A2_c_512_n 0.00985192f $X=5.675 $Y=0.935 $X2=0 $Y2=0
cc_354 N_A1_M1017_g N_A2_c_512_n 0.00985192f $X=6.105 $Y=0.935 $X2=0 $Y2=0
cc_355 N_A1_M1017_g N_A2_c_513_n 0.011445f $X=6.105 $Y=0.935 $X2=0 $Y2=0
cc_356 A1 N_A2_c_513_n 0.00183891f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_357 N_A1_M1022_g N_A2_M1014_g 0.0283223f $X=6.07 $Y=2.46 $X2=0 $Y2=0
cc_358 N_A1_c_460_n N_A2_M1014_g 0.011445f $X=6.105 $Y=1.615 $X2=0 $Y2=0
cc_359 N_A1_M1017_g N_A2_M1023_g 0.0119526f $X=6.105 $Y=0.935 $X2=0 $Y2=0
cc_360 N_A1_M1002_g N_A2_c_517_n 0.0302298f $X=5.675 $Y=0.935 $X2=0 $Y2=0
cc_361 N_A1_M1003_g N_VPWR_c_579_n 0.0117231f $X=5.62 $Y=2.46 $X2=0 $Y2=0
cc_362 N_A1_M1022_g N_VPWR_c_579_n 4.72395e-19 $X=6.07 $Y=2.46 $X2=0 $Y2=0
cc_363 N_A1_M1003_g N_VPWR_c_580_n 5.11214e-19 $X=5.62 $Y=2.46 $X2=0 $Y2=0
cc_364 N_A1_M1022_g N_VPWR_c_580_n 0.0128567f $X=6.07 $Y=2.46 $X2=0 $Y2=0
cc_365 N_A1_M1003_g N_VPWR_c_581_n 0.00475445f $X=5.62 $Y=2.46 $X2=0 $Y2=0
cc_366 N_A1_M1022_g N_VPWR_c_581_n 0.00460063f $X=6.07 $Y=2.46 $X2=0 $Y2=0
cc_367 N_A1_M1003_g N_VPWR_c_572_n 0.00938661f $X=5.62 $Y=2.46 $X2=0 $Y2=0
cc_368 N_A1_M1022_g N_VPWR_c_572_n 0.00908554f $X=6.07 $Y=2.46 $X2=0 $Y2=0
cc_369 N_A1_M1003_g N_A_517_392#_c_768_n 0.015087f $X=5.62 $Y=2.46 $X2=0 $Y2=0
cc_370 A1 N_A_517_392#_c_768_n 0.0378571f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_371 N_A1_M1022_g N_A_517_392#_c_738_n 0.0156329f $X=6.07 $Y=2.46 $X2=0 $Y2=0
cc_372 A1 N_A_517_392#_c_738_n 0.0111442f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_373 N_A1_c_460_n N_A_517_392#_c_738_n 8.30124e-19 $X=6.105 $Y=1.615 $X2=0
+ $Y2=0
cc_374 N_A1_M1003_g N_A_517_392#_c_742_n 0.0075793f $X=5.62 $Y=2.46 $X2=0 $Y2=0
cc_375 A1 N_A_517_392#_c_742_n 0.0230754f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_376 N_A1_c_460_n N_A_517_392#_c_742_n 0.00225438f $X=6.105 $Y=1.615 $X2=0
+ $Y2=0
cc_377 N_A1_M1017_g N_VGND_c_829_n 5.60436e-19 $X=6.105 $Y=0.935 $X2=0 $Y2=0
cc_378 N_A1_M1002_g N_VGND_c_838_n 9.15321e-19 $X=5.675 $Y=0.935 $X2=0 $Y2=0
cc_379 N_A1_M1017_g N_VGND_c_838_n 9.15321e-19 $X=6.105 $Y=0.935 $X2=0 $Y2=0
cc_380 N_A1_M1002_g N_A_1064_123#_c_927_n 0.00929401f $X=5.675 $Y=0.935 $X2=0
+ $Y2=0
cc_381 N_A1_M1017_g N_A_1064_123#_c_927_n 0.0116895f $X=6.105 $Y=0.935 $X2=0
+ $Y2=0
cc_382 A1 N_A_1064_123#_c_927_n 0.00154834f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_383 N_A1_M1017_g N_A_1064_123#_c_924_n 4.59247e-19 $X=6.105 $Y=0.935 $X2=0
+ $Y2=0
cc_384 N_A2_M1004_g N_VPWR_c_579_n 0.0118013f $X=4.815 $Y=2.46 $X2=0 $Y2=0
cc_385 N_A2_M1014_g N_VPWR_c_580_n 0.0158957f $X=6.52 $Y=2.46 $X2=0 $Y2=0
cc_386 N_A2_M1004_g N_VPWR_c_583_n 0.00475445f $X=4.815 $Y=2.46 $X2=0 $Y2=0
cc_387 N_A2_M1014_g N_VPWR_c_584_n 0.00460063f $X=6.52 $Y=2.46 $X2=0 $Y2=0
cc_388 N_A2_M1004_g N_VPWR_c_572_n 0.00938819f $X=4.815 $Y=2.46 $X2=0 $Y2=0
cc_389 N_A2_M1014_g N_VPWR_c_572_n 0.00912769f $X=6.52 $Y=2.46 $X2=0 $Y2=0
cc_390 N_A2_M1004_g N_A_517_392#_c_736_n 2.3305e-19 $X=4.815 $Y=2.46 $X2=0 $Y2=0
cc_391 N_A2_M1004_g N_A_517_392#_c_768_n 0.021249f $X=4.815 $Y=2.46 $X2=0 $Y2=0
cc_392 N_A2_c_509_n N_A_517_392#_c_768_n 0.00138191f $X=5.17 $Y=1.405 $X2=0
+ $Y2=0
cc_393 N_A2_M1014_g N_A_517_392#_c_738_n 0.0164962f $X=6.52 $Y=2.46 $X2=0 $Y2=0
cc_394 N_A2_M1014_g N_A_517_392#_c_739_n 0.00329219f $X=6.52 $Y=2.46 $X2=0 $Y2=0
cc_395 N_A2_M1014_g N_A_517_392#_c_740_n 4.78926e-19 $X=6.52 $Y=2.46 $X2=0 $Y2=0
cc_396 A2 N_VGND_M1013_s 0.00344879f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_397 N_A2_M1000_g N_VGND_c_828_n 0.00390703f $X=5.245 $Y=0.935 $X2=0 $Y2=0
cc_398 A2 N_VGND_c_828_n 0.0343402f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_399 N_A2_c_517_n N_VGND_c_828_n 0.0052481f $X=5.155 $Y=0.2 $X2=0 $Y2=0
cc_400 N_A2_c_512_n N_VGND_c_829_n 0.00811888f $X=6.46 $Y=0.2 $X2=0 $Y2=0
cc_401 N_A2_M1023_g N_VGND_c_829_n 0.026058f $X=6.535 $Y=0.935 $X2=0 $Y2=0
cc_402 A2 N_VGND_c_833_n 0.0257682f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_403 N_A2_c_517_n N_VGND_c_833_n 0.0403962f $X=5.155 $Y=0.2 $X2=0 $Y2=0
cc_404 N_A2_c_512_n N_VGND_c_838_n 0.0406735f $X=6.46 $Y=0.2 $X2=0 $Y2=0
cc_405 A2 N_VGND_c_838_n 0.0135719f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_406 N_A2_c_517_n N_VGND_c_838_n 0.0100036f $X=5.155 $Y=0.2 $X2=0 $Y2=0
cc_407 N_A2_M1000_g N_A_1064_123#_c_927_n 0.00405878f $X=5.245 $Y=0.935 $X2=0
+ $Y2=0
cc_408 N_A2_c_512_n N_A_1064_123#_c_927_n 0.00827463f $X=6.46 $Y=0.2 $X2=0 $Y2=0
cc_409 A2 N_A_1064_123#_c_927_n 0.00164856f $X=4.955 $Y=0.47 $X2=0 $Y2=0
cc_410 N_A2_c_512_n N_A_1064_123#_c_924_n 0.00275881f $X=6.46 $Y=0.2 $X2=0 $Y2=0
cc_411 N_VPWR_c_574_n N_X_c_671_n 0.0350591f $X=0.39 $Y=1.985 $X2=0 $Y2=0
cc_412 N_VPWR_c_575_n N_X_c_671_n 0.0109793f $X=1.125 $Y=3.33 $X2=0 $Y2=0
cc_413 N_VPWR_c_576_n N_X_c_671_n 0.0297232f $X=1.29 $Y=2.225 $X2=0 $Y2=0
cc_414 N_VPWR_c_572_n N_X_c_671_n 0.00901959f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_415 N_VPWR_M1011_s N_X_c_672_n 0.00165831f $X=1.155 $Y=1.84 $X2=0 $Y2=0
cc_416 N_VPWR_c_576_n N_X_c_672_n 0.0148589f $X=1.29 $Y=2.225 $X2=0 $Y2=0
cc_417 N_VPWR_c_578_n N_X_c_672_n 0.00322693f $X=2.19 $Y=1.985 $X2=0 $Y2=0
cc_418 N_VPWR_c_576_n N_X_c_673_n 0.0309857f $X=1.29 $Y=2.225 $X2=0 $Y2=0
cc_419 N_VPWR_c_577_n N_X_c_673_n 0.0144623f $X=2.105 $Y=3.33 $X2=0 $Y2=0
cc_420 N_VPWR_c_578_n N_X_c_673_n 0.0365151f $X=2.19 $Y=1.985 $X2=0 $Y2=0
cc_421 N_VPWR_c_572_n N_X_c_673_n 0.0118344f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_422 N_VPWR_c_574_n N_X_c_698_n 0.00326551f $X=0.39 $Y=1.985 $X2=0 $Y2=0
cc_423 N_VPWR_c_583_n N_A_517_392#_c_746_n 0.00348696f $X=4.88 $Y=3.33 $X2=0
+ $Y2=0
cc_424 N_VPWR_c_572_n N_A_517_392#_c_746_n 0.00804858f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_425 N_VPWR_c_579_n N_A_517_392#_c_736_n 0.0187075f $X=5.39 $Y=2.485 $X2=0
+ $Y2=0
cc_426 N_VPWR_c_583_n N_A_517_392#_c_736_n 0.00966867f $X=4.88 $Y=3.33 $X2=0
+ $Y2=0
cc_427 N_VPWR_c_572_n N_A_517_392#_c_736_n 0.007728f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_428 N_VPWR_M1004_s N_A_517_392#_c_768_n 0.0142317f $X=4.905 $Y=1.96 $X2=0
+ $Y2=0
cc_429 N_VPWR_c_579_n N_A_517_392#_c_768_n 0.0451464f $X=5.39 $Y=2.485 $X2=0
+ $Y2=0
cc_430 N_VPWR_c_579_n N_A_517_392#_c_737_n 0.0250291f $X=5.39 $Y=2.485 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_580_n N_A_517_392#_c_737_n 0.0266413f $X=6.295 $Y=2.375 $X2=0
+ $Y2=0
cc_432 N_VPWR_c_581_n N_A_517_392#_c_737_n 0.0103967f $X=6.13 $Y=3.33 $X2=0
+ $Y2=0
cc_433 N_VPWR_c_572_n N_A_517_392#_c_737_n 0.00860547f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_434 N_VPWR_M1022_d N_A_517_392#_c_738_n 0.00165831f $X=6.16 $Y=1.96 $X2=0
+ $Y2=0
cc_435 N_VPWR_c_580_n N_A_517_392#_c_738_n 0.0170259f $X=6.295 $Y=2.375 $X2=0
+ $Y2=0
cc_436 N_VPWR_c_580_n N_A_517_392#_c_740_n 0.0266615f $X=6.295 $Y=2.375 $X2=0
+ $Y2=0
cc_437 N_VPWR_c_584_n N_A_517_392#_c_740_n 0.0124046f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_438 N_VPWR_c_572_n N_A_517_392#_c_740_n 0.0102675f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_439 N_VPWR_c_578_n N_A_517_392#_c_741_n 0.021287f $X=2.19 $Y=1.985 $X2=0
+ $Y2=0
cc_440 N_VPWR_c_583_n N_A_517_392#_c_741_n 0.00679992f $X=4.88 $Y=3.33 $X2=0
+ $Y2=0
cc_441 N_VPWR_c_572_n N_A_517_392#_c_741_n 0.0101853f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_442 N_VPWR_c_583_n N_A_517_392#_c_762_n 7.51867e-19 $X=4.88 $Y=3.33 $X2=0
+ $Y2=0
cc_443 N_VPWR_c_572_n N_A_517_392#_c_762_n 0.0020158f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_444 N_VPWR_c_583_n N_A_605_392#_c_809_n 0.0530792f $X=4.88 $Y=3.33 $X2=0
+ $Y2=0
cc_445 N_VPWR_c_572_n N_A_605_392#_c_809_n 0.0433069f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_446 N_X_c_695_n N_VGND_M1007_s 0.00386728f $X=2.18 $Y=0.875 $X2=0 $Y2=0
cc_447 X N_VGND_M1007_s 3.57684e-19 $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_448 N_X_c_669_n N_VGND_M1007_s 0.00197831f $X=1.415 $Y=0.965 $X2=0 $Y2=0
cc_449 N_X_c_666_n N_VGND_c_823_n 0.0144939f $X=1.33 $Y=1.325 $X2=0 $Y2=0
cc_450 N_X_c_667_n N_VGND_c_823_n 0.00888458f $X=0.925 $Y=1.325 $X2=0 $Y2=0
cc_451 N_X_c_668_n N_VGND_c_823_n 0.0164567f $X=1.415 $Y=0.515 $X2=0 $Y2=0
cc_452 N_X_c_668_n N_VGND_c_824_n 0.00749631f $X=1.415 $Y=0.515 $X2=0 $Y2=0
cc_453 N_X_c_668_n N_VGND_c_825_n 0.0103637f $X=1.415 $Y=0.515 $X2=0 $Y2=0
cc_454 N_X_c_695_n N_VGND_c_825_n 0.0122752f $X=2.18 $Y=0.875 $X2=0 $Y2=0
cc_455 X N_VGND_c_825_n 0.00479967f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_456 N_X_c_699_n N_VGND_c_835_n 0.00408057f $X=2.275 $Y=0.745 $X2=0 $Y2=0
cc_457 N_X_c_668_n N_VGND_c_838_n 0.0062048f $X=1.415 $Y=0.515 $X2=0 $Y2=0
cc_458 N_X_c_695_n N_VGND_c_838_n 0.00594702f $X=2.18 $Y=0.875 $X2=0 $Y2=0
cc_459 N_X_c_699_n N_VGND_c_838_n 0.00596517f $X=2.275 $Y=0.745 $X2=0 $Y2=0
cc_460 X N_VGND_c_838_n 0.00681138f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_461 N_A_517_392#_c_746_n N_A_605_392#_M1010_d 0.00431381f $X=4.42 $Y=2.485
+ $X2=-0.19 $Y2=1.66
cc_462 N_A_517_392#_c_746_n N_A_605_392#_M1012_s 0.00422231f $X=4.42 $Y=2.485
+ $X2=0 $Y2=0
cc_463 N_A_517_392#_c_746_n N_A_605_392#_c_809_n 0.0655384f $X=4.42 $Y=2.485
+ $X2=0 $Y2=0
cc_464 N_A_517_392#_c_736_n N_A_605_392#_c_809_n 0.0101394f $X=4.585 $Y=2.825
+ $X2=0 $Y2=0
cc_465 N_A_517_392#_c_739_n N_VGND_c_829_n 0.0113f $X=6.77 $Y=2.12 $X2=0 $Y2=0
cc_466 N_A_517_392#_c_738_n N_A_1064_123#_c_925_n 0.00539705f $X=6.58 $Y=2.035
+ $X2=0 $Y2=0
cc_467 N_VGND_c_828_n N_A_1064_123#_c_927_n 0.00559098f $X=4.59 $Y=0.765 $X2=0
+ $Y2=0
cc_468 N_VGND_c_833_n N_A_1064_123#_c_927_n 0.0122684f $X=6.585 $Y=0 $X2=0 $Y2=0
cc_469 N_VGND_c_838_n N_A_1064_123#_c_927_n 0.0214259f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_470 N_VGND_c_829_n N_A_1064_123#_c_924_n 0.0096909f $X=6.75 $Y=0.76 $X2=0
+ $Y2=0
cc_471 N_VGND_c_833_n N_A_1064_123#_c_924_n 0.00374365f $X=6.585 $Y=0 $X2=0
+ $Y2=0
cc_472 N_VGND_c_838_n N_A_1064_123#_c_924_n 0.00464028f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_473 N_VGND_c_829_n N_A_1064_123#_c_925_n 0.0160983f $X=6.75 $Y=0.76 $X2=0
+ $Y2=0

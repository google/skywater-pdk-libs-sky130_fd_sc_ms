* File: sky130_fd_sc_ms__ha_4.pxi.spice
* Created: Fri Aug 28 17:37:31 2020
* 
x_PM_SKY130_FD_SC_MS__HA_4%A_435_99# N_A_435_99#_M1000_d N_A_435_99#_M1008_d
+ N_A_435_99#_M1029_d N_A_435_99#_c_196_n N_A_435_99#_M1023_g
+ N_A_435_99#_c_197_n N_A_435_99#_c_198_n N_A_435_99#_c_199_n
+ N_A_435_99#_M1028_g N_A_435_99#_M1001_g N_A_435_99#_M1006_g
+ N_A_435_99#_M1009_g N_A_435_99#_M1010_g N_A_435_99#_M1014_g
+ N_A_435_99#_M1012_g N_A_435_99#_M1018_g N_A_435_99#_M1032_g
+ N_A_435_99#_M1020_g N_A_435_99#_M1033_g N_A_435_99#_c_208_n
+ N_A_435_99#_c_209_n N_A_435_99#_c_237_p N_A_435_99#_c_220_n
+ N_A_435_99#_c_221_n N_A_435_99#_c_222_n N_A_435_99#_c_210_n
+ N_A_435_99#_c_285_p N_A_435_99#_c_223_n N_A_435_99#_c_224_n
+ N_A_435_99#_c_211_n PM_SKY130_FD_SC_MS__HA_4%A_435_99#
x_PM_SKY130_FD_SC_MS__HA_4%B N_B_M1002_g N_B_c_392_n N_B_M1019_g N_B_M1007_g
+ N_B_c_393_n N_B_M1021_g N_B_c_394_n N_B_c_386_n N_B_c_396_n N_B_c_397_n
+ N_B_c_398_n N_B_M1008_g N_B_M1000_g N_B_c_400_n N_B_c_388_n N_B_M1003_g
+ N_B_M1025_g N_B_c_390_n N_B_c_404_n B B PM_SKY130_FD_SC_MS__HA_4%B
x_PM_SKY130_FD_SC_MS__HA_4%A N_A_M1016_g N_A_M1013_g N_A_M1022_g N_A_c_521_n
+ N_A_M1017_g N_A_c_509_n N_A_c_510_n N_A_M1029_g N_A_M1004_g N_A_c_513_n
+ N_A_c_514_n N_A_M1011_g N_A_M1034_g N_A_c_516_n N_A_c_517_n A A A N_A_c_519_n
+ PM_SKY130_FD_SC_MS__HA_4%A
x_PM_SKY130_FD_SC_MS__HA_4%A_297_392# N_A_297_392#_M1023_d N_A_297_392#_M1019_d
+ N_A_297_392#_M1001_d N_A_297_392#_M1024_g N_A_297_392#_M1005_g
+ N_A_297_392#_M1027_g N_A_297_392#_M1015_g N_A_297_392#_M1031_g
+ N_A_297_392#_M1026_g N_A_297_392#_c_626_n N_A_297_392#_c_627_n
+ N_A_297_392#_M1030_g N_A_297_392#_M1035_g N_A_297_392#_c_639_n
+ N_A_297_392#_c_630_n N_A_297_392#_c_631_n N_A_297_392#_c_656_n
+ N_A_297_392#_c_658_n N_A_297_392#_c_660_n N_A_297_392#_c_641_n
+ N_A_297_392#_c_632_n N_A_297_392#_c_757_p N_A_297_392#_c_633_n
+ N_A_297_392#_c_642_n N_A_297_392#_c_634_n N_A_297_392#_c_643_n
+ N_A_297_392#_c_676_n N_A_297_392#_c_680_n PM_SKY130_FD_SC_MS__HA_4%A_297_392#
x_PM_SKY130_FD_SC_MS__HA_4%A_27_392# N_A_27_392#_M1016_s N_A_27_392#_M1017_s
+ N_A_27_392#_M1021_s N_A_27_392#_c_820_n N_A_27_392#_c_821_n
+ N_A_27_392#_c_822_n N_A_27_392#_c_823_n N_A_27_392#_c_840_n
+ N_A_27_392#_c_824_n N_A_27_392#_c_825_n N_A_27_392#_c_826_n
+ PM_SKY130_FD_SC_MS__HA_4%A_27_392#
x_PM_SKY130_FD_SC_MS__HA_4%VPWR N_VPWR_M1016_d N_VPWR_M1001_s N_VPWR_M1006_s
+ N_VPWR_M1025_s N_VPWR_M1034_s N_VPWR_M1014_s N_VPWR_M1020_s N_VPWR_M1027_s
+ N_VPWR_M1035_s N_VPWR_c_862_n N_VPWR_c_863_n N_VPWR_c_864_n N_VPWR_c_865_n
+ N_VPWR_c_866_n N_VPWR_c_867_n N_VPWR_c_868_n N_VPWR_c_869_n N_VPWR_c_870_n
+ N_VPWR_c_871_n N_VPWR_c_872_n N_VPWR_c_873_n N_VPWR_c_874_n N_VPWR_c_875_n
+ N_VPWR_c_876_n N_VPWR_c_877_n N_VPWR_c_878_n VPWR N_VPWR_c_879_n
+ N_VPWR_c_880_n N_VPWR_c_881_n N_VPWR_c_882_n N_VPWR_c_883_n N_VPWR_c_884_n
+ N_VPWR_c_885_n N_VPWR_c_886_n N_VPWR_c_887_n N_VPWR_c_888_n N_VPWR_c_861_n
+ PM_SKY130_FD_SC_MS__HA_4%VPWR
x_PM_SKY130_FD_SC_MS__HA_4%COUT N_COUT_M1010_s N_COUT_M1032_s N_COUT_M1009_d
+ N_COUT_M1018_d N_COUT_c_1015_n N_COUT_c_1012_n N_COUT_c_1013_n N_COUT_c_1014_n
+ N_COUT_c_1032_n COUT COUT COUT N_COUT_c_1041_n PM_SKY130_FD_SC_MS__HA_4%COUT
x_PM_SKY130_FD_SC_MS__HA_4%SUM N_SUM_M1005_s N_SUM_M1026_s N_SUM_M1024_d
+ N_SUM_M1031_d N_SUM_c_1070_n N_SUM_c_1071_n N_SUM_c_1063_n N_SUM_c_1064_n
+ N_SUM_c_1065_n N_SUM_c_1066_n N_SUM_c_1072_n N_SUM_c_1067_n N_SUM_c_1073_n
+ N_SUM_c_1068_n N_SUM_c_1069_n N_SUM_c_1075_n N_SUM_c_1076_n N_SUM_c_1117_n
+ N_SUM_c_1118_n SUM PM_SKY130_FD_SC_MS__HA_4%SUM
x_PM_SKY130_FD_SC_MS__HA_4%A_27_125# N_A_27_125#_M1013_d N_A_27_125#_M1022_d
+ N_A_27_125#_M1007_s N_A_27_125#_M1028_s N_A_27_125#_c_1152_n
+ N_A_27_125#_c_1153_n N_A_27_125#_c_1154_n N_A_27_125#_c_1155_n
+ N_A_27_125#_c_1156_n N_A_27_125#_c_1157_n N_A_27_125#_c_1158_n
+ N_A_27_125#_c_1159_n N_A_27_125#_c_1160_n N_A_27_125#_c_1161_n
+ PM_SKY130_FD_SC_MS__HA_4%A_27_125#
x_PM_SKY130_FD_SC_MS__HA_4%VGND N_VGND_M1013_s N_VGND_M1002_d N_VGND_M1004_d
+ N_VGND_M1010_d N_VGND_M1012_d N_VGND_M1033_d N_VGND_M1015_d N_VGND_M1030_d
+ N_VGND_c_1218_n N_VGND_c_1219_n N_VGND_c_1220_n N_VGND_c_1221_n
+ N_VGND_c_1222_n N_VGND_c_1223_n N_VGND_c_1224_n N_VGND_c_1225_n
+ N_VGND_c_1226_n N_VGND_c_1227_n N_VGND_c_1228_n N_VGND_c_1229_n
+ N_VGND_c_1230_n N_VGND_c_1231_n N_VGND_c_1232_n N_VGND_c_1233_n
+ N_VGND_c_1234_n N_VGND_c_1235_n VGND N_VGND_c_1236_n N_VGND_c_1237_n
+ N_VGND_c_1238_n N_VGND_c_1239_n N_VGND_c_1240_n N_VGND_c_1241_n
+ N_VGND_c_1242_n PM_SKY130_FD_SC_MS__HA_4%VGND
x_PM_SKY130_FD_SC_MS__HA_4%A_707_119# N_A_707_119#_M1000_s N_A_707_119#_M1003_s
+ N_A_707_119#_M1011_s N_A_707_119#_c_1344_n N_A_707_119#_c_1345_n
+ N_A_707_119#_c_1346_n N_A_707_119#_c_1347_n N_A_707_119#_c_1348_n
+ N_A_707_119#_c_1349_n N_A_707_119#_c_1350_n
+ PM_SKY130_FD_SC_MS__HA_4%A_707_119#
cc_1 VNB N_A_435_99#_c_196_n 0.0138943f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=1.34
cc_2 VNB N_A_435_99#_c_197_n 0.0163286f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.415
cc_3 VNB N_A_435_99#_c_198_n 0.00729893f $X=-0.19 $Y=-0.245 $X2=2.325 $Y2=1.415
cc_4 VNB N_A_435_99#_c_199_n 0.0156514f $X=-0.19 $Y=-0.245 $X2=2.72 $Y2=1.34
cc_5 VNB N_A_435_99#_M1009_g 5.57468e-19 $X=-0.19 $Y=-0.245 $X2=6.005 $Y2=2.4
cc_6 VNB N_A_435_99#_M1010_g 0.0248403f $X=-0.19 $Y=-0.245 $X2=6.3 $Y2=0.74
cc_7 VNB N_A_435_99#_M1014_g 5.31583e-19 $X=-0.19 $Y=-0.245 $X2=6.615 $Y2=2.4
cc_8 VNB N_A_435_99#_M1012_g 0.0213542f $X=-0.19 $Y=-0.245 $X2=6.73 $Y2=0.74
cc_9 VNB N_A_435_99#_M1018_g 4.76223e-19 $X=-0.19 $Y=-0.245 $X2=7.065 $Y2=2.4
cc_10 VNB N_A_435_99#_M1032_g 0.0205795f $X=-0.19 $Y=-0.245 $X2=7.16 $Y2=0.74
cc_11 VNB N_A_435_99#_M1020_g 4.55039e-19 $X=-0.19 $Y=-0.245 $X2=7.515 $Y2=2.4
cc_12 VNB N_A_435_99#_M1033_g 0.0210466f $X=-0.19 $Y=-0.245 $X2=7.59 $Y2=0.74
cc_13 VNB N_A_435_99#_c_208_n 0.00843023f $X=-0.19 $Y=-0.245 $X2=3.9 $Y2=1.57
cc_14 VNB N_A_435_99#_c_209_n 0.0609931f $X=-0.19 $Y=-0.245 $X2=3.24 $Y2=1.57
cc_15 VNB N_A_435_99#_c_210_n 0.00567831f $X=-0.19 $Y=-0.245 $X2=6.05 $Y2=1.485
cc_16 VNB N_A_435_99#_c_211_n 0.105428f $X=-0.19 $Y=-0.245 $X2=7.515 $Y2=1.485
cc_17 VNB N_B_M1002_g 0.0185323f $X=-0.19 $Y=-0.245 $X2=4.91 $Y2=2.05
cc_18 VNB N_B_M1007_g 0.0186662f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=1.34
cc_19 VNB N_B_c_386_n 0.0269801f $X=-0.19 $Y=-0.245 $X2=2.72 $Y2=0.945
cc_20 VNB N_B_M1000_g 0.025966f $X=-0.19 $Y=-0.245 $X2=6.005 $Y2=2.4
cc_21 VNB N_B_c_388_n 0.00653496f $X=-0.19 $Y=-0.245 $X2=6.3 $Y2=0.74
cc_22 VNB N_B_M1003_g 0.0231254f $X=-0.19 $Y=-0.245 $X2=6.615 $Y2=2.4
cc_23 VNB N_B_c_390_n 0.00674071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB B 0.0037323f $X=-0.19 $Y=-0.245 $X2=7.065 $Y2=2.4
cc_25 VNB N_A_M1013_g 0.0287386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_M1022_g 0.0316014f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=0.945
cc_27 VNB N_A_c_509_n 0.283484f $X=-0.19 $Y=-0.245 $X2=2.72 $Y2=0.945
cc_28 VNB N_A_c_510_n 0.0125033f $X=-0.19 $Y=-0.245 $X2=2.72 $Y2=0.945
cc_29 VNB N_A_M1029_g 9.04456e-19 $X=-0.19 $Y=-0.245 $X2=2.865 $Y2=2.315
cc_30 VNB N_A_M1004_g 0.0253437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_c_513_n 0.0195879f $X=-0.19 $Y=-0.245 $X2=6.005 $Y2=1.65
cc_32 VNB N_A_c_514_n 0.0163093f $X=-0.19 $Y=-0.245 $X2=6.005 $Y2=2.4
cc_33 VNB N_A_M1034_g 0.00188321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_c_516_n 0.0103239f $X=-0.19 $Y=-0.245 $X2=6.615 $Y2=2.4
cc_35 VNB N_A_c_517_n 0.0139766f $X=-0.19 $Y=-0.245 $X2=6.615 $Y2=2.4
cc_36 VNB A 0.0142582f $X=-0.19 $Y=-0.245 $X2=6.73 $Y2=0.74
cc_37 VNB N_A_c_519_n 0.0245972f $X=-0.19 $Y=-0.245 $X2=7.16 $Y2=0.74
cc_38 VNB N_A_297_392#_M1024_g 4.41828e-19 $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=0.945
cc_39 VNB N_A_297_392#_M1005_g 0.0219202f $X=-0.19 $Y=-0.245 $X2=2.72 $Y2=0.945
cc_40 VNB N_A_297_392#_M1027_g 4.78354e-19 $X=-0.19 $Y=-0.245 $X2=2.865
+ $Y2=2.315
cc_41 VNB N_A_297_392#_M1015_g 0.0226903f $X=-0.19 $Y=-0.245 $X2=3.315 $Y2=2.315
cc_42 VNB N_A_297_392#_M1031_g 5.61811e-19 $X=-0.19 $Y=-0.245 $X2=6.005 $Y2=2.4
cc_43 VNB N_A_297_392#_M1026_g 0.0237211f $X=-0.19 $Y=-0.245 $X2=6.3 $Y2=0.74
cc_44 VNB N_A_297_392#_c_626_n 0.0282531f $X=-0.19 $Y=-0.245 $X2=6.615 $Y2=1.65
cc_45 VNB N_A_297_392#_c_627_n 0.0577641f $X=-0.19 $Y=-0.245 $X2=6.615 $Y2=2.4
cc_46 VNB N_A_297_392#_M1030_g 0.0256152f $X=-0.19 $Y=-0.245 $X2=6.73 $Y2=1.32
cc_47 VNB N_A_297_392#_M1035_g 6.11644e-19 $X=-0.19 $Y=-0.245 $X2=7.065 $Y2=1.65
cc_48 VNB N_A_297_392#_c_630_n 0.00202173f $X=-0.19 $Y=-0.245 $X2=7.515 $Y2=1.65
cc_49 VNB N_A_297_392#_c_631_n 0.00324153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_297_392#_c_632_n 0.00477785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_297_392#_c_633_n 0.0237824f $X=-0.19 $Y=-0.245 $X2=4.23 $Y2=1.907
cc_52 VNB N_A_297_392#_c_634_n 0.00162343f $X=-0.19 $Y=-0.245 $X2=5.12 $Y2=1.985
cc_53 VNB N_VPWR_c_861_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_COUT_c_1012_n 0.00186123f $X=-0.19 $Y=-0.245 $X2=2.72 $Y2=0.945
cc_55 VNB N_COUT_c_1013_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=2.865 $Y2=2.315
cc_56 VNB N_COUT_c_1014_n 0.00541261f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_SUM_c_1063_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=2.865 $Y2=2.315
cc_58 VNB N_SUM_c_1064_n 0.00307912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_SUM_c_1065_n 0.00220472f $X=-0.19 $Y=-0.245 $X2=3.315 $Y2=1.735
cc_60 VNB N_SUM_c_1066_n 0.00327315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_SUM_c_1067_n 0.0154148f $X=-0.19 $Y=-0.245 $X2=6.3 $Y2=0.74
cc_62 VNB N_SUM_c_1068_n 0.0243971f $X=-0.19 $Y=-0.245 $X2=6.615 $Y2=2.4
cc_63 VNB N_SUM_c_1069_n 0.00241905f $X=-0.19 $Y=-0.245 $X2=6.73 $Y2=0.74
cc_64 VNB N_A_27_125#_c_1152_n 0.0221323f $X=-0.19 $Y=-0.245 $X2=2.72 $Y2=1.34
cc_65 VNB N_A_27_125#_c_1153_n 0.0027328f $X=-0.19 $Y=-0.245 $X2=2.72 $Y2=0.945
cc_66 VNB N_A_27_125#_c_1154_n 0.00952244f $X=-0.19 $Y=-0.245 $X2=2.865
+ $Y2=1.735
cc_67 VNB N_A_27_125#_c_1155_n 0.00244123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_27_125#_c_1156_n 0.00620491f $X=-0.19 $Y=-0.245 $X2=3.315
+ $Y2=2.315
cc_69 VNB N_A_27_125#_c_1157_n 0.00337282f $X=-0.19 $Y=-0.245 $X2=6.005 $Y2=2.4
cc_70 VNB N_A_27_125#_c_1158_n 0.0216937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_27_125#_c_1159_n 0.00432301f $X=-0.19 $Y=-0.245 $X2=6.3 $Y2=1.32
cc_72 VNB N_A_27_125#_c_1160_n 0.0134046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_27_125#_c_1161_n 0.00204143f $X=-0.19 $Y=-0.245 $X2=6.615 $Y2=2.4
cc_74 VNB N_VGND_c_1218_n 0.0181522f $X=-0.19 $Y=-0.245 $X2=6.005 $Y2=2.4
cc_75 VNB N_VGND_c_1219_n 0.00638216f $X=-0.19 $Y=-0.245 $X2=6.3 $Y2=0.74
cc_76 VNB N_VGND_c_1220_n 0.0151544f $X=-0.19 $Y=-0.245 $X2=6.615 $Y2=2.4
cc_77 VNB N_VGND_c_1221_n 0.0190588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1222_n 0.0178645f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1223_n 0.0026136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1224_n 0.002601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1225_n 0.00558127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1226_n 0.0142878f $X=-0.19 $Y=-0.245 $X2=7.59 $Y2=0.74
cc_83 VNB N_VGND_c_1227_n 0.029743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1228_n 0.0183144f $X=-0.19 $Y=-0.245 $X2=3.24 $Y2=1.57
cc_85 VNB N_VGND_c_1229_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=3.24 $Y2=1.57
cc_86 VNB N_VGND_c_1230_n 0.0172883f $X=-0.19 $Y=-0.245 $X2=4.115 $Y2=1.405
cc_87 VNB N_VGND_c_1231_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=4.115 $Y2=0.74
cc_88 VNB N_VGND_c_1232_n 0.016486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1233_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=4.955 $Y2=1.907
cc_90 VNB N_VGND_c_1234_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=5.88 $Y2=1.985
cc_91 VNB N_VGND_c_1235_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=5.12 $Y2=1.985
cc_92 VNB N_VGND_c_1236_n 0.0807918f $X=-0.19 $Y=-0.245 $X2=6.79 $Y2=1.485
cc_93 VNB N_VGND_c_1237_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=4.955 $Y2=1.985
cc_94 VNB N_VGND_c_1238_n 0.018855f $X=-0.19 $Y=-0.245 $X2=7.16 $Y2=1.485
cc_95 VNB N_VGND_c_1239_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1240_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1241_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1242_n 0.527831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_707_119#_c_1344_n 0.0130452f $X=-0.19 $Y=-0.245 $X2=2.25 $Y2=0.945
cc_100 VNB N_A_707_119#_c_1345_n 0.0106798f $X=-0.19 $Y=-0.245 $X2=2.325
+ $Y2=1.415
cc_101 VNB N_A_707_119#_c_1346_n 0.00422464f $X=-0.19 $Y=-0.245 $X2=2.72
+ $Y2=1.34
cc_102 VNB N_A_707_119#_c_1347_n 0.00269685f $X=-0.19 $Y=-0.245 $X2=2.865
+ $Y2=2.315
cc_103 VNB N_A_707_119#_c_1348_n 0.00636128f $X=-0.19 $Y=-0.245 $X2=2.865
+ $Y2=2.315
cc_104 VNB N_A_707_119#_c_1349_n 0.00152462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_707_119#_c_1350_n 0.0140492f $X=-0.19 $Y=-0.245 $X2=3.315
+ $Y2=2.315
cc_106 VPB N_A_435_99#_M1001_g 0.0186976f $X=-0.19 $Y=1.66 $X2=2.865 $Y2=2.315
cc_107 VPB N_A_435_99#_M1006_g 0.0179509f $X=-0.19 $Y=1.66 $X2=3.315 $Y2=2.315
cc_108 VPB N_A_435_99#_M1009_g 0.0261567f $X=-0.19 $Y=1.66 $X2=6.005 $Y2=2.4
cc_109 VPB N_A_435_99#_M1014_g 0.0234176f $X=-0.19 $Y=1.66 $X2=6.615 $Y2=2.4
cc_110 VPB N_A_435_99#_M1018_g 0.0215679f $X=-0.19 $Y=1.66 $X2=7.065 $Y2=2.4
cc_111 VPB N_A_435_99#_M1020_g 0.0213295f $X=-0.19 $Y=1.66 $X2=7.515 $Y2=2.4
cc_112 VPB N_A_435_99#_c_208_n 0.00428654f $X=-0.19 $Y=1.66 $X2=3.9 $Y2=1.57
cc_113 VPB N_A_435_99#_c_209_n 0.0100435f $X=-0.19 $Y=1.66 $X2=3.24 $Y2=1.57
cc_114 VPB N_A_435_99#_c_220_n 0.0104246f $X=-0.19 $Y=1.66 $X2=5.88 $Y2=1.985
cc_115 VPB N_A_435_99#_c_221_n 0.00184703f $X=-0.19 $Y=1.66 $X2=5.12 $Y2=1.985
cc_116 VPB N_A_435_99#_c_222_n 0.00193973f $X=-0.19 $Y=1.66 $X2=5.965 $Y2=1.82
cc_117 VPB N_A_435_99#_c_223_n 0.00404608f $X=-0.19 $Y=1.66 $X2=4.07 $Y2=1.907
cc_118 VPB N_A_435_99#_c_224_n 0.0105359f $X=-0.19 $Y=1.66 $X2=4.955 $Y2=1.985
cc_119 VPB N_B_c_392_n 0.0162877f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_B_c_393_n 0.0166049f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=0.945
cc_121 VPB N_B_c_394_n 0.0254305f $X=-0.19 $Y=1.66 $X2=2.72 $Y2=1.34
cc_122 VPB N_B_c_386_n 0.0225156f $X=-0.19 $Y=1.66 $X2=2.72 $Y2=0.945
cc_123 VPB N_B_c_396_n 0.0661267f $X=-0.19 $Y=1.66 $X2=2.865 $Y2=1.735
cc_124 VPB N_B_c_397_n 0.0891643f $X=-0.19 $Y=1.66 $X2=2.865 $Y2=2.315
cc_125 VPB N_B_c_398_n 0.0123634f $X=-0.19 $Y=1.66 $X2=2.865 $Y2=2.315
cc_126 VPB N_B_M1008_g 0.0303505f $X=-0.19 $Y=1.66 $X2=3.315 $Y2=2.315
cc_127 VPB N_B_c_400_n 0.041437f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_B_c_388_n 0.0157834f $X=-0.19 $Y=1.66 $X2=6.3 $Y2=0.74
cc_129 VPB N_B_M1025_g 0.0217152f $X=-0.19 $Y=1.66 $X2=6.73 $Y2=0.74
cc_130 VPB N_B_c_390_n 0.00761646f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_B_c_404_n 0.0087959f $X=-0.19 $Y=1.66 $X2=7.065 $Y2=1.65
cc_132 VPB B 5.62692e-19 $X=-0.19 $Y=1.66 $X2=7.065 $Y2=2.4
cc_133 VPB N_A_M1016_g 0.0304622f $X=-0.19 $Y=1.66 $X2=4.91 $Y2=2.05
cc_134 VPB N_A_c_521_n 0.0168597f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=1.415
cc_135 VPB N_A_M1029_g 0.0386086f $X=-0.19 $Y=1.66 $X2=2.865 $Y2=2.315
cc_136 VPB N_A_M1034_g 0.025438f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_c_516_n 0.00127149f $X=-0.19 $Y=1.66 $X2=6.615 $Y2=2.4
cc_138 VPB A 0.0121842f $X=-0.19 $Y=1.66 $X2=6.73 $Y2=0.74
cc_139 VPB N_A_c_519_n 0.0211223f $X=-0.19 $Y=1.66 $X2=7.16 $Y2=0.74
cc_140 VPB N_A_297_392#_M1024_g 0.0210788f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=0.945
cc_141 VPB N_A_297_392#_M1027_g 0.021618f $X=-0.19 $Y=1.66 $X2=2.865 $Y2=2.315
cc_142 VPB N_A_297_392#_M1031_g 0.024432f $X=-0.19 $Y=1.66 $X2=6.005 $Y2=2.4
cc_143 VPB N_A_297_392#_M1035_g 0.0276169f $X=-0.19 $Y=1.66 $X2=7.065 $Y2=1.65
cc_144 VPB N_A_297_392#_c_639_n 0.00704073f $X=-0.19 $Y=1.66 $X2=7.16 $Y2=1.32
cc_145 VPB N_A_297_392#_c_631_n 0.00458992f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_297_392#_c_641_n 0.00105386f $X=-0.19 $Y=1.66 $X2=3.24 $Y2=1.57
cc_147 VPB N_A_297_392#_c_642_n 0.00267377f $X=-0.19 $Y=1.66 $X2=5.12 $Y2=1.985
cc_148 VPB N_A_297_392#_c_643_n 5.40493e-19 $X=-0.19 $Y=1.66 $X2=5.965 $Y2=1.65
cc_149 VPB N_A_27_392#_c_820_n 0.0101511f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=1.34
cc_150 VPB N_A_27_392#_c_821_n 0.0340347f $X=-0.19 $Y=1.66 $X2=2.25 $Y2=0.945
cc_151 VPB N_A_27_392#_c_822_n 0.00236883f $X=-0.19 $Y=1.66 $X2=2.325 $Y2=1.415
cc_152 VPB N_A_27_392#_c_823_n 0.00206591f $X=-0.19 $Y=1.66 $X2=2.72 $Y2=0.945
cc_153 VPB N_A_27_392#_c_824_n 0.00614925f $X=-0.19 $Y=1.66 $X2=2.865 $Y2=2.315
cc_154 VPB N_A_27_392#_c_825_n 0.00160153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_27_392#_c_826_n 0.00525438f $X=-0.19 $Y=1.66 $X2=3.315 $Y2=2.315
cc_156 VPB N_VPWR_c_862_n 0.00521506f $X=-0.19 $Y=1.66 $X2=6.3 $Y2=1.32
cc_157 VPB N_VPWR_c_863_n 0.00898781f $X=-0.19 $Y=1.66 $X2=6.615 $Y2=1.65
cc_158 VPB N_VPWR_c_864_n 0.00328505f $X=-0.19 $Y=1.66 $X2=6.73 $Y2=1.32
cc_159 VPB N_VPWR_c_865_n 0.00490739f $X=-0.19 $Y=1.66 $X2=7.065 $Y2=1.65
cc_160 VPB N_VPWR_c_866_n 0.0231664f $X=-0.19 $Y=1.66 $X2=7.065 $Y2=2.4
cc_161 VPB N_VPWR_c_867_n 0.0139016f $X=-0.19 $Y=1.66 $X2=7.16 $Y2=0.74
cc_162 VPB N_VPWR_c_868_n 0.00329129f $X=-0.19 $Y=1.66 $X2=7.515 $Y2=2.4
cc_163 VPB N_VPWR_c_869_n 0.00261791f $X=-0.19 $Y=1.66 $X2=7.59 $Y2=0.74
cc_164 VPB N_VPWR_c_870_n 0.00329129f $X=-0.19 $Y=1.66 $X2=3.24 $Y2=1.57
cc_165 VPB N_VPWR_c_871_n 0.0119967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_872_n 0.0343838f $X=-0.19 $Y=1.66 $X2=4.115 $Y2=0.74
cc_167 VPB N_VPWR_c_873_n 0.0228504f $X=-0.19 $Y=1.66 $X2=4.955 $Y2=1.907
cc_168 VPB N_VPWR_c_874_n 0.00601644f $X=-0.19 $Y=1.66 $X2=4.23 $Y2=1.907
cc_169 VPB N_VPWR_c_875_n 0.0177589f $X=-0.19 $Y=1.66 $X2=5.12 $Y2=1.985
cc_170 VPB N_VPWR_c_876_n 0.00601644f $X=-0.19 $Y=1.66 $X2=5.12 $Y2=1.985
cc_171 VPB N_VPWR_c_877_n 0.0159778f $X=-0.19 $Y=1.66 $X2=5.965 $Y2=1.65
cc_172 VPB N_VPWR_c_878_n 0.00601644f $X=-0.19 $Y=1.66 $X2=5.965 $Y2=1.82
cc_173 VPB N_VPWR_c_879_n 0.0175377f $X=-0.19 $Y=1.66 $X2=6.11 $Y2=1.485
cc_174 VPB N_VPWR_c_880_n 0.0400623f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_881_n 0.0159813f $X=-0.19 $Y=1.66 $X2=3.24 $Y2=1.537
cc_176 VPB N_VPWR_c_882_n 0.0209137f $X=-0.19 $Y=1.66 $X2=6.615 $Y2=1.485
cc_177 VPB N_VPWR_c_883_n 0.0234703f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_884_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_885_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_886_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_887_n 0.00507883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_888_n 0.00853174f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_861_n 0.0920695f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_COUT_c_1015_n 0.0070956f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=1.415
cc_185 VPB COUT 0.00157509f $X=-0.19 $Y=1.66 $X2=6.005 $Y2=2.4
cc_186 VPB N_SUM_c_1070_n 0.00200827f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=1.415
cc_187 VPB N_SUM_c_1071_n 0.00233077f $X=-0.19 $Y=1.66 $X2=2.72 $Y2=1.34
cc_188 VPB N_SUM_c_1072_n 0.00332456f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_SUM_c_1073_n 0.00277699f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_SUM_c_1068_n 0.0226818f $X=-0.19 $Y=1.66 $X2=6.615 $Y2=2.4
cc_191 VPB N_SUM_c_1075_n 0.00338435f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_SUM_c_1076_n 0.0021278f $X=-0.19 $Y=1.66 $X2=7.065 $Y2=2.4
cc_193 VPB SUM 9.18137e-19 $X=-0.19 $Y=1.66 $X2=7.515 $Y2=1.65
cc_194 VPB N_A_707_119#_c_1349_n 0.00302006f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 N_A_435_99#_c_196_n N_B_M1007_g 0.0131498f $X=2.25 $Y=1.34 $X2=0 $Y2=0
cc_196 N_A_435_99#_c_198_n N_B_c_394_n 0.0155847f $X=2.325 $Y=1.415 $X2=0 $Y2=0
cc_197 N_A_435_99#_c_209_n N_B_c_394_n 0.0152784f $X=3.24 $Y=1.57 $X2=0 $Y2=0
cc_198 N_A_435_99#_c_198_n N_B_c_386_n 0.00195768f $X=2.325 $Y=1.415 $X2=0 $Y2=0
cc_199 N_A_435_99#_M1001_g N_B_c_396_n 0.0152784f $X=2.865 $Y=2.315 $X2=0 $Y2=0
cc_200 N_A_435_99#_M1001_g N_B_c_397_n 0.0123711f $X=2.865 $Y=2.315 $X2=0 $Y2=0
cc_201 N_A_435_99#_M1006_g N_B_c_397_n 0.0123711f $X=3.315 $Y=2.315 $X2=0 $Y2=0
cc_202 N_A_435_99#_M1006_g N_B_M1008_g 0.0239592f $X=3.315 $Y=2.315 $X2=0 $Y2=0
cc_203 N_A_435_99#_c_208_n N_B_M1008_g 0.00573983f $X=3.9 $Y=1.57 $X2=0 $Y2=0
cc_204 N_A_435_99#_c_223_n N_B_M1008_g 0.00672473f $X=4.07 $Y=1.907 $X2=0 $Y2=0
cc_205 N_A_435_99#_c_208_n N_B_M1000_g 0.00633468f $X=3.9 $Y=1.57 $X2=0 $Y2=0
cc_206 N_A_435_99#_c_209_n N_B_M1000_g 0.00541031f $X=3.24 $Y=1.57 $X2=0 $Y2=0
cc_207 N_A_435_99#_c_237_p N_B_M1000_g 0.0143629f $X=4.115 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A_435_99#_c_223_n N_B_M1000_g 0.00491066f $X=4.07 $Y=1.907 $X2=0 $Y2=0
cc_209 N_A_435_99#_c_223_n N_B_c_388_n 0.0138324f $X=4.07 $Y=1.907 $X2=0 $Y2=0
cc_210 N_A_435_99#_c_224_n N_B_c_388_n 0.00418849f $X=4.955 $Y=1.985 $X2=0 $Y2=0
cc_211 N_A_435_99#_c_237_p N_B_M1003_g 0.00998427f $X=4.115 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A_435_99#_c_223_n N_B_M1003_g 0.00276031f $X=4.07 $Y=1.907 $X2=0 $Y2=0
cc_213 N_A_435_99#_c_224_n N_B_M1025_g 0.00820544f $X=4.955 $Y=1.985 $X2=0 $Y2=0
cc_214 N_A_435_99#_c_208_n N_B_c_390_n 0.00808718f $X=3.9 $Y=1.57 $X2=0 $Y2=0
cc_215 N_A_435_99#_c_209_n N_B_c_390_n 0.0239592f $X=3.24 $Y=1.57 $X2=0 $Y2=0
cc_216 N_A_435_99#_c_223_n N_B_c_390_n 0.00256558f $X=4.07 $Y=1.907 $X2=0 $Y2=0
cc_217 N_A_435_99#_c_198_n B 0.00706672f $X=2.325 $Y=1.415 $X2=0 $Y2=0
cc_218 N_A_435_99#_c_196_n N_A_c_509_n 0.00737233f $X=2.25 $Y=1.34 $X2=0 $Y2=0
cc_219 N_A_435_99#_c_199_n N_A_c_509_n 0.00737233f $X=2.72 $Y=1.34 $X2=0 $Y2=0
cc_220 N_A_435_99#_c_221_n N_A_M1029_g 0.00232581f $X=5.12 $Y=1.985 $X2=0 $Y2=0
cc_221 N_A_435_99#_c_223_n N_A_M1029_g 0.00238841f $X=4.07 $Y=1.907 $X2=0 $Y2=0
cc_222 N_A_435_99#_c_224_n N_A_M1029_g 0.014982f $X=4.955 $Y=1.985 $X2=0 $Y2=0
cc_223 N_A_435_99#_c_237_p N_A_M1004_g 2.53475e-19 $X=4.115 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A_435_99#_c_221_n N_A_c_513_n 0.00376408f $X=5.12 $Y=1.985 $X2=0 $Y2=0
cc_225 N_A_435_99#_M1009_g N_A_M1034_g 0.0153028f $X=6.005 $Y=2.4 $X2=0 $Y2=0
cc_226 N_A_435_99#_c_220_n N_A_M1034_g 0.0168942f $X=5.88 $Y=1.985 $X2=0 $Y2=0
cc_227 N_A_435_99#_c_222_n N_A_M1034_g 0.00275668f $X=5.965 $Y=1.82 $X2=0 $Y2=0
cc_228 N_A_435_99#_c_223_n N_A_c_516_n 3.08349e-19 $X=4.07 $Y=1.907 $X2=0 $Y2=0
cc_229 N_A_435_99#_c_210_n N_A_c_517_n 0.00182743f $X=6.05 $Y=1.485 $X2=0 $Y2=0
cc_230 N_A_435_99#_c_211_n N_A_c_517_n 0.0183704f $X=7.515 $Y=1.485 $X2=0 $Y2=0
cc_231 N_A_435_99#_M1020_g N_A_297_392#_M1024_g 0.0280389f $X=7.515 $Y=2.4 $X2=0
+ $Y2=0
cc_232 N_A_435_99#_M1033_g N_A_297_392#_M1005_g 0.0317962f $X=7.59 $Y=0.74 $X2=0
+ $Y2=0
cc_233 N_A_435_99#_c_211_n N_A_297_392#_c_627_n 0.037891f $X=7.515 $Y=1.485
+ $X2=0 $Y2=0
cc_234 N_A_435_99#_c_197_n N_A_297_392#_c_639_n 0.00116202f $X=2.645 $Y=1.415
+ $X2=0 $Y2=0
cc_235 N_A_435_99#_c_198_n N_A_297_392#_c_639_n 7.88945e-19 $X=2.325 $Y=1.415
+ $X2=0 $Y2=0
cc_236 N_A_435_99#_c_196_n N_A_297_392#_c_630_n 3.39182e-19 $X=2.25 $Y=1.34
+ $X2=0 $Y2=0
cc_237 N_A_435_99#_c_199_n N_A_297_392#_c_630_n 0.00586917f $X=2.72 $Y=1.34
+ $X2=0 $Y2=0
cc_238 N_A_435_99#_c_196_n N_A_297_392#_c_631_n 0.00113236f $X=2.25 $Y=1.34
+ $X2=0 $Y2=0
cc_239 N_A_435_99#_c_197_n N_A_297_392#_c_631_n 0.00939344f $X=2.645 $Y=1.415
+ $X2=0 $Y2=0
cc_240 N_A_435_99#_c_199_n N_A_297_392#_c_631_n 0.00257225f $X=2.72 $Y=1.34
+ $X2=0 $Y2=0
cc_241 N_A_435_99#_c_208_n N_A_297_392#_c_631_n 0.0132865f $X=3.9 $Y=1.57 $X2=0
+ $Y2=0
cc_242 N_A_435_99#_c_209_n N_A_297_392#_c_631_n 0.0170184f $X=3.24 $Y=1.57 $X2=0
+ $Y2=0
cc_243 N_A_435_99#_M1001_g N_A_297_392#_c_656_n 0.0170496f $X=2.865 $Y=2.315
+ $X2=0 $Y2=0
cc_244 N_A_435_99#_c_209_n N_A_297_392#_c_656_n 0.00262599f $X=3.24 $Y=1.57
+ $X2=0 $Y2=0
cc_245 N_A_435_99#_M1006_g N_A_297_392#_c_658_n 0.0130928f $X=3.315 $Y=2.315
+ $X2=0 $Y2=0
cc_246 N_A_435_99#_c_208_n N_A_297_392#_c_658_n 0.0208597f $X=3.9 $Y=1.57 $X2=0
+ $Y2=0
cc_247 N_A_435_99#_M1008_d N_A_297_392#_c_660_n 0.00439536f $X=3.855 $Y=1.895
+ $X2=0 $Y2=0
cc_248 N_A_435_99#_M1029_d N_A_297_392#_c_660_n 0.00698844f $X=4.91 $Y=2.05
+ $X2=0 $Y2=0
cc_249 N_A_435_99#_M1009_g N_A_297_392#_c_660_n 0.0155313f $X=6.005 $Y=2.4 $X2=0
+ $Y2=0
cc_250 N_A_435_99#_M1014_g N_A_297_392#_c_660_n 0.0139057f $X=6.615 $Y=2.4 $X2=0
+ $Y2=0
cc_251 N_A_435_99#_M1018_g N_A_297_392#_c_660_n 0.0130823f $X=7.065 $Y=2.4 $X2=0
+ $Y2=0
cc_252 N_A_435_99#_M1020_g N_A_297_392#_c_660_n 0.0145517f $X=7.515 $Y=2.4 $X2=0
+ $Y2=0
cc_253 N_A_435_99#_c_220_n N_A_297_392#_c_660_n 0.0102837f $X=5.88 $Y=1.985
+ $X2=0 $Y2=0
cc_254 N_A_435_99#_c_221_n N_A_297_392#_c_660_n 0.0584005f $X=5.12 $Y=1.985
+ $X2=0 $Y2=0
cc_255 N_A_435_99#_c_285_p N_A_297_392#_c_660_n 0.00337845f $X=6.79 $Y=1.485
+ $X2=0 $Y2=0
cc_256 N_A_435_99#_c_223_n N_A_297_392#_c_660_n 0.00733564f $X=4.07 $Y=1.907
+ $X2=0 $Y2=0
cc_257 N_A_435_99#_c_224_n N_A_297_392#_c_660_n 0.0268397f $X=4.955 $Y=1.985
+ $X2=0 $Y2=0
cc_258 N_A_435_99#_c_211_n N_A_297_392#_c_660_n 9.58046e-19 $X=7.515 $Y=1.485
+ $X2=0 $Y2=0
cc_259 N_A_435_99#_M1020_g N_A_297_392#_c_641_n 0.00678981f $X=7.515 $Y=2.4
+ $X2=0 $Y2=0
cc_260 N_A_435_99#_c_211_n N_A_297_392#_c_632_n 0.00279232f $X=7.515 $Y=1.485
+ $X2=0 $Y2=0
cc_261 N_A_435_99#_c_197_n N_A_297_392#_c_634_n 0.00266209f $X=2.645 $Y=1.415
+ $X2=0 $Y2=0
cc_262 N_A_435_99#_c_199_n N_A_297_392#_c_634_n 0.00361003f $X=2.72 $Y=1.34
+ $X2=0 $Y2=0
cc_263 N_A_435_99#_M1001_g N_A_297_392#_c_676_n 0.00782021f $X=2.865 $Y=2.315
+ $X2=0 $Y2=0
cc_264 N_A_435_99#_M1006_g N_A_297_392#_c_676_n 0.0080397f $X=3.315 $Y=2.315
+ $X2=0 $Y2=0
cc_265 N_A_435_99#_c_208_n N_A_297_392#_c_676_n 0.0118089f $X=3.9 $Y=1.57 $X2=0
+ $Y2=0
cc_266 N_A_435_99#_c_209_n N_A_297_392#_c_676_n 0.00230862f $X=3.24 $Y=1.57
+ $X2=0 $Y2=0
cc_267 N_A_435_99#_M1008_d N_A_297_392#_c_680_n 0.00627358f $X=3.855 $Y=1.895
+ $X2=0 $Y2=0
cc_268 N_A_435_99#_c_223_n N_A_297_392#_c_680_n 0.0133856f $X=4.07 $Y=1.907
+ $X2=0 $Y2=0
cc_269 N_A_435_99#_c_220_n N_VPWR_M1034_s 0.00603299f $X=5.88 $Y=1.985 $X2=0
+ $Y2=0
cc_270 N_A_435_99#_M1001_g N_VPWR_c_863_n 0.01114f $X=2.865 $Y=2.315 $X2=0 $Y2=0
cc_271 N_A_435_99#_M1006_g N_VPWR_c_863_n 0.00152804f $X=3.315 $Y=2.315 $X2=0
+ $Y2=0
cc_272 N_A_435_99#_M1001_g N_VPWR_c_864_n 0.00105204f $X=2.865 $Y=2.315 $X2=0
+ $Y2=0
cc_273 N_A_435_99#_M1006_g N_VPWR_c_864_n 0.00904323f $X=3.315 $Y=2.315 $X2=0
+ $Y2=0
cc_274 N_A_435_99#_M1009_g N_VPWR_c_867_n 0.0190935f $X=6.005 $Y=2.4 $X2=0 $Y2=0
cc_275 N_A_435_99#_M1014_g N_VPWR_c_867_n 0.00191874f $X=6.615 $Y=2.4 $X2=0
+ $Y2=0
cc_276 N_A_435_99#_M1009_g N_VPWR_c_868_n 0.00192487f $X=6.005 $Y=2.4 $X2=0
+ $Y2=0
cc_277 N_A_435_99#_M1014_g N_VPWR_c_868_n 0.0117561f $X=6.615 $Y=2.4 $X2=0 $Y2=0
cc_278 N_A_435_99#_M1018_g N_VPWR_c_868_n 0.0107196f $X=7.065 $Y=2.4 $X2=0 $Y2=0
cc_279 N_A_435_99#_M1020_g N_VPWR_c_868_n 0.00125818f $X=7.515 $Y=2.4 $X2=0
+ $Y2=0
cc_280 N_A_435_99#_M1018_g N_VPWR_c_869_n 0.00125818f $X=7.065 $Y=2.4 $X2=0
+ $Y2=0
cc_281 N_A_435_99#_M1020_g N_VPWR_c_869_n 0.0106899f $X=7.515 $Y=2.4 $X2=0 $Y2=0
cc_282 N_A_435_99#_M1009_g N_VPWR_c_873_n 0.00460063f $X=6.005 $Y=2.4 $X2=0
+ $Y2=0
cc_283 N_A_435_99#_M1014_g N_VPWR_c_873_n 0.00460063f $X=6.615 $Y=2.4 $X2=0
+ $Y2=0
cc_284 N_A_435_99#_M1018_g N_VPWR_c_875_n 0.00460063f $X=7.065 $Y=2.4 $X2=0
+ $Y2=0
cc_285 N_A_435_99#_M1020_g N_VPWR_c_875_n 0.00460063f $X=7.515 $Y=2.4 $X2=0
+ $Y2=0
cc_286 N_A_435_99#_M1001_g N_VPWR_c_861_n 9.455e-19 $X=2.865 $Y=2.315 $X2=0
+ $Y2=0
cc_287 N_A_435_99#_M1006_g N_VPWR_c_861_n 9.455e-19 $X=3.315 $Y=2.315 $X2=0
+ $Y2=0
cc_288 N_A_435_99#_M1009_g N_VPWR_c_861_n 0.00462271f $X=6.005 $Y=2.4 $X2=0
+ $Y2=0
cc_289 N_A_435_99#_M1014_g N_VPWR_c_861_n 0.00462271f $X=6.615 $Y=2.4 $X2=0
+ $Y2=0
cc_290 N_A_435_99#_M1018_g N_VPWR_c_861_n 0.0046086f $X=7.065 $Y=2.4 $X2=0 $Y2=0
cc_291 N_A_435_99#_M1020_g N_VPWR_c_861_n 0.0046086f $X=7.515 $Y=2.4 $X2=0 $Y2=0
cc_292 N_A_435_99#_M1009_g N_COUT_c_1015_n 0.0028995f $X=6.005 $Y=2.4 $X2=0
+ $Y2=0
cc_293 N_A_435_99#_M1014_g N_COUT_c_1015_n 0.0146272f $X=6.615 $Y=2.4 $X2=0
+ $Y2=0
cc_294 N_A_435_99#_M1018_g N_COUT_c_1015_n 0.0205967f $X=7.065 $Y=2.4 $X2=0
+ $Y2=0
cc_295 N_A_435_99#_c_220_n N_COUT_c_1015_n 0.0287016f $X=5.88 $Y=1.985 $X2=0
+ $Y2=0
cc_296 N_A_435_99#_c_285_p N_COUT_c_1015_n 0.0574349f $X=6.79 $Y=1.485 $X2=0
+ $Y2=0
cc_297 N_A_435_99#_c_211_n N_COUT_c_1015_n 0.00813057f $X=7.515 $Y=1.485 $X2=0
+ $Y2=0
cc_298 N_A_435_99#_M1010_g N_COUT_c_1012_n 0.00335135f $X=6.3 $Y=0.74 $X2=0
+ $Y2=0
cc_299 N_A_435_99#_c_285_p N_COUT_c_1012_n 0.0192803f $X=6.79 $Y=1.485 $X2=0
+ $Y2=0
cc_300 N_A_435_99#_c_211_n N_COUT_c_1012_n 0.00269228f $X=7.515 $Y=1.485 $X2=0
+ $Y2=0
cc_301 N_A_435_99#_M1010_g N_COUT_c_1013_n 0.0067313f $X=6.3 $Y=0.74 $X2=0 $Y2=0
cc_302 N_A_435_99#_M1012_g N_COUT_c_1013_n 3.97481e-19 $X=6.73 $Y=0.74 $X2=0
+ $Y2=0
cc_303 N_A_435_99#_M1012_g N_COUT_c_1014_n 0.0147737f $X=6.73 $Y=0.74 $X2=0
+ $Y2=0
cc_304 N_A_435_99#_M1032_g N_COUT_c_1014_n 0.0163818f $X=7.16 $Y=0.74 $X2=0
+ $Y2=0
cc_305 N_A_435_99#_c_285_p N_COUT_c_1014_n 0.024649f $X=6.79 $Y=1.485 $X2=0
+ $Y2=0
cc_306 N_A_435_99#_c_211_n N_COUT_c_1014_n 0.00326012f $X=7.515 $Y=1.485 $X2=0
+ $Y2=0
cc_307 N_A_435_99#_M1032_g N_COUT_c_1032_n 0.001989f $X=7.16 $Y=0.74 $X2=0 $Y2=0
cc_308 N_A_435_99#_M1033_g N_COUT_c_1032_n 0.00705268f $X=7.59 $Y=0.74 $X2=0
+ $Y2=0
cc_309 N_A_435_99#_M1012_g COUT 9.18327e-19 $X=6.73 $Y=0.74 $X2=0 $Y2=0
cc_310 N_A_435_99#_M1018_g COUT 0.00462744f $X=7.065 $Y=2.4 $X2=0 $Y2=0
cc_311 N_A_435_99#_M1032_g COUT 0.00571358f $X=7.16 $Y=0.74 $X2=0 $Y2=0
cc_312 N_A_435_99#_M1020_g COUT 0.00447206f $X=7.515 $Y=2.4 $X2=0 $Y2=0
cc_313 N_A_435_99#_M1033_g COUT 0.005924f $X=7.59 $Y=0.74 $X2=0 $Y2=0
cc_314 N_A_435_99#_c_285_p COUT 0.0189686f $X=6.79 $Y=1.485 $X2=0 $Y2=0
cc_315 N_A_435_99#_c_211_n COUT 0.0227808f $X=7.515 $Y=1.485 $X2=0 $Y2=0
cc_316 N_A_435_99#_M1020_g N_COUT_c_1041_n 0.00800125f $X=7.515 $Y=2.4 $X2=0
+ $Y2=0
cc_317 N_A_435_99#_c_196_n N_A_27_125#_c_1157_n 0.00197658f $X=2.25 $Y=1.34
+ $X2=0 $Y2=0
cc_318 N_A_435_99#_c_196_n N_A_27_125#_c_1158_n 0.00371137f $X=2.25 $Y=1.34
+ $X2=0 $Y2=0
cc_319 N_A_435_99#_c_199_n N_A_27_125#_c_1158_n 0.00330783f $X=2.72 $Y=1.34
+ $X2=0 $Y2=0
cc_320 N_A_435_99#_c_199_n N_A_27_125#_c_1160_n 0.0155464f $X=2.72 $Y=1.34 $X2=0
+ $Y2=0
cc_321 N_A_435_99#_c_208_n N_A_27_125#_c_1160_n 0.00783057f $X=3.9 $Y=1.57 $X2=0
+ $Y2=0
cc_322 N_A_435_99#_c_209_n N_A_27_125#_c_1160_n 0.0110379f $X=3.24 $Y=1.57 $X2=0
+ $Y2=0
cc_323 N_A_435_99#_M1010_g N_VGND_c_1222_n 0.00511131f $X=6.3 $Y=0.74 $X2=0
+ $Y2=0
cc_324 N_A_435_99#_c_210_n N_VGND_c_1222_n 0.010681f $X=6.05 $Y=1.485 $X2=0
+ $Y2=0
cc_325 N_A_435_99#_c_285_p N_VGND_c_1222_n 0.00919629f $X=6.79 $Y=1.485 $X2=0
+ $Y2=0
cc_326 N_A_435_99#_c_211_n N_VGND_c_1222_n 0.0041377f $X=7.515 $Y=1.485 $X2=0
+ $Y2=0
cc_327 N_A_435_99#_M1010_g N_VGND_c_1223_n 4.53155e-19 $X=6.3 $Y=0.74 $X2=0
+ $Y2=0
cc_328 N_A_435_99#_M1012_g N_VGND_c_1223_n 0.00813302f $X=6.73 $Y=0.74 $X2=0
+ $Y2=0
cc_329 N_A_435_99#_M1032_g N_VGND_c_1223_n 0.0105568f $X=7.16 $Y=0.74 $X2=0
+ $Y2=0
cc_330 N_A_435_99#_M1033_g N_VGND_c_1223_n 0.00138519f $X=7.59 $Y=0.74 $X2=0
+ $Y2=0
cc_331 N_A_435_99#_M1032_g N_VGND_c_1224_n 0.00138519f $X=7.16 $Y=0.74 $X2=0
+ $Y2=0
cc_332 N_A_435_99#_M1033_g N_VGND_c_1224_n 0.0113816f $X=7.59 $Y=0.74 $X2=0
+ $Y2=0
cc_333 N_A_435_99#_M1032_g N_VGND_c_1232_n 0.00383152f $X=7.16 $Y=0.74 $X2=0
+ $Y2=0
cc_334 N_A_435_99#_M1033_g N_VGND_c_1232_n 0.00383152f $X=7.59 $Y=0.74 $X2=0
+ $Y2=0
cc_335 N_A_435_99#_M1010_g N_VGND_c_1237_n 0.00434272f $X=6.3 $Y=0.74 $X2=0
+ $Y2=0
cc_336 N_A_435_99#_M1012_g N_VGND_c_1237_n 0.00383152f $X=6.73 $Y=0.74 $X2=0
+ $Y2=0
cc_337 N_A_435_99#_M1010_g N_VGND_c_1242_n 0.00825283f $X=6.3 $Y=0.74 $X2=0
+ $Y2=0
cc_338 N_A_435_99#_M1012_g N_VGND_c_1242_n 0.0075754f $X=6.73 $Y=0.74 $X2=0
+ $Y2=0
cc_339 N_A_435_99#_M1032_g N_VGND_c_1242_n 0.0075754f $X=7.16 $Y=0.74 $X2=0
+ $Y2=0
cc_340 N_A_435_99#_M1033_g N_VGND_c_1242_n 0.0075754f $X=7.59 $Y=0.74 $X2=0
+ $Y2=0
cc_341 N_A_435_99#_c_208_n N_A_707_119#_c_1344_n 0.0218973f $X=3.9 $Y=1.57 $X2=0
+ $Y2=0
cc_342 N_A_435_99#_c_237_p N_A_707_119#_c_1345_n 0.0207073f $X=4.115 $Y=0.74
+ $X2=0 $Y2=0
cc_343 N_A_435_99#_c_237_p N_A_707_119#_c_1347_n 0.0351355f $X=4.115 $Y=0.74
+ $X2=0 $Y2=0
cc_344 N_A_435_99#_c_223_n N_A_707_119#_c_1347_n 0.00163629f $X=4.07 $Y=1.907
+ $X2=0 $Y2=0
cc_345 N_A_435_99#_c_220_n N_A_707_119#_c_1348_n 0.0181607f $X=5.88 $Y=1.985
+ $X2=0 $Y2=0
cc_346 N_A_435_99#_c_210_n N_A_707_119#_c_1348_n 0.015926f $X=6.05 $Y=1.485
+ $X2=0 $Y2=0
cc_347 N_A_435_99#_c_224_n N_A_707_119#_c_1348_n 0.0397923f $X=4.955 $Y=1.985
+ $X2=0 $Y2=0
cc_348 N_A_435_99#_c_211_n N_A_707_119#_c_1348_n 6.87859e-19 $X=7.515 $Y=1.485
+ $X2=0 $Y2=0
cc_349 N_A_435_99#_c_223_n N_A_707_119#_c_1349_n 0.0133289f $X=4.07 $Y=1.907
+ $X2=0 $Y2=0
cc_350 N_A_435_99#_c_224_n N_A_707_119#_c_1349_n 0.0224714f $X=4.955 $Y=1.985
+ $X2=0 $Y2=0
cc_351 N_A_435_99#_M1010_g N_A_707_119#_c_1350_n 0.00559358f $X=6.3 $Y=0.74
+ $X2=0 $Y2=0
cc_352 N_A_435_99#_c_210_n N_A_707_119#_c_1350_n 0.00906645f $X=6.05 $Y=1.485
+ $X2=0 $Y2=0
cc_353 N_A_435_99#_c_211_n N_A_707_119#_c_1350_n 3.53737e-19 $X=7.515 $Y=1.485
+ $X2=0 $Y2=0
cc_354 N_B_M1002_g N_A_M1022_g 0.0108461f $X=1.36 $Y=0.945 $X2=0 $Y2=0
cc_355 N_B_c_392_n N_A_c_521_n 0.00806011f $X=1.395 $Y=1.88 $X2=0 $Y2=0
cc_356 N_B_M1002_g N_A_c_509_n 0.00894529f $X=1.36 $Y=0.945 $X2=0 $Y2=0
cc_357 N_B_M1007_g N_A_c_509_n 0.00879826f $X=1.79 $Y=0.945 $X2=0 $Y2=0
cc_358 N_B_M1000_g N_A_c_509_n 0.00880809f $X=3.9 $Y=0.915 $X2=0 $Y2=0
cc_359 N_B_M1003_g N_A_c_509_n 0.00880809f $X=4.33 $Y=0.915 $X2=0 $Y2=0
cc_360 N_B_c_388_n N_A_M1029_g 0.0044794f $X=4.255 $Y=1.605 $X2=0 $Y2=0
cc_361 N_B_M1025_g N_A_M1029_g 0.0373678f $X=4.37 $Y=2.47 $X2=0 $Y2=0
cc_362 N_B_M1003_g N_A_M1004_g 0.0185653f $X=4.33 $Y=0.915 $X2=0 $Y2=0
cc_363 N_B_M1003_g N_A_c_516_n 0.0044794f $X=4.33 $Y=0.915 $X2=0 $Y2=0
cc_364 N_B_c_386_n A 0.0117291f $X=1.935 $Y=1.805 $X2=0 $Y2=0
cc_365 B A 0.0204071f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_366 N_B_c_386_n N_A_c_519_n 0.0264528f $X=1.935 $Y=1.805 $X2=0 $Y2=0
cc_367 N_B_c_393_n N_A_297_392#_c_639_n 0.0146579f $X=1.845 $Y=1.88 $X2=0 $Y2=0
cc_368 N_B_c_394_n N_A_297_392#_c_639_n 0.00353142f $X=2.28 $Y=1.805 $X2=0 $Y2=0
cc_369 N_B_c_396_n N_A_297_392#_c_639_n 0.0164254f $X=2.355 $Y=3.075 $X2=0 $Y2=0
cc_370 B N_A_297_392#_c_639_n 0.0398371f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_371 N_B_M1007_g N_A_297_392#_c_631_n 3.97112e-19 $X=1.79 $Y=0.945 $X2=0 $Y2=0
cc_372 N_B_c_394_n N_A_297_392#_c_631_n 0.00367419f $X=2.28 $Y=1.805 $X2=0 $Y2=0
cc_373 N_B_c_386_n N_A_297_392#_c_631_n 8.30845e-19 $X=1.935 $Y=1.805 $X2=0
+ $Y2=0
cc_374 B N_A_297_392#_c_631_n 0.0222825f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_375 N_B_M1008_g N_A_297_392#_c_658_n 0.0171639f $X=3.765 $Y=2.315 $X2=0 $Y2=0
cc_376 N_B_c_400_n N_A_297_392#_c_660_n 0.00266868f $X=4.28 $Y=3.15 $X2=0 $Y2=0
cc_377 N_B_M1025_g N_A_297_392#_c_660_n 0.0141516f $X=4.37 $Y=2.47 $X2=0 $Y2=0
cc_378 N_B_c_392_n N_A_297_392#_c_642_n 0.0111414f $X=1.395 $Y=1.88 $X2=0 $Y2=0
cc_379 N_B_c_386_n N_A_297_392#_c_642_n 0.00259573f $X=1.935 $Y=1.805 $X2=0
+ $Y2=0
cc_380 B N_A_297_392#_c_642_n 0.0143373f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_381 N_B_c_394_n N_A_297_392#_c_634_n 6.73123e-19 $X=2.28 $Y=1.805 $X2=0 $Y2=0
cc_382 N_B_c_396_n N_A_297_392#_c_643_n 0.00159405f $X=2.355 $Y=3.075 $X2=0
+ $Y2=0
cc_383 N_B_c_396_n N_A_297_392#_c_676_n 4.96612e-19 $X=2.355 $Y=3.075 $X2=0
+ $Y2=0
cc_384 N_B_M1008_g N_A_297_392#_c_676_n 0.00107343f $X=3.765 $Y=2.315 $X2=0
+ $Y2=0
cc_385 N_B_c_400_n N_A_297_392#_c_680_n 0.00298749f $X=4.28 $Y=3.15 $X2=0 $Y2=0
cc_386 N_B_M1025_g N_A_297_392#_c_680_n 0.00351821f $X=4.37 $Y=2.47 $X2=0 $Y2=0
cc_387 N_B_c_390_n N_A_297_392#_c_680_n 6.05565e-19 $X=3.825 $Y=1.605 $X2=0
+ $Y2=0
cc_388 N_B_c_392_n N_A_27_392#_c_824_n 0.0139961f $X=1.395 $Y=1.88 $X2=0 $Y2=0
cc_389 N_B_c_393_n N_A_27_392#_c_824_n 0.0136071f $X=1.845 $Y=1.88 $X2=0 $Y2=0
cc_390 N_B_c_396_n N_A_27_392#_c_824_n 0.00178843f $X=2.355 $Y=3.075 $X2=0 $Y2=0
cc_391 N_B_c_392_n N_A_27_392#_c_826_n 5.92432e-19 $X=1.395 $Y=1.88 $X2=0 $Y2=0
cc_392 N_B_c_393_n N_A_27_392#_c_826_n 0.00929817f $X=1.845 $Y=1.88 $X2=0 $Y2=0
cc_393 N_B_c_396_n N_A_27_392#_c_826_n 0.00793964f $X=2.355 $Y=3.075 $X2=0 $Y2=0
cc_394 N_B_c_396_n N_VPWR_c_863_n 0.00943712f $X=2.355 $Y=3.075 $X2=0 $Y2=0
cc_395 N_B_c_397_n N_VPWR_c_863_n 0.0228202f $X=3.675 $Y=3.15 $X2=0 $Y2=0
cc_396 N_B_c_397_n N_VPWR_c_864_n 0.0169345f $X=3.675 $Y=3.15 $X2=0 $Y2=0
cc_397 N_B_M1008_g N_VPWR_c_864_n 0.0185483f $X=3.765 $Y=2.315 $X2=0 $Y2=0
cc_398 N_B_M1025_g N_VPWR_c_864_n 0.00335233f $X=4.37 $Y=2.47 $X2=0 $Y2=0
cc_399 N_B_c_404_n N_VPWR_c_864_n 0.00476669f $X=3.765 $Y=3.15 $X2=0 $Y2=0
cc_400 N_B_M1008_g N_VPWR_c_865_n 0.00145241f $X=3.765 $Y=2.315 $X2=0 $Y2=0
cc_401 N_B_c_400_n N_VPWR_c_865_n 0.00778334f $X=4.28 $Y=3.15 $X2=0 $Y2=0
cc_402 N_B_M1025_g N_VPWR_c_865_n 0.0138637f $X=4.37 $Y=2.47 $X2=0 $Y2=0
cc_403 N_B_c_392_n N_VPWR_c_880_n 0.00333926f $X=1.395 $Y=1.88 $X2=0 $Y2=0
cc_404 N_B_c_393_n N_VPWR_c_880_n 0.00333896f $X=1.845 $Y=1.88 $X2=0 $Y2=0
cc_405 N_B_c_398_n N_VPWR_c_880_n 0.00757097f $X=2.43 $Y=3.15 $X2=0 $Y2=0
cc_406 N_B_c_397_n N_VPWR_c_881_n 0.0200847f $X=3.675 $Y=3.15 $X2=0 $Y2=0
cc_407 N_B_c_404_n N_VPWR_c_882_n 0.0273024f $X=3.765 $Y=3.15 $X2=0 $Y2=0
cc_408 N_B_c_392_n N_VPWR_c_861_n 0.00422798f $X=1.395 $Y=1.88 $X2=0 $Y2=0
cc_409 N_B_c_393_n N_VPWR_c_861_n 0.00423401f $X=1.845 $Y=1.88 $X2=0 $Y2=0
cc_410 N_B_c_397_n N_VPWR_c_861_n 0.0266924f $X=3.675 $Y=3.15 $X2=0 $Y2=0
cc_411 N_B_c_398_n N_VPWR_c_861_n 0.0114097f $X=2.43 $Y=3.15 $X2=0 $Y2=0
cc_412 N_B_c_400_n N_VPWR_c_861_n 0.0188444f $X=4.28 $Y=3.15 $X2=0 $Y2=0
cc_413 N_B_c_404_n N_VPWR_c_861_n 0.00904288f $X=3.765 $Y=3.15 $X2=0 $Y2=0
cc_414 N_B_M1002_g N_A_27_125#_c_1156_n 0.015945f $X=1.36 $Y=0.945 $X2=0 $Y2=0
cc_415 N_B_M1007_g N_A_27_125#_c_1156_n 0.0118929f $X=1.79 $Y=0.945 $X2=0 $Y2=0
cc_416 N_B_c_394_n N_A_27_125#_c_1156_n 0.00102103f $X=2.28 $Y=1.805 $X2=0 $Y2=0
cc_417 N_B_c_386_n N_A_27_125#_c_1156_n 0.00460258f $X=1.935 $Y=1.805 $X2=0
+ $Y2=0
cc_418 B N_A_27_125#_c_1156_n 0.0488126f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_419 N_B_M1002_g N_A_27_125#_c_1157_n 6.55263e-19 $X=1.36 $Y=0.945 $X2=0 $Y2=0
cc_420 N_B_M1007_g N_A_27_125#_c_1157_n 0.00945767f $X=1.79 $Y=0.945 $X2=0 $Y2=0
cc_421 N_B_M1000_g N_A_27_125#_c_1160_n 0.00165882f $X=3.9 $Y=0.915 $X2=0 $Y2=0
cc_422 N_B_M1002_g N_VGND_c_1219_n 0.0073425f $X=1.36 $Y=0.945 $X2=0 $Y2=0
cc_423 N_B_M1007_g N_VGND_c_1219_n 9.59856e-19 $X=1.79 $Y=0.945 $X2=0 $Y2=0
cc_424 N_B_M1002_g N_VGND_c_1242_n 7.97988e-19 $X=1.36 $Y=0.945 $X2=0 $Y2=0
cc_425 N_B_M1007_g N_VGND_c_1242_n 7.94319e-19 $X=1.79 $Y=0.945 $X2=0 $Y2=0
cc_426 N_B_M1000_g N_A_707_119#_c_1344_n 0.00320107f $X=3.9 $Y=0.915 $X2=0 $Y2=0
cc_427 N_B_c_390_n N_A_707_119#_c_1344_n 5.7345e-19 $X=3.825 $Y=1.605 $X2=0
+ $Y2=0
cc_428 N_B_M1000_g N_A_707_119#_c_1345_n 0.0076245f $X=3.9 $Y=0.915 $X2=0 $Y2=0
cc_429 N_B_M1003_g N_A_707_119#_c_1345_n 0.00750518f $X=4.33 $Y=0.915 $X2=0
+ $Y2=0
cc_430 N_B_M1003_g N_A_707_119#_c_1347_n 0.00665243f $X=4.33 $Y=0.915 $X2=0
+ $Y2=0
cc_431 N_B_M1003_g N_A_707_119#_c_1349_n 0.0021197f $X=4.33 $Y=0.915 $X2=0 $Y2=0
cc_432 N_A_M1029_g N_A_297_392#_c_660_n 0.0144762f $X=4.82 $Y=2.47 $X2=0 $Y2=0
cc_433 N_A_M1034_g N_A_297_392#_c_660_n 0.0145175f $X=5.345 $Y=2.26 $X2=0 $Y2=0
cc_434 A N_A_27_392#_c_820_n 0.023f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_435 N_A_M1016_g N_A_27_392#_c_822_n 0.0141975f $X=0.495 $Y=2.46 $X2=0 $Y2=0
cc_436 N_A_c_521_n N_A_27_392#_c_822_n 0.0128963f $X=0.945 $Y=1.875 $X2=0 $Y2=0
cc_437 A N_A_27_392#_c_822_n 0.0453755f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_438 N_A_c_519_n N_A_27_392#_c_822_n 0.00201785f $X=0.93 $Y=1.665 $X2=0 $Y2=0
cc_439 N_A_c_521_n N_A_27_392#_c_823_n 7.50501e-19 $X=0.945 $Y=1.875 $X2=0 $Y2=0
cc_440 A N_A_27_392#_c_823_n 0.0219786f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_441 N_A_M1016_g N_A_27_392#_c_840_n 4.43017e-19 $X=0.495 $Y=2.46 $X2=0 $Y2=0
cc_442 N_A_c_521_n N_A_27_392#_c_840_n 0.0105956f $X=0.945 $Y=1.875 $X2=0 $Y2=0
cc_443 N_A_c_521_n N_A_27_392#_c_825_n 0.00347836f $X=0.945 $Y=1.875 $X2=0 $Y2=0
cc_444 N_A_M1016_g N_VPWR_c_862_n 0.0152538f $X=0.495 $Y=2.46 $X2=0 $Y2=0
cc_445 N_A_c_521_n N_VPWR_c_862_n 0.00126302f $X=0.945 $Y=1.875 $X2=0 $Y2=0
cc_446 N_A_M1029_g N_VPWR_c_865_n 0.0148013f $X=4.82 $Y=2.47 $X2=0 $Y2=0
cc_447 N_A_M1034_g N_VPWR_c_865_n 6.94575e-19 $X=5.345 $Y=2.26 $X2=0 $Y2=0
cc_448 N_A_M1029_g N_VPWR_c_866_n 0.00526206f $X=4.82 $Y=2.47 $X2=0 $Y2=0
cc_449 N_A_M1034_g N_VPWR_c_866_n 0.00482866f $X=5.345 $Y=2.26 $X2=0 $Y2=0
cc_450 N_A_M1029_g N_VPWR_c_867_n 0.00569925f $X=4.82 $Y=2.47 $X2=0 $Y2=0
cc_451 N_A_M1034_g N_VPWR_c_867_n 0.00421725f $X=5.345 $Y=2.26 $X2=0 $Y2=0
cc_452 N_A_M1016_g N_VPWR_c_879_n 0.00460063f $X=0.495 $Y=2.46 $X2=0 $Y2=0
cc_453 N_A_c_521_n N_VPWR_c_880_n 0.00517089f $X=0.945 $Y=1.875 $X2=0 $Y2=0
cc_454 N_A_M1016_g N_VPWR_c_861_n 0.00912261f $X=0.495 $Y=2.46 $X2=0 $Y2=0
cc_455 N_A_c_521_n N_VPWR_c_861_n 0.00977588f $X=0.945 $Y=1.875 $X2=0 $Y2=0
cc_456 N_A_M1029_g N_VPWR_c_861_n 0.00527162f $X=4.82 $Y=2.47 $X2=0 $Y2=0
cc_457 N_A_M1034_g N_VPWR_c_861_n 0.00555093f $X=5.345 $Y=2.26 $X2=0 $Y2=0
cc_458 N_A_M1013_g N_A_27_125#_c_1152_n 4.43891e-19 $X=0.495 $Y=0.945 $X2=0
+ $Y2=0
cc_459 N_A_M1013_g N_A_27_125#_c_1153_n 0.0124643f $X=0.495 $Y=0.945 $X2=0 $Y2=0
cc_460 N_A_M1022_g N_A_27_125#_c_1153_n 0.0111806f $X=0.93 $Y=0.945 $X2=0 $Y2=0
cc_461 A N_A_27_125#_c_1153_n 0.0452882f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_462 N_A_c_519_n N_A_27_125#_c_1153_n 0.00280866f $X=0.93 $Y=1.665 $X2=0 $Y2=0
cc_463 A N_A_27_125#_c_1154_n 0.0212308f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_464 N_A_M1013_g N_A_27_125#_c_1155_n 5.76881e-19 $X=0.495 $Y=0.945 $X2=0
+ $Y2=0
cc_465 N_A_M1022_g N_A_27_125#_c_1155_n 0.00743339f $X=0.93 $Y=0.945 $X2=0 $Y2=0
cc_466 N_A_c_509_n N_A_27_125#_c_1155_n 0.0026496f $X=4.755 $Y=0.18 $X2=0 $Y2=0
cc_467 A N_A_27_125#_c_1156_n 0.00646543f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_468 N_A_c_509_n N_A_27_125#_c_1158_n 0.0189417f $X=4.755 $Y=0.18 $X2=0 $Y2=0
cc_469 N_A_c_509_n N_A_27_125#_c_1159_n 0.00772631f $X=4.755 $Y=0.18 $X2=0 $Y2=0
cc_470 N_A_M1022_g N_A_27_125#_c_1161_n 9.55648e-19 $X=0.93 $Y=0.945 $X2=0 $Y2=0
cc_471 A N_A_27_125#_c_1161_n 0.0218994f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_472 N_A_M1013_g N_VGND_c_1218_n 0.0104167f $X=0.495 $Y=0.945 $X2=0 $Y2=0
cc_473 N_A_c_510_n N_VGND_c_1218_n 0.013498f $X=1.005 $Y=0.18 $X2=0 $Y2=0
cc_474 N_A_M1022_g N_VGND_c_1219_n 0.00475281f $X=0.93 $Y=0.945 $X2=0 $Y2=0
cc_475 N_A_c_509_n N_VGND_c_1219_n 0.0203576f $X=4.755 $Y=0.18 $X2=0 $Y2=0
cc_476 N_A_c_509_n N_VGND_c_1220_n 0.0164781f $X=4.755 $Y=0.18 $X2=0 $Y2=0
cc_477 N_A_c_513_n N_VGND_c_1220_n 0.00455437f $X=5.255 $Y=1.47 $X2=0 $Y2=0
cc_478 N_A_c_514_n N_VGND_c_1220_n 0.0125021f $X=5.33 $Y=1.31 $X2=0 $Y2=0
cc_479 N_A_c_514_n N_VGND_c_1221_n 0.0035863f $X=5.33 $Y=1.31 $X2=0 $Y2=0
cc_480 N_A_c_514_n N_VGND_c_1222_n 0.00261122f $X=5.33 $Y=1.31 $X2=0 $Y2=0
cc_481 N_A_M1013_g N_VGND_c_1228_n 0.00345209f $X=0.495 $Y=0.945 $X2=0 $Y2=0
cc_482 N_A_c_510_n N_VGND_c_1230_n 0.0177193f $X=1.005 $Y=0.18 $X2=0 $Y2=0
cc_483 N_A_c_509_n N_VGND_c_1236_n 0.0773131f $X=4.755 $Y=0.18 $X2=0 $Y2=0
cc_484 N_A_M1013_g N_VGND_c_1242_n 0.00394323f $X=0.495 $Y=0.945 $X2=0 $Y2=0
cc_485 N_A_c_509_n N_VGND_c_1242_n 0.109515f $X=4.755 $Y=0.18 $X2=0 $Y2=0
cc_486 N_A_c_510_n N_VGND_c_1242_n 0.0106926f $X=1.005 $Y=0.18 $X2=0 $Y2=0
cc_487 N_A_c_514_n N_VGND_c_1242_n 0.00401353f $X=5.33 $Y=1.31 $X2=0 $Y2=0
cc_488 N_A_c_509_n N_A_707_119#_c_1345_n 0.0156098f $X=4.755 $Y=0.18 $X2=0 $Y2=0
cc_489 N_A_M1004_g N_A_707_119#_c_1345_n 0.00599831f $X=4.83 $Y=0.915 $X2=0
+ $Y2=0
cc_490 N_A_c_509_n N_A_707_119#_c_1346_n 0.00626586f $X=4.755 $Y=0.18 $X2=0
+ $Y2=0
cc_491 N_A_M1004_g N_A_707_119#_c_1347_n 0.01109f $X=4.83 $Y=0.915 $X2=0 $Y2=0
cc_492 N_A_c_514_n N_A_707_119#_c_1347_n 4.9686e-19 $X=5.33 $Y=1.31 $X2=0 $Y2=0
cc_493 N_A_c_516_n N_A_707_119#_c_1347_n 0.00685332f $X=4.73 $Y=1.46 $X2=0 $Y2=0
cc_494 N_A_c_513_n N_A_707_119#_c_1348_n 0.0144444f $X=5.255 $Y=1.47 $X2=0 $Y2=0
cc_495 N_A_c_516_n N_A_707_119#_c_1348_n 0.00979406f $X=4.73 $Y=1.46 $X2=0 $Y2=0
cc_496 N_A_c_517_n N_A_707_119#_c_1348_n 0.0143326f $X=5.255 $Y=1.31 $X2=0 $Y2=0
cc_497 N_A_c_516_n N_A_707_119#_c_1349_n 0.0040889f $X=4.73 $Y=1.46 $X2=0 $Y2=0
cc_498 N_A_c_514_n N_A_707_119#_c_1350_n 0.00688907f $X=5.33 $Y=1.31 $X2=0 $Y2=0
cc_499 N_A_297_392#_c_639_n N_A_27_392#_M1021_s 0.00226423f $X=2.5 $Y=2.04 $X2=0
+ $Y2=0
cc_500 N_A_297_392#_c_642_n N_A_27_392#_c_823_n 0.0064751f $X=1.62 $Y=2.12 $X2=0
+ $Y2=0
cc_501 N_A_297_392#_M1019_d N_A_27_392#_c_824_n 0.00165831f $X=1.485 $Y=1.96
+ $X2=0 $Y2=0
cc_502 N_A_297_392#_c_642_n N_A_27_392#_c_824_n 0.0139027f $X=1.62 $Y=2.12 $X2=0
+ $Y2=0
cc_503 N_A_297_392#_c_639_n N_A_27_392#_c_826_n 0.0219457f $X=2.5 $Y=2.04 $X2=0
+ $Y2=0
cc_504 N_A_297_392#_c_656_n N_VPWR_M1001_s 0.00132463f $X=2.925 $Y=2.015 $X2=0
+ $Y2=0
cc_505 N_A_297_392#_c_643_n N_VPWR_M1001_s 0.00228391f $X=2.585 $Y=2.015 $X2=0
+ $Y2=0
cc_506 N_A_297_392#_c_658_n N_VPWR_M1006_s 0.00425857f $X=3.9 $Y=2.25 $X2=0
+ $Y2=0
cc_507 N_A_297_392#_c_660_n N_VPWR_M1025_s 0.00388327f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_508 N_A_297_392#_c_660_n N_VPWR_M1034_s 0.00885391f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_509 N_A_297_392#_c_660_n N_VPWR_M1014_s 0.00323047f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_510 N_A_297_392#_c_660_n N_VPWR_M1020_s 0.00402005f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_511 N_A_297_392#_c_641_n N_VPWR_M1020_s 0.00444503f $X=7.81 $Y=2.32 $X2=0
+ $Y2=0
cc_512 N_A_297_392#_c_639_n N_VPWR_c_863_n 0.00140427f $X=2.5 $Y=2.04 $X2=0
+ $Y2=0
cc_513 N_A_297_392#_c_656_n N_VPWR_c_863_n 0.00420031f $X=2.925 $Y=2.015 $X2=0
+ $Y2=0
cc_514 N_A_297_392#_c_643_n N_VPWR_c_863_n 0.0105347f $X=2.585 $Y=2.015 $X2=0
+ $Y2=0
cc_515 N_A_297_392#_c_658_n N_VPWR_c_864_n 0.0170259f $X=3.9 $Y=2.25 $X2=0 $Y2=0
cc_516 N_A_297_392#_c_660_n N_VPWR_c_865_n 0.0166513f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_517 N_A_297_392#_c_660_n N_VPWR_c_867_n 0.0312856f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_518 N_A_297_392#_c_660_n N_VPWR_c_868_n 0.0166513f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_519 N_A_297_392#_M1024_g N_VPWR_c_869_n 0.00847469f $X=7.965 $Y=2.4 $X2=0
+ $Y2=0
cc_520 N_A_297_392#_M1027_g N_VPWR_c_869_n 4.09989e-19 $X=8.415 $Y=2.4 $X2=0
+ $Y2=0
cc_521 N_A_297_392#_c_660_n N_VPWR_c_869_n 0.0168473f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_522 N_A_297_392#_M1024_g N_VPWR_c_870_n 5.02386e-19 $X=7.965 $Y=2.4 $X2=0
+ $Y2=0
cc_523 N_A_297_392#_M1027_g N_VPWR_c_870_n 0.0124373f $X=8.415 $Y=2.4 $X2=0
+ $Y2=0
cc_524 N_A_297_392#_M1031_g N_VPWR_c_870_n 0.0147111f $X=8.865 $Y=2.4 $X2=0
+ $Y2=0
cc_525 N_A_297_392#_M1035_g N_VPWR_c_870_n 6.19991e-19 $X=9.575 $Y=2.4 $X2=0
+ $Y2=0
cc_526 N_A_297_392#_M1031_g N_VPWR_c_872_n 5.99329e-19 $X=8.865 $Y=2.4 $X2=0
+ $Y2=0
cc_527 N_A_297_392#_M1035_g N_VPWR_c_872_n 0.0149079f $X=9.575 $Y=2.4 $X2=0
+ $Y2=0
cc_528 N_A_297_392#_M1024_g N_VPWR_c_877_n 0.00460063f $X=7.965 $Y=2.4 $X2=0
+ $Y2=0
cc_529 N_A_297_392#_M1027_g N_VPWR_c_877_n 0.00460063f $X=8.415 $Y=2.4 $X2=0
+ $Y2=0
cc_530 N_A_297_392#_M1031_g N_VPWR_c_883_n 0.00460063f $X=8.865 $Y=2.4 $X2=0
+ $Y2=0
cc_531 N_A_297_392#_M1035_g N_VPWR_c_883_n 0.00460063f $X=9.575 $Y=2.4 $X2=0
+ $Y2=0
cc_532 N_A_297_392#_M1024_g N_VPWR_c_861_n 0.00908554f $X=7.965 $Y=2.4 $X2=0
+ $Y2=0
cc_533 N_A_297_392#_M1027_g N_VPWR_c_861_n 0.00908554f $X=8.415 $Y=2.4 $X2=0
+ $Y2=0
cc_534 N_A_297_392#_M1031_g N_VPWR_c_861_n 0.00910651f $X=8.865 $Y=2.4 $X2=0
+ $Y2=0
cc_535 N_A_297_392#_M1035_g N_VPWR_c_861_n 0.00910651f $X=9.575 $Y=2.4 $X2=0
+ $Y2=0
cc_536 N_A_297_392#_c_660_n N_VPWR_c_861_n 0.0800807f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_537 N_A_297_392#_c_680_n N_VPWR_c_861_n 0.00553057f $X=3.985 $Y=2.25 $X2=0
+ $Y2=0
cc_538 N_A_297_392#_c_660_n N_COUT_M1009_d 0.0108272f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_539 N_A_297_392#_c_660_n N_COUT_M1018_d 0.00472722f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_540 N_A_297_392#_c_660_n N_COUT_c_1015_n 0.0565079f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_541 N_A_297_392#_M1005_g N_COUT_c_1032_n 7.75513e-19 $X=8.02 $Y=0.74 $X2=0
+ $Y2=0
cc_542 N_A_297_392#_M1005_g COUT 9.08516e-19 $X=8.02 $Y=0.74 $X2=0 $Y2=0
cc_543 N_A_297_392#_c_627_n COUT 4.33563e-19 $X=9.025 $Y=1.485 $X2=0 $Y2=0
cc_544 N_A_297_392#_c_641_n COUT 0.0127061f $X=7.81 $Y=2.32 $X2=0 $Y2=0
cc_545 N_A_297_392#_c_632_n COUT 0.027912f $X=7.895 $Y=1.485 $X2=0 $Y2=0
cc_546 N_A_297_392#_M1024_g N_COUT_c_1041_n 3.00627e-19 $X=7.965 $Y=2.4 $X2=0
+ $Y2=0
cc_547 N_A_297_392#_c_660_n N_COUT_c_1041_n 0.0225105f $X=7.725 $Y=2.405 $X2=0
+ $Y2=0
cc_548 N_A_297_392#_c_641_n N_COUT_c_1041_n 0.0259638f $X=7.81 $Y=2.32 $X2=0
+ $Y2=0
cc_549 N_A_297_392#_c_627_n N_SUM_c_1070_n 0.00225438f $X=9.025 $Y=1.485 $X2=0
+ $Y2=0
cc_550 N_A_297_392#_c_641_n N_SUM_c_1070_n 0.011581f $X=7.81 $Y=2.32 $X2=0 $Y2=0
cc_551 N_A_297_392#_c_757_p N_SUM_c_1070_n 0.0193994f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_552 N_A_297_392#_M1024_g N_SUM_c_1071_n 4.039e-19 $X=7.965 $Y=2.4 $X2=0 $Y2=0
cc_553 N_A_297_392#_M1027_g N_SUM_c_1071_n 4.039e-19 $X=8.415 $Y=2.4 $X2=0 $Y2=0
cc_554 N_A_297_392#_M1005_g N_SUM_c_1063_n 3.97481e-19 $X=8.02 $Y=0.74 $X2=0
+ $Y2=0
cc_555 N_A_297_392#_M1015_g N_SUM_c_1063_n 0.00903544f $X=8.45 $Y=0.74 $X2=0
+ $Y2=0
cc_556 N_A_297_392#_M1026_g N_SUM_c_1063_n 6.75677e-19 $X=8.95 $Y=0.74 $X2=0
+ $Y2=0
cc_557 N_A_297_392#_M1015_g N_SUM_c_1064_n 0.0115433f $X=8.45 $Y=0.74 $X2=0
+ $Y2=0
cc_558 N_A_297_392#_M1026_g N_SUM_c_1064_n 0.0153874f $X=8.95 $Y=0.74 $X2=0
+ $Y2=0
cc_559 N_A_297_392#_c_627_n N_SUM_c_1064_n 0.00420549f $X=9.025 $Y=1.485 $X2=0
+ $Y2=0
cc_560 N_A_297_392#_c_757_p N_SUM_c_1064_n 0.0492199f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_561 N_A_297_392#_M1005_g N_SUM_c_1065_n 6.07621e-19 $X=8.02 $Y=0.74 $X2=0
+ $Y2=0
cc_562 N_A_297_392#_M1015_g N_SUM_c_1065_n 0.00110424f $X=8.45 $Y=0.74 $X2=0
+ $Y2=0
cc_563 N_A_297_392#_c_627_n N_SUM_c_1065_n 0.00252677f $X=9.025 $Y=1.485 $X2=0
+ $Y2=0
cc_564 N_A_297_392#_c_757_p N_SUM_c_1065_n 0.0209731f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_565 N_A_297_392#_M1026_g N_SUM_c_1066_n 0.00377577f $X=8.95 $Y=0.74 $X2=0
+ $Y2=0
cc_566 N_A_297_392#_M1030_g N_SUM_c_1066_n 5.54424e-19 $X=9.505 $Y=0.74 $X2=0
+ $Y2=0
cc_567 N_A_297_392#_M1031_g N_SUM_c_1072_n 0.0119155f $X=8.865 $Y=2.4 $X2=0
+ $Y2=0
cc_568 N_A_297_392#_M1035_g N_SUM_c_1072_n 0.0123461f $X=9.575 $Y=2.4 $X2=0
+ $Y2=0
cc_569 N_A_297_392#_M1030_g N_SUM_c_1067_n 0.015246f $X=9.505 $Y=0.74 $X2=0
+ $Y2=0
cc_570 N_A_297_392#_c_757_p N_SUM_c_1067_n 0.0177771f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_571 N_A_297_392#_c_633_n N_SUM_c_1067_n 0.00397982f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_572 N_A_297_392#_M1035_g N_SUM_c_1073_n 0.0288069f $X=9.575 $Y=2.4 $X2=0
+ $Y2=0
cc_573 N_A_297_392#_c_757_p N_SUM_c_1073_n 0.017083f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_574 N_A_297_392#_c_633_n N_SUM_c_1073_n 0.00171112f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_575 N_A_297_392#_M1030_g N_SUM_c_1068_n 0.00533837f $X=9.505 $Y=0.74 $X2=0
+ $Y2=0
cc_576 N_A_297_392#_M1035_g N_SUM_c_1068_n 0.0059715f $X=9.575 $Y=2.4 $X2=0
+ $Y2=0
cc_577 N_A_297_392#_c_757_p N_SUM_c_1068_n 0.0250942f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_578 N_A_297_392#_c_633_n N_SUM_c_1068_n 0.00951237f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_579 N_A_297_392#_c_626_n N_SUM_c_1069_n 0.00524152f $X=9.43 $Y=1.485 $X2=0
+ $Y2=0
cc_580 N_A_297_392#_c_757_p N_SUM_c_1069_n 0.0278321f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_581 N_A_297_392#_M1027_g N_SUM_c_1075_n 0.0196002f $X=8.415 $Y=2.4 $X2=0
+ $Y2=0
cc_582 N_A_297_392#_M1031_g N_SUM_c_1075_n 0.0217567f $X=8.865 $Y=2.4 $X2=0
+ $Y2=0
cc_583 N_A_297_392#_c_626_n N_SUM_c_1075_n 7.99111e-19 $X=9.43 $Y=1.485 $X2=0
+ $Y2=0
cc_584 N_A_297_392#_c_627_n N_SUM_c_1075_n 0.0021292f $X=9.025 $Y=1.485 $X2=0
+ $Y2=0
cc_585 N_A_297_392#_c_757_p N_SUM_c_1075_n 0.0574814f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_586 N_A_297_392#_c_626_n N_SUM_c_1076_n 0.00782931f $X=9.43 $Y=1.485 $X2=0
+ $Y2=0
cc_587 N_A_297_392#_c_757_p N_SUM_c_1076_n 0.0262158f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_588 N_A_297_392#_c_757_p N_SUM_c_1117_n 0.0032968f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_589 N_A_297_392#_M1031_g N_SUM_c_1118_n 0.00676779f $X=8.865 $Y=2.4 $X2=0
+ $Y2=0
cc_590 N_A_297_392#_c_757_p N_SUM_c_1118_n 0.00167912f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_591 N_A_297_392#_c_642_n N_A_27_125#_c_1156_n 0.00340883f $X=1.62 $Y=2.12
+ $X2=0 $Y2=0
cc_592 N_A_297_392#_c_634_n N_A_27_125#_c_1156_n 0.00167954f $X=2.505 $Y=1.285
+ $X2=0 $Y2=0
cc_593 N_A_297_392#_c_630_n N_A_27_125#_c_1157_n 0.00158095f $X=2.505 $Y=0.77
+ $X2=0 $Y2=0
cc_594 N_A_297_392#_c_630_n N_A_27_125#_c_1158_n 0.0258724f $X=2.505 $Y=0.77
+ $X2=0 $Y2=0
cc_595 N_A_297_392#_c_630_n N_A_27_125#_c_1160_n 0.0243921f $X=2.505 $Y=0.77
+ $X2=0 $Y2=0
cc_596 N_A_297_392#_c_656_n N_A_27_125#_c_1160_n 0.00208042f $X=2.925 $Y=2.015
+ $X2=0 $Y2=0
cc_597 N_A_297_392#_c_676_n N_A_27_125#_c_1160_n 0.00360966f $X=3.09 $Y=2.07
+ $X2=0 $Y2=0
cc_598 N_A_297_392#_M1005_g N_VGND_c_1224_n 0.00842225f $X=8.02 $Y=0.74 $X2=0
+ $Y2=0
cc_599 N_A_297_392#_M1015_g N_VGND_c_1224_n 4.51782e-19 $X=8.45 $Y=0.74 $X2=0
+ $Y2=0
cc_600 N_A_297_392#_c_632_n N_VGND_c_1224_n 0.00597123f $X=7.895 $Y=1.485 $X2=0
+ $Y2=0
cc_601 N_A_297_392#_c_757_p N_VGND_c_1224_n 0.00128723f $X=9.56 $Y=1.485 $X2=0
+ $Y2=0
cc_602 N_A_297_392#_M1015_g N_VGND_c_1225_n 0.00408259f $X=8.45 $Y=0.74 $X2=0
+ $Y2=0
cc_603 N_A_297_392#_M1026_g N_VGND_c_1225_n 0.00997407f $X=8.95 $Y=0.74 $X2=0
+ $Y2=0
cc_604 N_A_297_392#_M1030_g N_VGND_c_1225_n 6.10235e-19 $X=9.505 $Y=0.74 $X2=0
+ $Y2=0
cc_605 N_A_297_392#_M1030_g N_VGND_c_1227_n 0.00694336f $X=9.505 $Y=0.74 $X2=0
+ $Y2=0
cc_606 N_A_297_392#_M1005_g N_VGND_c_1234_n 0.00383152f $X=8.02 $Y=0.74 $X2=0
+ $Y2=0
cc_607 N_A_297_392#_M1015_g N_VGND_c_1234_n 0.00434272f $X=8.45 $Y=0.74 $X2=0
+ $Y2=0
cc_608 N_A_297_392#_M1026_g N_VGND_c_1238_n 0.00383152f $X=8.95 $Y=0.74 $X2=0
+ $Y2=0
cc_609 N_A_297_392#_M1030_g N_VGND_c_1238_n 0.00460063f $X=9.505 $Y=0.74 $X2=0
+ $Y2=0
cc_610 N_A_297_392#_M1005_g N_VGND_c_1242_n 0.0075754f $X=8.02 $Y=0.74 $X2=0
+ $Y2=0
cc_611 N_A_297_392#_M1015_g N_VGND_c_1242_n 0.00820718f $X=8.45 $Y=0.74 $X2=0
+ $Y2=0
cc_612 N_A_297_392#_M1026_g N_VGND_c_1242_n 0.00758657f $X=8.95 $Y=0.74 $X2=0
+ $Y2=0
cc_613 N_A_297_392#_M1030_g N_VGND_c_1242_n 0.00912119f $X=9.505 $Y=0.74 $X2=0
+ $Y2=0
cc_614 N_A_27_392#_c_822_n N_VPWR_M1016_d 0.00165831f $X=1.005 $Y=2.04 $X2=-0.19
+ $Y2=1.66
cc_615 N_A_27_392#_c_821_n N_VPWR_c_862_n 0.0242552f $X=0.27 $Y=2.8 $X2=0 $Y2=0
cc_616 N_A_27_392#_c_822_n N_VPWR_c_862_n 0.0148589f $X=1.005 $Y=2.04 $X2=0
+ $Y2=0
cc_617 N_A_27_392#_c_825_n N_VPWR_c_862_n 0.0103534f $X=1.255 $Y=2.99 $X2=0
+ $Y2=0
cc_618 N_A_27_392#_c_824_n N_VPWR_c_863_n 0.0117895f $X=1.905 $Y=2.99 $X2=0
+ $Y2=0
cc_619 N_A_27_392#_c_826_n N_VPWR_c_863_n 0.0326488f $X=2.07 $Y=2.38 $X2=0 $Y2=0
cc_620 N_A_27_392#_c_821_n N_VPWR_c_879_n 0.0116996f $X=0.27 $Y=2.8 $X2=0 $Y2=0
cc_621 N_A_27_392#_c_824_n N_VPWR_c_880_n 0.0644071f $X=1.905 $Y=2.99 $X2=0
+ $Y2=0
cc_622 N_A_27_392#_c_825_n N_VPWR_c_880_n 0.0178163f $X=1.255 $Y=2.99 $X2=0
+ $Y2=0
cc_623 N_A_27_392#_c_821_n N_VPWR_c_861_n 0.0101742f $X=0.27 $Y=2.8 $X2=0 $Y2=0
cc_624 N_A_27_392#_c_824_n N_VPWR_c_861_n 0.0356218f $X=1.905 $Y=2.99 $X2=0
+ $Y2=0
cc_625 N_A_27_392#_c_825_n N_VPWR_c_861_n 0.00958215f $X=1.255 $Y=2.99 $X2=0
+ $Y2=0
cc_626 N_A_27_392#_c_820_n N_A_27_125#_c_1154_n 3.57272e-19 $X=0.245 $Y=2.125
+ $X2=0 $Y2=0
cc_627 N_VPWR_M1014_s N_COUT_c_1015_n 0.00169665f $X=6.705 $Y=1.84 $X2=0 $Y2=0
cc_628 N_VPWR_c_869_n N_SUM_c_1071_n 0.0127556f $X=7.74 $Y=2.78 $X2=0 $Y2=0
cc_629 N_VPWR_c_870_n N_SUM_c_1071_n 0.0255132f $X=8.64 $Y=2.405 $X2=0 $Y2=0
cc_630 N_VPWR_c_877_n N_SUM_c_1071_n 0.0101736f $X=8.475 $Y=3.33 $X2=0 $Y2=0
cc_631 N_VPWR_c_861_n N_SUM_c_1071_n 0.0084208f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_632 N_VPWR_c_870_n N_SUM_c_1072_n 0.0359677f $X=8.64 $Y=2.405 $X2=0 $Y2=0
cc_633 N_VPWR_c_872_n N_SUM_c_1072_n 0.0406515f $X=9.8 $Y=2.415 $X2=0 $Y2=0
cc_634 N_VPWR_c_883_n N_SUM_c_1072_n 0.0146357f $X=9.635 $Y=3.33 $X2=0 $Y2=0
cc_635 N_VPWR_c_861_n N_SUM_c_1072_n 0.0121141f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_636 N_VPWR_M1035_s N_SUM_c_1073_n 4.81498e-19 $X=9.665 $Y=1.84 $X2=0 $Y2=0
cc_637 N_VPWR_c_872_n N_SUM_c_1073_n 0.0098937f $X=9.8 $Y=2.415 $X2=0 $Y2=0
cc_638 N_VPWR_M1035_s N_SUM_c_1068_n 0.00227995f $X=9.665 $Y=1.84 $X2=0 $Y2=0
cc_639 N_VPWR_c_872_n N_SUM_c_1068_n 0.0101282f $X=9.8 $Y=2.415 $X2=0 $Y2=0
cc_640 N_VPWR_M1027_s N_SUM_c_1075_n 0.00169251f $X=8.505 $Y=1.84 $X2=0 $Y2=0
cc_641 N_VPWR_c_870_n N_SUM_c_1075_n 0.0181933f $X=8.64 $Y=2.405 $X2=0 $Y2=0
cc_642 N_VPWR_c_872_n N_SUM_c_1117_n 4.31246e-19 $X=9.8 $Y=2.415 $X2=0 $Y2=0
cc_643 N_VPWR_c_870_n N_SUM_c_1118_n 0.00182758f $X=8.64 $Y=2.405 $X2=0 $Y2=0
cc_644 N_VPWR_M1035_s SUM 0.00184365f $X=9.665 $Y=1.84 $X2=0 $Y2=0
cc_645 N_VPWR_c_872_n SUM 0.00488527f $X=9.8 $Y=2.415 $X2=0 $Y2=0
cc_646 N_COUT_c_1032_n N_SUM_c_1065_n 0.00260272f $X=7.382 $Y=1.13 $X2=0 $Y2=0
cc_647 COUT N_SUM_c_1065_n 6.38315e-19 $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_648 N_COUT_c_1014_n N_VGND_M1012_d 0.00178571f $X=7.21 $Y=1.005 $X2=0 $Y2=0
cc_649 N_COUT_c_1012_n N_VGND_c_1222_n 0.0107873f $X=6.475 $Y=0.88 $X2=0 $Y2=0
cc_650 N_COUT_c_1013_n N_VGND_c_1222_n 0.0188983f $X=6.515 $Y=0.515 $X2=0 $Y2=0
cc_651 N_COUT_c_1013_n N_VGND_c_1223_n 0.0136308f $X=6.515 $Y=0.515 $X2=0 $Y2=0
cc_652 N_COUT_c_1014_n N_VGND_c_1223_n 0.0175375f $X=7.21 $Y=1.005 $X2=0 $Y2=0
cc_653 N_COUT_c_1013_n N_VGND_c_1237_n 0.0109942f $X=6.515 $Y=0.515 $X2=0 $Y2=0
cc_654 N_COUT_c_1013_n N_VGND_c_1242_n 0.00904371f $X=6.515 $Y=0.515 $X2=0 $Y2=0
cc_655 N_SUM_c_1064_n N_VGND_M1015_d 0.00250873f $X=9.07 $Y=1.065 $X2=0 $Y2=0
cc_656 N_SUM_c_1067_n N_VGND_M1030_d 0.00317529f $X=9.825 $Y=1.065 $X2=0 $Y2=0
cc_657 N_SUM_c_1063_n N_VGND_c_1224_n 0.0136308f $X=8.235 $Y=0.515 $X2=0 $Y2=0
cc_658 N_SUM_c_1063_n N_VGND_c_1225_n 0.0173318f $X=8.235 $Y=0.515 $X2=0 $Y2=0
cc_659 N_SUM_c_1064_n N_VGND_c_1225_n 0.0210288f $X=9.07 $Y=1.065 $X2=0 $Y2=0
cc_660 N_SUM_c_1066_n N_VGND_c_1225_n 0.0180508f $X=9.235 $Y=0.515 $X2=0 $Y2=0
cc_661 N_SUM_c_1066_n N_VGND_c_1227_n 0.0157236f $X=9.235 $Y=0.515 $X2=0 $Y2=0
cc_662 N_SUM_c_1067_n N_VGND_c_1227_n 0.0206457f $X=9.825 $Y=1.065 $X2=0 $Y2=0
cc_663 N_SUM_c_1063_n N_VGND_c_1234_n 0.0109942f $X=8.235 $Y=0.515 $X2=0 $Y2=0
cc_664 N_SUM_c_1066_n N_VGND_c_1238_n 0.0146357f $X=9.235 $Y=0.515 $X2=0 $Y2=0
cc_665 N_SUM_c_1063_n N_VGND_c_1242_n 0.00904371f $X=8.235 $Y=0.515 $X2=0 $Y2=0
cc_666 N_SUM_c_1066_n N_VGND_c_1242_n 0.0121141f $X=9.235 $Y=0.515 $X2=0 $Y2=0
cc_667 N_A_27_125#_c_1153_n N_VGND_M1013_s 0.00177524f $X=0.98 $Y=1.2 $X2=-0.19
+ $Y2=-0.245
cc_668 N_A_27_125#_c_1156_n N_VGND_M1002_d 0.00176461f $X=1.84 $Y=1.2 $X2=0
+ $Y2=0
cc_669 N_A_27_125#_c_1152_n N_VGND_c_1218_n 0.0124064f $X=0.28 $Y=0.77 $X2=0
+ $Y2=0
cc_670 N_A_27_125#_c_1153_n N_VGND_c_1218_n 0.015373f $X=0.98 $Y=1.2 $X2=0 $Y2=0
cc_671 N_A_27_125#_c_1155_n N_VGND_c_1218_n 0.0237383f $X=1.145 $Y=0.77 $X2=0
+ $Y2=0
cc_672 N_A_27_125#_c_1155_n N_VGND_c_1219_n 0.0124064f $X=1.145 $Y=0.77 $X2=0
+ $Y2=0
cc_673 N_A_27_125#_c_1156_n N_VGND_c_1219_n 0.0152916f $X=1.84 $Y=1.2 $X2=0
+ $Y2=0
cc_674 N_A_27_125#_c_1157_n N_VGND_c_1219_n 0.0257313f $X=2.005 $Y=0.77 $X2=0
+ $Y2=0
cc_675 N_A_27_125#_c_1159_n N_VGND_c_1219_n 0.0141601f $X=2.17 $Y=0.35 $X2=0
+ $Y2=0
cc_676 N_A_27_125#_c_1152_n N_VGND_c_1228_n 0.00535163f $X=0.28 $Y=0.77 $X2=0
+ $Y2=0
cc_677 N_A_27_125#_c_1155_n N_VGND_c_1230_n 0.00529024f $X=1.145 $Y=0.77 $X2=0
+ $Y2=0
cc_678 N_A_27_125#_c_1158_n N_VGND_c_1236_n 0.0627959f $X=2.84 $Y=0.35 $X2=0
+ $Y2=0
cc_679 N_A_27_125#_c_1159_n N_VGND_c_1236_n 0.0222408f $X=2.17 $Y=0.35 $X2=0
+ $Y2=0
cc_680 N_A_27_125#_c_1152_n N_VGND_c_1242_n 0.00769355f $X=0.28 $Y=0.77 $X2=0
+ $Y2=0
cc_681 N_A_27_125#_c_1155_n N_VGND_c_1242_n 0.00666603f $X=1.145 $Y=0.77 $X2=0
+ $Y2=0
cc_682 N_A_27_125#_c_1158_n N_VGND_c_1242_n 0.0338116f $X=2.84 $Y=0.35 $X2=0
+ $Y2=0
cc_683 N_A_27_125#_c_1159_n N_VGND_c_1242_n 0.0114525f $X=2.17 $Y=0.35 $X2=0
+ $Y2=0
cc_684 N_A_27_125#_c_1160_n N_A_707_119#_c_1344_n 0.0372071f $X=3.005 $Y=0.77
+ $X2=0 $Y2=0
cc_685 N_A_27_125#_c_1158_n N_A_707_119#_c_1346_n 0.00679393f $X=2.84 $Y=0.35
+ $X2=0 $Y2=0
cc_686 N_A_27_125#_c_1160_n N_A_707_119#_c_1346_n 0.00265323f $X=3.005 $Y=0.77
+ $X2=0 $Y2=0
cc_687 N_VGND_c_1220_n N_A_707_119#_c_1345_n 0.0142636f $X=5.115 $Y=0.74 $X2=0
+ $Y2=0
cc_688 N_VGND_c_1236_n N_A_707_119#_c_1345_n 0.048346f $X=4.95 $Y=0 $X2=0 $Y2=0
cc_689 N_VGND_c_1242_n N_A_707_119#_c_1345_n 0.0326371f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_690 N_VGND_c_1236_n N_A_707_119#_c_1346_n 0.0134803f $X=4.95 $Y=0 $X2=0 $Y2=0
cc_691 N_VGND_c_1242_n N_A_707_119#_c_1346_n 0.00875888f $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_692 N_VGND_c_1220_n N_A_707_119#_c_1347_n 0.0341802f $X=5.115 $Y=0.74 $X2=0
+ $Y2=0
cc_693 N_VGND_c_1220_n N_A_707_119#_c_1348_n 0.0263226f $X=5.115 $Y=0.74 $X2=0
+ $Y2=0
cc_694 N_VGND_c_1220_n N_A_707_119#_c_1350_n 0.025828f $X=5.115 $Y=0.74 $X2=0
+ $Y2=0
cc_695 N_VGND_c_1221_n N_A_707_119#_c_1350_n 0.00571886f $X=5.92 $Y=0 $X2=0
+ $Y2=0
cc_696 N_VGND_c_1222_n N_A_707_119#_c_1350_n 0.0382129f $X=6.085 $Y=0.515 $X2=0
+ $Y2=0
cc_697 N_VGND_c_1242_n N_A_707_119#_c_1350_n 0.00786368f $X=9.84 $Y=0 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__ebufn_2.pxi.spice
* Created: Wed Sep  2 12:07:38 2020
* 
x_PM_SKY130_FD_SC_MS__EBUFN_2%A_84_48# N_A_84_48#_M1000_d N_A_84_48#_M1010_d
+ N_A_84_48#_M1008_g N_A_84_48#_M1005_g N_A_84_48#_M1009_g N_A_84_48#_M1007_g
+ N_A_84_48#_c_86_n N_A_84_48#_c_93_n N_A_84_48#_c_94_n N_A_84_48#_c_111_p
+ N_A_84_48#_c_87_n N_A_84_48#_c_95_n N_A_84_48#_c_88_n N_A_84_48#_c_96_n
+ N_A_84_48#_c_89_n N_A_84_48#_c_90_n PM_SKY130_FD_SC_MS__EBUFN_2%A_84_48#
x_PM_SKY130_FD_SC_MS__EBUFN_2%A_283_48# N_A_283_48#_M1011_s N_A_283_48#_M1001_s
+ N_A_283_48#_c_196_n N_A_283_48#_M1002_g N_A_283_48#_c_197_n
+ N_A_283_48#_c_198_n N_A_283_48#_c_199_n N_A_283_48#_M1003_g
+ N_A_283_48#_c_200_n N_A_283_48#_c_201_n N_A_283_48#_c_202_n
+ N_A_283_48#_c_206_n N_A_283_48#_c_207_n N_A_283_48#_c_203_n
+ N_A_283_48#_c_204_n PM_SKY130_FD_SC_MS__EBUFN_2%A_283_48#
x_PM_SKY130_FD_SC_MS__EBUFN_2%TE_B N_TE_B_c_275_n N_TE_B_M1004_g N_TE_B_c_268_n
+ N_TE_B_c_269_n N_TE_B_c_278_n N_TE_B_M1006_g N_TE_B_c_270_n N_TE_B_M1001_g
+ N_TE_B_M1011_g N_TE_B_c_272_n TE_B N_TE_B_c_274_n N_TE_B_c_282_n
+ PM_SKY130_FD_SC_MS__EBUFN_2%TE_B
x_PM_SKY130_FD_SC_MS__EBUFN_2%A N_A_M1000_g N_A_M1010_g A N_A_c_356_n
+ N_A_c_357_n PM_SKY130_FD_SC_MS__EBUFN_2%A
x_PM_SKY130_FD_SC_MS__EBUFN_2%A_33_368# N_A_33_368#_M1005_d N_A_33_368#_M1007_d
+ N_A_33_368#_M1006_s N_A_33_368#_c_391_n N_A_33_368#_c_392_n
+ N_A_33_368#_c_393_n N_A_33_368#_c_402_n N_A_33_368#_c_394_n
+ N_A_33_368#_c_395_n PM_SKY130_FD_SC_MS__EBUFN_2%A_33_368#
x_PM_SKY130_FD_SC_MS__EBUFN_2%Z N_Z_M1008_d N_Z_M1005_s N_Z_c_440_n N_Z_c_435_n
+ N_Z_c_448_n N_Z_c_436_n N_Z_c_438_n Z Z PM_SKY130_FD_SC_MS__EBUFN_2%Z
x_PM_SKY130_FD_SC_MS__EBUFN_2%VPWR N_VPWR_M1004_d N_VPWR_M1001_d N_VPWR_c_476_n
+ VPWR N_VPWR_c_477_n N_VPWR_c_478_n N_VPWR_c_479_n N_VPWR_c_475_n
+ N_VPWR_c_481_n N_VPWR_c_482_n PM_SKY130_FD_SC_MS__EBUFN_2%VPWR
x_PM_SKY130_FD_SC_MS__EBUFN_2%A_27_74# N_A_27_74#_M1008_s N_A_27_74#_M1009_s
+ N_A_27_74#_M1003_s N_A_27_74#_c_522_n N_A_27_74#_c_523_n N_A_27_74#_c_524_n
+ N_A_27_74#_c_525_n N_A_27_74#_c_526_n N_A_27_74#_c_527_n
+ PM_SKY130_FD_SC_MS__EBUFN_2%A_27_74#
x_PM_SKY130_FD_SC_MS__EBUFN_2%VGND N_VGND_M1002_d N_VGND_M1011_d N_VGND_c_563_n
+ N_VGND_c_564_n N_VGND_c_565_n N_VGND_c_566_n VGND N_VGND_c_567_n
+ N_VGND_c_568_n N_VGND_c_569_n N_VGND_c_570_n PM_SKY130_FD_SC_MS__EBUFN_2%VGND
cc_1 VNB N_A_84_48#_M1008_g 0.0267131f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_84_48#_M1005_g 0.00237661f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_3 VNB N_A_84_48#_M1009_g 0.0219916f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_4 VNB N_A_84_48#_M1007_g 0.0017025f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.4
cc_5 VNB N_A_84_48#_c_86_n 0.006822f $X=-0.19 $Y=-0.245 $X2=1.965 $Y2=1.465
cc_6 VNB N_A_84_48#_c_87_n 0.0227309f $X=-0.19 $Y=-0.245 $X2=4.005 $Y2=0.515
cc_7 VNB N_A_84_48#_c_88_n 0.0131174f $X=-0.19 $Y=-0.245 $X2=4.022 $Y2=1.03
cc_8 VNB N_A_84_48#_c_89_n 0.0300599f $X=-0.19 $Y=-0.245 $X2=4.04 $Y2=1.95
cc_9 VNB N_A_84_48#_c_90_n 0.0686298f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.465
cc_10 VNB N_A_283_48#_c_196_n 0.0157819f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.3
cc_11 VNB N_A_283_48#_c_197_n 0.0100196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_283_48#_c_198_n 0.00785843f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.63
cc_13 VNB N_A_283_48#_c_199_n 0.0180733f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_14 VNB N_A_283_48#_c_200_n 0.0317356f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.3
cc_15 VNB N_A_283_48#_c_201_n 0.00411221f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_16 VNB N_A_283_48#_c_202_n 0.00429685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_283_48#_c_203_n 0.0713883f $X=-0.19 $Y=-0.245 $X2=3.875 $Y2=2.325
cc_18 VNB N_A_283_48#_c_204_n 0.0105673f $X=-0.19 $Y=-0.245 $X2=4.022 $Y2=0.515
cc_19 VNB N_TE_B_c_268_n 0.00902204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_TE_B_c_269_n 0.00498041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_TE_B_c_270_n 0.0200546f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_22 VNB N_TE_B_M1011_g 0.0337994f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_23 VNB N_TE_B_c_272_n 0.00445378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB TE_B 0.00265516f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=1.63
cc_25 VNB N_TE_B_c_274_n 0.0296433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_M1000_g 0.0382437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_c_356_n 0.0294963f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_28 VNB N_A_c_357_n 0.00603075f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_29 VNB N_Z_c_435_n 0.00143713f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_30 VNB N_Z_c_436_n 0.00185767f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_31 VNB N_VPWR_c_475_n 0.183584f $X=-0.19 $Y=-0.245 $X2=2.05 $Y2=2.24
cc_32 VNB N_A_27_74#_c_522_n 0.0362285f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_33 VNB N_A_27_74#_c_523_n 0.00655758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_27_74#_c_524_n 0.00931596f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.3
cc_35 VNB N_A_27_74#_c_525_n 0.00423028f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.4
cc_36 VNB N_A_27_74#_c_526_n 0.00276453f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.4
cc_37 VNB N_A_27_74#_c_527_n 0.00206817f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.465
cc_38 VNB N_VGND_c_563_n 0.00563933f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_39 VNB N_VGND_c_564_n 0.0167127f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.4
cc_40 VNB N_VGND_c_565_n 0.0408183f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_41 VNB N_VGND_c_566_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_42 VNB N_VGND_c_567_n 0.039031f $X=-0.19 $Y=-0.245 $X2=1.035 $Y2=2.4
cc_43 VNB N_VGND_c_568_n 0.0199919f $X=-0.19 $Y=-0.245 $X2=4.04 $Y2=2.41
cc_44 VNB N_VGND_c_569_n 0.261479f $X=-0.19 $Y=-0.245 $X2=4.04 $Y2=2.715
cc_45 VNB N_VGND_c_570_n 0.00462376f $X=-0.19 $Y=-0.245 $X2=4.12 $Y2=1.03
cc_46 VPB N_A_84_48#_M1005_g 0.0291781f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.4
cc_47 VPB N_A_84_48#_M1007_g 0.0226878f $X=-0.19 $Y=1.66 $X2=1.035 $Y2=2.4
cc_48 VPB N_A_84_48#_c_93_n 0.00109674f $X=-0.19 $Y=1.66 $X2=2.05 $Y2=2.24
cc_49 VPB N_A_84_48#_c_94_n 0.0124138f $X=-0.19 $Y=1.66 $X2=3.875 $Y2=2.325
cc_50 VPB N_A_84_48#_c_95_n 0.0202496f $X=-0.19 $Y=1.66 $X2=4.04 $Y2=2.715
cc_51 VPB N_A_84_48#_c_96_n 0.0174668f $X=-0.19 $Y=1.66 $X2=4.04 $Y2=2.035
cc_52 VPB N_A_84_48#_c_89_n 0.0125498f $X=-0.19 $Y=1.66 $X2=4.04 $Y2=1.95
cc_53 VPB N_A_283_48#_c_202_n 0.00178921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_283_48#_c_206_n 0.00323181f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.465
cc_55 VPB N_A_283_48#_c_207_n 0.0043156f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.465
cc_56 VPB N_TE_B_c_275_n 0.0202238f $X=-0.19 $Y=1.66 $X2=3.865 $Y2=0.37
cc_57 VPB N_TE_B_c_268_n 0.0130416f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_TE_B_c_269_n 0.00264715f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_TE_B_c_278_n 0.0241245f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_TE_B_c_270_n 0.021231f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_61 VPB N_TE_B_c_272_n 0.00124171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_TE_B_c_274_n 0.00557786f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_TE_B_c_282_n 0.0218596f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.465
cc_64 VPB N_A_M1010_g 0.0265693f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.3
cc_65 VPB N_A_c_356_n 0.00692757f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.4
cc_66 VPB N_A_c_357_n 0.00469509f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.4
cc_67 VPB N_A_33_368#_c_391_n 0.0297839f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.4
cc_68 VPB N_A_33_368#_c_392_n 0.00265439f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_33_368#_c_393_n 0.00965867f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.3
cc_70 VPB N_A_33_368#_c_394_n 0.00238711f $X=-0.19 $Y=1.66 $X2=1.035 $Y2=1.63
cc_71 VPB N_A_33_368#_c_395_n 0.00901991f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.465
cc_72 VPB N_Z_c_435_n 9.10919e-19 $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.4
cc_73 VPB N_Z_c_438_n 0.00234957f $X=-0.19 $Y=1.66 $X2=1.035 $Y2=2.4
cc_74 VPB Z 0.0040183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_476_n 0.0190046f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_76 VPB N_VPWR_c_477_n 0.0416737f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.4
cc_77 VPB N_VPWR_c_478_n 0.0350409f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_479_n 0.0196898f $X=-0.19 $Y=1.66 $X2=2.05 $Y2=1.63
cc_79 VPB N_VPWR_c_475_n 0.088056f $X=-0.19 $Y=1.66 $X2=2.05 $Y2=2.24
cc_80 VPB N_VPWR_c_481_n 0.0138146f $X=-0.19 $Y=1.66 $X2=4.022 $Y2=0.848
cc_81 VPB N_VPWR_c_482_n 0.00920679f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 N_A_84_48#_c_94_n N_A_283_48#_M1001_s 0.011598f $X=3.875 $Y=2.325 $X2=0
+ $Y2=0
cc_83 N_A_84_48#_M1009_g N_A_283_48#_c_196_n 0.025089f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_84 N_A_84_48#_c_86_n N_A_283_48#_c_197_n 0.00720366f $X=1.965 $Y=1.465 $X2=0
+ $Y2=0
cc_85 N_A_84_48#_c_86_n N_A_283_48#_c_198_n 0.00475854f $X=1.965 $Y=1.465 $X2=0
+ $Y2=0
cc_86 N_A_84_48#_c_90_n N_A_283_48#_c_198_n 0.00230752f $X=1.035 $Y=1.465 $X2=0
+ $Y2=0
cc_87 N_A_84_48#_c_86_n N_A_283_48#_c_200_n 0.00411929f $X=1.965 $Y=1.465 $X2=0
+ $Y2=0
cc_88 N_A_84_48#_c_86_n N_A_283_48#_c_201_n 0.00414715f $X=1.965 $Y=1.465 $X2=0
+ $Y2=0
cc_89 N_A_84_48#_c_86_n N_A_283_48#_c_202_n 0.0208807f $X=1.965 $Y=1.465 $X2=0
+ $Y2=0
cc_90 N_A_84_48#_c_93_n N_A_283_48#_c_202_n 0.009984f $X=2.05 $Y=2.24 $X2=0
+ $Y2=0
cc_91 N_A_84_48#_c_93_n N_A_283_48#_c_206_n 0.0143324f $X=2.05 $Y=2.24 $X2=0
+ $Y2=0
cc_92 N_A_84_48#_c_94_n N_A_283_48#_c_206_n 0.0274686f $X=3.875 $Y=2.325 $X2=0
+ $Y2=0
cc_93 N_A_84_48#_c_94_n N_A_283_48#_c_207_n 0.0241284f $X=3.875 $Y=2.325 $X2=0
+ $Y2=0
cc_94 N_A_84_48#_c_93_n N_TE_B_c_275_n 0.0038583f $X=2.05 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_95 N_A_84_48#_c_111_p N_TE_B_c_275_n 0.00277024f $X=2.135 $Y=2.325 $X2=-0.19
+ $Y2=-0.245
cc_96 N_A_84_48#_c_86_n N_TE_B_c_268_n 0.0154854f $X=1.965 $Y=1.465 $X2=0 $Y2=0
cc_97 N_A_84_48#_c_93_n N_TE_B_c_268_n 0.00502138f $X=2.05 $Y=2.24 $X2=0 $Y2=0
cc_98 N_A_84_48#_M1007_g N_TE_B_c_269_n 0.0307073f $X=1.035 $Y=2.4 $X2=0 $Y2=0
cc_99 N_A_84_48#_c_86_n N_TE_B_c_269_n 0.00589245f $X=1.965 $Y=1.465 $X2=0 $Y2=0
cc_100 N_A_84_48#_c_90_n N_TE_B_c_269_n 0.00306818f $X=1.035 $Y=1.465 $X2=0
+ $Y2=0
cc_101 N_A_84_48#_c_93_n N_TE_B_c_278_n 0.0180787f $X=2.05 $Y=2.24 $X2=0 $Y2=0
cc_102 N_A_84_48#_c_94_n N_TE_B_c_278_n 0.0119405f $X=3.875 $Y=2.325 $X2=0 $Y2=0
cc_103 N_A_84_48#_c_111_p N_TE_B_c_278_n 0.00370027f $X=2.135 $Y=2.325 $X2=0
+ $Y2=0
cc_104 N_A_84_48#_c_94_n N_TE_B_c_270_n 0.00288155f $X=3.875 $Y=2.325 $X2=0
+ $Y2=0
cc_105 N_A_84_48#_c_87_n N_TE_B_M1011_g 2.21897e-19 $X=4.005 $Y=0.515 $X2=0
+ $Y2=0
cc_106 N_A_84_48#_c_86_n N_TE_B_c_272_n 0.00209554f $X=1.965 $Y=1.465 $X2=0
+ $Y2=0
cc_107 N_A_84_48#_c_93_n N_TE_B_c_272_n 0.0022263f $X=2.05 $Y=2.24 $X2=0 $Y2=0
cc_108 N_A_84_48#_c_94_n TE_B 0.00450693f $X=3.875 $Y=2.325 $X2=0 $Y2=0
cc_109 N_A_84_48#_c_94_n N_TE_B_c_282_n 0.0210391f $X=3.875 $Y=2.325 $X2=0 $Y2=0
cc_110 N_A_84_48#_c_96_n N_TE_B_c_282_n 0.00222056f $X=4.04 $Y=2.035 $X2=0 $Y2=0
cc_111 N_A_84_48#_c_87_n N_A_M1000_g 0.00575762f $X=4.005 $Y=0.515 $X2=0 $Y2=0
cc_112 N_A_84_48#_c_88_n N_A_M1000_g 0.00293996f $X=4.022 $Y=1.03 $X2=0 $Y2=0
cc_113 N_A_84_48#_c_89_n N_A_M1000_g 0.009227f $X=4.04 $Y=1.95 $X2=0 $Y2=0
cc_114 N_A_84_48#_c_94_n N_A_M1010_g 0.0158595f $X=3.875 $Y=2.325 $X2=0 $Y2=0
cc_115 N_A_84_48#_c_95_n N_A_M1010_g 0.00802093f $X=4.04 $Y=2.715 $X2=0 $Y2=0
cc_116 N_A_84_48#_c_96_n N_A_M1010_g 0.00878771f $X=4.04 $Y=2.035 $X2=0 $Y2=0
cc_117 N_A_84_48#_c_94_n N_A_c_356_n 7.45189e-19 $X=3.875 $Y=2.325 $X2=0 $Y2=0
cc_118 N_A_84_48#_c_88_n N_A_c_356_n 0.00163857f $X=4.022 $Y=1.03 $X2=0 $Y2=0
cc_119 N_A_84_48#_c_89_n N_A_c_356_n 0.0132753f $X=4.04 $Y=1.95 $X2=0 $Y2=0
cc_120 N_A_84_48#_c_94_n N_A_c_357_n 0.0129246f $X=3.875 $Y=2.325 $X2=0 $Y2=0
cc_121 N_A_84_48#_c_88_n N_A_c_357_n 0.00112892f $X=4.022 $Y=1.03 $X2=0 $Y2=0
cc_122 N_A_84_48#_c_89_n N_A_c_357_n 0.0326294f $X=4.04 $Y=1.95 $X2=0 $Y2=0
cc_123 N_A_84_48#_c_94_n N_A_33_368#_M1006_s 0.00672062f $X=3.875 $Y=2.325 $X2=0
+ $Y2=0
cc_124 N_A_84_48#_M1005_g N_A_33_368#_c_391_n 0.0151195f $X=0.535 $Y=2.4 $X2=0
+ $Y2=0
cc_125 N_A_84_48#_M1007_g N_A_33_368#_c_391_n 2.72638e-19 $X=1.035 $Y=2.4 $X2=0
+ $Y2=0
cc_126 N_A_84_48#_M1005_g N_A_33_368#_c_392_n 0.0118818f $X=0.535 $Y=2.4 $X2=0
+ $Y2=0
cc_127 N_A_84_48#_M1007_g N_A_33_368#_c_392_n 0.0135121f $X=1.035 $Y=2.4 $X2=0
+ $Y2=0
cc_128 N_A_84_48#_M1005_g N_A_33_368#_c_393_n 0.00291744f $X=0.535 $Y=2.4 $X2=0
+ $Y2=0
cc_129 N_A_84_48#_c_94_n N_A_33_368#_c_402_n 0.00538854f $X=3.875 $Y=2.325 $X2=0
+ $Y2=0
cc_130 N_A_84_48#_c_111_p N_A_33_368#_c_402_n 0.00870963f $X=2.135 $Y=2.325
+ $X2=0 $Y2=0
cc_131 N_A_84_48#_M1007_g N_A_33_368#_c_394_n 4.1224e-19 $X=1.035 $Y=2.4 $X2=0
+ $Y2=0
cc_132 N_A_84_48#_c_111_p N_A_33_368#_c_394_n 0.00326691f $X=2.135 $Y=2.325
+ $X2=0 $Y2=0
cc_133 N_A_84_48#_c_94_n N_A_33_368#_c_395_n 0.0210366f $X=3.875 $Y=2.325 $X2=0
+ $Y2=0
cc_134 N_A_84_48#_M1008_g N_Z_c_440_n 0.00439897f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A_84_48#_M1009_g N_Z_c_440_n 0.00388974f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A_84_48#_M1008_g N_Z_c_435_n 0.00866774f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_137 N_A_84_48#_M1005_g N_Z_c_435_n 0.00947478f $X=0.535 $Y=2.4 $X2=0 $Y2=0
cc_138 N_A_84_48#_M1009_g N_Z_c_435_n 0.0025553f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A_84_48#_M1007_g N_Z_c_435_n 0.0023381f $X=1.035 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A_84_48#_c_86_n N_Z_c_435_n 0.0249855f $X=1.965 $Y=1.465 $X2=0 $Y2=0
cc_141 N_A_84_48#_c_90_n N_Z_c_435_n 0.0232163f $X=1.035 $Y=1.465 $X2=0 $Y2=0
cc_142 N_A_84_48#_M1007_g N_Z_c_448_n 0.00842746f $X=1.035 $Y=2.4 $X2=0 $Y2=0
cc_143 N_A_84_48#_M1008_g N_Z_c_436_n 0.00379299f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A_84_48#_M1009_g N_Z_c_436_n 0.00426649f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A_84_48#_c_90_n N_Z_c_436_n 0.00165838f $X=1.035 $Y=1.465 $X2=0 $Y2=0
cc_146 N_A_84_48#_M1005_g N_Z_c_438_n 0.0140517f $X=0.535 $Y=2.4 $X2=0 $Y2=0
cc_147 N_A_84_48#_M1007_g N_Z_c_438_n 0.00191449f $X=1.035 $Y=2.4 $X2=0 $Y2=0
cc_148 N_A_84_48#_c_86_n N_Z_c_438_n 0.00829947f $X=1.965 $Y=1.465 $X2=0 $Y2=0
cc_149 N_A_84_48#_c_90_n N_Z_c_438_n 0.0045978f $X=1.035 $Y=1.465 $X2=0 $Y2=0
cc_150 N_A_84_48#_M1007_g Z 0.0186905f $X=1.035 $Y=2.4 $X2=0 $Y2=0
cc_151 N_A_84_48#_c_86_n Z 0.0647541f $X=1.965 $Y=1.465 $X2=0 $Y2=0
cc_152 N_A_84_48#_c_93_n Z 0.028433f $X=2.05 $Y=2.24 $X2=0 $Y2=0
cc_153 N_A_84_48#_c_90_n Z 0.00182536f $X=1.035 $Y=1.465 $X2=0 $Y2=0
cc_154 N_A_84_48#_c_93_n N_VPWR_M1004_d 0.00395544f $X=2.05 $Y=2.24 $X2=-0.19
+ $Y2=-0.245
cc_155 N_A_84_48#_c_111_p N_VPWR_M1004_d 0.00305157f $X=2.135 $Y=2.325 $X2=-0.19
+ $Y2=-0.245
cc_156 N_A_84_48#_c_94_n N_VPWR_M1001_d 0.0145572f $X=3.875 $Y=2.325 $X2=0 $Y2=0
cc_157 N_A_84_48#_c_94_n N_VPWR_c_476_n 0.0275977f $X=3.875 $Y=2.325 $X2=0 $Y2=0
cc_158 N_A_84_48#_c_95_n N_VPWR_c_476_n 0.0102171f $X=4.04 $Y=2.715 $X2=0 $Y2=0
cc_159 N_A_84_48#_M1005_g N_VPWR_c_477_n 0.00333896f $X=0.535 $Y=2.4 $X2=0 $Y2=0
cc_160 N_A_84_48#_M1007_g N_VPWR_c_477_n 0.00333926f $X=1.035 $Y=2.4 $X2=0 $Y2=0
cc_161 N_A_84_48#_c_95_n N_VPWR_c_479_n 0.00975961f $X=4.04 $Y=2.715 $X2=0 $Y2=0
cc_162 N_A_84_48#_M1005_g N_VPWR_c_475_n 0.00427015f $X=0.535 $Y=2.4 $X2=0 $Y2=0
cc_163 N_A_84_48#_M1007_g N_VPWR_c_475_n 0.00423742f $X=1.035 $Y=2.4 $X2=0 $Y2=0
cc_164 N_A_84_48#_c_95_n N_VPWR_c_475_n 0.0111753f $X=4.04 $Y=2.715 $X2=0 $Y2=0
cc_165 N_A_84_48#_M1008_g N_A_27_74#_c_522_n 0.0015901f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_166 N_A_84_48#_M1008_g N_A_27_74#_c_523_n 0.0129836f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_167 N_A_84_48#_M1009_g N_A_27_74#_c_523_n 0.013442f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_168 N_A_84_48#_c_86_n N_A_27_74#_c_525_n 0.0582054f $X=1.965 $Y=1.465 $X2=0
+ $Y2=0
cc_169 N_A_84_48#_M1009_g N_A_27_74#_c_526_n 0.00109932f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_170 N_A_84_48#_c_86_n N_A_27_74#_c_526_n 0.0285318f $X=1.965 $Y=1.465 $X2=0
+ $Y2=0
cc_171 N_A_84_48#_c_90_n N_A_27_74#_c_526_n 0.00404284f $X=1.035 $Y=1.465 $X2=0
+ $Y2=0
cc_172 N_A_84_48#_M1009_g N_VGND_c_563_n 2.65335e-19 $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_173 N_A_84_48#_c_87_n N_VGND_c_564_n 0.0259022f $X=4.005 $Y=0.515 $X2=0 $Y2=0
cc_174 N_A_84_48#_M1008_g N_VGND_c_567_n 0.00278271f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_175 N_A_84_48#_M1009_g N_VGND_c_567_n 0.00278271f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_176 N_A_84_48#_c_87_n N_VGND_c_568_n 0.0161257f $X=4.005 $Y=0.515 $X2=0 $Y2=0
cc_177 N_A_84_48#_M1008_g N_VGND_c_569_n 0.00357086f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_178 N_A_84_48#_M1009_g N_VGND_c_569_n 0.00354644f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_179 N_A_84_48#_c_87_n N_VGND_c_569_n 0.013291f $X=4.005 $Y=0.515 $X2=0 $Y2=0
cc_180 N_A_283_48#_c_197_n N_TE_B_c_268_n 0.0182548f $X=1.85 $Y=1.26 $X2=0 $Y2=0
cc_181 N_A_283_48#_c_198_n N_TE_B_c_269_n 0.0182548f $X=1.565 $Y=1.26 $X2=0
+ $Y2=0
cc_182 N_A_283_48#_c_202_n N_TE_B_c_278_n 0.00205978f $X=2.56 $Y=1.17 $X2=0
+ $Y2=0
cc_183 N_A_283_48#_c_206_n N_TE_B_c_278_n 0.00566976f $X=2.725 $Y=1.945 $X2=0
+ $Y2=0
cc_184 N_A_283_48#_c_200_n N_TE_B_c_270_n 0.0182548f $X=2.395 $Y=1.26 $X2=0
+ $Y2=0
cc_185 N_A_283_48#_c_202_n N_TE_B_c_270_n 0.0221236f $X=2.56 $Y=1.17 $X2=0 $Y2=0
cc_186 N_A_283_48#_c_207_n N_TE_B_c_270_n 0.00982869f $X=2.94 $Y=1.985 $X2=0
+ $Y2=0
cc_187 N_A_283_48#_c_204_n N_TE_B_c_270_n 0.00656082f $X=3.005 $Y=0.515 $X2=0
+ $Y2=0
cc_188 N_A_283_48#_c_202_n N_TE_B_M1011_g 0.00109888f $X=2.56 $Y=1.17 $X2=0
+ $Y2=0
cc_189 N_A_283_48#_c_203_n N_TE_B_M1011_g 0.0183842f $X=2.56 $Y=0.49 $X2=0 $Y2=0
cc_190 N_A_283_48#_c_204_n N_TE_B_M1011_g 0.00832294f $X=3.005 $Y=0.515 $X2=0
+ $Y2=0
cc_191 N_A_283_48#_c_201_n N_TE_B_c_272_n 0.0182548f $X=1.925 $Y=1.26 $X2=0
+ $Y2=0
cc_192 N_A_283_48#_c_202_n TE_B 0.0283543f $X=2.56 $Y=1.17 $X2=0 $Y2=0
cc_193 N_A_283_48#_c_207_n TE_B 0.0109882f $X=2.94 $Y=1.985 $X2=0 $Y2=0
cc_194 N_A_283_48#_c_203_n TE_B 0.00125277f $X=2.56 $Y=0.49 $X2=0 $Y2=0
cc_195 N_A_283_48#_c_204_n TE_B 0.015386f $X=3.005 $Y=0.515 $X2=0 $Y2=0
cc_196 N_A_283_48#_c_200_n N_TE_B_c_274_n 8.25111e-19 $X=2.395 $Y=1.26 $X2=0
+ $Y2=0
cc_197 N_A_283_48#_c_202_n N_TE_B_c_274_n 0.00529176f $X=2.56 $Y=1.17 $X2=0
+ $Y2=0
cc_198 N_A_283_48#_c_204_n N_TE_B_c_274_n 8.62818e-19 $X=3.005 $Y=0.515 $X2=0
+ $Y2=0
cc_199 N_A_283_48#_c_202_n N_TE_B_c_282_n 0.00293513f $X=2.56 $Y=1.17 $X2=0
+ $Y2=0
cc_200 N_A_283_48#_c_207_n N_TE_B_c_282_n 0.00720423f $X=2.94 $Y=1.985 $X2=0
+ $Y2=0
cc_201 N_A_283_48#_c_207_n N_A_M1010_g 0.00107664f $X=2.94 $Y=1.985 $X2=0 $Y2=0
cc_202 N_A_283_48#_c_206_n N_A_33_368#_M1006_s 0.00497033f $X=2.725 $Y=1.945
+ $X2=0 $Y2=0
cc_203 N_A_283_48#_c_198_n Z 2.17732e-19 $X=1.565 $Y=1.26 $X2=0 $Y2=0
cc_204 N_A_283_48#_c_196_n N_A_27_74#_c_523_n 0.00148915f $X=1.49 $Y=1.185 $X2=0
+ $Y2=0
cc_205 N_A_283_48#_c_196_n N_A_27_74#_c_525_n 0.0147594f $X=1.49 $Y=1.185 $X2=0
+ $Y2=0
cc_206 N_A_283_48#_c_197_n N_A_27_74#_c_525_n 0.00230303f $X=1.85 $Y=1.26 $X2=0
+ $Y2=0
cc_207 N_A_283_48#_c_199_n N_A_27_74#_c_525_n 0.012029f $X=1.925 $Y=1.185 $X2=0
+ $Y2=0
cc_208 N_A_283_48#_c_200_n N_A_27_74#_c_525_n 0.00522989f $X=2.395 $Y=1.26 $X2=0
+ $Y2=0
cc_209 N_A_283_48#_c_202_n N_A_27_74#_c_525_n 0.00994473f $X=2.56 $Y=1.17 $X2=0
+ $Y2=0
cc_210 N_A_283_48#_c_203_n N_A_27_74#_c_525_n 0.0012571f $X=2.56 $Y=0.49 $X2=0
+ $Y2=0
cc_211 N_A_283_48#_c_204_n N_A_27_74#_c_525_n 0.00428282f $X=3.005 $Y=0.515
+ $X2=0 $Y2=0
cc_212 N_A_283_48#_c_196_n N_A_27_74#_c_527_n 6.17395e-19 $X=1.49 $Y=1.185 $X2=0
+ $Y2=0
cc_213 N_A_283_48#_c_199_n N_A_27_74#_c_527_n 0.00883931f $X=1.925 $Y=1.185
+ $X2=0 $Y2=0
cc_214 N_A_283_48#_c_203_n N_A_27_74#_c_527_n 0.00224515f $X=2.56 $Y=0.49 $X2=0
+ $Y2=0
cc_215 N_A_283_48#_c_204_n N_A_27_74#_c_527_n 0.0492585f $X=3.005 $Y=0.515 $X2=0
+ $Y2=0
cc_216 N_A_283_48#_c_196_n N_VGND_c_563_n 0.00803879f $X=1.49 $Y=1.185 $X2=0
+ $Y2=0
cc_217 N_A_283_48#_c_199_n N_VGND_c_563_n 0.00291064f $X=1.925 $Y=1.185 $X2=0
+ $Y2=0
cc_218 N_A_283_48#_c_204_n N_VGND_c_563_n 7.47461e-19 $X=3.005 $Y=0.515 $X2=0
+ $Y2=0
cc_219 N_A_283_48#_c_204_n N_VGND_c_564_n 0.0305673f $X=3.005 $Y=0.515 $X2=0
+ $Y2=0
cc_220 N_A_283_48#_c_199_n N_VGND_c_565_n 0.00434272f $X=1.925 $Y=1.185 $X2=0
+ $Y2=0
cc_221 N_A_283_48#_c_203_n N_VGND_c_565_n 0.00804684f $X=2.56 $Y=0.49 $X2=0
+ $Y2=0
cc_222 N_A_283_48#_c_204_n N_VGND_c_565_n 0.0371632f $X=3.005 $Y=0.515 $X2=0
+ $Y2=0
cc_223 N_A_283_48#_c_196_n N_VGND_c_567_n 0.00398535f $X=1.49 $Y=1.185 $X2=0
+ $Y2=0
cc_224 N_A_283_48#_c_196_n N_VGND_c_569_n 0.0078875f $X=1.49 $Y=1.185 $X2=0
+ $Y2=0
cc_225 N_A_283_48#_c_199_n N_VGND_c_569_n 0.00825333f $X=1.925 $Y=1.185 $X2=0
+ $Y2=0
cc_226 N_A_283_48#_c_203_n N_VGND_c_569_n 0.0114187f $X=2.56 $Y=0.49 $X2=0 $Y2=0
cc_227 N_A_283_48#_c_204_n N_VGND_c_569_n 0.0286628f $X=3.005 $Y=0.515 $X2=0
+ $Y2=0
cc_228 N_TE_B_M1011_g N_A_M1000_g 0.0255424f $X=3.22 $Y=0.69 $X2=0 $Y2=0
cc_229 TE_B N_A_M1000_g 9.57049e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_230 N_TE_B_c_274_n N_A_M1010_g 0.00109605f $X=3.13 $Y=1.485 $X2=0 $Y2=0
cc_231 N_TE_B_c_282_n N_A_M1010_g 0.0294302f $X=3.13 $Y=1.725 $X2=0 $Y2=0
cc_232 TE_B N_A_c_356_n 3.46758e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_233 N_TE_B_c_274_n N_A_c_356_n 0.0177927f $X=3.13 $Y=1.485 $X2=0 $Y2=0
cc_234 TE_B N_A_c_357_n 0.0220909f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_235 N_TE_B_c_274_n N_A_c_357_n 0.00384747f $X=3.13 $Y=1.485 $X2=0 $Y2=0
cc_236 N_TE_B_c_282_n N_A_c_357_n 0.00133862f $X=3.13 $Y=1.725 $X2=0 $Y2=0
cc_237 N_TE_B_c_275_n N_A_33_368#_c_402_n 0.0120453f $X=1.535 $Y=1.725 $X2=0
+ $Y2=0
cc_238 N_TE_B_c_278_n N_A_33_368#_c_402_n 0.0106713f $X=2.155 $Y=1.725 $X2=0
+ $Y2=0
cc_239 N_TE_B_c_275_n N_A_33_368#_c_394_n 0.0138313f $X=1.535 $Y=1.725 $X2=0
+ $Y2=0
cc_240 N_TE_B_c_278_n N_A_33_368#_c_394_n 0.00170449f $X=2.155 $Y=1.725 $X2=0
+ $Y2=0
cc_241 N_TE_B_c_275_n N_A_33_368#_c_395_n 8.44357e-19 $X=1.535 $Y=1.725 $X2=0
+ $Y2=0
cc_242 N_TE_B_c_278_n N_A_33_368#_c_395_n 0.0065863f $X=2.155 $Y=1.725 $X2=0
+ $Y2=0
cc_243 N_TE_B_c_282_n N_A_33_368#_c_395_n 0.0101219f $X=3.13 $Y=1.725 $X2=0
+ $Y2=0
cc_244 N_TE_B_c_275_n N_Z_c_448_n 7.23397e-19 $X=1.535 $Y=1.725 $X2=0 $Y2=0
cc_245 N_TE_B_c_275_n Z 0.0206424f $X=1.535 $Y=1.725 $X2=0 $Y2=0
cc_246 N_TE_B_c_268_n Z 0.00175072f $X=2.065 $Y=1.65 $X2=0 $Y2=0
cc_247 N_TE_B_c_278_n Z 0.00122241f $X=2.155 $Y=1.725 $X2=0 $Y2=0
cc_248 N_TE_B_c_282_n N_VPWR_c_476_n 0.0234552f $X=3.13 $Y=1.725 $X2=0 $Y2=0
cc_249 N_TE_B_c_275_n N_VPWR_c_477_n 0.00376977f $X=1.535 $Y=1.725 $X2=0 $Y2=0
cc_250 N_TE_B_c_278_n N_VPWR_c_478_n 0.00379565f $X=2.155 $Y=1.725 $X2=0 $Y2=0
cc_251 N_TE_B_c_282_n N_VPWR_c_478_n 0.00492916f $X=3.13 $Y=1.725 $X2=0 $Y2=0
cc_252 N_TE_B_c_275_n N_VPWR_c_475_n 0.00470119f $X=1.535 $Y=1.725 $X2=0 $Y2=0
cc_253 N_TE_B_c_278_n N_VPWR_c_475_n 0.00475768f $X=2.155 $Y=1.725 $X2=0 $Y2=0
cc_254 N_TE_B_c_282_n N_VPWR_c_475_n 0.00511769f $X=3.13 $Y=1.725 $X2=0 $Y2=0
cc_255 N_TE_B_c_275_n N_VPWR_c_481_n 0.00184805f $X=1.535 $Y=1.725 $X2=0 $Y2=0
cc_256 N_TE_B_c_278_n N_VPWR_c_481_n 0.00365882f $X=2.155 $Y=1.725 $X2=0 $Y2=0
cc_257 N_TE_B_c_268_n N_A_27_74#_c_525_n 3.0146e-19 $X=2.065 $Y=1.65 $X2=0 $Y2=0
cc_258 N_TE_B_c_269_n N_A_27_74#_c_525_n 4.06922e-19 $X=1.625 $Y=1.65 $X2=0
+ $Y2=0
cc_259 N_TE_B_M1011_g N_VGND_c_564_n 0.00678145f $X=3.22 $Y=0.69 $X2=0 $Y2=0
cc_260 N_TE_B_M1011_g N_VGND_c_565_n 0.00432591f $X=3.22 $Y=0.69 $X2=0 $Y2=0
cc_261 N_TE_B_M1011_g N_VGND_c_569_n 0.00822267f $X=3.22 $Y=0.69 $X2=0 $Y2=0
cc_262 N_A_M1010_g N_VPWR_c_476_n 0.00555154f $X=3.815 $Y=2.34 $X2=0 $Y2=0
cc_263 N_A_M1010_g N_VPWR_c_479_n 0.00567889f $X=3.815 $Y=2.34 $X2=0 $Y2=0
cc_264 N_A_M1010_g N_VPWR_c_475_n 0.00610055f $X=3.815 $Y=2.34 $X2=0 $Y2=0
cc_265 N_A_M1000_g N_VGND_c_564_n 0.0072585f $X=3.79 $Y=0.69 $X2=0 $Y2=0
cc_266 N_A_c_356_n N_VGND_c_564_n 9.25785e-19 $X=3.7 $Y=1.515 $X2=0 $Y2=0
cc_267 N_A_c_357_n N_VGND_c_564_n 0.00897894f $X=3.7 $Y=1.515 $X2=0 $Y2=0
cc_268 N_A_M1000_g N_VGND_c_568_n 0.00434272f $X=3.79 $Y=0.69 $X2=0 $Y2=0
cc_269 N_A_M1000_g N_VGND_c_569_n 0.00825084f $X=3.79 $Y=0.69 $X2=0 $Y2=0
cc_270 N_A_33_368#_c_392_n N_Z_M1005_s 0.00218982f $X=1.145 $Y=2.99 $X2=0 $Y2=0
cc_271 N_A_33_368#_c_392_n N_Z_c_448_n 0.0177084f $X=1.145 $Y=2.99 $X2=0 $Y2=0
cc_272 N_A_33_368#_M1007_d Z 0.00223902f $X=1.125 $Y=1.84 $X2=0 $Y2=0
cc_273 N_A_33_368#_c_402_n Z 0.00946115f $X=2.215 $Y=2.665 $X2=0 $Y2=0
cc_274 N_A_33_368#_c_394_n Z 0.0198996f $X=1.31 $Y=2.44 $X2=0 $Y2=0
cc_275 N_A_33_368#_c_402_n N_VPWR_M1004_d 0.0128526f $X=2.215 $Y=2.665 $X2=-0.19
+ $Y2=1.66
cc_276 N_A_33_368#_c_392_n N_VPWR_c_477_n 0.0421734f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_277 N_A_33_368#_c_393_n N_VPWR_c_477_n 0.0235512f $X=0.475 $Y=2.99 $X2=0
+ $Y2=0
cc_278 N_A_33_368#_c_402_n N_VPWR_c_477_n 0.00341791f $X=2.215 $Y=2.665 $X2=0
+ $Y2=0
cc_279 N_A_33_368#_c_394_n N_VPWR_c_477_n 0.0234113f $X=1.31 $Y=2.44 $X2=0 $Y2=0
cc_280 N_A_33_368#_c_402_n N_VPWR_c_478_n 0.00341061f $X=2.215 $Y=2.665 $X2=0
+ $Y2=0
cc_281 N_A_33_368#_c_395_n N_VPWR_c_478_n 0.0140093f $X=2.38 $Y=2.665 $X2=0
+ $Y2=0
cc_282 N_A_33_368#_c_392_n N_VPWR_c_475_n 0.0236854f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_283 N_A_33_368#_c_393_n N_VPWR_c_475_n 0.0126924f $X=0.475 $Y=2.99 $X2=0
+ $Y2=0
cc_284 N_A_33_368#_c_402_n N_VPWR_c_475_n 0.0124404f $X=2.215 $Y=2.665 $X2=0
+ $Y2=0
cc_285 N_A_33_368#_c_394_n N_VPWR_c_475_n 0.0126192f $X=1.31 $Y=2.44 $X2=0 $Y2=0
cc_286 N_A_33_368#_c_395_n N_VPWR_c_475_n 0.0117657f $X=2.38 $Y=2.665 $X2=0
+ $Y2=0
cc_287 N_A_33_368#_c_402_n N_VPWR_c_481_n 0.0243979f $X=2.215 $Y=2.665 $X2=0
+ $Y2=0
cc_288 N_A_33_368#_c_394_n N_VPWR_c_481_n 0.00916478f $X=1.31 $Y=2.44 $X2=0
+ $Y2=0
cc_289 N_A_33_368#_c_395_n N_VPWR_c_481_n 0.00263112f $X=2.38 $Y=2.665 $X2=0
+ $Y2=0
cc_290 Z N_VPWR_M1004_d 0.00472472f $X=1.595 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_291 N_Z_c_440_n N_A_27_74#_c_522_n 0.0201328f $X=0.71 $Y=0.78 $X2=0 $Y2=0
cc_292 N_Z_M1008_d N_A_27_74#_c_523_n 0.00184993f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_293 N_Z_c_440_n N_A_27_74#_c_523_n 0.0149881f $X=0.71 $Y=0.78 $X2=0 $Y2=0
cc_294 N_Z_c_436_n N_A_27_74#_c_526_n 0.00732422f $X=0.705 $Y=1.13 $X2=0 $Y2=0
cc_295 N_A_27_74#_c_525_n N_VGND_M1002_d 0.00181776f $X=1.975 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_296 N_A_27_74#_c_523_n N_VGND_c_563_n 0.0114567f $X=1.045 $Y=0.34 $X2=0 $Y2=0
cc_297 N_A_27_74#_c_525_n N_VGND_c_563_n 0.0153175f $X=1.975 $Y=1.045 $X2=0
+ $Y2=0
cc_298 N_A_27_74#_c_527_n N_VGND_c_563_n 0.0158413f $X=2.14 $Y=0.515 $X2=0 $Y2=0
cc_299 N_A_27_74#_c_527_n N_VGND_c_565_n 0.0109942f $X=2.14 $Y=0.515 $X2=0 $Y2=0
cc_300 N_A_27_74#_c_523_n N_VGND_c_567_n 0.0665295f $X=1.045 $Y=0.34 $X2=0 $Y2=0
cc_301 N_A_27_74#_c_524_n N_VGND_c_567_n 0.0179217f $X=0.365 $Y=0.34 $X2=0 $Y2=0
cc_302 N_A_27_74#_c_523_n N_VGND_c_569_n 0.0370229f $X=1.045 $Y=0.34 $X2=0 $Y2=0
cc_303 N_A_27_74#_c_524_n N_VGND_c_569_n 0.00971942f $X=0.365 $Y=0.34 $X2=0
+ $Y2=0
cc_304 N_A_27_74#_c_527_n N_VGND_c_569_n 0.00904371f $X=2.14 $Y=0.515 $X2=0
+ $Y2=0

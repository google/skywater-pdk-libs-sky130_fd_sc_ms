* File: sky130_fd_sc_ms__o211ai_1.pex.spice
* Created: Wed Sep  2 12:20:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O211AI_1%A1 3 7 9 13 16
r28 15 16 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.505 $Y=1.465
+ $X2=0.515 $Y2=1.465
r29 12 15 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=0.27 $Y=1.465
+ $X2=0.505 $Y2=1.465
r30 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r31 9 13 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.27 $Y=1.665 $X2=0.27
+ $Y2=1.465
r32 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.3
+ $X2=0.515 $Y2=1.465
r33 5 7 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.515 $Y=1.3 $X2=0.515
+ $Y2=0.74
r34 1 15 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=1.465
r35 1 3 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O211AI_1%A2 3 7 9 10 11 12 19 25
r40 23 25 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.72 $Y=1.63
+ $X2=0.72 $Y2=1.665
r41 19 22 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.465 $X2=1
+ $Y2=1.63
r42 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=1.465 $X2=1
+ $Y2=1.3
r43 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.465
+ $X2=1 $Y2=1.465
r44 11 12 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=2.405
+ $X2=0.72 $Y2=2.775
r45 10 11 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=2.035
+ $X2=0.72 $Y2=2.405
r46 9 20 11.2739 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=0.72 $Y=1.465 $X2=1
+ $Y2=1.465
r47 9 23 2.35376 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.72 $Y=1.465
+ $X2=0.72 $Y2=1.63
r48 9 10 17.2866 $w=2.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.72 $Y=1.69
+ $X2=0.72 $Y2=2.035
r49 9 25 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.72 $Y=1.69 $X2=0.72
+ $Y2=1.665
r50 7 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.015 $Y=0.74
+ $X2=1.015 $Y2=1.3
r51 3 22 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.925 $Y=2.4
+ $X2=0.925 $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_MS__O211AI_1%B1 3 7 9 10 11 17 29
c40 3 0 1.83455e-19 $X=1.48 $Y=0.74
r41 21 29 0.250531 $w=2.28e-07 $l=5e-09 $layer=LI1_cond $X=1.68 $Y=1.3 $X2=1.68
+ $Y2=1.295
r42 17 20 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.57 $Y=1.465
+ $X2=1.57 $Y2=1.63
r43 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.57 $Y=1.465
+ $X2=1.57 $Y2=1.3
r44 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.57
+ $Y=1.465 $X2=1.57 $Y2=1.465
r45 11 18 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=1.68 $Y=1.465
+ $X2=1.57 $Y2=1.465
r46 11 21 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=1.465
+ $X2=1.68 $Y2=1.3
r47 11 29 2.00425 $w=2.28e-07 $l=4e-08 $layer=LI1_cond $X=1.68 $Y=1.255 $X2=1.68
+ $Y2=1.295
r48 10 11 16.5351 $w=2.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.68 $Y=0.925
+ $X2=1.68 $Y2=1.255
r49 9 10 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=0.555
+ $X2=1.68 $Y2=0.925
r50 7 20 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.645 $Y=2.4
+ $X2=1.645 $Y2=1.63
r51 3 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.48 $Y=0.74 $X2=1.48
+ $Y2=1.3
.ends

.subckt PM_SKY130_FD_SC_MS__O211AI_1%C1 3 6 8 11 13
r33 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.14 $Y=1.385
+ $X2=2.14 $Y2=1.55
r34 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.14 $Y=1.385
+ $X2=2.14 $Y2=1.22
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.385 $X2=2.14 $Y2=1.385
r36 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.14 $Y=1.295 $X2=2.14
+ $Y2=1.385
r37 6 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.145 $Y=2.4
+ $X2=2.145 $Y2=1.55
r38 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.05 $Y=0.74 $X2=2.05
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__O211AI_1%VPWR 1 2 7 9 15 18 19 20 30 31
r32 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r34 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r35 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r36 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r37 24 27 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r38 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 22 34 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r40 22 24 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 20 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 20 25 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 18 27 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.705 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.705 $Y=3.33
+ $X2=1.87 $Y2=3.33
r45 17 30 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=1.87 $Y2=3.33
r47 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.87 $Y=3.245
+ $X2=1.87 $Y2=3.33
r48 13 15 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=1.87 $Y=3.245
+ $X2=1.87 $Y2=2.305
r49 9 12 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=0.24 $Y=2.115 $X2=0.24
+ $Y2=2.815
r50 7 34 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r51 7 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245 $X2=0.24
+ $Y2=2.815
r52 2 15 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=1.735
+ $Y=1.84 $X2=1.87 $Y2=2.305
r53 1 12 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r54 1 9 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__O211AI_1%Y 1 2 3 12 16 17 20 25 26 27 28 37
r46 28 37 1.61576 $w=5.68e-07 $l=7.7e-08 $layer=LI1_cond $X=2.605 $Y=0.725
+ $X2=2.682 $Y2=0.725
r47 27 28 9.3378 $w=5.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.16 $Y=0.725
+ $X2=2.605 $Y2=0.725
r48 25 26 2.59952 $w=3.7e-07 $l=2.33666e-07 $layer=LI1_cond $X=2.682 $Y=1.8
+ $X2=2.487 $Y2=1.885
r49 24 37 7.81285 $w=1.75e-07 $l=2.85e-07 $layer=LI1_cond $X=2.682 $Y=1.01
+ $X2=2.682 $Y2=0.725
r50 24 25 50.0675 $w=1.73e-07 $l=7.9e-07 $layer=LI1_cond $X=2.682 $Y=1.01
+ $X2=2.682 $Y2=1.8
r51 20 22 17.5707 $w=5.63e-07 $l=8.3e-07 $layer=LI1_cond $X=2.487 $Y=1.985
+ $X2=2.487 $Y2=2.815
r52 18 26 2.59952 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.487 $Y=1.97
+ $X2=2.487 $Y2=1.885
r53 18 20 0.317543 $w=5.63e-07 $l=1.5e-08 $layer=LI1_cond $X=2.487 $Y=1.97
+ $X2=2.487 $Y2=1.985
r54 16 26 4.24538 $w=1.7e-07 $l=2.82e-07 $layer=LI1_cond $X=2.205 $Y=1.885
+ $X2=2.487 $Y2=1.885
r55 16 17 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.205 $Y=1.885
+ $X2=1.455 $Y2=1.885
r56 12 14 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.29 $Y=1.985
+ $X2=1.29 $Y2=2.815
r57 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.29 $Y=1.97
+ $X2=1.455 $Y2=1.885
r58 10 12 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.29 $Y=1.97
+ $X2=1.29 $Y2=1.985
r59 3 22 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.235
+ $Y=1.84 $X2=2.37 $Y2=2.815
r60 3 20 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.235
+ $Y=1.84 $X2=2.37 $Y2=1.985
r61 2 14 400 $w=1.7e-07 $l=1.10397e-06 $layer=licon1_PDIFF $count=1 $X=1.015
+ $Y=1.84 $X2=1.29 $Y2=2.815
r62 2 12 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=1.015
+ $Y=1.84 $X2=1.29 $Y2=1.985
r63 1 28 45.5 $w=1.7e-07 $l=5.67098e-07 $layer=licon1_NDIFF $count=4 $X=2.125
+ $Y=0.37 $X2=2.605 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_MS__O211AI_1%A_31_74# 1 2 9 11 12 15
c26 11 0 1.83455e-19 $X=1.145 $Y=1.045
r27 13 15 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=1.27 $Y=0.96
+ $X2=1.27 $Y2=0.515
r28 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.145 $Y=1.045
+ $X2=1.27 $Y2=0.96
r29 11 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.145 $Y=1.045
+ $X2=0.465 $Y2=1.045
r30 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.3 $Y=0.96
+ $X2=0.465 $Y2=1.045
r31 7 9 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.3 $Y=0.96 $X2=0.3
+ $Y2=0.515
r32 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.09
+ $Y=0.37 $X2=1.23 $Y2=0.515
r33 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.155
+ $Y=0.37 $X2=0.3 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O211AI_1%VGND 1 6 8 10 20 21 24
r28 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r29 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r30 18 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r31 17 20 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r32 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r33 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=0 $X2=0.8
+ $Y2=0
r34 15 17 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.965 $Y=0 $X2=1.2
+ $Y2=0
r35 13 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r36 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r37 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.635 $Y=0 $X2=0.8
+ $Y2=0
r38 10 12 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=0 $X2=0.24
+ $Y2=0
r39 8 21 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.64
+ $Y2=0
r40 8 18 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r41 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=0.085 $X2=0.8
+ $Y2=0
r42 4 6 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=0.8 $Y=0.085 $X2=0.8
+ $Y2=0.615
r43 1 6 182 $w=1.7e-07 $l=3.33879e-07 $layer=licon1_NDIFF $count=1 $X=0.59
+ $Y=0.37 $X2=0.8 $Y2=0.615
.ends


* File: sky130_fd_sc_ms__o41ai_1.spice
* Created: Fri Aug 28 18:05:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o41ai_1.pex.spice"
.subckt sky130_fd_sc_ms__o41ai_1  VNB VPB B1 A4 A3 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1009 N_A_157_74#_M1009_d N_B1_M1009_g N_Y_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.14615 AS=0.2109 PD=1.135 PS=2.05 NRD=18.648 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.3 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_A4_M1008_g N_A_157_74#_M1009_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.16095 AS=0.14615 PD=1.175 PS=1.135 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.8 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1003 N_A_157_74#_M1003_d N_A3_M1003_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.16095 PD=1.02 PS=1.175 NRD=0 NRS=13.776 M=1 R=4.93333
+ SA=75001.3 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g N_A_157_74#_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.8
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1000 N_A_157_74#_M1000_d N_A1_M1000_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.3
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_Y_M1006_d N_B1_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.56 PD=1.44 PS=3.24 NRD=7.8997 NRS=4.6886 M=1 R=6.22222
+ SA=90000.4 SB=90002.3 A=0.2016 P=2.6 MULT=1
MM1005 A_263_368# N_A4_M1005_g N_Y_M1006_d VPB PSHORT L=0.18 W=1.12 AD=0.1736
+ AS=0.1792 PD=1.43 PS=1.44 NRD=17.5724 NRS=0 M=1 R=6.22222 SA=90000.9
+ SB=90001.8 A=0.2016 P=2.6 MULT=1
MM1002 A_361_368# N_A3_M1002_g A_263_368# VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.1736 PD=1.51 PS=1.43 NRD=24.6053 NRS=17.5724 M=1 R=6.22222 SA=90001.4
+ SB=90001.3 A=0.2016 P=2.6 MULT=1
MM1001 A_475_368# N_A2_M1001_g A_361_368# VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.2184 PD=1.51 PS=1.51 NRD=24.6053 NRS=24.6053 M=1 R=6.22222 SA=90002
+ SB=90000.8 A=0.2016 P=2.6 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g A_475_368# VPB PSHORT L=0.18 W=1.12 AD=0.3136
+ AS=0.2184 PD=2.8 PS=1.51 NRD=0 NRS=24.6053 M=1 R=6.22222 SA=90002.5 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__o41ai_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__sedfxbp_2.pex.spice
* Created: Fri Aug 28 18:15:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SEDFXBP_2%D 3 7 11 12 17 18 20 22
c40 22 0 2.19166e-19 $X=0.54 $Y=1.99
c41 17 0 8.95046e-20 $X=0.54 $Y=1.145
r42 20 22 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.825
+ $X2=0.54 $Y2=1.99
r43 20 21 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.54
+ $Y=1.825 $X2=0.54 $Y2=1.825
r44 17 20 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=0.54 $Y=1.145
+ $X2=0.54 $Y2=1.825
r45 17 18 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.54
+ $Y=1.145 $X2=0.54 $Y2=1.145
r46 12 21 4.49734 $w=4.08e-07 $l=1.6e-07 $layer=LI1_cond $X=0.63 $Y=1.665
+ $X2=0.63 $Y2=1.825
r47 11 12 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.63 $Y=1.295
+ $X2=0.63 $Y2=1.665
r48 11 18 4.21625 $w=4.08e-07 $l=1.5e-07 $layer=LI1_cond $X=0.63 $Y=1.295
+ $X2=0.63 $Y2=1.145
r49 10 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=0.98
+ $X2=0.54 $Y2=1.145
r50 7 10 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.63 $Y=0.58 $X2=0.63
+ $Y2=0.98
r51 3 22 252.661 $w=1.8e-07 $l=6.5e-07 $layer=POLY_cond $X=0.585 $Y=2.64
+ $X2=0.585 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_2%A_183_290# 1 2 9 13 16 20 21 22 23 24 25
+ 28 32 34 38 39 41
c109 39 0 2.64211e-20 $X=2.47 $Y=1.68
c110 25 0 3.35759e-20 $X=1.335 $Y=2.035
c111 23 0 8.95046e-20 $X=1.335 $Y=1.195
r112 39 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.47 $Y=1.68
+ $X2=2.47 $Y2=1.515
r113 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.47
+ $Y=1.68 $X2=2.47 $Y2=1.68
r114 36 38 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=2.47 $Y=1.95
+ $X2=2.47 $Y2=1.68
r115 35 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=2.035
+ $X2=1.91 $Y2=2.035
r116 34 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.305 $Y=2.035
+ $X2=2.47 $Y2=1.95
r117 34 35 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.305 $Y=2.035
+ $X2=1.995 $Y2=2.035
r118 30 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.91 $Y=2.12
+ $X2=1.91 $Y2=2.035
r119 30 32 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.91 $Y=2.12
+ $X2=1.91 $Y2=2.51
r120 26 28 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.845 $Y=1.11
+ $X2=1.845 $Y2=0.775
r121 24 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.825 $Y=2.035
+ $X2=1.91 $Y2=2.035
r122 24 25 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.825 $Y=2.035
+ $X2=1.335 $Y2=2.035
r123 22 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.68 $Y=1.195
+ $X2=1.845 $Y2=1.11
r124 22 23 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.68 $Y=1.195
+ $X2=1.335 $Y2=1.195
r125 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.17
+ $Y=1.615 $X2=1.17 $Y2=1.615
r126 18 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.17 $Y=1.95
+ $X2=1.335 $Y2=2.035
r127 18 20 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.17 $Y=1.95
+ $X2=1.17 $Y2=1.615
r128 17 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.17 $Y=1.28
+ $X2=1.335 $Y2=1.195
r129 17 20 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.17 $Y=1.28
+ $X2=1.17 $Y2=1.615
r130 15 21 39.0632 $w=4.2e-07 $l=2.95e-07 $layer=POLY_cond $X=1.125 $Y=1.91
+ $X2=1.125 $Y2=1.615
r131 15 16 46.3397 $w=4.2e-07 $l=2.1e-07 $layer=POLY_cond $X=1.125 $Y=1.91
+ $X2=1.125 $Y2=2.12
r132 13 45 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.56 $Y=0.775
+ $X2=2.56 $Y2=1.515
r133 9 16 202.129 $w=1.8e-07 $l=5.2e-07 $layer=POLY_cond $X=1.005 $Y=2.64
+ $X2=1.005 $Y2=2.12
r134 2 32 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=1.765
+ $Y=2.31 $X2=1.91 $Y2=2.51
r135 1 28 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.7
+ $Y=0.565 $X2=1.845 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_2%DE 3 5 6 9 12 13 15 16 18 19 20 21 23 24
+ 28 31 33
c89 19 0 1.42059e-19 $X=2.725 $Y=2.16
r90 31 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.74 $Y=1.615
+ $X2=1.74 $Y2=1.78
r91 31 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.74 $Y=1.615
+ $X2=1.74 $Y2=1.45
r92 28 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.74
+ $Y=1.615 $X2=1.74 $Y2=1.615
r93 21 23 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.815 $Y=2.235
+ $X2=2.815 $Y2=2.63
r94 19 21 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.725 $Y=2.16
+ $X2=2.815 $Y2=2.235
r95 19 20 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.725 $Y=2.16
+ $X2=2.225 $Y2=2.16
r96 16 20 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.135 $Y=2.16
+ $X2=2.225 $Y2=2.16
r97 16 25 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=2.135 $Y=2.16
+ $X2=1.83 $Y2=2.16
r98 16 18 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.135 $Y=2.235
+ $X2=2.135 $Y2=2.63
r99 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.06 $Y=1.06 $X2=2.06
+ $Y2=0.775
r100 12 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.83 $Y=2.085
+ $X2=1.83 $Y2=2.16
r101 12 34 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=1.83 $Y=2.085
+ $X2=1.83 $Y2=1.78
r102 10 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.725 $Y=1.135
+ $X2=1.65 $Y2=1.135
r103 9 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.985 $Y=1.135
+ $X2=2.06 $Y2=1.06
r104 9 10 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.985 $Y=1.135
+ $X2=1.725 $Y2=1.135
r105 7 24 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.65 $Y=1.21
+ $X2=1.65 $Y2=1.135
r106 7 33 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.65 $Y=1.21
+ $X2=1.65 $Y2=1.45
r107 5 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.575 $Y=1.135
+ $X2=1.65 $Y2=1.135
r108 5 6 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.575 $Y=1.135
+ $X2=1.095 $Y2=1.135
r109 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.02 $Y=1.06
+ $X2=1.095 $Y2=1.135
r110 1 3 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.02 $Y=1.06 $X2=1.02
+ $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_2%A_575_87# 1 2 9 13 15 17 18 19 22 28 32 36
+ 40 42 45 47 49 53 56 57 60 61 65 68 69 75 82 83 86 91
c287 82 0 1.42059e-19 $X=3.04 $Y=1.68
c288 75 0 1.80649e-19 $X=15.12 $Y=1.665
c289 68 0 2.55325e-20 $X=14.975 $Y=1.665
c290 57 0 1.50731e-19 $X=15.995 $Y=2.405
c291 19 0 4.92549e-20 $X=13.345 $Y=0.94
c292 13 0 1.75904e-19 $X=3.205 $Y=2.63
r293 99 100 3.23498 $w=7.09e-07 $l=1.88e-07 $layer=LI1_cond $X=14.855 $Y=2.217
+ $X2=14.855 $Y2=2.405
r294 98 99 3.9921 $w=7.09e-07 $l=2.32e-07 $layer=LI1_cond $X=14.855 $Y=1.985
+ $X2=14.855 $Y2=2.217
r295 88 89 2.91239 $w=3.31e-07 $l=2e-08 $layer=POLY_cond $X=16.305 $Y=1.467
+ $X2=16.325 $Y2=1.467
r296 81 83 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.04 $Y=1.68
+ $X2=3.205 $Y2=1.68
r297 81 82 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.04
+ $Y=1.68 $X2=3.04 $Y2=1.68
r298 78 81 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.95 $Y=1.68 $X2=3.04
+ $Y2=1.68
r299 76 98 5.50635 $w=7.09e-07 $l=3.2e-07 $layer=LI1_cond $X=14.855 $Y=1.665
+ $X2=14.855 $Y2=1.985
r300 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=1.665
+ $X2=15.12 $Y2=1.665
r301 71 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.665
+ $X2=3.12 $Y2=1.665
r302 69 71 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=1.665
+ $X2=3.12 $Y2=1.665
r303 68 75 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.975 $Y=1.665
+ $X2=15.12 $Y2=1.665
r304 68 69 14.4925 $w=1.4e-07 $l=1.171e-05 $layer=MET1_cond $X=14.975 $Y=1.665
+ $X2=3.265 $Y2=1.665
r305 66 91 49.5106 $w=3.31e-07 $l=3.4e-07 $layer=POLY_cond $X=16.395 $Y=1.467
+ $X2=16.735 $Y2=1.467
r306 66 89 10.1934 $w=3.31e-07 $l=7e-08 $layer=POLY_cond $X=16.395 $Y=1.467
+ $X2=16.325 $Y2=1.467
r307 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=16.395
+ $Y=1.465 $X2=16.395 $Y2=1.465
r308 62 65 10.4924 $w=3.33e-07 $l=3.05e-07 $layer=LI1_cond $X=16.09 $Y=1.467
+ $X2=16.395 $Y2=1.467
r309 59 62 4.05585 $w=1.9e-07 $l=1.68e-07 $layer=LI1_cond $X=16.09 $Y=1.635
+ $X2=16.09 $Y2=1.467
r310 59 60 39.9856 $w=1.88e-07 $l=6.85e-07 $layer=LI1_cond $X=16.09 $Y=1.635
+ $X2=16.09 $Y2=2.32
r311 58 100 9.40575 $w=1.7e-07 $l=3.8e-07 $layer=LI1_cond $X=15.235 $Y=2.405
+ $X2=14.855 $Y2=2.405
r312 57 60 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=15.995 $Y=2.405
+ $X2=16.09 $Y2=2.32
r313 57 58 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=15.995 $Y=2.405
+ $X2=15.235 $Y2=2.405
r314 56 76 10.2197 $w=7.09e-07 $l=1.5906e-07 $layer=LI1_cond $X=14.75 $Y=1.55
+ $X2=14.855 $Y2=1.665
r315 56 61 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=14.75 $Y=1.55
+ $X2=14.75 $Y2=1.13
r316 51 61 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=14.67 $Y=0.965
+ $X2=14.67 $Y2=1.13
r317 51 53 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=14.67 $Y=0.965
+ $X2=14.67 $Y2=0.515
r318 47 100 4.4124 $w=7.09e-07 $l=2.38747e-07 $layer=LI1_cond $X=14.655 $Y=2.49
+ $X2=14.855 $Y2=2.405
r319 47 49 10.404 $w=3.58e-07 $l=3.25e-07 $layer=LI1_cond $X=14.655 $Y=2.49
+ $X2=14.655 $Y2=2.815
r320 45 87 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.75 $Y=2.215
+ $X2=13.75 $Y2=2.38
r321 45 86 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.75 $Y=2.215
+ $X2=13.75 $Y2=2.05
r322 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.75
+ $Y=2.215 $X2=13.75 $Y2=2.215
r323 42 99 5.32966 $w=3.25e-07 $l=3.8e-07 $layer=LI1_cond $X=14.475 $Y=2.217
+ $X2=14.855 $Y2=2.217
r324 42 44 25.7083 $w=3.23e-07 $l=7.25e-07 $layer=LI1_cond $X=14.475 $Y=2.217
+ $X2=13.75 $Y2=2.217
r325 38 91 5.82477 $w=3.31e-07 $l=4e-08 $layer=POLY_cond $X=16.775 $Y=1.467
+ $X2=16.735 $Y2=1.467
r326 38 40 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=16.775 $Y=1.63
+ $X2=16.775 $Y2=2.4
r327 34 91 21.295 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=16.735 $Y=1.3
+ $X2=16.735 $Y2=1.467
r328 34 36 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=16.735 $Y=1.3
+ $X2=16.735 $Y2=0.74
r329 30 89 17.0024 $w=1.8e-07 $l=1.68e-07 $layer=POLY_cond $X=16.325 $Y=1.635
+ $X2=16.325 $Y2=1.467
r330 30 32 297.363 $w=1.8e-07 $l=7.65e-07 $layer=POLY_cond $X=16.325 $Y=1.635
+ $X2=16.325 $Y2=2.4
r331 26 88 21.295 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=16.305 $Y=1.3
+ $X2=16.305 $Y2=1.467
r332 26 28 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=16.305 $Y=1.3
+ $X2=16.305 $Y2=0.74
r333 24 86 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=13.84 $Y=1.015
+ $X2=13.84 $Y2=2.05
r334 22 87 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=13.705 $Y=2.75
+ $X2=13.705 $Y2=2.38
r335 18 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.765 $Y=0.94
+ $X2=13.84 $Y2=1.015
r336 18 19 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=13.765 $Y=0.94
+ $X2=13.345 $Y2=0.94
r337 15 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.27 $Y=0.865
+ $X2=13.345 $Y2=0.94
r338 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=13.27 $Y=0.865
+ $X2=13.27 $Y2=0.58
r339 11 83 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=1.845
+ $X2=3.205 $Y2=1.68
r340 11 13 305.137 $w=1.8e-07 $l=7.85e-07 $layer=POLY_cond $X=3.205 $Y=1.845
+ $X2=3.205 $Y2=2.63
r341 7 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.515
+ $X2=2.95 $Y2=1.68
r342 7 9 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.95 $Y=1.515
+ $X2=2.95 $Y2=0.775
r343 2 98 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=14.505
+ $Y=1.84 $X2=14.64 $Y2=1.985
r344 2 49 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=14.505
+ $Y=1.84 $X2=14.64 $Y2=2.815
r345 1 53 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.53
+ $Y=0.37 $X2=14.67 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_2%A_661_87# 1 2 7 9 10 11 14 18 20 21 24 27
+ 30 32 36 37 40 45 48 49
c108 48 0 1.27569e-19 $X=5.97 $Y=1.58
r109 48 51 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=5.97 $Y=1.58
+ $X2=5.97 $Y2=1.765
r110 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.97
+ $Y=1.58 $X2=5.97 $Y2=1.58
r111 42 45 5.37015 $w=4.88e-07 $l=2.2e-07 $layer=LI1_cond $X=4.22 $Y=2.49
+ $X2=4.44 $Y2=2.49
r112 39 41 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.18 $Y=1.89
+ $X2=4.18 $Y2=2.055
r113 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.18
+ $Y=1.89 $X2=4.18 $Y2=1.89
r114 37 39 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=4.18 $Y=1.765
+ $X2=4.18 $Y2=1.89
r115 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.18
+ $Y=0.53 $X2=4.18 $Y2=0.53
r116 33 37 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.305 $Y=1.765
+ $X2=4.18 $Y2=1.765
r117 32 51 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.805 $Y=1.765
+ $X2=5.97 $Y2=1.765
r118 32 33 97.861 $w=1.68e-07 $l=1.5e-06 $layer=LI1_cond $X=5.805 $Y=1.765
+ $X2=4.305 $Y2=1.765
r119 28 35 3.15958 $w=4.05e-07 $l=1.75e-07 $layer=LI1_cond $X=4.305 $Y=0.807
+ $X2=4.18 $Y2=0.687
r120 28 30 9.10572 $w=4.03e-07 $l=3.2e-07 $layer=LI1_cond $X=4.305 $Y=0.807
+ $X2=4.625 $Y2=0.807
r121 27 42 7.03003 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=4.22 $Y=2.245
+ $X2=4.22 $Y2=2.49
r122 27 41 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.22 $Y=2.245
+ $X2=4.22 $Y2=2.055
r123 25 40 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=4.18 $Y=1.21
+ $X2=4.18 $Y2=1.89
r124 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.18
+ $Y=1.21 $X2=4.18 $Y2=1.21
r125 22 37 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=4.18 $Y=1.68
+ $X2=4.18 $Y2=1.765
r126 22 24 21.6659 $w=2.48e-07 $l=4.7e-07 $layer=LI1_cond $X=4.18 $Y=1.68
+ $X2=4.18 $Y2=1.21
r127 21 35 4.16548 $w=2.5e-07 $l=3.23e-07 $layer=LI1_cond $X=4.18 $Y=1.01
+ $X2=4.18 $Y2=0.687
r128 21 24 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=4.18 $Y=1.01 $X2=4.18
+ $Y2=1.21
r129 19 49 36.0236 $w=4.4e-07 $l=2.85e-07 $layer=POLY_cond $X=5.915 $Y=1.865
+ $X2=5.915 $Y2=1.58
r130 19 20 47.7869 $w=4.4e-07 $l=2.2e-07 $layer=POLY_cond $X=5.915 $Y=1.865
+ $X2=5.915 $Y2=2.085
r131 18 25 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.18 $Y=1.135
+ $X2=4.18 $Y2=1.21
r132 16 36 92.6765 $w=3.3e-07 $l=5.3e-07 $layer=POLY_cond $X=4.18 $Y=1.06
+ $X2=4.18 $Y2=0.53
r133 16 18 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.18 $Y=1.06
+ $X2=4.18 $Y2=1.135
r134 14 20 194.355 $w=1.8e-07 $l=5e-07 $layer=POLY_cond $X=5.785 $Y=2.585
+ $X2=5.785 $Y2=2.085
r135 10 18 16.9349 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.015 $Y=1.135
+ $X2=4.18 $Y2=1.135
r136 10 11 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.015 $Y=1.135
+ $X2=3.455 $Y2=1.135
r137 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.38 $Y=1.06
+ $X2=3.455 $Y2=1.135
r138 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.38 $Y=1.06 $X2=3.38
+ $Y2=0.775
r139 2 45 600 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_PDIFF $count=1 $X=4.295
+ $Y=2.265 $X2=4.44 $Y2=2.49
r140 1 30 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=4.48
+ $Y=0.625 $X2=4.625 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_2%SCD 3 7 9 12
r41 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.29 $Y=1.345
+ $X2=5.29 $Y2=1.51
r42 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.29 $Y=1.345
+ $X2=5.29 $Y2=1.18
r43 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.29
+ $Y=1.345 $X2=5.29 $Y2=1.345
r44 9 13 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=5.52 $Y=1.345
+ $X2=5.29 $Y2=1.345
r45 7 14 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=5.38 $Y=0.835
+ $X2=5.38 $Y2=1.18
r46 3 15 417.863 $w=1.8e-07 $l=1.075e-06 $layer=POLY_cond $X=5.365 $Y=2.585
+ $X2=5.365 $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_2%SCE 1 3 4 5 9 13 14 15 18 20 23 24
c75 18 0 1.27569e-19 $X=5.77 $Y=0.835
c76 1 0 3.25608e-19 $X=3.655 $Y=3.025
r77 23 26 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.75 $Y=1.345
+ $X2=4.75 $Y2=1.51
r78 23 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.75 $Y=1.345
+ $X2=4.75 $Y2=1.18
r79 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.75
+ $Y=1.345 $X2=4.75 $Y2=1.345
r80 20 24 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.56 $Y=1.345
+ $X2=4.75 $Y2=1.345
r81 16 18 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.77 $Y=0.255
+ $X2=5.77 $Y2=0.835
r82 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.695 $Y=0.18
+ $X2=5.77 $Y2=0.255
r83 14 15 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=5.695 $Y=0.18
+ $X2=4.915 $Y2=0.18
r84 13 25 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=4.84 $Y=0.835
+ $X2=4.84 $Y2=1.18
r85 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.84 $Y=0.255
+ $X2=4.915 $Y2=0.18
r86 10 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.84 $Y=0.255
+ $X2=4.84 $Y2=0.835
r87 9 26 417.863 $w=1.8e-07 $l=1.075e-06 $layer=POLY_cond $X=4.675 $Y=2.585
+ $X2=4.675 $Y2=1.51
r88 7 9 171.032 $w=1.8e-07 $l=4.4e-07 $layer=POLY_cond $X=4.675 $Y=3.025
+ $X2=4.675 $Y2=2.585
r89 4 7 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.585 $Y=3.1
+ $X2=4.675 $Y2=3.025
r90 4 5 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.585 $Y=3.1 $X2=3.745
+ $Y2=3.1
r91 1 5 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.655 $Y=3.025
+ $X2=3.745 $Y2=3.1
r92 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.655 $Y=3.025
+ $X2=3.655 $Y2=2.63
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_2%CLK 3 7 8 11 13
r39 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.87 $Y=1.385
+ $X2=6.87 $Y2=1.55
r40 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.87 $Y=1.385
+ $X2=6.87 $Y2=1.22
r41 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.87
+ $Y=1.385 $X2=6.87 $Y2=1.385
r42 8 12 3.05058 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=6.875 $Y=1.295
+ $X2=6.875 $Y2=1.385
r43 7 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.865 $Y=0.74
+ $X2=6.865 $Y2=1.22
r44 3 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=6.795 $Y=2.4
+ $X2=6.795 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_2%A_1586_74# 1 2 9 11 13 16 20 24 26 27 28
+ 34 37 40 41 43 46 47 48 50 51 52 53 55 58 60 61 64 66 67 70 74 84
c232 84 0 5.95143e-20 $X=12.37 $Y=1.635
c233 70 0 9.34686e-20 $X=13.36 $Y=1.215
c234 64 0 1.96976e-19 $X=8.89 $Y=2.14
c235 60 0 1.82067e-19 $X=8.89 $Y=1.98
c236 37 0 1.94394e-19 $X=9.65 $Y=0.85
c237 20 0 2.68352e-19 $X=13.285 $Y=2.75
r238 74 88 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.36 $Y=1.39
+ $X2=13.36 $Y2=1.555
r239 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.36
+ $Y=1.39 $X2=13.36 $Y2=1.39
r240 70 73 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=13.36 $Y=1.215
+ $X2=13.36 $Y2=1.39
r241 68 69 15.5982 $w=2.19e-07 $l=2.8e-07 $layer=LI1_cond $X=12.23 $Y=0.935
+ $X2=12.23 $Y2=1.215
r242 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.89
+ $Y=2.14 $X2=8.89 $Y2=2.14
r243 60 63 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=8.89 $Y=1.98
+ $X2=8.89 $Y2=2.14
r244 60 61 8.28756 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=8.89 $Y=1.98
+ $X2=8.89 $Y2=1.82
r245 59 69 2.22295 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=12.38 $Y=1.215
+ $X2=12.23 $Y2=1.215
r246 58 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.195 $Y=1.215
+ $X2=13.36 $Y2=1.215
r247 58 59 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=13.195 $Y=1.215
+ $X2=12.38 $Y2=1.215
r248 56 84 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=12.26 $Y=1.635
+ $X2=12.37 $Y2=1.635
r249 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.26
+ $Y=1.635 $X2=12.26 $Y2=1.635
r250 53 69 4.36852 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.23 $Y=1.3 $X2=12.23
+ $Y2=1.215
r251 53 55 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=12.23 $Y=1.3
+ $X2=12.23 $Y2=1.635
r252 51 68 2.22295 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=12.08 $Y=0.935
+ $X2=12.23 $Y2=0.935
r253 51 52 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=12.08 $Y=0.935
+ $X2=11.54 $Y2=0.935
r254 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.455 $Y=0.85
+ $X2=11.54 $Y2=0.935
r255 49 50 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=11.455 $Y=0.425
+ $X2=11.455 $Y2=0.85
r256 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.37 $Y=0.34
+ $X2=11.455 $Y2=0.425
r257 47 48 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=11.37 $Y=0.34
+ $X2=10.86 $Y2=0.34
r258 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.775 $Y=0.425
+ $X2=10.86 $Y2=0.34
r259 45 46 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=10.775 $Y=0.425
+ $X2=10.775 $Y2=0.85
r260 44 67 2.45049 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=9.855 $Y=0.935
+ $X2=9.71 $Y2=0.935
r261 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.69 $Y=0.935
+ $X2=10.775 $Y2=0.85
r262 43 44 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=10.69 $Y=0.935
+ $X2=9.855 $Y2=0.935
r263 41 78 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.69 $Y=1.18
+ $X2=9.525 $Y2=1.18
r264 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.69
+ $Y=1.18 $X2=9.69 $Y2=1.18
r265 38 67 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.71 $Y=1.02
+ $X2=9.71 $Y2=0.935
r266 38 40 6.35831 $w=2.88e-07 $l=1.6e-07 $layer=LI1_cond $X=9.71 $Y=1.02
+ $X2=9.71 $Y2=1.18
r267 37 67 3.98977 $w=2.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=9.65 $Y=0.85
+ $X2=9.71 $Y2=0.935
r268 36 37 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=9.65 $Y=0.425
+ $X2=9.65 $Y2=0.85
r269 35 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.055 $Y=0.34
+ $X2=8.97 $Y2=0.34
r270 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.565 $Y=0.34
+ $X2=9.65 $Y2=0.425
r271 34 35 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.565 $Y=0.34
+ $X2=9.055 $Y2=0.34
r272 32 66 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.97 $Y=0.425
+ $X2=8.97 $Y2=0.34
r273 32 61 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=8.97 $Y=0.425
+ $X2=8.97 $Y2=1.82
r274 28 60 0.903439 $w=3.2e-07 $l=1.65e-07 $layer=LI1_cond $X=8.725 $Y=1.98
+ $X2=8.89 $Y2=1.98
r275 28 30 11.3444 $w=3.18e-07 $l=3.15e-07 $layer=LI1_cond $X=8.725 $Y=1.98
+ $X2=8.41 $Y2=1.98
r276 26 66 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.885 $Y=0.34
+ $X2=8.97 $Y2=0.34
r277 26 27 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=8.885 $Y=0.34
+ $X2=8.235 $Y2=0.34
r278 22 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.07 $Y=0.425
+ $X2=8.235 $Y2=0.34
r279 22 24 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=8.07 $Y=0.425
+ $X2=8.07 $Y2=0.515
r280 20 88 464.508 $w=1.8e-07 $l=1.195e-06 $layer=POLY_cond $X=13.285 $Y=2.75
+ $X2=13.285 $Y2=1.555
r281 14 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.37 $Y=1.47
+ $X2=12.37 $Y2=1.635
r282 14 16 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=12.37 $Y=1.47
+ $X2=12.37 $Y2=0.69
r283 11 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.525 $Y=1.015
+ $X2=9.525 $Y2=1.18
r284 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.525 $Y=1.015
+ $X2=9.525 $Y2=0.695
r285 7 64 57.4258 $w=2.56e-07 $l=3.78616e-07 $layer=POLY_cond $X=9.195 $Y=2.305
+ $X2=8.89 $Y2=2.14
r286 7 9 172.976 $w=1.8e-07 $l=4.45e-07 $layer=POLY_cond $X=9.195 $Y=2.305
+ $X2=9.195 $Y2=2.75
r287 2 30 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=8.275
+ $Y=1.84 $X2=8.41 $Y2=2.02
r288 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.93
+ $Y=0.37 $X2=8.07 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_2%A_1377_368# 1 2 11 13 15 17 18 22 24 30 34
+ 38 40 41 42 48 51 53 57 58 59 63 64 69 70 75 77
c191 77 0 1.82067e-19 $X=9.69 $Y=2.03
c192 70 0 9.34686e-20 $X=12.82 $Y=1.635
c193 69 0 1.09438e-19 $X=12.82 $Y=1.635
c194 63 0 1.96976e-19 $X=9.69 $Y=2.195
c195 48 0 1.58914e-19 $X=12.55 $Y=2.475
c196 22 0 1.94394e-19 $X=8.845 $Y=0.695
r197 70 81 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.82 $Y=1.635
+ $X2=12.82 $Y2=1.8
r198 70 80 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.82 $Y=1.635
+ $X2=12.82 $Y2=1.47
r199 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.82
+ $Y=1.635 $X2=12.82 $Y2=1.635
r200 66 69 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=12.635 $Y=1.635
+ $X2=12.82 $Y2=1.635
r201 64 78 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.69 $Y=2.195
+ $X2=9.69 $Y2=2.36
r202 64 77 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.69 $Y=2.195
+ $X2=9.69 $Y2=2.03
r203 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.69
+ $Y=2.195 $X2=9.69 $Y2=2.195
r204 57 60 9.0362 $w=4.38e-07 $l=3.45e-07 $layer=LI1_cond $X=7.435 $Y=1.635
+ $X2=7.435 $Y2=1.98
r205 57 59 8.83531 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=7.435 $Y=1.635
+ $X2=7.435 $Y2=1.47
r206 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.49
+ $Y=1.635 $X2=7.49 $Y2=1.635
r207 55 59 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=7.3 $Y=1.01 $X2=7.3
+ $Y2=1.47
r208 53 55 17.7356 $w=4.68e-07 $l=4.95e-07 $layer=LI1_cond $X=7.15 $Y=0.515
+ $X2=7.15 $Y2=1.01
r209 50 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.635 $Y=1.8
+ $X2=12.635 $Y2=1.635
r210 50 51 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=12.635 $Y=1.8
+ $X2=12.635 $Y2=2.39
r211 49 63 11.8611 $w=2.88e-07 $l=3.58887e-07 $layer=LI1_cond $X=9.925 $Y=2.475
+ $X2=9.745 $Y2=2.195
r212 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.55 $Y=2.475
+ $X2=12.635 $Y2=2.39
r213 48 49 171.257 $w=1.68e-07 $l=2.625e-06 $layer=LI1_cond $X=12.55 $Y=2.475
+ $X2=9.925 $Y2=2.475
r214 42 60 2.60351 $w=3.2e-07 $l=2.2e-07 $layer=LI1_cond $X=7.215 $Y=1.98
+ $X2=7.435 $Y2=1.98
r215 42 44 7.0227 $w=3.18e-07 $l=1.95e-07 $layer=LI1_cond $X=7.215 $Y=1.98
+ $X2=7.02 $Y2=1.98
r216 38 80 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=12.88 $Y=0.58
+ $X2=12.88 $Y2=1.47
r217 34 81 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=12.75 $Y=2.46
+ $X2=12.75 $Y2=1.8
r218 30 78 151.597 $w=1.8e-07 $l=3.9e-07 $layer=POLY_cond $X=9.645 $Y=2.75
+ $X2=9.645 $Y2=2.36
r219 26 77 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=9.6 $Y=1.735
+ $X2=9.6 $Y2=2.03
r220 25 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.92 $Y=1.66
+ $X2=8.845 $Y2=1.66
r221 24 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.525 $Y=1.66
+ $X2=9.6 $Y2=1.735
r222 24 25 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=9.525 $Y=1.66
+ $X2=8.92 $Y2=1.66
r223 20 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.845 $Y=1.585
+ $X2=8.845 $Y2=1.66
r224 20 22 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=8.845 $Y=1.585
+ $X2=8.845 $Y2=0.695
r225 19 40 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.275 $Y=1.66
+ $X2=8.185 $Y2=1.66
r226 18 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.77 $Y=1.66
+ $X2=8.845 $Y2=1.66
r227 18 19 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=8.77 $Y=1.66
+ $X2=8.275 $Y2=1.66
r228 15 40 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=8.185 $Y=1.735
+ $X2=8.185 $Y2=1.66
r229 15 17 178.072 $w=1.8e-07 $l=6.65e-07 $layer=POLY_cond $X=8.185 $Y=1.735
+ $X2=8.185 $Y2=2.4
r230 13 40 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.095 $Y=1.66
+ $X2=8.185 $Y2=1.66
r231 13 75 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.095 $Y=1.66
+ $X2=7.93 $Y2=1.66
r232 9 75 28.1815 $w=2.65e-07 $l=7.5e-08 $layer=POLY_cond $X=7.855 $Y=1.602
+ $X2=7.93 $Y2=1.602
r233 9 58 82.6235 $w=2.65e-07 $l=3.65e-07 $layer=POLY_cond $X=7.855 $Y=1.602
+ $X2=7.49 $Y2=1.602
r234 9 11 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=7.855 $Y=1.47
+ $X2=7.855 $Y2=0.74
r235 2 44 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=6.885
+ $Y=1.84 $X2=7.02 $Y2=2.02
r236 1 53 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.94
+ $Y=0.37 $X2=7.08 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_2%A_2013_71# 1 2 9 13 17 19 21 23 24 26 32
+ 35 36 38 39 41 45
c113 45 0 2.55325e-20 $X=10.23 $Y=1.355
c114 41 0 1.43495e-19 $X=10.23 $Y=1.275
c115 38 0 5.95143e-20 $X=11.72 $Y=1.355
r116 47 48 9.1748 $w=2.46e-07 $l=1.85e-07 $layer=LI1_cond $X=11.115 $Y=1.355
+ $X2=11.3 $Y2=1.355
r117 45 51 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.23 $Y=1.355
+ $X2=10.23 $Y2=1.52
r118 45 50 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.23 $Y=1.355
+ $X2=10.23 $Y2=1.19
r119 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.23
+ $Y=1.355 $X2=10.23 $Y2=1.355
r120 41 44 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=10.23 $Y=1.275
+ $X2=10.23 $Y2=1.355
r121 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.72
+ $Y=1.355 $X2=11.72 $Y2=1.355
r122 36 48 3.95924 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.385 $Y=1.355
+ $X2=11.3 $Y2=1.355
r123 36 38 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=11.385 $Y=1.355
+ $X2=11.72 $Y2=1.355
r124 34 48 2.90119 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.3 $Y=1.52
+ $X2=11.3 $Y2=1.355
r125 34 35 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=11.3 $Y=1.52
+ $X2=11.3 $Y2=2.05
r126 30 47 2.90119 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.115 $Y=1.19
+ $X2=11.115 $Y2=1.355
r127 30 32 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=11.115 $Y=1.19
+ $X2=11.115 $Y2=0.805
r128 26 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.215 $Y=2.135
+ $X2=11.3 $Y2=2.05
r129 26 28 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=11.215 $Y=2.135
+ $X2=10.925 $Y2=2.135
r130 25 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.395 $Y=1.275
+ $X2=10.23 $Y2=1.275
r131 24 47 5.39088 $w=2.46e-07 $l=1.18427e-07 $layer=LI1_cond $X=11.03 $Y=1.275
+ $X2=11.115 $Y2=1.355
r132 24 25 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=11.03 $Y=1.275
+ $X2=10.395 $Y2=1.275
r133 21 23 134.96 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=12.01 $Y=1.11
+ $X2=12.01 $Y2=0.69
r134 17 21 37.9597 $w=2.73e-07 $l=3.7229e-07 $layer=POLY_cond $X=11.795 $Y=1.39
+ $X2=12.01 $Y2=1.11
r135 17 39 13.2418 $w=2.73e-07 $l=7.5e-08 $layer=POLY_cond $X=11.795 $Y=1.39
+ $X2=11.72 $Y2=1.39
r136 17 19 365.387 $w=1.8e-07 $l=9.4e-07 $layer=POLY_cond $X=11.795 $Y=1.52
+ $X2=11.795 $Y2=2.46
r137 13 51 478.113 $w=1.8e-07 $l=1.23e-06 $layer=POLY_cond $X=10.155 $Y=2.75
+ $X2=10.155 $Y2=1.52
r138 9 50 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.14 $Y=0.695
+ $X2=10.14 $Y2=1.19
r139 2 28 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.79
+ $Y=1.99 $X2=10.925 $Y2=2.135
r140 1 32 182 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_NDIFF $count=1 $X=10.975
+ $Y=0.37 $X2=11.115 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_2%A_1784_97# 1 2 9 13 17 21 23 25 26 29 37
c88 37 0 1.43495e-19 $X=10.9 $Y=1.665
r89 30 37 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=10.775 $Y=1.665
+ $X2=10.9 $Y2=1.665
r90 30 34 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=10.775 $Y=1.665
+ $X2=10.7 $Y2=1.665
r91 29 32 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=10.775 $Y=1.665
+ $X2=10.775 $Y2=1.775
r92 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.775
+ $Y=1.665 $X2=10.775 $Y2=1.665
r93 25 26 10.4318 $w=3.58e-07 $l=2.25e-07 $layer=LI1_cond $X=9.405 $Y=2.755
+ $X2=9.405 $Y2=2.53
r94 22 23 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.395 $Y=1.775
+ $X2=9.31 $Y2=1.775
r95 21 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.61 $Y=1.775
+ $X2=10.775 $Y2=1.775
r96 21 22 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=10.61 $Y=1.775
+ $X2=9.395 $Y2=1.775
r97 19 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.31 $Y=1.86 $X2=9.31
+ $Y2=1.775
r98 19 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.31 $Y=1.86
+ $X2=9.31 $Y2=2.53
r99 15 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.31 $Y=1.69 $X2=9.31
+ $Y2=1.775
r100 15 17 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=9.31 $Y=1.69
+ $X2=9.31 $Y2=0.76
r101 11 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.9 $Y=1.5
+ $X2=10.9 $Y2=1.665
r102 11 13 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=10.9 $Y=1.5 $X2=10.9
+ $Y2=0.69
r103 7 34 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.7 $Y=1.83
+ $X2=10.7 $Y2=1.665
r104 7 9 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=10.7 $Y=1.83 $X2=10.7
+ $Y2=2.41
r105 2 25 600 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=9.285
+ $Y=2.54 $X2=9.42 $Y2=2.755
r106 1 17 182 $w=1.7e-07 $l=5.09264e-07 $layer=licon1_NDIFF $count=1 $X=8.92
+ $Y=0.485 $X2=9.31 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_2%A_2489_74# 1 2 9 13 15 19 23 27 31 35 37
+ 39 41 44 45 46 48 49 51 52 59
c152 51 0 1.80649e-19 $X=14.33 $Y=1.465
c153 46 0 4.92549e-20 $X=13.325 $Y=1.8
c154 37 0 1.45871e-19 $X=12.585 $Y=0.77
c155 15 0 1.50731e-19 $X=15.335 $Y=1.465
r156 57 59 6.89045 $w=4.58e-07 $l=2.65e-07 $layer=LI1_cond $X=12.975 $Y=2.75
+ $X2=13.24 $Y2=2.75
r157 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.33
+ $Y=1.465 $X2=14.33 $Y2=1.465
r158 49 62 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=13.78 $Y=1.465
+ $X2=13.78 $Y2=1.8
r159 49 51 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=13.865 $Y=1.465
+ $X2=14.33 $Y2=1.465
r160 48 49 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=13.78 $Y=1.3
+ $X2=13.78 $Y2=1.465
r161 47 48 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=13.78 $Y=0.94
+ $X2=13.78 $Y2=1.3
r162 45 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.695 $Y=1.8
+ $X2=13.78 $Y2=1.8
r163 45 46 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=13.695 $Y=1.8
+ $X2=13.325 $Y2=1.8
r164 44 59 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=13.24 $Y=2.52
+ $X2=13.24 $Y2=2.75
r165 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.24 $Y=1.885
+ $X2=13.325 $Y2=1.8
r166 43 44 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=13.24 $Y=1.885
+ $X2=13.24 $Y2=2.52
r167 42 55 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.75 $Y=0.855
+ $X2=12.585 $Y2=0.855
r168 41 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.695 $Y=0.855
+ $X2=13.78 $Y2=0.94
r169 41 42 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=13.695 $Y=0.855
+ $X2=12.75 $Y2=0.855
r170 37 55 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.585 $Y=0.77
+ $X2=12.585 $Y2=0.855
r171 37 39 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=12.585 $Y=0.77
+ $X2=12.585 $Y2=0.515
r172 34 35 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=15.445 $Y=1.465
+ $X2=15.875 $Y2=1.465
r173 33 34 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=15.425 $Y=1.465
+ $X2=15.445 $Y2=1.465
r174 29 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.875 $Y=1.3
+ $X2=15.875 $Y2=1.465
r175 29 31 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=15.875 $Y=1.3
+ $X2=15.875 $Y2=0.74
r176 25 35 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=15.875 $Y=1.63
+ $X2=15.875 $Y2=1.465
r177 25 27 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=15.875 $Y=1.63
+ $X2=15.875 $Y2=2.4
r178 21 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.445 $Y=1.3
+ $X2=15.445 $Y2=1.465
r179 21 23 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=15.445 $Y=1.3
+ $X2=15.445 $Y2=0.74
r180 17 33 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=15.425 $Y=1.63
+ $X2=15.425 $Y2=1.465
r181 17 19 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=15.425 $Y=1.63
+ $X2=15.425 $Y2=2.4
r182 16 52 3.90195 $w=3.3e-07 $l=1.83e-07 $layer=POLY_cond $X=14.53 $Y=1.465
+ $X2=14.347 $Y2=1.465
r183 15 33 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=15.335 $Y=1.465
+ $X2=15.425 $Y2=1.465
r184 15 16 140.763 $w=3.3e-07 $l=8.05e-07 $layer=POLY_cond $X=15.335 $Y=1.465
+ $X2=14.53 $Y2=1.465
r185 11 52 34.7346 $w=1.65e-07 $l=2.12238e-07 $layer=POLY_cond $X=14.455 $Y=1.3
+ $X2=14.347 $Y2=1.465
r186 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=14.455 $Y=1.3
+ $X2=14.455 $Y2=0.74
r187 7 52 34.7346 $w=1.65e-07 $l=1.96074e-07 $layer=POLY_cond $X=14.415 $Y=1.63
+ $X2=14.347 $Y2=1.465
r188 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=14.415 $Y=1.63
+ $X2=14.415 $Y2=2.4
r189 2 57 600 $w=1.7e-07 $l=8.54839e-07 $layer=licon1_PDIFF $count=1 $X=12.84
+ $Y=1.96 $X2=12.975 $Y2=2.75
r190 1 55 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=12.445
+ $Y=0.37 $X2=12.585 $Y2=0.855
r191 1 39 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=12.445
+ $Y=0.37 $X2=12.585 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_2%A_32_74# 1 2 3 4 14 17 19 22 23 24 26 27
+ 28 31 36 40 42 45 48
c115 48 0 3.25608e-19 $X=3.43 $Y=2.455
c116 28 0 2.64211e-20 $X=2.335 $Y=2.375
c117 19 0 1.8559e-19 $X=1.485 $Y=2.375
r118 37 40 9.10802 $w=3.08e-07 $l=2.45e-07 $layer=LI1_cond $X=0.17 $Y=0.575
+ $X2=0.415 $Y2=0.575
r119 36 48 4.06715 $w=2.25e-07 $l=1.09087e-07 $layer=LI1_cond $X=3.46 $Y=2.29
+ $X2=3.405 $Y2=2.375
r120 35 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=1.345
+ $X2=3.46 $Y2=1.26
r121 35 36 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=3.46 $Y=1.345
+ $X2=3.46 $Y2=2.29
r122 29 45 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.165 $Y=1.26
+ $X2=3.46 $Y2=1.26
r123 29 31 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=3.165 $Y=1.175
+ $X2=3.165 $Y2=0.775
r124 27 48 2.36881 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.265 $Y=2.375
+ $X2=3.405 $Y2=2.375
r125 27 28 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.265 $Y=2.375
+ $X2=2.335 $Y2=2.375
r126 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.25 $Y=2.46
+ $X2=2.335 $Y2=2.375
r127 25 26 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.25 $Y=2.46
+ $X2=2.25 $Y2=2.905
r128 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.165 $Y=2.99
+ $X2=2.25 $Y2=2.905
r129 23 24 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.165 $Y=2.99
+ $X2=1.655 $Y2=2.99
r130 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.57 $Y=2.905
+ $X2=1.655 $Y2=2.99
r131 21 22 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.57 $Y=2.46
+ $X2=1.57 $Y2=2.905
r132 20 42 3.51065 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.525 $Y=2.375
+ $X2=0.305 $Y2=2.375
r133 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.485 $Y=2.375
+ $X2=1.57 $Y2=2.46
r134 19 20 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.485 $Y=2.375
+ $X2=0.525 $Y2=2.375
r135 15 42 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.305 $Y=2.46
+ $X2=0.305 $Y2=2.375
r136 15 17 0.130959 $w=4.38e-07 $l=5e-09 $layer=LI1_cond $X=0.305 $Y=2.46
+ $X2=0.305 $Y2=2.465
r137 14 42 3.10218 $w=3.05e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.17 $Y=2.29
+ $X2=0.305 $Y2=2.375
r138 13 37 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.17 $Y=0.73
+ $X2=0.17 $Y2=0.575
r139 13 14 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=0.17 $Y=0.73
+ $X2=0.17 $Y2=2.29
r140 4 48 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.295
+ $Y=2.31 $X2=3.43 $Y2=2.455
r141 3 17 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.215
+ $Y=2.32 $X2=0.36 $Y2=2.465
r142 2 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.025
+ $Y=0.565 $X2=3.165 $Y2=0.775
r143 1 40 182 $w=1.7e-07 $l=3.46194e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.37 $X2=0.415 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_2%VPWR 1 2 3 4 5 6 7 8 9 10 11 36 40 44 48
+ 52 56 60 64 68 72 74 76 79 80 82 83 84 86 91 96 108 112 124 131 136 141 147
+ 150 153 156 159 162 165 168 172
r199 171 172 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.04 $Y=3.33
+ $X2=17.04 $Y2=3.33
r200 168 169 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.08 $Y=3.33
+ $X2=16.08 $Y2=3.33
r201 165 166 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r202 162 163 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r203 159 160 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r204 156 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r205 153 154 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r206 150 151 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r207 147 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r208 145 172 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.56 $Y=3.33
+ $X2=17.04 $Y2=3.33
r209 145 169 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.56 $Y=3.33
+ $X2=16.08 $Y2=3.33
r210 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.56 $Y=3.33
+ $X2=16.56 $Y2=3.33
r211 142 168 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.265 $Y=3.33
+ $X2=16.1 $Y2=3.33
r212 142 144 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=16.265 $Y=3.33
+ $X2=16.56 $Y2=3.33
r213 141 171 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=16.835 $Y=3.33
+ $X2=17.057 $Y2=3.33
r214 141 144 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=16.835 $Y=3.33
+ $X2=16.56 $Y2=3.33
r215 140 169 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=16.08 $Y2=3.33
r216 140 166 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=15.12 $Y2=3.33
r217 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r218 137 165 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.365 $Y=3.33
+ $X2=15.2 $Y2=3.33
r219 137 139 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=15.365 $Y=3.33
+ $X2=15.6 $Y2=3.33
r220 136 168 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.935 $Y=3.33
+ $X2=16.1 $Y2=3.33
r221 136 139 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=15.935 $Y=3.33
+ $X2=15.6 $Y2=3.33
r222 135 166 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=15.12 $Y2=3.33
r223 135 163 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=14.16 $Y2=3.33
r224 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r225 132 162 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=14.305 $Y=3.33
+ $X2=14.035 $Y2=3.33
r226 132 134 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=14.305 $Y=3.33
+ $X2=14.64 $Y2=3.33
r227 131 165 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.035 $Y=3.33
+ $X2=15.2 $Y2=3.33
r228 131 134 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=15.035 $Y=3.33
+ $X2=14.64 $Y2=3.33
r229 130 163 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.16 $Y2=3.33
r230 129 130 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r231 127 130 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=13.68 $Y2=3.33
r232 126 129 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=11.76 $Y=3.33
+ $X2=13.68 $Y2=3.33
r233 126 127 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r234 124 162 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=13.765 $Y=3.33
+ $X2=14.035 $Y2=3.33
r235 124 129 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=13.765 $Y=3.33
+ $X2=13.68 $Y2=3.33
r236 123 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r237 123 160 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.32 $Y2=3.33
r238 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r239 120 159 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.555 $Y=3.33
+ $X2=10.39 $Y2=3.33
r240 120 122 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=10.555 $Y=3.33
+ $X2=11.28 $Y2=3.33
r241 119 160 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r242 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r243 116 157 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r244 115 118 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=9.84 $Y2=3.33
r245 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r246 113 156 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.125 $Y=3.33
+ $X2=7.96 $Y2=3.33
r247 113 115 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.125 $Y=3.33
+ $X2=8.4 $Y2=3.33
r248 112 159 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.225 $Y=3.33
+ $X2=10.39 $Y2=3.33
r249 112 118 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.225 $Y=3.33
+ $X2=9.84 $Y2=3.33
r250 111 157 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r251 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r252 108 156 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.795 $Y=3.33
+ $X2=7.96 $Y2=3.33
r253 108 110 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.795 $Y=3.33
+ $X2=7.44 $Y2=3.33
r254 107 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r255 106 107 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r256 104 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r257 104 154 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r258 103 106 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r259 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r260 101 153 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.305 $Y=3.33
+ $X2=5.17 $Y2=3.33
r261 101 103 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.305 $Y=3.33
+ $X2=5.52 $Y2=3.33
r262 100 154 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=5.04 $Y2=3.33
r263 100 151 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r264 99 100 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r265 97 150 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=2.63 $Y2=3.33
r266 97 99 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=3.12 $Y2=3.33
r267 96 153 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=5.17 $Y2=3.33
r268 96 99 124.936 $w=1.68e-07 $l=1.915e-06 $layer=LI1_cond $X=5.035 $Y=3.33
+ $X2=3.12 $Y2=3.33
r269 95 151 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r270 95 148 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r271 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r272 92 147 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.315 $Y=3.33
+ $X2=1.19 $Y2=3.33
r273 92 94 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=1.315 $Y=3.33
+ $X2=2.16 $Y2=3.33
r274 91 150 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.63 $Y2=3.33
r275 91 94 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.16 $Y2=3.33
r276 89 148 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r277 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r278 86 147 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.19 $Y2=3.33
r279 86 88 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.72 $Y2=3.33
r280 84 119 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=8.64 $Y=3.33
+ $X2=9.84 $Y2=3.33
r281 84 116 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=8.64 $Y=3.33
+ $X2=8.4 $Y2=3.33
r282 82 122 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=11.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r283 82 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.32 $Y=3.33
+ $X2=11.485 $Y2=3.33
r284 81 126 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=11.65 $Y=3.33
+ $X2=11.76 $Y2=3.33
r285 81 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.65 $Y=3.33
+ $X2=11.485 $Y2=3.33
r286 79 106 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.485 $Y=3.33
+ $X2=6.48 $Y2=3.33
r287 79 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.485 $Y=3.33
+ $X2=6.61 $Y2=3.33
r288 78 110 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=6.735 $Y=3.33
+ $X2=7.44 $Y2=3.33
r289 78 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.735 $Y=3.33
+ $X2=6.61 $Y2=3.33
r290 74 171 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=17 $Y=3.245
+ $X2=17.057 $Y2=3.33
r291 74 76 34.7479 $w=3.28e-07 $l=9.95e-07 $layer=LI1_cond $X=17 $Y=3.245 $X2=17
+ $Y2=2.25
r292 70 168 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=16.1 $Y=3.245
+ $X2=16.1 $Y2=3.33
r293 70 72 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=16.1 $Y=3.245
+ $X2=16.1 $Y2=2.78
r294 66 165 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.2 $Y=3.245
+ $X2=15.2 $Y2=3.33
r295 66 68 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=15.2 $Y=3.245
+ $X2=15.2 $Y2=2.78
r296 62 162 2.26835 $w=5.4e-07 $l=8.5e-08 $layer=LI1_cond $X=14.035 $Y=3.245
+ $X2=14.035 $Y2=3.33
r297 62 64 9.52433 $w=5.38e-07 $l=4.3e-07 $layer=LI1_cond $X=14.035 $Y=3.245
+ $X2=14.035 $Y2=2.815
r298 58 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.485 $Y=3.245
+ $X2=11.485 $Y2=3.33
r299 58 60 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=11.485 $Y=3.245
+ $X2=11.485 $Y2=2.895
r300 54 159 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.39 $Y=3.245
+ $X2=10.39 $Y2=3.33
r301 54 56 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.39 $Y=3.245
+ $X2=10.39 $Y2=2.815
r302 50 156 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.96 $Y=3.245
+ $X2=7.96 $Y2=3.33
r303 50 52 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.96 $Y=3.245
+ $X2=7.96 $Y2=2.815
r304 46 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.61 $Y=3.245
+ $X2=6.61 $Y2=3.33
r305 46 48 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6.61 $Y=3.245
+ $X2=6.61 $Y2=2.815
r306 42 153 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.17 $Y=3.245
+ $X2=5.17 $Y2=3.33
r307 42 44 20.7013 $w=2.68e-07 $l=4.85e-07 $layer=LI1_cond $X=5.17 $Y=3.245
+ $X2=5.17 $Y2=2.76
r308 38 150 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=3.245
+ $X2=2.63 $Y2=3.33
r309 38 40 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=2.63 $Y=3.245
+ $X2=2.63 $Y2=2.8
r310 34 147 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=3.245
+ $X2=1.19 $Y2=3.33
r311 34 36 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=1.19 $Y=3.245
+ $X2=1.19 $Y2=2.805
r312 11 76 300 $w=1.7e-07 $l=4.72705e-07 $layer=licon1_PDIFF $count=2 $X=16.865
+ $Y=1.84 $X2=17 $Y2=2.25
r313 10 72 600 $w=1.7e-07 $l=1.00524e-06 $layer=licon1_PDIFF $count=1 $X=15.965
+ $Y=1.84 $X2=16.1 $Y2=2.78
r314 9 68 600 $w=1.7e-07 $l=1.0099e-06 $layer=licon1_PDIFF $count=1 $X=15.055
+ $Y=1.84 $X2=15.2 $Y2=2.78
r315 8 64 600 $w=1.7e-07 $l=3.76331e-07 $layer=licon1_PDIFF $count=1 $X=13.795
+ $Y=2.54 $X2=14.035 $Y2=2.815
r316 7 60 600 $w=1.7e-07 $l=1.00489e-06 $layer=licon1_PDIFF $count=1 $X=11.34
+ $Y=1.96 $X2=11.485 $Y2=2.895
r317 6 56 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=10.245
+ $Y=2.54 $X2=10.39 $Y2=2.815
r318 5 52 600 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=7.815
+ $Y=1.84 $X2=7.96 $Y2=2.815
r319 4 48 600 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=6.425
+ $Y=1.84 $X2=6.57 $Y2=2.815
r320 3 44 600 $w=1.7e-07 $l=6.52457e-07 $layer=licon1_PDIFF $count=1 $X=4.765
+ $Y=2.265 $X2=5.13 $Y2=2.76
r321 2 40 600 $w=1.7e-07 $l=6.47263e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=2.31 $X2=2.59 $Y2=2.8
r322 1 36 600 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=2.32 $X2=1.23 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_2%A_691_113# 1 2 3 4 5 6 21 24 25 26 28 29
+ 30 33 36 37 38 40 41 42 43 47 49 53 56 59 62 67 68
c181 21 0 1.75904e-19 $X=3.84 $Y=2.415
r182 68 70 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.38 $Y=2.395
+ $X2=8.38 $Y2=2.565
r183 58 59 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=3.8 $Y=1.005
+ $X2=3.8 $Y2=2.29
r184 56 58 10.5346 $w=3.83e-07 $l=2.3e-07 $layer=LI1_cond $X=3.692 $Y=0.775
+ $X2=3.692 $Y2=1.005
r185 51 53 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=8.93 $Y=2.65 $X2=8.93
+ $Y2=2.75
r186 50 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.465 $Y=2.565
+ $X2=8.38 $Y2=2.565
r187 49 51 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.805 $Y=2.565
+ $X2=8.93 $Y2=2.65
r188 49 50 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=8.805 $Y=2.565
+ $X2=8.465 $Y2=2.565
r189 45 47 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=8.59 $Y=1.48
+ $X2=8.59 $Y2=0.76
r190 44 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.075 $Y=2.395
+ $X2=7.99 $Y2=2.395
r191 43 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.295 $Y=2.395
+ $X2=8.38 $Y2=2.395
r192 43 44 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.295 $Y=2.395
+ $X2=8.075 $Y2=2.395
r193 41 45 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.465 $Y=1.565
+ $X2=8.59 $Y2=1.48
r194 41 42 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=8.465 $Y=1.565
+ $X2=8.075 $Y2=1.565
r195 40 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.99 $Y=2.31
+ $X2=7.99 $Y2=2.395
r196 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.99 $Y=1.65
+ $X2=8.075 $Y2=1.565
r197 39 40 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=7.99 $Y=1.65
+ $X2=7.99 $Y2=2.31
r198 37 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.905 $Y=2.395
+ $X2=7.99 $Y2=2.395
r199 37 38 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=7.905 $Y=2.395
+ $X2=6.475 $Y2=2.395
r200 36 38 8.2443 $w=5.49e-07 $l=1.77482e-07 $layer=LI1_cond $X=6.39 $Y=2.255
+ $X2=6.475 $Y2=2.395
r201 36 65 8.44444 $w=5.49e-07 $l=5.21248e-07 $layer=LI1_cond $X=6.39 $Y=2.255
+ $X2=6.01 $Y2=2.59
r202 35 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.39 $Y=1.26
+ $X2=6.39 $Y2=1.175
r203 35 36 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=6.39 $Y=1.26
+ $X2=6.39 $Y2=2.255
r204 31 62 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.985 $Y=1.175
+ $X2=6.39 $Y2=1.175
r205 31 33 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.985 $Y=1.09
+ $X2=5.985 $Y2=0.835
r206 29 65 10.0221 $w=5.49e-07 $l=3.22102e-07 $layer=LI1_cond $X=5.845 $Y=2.34
+ $X2=6.01 $Y2=2.59
r207 29 30 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=5.845 $Y=2.34
+ $X2=4.865 $Y2=2.34
r208 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.78 $Y=2.425
+ $X2=4.865 $Y2=2.34
r209 27 28 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.78 $Y=2.425
+ $X2=4.78 $Y2=2.905
r210 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.695 $Y=2.99
+ $X2=4.78 $Y2=2.905
r211 25 26 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.695 $Y=2.99
+ $X2=3.965 $Y2=2.99
r212 22 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.84 $Y=2.905
+ $X2=3.965 $Y2=2.99
r213 22 24 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=3.84 $Y=2.905
+ $X2=3.84 $Y2=2.455
r214 21 59 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=3.84 $Y=2.415
+ $X2=3.84 $Y2=2.29
r215 21 24 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=3.84 $Y=2.415
+ $X2=3.84 $Y2=2.455
r216 6 53 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=8.825
+ $Y=2.54 $X2=8.97 $Y2=2.75
r217 5 65 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=5.875
+ $Y=2.265 $X2=6.01 $Y2=2.42
r218 4 24 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.745
+ $Y=2.31 $X2=3.88 $Y2=2.455
r219 3 47 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=8.485
+ $Y=0.485 $X2=8.63 $Y2=0.76
r220 2 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.845
+ $Y=0.625 $X2=5.985 $Y2=0.835
r221 1 56 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=3.455
+ $Y=0.565 $X2=3.665 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_2%Q 1 2 7 8 9 10 11
r19 10 11 10.8465 $w=3.38e-07 $l=3.2e-07 $layer=LI1_cond $X=15.655 $Y=1.665
+ $X2=15.655 $Y2=1.985
r20 9 10 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=15.655 $Y=1.295
+ $X2=15.655 $Y2=1.665
r21 8 9 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=15.655 $Y=0.925
+ $X2=15.655 $Y2=1.295
r22 7 8 13.8971 $w=3.38e-07 $l=4.1e-07 $layer=LI1_cond $X=15.655 $Y=0.515
+ $X2=15.655 $Y2=0.925
r23 2 11 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=15.515
+ $Y=1.84 $X2=15.65 $Y2=1.985
r24 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=15.52
+ $Y=0.37 $X2=15.66 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_2%Q_N 1 2 7 8 9 10 11 12 13 28 32
r33 29 32 0.501062 $w=2.28e-07 $l=1e-08 $layer=LI1_cond $X=16.55 $Y=1.975
+ $X2=16.55 $Y2=1.985
r34 21 28 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=16.52 $Y=0.96
+ $X2=16.52 $Y2=0.925
r35 12 13 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=16.55 $Y=2.405
+ $X2=16.55 $Y2=2.775
r36 11 29 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=16.56 $Y=1.89
+ $X2=16.55 $Y2=1.89
r37 11 12 17.938 $w=2.28e-07 $l=3.58e-07 $layer=LI1_cond $X=16.55 $Y=2.047
+ $X2=16.55 $Y2=2.405
r38 11 32 3.10659 $w=2.28e-07 $l=6.2e-08 $layer=LI1_cond $X=16.55 $Y=2.047
+ $X2=16.55 $Y2=1.985
r39 10 21 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=16.56 $Y=1.045
+ $X2=16.52 $Y2=1.045
r40 10 28 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=16.52 $Y=0.9
+ $X2=16.52 $Y2=0.925
r41 9 10 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=16.52 $Y=0.515
+ $X2=16.52 $Y2=0.9
r42 8 11 24.2695 $w=1.68e-07 $l=3.72e-07 $layer=LI1_cond $X=16.932 $Y=1.89
+ $X2=16.56 $Y2=1.89
r43 7 10 24.2695 $w=1.68e-07 $l=3.72e-07 $layer=LI1_cond $X=16.932 $Y=1.045
+ $X2=16.56 $Y2=1.045
r44 7 8 17.3624 $w=4.63e-07 $l=6.75e-07 $layer=LI1_cond $X=16.932 $Y=1.13
+ $X2=16.932 $Y2=1.805
r45 2 32 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=16.415
+ $Y=1.84 $X2=16.55 $Y2=1.985
r46 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=16.38
+ $Y=0.37 $X2=16.52 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXBP_2%VGND 1 2 3 4 5 6 7 8 9 10 11 36 40 44 48
+ 52 56 60 62 63 68 70 74 76 80 82 84 87 88 90 91 93 94 96 105 109 118 122 134
+ 140 143 146 149 152 155 159 162 166
r220 165 166 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.04 $Y=0
+ $X2=17.04 $Y2=0
r221 162 163 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.08 $Y=0
+ $X2=16.08 $Y2=0
r222 160 163 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.12 $Y=0
+ $X2=16.08 $Y2=0
r223 159 160 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r224 156 160 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=15.12 $Y2=0
r225 155 156 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r226 152 153 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r227 149 150 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r228 146 147 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r229 143 144 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r230 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r231 138 166 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.56 $Y=0
+ $X2=17.04 $Y2=0
r232 138 163 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.56 $Y=0
+ $X2=16.08 $Y2=0
r233 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.56 $Y=0
+ $X2=16.56 $Y2=0
r234 135 162 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.175 $Y=0
+ $X2=16.09 $Y2=0
r235 135 137 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=16.175 $Y=0
+ $X2=16.56 $Y2=0
r236 134 165 4.03428 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=16.855 $Y=0
+ $X2=17.067 $Y2=0
r237 134 137 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=16.855 $Y=0
+ $X2=16.56 $Y2=0
r238 133 156 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=14.16 $Y2=0
r239 132 133 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r240 130 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=13.2 $Y2=0
r241 130 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r242 129 132 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=12.24 $Y=0
+ $X2=13.2 $Y2=0
r243 129 130 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r244 127 152 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.96 $Y=0
+ $X2=11.835 $Y2=0
r245 127 129 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=11.96 $Y=0
+ $X2=12.24 $Y2=0
r246 126 153 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.76 $Y2=0
r247 126 150 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r248 125 126 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r249 123 149 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.52 $Y=0
+ $X2=10.395 $Y2=0
r250 123 125 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.52 $Y=0
+ $X2=10.8 $Y2=0
r251 122 152 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.71 $Y=0
+ $X2=11.835 $Y2=0
r252 122 125 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=11.71 $Y=0
+ $X2=10.8 $Y2=0
r253 120 121 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r254 118 149 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.27 $Y=0
+ $X2=10.395 $Y2=0
r255 118 120 153.316 $w=1.68e-07 $l=2.35e-06 $layer=LI1_cond $X=10.27 $Y=0
+ $X2=7.92 $Y2=0
r256 117 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r257 117 147 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.48 $Y2=0
r258 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r259 114 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.745 $Y=0
+ $X2=6.58 $Y2=0
r260 114 116 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.745 $Y=0
+ $X2=7.44 $Y2=0
r261 113 147 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=6.48 $Y2=0
r262 113 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=5.04 $Y2=0
r263 112 113 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r264 110 143 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.29 $Y=0
+ $X2=5.125 $Y2=0
r265 110 112 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.29 $Y=0
+ $X2=5.52 $Y2=0
r266 109 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.415 $Y=0
+ $X2=6.58 $Y2=0
r267 109 112 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=6.415 $Y=0
+ $X2=5.52 $Y2=0
r268 108 144 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=5.04 $Y2=0
r269 107 108 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r270 105 143 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.96 $Y=0
+ $X2=5.125 $Y2=0
r271 105 107 151.358 $w=1.68e-07 $l=2.32e-06 $layer=LI1_cond $X=4.96 $Y=0
+ $X2=2.64 $Y2=0
r272 104 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=2.64 $Y2=0
r273 104 141 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.2 $Y2=0
r274 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r275 101 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.4 $Y=0
+ $X2=1.235 $Y2=0
r276 101 103 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=1.4 $Y=0 $X2=2.16
+ $Y2=0
r277 99 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r278 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r279 96 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.07 $Y=0
+ $X2=1.235 $Y2=0
r280 96 98 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.07 $Y=0 $X2=0.72
+ $Y2=0
r281 94 150 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=8.64 $Y=0
+ $X2=10.32 $Y2=0
r282 94 121 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=8.64 $Y=0
+ $X2=7.92 $Y2=0
r283 93 132 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=13.32 $Y=0
+ $X2=13.2 $Y2=0
r284 90 116 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.555 $Y=0
+ $X2=7.44 $Y2=0
r285 90 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.555 $Y=0 $X2=7.64
+ $Y2=0
r286 89 120 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=7.725 $Y=0
+ $X2=7.92 $Y2=0
r287 89 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.725 $Y=0 $X2=7.64
+ $Y2=0
r288 87 103 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.16
+ $Y2=0
r289 87 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.18 $Y=0 $X2=2.345
+ $Y2=0
r290 86 107 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.51 $Y=0 $X2=2.64
+ $Y2=0
r291 86 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.51 $Y=0 $X2=2.345
+ $Y2=0
r292 82 165 3.17794 $w=2.6e-07 $l=1.19143e-07 $layer=LI1_cond $X=16.985 $Y=0.085
+ $X2=17.067 $Y2=0
r293 82 84 23.9354 $w=2.58e-07 $l=5.4e-07 $layer=LI1_cond $X=16.985 $Y=0.085
+ $X2=16.985 $Y2=0.625
r294 78 162 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.09 $Y=0.085
+ $X2=16.09 $Y2=0
r295 78 80 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=16.09 $Y=0.085
+ $X2=16.09 $Y2=0.515
r296 77 159 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.315 $Y=0
+ $X2=15.19 $Y2=0
r297 76 162 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.005 $Y=0
+ $X2=16.09 $Y2=0
r298 76 77 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=16.005 $Y=0
+ $X2=15.315 $Y2=0
r299 72 159 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=15.19 $Y=0.085
+ $X2=15.19 $Y2=0
r300 72 74 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=15.19 $Y=0.085
+ $X2=15.19 $Y2=0.515
r301 71 155 3.47156 $w=4.27e-07 $l=3.17402e-07 $layer=LI1_cond $X=14.335 $Y=0
+ $X2=14.2 $Y2=0.257
r302 70 159 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.065 $Y=0
+ $X2=15.19 $Y2=0
r303 70 71 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=15.065 $Y=0
+ $X2=14.335 $Y2=0
r304 66 155 3.03886 $w=2.7e-07 $l=3.43e-07 $layer=LI1_cond $X=14.2 $Y=0.6
+ $X2=14.2 $Y2=0.257
r305 66 68 15.1525 $w=2.68e-07 $l=3.55e-07 $layer=LI1_cond $X=14.2 $Y=0.6
+ $X2=14.2 $Y2=0.955
r306 63 93 13.7992 $w=6.83e-07 $l=3.42e-07 $layer=LI1_cond $X=13.662 $Y=0.257
+ $X2=13.32 $Y2=0.257
r307 63 65 3.19536 $w=6.83e-07 $l=1.83e-07 $layer=LI1_cond $X=13.662 $Y=0.257
+ $X2=13.845 $Y2=0.257
r308 62 155 3.47156 $w=4.27e-07 $l=1.35e-07 $layer=LI1_cond $X=14.065 $Y=0.257
+ $X2=14.2 $Y2=0.257
r309 62 65 3.84142 $w=6.83e-07 $l=2.2e-07 $layer=LI1_cond $X=14.065 $Y=0.257
+ $X2=13.845 $Y2=0.257
r310 58 152 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.835 $Y=0.085
+ $X2=11.835 $Y2=0
r311 58 60 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.835 $Y=0.085
+ $X2=11.835 $Y2=0.515
r312 54 149 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.395 $Y=0.085
+ $X2=10.395 $Y2=0
r313 54 56 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.395 $Y=0.085
+ $X2=10.395 $Y2=0.515
r314 50 91 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.64 $Y=0.085
+ $X2=7.64 $Y2=0
r315 50 52 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=7.64 $Y=0.085
+ $X2=7.64 $Y2=0.515
r316 46 146 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.58 $Y=0.085
+ $X2=6.58 $Y2=0
r317 46 48 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.58 $Y=0.085
+ $X2=6.58 $Y2=0.495
r318 42 143 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.125 $Y=0.085
+ $X2=5.125 $Y2=0
r319 42 44 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=5.125 $Y=0.085
+ $X2=5.125 $Y2=0.805
r320 38 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.345 $Y=0.085
+ $X2=2.345 $Y2=0
r321 38 40 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=2.345 $Y=0.085
+ $X2=2.345 $Y2=0.775
r322 34 140 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=0.085
+ $X2=1.235 $Y2=0
r323 34 36 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.235 $Y=0.085
+ $X2=1.235 $Y2=0.58
r324 11 84 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=16.81
+ $Y=0.37 $X2=16.95 $Y2=0.625
r325 10 80 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=15.95
+ $Y=0.37 $X2=16.09 $Y2=0.515
r326 9 74 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=15.085
+ $Y=0.37 $X2=15.23 $Y2=0.515
r327 8 155 182 $w=1.7e-07 $l=9.6478e-07 $layer=licon1_NDIFF $count=1 $X=13.345
+ $Y=0.37 $X2=14.24 $Y2=0.515
r328 8 68 182 $w=1.7e-07 $l=1.15091e-06 $layer=licon1_NDIFF $count=1 $X=13.345
+ $Y=0.37 $X2=14.24 $Y2=0.955
r329 8 65 91 $w=1.7e-07 $l=5.67891e-07 $layer=licon1_NDIFF $count=2 $X=13.345
+ $Y=0.37 $X2=13.845 $Y2=0.515
r330 7 60 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=11.65
+ $Y=0.37 $X2=11.795 $Y2=0.515
r331 6 56 182 $w=1.7e-07 $l=2.34521e-07 $layer=licon1_NDIFF $count=1 $X=10.215
+ $Y=0.485 $X2=10.435 $Y2=0.515
r332 5 52 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=7.495
+ $Y=0.37 $X2=7.64 $Y2=0.515
r333 4 48 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=6.435
+ $Y=0.37 $X2=6.58 $Y2=0.495
r334 3 44 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=4.915
+ $Y=0.625 $X2=5.125 $Y2=0.805
r335 2 40 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=2.135
+ $Y=0.565 $X2=2.345 $Y2=0.775
r336 1 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.37 $X2=1.235 $Y2=0.58
.ends


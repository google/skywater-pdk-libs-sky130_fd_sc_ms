* File: sky130_fd_sc_ms__a311oi_4.pex.spice
* Created: Fri Aug 28 17:06:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A311OI_4%A3 3 7 11 15 19 23 27 31 33 34 35 51 53
c73 31 0 1.47716e-19 $X=1.845 $Y=2.4
c74 19 0 1.47716e-19 $X=1.395 $Y=2.4
c75 11 0 1.53462e-19 $X=0.945 $Y=2.4
r76 52 53 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.82 $Y=1.515
+ $X2=1.845 $Y2=1.515
r77 50 52 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=1.71 $Y=1.515
+ $X2=1.82 $Y2=1.515
r78 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.71
+ $Y=1.515 $X2=1.71 $Y2=1.515
r79 48 50 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=1.395 $Y=1.515
+ $X2=1.71 $Y2=1.515
r80 47 48 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=1.39 $Y=1.515
+ $X2=1.395 $Y2=1.515
r81 46 47 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.96 $Y=1.515
+ $X2=1.39 $Y2=1.515
r82 45 46 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.945 $Y=1.515
+ $X2=0.96 $Y2=1.515
r83 43 45 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=0.69 $Y=1.515
+ $X2=0.945 $Y2=1.515
r84 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.69
+ $Y=1.515 $X2=0.69 $Y2=1.515
r85 41 43 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.53 $Y=1.515
+ $X2=0.69 $Y2=1.515
r86 39 41 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=0.495 $Y=1.515
+ $X2=0.53 $Y2=1.515
r87 35 51 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=1.68 $Y=1.565 $X2=1.71
+ $Y2=1.565
r88 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.68 $Y2=1.565
r89 33 34 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r90 33 44 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=0.72 $Y=1.565 $X2=0.69
+ $Y2=1.565
r91 29 53 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.68
+ $X2=1.845 $Y2=1.515
r92 29 31 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.845 $Y=1.68
+ $X2=1.845 $Y2=2.4
r93 25 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.82 $Y=1.35
+ $X2=1.82 $Y2=1.515
r94 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.82 $Y=1.35
+ $X2=1.82 $Y2=0.74
r95 21 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.39 $Y=1.35
+ $X2=1.39 $Y2=1.515
r96 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.39 $Y=1.35
+ $X2=1.39 $Y2=0.74
r97 17 48 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.395 $Y=1.68
+ $X2=1.395 $Y2=1.515
r98 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.395 $Y=1.68
+ $X2=1.395 $Y2=2.4
r99 13 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.35
+ $X2=0.96 $Y2=1.515
r100 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.96 $Y=1.35
+ $X2=0.96 $Y2=0.74
r101 9 45 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=1.68
+ $X2=0.945 $Y2=1.515
r102 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.945 $Y=1.68
+ $X2=0.945 $Y2=2.4
r103 5 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.35
+ $X2=0.53 $Y2=1.515
r104 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.53 $Y=1.35 $X2=0.53
+ $Y2=0.74
r105 1 39 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.68
+ $X2=0.495 $Y2=1.515
r106 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.495 $Y=1.68
+ $X2=0.495 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_4%A2 3 7 11 15 19 23 27 31 33 34 35 36 53
c80 31 0 1.47716e-19 $X=3.645 $Y=2.4
c81 23 0 1.47716e-19 $X=3.195 $Y=2.4
c82 15 0 1.47716e-19 $X=2.745 $Y=2.4
c83 7 0 1.47716e-19 $X=2.295 $Y=2.4
r84 53 54 15.5245 $w=3.26e-07 $l=1.05e-07 $layer=POLY_cond $X=3.54 $Y=1.515
+ $X2=3.645 $Y2=1.515
r85 51 53 22.1779 $w=3.26e-07 $l=1.5e-07 $layer=POLY_cond $X=3.39 $Y=1.515
+ $X2=3.54 $Y2=1.515
r86 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.39
+ $Y=1.515 $X2=3.39 $Y2=1.515
r87 49 51 28.8313 $w=3.26e-07 $l=1.95e-07 $layer=POLY_cond $X=3.195 $Y=1.515
+ $X2=3.39 $Y2=1.515
r88 48 49 12.5675 $w=3.26e-07 $l=8.5e-08 $layer=POLY_cond $X=3.11 $Y=1.515
+ $X2=3.195 $Y2=1.515
r89 47 48 53.9663 $w=3.26e-07 $l=3.65e-07 $layer=POLY_cond $X=2.745 $Y=1.515
+ $X2=3.11 $Y2=1.515
r90 46 47 9.61043 $w=3.26e-07 $l=6.5e-08 $layer=POLY_cond $X=2.68 $Y=1.515
+ $X2=2.745 $Y2=1.515
r91 44 46 45.8344 $w=3.26e-07 $l=3.1e-07 $layer=POLY_cond $X=2.37 $Y=1.515
+ $X2=2.68 $Y2=1.515
r92 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.37
+ $Y=1.515 $X2=2.37 $Y2=1.515
r93 42 44 11.089 $w=3.26e-07 $l=7.5e-08 $layer=POLY_cond $X=2.295 $Y=1.515
+ $X2=2.37 $Y2=1.515
r94 41 42 6.65337 $w=3.26e-07 $l=4.5e-08 $layer=POLY_cond $X=2.25 $Y=1.515
+ $X2=2.295 $Y2=1.515
r95 36 52 5.62821 $w=4.28e-07 $l=2.1e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.39 $Y2=1.565
r96 35 52 7.23627 $w=4.28e-07 $l=2.7e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.39 $Y2=1.565
r97 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.12 $Y2=1.565
r98 34 45 7.23627 $w=4.28e-07 $l=2.7e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.37 $Y2=1.565
r99 33 45 5.62821 $w=4.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.37 $Y2=1.565
r100 29 54 16.6478 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.645 $Y=1.68
+ $X2=3.645 $Y2=1.515
r101 29 31 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.645 $Y=1.68
+ $X2=3.645 $Y2=2.4
r102 25 53 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.54 $Y=1.35
+ $X2=3.54 $Y2=1.515
r103 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.54 $Y=1.35
+ $X2=3.54 $Y2=0.74
r104 21 49 16.6478 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.195 $Y=1.68
+ $X2=3.195 $Y2=1.515
r105 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.195 $Y=1.68
+ $X2=3.195 $Y2=2.4
r106 17 48 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.11 $Y=1.35
+ $X2=3.11 $Y2=1.515
r107 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.11 $Y=1.35
+ $X2=3.11 $Y2=0.74
r108 13 47 16.6478 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.745 $Y=1.68
+ $X2=2.745 $Y2=1.515
r109 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.745 $Y=1.68
+ $X2=2.745 $Y2=2.4
r110 9 46 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.35
+ $X2=2.68 $Y2=1.515
r111 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.68 $Y=1.35
+ $X2=2.68 $Y2=0.74
r112 5 42 16.6478 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=1.68
+ $X2=2.295 $Y2=1.515
r113 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.295 $Y=1.68
+ $X2=2.295 $Y2=2.4
r114 1 41 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.35
+ $X2=2.25 $Y2=1.515
r115 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.25 $Y=1.35 $X2=2.25
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_4%A1 3 5 6 9 13 17 21 25 29 33 35 36 49
c82 49 0 1.98771e-19 $X=5.91 $Y=1.515
c83 33 0 8.65694e-20 $X=6 $Y=0.74
c84 25 0 1.53462e-19 $X=5.445 $Y=2.4
r85 49 51 13.9935 $w=3.1e-07 $l=9e-08 $layer=POLY_cond $X=5.91 $Y=1.515 $X2=6
+ $Y2=1.515
r86 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.91
+ $Y=1.515 $X2=5.91 $Y2=1.515
r87 47 49 52.8645 $w=3.1e-07 $l=3.4e-07 $layer=POLY_cond $X=5.57 $Y=1.515
+ $X2=5.91 $Y2=1.515
r88 46 47 19.4355 $w=3.1e-07 $l=1.25e-07 $layer=POLY_cond $X=5.445 $Y=1.515
+ $X2=5.57 $Y2=1.515
r89 44 46 38.0935 $w=3.1e-07 $l=2.45e-07 $layer=POLY_cond $X=5.2 $Y=1.515
+ $X2=5.445 $Y2=1.515
r90 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.2
+ $Y=1.515 $X2=5.2 $Y2=1.515
r91 42 44 9.32903 $w=3.1e-07 $l=6e-08 $layer=POLY_cond $X=5.14 $Y=1.515 $X2=5.2
+ $Y2=1.515
r92 41 42 22.5452 $w=3.1e-07 $l=1.45e-07 $layer=POLY_cond $X=4.995 $Y=1.515
+ $X2=5.14 $Y2=1.515
r93 40 41 44.3129 $w=3.1e-07 $l=2.85e-07 $layer=POLY_cond $X=4.71 $Y=1.515
+ $X2=4.995 $Y2=1.515
r94 36 50 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=6 $Y=1.565 $X2=5.91
+ $Y2=1.565
r95 35 50 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.91 $Y2=1.565
r96 35 45 8.57632 $w=4.28e-07 $l=3.2e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.2 $Y2=1.565
r97 31 51 19.7411 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6 $Y=1.35 $X2=6
+ $Y2=1.515
r98 31 33 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6 $Y=1.35 $X2=6
+ $Y2=0.74
r99 27 47 19.7411 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.57 $Y=1.35
+ $X2=5.57 $Y2=1.515
r100 27 29 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.57 $Y=1.35
+ $X2=5.57 $Y2=0.74
r101 23 46 15.4789 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.445 $Y=1.68
+ $X2=5.445 $Y2=1.515
r102 23 25 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.445 $Y=1.68
+ $X2=5.445 $Y2=2.4
r103 19 42 19.7411 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.14 $Y=1.35
+ $X2=5.14 $Y2=1.515
r104 19 21 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.14 $Y=1.35
+ $X2=5.14 $Y2=0.74
r105 15 41 15.4789 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.995 $Y=1.68
+ $X2=4.995 $Y2=1.515
r106 15 17 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.995 $Y=1.68
+ $X2=4.995 $Y2=2.4
r107 11 40 19.7411 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.71 $Y=1.35
+ $X2=4.71 $Y2=1.515
r108 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.71 $Y=1.35
+ $X2=4.71 $Y2=0.74
r109 7 40 25.6548 $w=3.1e-07 $l=2.33345e-07 $layer=POLY_cond $X=4.545 $Y=1.68
+ $X2=4.71 $Y2=1.515
r110 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.545 $Y=1.68
+ $X2=4.545 $Y2=2.4
r111 5 7 26.8705 $w=3.1e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.455 $Y=1.605
+ $X2=4.545 $Y2=1.68
r112 5 6 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.455 $Y=1.605
+ $X2=4.185 $Y2=1.605
r113 1 6 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.095 $Y=1.68
+ $X2=4.185 $Y2=1.605
r114 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.095 $Y=1.68
+ $X2=4.095 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_4%B1 3 7 11 15 19 23 25 26 39 41
c80 41 0 2.85341e-19 $X=7.32 $Y=1.415
c81 23 0 1.70682e-19 $X=7.765 $Y=2.4
c82 7 0 1.0484e-19 $X=6.43 $Y=0.74
r83 39 40 8.25857 $w=3.21e-07 $l=5.5e-08 $layer=POLY_cond $X=7.71 $Y=1.485
+ $X2=7.765 $Y2=1.485
r84 37 39 13.514 $w=3.21e-07 $l=9e-08 $layer=POLY_cond $X=7.62 $Y=1.485 $X2=7.71
+ $Y2=1.485
r85 37 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.62
+ $Y=1.485 $X2=7.62 $Y2=1.485
r86 35 37 45.7975 $w=3.21e-07 $l=3.05e-07 $layer=POLY_cond $X=7.315 $Y=1.485
+ $X2=7.62 $Y2=1.485
r87 33 35 56.3084 $w=3.21e-07 $l=3.75e-07 $layer=POLY_cond $X=6.94 $Y=1.485
+ $X2=7.315 $Y2=1.485
r88 33 34 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.94
+ $Y=1.485 $X2=6.94 $Y2=1.485
r89 31 33 11.2617 $w=3.21e-07 $l=7.5e-08 $layer=POLY_cond $X=6.865 $Y=1.485
+ $X2=6.94 $Y2=1.485
r90 30 31 65.3178 $w=3.21e-07 $l=4.35e-07 $layer=POLY_cond $X=6.43 $Y=1.485
+ $X2=6.865 $Y2=1.485
r91 29 30 2.25234 $w=3.21e-07 $l=1.5e-08 $layer=POLY_cond $X=6.415 $Y=1.485
+ $X2=6.43 $Y2=1.485
r92 26 38 5.49 $w=4e-07 $l=1.8e-07 $layer=LI1_cond $X=7.44 $Y=1.415 $X2=7.62
+ $Y2=1.415
r93 26 41 3.4204 $w=4.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.44 $Y=1.415 $X2=7.32
+ $Y2=1.415
r94 25 41 9.16145 $w=4.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.96 $Y=1.415
+ $X2=7.32 $Y2=1.415
r95 25 34 0.50897 $w=4.68e-07 $l=2e-08 $layer=LI1_cond $X=6.96 $Y=1.415 $X2=6.94
+ $Y2=1.415
r96 21 40 16.2883 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.765 $Y=1.65
+ $X2=7.765 $Y2=1.485
r97 21 23 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=7.765 $Y=1.65
+ $X2=7.765 $Y2=2.4
r98 17 39 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.71 $Y=1.32
+ $X2=7.71 $Y2=1.485
r99 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.71 $Y=1.32
+ $X2=7.71 $Y2=0.74
r100 13 35 16.2883 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.315 $Y=1.65
+ $X2=7.315 $Y2=1.485
r101 13 15 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=7.315 $Y=1.65
+ $X2=7.315 $Y2=2.4
r102 9 31 16.2883 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.865 $Y=1.65
+ $X2=6.865 $Y2=1.485
r103 9 11 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=6.865 $Y=1.65
+ $X2=6.865 $Y2=2.4
r104 5 30 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.43 $Y=1.32
+ $X2=6.43 $Y2=1.485
r105 5 7 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.43 $Y=1.32 $X2=6.43
+ $Y2=0.74
r106 1 29 16.2883 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.415 $Y=1.65
+ $X2=6.415 $Y2=1.485
r107 1 3 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=6.415 $Y=1.65
+ $X2=6.415 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_4%C1 1 3 6 8 10 13 17 19 23 25 26 39 41 42 51
c76 1 0 1.44963e-19 $X=8.14 $Y=1.22
r77 42 51 2.36628 $w=3.7e-07 $l=7e-08 $layer=LI1_cond $X=8.47 $Y=1.365 $X2=8.4
+ $Y2=1.365
r78 40 41 19.2659 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.115 $Y=1.385
+ $X2=9.205 $Y2=1.385
r79 38 40 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=8.91 $Y=1.385
+ $X2=9.115 $Y2=1.385
r80 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.91
+ $Y=1.385 $X2=8.91 $Y2=1.385
r81 36 38 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=8.665 $Y=1.385
+ $X2=8.91 $Y2=1.385
r82 34 36 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=8.57 $Y=1.385
+ $X2=8.665 $Y2=1.385
r83 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.57
+ $Y=1.385 $X2=8.57 $Y2=1.385
r84 32 34 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=8.215 $Y=1.385
+ $X2=8.57 $Y2=1.385
r85 30 32 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.14 $Y=1.385
+ $X2=8.215 $Y2=1.385
r86 26 39 0.934413 $w=3.68e-07 $l=3e-08 $layer=LI1_cond $X=8.88 $Y=1.365
+ $X2=8.91 $Y2=1.365
r87 26 35 9.6556 $w=3.68e-07 $l=3.1e-07 $layer=LI1_cond $X=8.88 $Y=1.365
+ $X2=8.57 $Y2=1.365
r88 25 51 0.28046 $w=3.48e-07 $l=8e-09 $layer=LI1_cond $X=8.392 $Y=1.365 $X2=8.4
+ $Y2=1.365
r89 25 35 2.89668 $w=3.68e-07 $l=9.3e-08 $layer=LI1_cond $X=8.477 $Y=1.365
+ $X2=8.57 $Y2=1.365
r90 25 42 0.21803 $w=3.68e-07 $l=7e-09 $layer=LI1_cond $X=8.477 $Y=1.365
+ $X2=8.47 $Y2=1.365
r91 21 23 361.5 $w=1.8e-07 $l=9.3e-07 $layer=POLY_cond $X=9.565 $Y=1.47
+ $X2=9.565 $Y2=2.4
r92 19 21 27.8695 $w=2.5e-07 $l=1.63936e-07 $layer=POLY_cond $X=9.475 $Y=1.345
+ $X2=9.565 $Y2=1.47
r93 19 41 67.0825 $w=2.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.475 $Y=1.345
+ $X2=9.205 $Y2=1.345
r94 15 40 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.115 $Y=1.55
+ $X2=9.115 $Y2=1.385
r95 15 17 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=9.115 $Y=1.55
+ $X2=9.115 $Y2=2.4
r96 11 36 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.665 $Y=1.55
+ $X2=8.665 $Y2=1.385
r97 11 13 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=8.665 $Y=1.55
+ $X2=8.665 $Y2=2.4
r98 8 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.57 $Y=1.22
+ $X2=8.57 $Y2=1.385
r99 8 10 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.57 $Y=1.22 $X2=8.57
+ $Y2=0.74
r100 4 32 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.215 $Y=1.55
+ $X2=8.215 $Y2=1.385
r101 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=8.215 $Y=1.55
+ $X2=8.215 $Y2=2.4
r102 1 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.14 $Y=1.22
+ $X2=8.14 $Y2=1.385
r103 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.14 $Y=1.22 $X2=8.14
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_4%VPWR 1 2 3 4 5 6 7 22 24 30 34 38 42 46 48
+ 52 55 56 58 59 61 62 63 64 65 67 90 91 97 100
r141 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r142 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r143 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r144 90 91 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r145 88 91 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=6 $Y=3.33 $X2=9.84
+ $Y2=3.33
r146 88 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r147 87 90 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=9.84
+ $Y2=3.33
r148 87 88 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6 $Y=3.33
+ $X2=6 $Y2=3.33
r149 85 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.835 $Y=3.33
+ $X2=5.67 $Y2=3.33
r150 85 87 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.835 $Y=3.33
+ $X2=6 $Y2=3.33
r151 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r152 81 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r153 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r154 78 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r155 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r156 75 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r157 75 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r158 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r159 72 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.17 $Y2=3.33
r160 72 74 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.68 $Y2=3.33
r161 71 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r162 71 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r163 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r164 68 94 4.02368 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.177 $Y2=3.33
r165 68 70 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.72 $Y2=3.33
r166 67 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.17 $Y2=3.33
r167 67 70 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.72 $Y2=3.33
r168 65 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r169 65 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r170 63 83 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.605 $Y=3.33
+ $X2=4.56 $Y2=3.33
r171 63 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.605 $Y=3.33
+ $X2=4.73 $Y2=3.33
r172 61 80 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=3.6 $Y2=3.33
r173 61 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=3.87 $Y2=3.33
r174 60 83 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=4.035 $Y=3.33
+ $X2=4.56 $Y2=3.33
r175 60 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.035 $Y=3.33
+ $X2=3.87 $Y2=3.33
r176 58 77 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=2.64 $Y2=3.33
r177 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=3.33
+ $X2=2.97 $Y2=3.33
r178 57 80 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.135 $Y=3.33
+ $X2=3.6 $Y2=3.33
r179 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.135 $Y=3.33
+ $X2=2.97 $Y2=3.33
r180 55 74 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=1.68 $Y2=3.33
r181 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=2.07 $Y2=3.33
r182 54 77 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.235 $Y=3.33
+ $X2=2.64 $Y2=3.33
r183 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=3.33
+ $X2=2.07 $Y2=3.33
r184 50 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.67 $Y=3.245
+ $X2=5.67 $Y2=3.33
r185 50 52 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=5.67 $Y=3.245
+ $X2=5.67 $Y2=2.455
r186 49 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=4.73 $Y2=3.33
r187 48 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.505 $Y=3.33
+ $X2=5.67 $Y2=3.33
r188 48 49 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.505 $Y=3.33
+ $X2=4.855 $Y2=3.33
r189 44 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.73 $Y=3.245
+ $X2=4.73 $Y2=3.33
r190 44 46 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=4.73 $Y=3.245
+ $X2=4.73 $Y2=2.455
r191 40 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.87 $Y=3.245
+ $X2=3.87 $Y2=3.33
r192 40 42 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=3.87 $Y=3.245
+ $X2=3.87 $Y2=2.455
r193 36 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=3.245
+ $X2=2.97 $Y2=3.33
r194 36 38 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.97 $Y=3.245
+ $X2=2.97 $Y2=2.455
r195 32 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=3.245
+ $X2=2.07 $Y2=3.33
r196 32 34 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.07 $Y=3.245
+ $X2=2.07 $Y2=2.455
r197 28 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=3.33
r198 28 30 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=2.455
r199 24 27 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.23 $Y=1.985
+ $X2=0.23 $Y2=2.815
r200 22 94 3.11948 $w=2.5e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.23 $Y=3.245
+ $X2=0.177 $Y2=3.33
r201 22 27 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.23 $Y=3.245
+ $X2=0.23 $Y2=2.815
r202 7 52 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=5.535
+ $Y=1.84 $X2=5.67 $Y2=2.455
r203 6 46 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=4.635
+ $Y=1.84 $X2=4.77 $Y2=2.455
r204 5 42 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=3.735
+ $Y=1.84 $X2=3.87 $Y2=2.455
r205 4 38 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=2.835
+ $Y=1.84 $X2=2.97 $Y2=2.455
r206 3 34 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.935
+ $Y=1.84 $X2=2.07 $Y2=2.455
r207 2 30 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.035
+ $Y=1.84 $X2=1.17 $Y2=2.455
r208 1 27 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=2.815
r209 1 24 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.27 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_4%A_117_368# 1 2 3 4 5 6 7 8 25 27 29 33 35
+ 39 41 45 47 51 53 57 59 63 65 67 69 74 76 78 80 82 84
c108 67 0 1.70682e-19 $X=7.54 $Y=2.15
c109 57 0 1.53462e-19 $X=5.22 $Y=2.815
c110 45 0 2.95431e-19 $X=3.42 $Y=2.815
c111 39 0 2.95431e-19 $X=2.52 $Y=2.815
c112 33 0 2.95431e-19 $X=1.62 $Y=2.815
c113 27 0 1.53462e-19 $X=0.72 $Y=2.815
r114 67 86 4.18573 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.54 $Y=2.15
+ $X2=7.54 $Y2=1.985
r115 67 69 21.0446 $w=2.28e-07 $l=4.2e-07 $layer=LI1_cond $X=7.54 $Y=2.15
+ $X2=7.54 $Y2=2.57
r116 66 84 4.81705 $w=2.5e-07 $l=1.4e-07 $layer=LI1_cond $X=6.755 $Y=1.985
+ $X2=6.615 $Y2=1.985
r117 65 86 2.91733 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=7.425 $Y=1.985
+ $X2=7.54 $Y2=1.985
r118 65 66 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=7.425 $Y=1.985
+ $X2=6.755 $Y2=1.985
r119 61 84 1.64447 $w=2.3e-07 $l=1.77059e-07 $layer=LI1_cond $X=6.64 $Y=2.15
+ $X2=6.615 $Y2=1.985
r120 61 63 21.0446 $w=2.28e-07 $l=4.2e-07 $layer=LI1_cond $X=6.64 $Y=2.15
+ $X2=6.64 $Y2=2.57
r121 60 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.305 $Y=2.035
+ $X2=5.18 $Y2=2.035
r122 59 84 4.81705 $w=2.5e-07 $l=1.63095e-07 $layer=LI1_cond $X=6.475 $Y=2.035
+ $X2=6.615 $Y2=1.985
r123 59 60 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=6.475 $Y=2.035
+ $X2=5.305 $Y2=2.035
r124 55 82 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.18 $Y=2.12
+ $X2=5.18 $Y2=2.035
r125 55 57 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=5.18 $Y=2.12
+ $X2=5.18 $Y2=2.815
r126 54 80 5.16603 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=4.405 $Y=2.035
+ $X2=4.32 $Y2=1.97
r127 53 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.055 $Y=2.035
+ $X2=5.18 $Y2=2.035
r128 53 54 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.055 $Y=2.035
+ $X2=4.405 $Y2=2.035
r129 49 80 1.34256 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.32 $Y=2.12
+ $X2=4.32 $Y2=1.97
r130 49 51 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.32 $Y=2.12
+ $X2=4.32 $Y2=2.4
r131 48 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.505 $Y=2.035
+ $X2=3.42 $Y2=2.035
r132 47 80 5.16603 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=4.235 $Y=2.035
+ $X2=4.32 $Y2=1.97
r133 47 48 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.235 $Y=2.035
+ $X2=3.505 $Y2=2.035
r134 43 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=2.12
+ $X2=3.42 $Y2=2.035
r135 43 45 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.42 $Y=2.12
+ $X2=3.42 $Y2=2.815
r136 42 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.605 $Y=2.035
+ $X2=2.52 $Y2=2.035
r137 41 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=2.035
+ $X2=3.42 $Y2=2.035
r138 41 42 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.335 $Y=2.035
+ $X2=2.605 $Y2=2.035
r139 37 76 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.52 $Y=2.12
+ $X2=2.52 $Y2=2.035
r140 37 39 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.52 $Y=2.12
+ $X2=2.52 $Y2=2.815
r141 36 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=2.035
+ $X2=1.62 $Y2=2.035
r142 35 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.435 $Y=2.035
+ $X2=2.52 $Y2=2.035
r143 35 36 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.435 $Y=2.035
+ $X2=1.705 $Y2=2.035
r144 31 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=2.12
+ $X2=1.62 $Y2=2.035
r145 31 33 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.62 $Y=2.12
+ $X2=1.62 $Y2=2.815
r146 30 72 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.805 $Y=2.035
+ $X2=0.68 $Y2=2.035
r147 29 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=2.035
+ $X2=1.62 $Y2=2.035
r148 29 30 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.535 $Y=2.035
+ $X2=0.805 $Y2=2.035
r149 25 72 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.12
+ $X2=0.68 $Y2=2.035
r150 25 27 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=0.68 $Y=2.12
+ $X2=0.68 $Y2=2.815
r151 8 86 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.405
+ $Y=1.84 $X2=7.54 $Y2=1.985
r152 8 69 600 $w=1.7e-07 $l=7.94638e-07 $layer=licon1_PDIFF $count=1 $X=7.405
+ $Y=1.84 $X2=7.54 $Y2=2.57
r153 7 84 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.505
+ $Y=1.84 $X2=6.64 $Y2=1.985
r154 7 63 600 $w=1.7e-07 $l=7.94638e-07 $layer=licon1_PDIFF $count=1 $X=6.505
+ $Y=1.84 $X2=6.64 $Y2=2.57
r155 6 82 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=5.085
+ $Y=1.84 $X2=5.22 $Y2=2.115
r156 6 57 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.085
+ $Y=1.84 $X2=5.22 $Y2=2.815
r157 5 80 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.185
+ $Y=1.84 $X2=4.32 $Y2=1.985
r158 5 51 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=4.185
+ $Y=1.84 $X2=4.32 $Y2=2.4
r159 4 78 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=3.285
+ $Y=1.84 $X2=3.42 $Y2=2.115
r160 4 45 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.285
+ $Y=1.84 $X2=3.42 $Y2=2.815
r161 3 76 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=1.84 $X2=2.52 $Y2=2.115
r162 3 39 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=1.84 $X2=2.52 $Y2=2.815
r163 2 74 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.84 $X2=1.62 $Y2=2.115
r164 2 33 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.84 $X2=1.62 $Y2=2.815
r165 1 72 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.72 $Y2=2.115
r166 1 27 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.72 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_4%A_1213_368# 1 2 3 4 5 18 20 21 24 26 30 34
+ 38 40 44 48 49 50
r80 44 47 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=9.79 $Y=1.985
+ $X2=9.79 $Y2=2.815
r81 42 47 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=9.79 $Y=2.905 $X2=9.79
+ $Y2=2.815
r82 41 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.055 $Y=2.99
+ $X2=8.89 $Y2=2.99
r83 40 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.625 $Y=2.99
+ $X2=9.79 $Y2=2.905
r84 40 41 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=9.625 $Y=2.99
+ $X2=9.055 $Y2=2.99
r85 36 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.89 $Y=2.905
+ $X2=8.89 $Y2=2.99
r86 36 38 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=8.89 $Y=2.905
+ $X2=8.89 $Y2=2.225
r87 35 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.155 $Y=2.99
+ $X2=7.99 $Y2=2.99
r88 34 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.725 $Y=2.99
+ $X2=8.89 $Y2=2.99
r89 34 35 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.725 $Y=2.99
+ $X2=8.155 $Y2=2.99
r90 30 33 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=7.99 $Y=1.985
+ $X2=7.99 $Y2=2.815
r91 28 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.99 $Y=2.905
+ $X2=7.99 $Y2=2.99
r92 28 33 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=7.99 $Y=2.905 $X2=7.99
+ $Y2=2.815
r93 27 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.255 $Y=2.99
+ $X2=7.09 $Y2=2.99
r94 26 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.825 $Y=2.99
+ $X2=7.99 $Y2=2.99
r95 26 27 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=7.825 $Y=2.99
+ $X2=7.255 $Y2=2.99
r96 22 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.09 $Y=2.905
+ $X2=7.09 $Y2=2.99
r97 22 24 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=7.09 $Y=2.905 $X2=7.09
+ $Y2=2.405
r98 20 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.925 $Y=2.99
+ $X2=7.09 $Y2=2.99
r99 20 21 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=6.925 $Y=2.99
+ $X2=6.355 $Y2=2.99
r100 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.19 $Y=2.905
+ $X2=6.355 $Y2=2.99
r101 16 18 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=6.19 $Y=2.905
+ $X2=6.19 $Y2=2.405
r102 5 47 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.655
+ $Y=1.84 $X2=9.79 $Y2=2.815
r103 5 44 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.655
+ $Y=1.84 $X2=9.79 $Y2=1.985
r104 4 38 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=8.755
+ $Y=1.84 $X2=8.89 $Y2=2.225
r105 3 33 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.855
+ $Y=1.84 $X2=7.99 $Y2=2.815
r106 3 30 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.855
+ $Y=1.84 $X2=7.99 $Y2=1.985
r107 2 24 300 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=2 $X=6.955
+ $Y=1.84 $X2=7.09 $Y2=2.405
r108 1 18 300 $w=1.7e-07 $l=6.2438e-07 $layer=licon1_PDIFF $count=2 $X=6.065
+ $Y=1.84 $X2=6.19 $Y2=2.405
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_4%Y 1 2 3 4 5 6 7 22 28 30 34 40 42 43 45 48
+ 53 55 56 57 58 59 60 72 79 80
c91 34 0 1.44963e-19 $X=7.925 $Y=0.515
r92 79 80 4.36053 $w=6.58e-07 $l=6.5e-08 $layer=LI1_cond $X=9.36 $Y=0.68
+ $X2=9.425 $Y2=0.68
r93 71 72 9.09709 $w=6.58e-07 $l=8.5e-08 $layer=LI1_cond $X=8.785 $Y=0.68
+ $X2=8.7 $Y2=0.68
r94 59 79 0.181224 $w=6.58e-07 $l=1e-08 $layer=LI1_cond $X=9.35 $Y=0.68 $X2=9.36
+ $Y2=0.68
r95 59 76 0.181224 $w=6.58e-07 $l=1e-08 $layer=LI1_cond $X=9.35 $Y=0.68 $X2=9.34
+ $Y2=0.68
r96 59 60 14.5856 $w=3.18e-07 $l=4.05e-07 $layer=LI1_cond $X=9.435 $Y=0.51
+ $X2=9.84 $Y2=0.51
r97 59 80 0.360138 $w=3.18e-07 $l=1e-08 $layer=LI1_cond $X=9.435 $Y=0.51
+ $X2=9.425 $Y2=0.51
r98 58 76 8.3363 $w=6.58e-07 $l=4.6e-07 $layer=LI1_cond $X=8.88 $Y=0.68 $X2=9.34
+ $Y2=0.68
r99 58 71 1.72163 $w=6.58e-07 $l=9.5e-08 $layer=LI1_cond $X=8.88 $Y=0.68
+ $X2=8.785 $Y2=0.68
r100 51 53 5.88189 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.495 $Y=0.95
+ $X2=4.66 $Y2=0.95
r101 46 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.34 $Y=1.89
+ $X2=9.34 $Y2=1.805
r102 46 48 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=9.34 $Y=1.89
+ $X2=9.34 $Y2=1.985
r103 45 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.34 $Y=1.72
+ $X2=9.34 $Y2=1.805
r104 44 76 8.93547 $w=1.7e-07 $l=3.3e-07 $layer=LI1_cond $X=9.34 $Y=1.01
+ $X2=9.34 $Y2=0.68
r105 44 45 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=9.34 $Y=1.01
+ $X2=9.34 $Y2=1.72
r106 42 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.255 $Y=1.805
+ $X2=9.34 $Y2=1.805
r107 42 43 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=9.255 $Y=1.805
+ $X2=8.525 $Y2=1.805
r108 38 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.44 $Y=1.89
+ $X2=8.525 $Y2=1.805
r109 38 40 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=8.44 $Y=1.89
+ $X2=8.44 $Y2=1.985
r110 37 56 7.02821 $w=1.7e-07 $l=1.34629e-07 $layer=LI1_cond $X=8.01 $Y=0.925
+ $X2=7.885 $Y2=0.945
r111 37 72 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.01 $Y=0.925
+ $X2=8.7 $Y2=0.925
r112 32 56 0.00168595 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=7.885 $Y=0.84
+ $X2=7.885 $Y2=0.945
r113 32 34 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=7.885 $Y=0.84
+ $X2=7.885 $Y2=0.515
r114 31 55 5.63431 $w=2.25e-07 $l=1.52069e-07 $layer=LI1_cond $X=6.38 $Y=0.925
+ $X2=6.255 $Y2=0.985
r115 30 56 7.02821 $w=1.7e-07 $l=1.34629e-07 $layer=LI1_cond $X=7.76 $Y=0.925
+ $X2=7.885 $Y2=0.945
r116 30 31 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=7.76 $Y=0.925
+ $X2=6.38 $Y2=0.925
r117 26 55 0.966048 $w=2.5e-07 $l=1.45e-07 $layer=LI1_cond $X=6.255 $Y=0.84
+ $X2=6.255 $Y2=0.985
r118 26 28 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=6.255 $Y=0.84
+ $X2=6.255 $Y2=0.515
r119 25 53 28.6053 $w=2.78e-07 $l=6.95e-07 $layer=LI1_cond $X=5.355 $Y=0.99
+ $X2=4.66 $Y2=0.99
r120 22 55 5.63431 $w=2.25e-07 $l=1.27475e-07 $layer=LI1_cond $X=6.13 $Y=0.99
+ $X2=6.255 $Y2=0.985
r121 22 25 31.898 $w=2.78e-07 $l=7.75e-07 $layer=LI1_cond $X=6.13 $Y=0.99
+ $X2=5.355 $Y2=0.99
r122 7 48 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=9.205
+ $Y=1.84 $X2=9.34 $Y2=1.985
r123 6 40 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=8.305
+ $Y=1.84 $X2=8.44 $Y2=1.985
r124 5 71 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=8.645
+ $Y=0.37 $X2=8.785 $Y2=0.925
r125 5 71 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=8.645
+ $Y=0.37 $X2=8.785 $Y2=0.515
r126 4 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.785
+ $Y=0.37 $X2=7.925 $Y2=0.515
r127 3 55 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=6.075
+ $Y=0.37 $X2=6.215 $Y2=0.965
r128 3 28 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.075
+ $Y=0.37 $X2=6.215 $Y2=0.515
r129 2 25 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=5.215
+ $Y=0.37 $X2=5.355 $Y2=0.95
r130 1 51 182 $w=1.7e-07 $l=6.39453e-07 $layer=licon1_NDIFF $count=1 $X=4.37
+ $Y=0.37 $X2=4.495 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_4%A_34_74# 1 2 3 4 5 18 20 21 24 26 30 34 36
+ 37 40 41 43
r74 43 45 4.43516 $w=3.28e-07 $l=1.27e-07 $layer=LI1_cond $X=3.755 $Y=0.95
+ $X2=3.755 $Y2=1.077
r75 39 41 7.51706 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=0.975
+ $X2=3.06 $Y2=0.975
r76 39 40 7.51706 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=0.975
+ $X2=2.73 $Y2=0.975
r77 34 45 3.54104 $w=2.05e-07 $l=1.65e-07 $layer=LI1_cond $X=3.59 $Y=1.077
+ $X2=3.755 $Y2=1.077
r78 34 41 28.6741 $w=2.03e-07 $l=5.3e-07 $layer=LI1_cond $X=3.59 $Y=1.077
+ $X2=3.06 $Y2=1.077
r79 33 37 4.7579 $w=1.87e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=1.077
+ $X2=2.035 $Y2=1.077
r80 33 40 33.0022 $w=2.03e-07 $l=6.1e-07 $layer=LI1_cond $X=2.12 $Y=1.077
+ $X2=2.73 $Y2=1.077
r81 28 37 1.69765 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=2.035 $Y=0.975
+ $X2=2.035 $Y2=1.077
r82 28 30 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.035 $Y=0.975
+ $X2=2.035 $Y2=0.515
r83 27 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.26 $Y=1.095
+ $X2=1.135 $Y2=1.095
r84 26 37 4.7579 $w=1.87e-07 $l=9.35682e-08 $layer=LI1_cond $X=1.95 $Y=1.095
+ $X2=2.035 $Y2=1.077
r85 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.95 $Y=1.095
+ $X2=1.26 $Y2=1.095
r86 22 36 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=1.01
+ $X2=1.135 $Y2=1.095
r87 22 24 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.135 $Y=1.01
+ $X2=1.135 $Y2=0.515
r88 20 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.01 $Y=1.095
+ $X2=1.135 $Y2=1.095
r89 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.01 $Y=1.095
+ $X2=0.4 $Y2=1.095
r90 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.275 $Y=1.01
+ $X2=0.4 $Y2=1.095
r91 16 18 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.275 $Y=1.01
+ $X2=0.275 $Y2=0.515
r92 5 43 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=3.615
+ $Y=0.37 $X2=3.755 $Y2=0.95
r93 4 39 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=2.755
+ $Y=0.37 $X2=2.895 $Y2=0.95
r94 3 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.895
+ $Y=0.37 $X2=2.035 $Y2=0.515
r95 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.035
+ $Y=0.37 $X2=1.175 $Y2=0.515
r96 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.17
+ $Y=0.37 $X2=0.315 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_4%VGND 1 2 3 4 15 19 23 25 27 32 45 55 56 59
+ 62 66 72 74
r89 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r90 70 72 10.9168 $w=7.53e-07 $l=1.5e-07 $layer=LI1_cond $X=7.44 $Y=0.292
+ $X2=7.59 $Y2=0.292
r91 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r92 68 70 0.237631 $w=7.53e-07 $l=1.5e-08 $layer=LI1_cond $X=7.425 $Y=0.292
+ $X2=7.44 $Y2=0.292
r93 65 68 11.2479 $w=7.53e-07 $l=7.1e-07 $layer=LI1_cond $X=6.715 $Y=0.292
+ $X2=7.425 $Y2=0.292
r94 65 66 11.1544 $w=7.53e-07 $l=1.65e-07 $layer=LI1_cond $X=6.715 $Y=0.292
+ $X2=6.55 $Y2=0.292
r95 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r96 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r97 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r98 53 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r99 53 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r100 52 55 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r101 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r102 50 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.52 $Y=0 $X2=8.355
+ $Y2=0
r103 50 52 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.52 $Y=0 $X2=8.88
+ $Y2=0
r104 49 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r105 49 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r106 48 72 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.92 $Y=0 $X2=7.59
+ $Y2=0
r107 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r108 45 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.19 $Y=0 $X2=8.355
+ $Y2=0
r109 45 48 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.19 $Y=0 $X2=7.92
+ $Y2=0
r110 44 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r111 43 66 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=6.48 $Y=0 $X2=6.55
+ $Y2=0
r112 43 44 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r113 41 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r114 40 43 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=6.48
+ $Y2=0
r115 40 41 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r116 38 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.77 $Y=0 $X2=1.605
+ $Y2=0
r117 38 40 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.77 $Y=0 $X2=2.16
+ $Y2=0
r118 36 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r119 36 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r120 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r121 33 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.705
+ $Y2=0
r122 33 35 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=1.2
+ $Y2=0
r123 32 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.44 $Y=0 $X2=1.605
+ $Y2=0
r124 32 35 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r125 30 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r126 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r127 27 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.58 $Y=0 $X2=0.705
+ $Y2=0
r128 27 29 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.58 $Y=0 $X2=0.24
+ $Y2=0
r129 25 44 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.48 $Y2=0
r130 25 41 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=2.16 $Y2=0
r131 21 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.355 $Y=0.085
+ $X2=8.355 $Y2=0
r132 21 23 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=8.355 $Y=0.085
+ $X2=8.355 $Y2=0.55
r133 17 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=0.085
+ $X2=1.605 $Y2=0
r134 17 19 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.605 $Y=0.085
+ $X2=1.605 $Y2=0.675
r135 13 59 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0
r136 13 15 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.675
r137 4 23 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=8.215
+ $Y=0.37 $X2=8.355 $Y2=0.55
r138 3 68 121.333 $w=1.7e-07 $l=1.00598e-06 $layer=licon1_NDIFF $count=1
+ $X=6.505 $Y=0.37 $X2=7.425 $Y2=0.55
r139 3 65 121.333 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1
+ $X=6.505 $Y=0.37 $X2=6.715 $Y2=0.55
r140 2 19 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.465
+ $Y=0.37 $X2=1.605 $Y2=0.675
r141 1 15 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=0.605
+ $Y=0.37 $X2=0.745 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_MS__A311OI_4%A_465_74# 1 2 3 4 22 25 26 28 29
c37 28 0 1.0484e-19 $X=5.785 $Y=0.515
r38 28 29 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.785 $Y=0.515
+ $X2=5.62 $Y2=0.515
r39 24 26 4.02231 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.325 $Y=0.515
+ $X2=3.42 $Y2=0.515
r40 24 25 4.02231 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.325 $Y=0.515
+ $X2=3.23 $Y2=0.515
r41 22 25 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=2.56 $Y=0.475
+ $X2=3.23 $Y2=0.475
r42 20 22 4.02231 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.465 $Y=0.515
+ $X2=2.56 $Y2=0.515
r43 18 29 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=4.925 $Y=0.475
+ $X2=5.62 $Y2=0.475
r44 18 26 69.3771 $w=2.48e-07 $l=1.505e-06 $layer=LI1_cond $X=4.925 $Y=0.475
+ $X2=3.42 $Y2=0.475
r45 4 28 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.645
+ $Y=0.37 $X2=5.785 $Y2=0.515
r46 3 18 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.785
+ $Y=0.37 $X2=4.925 $Y2=0.515
r47 2 24 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.185
+ $Y=0.37 $X2=3.325 $Y2=0.515
r48 1 20 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.37 $X2=2.465 $Y2=0.515
.ends


* File: sky130_fd_sc_ms__a2bb2o_4.spice
* Created: Fri Aug 28 17:04:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a2bb2o_4.pex.spice"
.subckt sky130_fd_sc_ms__a2bb2o_4  VNB VPB A1_N A2_N B2 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_162_48#_M1000_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_162_48#_M1007_g N_X_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1007_d N_A_162_48#_M1010_g N_X_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1021_d N_A_162_48#_M1021_g N_X_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=1.36203 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1014 N_A_586_94#_M1014_d N_A1_N_M1014_g N_VGND_M1021_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.17797 NRD=0 NRS=46.872 M=1 R=4.26667
+ SA=75002.2 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1022 N_VGND_M1022_d N_A2_N_M1022_g N_A_586_94#_M1014_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.309101 AS=0.0896 PD=1.61391 PS=0.92 NRD=53.436 NRS=0 M=1 R=4.26667
+ SA=75002.6 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1017 N_A_162_48#_M1017_d N_A_586_94#_M1017_g N_VGND_M1022_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1961 AS=0.357399 PD=2.01 PS=1.86609 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_A_1009_74#_M1001_d N_B2_M1001_g N_A_162_48#_M1001_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1011 N_A_1009_74#_M1011_d N_B2_M1011_g N_A_162_48#_M1001_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1005 N_A_1009_74#_M1011_d N_B1_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1024 PD=0.92 PS=0.96 NRD=0 NRS=3.744 M=1 R=4.26667 SA=75001.1
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1008 N_A_1009_74#_M1008_d N_B1_M1008_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1696 AS=0.1024 PD=1.81 PS=0.96 NRD=0 NRS=3.744 M=1 R=4.26667 SA=75001.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1012 N_X_M1012_d N_A_162_48#_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1016 N_X_M1012_d N_A_162_48#_M1016_g N_VPWR_M1016_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90002 A=0.2016 P=2.6 MULT=1
MM1018 N_X_M1018_d N_A_162_48#_M1018_g N_VPWR_M1016_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1020 N_X_M1018_d N_A_162_48#_M1020_g N_VPWR_M1020_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2016 PD=1.39 PS=1.48 NRD=0 NRS=11.426 M=1 R=6.22222 SA=90001.5
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1002 A_586_368# N_A1_N_M1002_g N_VPWR_M1020_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1176 AS=0.2016 PD=1.33 PS=1.48 NRD=8.7862 NRS=2.6201 M=1 R=6.22222
+ SA=90002.1 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1006 N_A_586_94#_M1006_d N_A2_N_M1006_g A_586_368# VPB PSHORT L=0.18 W=1.12
+ AD=0.2912 AS=0.1176 PD=2.76 PS=1.33 NRD=0 NRS=8.7862 M=1 R=6.22222 SA=90002.4
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1003 N_A_162_48#_M1003_d N_A_586_94#_M1003_g N_A_820_392#_M1003_s VPB PSHORT
+ L=0.18 W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90002.4 A=0.18 P=2.36 MULT=1
MM1004 N_A_162_48#_M1003_d N_A_586_94#_M1004_g N_A_820_392#_M1004_s VPB PSHORT
+ L=0.18 W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.6 SB=90002 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_B2_M1009_g N_A_820_392#_M1004_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.1
+ SB=90001.5 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1009_d N_B2_M1013_g N_A_820_392#_M1013_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.5
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1015 N_VPWR_M1015_d N_B1_M1015_g N_A_820_392#_M1013_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90002
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1019 N_VPWR_M1015_d N_B1_M1019_g N_A_820_392#_M1019_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=5.55556 SA=90002.4
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX23_noxref VNB VPB NWDIODE A=14.0988 P=18.88
*
.include "sky130_fd_sc_ms__a2bb2o_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__a221o_1.pex.spice
* Created: Fri Aug 28 17:00:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A221O_1%A_148_260# 1 2 3 12 16 18 19 22 24 28 35 36
+ 38
r87 35 44 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.465
+ $X2=0.905 $Y2=1.63
r88 35 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.465
+ $X2=0.905 $Y2=1.3
r89 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.905
+ $Y=1.465 $X2=0.905 $Y2=1.465
r90 28 30 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.05 $Y=2.105
+ $X2=4.05 $Y2=2.815
r91 28 41 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=4.05 $Y=2.105
+ $X2=4.05 $Y2=1.285
r92 25 36 10.4332 $w=1.7e-07 $l=5.26498e-07 $layer=LI1_cond $X=2.86 $Y=1.2
+ $X2=2.42 $Y2=1.01
r93 24 41 2.83394 $w=3.53e-07 $l=8.5e-08 $layer=LI1_cond $X=4.037 $Y=1.2
+ $X2=4.037 $Y2=1.285
r94 24 38 6.33032 $w=3.53e-07 $l=1.95e-07 $layer=LI1_cond $X=4.037 $Y=1.2
+ $X2=4.037 $Y2=1.005
r95 24 25 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=3.86 $Y=1.2 $X2=2.86
+ $Y2=1.2
r96 20 36 1.73497 $w=4.4e-07 $l=2.2e-07 $layer=LI1_cond $X=2.64 $Y=1.01 $X2=2.42
+ $Y2=1.01
r97 20 22 12.834 $w=4.38e-07 $l=4.9e-07 $layer=LI1_cond $X=2.64 $Y=1.01 $X2=2.64
+ $Y2=0.52
r98 19 34 13.8043 $w=3.27e-07 $l=4.72345e-07 $layer=LI1_cond $X=1.205 $Y=1.095
+ $X2=0.972 $Y2=1.465
r99 18 36 10.4332 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.42 $Y=1.095
+ $X2=2.42 $Y2=1.01
r100 18 19 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=2.42 $Y=1.095
+ $X2=1.205 $Y2=1.095
r101 16 43 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.995 $Y=0.74
+ $X2=0.995 $Y2=1.3
r102 12 44 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.96 $Y=2.4
+ $X2=0.96 $Y2=1.63
r103 3 30 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.915
+ $Y=1.96 $X2=4.05 $Y2=2.815
r104 3 28 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.915
+ $Y=1.96 $X2=4.05 $Y2=2.105
r105 2 38 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.615 $X2=4.025 $Y2=1.005
r106 1 22 91 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=2 $X=2.445
+ $Y=0.395 $X2=2.64 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_1%A2 1 3 5 7 9 10
c42 3 0 1.75411e-19 $X=1.475 $Y=2.46
c43 1 0 1.57005e-19 $X=1.475 $Y=1.68
r44 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.46
+ $Y=1.515 $X2=1.46 $Y2=1.515
r45 10 15 5.89622 $w=4.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.46 $Y2=1.565
r46 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.01 $Y=1.11 $X2=2.01
+ $Y2=0.715
r47 6 14 56.4043 $w=2.82e-07 $l=4.04166e-07 $layer=POLY_cond $X=1.625 $Y=1.185
+ $X2=1.46 $Y2=1.515
r48 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.935 $Y=1.185
+ $X2=2.01 $Y2=1.11
r49 5 6 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=1.935 $Y=1.185
+ $X2=1.625 $Y2=1.185
r50 1 14 34.4858 $w=2.82e-07 $l=1.72337e-07 $layer=POLY_cond $X=1.475 $Y=1.68
+ $X2=1.46 $Y2=1.515
r51 1 3 303.194 $w=1.8e-07 $l=7.8e-07 $layer=POLY_cond $X=1.475 $Y=1.68
+ $X2=1.475 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_1%A1 3 7 9 16
c37 9 0 4.22091e-19 $X=2.16 $Y=1.665
c38 3 0 1.53462e-19 $X=1.925 $Y=2.46
r39 14 16 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=2.13 $Y=1.635
+ $X2=2.37 $Y2=1.635
r40 11 14 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.925 $Y=1.635
+ $X2=2.13 $Y2=1.635
r41 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.635 $X2=2.13 $Y2=1.635
r42 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.37 $Y=1.47
+ $X2=2.37 $Y2=1.635
r43 5 7 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.37 $Y=1.47 $X2=2.37
+ $Y2=0.715
r44 1 11 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.8
+ $X2=1.925 $Y2=1.635
r45 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.925 $Y=1.8 $X2=1.925
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_1%B1 3 7 9 12 13
c36 3 0 8.9675e-20 $X=2.895 $Y=2.46
r37 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.82 $Y=1.615
+ $X2=2.82 $Y2=1.78
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.82 $Y=1.615
+ $X2=2.82 $Y2=1.45
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.82
+ $Y=1.615 $X2=2.82 $Y2=1.615
r40 9 13 6.38276 $w=3.23e-07 $l=1.8e-07 $layer=LI1_cond $X=2.64 $Y=1.617
+ $X2=2.82 $Y2=1.617
r41 7 14 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=2.91 $Y=0.715
+ $X2=2.91 $Y2=1.45
r42 3 15 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=2.895 $Y=2.46
+ $X2=2.895 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_1%B2 3 7 9 12
c37 7 0 7.73749e-20 $X=3.345 $Y=2.46
c38 3 0 1.47272e-19 $X=3.27 $Y=0.715
r39 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.36 $Y=1.615
+ $X2=3.36 $Y2=1.78
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.36 $Y=1.615
+ $X2=3.36 $Y2=1.45
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.36
+ $Y=1.615 $X2=3.36 $Y2=1.615
r42 9 13 8.51035 $w=3.23e-07 $l=2.4e-07 $layer=LI1_cond $X=3.6 $Y=1.617 $X2=3.36
+ $Y2=1.617
r43 7 15 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=3.345 $Y=2.46
+ $X2=3.345 $Y2=1.78
r44 3 14 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=3.27 $Y=0.715
+ $X2=3.27 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_1%C1 4 5 7 10 15 16
c27 16 0 1.47272e-19 $X=4.03 $Y=0.34
c28 7 0 7.75124e-20 $X=3.825 $Y=2.46
r29 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.03
+ $Y=0.34 $X2=4.03 $Y2=0.34
r30 12 15 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=3.81 $Y=0.34
+ $X2=4.03 $Y2=0.34
r31 10 16 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=4.03 $Y=0.555
+ $X2=4.03 $Y2=0.34
r32 5 9 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.825 $Y=1.42 $X2=3.825
+ $Y2=1.33
r33 5 7 404.258 $w=1.8e-07 $l=1.04e-06 $layer=POLY_cond $X=3.825 $Y=1.42
+ $X2=3.825 $Y2=2.46
r34 4 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.81 $Y=0.935
+ $X2=3.81 $Y2=1.33
r35 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.81 $Y=0.505
+ $X2=3.81 $Y2=0.34
r36 1 4 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.81 $Y=0.505 $X2=3.81
+ $Y2=0.935
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_1%X 1 2 12 14 15 16 27 28
r21 27 28 5.7419 $w=7.73e-07 $l=1.65e-07 $layer=LI1_cond $X=0.512 $Y=1.985
+ $X2=0.512 $Y2=1.82
r22 15 16 5.71031 $w=7.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.512 $Y=2.405
+ $X2=0.512 $Y2=2.775
r23 14 15 5.71031 $w=7.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.512 $Y=2.035
+ $X2=0.512 $Y2=2.405
r24 14 27 0.771663 $w=7.73e-07 $l=5e-08 $layer=LI1_cond $X=0.512 $Y=2.035
+ $X2=0.512 $Y2=1.985
r25 9 12 7.17647 $w=7.78e-07 $l=4.68e-07 $layer=LI1_cond $X=0.312 $Y=0.74
+ $X2=0.78 $Y2=0.74
r26 7 9 5.04298 $w=3.75e-07 $l=3.9e-07 $layer=LI1_cond $X=0.312 $Y=1.13
+ $X2=0.312 $Y2=0.74
r27 7 28 21.205 $w=3.73e-07 $l=6.9e-07 $layer=LI1_cond $X=0.312 $Y=1.13
+ $X2=0.312 $Y2=1.82
r28 2 16 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.84 $X2=0.735 $Y2=2.815
r29 2 27 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.84 $X2=0.735 $Y2=1.985
r30 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.655
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_1%VPWR 1 2 9 15 17 19 24 34 35 38 41
r46 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r47 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r48 32 35 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r49 31 34 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r50 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 29 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=2.15 $Y2=3.33
r52 29 31 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r54 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 25 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.35 $Y=3.33
+ $X2=1.225 $Y2=3.33
r56 25 27 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.35 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 24 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=2.15 $Y2=3.33
r58 24 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=1.68 $Y2=3.33
r59 22 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r60 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 19 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.1 $Y=3.33
+ $X2=1.225 $Y2=3.33
r62 19 21 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.1 $Y=3.33 $X2=0.72
+ $Y2=3.33
r63 17 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r64 17 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 17 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r66 13 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=3.245
+ $X2=2.15 $Y2=3.33
r67 13 15 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.15 $Y=3.245
+ $X2=2.15 $Y2=2.475
r68 9 12 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=1.225 $Y=2.115
+ $X2=1.225 $Y2=2.815
r69 7 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=3.245
+ $X2=1.225 $Y2=3.33
r70 7 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=1.225 $Y=3.245
+ $X2=1.225 $Y2=2.815
r71 2 15 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=2.015
+ $Y=1.96 $X2=2.15 $Y2=2.475
r72 1 12 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.84 $X2=1.185 $Y2=2.815
r73 1 9 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.84 $X2=1.185 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_1%A_313_392# 1 2 7 9 11 18
c33 9 0 1.53462e-19 $X=1.7 $Y=2.815
r34 12 16 4.19273 $w=1.7e-07 $l=1.29904e-07 $layer=LI1_cond $X=1.785 $Y=2.055
+ $X2=1.66 $Y2=2.045
r35 11 18 5.03363 $w=1.7e-07 $l=1.69926e-07 $layer=LI1_cond $X=2.955 $Y=2.055
+ $X2=3.12 $Y2=2.045
r36 11 12 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=2.955 $Y=2.055
+ $X2=1.785 $Y2=2.055
r37 7 16 2.95044 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=1.66 $Y=2.14 $X2=1.66
+ $Y2=2.045
r38 7 9 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.66 $Y=2.14 $X2=1.66
+ $Y2=2.815
r39 2 18 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=2.985
+ $Y=1.96 $X2=3.12 $Y2=2.115
r40 1 16 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=1.565
+ $Y=1.96 $X2=1.7 $Y2=2.115
r41 1 9 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.565
+ $Y=1.96 $X2=1.7 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_1%A_509_392# 1 2 9 11 12 15
c23 15 0 1.54887e-19 $X=3.585 $Y=2.115
r24 15 18 38.8182 $w=1.98e-07 $l=7e-07 $layer=LI1_cond $X=3.585 $Y=2.115
+ $X2=3.585 $Y2=2.815
r25 13 18 4.99091 $w=1.98e-07 $l=9e-08 $layer=LI1_cond $X=3.585 $Y=2.905
+ $X2=3.585 $Y2=2.815
r26 11 13 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.485 $Y=2.99
+ $X2=3.585 $Y2=2.905
r27 11 12 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.485 $Y=2.99
+ $X2=2.785 $Y2=2.99
r28 7 12 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.645 $Y=2.905
+ $X2=2.785 $Y2=2.99
r29 7 9 17.6982 $w=2.78e-07 $l=4.3e-07 $layer=LI1_cond $X=2.645 $Y=2.905
+ $X2=2.645 $Y2=2.475
r30 2 18 400 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=3.435
+ $Y=1.96 $X2=3.585 $Y2=2.815
r31 2 15 400 $w=1.7e-07 $l=2.17428e-07 $layer=licon1_PDIFF $count=1 $X=3.435
+ $Y=1.96 $X2=3.585 $Y2=2.115
r32 1 9 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=2.545
+ $Y=1.96 $X2=2.67 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_MS__A221O_1%VGND 1 2 9 11 18 28 29 34 42 44
r43 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r44 41 42 12.4865 $w=9.23e-07 $l=1.7e-07 $layer=LI1_cond $X=1.795 $Y=0.377
+ $X2=1.965 $Y2=0.377
r45 38 41 1.51676 $w=9.23e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=0.377
+ $X2=1.795 $Y2=0.377
r46 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r47 36 38 6.19892 $w=9.23e-07 $l=4.7e-07 $layer=LI1_cond $X=1.21 $Y=0.377
+ $X2=1.68 $Y2=0.377
r48 33 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r49 32 36 0.131892 $w=9.23e-07 $l=1e-08 $layer=LI1_cond $X=1.2 $Y=0.377 $X2=1.21
+ $Y2=0.377
r50 32 34 12.2887 $w=9.23e-07 $l=1.55e-07 $layer=LI1_cond $X=1.2 $Y=0.377
+ $X2=1.045 $Y2=0.377
r51 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r52 29 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r53 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r54 26 44 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.69 $Y=0 $X2=3.505
+ $Y2=0
r55 26 28 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.69 $Y=0 $X2=4.08
+ $Y2=0
r56 25 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r57 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r58 21 24 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r59 21 42 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=1.965
+ $Y2=0
r60 18 44 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.32 $Y=0 $X2=3.505
+ $Y2=0
r61 18 24 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.32 $Y=0 $X2=3.12
+ $Y2=0
r62 16 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r63 15 34 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.045
+ $Y2=0
r64 15 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r65 11 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r66 11 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r67 11 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r68 7 44 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.505 $Y=0.085
+ $X2=3.505 $Y2=0
r69 7 9 13.549 $w=3.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.505 $Y=0.085
+ $X2=3.505 $Y2=0.52
r70 2 9 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=3.345
+ $Y=0.395 $X2=3.505 $Y2=0.52
r71 1 41 182 $w=1.7e-07 $l=8.64147e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.795 $Y2=0.675
r72 1 36 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.21 $Y2=0.675
.ends


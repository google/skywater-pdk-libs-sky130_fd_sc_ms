* File: sky130_fd_sc_ms__mux4_2.spice
* Created: Wed Sep  2 12:12:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__mux4_2.pex.spice"
.subckt sky130_fd_sc_ms__mux4_2  VNB VPB S0 A1 A0 A3 A2 S1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* S1	S1
* A2	A2
* A3	A3
* A0	A0
* A1	A1
* S0	S0
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_S0_M1000_g N_A_31_94#_M1000_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.172012 AS=0.1824 PD=1.18261 PS=1.85 NRD=48.276 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75005.8 A=0.096 P=1.58 MULT=1
MM1013 A_255_74# N_A1_M1013_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.198888 PD=0.98 PS=1.36739 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.8
+ SB=75005.1 A=0.111 P=1.78 MULT=1
MM1011 N_A_333_74#_M1011_d N_S0_M1011_g A_255_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.2664 AS=0.0888 PD=1.46 PS=0.98 NRD=44.592 NRS=10.536 M=1 R=4.93333
+ SA=75001.2 SB=75004.7 A=0.111 P=1.78 MULT=1
MM1014 A_507_74# N_A_31_94#_M1014_g N_A_333_74#_M1011_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2886 AS=0.2664 PD=1.52 PS=1.46 NRD=54.324 NRS=26.748 M=1 R=4.93333
+ SA=75002.1 SB=75003.8 A=0.111 P=1.78 MULT=1
MM1024 N_VGND_M1024_d N_A0_M1024_g A_507_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1998
+ AS=0.2886 PD=1.28 PS=1.52 NRD=7.296 NRS=54.324 M=1 R=4.93333 SA=75003
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1020 A_831_74# N_A3_M1020_g N_VGND_M1024_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.1998 PD=0.98 PS=1.28 NRD=10.536 NRS=34.86 M=1 R=4.93333 SA=75003.7
+ SB=75002.2 A=0.111 P=1.78 MULT=1
MM1016 N_A_909_74#_M1016_d N_S0_M1016_g A_831_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1998 AS=0.0888 PD=1.28 PS=0.98 NRD=27.564 NRS=10.536 M=1 R=4.93333
+ SA=75004.1 SB=75001.8 A=0.111 P=1.78 MULT=1
MM1004 A_1047_74# N_A_31_94#_M1004_g N_A_909_74#_M1016_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2886 AS=0.1998 PD=1.52 PS=1.28 NRD=54.324 NRS=14.592 M=1 R=4.93333
+ SA=75004.8 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_A2_M1012_g A_1047_74# VNB NLOWVT L=0.15 W=0.74 AD=0.2072
+ AS=0.2886 PD=2.04 PS=1.52 NRD=0 NRS=54.324 M=1 R=4.93333 SA=75005.7 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1010 N_A_1429_74#_M1010_d N_S1_M1010_g N_A_909_74#_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.151475 AS=0.2072 PD=1.325 PS=2.04 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1007 N_A_333_74#_M1007_d N_A_1500_94#_M1007_g N_A_1429_74#_M1010_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.151475 PD=2.05 PS=1.325 NRD=0 NRS=24.264 M=1
+ R=4.93333 SA=75000.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_S1_M1009_g N_A_1500_94#_M1009_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.232858 AS=0.276725 PD=1.37275 PS=2.15 NRD=86.712 NRS=26.244 M=1 R=4.26667
+ SA=75000.4 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1022 N_X_M1022_d N_A_1429_74#_M1022_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.269242 PD=1.02 PS=1.58725 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1025 N_X_M1022_d N_A_1429_74#_M1025_g N_VGND_M1025_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VPWR_M1001_d N_S0_M1001_g N_A_31_94#_M1001_s VPB PSHORT L=0.18 W=1
+ AD=0.21 AS=0.28 PD=1.42 PS=2.56 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90005.6 A=0.18 P=2.36 MULT=1
MM1026 A_267_392# N_A1_M1026_g N_VPWR_M1001_d VPB PSHORT L=0.18 W=1 AD=0.435
+ AS=0.21 PD=1.87 PS=1.42 NRD=74.8403 NRS=18.715 M=1 R=5.55556 SA=90000.8
+ SB=90005 A=0.18 P=2.36 MULT=1
MM1023 N_A_333_74#_M1023_d N_A_31_94#_M1023_g A_267_392# VPB PSHORT L=0.18 W=1
+ AD=0.27 AS=0.435 PD=1.54 PS=1.87 NRD=26.5753 NRS=74.8403 M=1 R=5.55556
+ SA=90001.8 SB=90004 A=0.18 P=2.36 MULT=1
MM1008 A_621_392# N_S0_M1008_g N_A_333_74#_M1023_d VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.27 PD=1.24 PS=1.54 NRD=12.7853 NRS=24.6053 M=1 R=5.55556 SA=90002.6
+ SB=90003.3 A=0.18 P=2.36 MULT=1
MM1017 N_VPWR_M1017_d N_A0_M1017_g A_621_392# VPB PSHORT L=0.18 W=1 AD=0.255
+ AS=0.12 PD=1.51 PS=1.24 NRD=22.6353 NRS=12.7853 M=1 R=5.55556 SA=90003
+ SB=90002.9 A=0.18 P=2.36 MULT=1
MM1018 A_843_392# N_A3_M1018_g N_VPWR_M1017_d VPB PSHORT L=0.18 W=1 AD=0.345
+ AS=0.255 PD=1.69 PS=1.51 NRD=57.1103 NRS=22.6353 M=1 R=5.55556 SA=90003.7
+ SB=90002.2 A=0.18 P=2.36 MULT=1
MM1005 N_A_909_74#_M1005_d N_A_31_94#_M1005_g A_843_392# VPB PSHORT L=0.18 W=1
+ AD=0.255 AS=0.345 PD=1.51 PS=1.69 NRD=22.6353 NRS=57.1103 M=1 R=5.55556
+ SA=90004.5 SB=90001.3 A=0.18 P=2.36 MULT=1
MM1002 A_1155_392# N_S0_M1002_g N_A_909_74#_M1005_d VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.255 PD=1.24 PS=1.51 NRD=12.7853 NRS=22.6353 M=1 R=5.55556
+ SA=90005.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1019 N_VPWR_M1019_d N_A2_M1019_g A_1155_392# VPB PSHORT L=0.18 W=1 AD=0.28
+ AS=0.12 PD=2.56 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556 SA=90005.6 SB=90000.2
+ A=0.18 P=2.36 MULT=1
MM1003 N_A_1429_74#_M1003_d N_S1_M1003_g N_A_333_74#_M1003_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.305 PD=1.27 PS=2.61 NRD=0 NRS=1.9503 M=1 R=5.55556
+ SA=90000.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1006 N_A_909_74#_M1006_d N_A_1500_94#_M1006_g N_A_1429_74#_M1003_d VPB PSHORT
+ L=0.18 W=1 AD=0.275 AS=0.135 PD=2.55 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.7 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1027 N_VPWR_M1027_d N_S1_M1027_g N_A_1500_94#_M1027_s VPB PSHORT L=0.18 W=1
+ AD=0.348113 AS=0.41 PD=1.7217 PS=2.82 NRD=85.0252 NRS=25.5903 M=1 R=5.55556
+ SA=90000.3 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1015 N_X_M1015_d N_A_1429_74#_M1015_g N_VPWR_M1027_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.389887 PD=1.39 PS=1.9283 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1021 N_X_M1015_d N_A_1429_74#_M1021_g N_VPWR_M1021_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.308 PD=1.39 PS=2.79 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX28_noxref VNB VPB NWDIODE A=20.2119 P=25.8
c_1339 A_507_74# 0 1.87351e-19 $X=2.535 $Y=0.37
*
.include "sky130_fd_sc_ms__mux4_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__bufinv_16.spice
* Created: Fri Aug 28 17:16:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__bufinv_16.pex.spice"
.subckt sky130_fd_sc_ms__bufinv_16  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_A_27_74#_M1000_d N_A_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1258 PD=2.05 PS=1.08 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75011.2 A=0.111 P=1.78 MULT=1
MM1035 N_A_27_74#_M1035_d N_A_M1035_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1258 PD=1.02 PS=1.08 NRD=0 NRS=9.72 M=1 R=4.93333 SA=75000.7
+ SB=75010.7 A=0.111 P=1.78 MULT=1
MM1047 N_A_27_74#_M1035_d N_A_M1047_g N_VGND_M1047_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75010.3 A=0.111 P=1.78 MULT=1
MM1011 N_A_384_74#_M1011_d N_A_27_74#_M1011_g N_VGND_M1047_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75009.9 A=0.111 P=1.78 MULT=1
MM1015 N_A_384_74#_M1011_d N_A_27_74#_M1015_g N_VGND_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002
+ SB=75009.4 A=0.111 P=1.78 MULT=1
MM1018 N_A_384_74#_M1018_d N_A_27_74#_M1018_g N_VGND_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75009 A=0.111 P=1.78 MULT=1
MM1026 N_A_384_74#_M1018_d N_A_27_74#_M1026_g N_VGND_M1026_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.9 SB=75008.6 A=0.111 P=1.78 MULT=1
MM1048 N_A_384_74#_M1048_d N_A_27_74#_M1048_g N_VGND_M1026_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75003.3 SB=75008.1 A=0.111 P=1.78 MULT=1
MM1049 N_A_384_74#_M1048_d N_A_27_74#_M1049_g N_VGND_M1049_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.8 SB=75007.6 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1049_s N_A_384_74#_M1003_g N_Y_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75004.3
+ SB=75007.2 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_384_74#_M1007_g N_Y_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.7
+ SB=75006.7 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1007_d N_A_384_74#_M1013_g N_Y_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.1
+ SB=75006.3 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1021_d N_A_384_74#_M1021_g N_Y_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.6
+ SB=75005.9 A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1021_d N_A_384_74#_M1022_g N_Y_M1022_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75006.1
+ SB=75005.4 A=0.111 P=1.78 MULT=1
MM1023 N_VGND_M1023_d N_A_384_74#_M1023_g N_Y_M1022_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75006.5
+ SB=75004.9 A=0.111 P=1.78 MULT=1
MM1027 N_VGND_M1023_d N_A_384_74#_M1027_g N_Y_M1027_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75007
+ SB=75004.4 A=0.111 P=1.78 MULT=1
MM1028 N_VGND_M1028_d N_A_384_74#_M1028_g N_Y_M1027_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75007.4
+ SB=75004 A=0.111 P=1.78 MULT=1
MM1032 N_VGND_M1028_d N_A_384_74#_M1032_g N_Y_M1032_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75007.9
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1036 N_VGND_M1036_d N_A_384_74#_M1036_g N_Y_M1032_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75008.4
+ SB=75003.1 A=0.111 P=1.78 MULT=1
MM1038 N_VGND_M1036_d N_A_384_74#_M1038_g N_Y_M1038_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75008.9
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1039 N_VGND_M1039_d N_A_384_74#_M1039_g N_Y_M1038_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75009.3
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1041 N_VGND_M1039_d N_A_384_74#_M1041_g N_Y_M1041_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75009.8
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1042 N_VGND_M1042_d N_A_384_74#_M1042_g N_Y_M1041_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75010.2
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1044 N_VGND_M1042_d N_A_384_74#_M1044_g N_Y_M1044_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75010.7
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1046 N_VGND_M1046_d N_A_384_74#_M1046_g N_Y_M1044_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.1036 PD=2.19 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75011.1
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_A_27_74#_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90011.2 A=0.2016 P=2.6 MULT=1
MM1002 N_VPWR_M1001_d N_A_M1002_g N_A_27_74#_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90010.7 A=0.2016 P=2.6 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g N_A_27_74#_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90010.3 A=0.2016 P=2.6 MULT=1
MM1009 N_A_384_74#_M1009_d N_A_27_74#_M1009_g N_VPWR_M1005_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1624 AS=0.1512 PD=1.41 PS=1.39 NRD=2.6201 NRS=0 M=1 R=6.22222
+ SA=90001.5 SB=90009.8 A=0.2016 P=2.6 MULT=1
MM1016 N_A_384_74#_M1009_d N_A_27_74#_M1016_g N_VPWR_M1016_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1624 AS=0.1512 PD=1.41 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90009.3 A=0.2016 P=2.6 MULT=1
MM1019 N_A_384_74#_M1019_d N_A_27_74#_M1019_g N_VPWR_M1016_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90002.5 SB=90008.9 A=0.2016 P=2.6 MULT=1
MM1025 N_A_384_74#_M1019_d N_A_27_74#_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90002.9 SB=90008.4 A=0.2016 P=2.6 MULT=1
MM1029 N_A_384_74#_M1029_d N_A_27_74#_M1029_g N_VPWR_M1025_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90003.4 SB=90008 A=0.2016 P=2.6 MULT=1
MM1033 N_A_384_74#_M1029_d N_A_27_74#_M1033_g N_VPWR_M1033_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90003.8 SB=90007.5 A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1004_d N_A_384_74#_M1004_g N_VPWR_M1033_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.3
+ SB=90007.1 A=0.2016 P=2.6 MULT=1
MM1006 N_Y_M1004_d N_A_384_74#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.7
+ SB=90006.6 A=0.2016 P=2.6 MULT=1
MM1008 N_Y_M1008_d N_A_384_74#_M1008_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90005.2
+ SB=90006.2 A=0.2016 P=2.6 MULT=1
MM1010 N_Y_M1008_d N_A_384_74#_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90005.6
+ SB=90005.7 A=0.2016 P=2.6 MULT=1
MM1012 N_Y_M1012_d N_A_384_74#_M1012_g N_VPWR_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90006.1
+ SB=90005.3 A=0.2016 P=2.6 MULT=1
MM1014 N_Y_M1012_d N_A_384_74#_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90006.5
+ SB=90004.8 A=0.2016 P=2.6 MULT=1
MM1017 N_Y_M1017_d N_A_384_74#_M1017_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90007
+ SB=90004.4 A=0.2016 P=2.6 MULT=1
MM1020 N_Y_M1017_d N_A_384_74#_M1020_g N_VPWR_M1020_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90007.4
+ SB=90003.9 A=0.2016 P=2.6 MULT=1
MM1024 N_Y_M1024_d N_A_384_74#_M1024_g N_VPWR_M1020_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90007.9
+ SB=90003.5 A=0.2016 P=2.6 MULT=1
MM1030 N_Y_M1024_d N_A_384_74#_M1030_g N_VPWR_M1030_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90008.3
+ SB=90003 A=0.2016 P=2.6 MULT=1
MM1031 N_Y_M1031_d N_A_384_74#_M1031_g N_VPWR_M1030_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90008.8
+ SB=90002.5 A=0.2016 P=2.6 MULT=1
MM1034 N_Y_M1031_d N_A_384_74#_M1034_g N_VPWR_M1034_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90009.3
+ SB=90002.1 A=0.2016 P=2.6 MULT=1
MM1037 N_Y_M1037_d N_A_384_74#_M1037_g N_VPWR_M1034_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90009.8
+ SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1040 N_Y_M1037_d N_A_384_74#_M1040_g N_VPWR_M1040_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1568 PD=1.39 PS=1.4 NRD=0 NRS=0 M=1 R=6.22222 SA=90010.2
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1043 N_Y_M1043_d N_A_384_74#_M1043_g N_VPWR_M1040_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1736 AS=0.1568 PD=1.43 PS=1.4 NRD=6.1464 NRS=0.8668 M=1 R=6.22222
+ SA=90010.7 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1045 N_Y_M1043_d N_A_384_74#_M1045_g N_VPWR_M1045_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1736 AS=0.3136 PD=1.43 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90011.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX50_noxref VNB VPB NWDIODE A=23.0268 P=28.48
*
.include "sky130_fd_sc_ms__bufinv_16.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__ebufn_4.spice
* Created: Fri Aug 28 17:32:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__ebufn_4.pex.spice"
.subckt sky130_fd_sc_ms__ebufn_4  VNB VPB A TE_B VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* TE_B	TE_B
* A	A
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_27_368#_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1011 N_A_208_74#_M1011_d N_TE_B_M1011_g N_VGND_M1004_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_208_74#_M1007_g N_A_378_74#_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2072 PD=1.02 PS=2.04 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75003.2 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1007_d N_A_208_74#_M1008_g N_A_378_74#_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75002.8 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_A_208_74#_M1009_g N_A_378_74#_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75002.4 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1009_d N_A_208_74#_M1015_g N_A_378_74#_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1005 N_A_378_74#_M1015_s N_A_27_368#_M1005_g N_Z_M1005_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.9 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1012 N_A_378_74#_M1012_d N_A_27_368#_M1012_g N_Z_M1005_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1014 N_A_378_74#_M1012_d N_A_27_368#_M1014_g N_Z_M1014_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.111 PD=1.02 PS=1.04 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1018 N_A_378_74#_M1018_d N_A_27_368#_M1018_g N_Z_M1014_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2035 AS=0.111 PD=2.03 PS=1.04 NRD=0 NRS=3.24 M=1 R=4.93333
+ SA=75003.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_A_27_368#_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1652 AS=0.3136 PD=1.415 PS=2.8 NRD=0.8668 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1001 N_A_208_74#_M1001_d N_TE_B_M1001_g N_VPWR_M1006_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.1652 PD=2.8 PS=1.415 NRD=0 NRS=1.7533 M=1 R=6.22222
+ SA=90000.7 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1013 N_VPWR_M1013_d N_TE_B_M1013_g N_A_348_368#_M1013_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003.3 A=0.2016 P=2.6 MULT=1
MM1016 N_VPWR_M1013_d N_TE_B_M1016_g N_A_348_368#_M1016_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90002.9 A=0.2016 P=2.6 MULT=1
MM1017 N_VPWR_M1017_d N_TE_B_M1017_g N_A_348_368#_M1016_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.1 SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1019 N_VPWR_M1017_d N_TE_B_M1019_g N_A_348_368#_M1019_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.5 SB=90002 A=0.2016 P=2.6 MULT=1
MM1000 N_Z_M1000_d N_A_27_368#_M1000_g N_A_348_368#_M1019_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1002 N_Z_M1000_d N_A_27_368#_M1002_g N_A_348_368#_M1002_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90002.4 SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1003 N_Z_M1003_d N_A_27_368#_M1003_g N_A_348_368#_M1002_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90002.9 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1010 N_Z_M1003_d N_A_27_368#_M1010_g N_A_348_368#_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.308 PD=1.39 PS=2.79 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.3
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ms__ebufn_4.pxi.spice"
*
.ends
*
*

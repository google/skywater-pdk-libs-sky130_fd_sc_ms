* File: sky130_fd_sc_ms__a21bo_2.pex.spice
* Created: Wed Sep  2 11:50:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A21BO_2%B1_N 3 5 7 8 12 15
r30 14 15 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=0.51 $Y=1.385
+ $X2=0.65 $Y2=1.385
r31 11 14 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.345 $Y=1.385
+ $X2=0.51 $Y2=1.385
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.345
+ $Y=1.385 $X2=0.345 $Y2=1.385
r33 8 12 3.27045 $w=3.68e-07 $l=1.05e-07 $layer=LI1_cond $X=0.24 $Y=1.365
+ $X2=0.345 $Y2=1.365
r34 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.65 $Y=1.22
+ $X2=0.65 $Y2=1.385
r35 5 7 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.65 $Y=1.22 $X2=0.65
+ $Y2=0.835
r36 1 14 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.55
+ $X2=0.51 $Y2=1.385
r37 1 3 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=0.51 $Y=1.55 $X2=0.51
+ $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_2%A_187_244# 1 2 9 11 13 16 18 20 21 22 26 29
+ 34 36 37
r97 39 40 61.307 $w=2.28e-07 $l=2.9e-07 $layer=POLY_cond $X=1.185 $Y=1.37
+ $X2=1.475 $Y2=1.37
r98 34 42 19.0263 $w=2.28e-07 $l=9e-08 $layer=POLY_cond $X=1.525 $Y=1.37
+ $X2=1.615 $Y2=1.37
r99 34 40 10.5702 $w=2.28e-07 $l=5e-08 $layer=POLY_cond $X=1.525 $Y=1.37
+ $X2=1.475 $Y2=1.37
r100 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.525
+ $Y=1.385 $X2=1.525 $Y2=1.385
r101 27 37 3.70735 $w=2.5e-07 $l=1.06325e-07 $layer=LI1_cond $X=2.645 $Y=0.92
+ $X2=2.597 $Y2=1.005
r102 27 29 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=2.645 $Y=0.92
+ $X2=2.645 $Y2=0.515
r103 26 36 21.6337 $w=2.9e-07 $l=5.41249e-07 $layer=LI1_cond $X=2.47 $Y=1.76
+ $X2=2.305 $Y2=2.225
r104 25 37 3.70735 $w=2.5e-07 $l=1.64085e-07 $layer=LI1_cond $X=2.47 $Y=1.09
+ $X2=2.597 $Y2=1.005
r105 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.47 $Y=1.09
+ $X2=2.47 $Y2=1.76
r106 22 33 16.7365 $w=2.77e-07 $l=4.64586e-07 $layer=LI1_cond $X=1.735 $Y=1.005
+ $X2=1.547 $Y2=1.385
r107 21 37 2.76166 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.385 $Y=1.005
+ $X2=2.597 $Y2=1.005
r108 21 22 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.385 $Y=1.005
+ $X2=1.735 $Y2=1.005
r109 18 42 12.5943 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.615 $Y=1.22
+ $X2=1.615 $Y2=1.37
r110 18 20 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.615 $Y=1.22
+ $X2=1.615 $Y2=0.74
r111 14 40 8.39207 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=1.475 $Y=1.55
+ $X2=1.475 $Y2=1.37
r112 14 16 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.475 $Y=1.55
+ $X2=1.475 $Y2=2.4
r113 11 39 12.5943 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.185 $Y=1.22
+ $X2=1.185 $Y2=1.37
r114 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.185 $Y=1.22
+ $X2=1.185 $Y2=0.74
r115 7 39 33.8246 $w=2.28e-07 $l=1.6e-07 $layer=POLY_cond $X=1.025 $Y=1.37
+ $X2=1.185 $Y2=1.37
r116 7 9 400.371 $w=1.8e-07 $l=1.03e-06 $layer=POLY_cond $X=1.025 $Y=1.37
+ $X2=1.025 $Y2=2.4
r117 2 36 300 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_PDIFF $count=2 $X=2.095
+ $Y=1.96 $X2=2.22 $Y2=2.225
r118 1 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.505
+ $Y=0.37 $X2=2.645 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_2%A_32_368# 1 2 9 13 15 17 18 19 22 24 25 27
+ 28 30 31 33 35
c98 13 0 1.81275e-19 $X=2.445 $Y=1.82
r99 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.065
+ $Y=1.425 $X2=2.065 $Y2=1.425
r100 30 37 19.1478 $w=3.24e-07 $l=5.57333e-07 $layer=LI1_cond $X=1.707 $Y=1.89
+ $X2=1.91 $Y2=1.425
r101 30 31 18.9357 $w=2.03e-07 $l=3.5e-07 $layer=LI1_cond $X=1.707 $Y=1.89
+ $X2=1.707 $Y2=2.24
r102 29 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=2.325
+ $X2=0.765 $Y2=2.325
r103 28 31 6.89401 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=1.605 $Y=2.325
+ $X2=1.707 $Y2=2.24
r104 28 29 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.605 $Y=2.325
+ $X2=0.85 $Y2=2.325
r105 27 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=2.24
+ $X2=0.765 $Y2=2.325
r106 26 33 11.8412 $w=3.4e-07 $l=4.31799e-07 $layer=LI1_cond $X=0.765 $Y=1.01
+ $X2=0.435 $Y2=0.775
r107 26 27 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=0.765 $Y=1.01
+ $X2=0.765 $Y2=2.24
r108 24 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=2.325
+ $X2=0.765 $Y2=2.325
r109 24 25 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.68 $Y=2.325
+ $X2=0.45 $Y2=2.325
r110 20 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.285 $Y=2.24
+ $X2=0.45 $Y2=2.325
r111 20 22 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=0.285 $Y=2.24
+ $X2=0.285 $Y2=1.985
r112 17 38 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=2.355 $Y=1.425
+ $X2=2.065 $Y2=1.425
r113 17 18 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.355 $Y=1.425
+ $X2=2.43 $Y2=1.425
r114 13 19 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.445 $Y=1.82
+ $X2=2.445 $Y2=1.73
r115 13 15 248.774 $w=1.8e-07 $l=6.4e-07 $layer=POLY_cond $X=2.445 $Y=1.82
+ $X2=2.445 $Y2=2.46
r116 11 18 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.43 $Y=1.59
+ $X2=2.43 $Y2=1.425
r117 11 19 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=2.43 $Y=1.59
+ $X2=2.43 $Y2=1.73
r118 7 18 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.43 $Y=1.26
+ $X2=2.43 $Y2=1.425
r119 7 9 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.43 $Y=1.26 $X2=2.43
+ $Y2=0.74
r120 2 22 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.16
+ $Y=1.84 $X2=0.285 $Y2=1.985
r121 1 33 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=0.31
+ $Y=0.56 $X2=0.435 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_2%A1 3 7 9 12 13
c40 13 0 1.81275e-19 $X=2.88 $Y=1.425
c41 12 0 2.3968e-19 $X=2.88 $Y=1.425
c42 7 0 1.3104e-19 $X=2.895 $Y=2.46
r43 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.88 $Y=1.425
+ $X2=2.88 $Y2=1.59
r44 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.88 $Y=1.425
+ $X2=2.88 $Y2=1.26
r45 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.88
+ $Y=1.425 $X2=2.88 $Y2=1.425
r46 9 13 5.6286 $w=5.08e-07 $l=2.4e-07 $layer=LI1_cond $X=2.98 $Y=1.665 $X2=2.98
+ $Y2=1.425
r47 7 15 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=2.895 $Y=2.46
+ $X2=2.895 $Y2=1.59
r48 3 14 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.86 $Y=0.74 $X2=2.86
+ $Y2=1.26
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_2%A2 3 7 9 15
c26 9 0 2.30057e-19 $X=3.6 $Y=1.665
r27 13 15 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.345 $Y=1.615
+ $X2=3.57 $Y2=1.615
r28 11 13 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.33 $Y=1.615
+ $X2=3.345 $Y2=1.615
r29 9 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.615 $X2=3.57 $Y2=1.615
r30 5 13 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.345 $Y=1.78
+ $X2=3.345 $Y2=1.615
r31 5 7 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=3.345 $Y=1.78
+ $X2=3.345 $Y2=2.46
r32 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.33 $Y=1.45
+ $X2=3.33 $Y2=1.615
r33 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.33 $Y=1.45 $X2=3.33
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_2%VPWR 1 2 3 12 16 20 22 24 29 34 41 42 45 48
+ 51
r58 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r59 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 42 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r62 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r63 39 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.205 $Y=3.33
+ $X2=3.08 $Y2=3.33
r64 39 41 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.205 $Y=3.33
+ $X2=3.6 $Y2=3.33
r65 38 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r66 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r67 35 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=3.33
+ $X2=1.7 $Y2=3.33
r68 35 37 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.865 $Y=3.33
+ $X2=2.64 $Y2=3.33
r69 34 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.955 $Y=3.33
+ $X2=3.08 $Y2=3.33
r70 34 37 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.955 $Y=3.33
+ $X2=2.64 $Y2=3.33
r71 33 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r72 33 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r73 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r74 30 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=0.8 $Y2=3.33
r75 30 32 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=1.2 $Y2=3.33
r76 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.535 $Y=3.33
+ $X2=1.7 $Y2=3.33
r77 29 32 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.535 $Y=3.33
+ $X2=1.2 $Y2=3.33
r78 27 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r79 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r80 24 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.8 $Y2=3.33
r81 24 26 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.24 $Y2=3.33
r82 22 38 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r83 22 49 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r84 18 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.08 $Y2=3.33
r85 18 20 24.6623 $w=2.48e-07 $l=5.35e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.08 $Y2=2.71
r86 14 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=3.245 $X2=1.7
+ $Y2=3.33
r87 14 16 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=1.7 $Y=3.245 $X2=1.7
+ $Y2=2.745
r88 10 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=3.245 $X2=0.8
+ $Y2=3.33
r89 10 12 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=0.8 $Y=3.245 $X2=0.8
+ $Y2=2.745
r90 3 20 600 $w=1.7e-07 $l=8.14709e-07 $layer=licon1_PDIFF $count=1 $X=2.985
+ $Y=1.96 $X2=3.12 $Y2=2.71
r91 2 16 600 $w=1.7e-07 $l=9.70155e-07 $layer=licon1_PDIFF $count=1 $X=1.565
+ $Y=1.84 $X2=1.7 $Y2=2.745
r92 1 12 600 $w=1.7e-07 $l=1.00001e-06 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.84 $X2=0.8 $Y2=2.745
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_2%X 1 2 7 8 12 14
r35 14 17 13.9908 $w=3.27e-07 $l=3.75e-07 $layer=LI1_cond $X=1.292 $Y=0.925
+ $X2=1.292 $Y2=0.55
r36 9 12 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=1.105 $Y=1.945
+ $X2=1.25 $Y2=1.945
r37 8 9 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.105 $Y=1.82
+ $X2=1.105 $Y2=1.945
r38 7 14 7.09126 $w=3.27e-07 $l=2.37643e-07 $layer=LI1_cond $X=1.105 $Y=1.04
+ $X2=1.292 $Y2=0.925
r39 7 8 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=1.105 $Y=1.04
+ $X2=1.105 $Y2=1.82
r40 2 12 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.115
+ $Y=1.84 $X2=1.25 $Y2=1.985
r41 1 17 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.26 $Y=0.37
+ $X2=1.4 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_2%A_507_392# 1 2 9 11 13 16
c25 9 0 1.40663e-19 $X=3.405 $Y=2.185
r26 11 18 3.10647 $w=3.3e-07 $l=1.6e-07 $layer=LI1_cond $X=3.57 $Y=2.27 $X2=3.57
+ $Y2=2.11
r27 11 13 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=3.57 $Y=2.27
+ $X2=3.57 $Y2=2.815
r28 10 16 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=2.185
+ $X2=2.67 $Y2=2.185
r29 9 18 4.65971 $w=1.7e-07 $l=1.98997e-07 $layer=LI1_cond $X=3.405 $Y=2.185
+ $X2=3.57 $Y2=2.11
r30 9 10 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.405 $Y=2.185
+ $X2=2.755 $Y2=2.185
r31 2 18 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=3.435
+ $Y=1.96 $X2=3.57 $Y2=2.115
r32 2 13 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.435
+ $Y=1.96 $X2=3.57 $Y2=2.815
r33 1 16 300 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_PDIFF $count=2 $X=2.535
+ $Y=1.96 $X2=2.67 $Y2=2.265
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_2%VGND 1 2 3 12 16 18 20 23 24 25 31 35 41 45
r49 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r50 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r51 39 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r52 39 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r53 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r54 36 41 12.2593 $w=1.7e-07 $l=2.88e-07 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.022
+ $Y2=0
r55 36 38 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.31 $Y=0 $X2=3.12
+ $Y2=0
r56 35 44 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.38 $Y=0 $X2=3.61
+ $Y2=0
r57 35 38 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.38 $Y=0 $X2=3.12
+ $Y2=0
r58 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r59 31 41 12.2593 $w=1.7e-07 $l=2.87e-07 $layer=LI1_cond $X=1.735 $Y=0 $X2=2.022
+ $Y2=0
r60 31 33 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.735 $Y=0 $X2=1.68
+ $Y2=0
r61 29 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r62 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r63 25 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r64 25 34 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r65 23 28 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=0 $X2=0.72
+ $Y2=0
r66 23 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.805 $Y=0 $X2=0.93
+ $Y2=0
r67 22 33 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.68
+ $Y2=0
r68 22 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=0.93
+ $Y2=0
r69 18 44 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=3.545 $Y=0.085
+ $X2=3.61 $Y2=0
r70 18 20 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.545 $Y=0.085
+ $X2=3.545 $Y2=0.515
r71 14 41 2.42056 $w=5.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.022 $Y=0.085
+ $X2=2.022 $Y2=0
r72 14 16 10.4007 $w=5.73e-07 $l=5e-07 $layer=LI1_cond $X=2.022 $Y=0.085
+ $X2=2.022 $Y2=0.585
r73 10 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.93 $Y=0.085
+ $X2=0.93 $Y2=0
r74 10 12 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=0.93 $Y=0.085
+ $X2=0.93 $Y2=0.505
r75 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.405
+ $Y=0.37 $X2=3.545 $Y2=0.515
r76 2 16 91 $w=1.7e-07 $l=6.23298e-07 $layer=licon1_NDIFF $count=2 $X=1.69
+ $Y=0.37 $X2=2.215 $Y2=0.585
r77 1 12 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.725
+ $Y=0.56 $X2=0.97 $Y2=0.505
.ends


* NGSPICE file created from sky130_fd_sc_ms__clkinv_8.ext - technology: sky130A

.subckt sky130_fd_sc_ms__clkinv_8 A VGND VNB VPB VPWR Y
M1000 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=1.2264e+12p pd=9.2e+06u as=7.77e+11p ps=7.9e+06u
M1001 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.8144e+12p pd=1.668e+07u as=2.4472e+12p ps=2.005e+07u
M1003 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Y A VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A Y VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y A VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


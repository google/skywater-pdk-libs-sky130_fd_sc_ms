* File: sky130_fd_sc_ms__sedfxtp_4.spice
* Created: Wed Sep  2 12:32:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sedfxtp_4.pex.spice"
.subckt sky130_fd_sc_ms__sedfxtp_4  VNB VPB D DE SCD SCE CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCE	SCE
* SCD	SCD
* DE	DE
* D	D
* VPB	VPB
* VNB	VNB
MM1002 A_135_74# N_D_M1002_g N_A_37_464#_M1002_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_DE_M1026_g A_135_74# VNB NLOWVT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_DE_M1006_g N_A_177_290#_M1006_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1034 A_497_113# N_A_177_290#_M1034_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1018 N_A_37_464#_M1018_d N_A_545_87#_M1018_g A_497_113# VNB NLOWVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1019 N_A_661_113#_M1019_d N_A_631_87#_M1019_g N_A_37_464#_M1018_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.21 AS=0.0588 PD=1.84 PS=0.7 NRD=39.996 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75000.4 A=0.063 P=1.14 MULT=1
MM1043 N_VGND_M1043_d N_SCE_M1043_g N_A_631_87#_M1043_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1007 A_1044_125# N_SCD_M1007_g N_VGND_M1043_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_A_661_113#_M1003_d N_SCE_M1003_g A_1044_125# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1176 AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1020 N_A_1313_74#_M1020_d N_CLK_M1020_g N_VGND_M1020_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2072 AS=0.2109 PD=2.04 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_A_1510_74#_M1011_d N_A_1313_74#_M1011_g N_VGND_M1011_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2072 AS=0.2109 PD=2.04 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1038 N_A_1756_97#_M1038_d N_A_1313_74#_M1038_g N_A_661_113#_M1038_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.083475 AS=0.2226 PD=0.87 PS=1.9 NRD=0 NRS=71.424 M=1 R=2.8
+ SA=75000.5 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1031 A_1858_79# N_A_1510_74#_M1031_g N_A_1756_97#_M1038_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.08925 AS=0.083475 PD=0.845 PS=0.87 NRD=45 NRS=24.276 M=1 R=2.8
+ SA=75000.8 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_A_1943_53#_M1025_g A_1858_79# VNB NLOWVT L=0.15 W=0.42
+ AD=0.109992 AS=0.08925 PD=0.92717 PS=0.845 NRD=0 NRS=45 M=1 R=2.8 SA=75001.4
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1046 N_A_1943_53#_M1046_d N_A_1756_97#_M1046_g N_VGND_M1025_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.167608 PD=1.85 PS=1.41283 NRD=0 NRS=46.872 M=1
+ R=4.26667 SA=75001.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1047 A_2331_74# N_A_1943_53#_M1047_g N_VGND_M1047_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1824 PD=0.85 PS=1.85 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1022 N_A_2403_74#_M1022_d N_A_1510_74#_M1022_g A_2331_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.115623 AS=0.0672 PD=1.16528 PS=0.85 NRD=8.436 NRS=9.372 M=1
+ R=4.26667 SA=75000.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1013 A_2498_74# N_A_1313_74#_M1013_g N_A_2403_74#_M1022_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0758774 PD=0.66 PS=0.764717 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75001 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_A_545_87#_M1014_g A_2498_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.21 AS=0.0504 PD=1.42 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1016 N_A_545_87#_M1016_d N_A_2403_74#_M1016_g N_VGND_M1014_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.21 PD=1.41 PS=1.42 NRD=0 NRS=19.992 M=1 R=2.8 SA=75002.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 N_Q_M1017_d N_A_2403_74#_M1017_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1037 N_Q_M1017_d N_A_2403_74#_M1037_g N_VGND_M1037_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1040 N_Q_M1040_d N_A_2403_74#_M1040_g N_VGND_M1037_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10915 AS=0.1295 PD=1.035 PS=1.09 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1041 N_Q_M1040_d N_A_2403_74#_M1041_g N_VGND_M1041_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10915 AS=0.1998 PD=1.035 PS=2.02 NRD=1.62 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 A_129_464# N_D_M1004_g N_A_37_464#_M1004_s VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.1792 PD=0.88 PS=1.84 NRD=19.9955 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1009 N_VPWR_M1009_d N_A_177_290#_M1009_g A_129_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.1792 AS=0.0768 PD=1.84 PS=0.88 NRD=0 NRS=19.9955 M=1 R=3.55556 SA=90000.6
+ SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1029 N_VPWR_M1029_d N_DE_M1029_g N_A_177_290#_M1029_s VPB PSHORT L=0.18 W=0.64
+ AD=0.16 AS=0.1792 PD=1.14 PS=1.84 NRD=69.2455 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90001.7 A=0.1152 P=1.64 MULT=1
MM1001 A_575_463# N_DE_M1001_g N_VPWR_M1029_d VPB PSHORT L=0.18 W=0.64 AD=0.0672
+ AS=0.16 PD=0.85 PS=1.14 NRD=15.3857 NRS=0 M=1 R=3.55556 SA=90000.9 SB=90001
+ A=0.1152 P=1.64 MULT=1
MM1023 N_A_37_464#_M1023_d N_A_545_87#_M1023_g A_575_463# VPB PSHORT L=0.18
+ W=0.64 AD=0.0864 AS=0.0672 PD=0.91 PS=0.85 NRD=0 NRS=15.3857 M=1 R=3.55556
+ SA=90001.3 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1027 N_A_661_113#_M1027_d N_SCE_M1027_g N_A_37_464#_M1023_d VPB PSHORT L=0.18
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=3.55556 SA=90001.7
+ SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1024 N_VPWR_M1024_d N_SCE_M1024_g N_A_631_87#_M1024_s VPB PSHORT L=0.18 W=0.64
+ AD=0.16 AS=0.1696 PD=1.14 PS=1.81 NRD=69.2455 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90001.2 A=0.1152 P=1.64 MULT=1
MM1005 A_1074_455# N_SCD_M1005_g N_VPWR_M1024_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0672 AS=0.16 PD=0.85 PS=1.14 NRD=15.3857 NRS=0 M=1 R=3.55556 SA=90000.9
+ SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1028 N_A_661_113#_M1028_d N_A_631_87#_M1028_g A_1074_455# VPB PSHORT L=0.18
+ W=0.64 AD=0.1696 AS=0.0672 PD=1.81 PS=0.85 NRD=0 NRS=15.3857 M=1 R=3.55556
+ SA=90001.2 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1010 N_A_1313_74#_M1010_d N_CLK_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.2912 AS=0.2968 PD=2.76 PS=2.77 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1015 N_A_1510_74#_M1015_d N_A_1313_74#_M1015_g N_VPWR_M1015_s VPB PSHORT
+ L=0.18 W=1.12 AD=0.2912 AS=0.2912 PD=2.76 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1033 N_A_1756_97#_M1033_d N_A_1510_74#_M1033_g N_A_661_113#_M1033_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90001.5 A=0.0756 P=1.2 MULT=1
MM1042 A_1902_508# N_A_1313_74#_M1042_g N_A_1756_97#_M1033_d VPB PSHORT L=0.18
+ W=0.42 AD=0.063 AS=0.0567 PD=0.72 PS=0.69 NRD=44.5417 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90001 A=0.0756 P=1.2 MULT=1
MM1036 N_VPWR_M1036_d N_A_1943_53#_M1036_g A_1902_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.0894833 AS=0.063 PD=0.87 PS=0.72 NRD=0 NRS=44.5417 M=1 R=2.33333
+ SA=90001.1 SB=90000.5 A=0.0756 P=1.2 MULT=1
MM1021 N_A_1943_53#_M1021_d N_A_1756_97#_M1021_g N_VPWR_M1036_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2184 AS=0.178967 PD=2.2 PS=1.74 NRD=0 NRS=15.2281 M=1
+ R=4.66667 SA=90000.7 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1044 A_2295_392# N_A_1943_53#_M1044_g N_VPWR_M1044_s VPB PSHORT L=0.18 W=1
+ AD=0.39 AS=0.26 PD=1.78 PS=2.52 NRD=65.9753 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.8 A=0.18 P=2.36 MULT=1
MM1035 N_A_2403_74#_M1035_d N_A_1313_74#_M1035_g A_2295_392# VPB PSHORT L=0.18
+ W=1 AD=0.199718 AS=0.39 PD=1.87324 PS=1.78 NRD=10.8153 NRS=65.9753 M=1
+ R=5.55556 SA=90001.1 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1000 A_2589_508# N_A_1510_74#_M1000_g N_A_2403_74#_M1035_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0838817 PD=0.66 PS=0.786761 NRD=30.4759 NRS=0 M=1
+ R=2.33333 SA=90001.6 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1008 N_VPWR_M1008_d N_A_545_87#_M1008_g A_2589_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.109992 AS=0.0504 PD=0.92717 PS=0.66 NRD=46.886 NRS=30.4759 M=1 R=2.33333
+ SA=90002.1 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1030 N_A_545_87#_M1030_d N_A_2403_74#_M1030_g N_VPWR_M1008_d VPB PSHORT L=0.18
+ W=0.64 AD=0.1664 AS=0.167608 PD=1.8 PS=1.41283 NRD=0 NRS=46.1571 M=1 R=3.55556
+ SA=90001.9 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1012 N_Q_M1012_d N_A_2403_74#_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1032 N_Q_M1012_d N_A_2403_74#_M1032_g N_VPWR_M1032_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1039 N_Q_M1039_d N_A_2403_74#_M1039_g N_VPWR_M1032_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1045 N_Q_M1039_d N_A_2403_74#_M1045_g N_VPWR_M1045_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3024 PD=1.39 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX48_noxref VNB VPB NWDIODE A=31.9921 P=38.15
c_177 VNB 0 1.36415e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__sedfxtp_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__a211oi_4.pex.spice
* Created: Fri Aug 28 16:57:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A211OI_4%A2 3 7 11 15 19 23 27 31 33 34 35 36 37 57
c81 31 0 2.04552e-19 $X=2.09 $Y=0.74
r82 56 57 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=2.085 $Y=1.515
+ $X2=2.09 $Y2=1.515
r83 54 56 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=1.83 $Y=1.515
+ $X2=2.085 $Y2=1.515
r84 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.83
+ $Y=1.515 $X2=1.83 $Y2=1.515
r85 52 54 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=1.66 $Y=1.515
+ $X2=1.83 $Y2=1.515
r86 51 52 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.635 $Y=1.515
+ $X2=1.66 $Y2=1.515
r87 50 51 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=1.23 $Y=1.515
+ $X2=1.635 $Y2=1.515
r88 49 50 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=1.185 $Y=1.515
+ $X2=1.23 $Y2=1.515
r89 47 49 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=0.81 $Y=1.515
+ $X2=1.185 $Y2=1.515
r90 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.81
+ $Y=1.515 $X2=0.81 $Y2=1.515
r91 45 47 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.8 $Y=1.515 $X2=0.81
+ $Y2=1.515
r92 43 45 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=0.735 $Y=1.515
+ $X2=0.8 $Y2=1.515
r93 37 55 8.84433 $w=4.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=1.83 $Y2=1.565
r94 36 55 4.02015 $w=4.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.83 $Y2=1.565
r95 35 36 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.68 $Y2=1.565
r96 35 48 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=0.81 $Y2=1.565
r97 34 48 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=0.72 $Y=1.565 $X2=0.81
+ $Y2=1.565
r98 33 34 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.72 $Y2=1.565
r99 29 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.09 $Y=1.35
+ $X2=2.09 $Y2=1.515
r100 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.09 $Y=1.35
+ $X2=2.09 $Y2=0.74
r101 25 56 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.085 $Y=1.68
+ $X2=2.085 $Y2=1.515
r102 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.085 $Y=1.68
+ $X2=2.085 $Y2=2.4
r103 21 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.66 $Y=1.35
+ $X2=1.66 $Y2=1.515
r104 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.66 $Y=1.35
+ $X2=1.66 $Y2=0.74
r105 17 51 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.635 $Y=1.68
+ $X2=1.635 $Y2=1.515
r106 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.635 $Y=1.68
+ $X2=1.635 $Y2=2.4
r107 13 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.23 $Y=1.35
+ $X2=1.23 $Y2=1.515
r108 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.23 $Y=1.35
+ $X2=1.23 $Y2=0.74
r109 9 49 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.185 $Y=1.68
+ $X2=1.185 $Y2=1.515
r110 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.185 $Y=1.68
+ $X2=1.185 $Y2=2.4
r111 5 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.8 $Y=1.35 $X2=0.8
+ $Y2=1.515
r112 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.8 $Y=1.35 $X2=0.8
+ $Y2=0.74
r113 1 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.735 $Y=1.68
+ $X2=0.735 $Y2=1.515
r114 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.735 $Y=1.68
+ $X2=0.735 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A211OI_4%A1 3 7 11 15 19 23 27 31 33 34 35 51 53
r73 52 53 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.81 $Y=1.515
+ $X2=3.885 $Y2=1.515
r74 50 52 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=3.69 $Y=1.515
+ $X2=3.81 $Y2=1.515
r75 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.69
+ $Y=1.515 $X2=3.69 $Y2=1.515
r76 48 50 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=3.435 $Y=1.515
+ $X2=3.69 $Y2=1.515
r77 47 48 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=3.38 $Y=1.515
+ $X2=3.435 $Y2=1.515
r78 46 47 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=2.985 $Y=1.515
+ $X2=3.38 $Y2=1.515
r79 45 46 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=2.95 $Y=1.515
+ $X2=2.985 $Y2=1.515
r80 43 45 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=2.67 $Y=1.515
+ $X2=2.95 $Y2=1.515
r81 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.67
+ $Y=1.515 $X2=2.67 $Y2=1.515
r82 41 43 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.535 $Y=1.515
+ $X2=2.67 $Y2=1.515
r83 39 41 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.52 $Y=1.515
+ $X2=2.535 $Y2=1.515
r84 35 51 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=3.6 $Y=1.565 $X2=3.69
+ $Y2=1.565
r85 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.6 $Y2=1.565
r86 34 44 12.0604 $w=4.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=2.67 $Y2=1.565
r87 33 44 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=2.64 $Y=1.565 $X2=2.67
+ $Y2=1.565
r88 29 53 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.885 $Y=1.68
+ $X2=3.885 $Y2=1.515
r89 29 31 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.885 $Y=1.68
+ $X2=3.885 $Y2=2.4
r90 25 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.81 $Y=1.35
+ $X2=3.81 $Y2=1.515
r91 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.81 $Y=1.35
+ $X2=3.81 $Y2=0.74
r92 21 48 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.435 $Y=1.68
+ $X2=3.435 $Y2=1.515
r93 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.435 $Y=1.68
+ $X2=3.435 $Y2=2.4
r94 17 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.38 $Y=1.35
+ $X2=3.38 $Y2=1.515
r95 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.38 $Y=1.35
+ $X2=3.38 $Y2=0.74
r96 13 46 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.985 $Y=1.68
+ $X2=2.985 $Y2=1.515
r97 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.985 $Y=1.68
+ $X2=2.985 $Y2=2.4
r98 9 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.35
+ $X2=2.95 $Y2=1.515
r99 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.95 $Y=1.35 $X2=2.95
+ $Y2=0.74
r100 5 41 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.535 $Y=1.68
+ $X2=2.535 $Y2=1.515
r101 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.535 $Y=1.68
+ $X2=2.535 $Y2=2.4
r102 1 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.52 $Y=1.35
+ $X2=2.52 $Y2=1.515
r103 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.52 $Y=1.35 $X2=2.52
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A211OI_4%B1 3 7 11 15 19 23 25 26 27 28 43
c76 28 0 7.2903e-20 $X=6 $Y=1.665
r77 43 44 2.19757 $w=3.29e-07 $l=1.5e-08 $layer=POLY_cond $X=6.19 $Y=1.465
+ $X2=6.205 $Y2=1.465
r78 41 43 35.1611 $w=3.29e-07 $l=2.4e-07 $layer=POLY_cond $X=5.95 $Y=1.465
+ $X2=6.19 $Y2=1.465
r79 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.95
+ $Y=1.465 $X2=5.95 $Y2=1.465
r80 39 41 27.8359 $w=3.29e-07 $l=1.9e-07 $layer=POLY_cond $X=5.76 $Y=1.465
+ $X2=5.95 $Y2=1.465
r81 38 39 0.732523 $w=3.29e-07 $l=5e-09 $layer=POLY_cond $X=5.755 $Y=1.465
+ $X2=5.76 $Y2=1.465
r82 37 38 65.9271 $w=3.29e-07 $l=4.5e-07 $layer=POLY_cond $X=5.305 $Y=1.465
+ $X2=5.755 $Y2=1.465
r83 35 37 54.9392 $w=3.29e-07 $l=3.75e-07 $layer=POLY_cond $X=4.93 $Y=1.465
+ $X2=5.305 $Y2=1.465
r84 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.93
+ $Y=1.465 $X2=4.93 $Y2=1.465
r85 33 35 10.9878 $w=3.29e-07 $l=7.5e-08 $layer=POLY_cond $X=4.855 $Y=1.465
+ $X2=4.93 $Y2=1.465
r86 28 42 1.24592 $w=4.78e-07 $l=5e-08 $layer=LI1_cond $X=6 $Y=1.54 $X2=5.95
+ $Y2=1.54
r87 27 42 10.7149 $w=4.78e-07 $l=4.3e-07 $layer=LI1_cond $X=5.52 $Y=1.54
+ $X2=5.95 $Y2=1.54
r88 26 27 11.9608 $w=4.78e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.54
+ $X2=5.52 $Y2=1.54
r89 26 36 2.74101 $w=4.78e-07 $l=1.1e-07 $layer=LI1_cond $X=5.04 $Y=1.54
+ $X2=4.93 $Y2=1.54
r90 25 36 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=4.56 $Y=1.54
+ $X2=4.93 $Y2=1.54
r91 21 44 16.8611 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.205 $Y=1.63
+ $X2=6.205 $Y2=1.465
r92 21 23 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=6.205 $Y=1.63
+ $X2=6.205 $Y2=2.4
r93 17 43 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.19 $Y=1.3
+ $X2=6.19 $Y2=1.465
r94 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.19 $Y=1.3 $X2=6.19
+ $Y2=0.74
r95 13 39 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.76 $Y=1.3
+ $X2=5.76 $Y2=1.465
r96 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.76 $Y=1.3 $X2=5.76
+ $Y2=0.74
r97 9 38 16.8611 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.755 $Y=1.63
+ $X2=5.755 $Y2=1.465
r98 9 11 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=5.755 $Y=1.63
+ $X2=5.755 $Y2=2.4
r99 5 37 16.8611 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.305 $Y=1.63
+ $X2=5.305 $Y2=1.465
r100 5 7 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=5.305 $Y=1.63
+ $X2=5.305 $Y2=2.4
r101 1 33 16.8611 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.855 $Y=1.63
+ $X2=4.855 $Y2=1.465
r102 1 3 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.855 $Y=1.63
+ $X2=4.855 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A211OI_4%C1 3 7 11 15 19 23 25 26 27 43
c62 7 0 7.2903e-20 $X=6.655 $Y=2.4
r63 42 43 72.1303 $w=3.6e-07 $l=4.5e-07 $layer=POLY_cond $X=7.555 $Y=1.5
+ $X2=8.005 $Y2=1.5
r64 40 42 26.4478 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=7.39 $Y=1.5
+ $X2=7.555 $Y2=1.5
r65 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.39
+ $Y=1.515 $X2=7.39 $Y2=1.515
r66 38 40 45.6825 $w=3.6e-07 $l=2.85e-07 $layer=POLY_cond $X=7.105 $Y=1.5
+ $X2=7.39 $Y2=1.5
r67 37 38 8.81592 $w=3.6e-07 $l=5.5e-08 $layer=POLY_cond $X=7.05 $Y=1.5
+ $X2=7.105 $Y2=1.5
r68 35 37 54.4984 $w=3.6e-07 $l=3.4e-07 $layer=POLY_cond $X=6.71 $Y=1.5 $X2=7.05
+ $Y2=1.5
r69 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.71
+ $Y=1.515 $X2=6.71 $Y2=1.515
r70 33 35 8.81592 $w=3.6e-07 $l=5.5e-08 $layer=POLY_cond $X=6.655 $Y=1.5
+ $X2=6.71 $Y2=1.5
r71 31 33 5.61013 $w=3.6e-07 $l=3.5e-08 $layer=POLY_cond $X=6.62 $Y=1.5
+ $X2=6.655 $Y2=1.5
r72 27 41 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=7.44 $Y=1.565 $X2=7.39
+ $Y2=1.565
r73 26 41 11.5244 $w=4.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.39 $Y2=1.565
r74 26 36 6.70025 $w=4.28e-07 $l=2.5e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=6.71 $Y2=1.565
r75 25 36 6.16423 $w=4.28e-07 $l=2.3e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.71 $Y2=1.565
r76 21 43 18.9685 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=8.005 $Y=1.68
+ $X2=8.005 $Y2=1.5
r77 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.005 $Y=1.68
+ $X2=8.005 $Y2=2.4
r78 17 42 18.9685 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=7.555 $Y=1.68
+ $X2=7.555 $Y2=1.5
r79 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.555 $Y=1.68
+ $X2=7.555 $Y2=2.4
r80 13 38 18.9685 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=7.105 $Y=1.68
+ $X2=7.105 $Y2=1.5
r81 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.105 $Y=1.68
+ $X2=7.105 $Y2=2.4
r82 9 37 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.05 $Y=1.32 $X2=7.05
+ $Y2=1.5
r83 9 11 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.05 $Y=1.32 $X2=7.05
+ $Y2=0.74
r84 5 33 18.9685 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=6.655 $Y=1.68
+ $X2=6.655 $Y2=1.5
r85 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.655 $Y=1.68
+ $X2=6.655 $Y2=2.4
r86 1 31 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.62 $Y=1.32 $X2=6.62
+ $Y2=1.5
r87 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.62 $Y=1.32 $X2=6.62
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A211OI_4%A_77_368# 1 2 3 4 5 6 7 22 24 26 30 32 36
+ 38 42 44 48 50 54 56 58 60 65 67 69 71 73
r93 58 75 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.02 $Y=2.12 $X2=6.02
+ $Y2=2.035
r94 58 60 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=6.02 $Y=2.12 $X2=6.02
+ $Y2=2.57
r95 57 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.165 $Y=2.035
+ $X2=5.08 $Y2=2.035
r96 56 75 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.895 $Y=2.035
+ $X2=6.02 $Y2=2.035
r97 56 57 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.895 $Y=2.035
+ $X2=5.165 $Y2=2.035
r98 52 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.08 $Y=2.12 $X2=5.08
+ $Y2=2.035
r99 52 54 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=5.08 $Y=2.12
+ $X2=5.08 $Y2=2.57
r100 51 71 7.02821 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=4.275 $Y=2.035
+ $X2=4.15 $Y2=1.97
r101 50 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.995 $Y=2.035
+ $X2=5.08 $Y2=2.035
r102 50 51 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=4.995 $Y=2.035
+ $X2=4.275 $Y2=2.035
r103 46 71 0.00168595 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=4.15 $Y=2.12
+ $X2=4.15 $Y2=1.97
r104 46 48 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=4.15 $Y=2.12
+ $X2=4.15 $Y2=2.4
r105 45 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.295 $Y=2.035
+ $X2=3.21 $Y2=2.035
r106 44 71 7.02821 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=4.025 $Y=2.035
+ $X2=4.15 $Y2=1.97
r107 44 45 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.025 $Y=2.035
+ $X2=3.295 $Y2=2.035
r108 40 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.21 $Y=2.12
+ $X2=3.21 $Y2=2.035
r109 40 42 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.21 $Y=2.12
+ $X2=3.21 $Y2=2.445
r110 39 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.395 $Y=2.035
+ $X2=2.31 $Y2=2.035
r111 38 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.125 $Y=2.035
+ $X2=3.21 $Y2=2.035
r112 38 39 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.125 $Y=2.035
+ $X2=2.395 $Y2=2.035
r113 34 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.31 $Y=2.12
+ $X2=2.31 $Y2=2.035
r114 34 36 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.31 $Y=2.12
+ $X2=2.31 $Y2=2.445
r115 33 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.495 $Y=2.035
+ $X2=1.37 $Y2=2.035
r116 32 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=2.035
+ $X2=2.31 $Y2=2.035
r117 32 33 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.225 $Y=2.035
+ $X2=1.495 $Y2=2.035
r118 28 65 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.37 $Y=2.12
+ $X2=1.37 $Y2=2.035
r119 28 30 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=1.37 $Y=2.12
+ $X2=1.37 $Y2=2.445
r120 27 63 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.675 $Y=2.035
+ $X2=0.51 $Y2=2.035
r121 26 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.245 $Y=2.035
+ $X2=1.37 $Y2=2.035
r122 26 27 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.245 $Y=2.035
+ $X2=0.675 $Y2=2.035
r123 22 63 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.51 $Y=2.12 $X2=0.51
+ $Y2=2.035
r124 22 24 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.51 $Y=2.12
+ $X2=0.51 $Y2=2.815
r125 7 75 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=5.845
+ $Y=1.84 $X2=5.98 $Y2=2.035
r126 7 60 600 $w=1.7e-07 $l=7.94638e-07 $layer=licon1_PDIFF $count=1 $X=5.845
+ $Y=1.84 $X2=5.98 $Y2=2.57
r127 6 73 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=4.945
+ $Y=1.84 $X2=5.08 $Y2=2.035
r128 6 54 600 $w=1.7e-07 $l=7.94638e-07 $layer=licon1_PDIFF $count=1 $X=4.945
+ $Y=1.84 $X2=5.08 $Y2=2.57
r129 5 71 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.975
+ $Y=1.84 $X2=4.11 $Y2=1.985
r130 5 48 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=3.975
+ $Y=1.84 $X2=4.11 $Y2=2.4
r131 4 69 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=3.075
+ $Y=1.84 $X2=3.21 $Y2=2.035
r132 4 42 300 $w=1.7e-07 $l=6.69104e-07 $layer=licon1_PDIFF $count=2 $X=3.075
+ $Y=1.84 $X2=3.21 $Y2=2.445
r133 3 67 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=2.175
+ $Y=1.84 $X2=2.31 $Y2=2.035
r134 3 36 300 $w=1.7e-07 $l=6.69104e-07 $layer=licon1_PDIFF $count=2 $X=2.175
+ $Y=1.84 $X2=2.31 $Y2=2.445
r135 2 65 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=1.275
+ $Y=1.84 $X2=1.41 $Y2=2.035
r136 2 30 300 $w=1.7e-07 $l=6.69104e-07 $layer=licon1_PDIFF $count=2 $X=1.275
+ $Y=1.84 $X2=1.41 $Y2=2.445
r137 1 63 400 $w=1.7e-07 $l=2.498e-07 $layer=licon1_PDIFF $count=1 $X=0.385
+ $Y=1.84 $X2=0.51 $Y2=2.035
r138 1 24 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.385
+ $Y=1.84 $X2=0.51 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__A211OI_4%VPWR 1 2 3 4 15 19 21 25 29 32 33 34 35 36
+ 45 55 56 59 62
r103 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r104 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r105 55 56 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r106 53 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r107 52 55 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=8.4 $Y2=3.33
r108 52 53 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r109 50 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.825 $Y=3.33
+ $X2=3.66 $Y2=3.33
r110 50 52 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.825 $Y=3.33
+ $X2=4.08 $Y2=3.33
r111 49 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r112 49 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r113 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r114 46 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.925 $Y=3.33
+ $X2=2.76 $Y2=3.33
r115 46 48 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.925 $Y=3.33
+ $X2=3.12 $Y2=3.33
r116 45 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.495 $Y=3.33
+ $X2=3.66 $Y2=3.33
r117 45 48 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.495 $Y=3.33
+ $X2=3.12 $Y2=3.33
r118 44 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r119 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r120 40 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r121 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r122 36 56 1.13724 $w=4.9e-07 $l=4.08e-06 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=8.4 $Y2=3.33
r123 36 53 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r124 34 43 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.695 $Y=3.33
+ $X2=1.68 $Y2=3.33
r125 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.695 $Y=3.33
+ $X2=1.86 $Y2=3.33
r126 32 39 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.875 $Y=3.33
+ $X2=0.72 $Y2=3.33
r127 32 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.875 $Y=3.33
+ $X2=0.96 $Y2=3.33
r128 31 43 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.045 $Y=3.33
+ $X2=1.68 $Y2=3.33
r129 31 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.045 $Y=3.33
+ $X2=0.96 $Y2=3.33
r130 27 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.66 $Y=3.245
+ $X2=3.66 $Y2=3.33
r131 27 29 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=3.66 $Y=3.245
+ $X2=3.66 $Y2=2.41
r132 23 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.76 $Y=3.245
+ $X2=2.76 $Y2=3.33
r133 23 25 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=2.76 $Y=3.245
+ $X2=2.76 $Y2=2.41
r134 22 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=1.86 $Y2=3.33
r135 21 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.595 $Y=3.33
+ $X2=2.76 $Y2=3.33
r136 21 22 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.595 $Y=3.33
+ $X2=2.025 $Y2=3.33
r137 17 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.86 $Y=3.245
+ $X2=1.86 $Y2=3.33
r138 17 19 29.1603 $w=3.28e-07 $l=8.35e-07 $layer=LI1_cond $X=1.86 $Y=3.245
+ $X2=1.86 $Y2=2.41
r139 13 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.96 $Y=3.245
+ $X2=0.96 $Y2=3.33
r140 13 15 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.96 $Y=3.245
+ $X2=0.96 $Y2=2.455
r141 4 29 300 $w=1.7e-07 $l=6.33916e-07 $layer=licon1_PDIFF $count=2 $X=3.525
+ $Y=1.84 $X2=3.66 $Y2=2.41
r142 3 25 300 $w=1.7e-07 $l=6.33916e-07 $layer=licon1_PDIFF $count=2 $X=2.625
+ $Y=1.84 $X2=2.76 $Y2=2.41
r143 2 19 300 $w=1.7e-07 $l=6.33916e-07 $layer=licon1_PDIFF $count=2 $X=1.725
+ $Y=1.84 $X2=1.86 $Y2=2.41
r144 1 15 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=0.825
+ $Y=1.84 $X2=0.96 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__A211OI_4%A_901_368# 1 2 3 4 5 18 20 21 24 26 30 34
+ 38 40 44 46 47 48
r75 42 44 21.652 $w=3.28e-07 $l=6.2e-07 $layer=LI1_cond $X=8.23 $Y=2.905
+ $X2=8.23 $Y2=2.285
r76 41 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.495 $Y=2.99
+ $X2=7.33 $Y2=2.99
r77 40 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.065 $Y=2.99
+ $X2=8.23 $Y2=2.905
r78 40 41 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.065 $Y=2.99
+ $X2=7.495 $Y2=2.99
r79 36 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.33 $Y=2.905
+ $X2=7.33 $Y2=2.99
r80 36 38 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=7.33 $Y=2.905
+ $X2=7.33 $Y2=2.455
r81 35 47 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=6.595 $Y=2.99
+ $X2=6.455 $Y2=2.99
r82 34 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.165 $Y=2.99
+ $X2=7.33 $Y2=2.99
r83 34 35 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=7.165 $Y=2.99
+ $X2=6.595 $Y2=2.99
r84 30 33 28.8111 $w=2.78e-07 $l=7e-07 $layer=LI1_cond $X=6.455 $Y=2.115
+ $X2=6.455 $Y2=2.815
r85 28 47 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.455 $Y=2.905
+ $X2=6.455 $Y2=2.99
r86 28 33 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=6.455 $Y=2.905
+ $X2=6.455 $Y2=2.815
r87 27 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.695 $Y=2.99
+ $X2=5.53 $Y2=2.99
r88 26 47 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=6.315 $Y=2.99
+ $X2=6.455 $Y2=2.99
r89 26 27 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=6.315 $Y=2.99
+ $X2=5.695 $Y2=2.99
r90 22 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.53 $Y=2.905
+ $X2=5.53 $Y2=2.99
r91 22 24 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=5.53 $Y=2.905
+ $X2=5.53 $Y2=2.395
r92 20 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.365 $Y=2.99
+ $X2=5.53 $Y2=2.99
r93 20 21 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.365 $Y=2.99
+ $X2=4.795 $Y2=2.99
r94 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.63 $Y=2.905
+ $X2=4.795 $Y2=2.99
r95 16 18 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=4.63 $Y=2.905
+ $X2=4.63 $Y2=2.395
r96 5 44 300 $w=1.7e-07 $l=5.08035e-07 $layer=licon1_PDIFF $count=2 $X=8.095
+ $Y=1.84 $X2=8.23 $Y2=2.285
r97 4 38 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=7.195
+ $Y=1.84 $X2=7.33 $Y2=2.455
r98 3 33 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=1.84 $X2=6.43 $Y2=2.815
r99 3 30 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=1.84 $X2=6.43 $Y2=2.115
r100 2 24 300 $w=1.7e-07 $l=6.1883e-07 $layer=licon1_PDIFF $count=2 $X=5.395
+ $Y=1.84 $X2=5.53 $Y2=2.395
r101 1 18 300 $w=1.7e-07 $l=6.14329e-07 $layer=licon1_PDIFF $count=2 $X=4.505
+ $Y=1.84 $X2=4.63 $Y2=2.395
.ends

.subckt PM_SKY130_FD_SC_MS__A211OI_4%Y 1 2 3 4 5 6 7 22 26 30 32 36 38 42 48 49
+ 50 52 53 54 55 56 57 58 59 60
c73 22 0 4.29123e-20 $X=3.588 $Y=0.957
r74 56 60 11.6415 $w=1.7e-07 $l=5.53e-07 $layer=LI1_cond $X=7.847 $Y=1.665
+ $X2=8.4 $Y2=1.665
r75 55 56 4.56883 $w=9.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.847 $Y=1.295
+ $X2=7.847 $Y2=1.665
r76 55 59 11.6415 $w=1.7e-07 $l=5.53e-07 $layer=LI1_cond $X=7.847 $Y=1.295
+ $X2=8.4 $Y2=1.295
r77 55 77 2.46964 $w=9.88e-07 $l=2e-07 $layer=LI1_cond $X=7.847 $Y=1.295
+ $X2=7.847 $Y2=1.095
r78 54 77 2.09919 $w=9.88e-07 $l=1.7e-07 $layer=LI1_cond $X=7.847 $Y=0.925
+ $X2=7.847 $Y2=1.095
r79 54 58 11.6415 $w=1.7e-07 $l=5.53e-07 $layer=LI1_cond $X=7.847 $Y=0.925
+ $X2=8.4 $Y2=0.925
r80 53 54 4.56883 $w=9.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.847 $Y=0.555
+ $X2=7.847 $Y2=0.925
r81 53 57 11.6415 $w=1.7e-07 $l=5.53e-07 $layer=LI1_cond $X=7.847 $Y=0.555
+ $X2=8.4 $Y2=0.555
r82 53 70 0.493927 $w=9.88e-07 $l=4e-08 $layer=LI1_cond $X=7.847 $Y=0.555
+ $X2=7.847 $Y2=0.515
r83 47 48 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=0.957
+ $X2=3.76 $Y2=0.957
r84 43 52 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.965 $Y=2.035
+ $X2=6.88 $Y2=2.035
r85 42 56 4.56883 $w=9.88e-07 $l=3.7e-07 $layer=LI1_cond $X=7.847 $Y=2.035
+ $X2=7.847 $Y2=1.665
r86 42 43 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=7.695 $Y=2.035
+ $X2=6.965 $Y2=2.035
r87 39 50 5.16603 $w=1.7e-07 $l=9.66954e-08 $layer=LI1_cond $X=6.49 $Y=1.095
+ $X2=6.405 $Y2=1.07
r88 38 77 11.6415 $w=1.7e-07 $l=6.67e-07 $layer=LI1_cond $X=7.18 $Y=1.095
+ $X2=7.847 $Y2=1.095
r89 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.18 $Y=1.095
+ $X2=6.49 $Y2=1.095
r90 34 50 1.34256 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=6.405 $Y=0.96
+ $X2=6.405 $Y2=1.07
r91 34 36 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=6.405 $Y=0.96
+ $X2=6.405 $Y2=0.515
r92 33 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.63 $Y=1.045
+ $X2=5.505 $Y2=1.045
r93 32 50 5.16603 $w=1.7e-07 $l=9.66954e-08 $layer=LI1_cond $X=6.32 $Y=1.045
+ $X2=6.405 $Y2=1.07
r94 32 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.32 $Y=1.045
+ $X2=5.63 $Y2=1.045
r95 28 49 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.505 $Y=0.96
+ $X2=5.505 $Y2=1.045
r96 28 30 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=5.505 $Y=0.96
+ $X2=5.505 $Y2=0.515
r97 26 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.38 $Y=1.045
+ $X2=5.505 $Y2=1.045
r98 26 48 105.69 $w=1.68e-07 $l=1.62e-06 $layer=LI1_cond $X=5.38 $Y=1.045
+ $X2=3.76 $Y2=1.045
r99 22 47 0.233829 $w=3.43e-07 $l=7e-09 $layer=LI1_cond $X=3.588 $Y=0.957
+ $X2=3.595 $Y2=0.957
r100 22 24 28.4937 $w=3.43e-07 $l=8.53e-07 $layer=LI1_cond $X=3.588 $Y=0.957
+ $X2=2.735 $Y2=0.957
r101 7 42 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=7.645
+ $Y=1.84 $X2=7.78 $Y2=2.115
r102 6 52 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=6.745
+ $Y=1.84 $X2=6.88 $Y2=2.115
r103 5 70 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.125
+ $Y=0.37 $X2=7.265 $Y2=0.515
r104 4 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.265
+ $Y=0.37 $X2=6.405 $Y2=0.515
r105 3 30 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=5.42
+ $Y=0.37 $X2=5.545 $Y2=0.515
r106 2 47 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=3.455
+ $Y=0.37 $X2=3.595 $Y2=0.95
r107 1 24 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=2.595
+ $Y=0.37 $X2=2.735 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_MS__A211OI_4%A_92_74# 1 2 3 4 5 18 20 21 24 26 28 36 38
c51 28 0 1.6164e-19 $X=2.305 $Y=0.615
r52 34 36 37.4 $w=2.63e-07 $l=8.6e-07 $layer=LI1_cond $X=3.165 $Y=0.482
+ $X2=4.025 $Y2=0.482
r53 32 40 2.82608 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.39 $Y=0.482
+ $X2=2.305 $Y2=0.482
r54 32 34 33.7035 $w=2.63e-07 $l=7.75e-07 $layer=LI1_cond $X=2.39 $Y=0.482
+ $X2=3.165 $Y2=0.482
r55 29 31 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.305 $Y=1.01
+ $X2=2.305 $Y2=0.965
r56 28 40 4.42198 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=2.305 $Y=0.615
+ $X2=2.305 $Y2=0.482
r57 28 31 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.305 $Y=0.615
+ $X2=2.305 $Y2=0.965
r58 27 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.53 $Y=1.095
+ $X2=1.445 $Y2=1.095
r59 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.22 $Y=1.095
+ $X2=2.305 $Y2=1.01
r60 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.22 $Y=1.095
+ $X2=1.53 $Y2=1.095
r61 22 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.445 $Y=1.01
+ $X2=1.445 $Y2=1.095
r62 22 24 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.445 $Y=1.01
+ $X2=1.445 $Y2=0.515
r63 20 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.36 $Y=1.095
+ $X2=1.445 $Y2=1.095
r64 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.36 $Y=1.095
+ $X2=0.67 $Y2=1.095
r65 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.545 $Y=1.01
+ $X2=0.67 $Y2=1.095
r66 16 18 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.545 $Y=1.01
+ $X2=0.545 $Y2=0.515
r67 5 36 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.37 $X2=4.025 $Y2=0.515
r68 4 34 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.025
+ $Y=0.37 $X2=3.165 $Y2=0.515
r69 3 40 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.165
+ $Y=0.37 $X2=2.305 $Y2=0.515
r70 3 31 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=2.165
+ $Y=0.37 $X2=2.305 $Y2=0.965
r71 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.305
+ $Y=0.37 $X2=1.445 $Y2=0.515
r72 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.46
+ $Y=0.37 $X2=0.585 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A211OI_4%VGND 1 2 3 4 15 19 23 27 30 31 33 34 35 44
+ 51 58 59 62 65
r81 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r82 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r83 59 66 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.4 $Y=0 $X2=6.96
+ $Y2=0
r84 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r85 56 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7 $Y=0 $X2=6.835
+ $Y2=0
r86 56 58 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=7 $Y=0 $X2=8.4 $Y2=0
r87 55 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r88 55 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r89 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r90 52 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.14 $Y=0 $X2=5.975
+ $Y2=0
r91 52 54 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.14 $Y=0 $X2=6.48
+ $Y2=0
r92 51 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.67 $Y=0 $X2=6.835
+ $Y2=0
r93 51 54 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=6.67 $Y=0 $X2=6.48
+ $Y2=0
r94 50 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r95 49 50 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r96 46 49 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=5.52
+ $Y2=0
r97 46 47 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r98 44 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.81 $Y=0 $X2=5.975
+ $Y2=0
r99 44 49 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.81 $Y=0 $X2=5.52
+ $Y2=0
r100 43 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r101 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r102 39 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r103 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r104 35 50 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.32 $Y=0 $X2=5.52
+ $Y2=0
r105 35 47 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=2.16 $Y2=0
r106 33 42 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.71 $Y=0 $X2=1.68
+ $Y2=0
r107 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.71 $Y=0 $X2=1.875
+ $Y2=0
r108 32 46 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.04 $Y=0 $X2=2.16
+ $Y2=0
r109 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.04 $Y=0 $X2=1.875
+ $Y2=0
r110 30 38 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.85 $Y=0 $X2=0.72
+ $Y2=0
r111 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.85 $Y=0 $X2=1.015
+ $Y2=0
r112 29 42 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=1.18 $Y=0 $X2=1.68
+ $Y2=0
r113 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.18 $Y=0 $X2=1.015
+ $Y2=0
r114 25 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.835 $Y=0.085
+ $X2=6.835 $Y2=0
r115 25 27 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=6.835 $Y=0.085
+ $X2=6.835 $Y2=0.675
r116 21 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.975 $Y=0.085
+ $X2=5.975 $Y2=0
r117 21 23 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=5.975 $Y=0.085
+ $X2=5.975 $Y2=0.625
r118 17 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=0.085
+ $X2=1.875 $Y2=0
r119 17 19 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.875 $Y=0.085
+ $X2=1.875 $Y2=0.675
r120 13 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=0.085
+ $X2=1.015 $Y2=0
r121 13 15 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.015 $Y=0.085
+ $X2=1.015 $Y2=0.675
r122 4 27 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=6.695
+ $Y=0.37 $X2=6.835 $Y2=0.675
r123 3 23 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=5.835
+ $Y=0.37 $X2=5.975 $Y2=0.625
r124 2 19 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.735
+ $Y=0.37 $X2=1.875 $Y2=0.675
r125 1 15 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=0.875
+ $Y=0.37 $X2=1.015 $Y2=0.675
.ends


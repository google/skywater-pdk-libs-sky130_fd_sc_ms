* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and3_4 A B C VGND VNB VPB VPWR X
M1000 a_686_74# B a_489_74# VNB nlowvt w=640000u l=150000u
+  ad=5.76e+11p pd=5.64e+06u as=3.84e+11p ps=3.76e+06u
M1001 VPWR B a_83_260# VPB pshort w=840000u l=180000u
+  ad=2.184e+12p pd=1.636e+07u as=7.14e+11p ps=6.74e+06u
M1002 a_489_74# B a_686_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_83_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1004 VPWR a_83_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_83_260# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_83_260# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_83_260# C VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR C a_83_260# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_489_74# C VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=9.013e+11p ps=8.26e+06u
M1010 a_83_260# A a_686_74# VNB nlowvt w=640000u l=150000u
+  ad=2.368e+11p pd=2.02e+06u as=0p ps=0u
M1011 VGND a_83_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.144e+11p ps=4.08e+06u
M1012 a_83_260# A VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_83_260# B VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND C a_489_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_83_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR A a_83_260# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_83_260# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_83_260# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_686_74# A a_83_260# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_ms__o41ai_4.pxi.spice
* Created: Wed Sep  2 12:27:23 2020
* 
x_PM_SKY130_FD_SC_MS__O41AI_4%B1 N_B1_M1004_g N_B1_c_156_n N_B1_M1009_g
+ N_B1_c_157_n N_B1_M1010_g N_B1_M1008_g N_B1_c_159_n N_B1_M1029_g N_B1_c_160_n
+ N_B1_c_161_n N_B1_c_162_n N_B1_M1030_g B1 B1 N_B1_c_163_n
+ PM_SKY130_FD_SC_MS__O41AI_4%B1
x_PM_SKY130_FD_SC_MS__O41AI_4%A4 N_A4_c_230_n N_A4_M1015_g N_A4_c_223_n
+ N_A4_M1000_g N_A4_c_231_n N_A4_M1018_g N_A4_c_232_n N_A4_M1020_g N_A4_c_224_n
+ N_A4_M1007_g N_A4_c_233_n N_A4_M1023_g N_A4_c_225_n N_A4_M1012_g N_A4_c_226_n
+ N_A4_c_227_n N_A4_c_228_n N_A4_M1017_g A4 A4 N_A4_c_229_n
+ PM_SKY130_FD_SC_MS__O41AI_4%A4
x_PM_SKY130_FD_SC_MS__O41AI_4%A3 N_A3_c_335_n N_A3_M1003_g N_A3_c_327_n
+ N_A3_c_328_n N_A3_c_329_n N_A3_M1001_g N_A3_c_338_n N_A3_M1021_g N_A3_c_339_n
+ N_A3_M1024_g N_A3_c_330_n N_A3_M1031_g N_A3_c_340_n N_A3_M1028_g N_A3_c_331_n
+ N_A3_M1034_g N_A3_c_332_n N_A3_M1037_g A3 A3 A3 A3 N_A3_c_334_n
+ PM_SKY130_FD_SC_MS__O41AI_4%A3
x_PM_SKY130_FD_SC_MS__O41AI_4%A2 N_A2_c_430_n N_A2_M1002_g N_A2_M1013_g
+ N_A2_c_432_n N_A2_M1011_g N_A2_M1016_g N_A2_c_434_n N_A2_M1014_g N_A2_M1019_g
+ N_A2_c_436_n N_A2_M1027_g N_A2_M1022_g A2 A2 A2 A2 N_A2_c_439_n
+ PM_SKY130_FD_SC_MS__O41AI_4%A2
x_PM_SKY130_FD_SC_MS__O41AI_4%A1 N_A1_M1025_g N_A1_c_528_n N_A1_M1005_g
+ N_A1_M1026_g N_A1_c_530_n N_A1_M1006_g N_A1_M1035_g N_A1_c_532_n N_A1_M1032_g
+ N_A1_c_533_n N_A1_M1036_g N_A1_c_535_n N_A1_M1033_g A1 A1 A1 A1
+ PM_SKY130_FD_SC_MS__O41AI_4%A1
x_PM_SKY130_FD_SC_MS__O41AI_4%VPWR N_VPWR_M1004_d N_VPWR_M1008_d N_VPWR_M1025_d
+ N_VPWR_M1035_d N_VPWR_c_609_n N_VPWR_c_610_n N_VPWR_c_611_n N_VPWR_c_612_n
+ N_VPWR_c_613_n VPWR N_VPWR_c_614_n N_VPWR_c_615_n N_VPWR_c_616_n
+ N_VPWR_c_617_n N_VPWR_c_608_n N_VPWR_c_619_n N_VPWR_c_620_n N_VPWR_c_621_n
+ PM_SKY130_FD_SC_MS__O41AI_4%VPWR
x_PM_SKY130_FD_SC_MS__O41AI_4%Y N_Y_M1009_s N_Y_M1029_s N_Y_M1004_s N_Y_M1015_d
+ N_Y_M1020_d N_Y_c_716_n N_Y_c_724_n N_Y_c_717_n N_Y_c_718_n N_Y_c_734_n
+ N_Y_c_715_n N_Y_c_720_n N_Y_c_741_n N_Y_c_721_n N_Y_c_749_n Y Y N_Y_c_759_n
+ PM_SKY130_FD_SC_MS__O41AI_4%Y
x_PM_SKY130_FD_SC_MS__O41AI_4%A_339_368# N_A_339_368#_M1015_s
+ N_A_339_368#_M1018_s N_A_339_368#_M1023_s N_A_339_368#_M1021_d
+ N_A_339_368#_M1028_d N_A_339_368#_c_795_n N_A_339_368#_c_796_n
+ N_A_339_368#_c_797_n N_A_339_368#_c_813_n N_A_339_368#_c_798_n
+ N_A_339_368#_c_799_n N_A_339_368#_c_800_n N_A_339_368#_c_830_n
+ N_A_339_368#_c_801_n N_A_339_368#_c_802_n N_A_339_368#_c_803_n
+ N_A_339_368#_c_804_n N_A_339_368#_c_805_n
+ PM_SKY130_FD_SC_MS__O41AI_4%A_339_368#
x_PM_SKY130_FD_SC_MS__O41AI_4%A_791_368# N_A_791_368#_M1003_s
+ N_A_791_368#_M1024_s N_A_791_368#_M1013_d N_A_791_368#_M1019_d
+ N_A_791_368#_c_918_n N_A_791_368#_c_893_n N_A_791_368#_c_889_n
+ N_A_791_368#_c_922_n N_A_791_368#_c_890_n N_A_791_368#_c_929_p
+ N_A_791_368#_c_891_n N_A_791_368#_c_932_p N_A_791_368#_c_903_n
+ N_A_791_368#_c_892_n PM_SKY130_FD_SC_MS__O41AI_4%A_791_368#
x_PM_SKY130_FD_SC_MS__O41AI_4%A_1191_368# N_A_1191_368#_M1013_s
+ N_A_1191_368#_M1016_s N_A_1191_368#_M1022_s N_A_1191_368#_M1026_s
+ N_A_1191_368#_M1036_s N_A_1191_368#_c_935_n N_A_1191_368#_c_936_n
+ N_A_1191_368#_c_937_n N_A_1191_368#_c_953_n N_A_1191_368#_c_938_n
+ N_A_1191_368#_c_959_n N_A_1191_368#_c_939_n N_A_1191_368#_c_940_n
+ N_A_1191_368#_c_941_n N_A_1191_368#_c_942_n N_A_1191_368#_c_943_n
+ N_A_1191_368#_c_944_n N_A_1191_368#_c_945_n
+ PM_SKY130_FD_SC_MS__O41AI_4%A_1191_368#
x_PM_SKY130_FD_SC_MS__O41AI_4%A_27_74# N_A_27_74#_M1009_d N_A_27_74#_M1010_d
+ N_A_27_74#_M1030_d N_A_27_74#_M1007_s N_A_27_74#_M1017_s N_A_27_74#_M1031_s
+ N_A_27_74#_M1037_s N_A_27_74#_M1011_d N_A_27_74#_M1027_d N_A_27_74#_M1006_d
+ N_A_27_74#_M1033_d N_A_27_74#_c_1016_n N_A_27_74#_c_1017_n N_A_27_74#_c_1018_n
+ N_A_27_74#_c_1019_n N_A_27_74#_c_1047_n N_A_27_74#_c_1048_n
+ N_A_27_74#_c_1052_n N_A_27_74#_c_1020_n N_A_27_74#_c_1021_n
+ N_A_27_74#_c_1022_n N_A_27_74#_c_1063_n N_A_27_74#_c_1023_n
+ N_A_27_74#_c_1024_n N_A_27_74#_c_1079_n N_A_27_74#_c_1025_n
+ N_A_27_74#_c_1086_n N_A_27_74#_c_1026_n N_A_27_74#_c_1099_n
+ N_A_27_74#_c_1027_n N_A_27_74#_c_1105_n N_A_27_74#_c_1028_n
+ N_A_27_74#_c_1115_n N_A_27_74#_c_1029_n N_A_27_74#_c_1123_n
+ N_A_27_74#_c_1030_n N_A_27_74#_c_1031_n N_A_27_74#_c_1032_n
+ N_A_27_74#_c_1068_n N_A_27_74#_c_1070_n N_A_27_74#_c_1093_n
+ N_A_27_74#_c_1096_n N_A_27_74#_c_1111_n N_A_27_74#_c_1113_n
+ N_A_27_74#_c_1129_n PM_SKY130_FD_SC_MS__O41AI_4%A_27_74#
x_PM_SKY130_FD_SC_MS__O41AI_4%VGND N_VGND_M1000_d N_VGND_M1012_d N_VGND_M1001_d
+ N_VGND_M1034_d N_VGND_M1002_s N_VGND_M1014_s N_VGND_M1005_s N_VGND_M1032_s
+ N_VGND_c_1206_n N_VGND_c_1207_n N_VGND_c_1208_n N_VGND_c_1209_n
+ N_VGND_c_1210_n N_VGND_c_1211_n N_VGND_c_1212_n N_VGND_c_1213_n
+ N_VGND_c_1214_n N_VGND_c_1215_n N_VGND_c_1216_n VGND N_VGND_c_1217_n
+ N_VGND_c_1218_n N_VGND_c_1219_n N_VGND_c_1220_n N_VGND_c_1221_n
+ N_VGND_c_1222_n N_VGND_c_1223_n N_VGND_c_1224_n N_VGND_c_1225_n
+ N_VGND_c_1226_n N_VGND_c_1227_n N_VGND_c_1228_n N_VGND_c_1229_n
+ PM_SKY130_FD_SC_MS__O41AI_4%VGND
cc_1 VNB N_B1_M1004_g 0.00959774f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_B1_c_156_n 0.0185832f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.185
cc_3 VNB N_B1_c_157_n 0.0143157f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.185
cc_4 VNB N_B1_M1008_g 0.00713352f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.4
cc_5 VNB N_B1_c_159_n 0.0149371f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.185
cc_6 VNB N_B1_c_160_n 0.0298945f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.26
cc_7 VNB N_B1_c_161_n 0.09435f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=1.26
cc_8 VNB N_B1_c_162_n 0.0152736f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.185
cc_9 VNB N_B1_c_163_n 0.0259935f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.385
cc_10 VNB N_A4_c_223_n 0.0173669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A4_c_224_n 0.0173529f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.4
cc_12 VNB N_A4_c_225_n 0.0151591f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=1.26
cc_13 VNB N_A4_c_226_n 0.0185585f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=0.74
cc_14 VNB N_A4_c_227_n 0.120341f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_15 VNB N_A4_c_228_n 0.0151037f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_16 VNB N_A4_c_229_n 0.0115136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A3_c_327_n 0.0124747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A3_c_328_n 0.00656097f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.185
cc_19 VNB N_A3_c_329_n 0.0178826f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_20 VNB N_A3_c_330_n 0.0168239f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.185
cc_21 VNB N_A3_c_331_n 0.0173859f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=0.74
cc_22 VNB N_A3_c_332_n 0.0171629f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_23 VNB A3 0.0173798f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.367
cc_24 VNB N_A3_c_334_n 0.113711f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.365
cc_25 VNB N_A2_c_430_n 0.0180414f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.55
cc_26 VNB N_A2_M1013_g 0.00916985f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_27 VNB N_A2_c_432_n 0.0168231f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.185
cc_28 VNB N_A2_M1016_g 0.0057996f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.4
cc_29 VNB N_A2_c_434_n 0.0165146f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=1.185
cc_30 VNB N_A2_M1019_g 0.0057996f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.185
cc_31 VNB N_A2_c_436_n 0.0179931f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=0.74
cc_32 VNB N_A2_M1022_g 0.00599907f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=1.367
cc_33 VNB A2 0.0177499f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.367
cc_34 VNB N_A2_c_439_n 0.0877756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A1_M1025_g 0.00108424f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_36 VNB N_A1_c_528_n 0.0181973f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.185
cc_37 VNB N_A1_M1026_g 0.00602065f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_38 VNB N_A1_c_530_n 0.0175147f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.4
cc_39 VNB N_A1_M1035_g 0.00602065f $X=-0.19 $Y=-0.245 $X2=1.355 $Y2=0.74
cc_40 VNB N_A1_c_532_n 0.0173888f $X=-0.19 $Y=-0.245 $X2=1.43 $Y2=1.26
cc_41 VNB N_A1_c_533_n 0.100419f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=0.74
cc_42 VNB N_A1_M1036_g 0.0093909f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_43 VNB N_A1_c_535_n 0.0228112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB A1 0.0307917f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.367
cc_45 VNB N_VPWR_c_608_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_Y_c_715_n 0.00830153f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=1.367
cc_47 VNB N_A_27_74#_c_1016_n 0.0226322f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.367
cc_48 VNB N_A_27_74#_c_1017_n 0.00199363f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.365
cc_49 VNB N_A_27_74#_c_1018_n 0.00971634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_27_74#_c_1019_n 0.00502562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_27_74#_c_1020_n 0.0028074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_27_74#_c_1021_n 6.81442e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_27_74#_c_1022_n 0.00753795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_27_74#_c_1023_n 0.00240128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_27_74#_c_1024_n 0.00140577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_27_74#_c_1025_n 0.00206561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_27_74#_c_1026_n 0.00206561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_27_74#_c_1027_n 0.00178829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_27_74#_c_1028_n 0.00253253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_27_74#_c_1029_n 0.0024006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_27_74#_c_1030_n 0.0075085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_27_74#_c_1031_n 0.0203664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_27_74#_c_1032_n 0.00202117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1206_n 0.00933987f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=1.367
cc_65 VNB N_VGND_c_1207_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=1.385
cc_66 VNB N_VGND_c_1208_n 0.00578139f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.367
cc_67 VNB N_VGND_c_1209_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.385
cc_68 VNB N_VGND_c_1210_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1211_n 0.00485164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1212_n 0.00498382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1213_n 0.00528272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1214_n 0.00571618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1215_n 0.0189539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1216_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1217_n 0.0809332f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1218_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1219_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1220_n 0.018048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1221_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1222_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1223_n 0.507588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1224_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1225_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1226_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1227_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1228_n 0.00617178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1229_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VPB N_B1_M1004_g 0.0301521f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_89 VPB N_B1_M1008_g 0.0263526f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.4
cc_90 VPB N_A4_c_230_n 0.020867f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.55
cc_91 VPB N_A4_c_231_n 0.0170611f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_92 VPB N_A4_c_232_n 0.0170611f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_93 VPB N_A4_c_233_n 0.0175526f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.74
cc_94 VPB N_A4_c_227_n 0.0211094f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_95 VPB N_A3_c_335_n 0.018911f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.55
cc_96 VPB N_A3_c_327_n 0.00798007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A3_c_328_n 0.00251844f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.185
cc_98 VPB N_A3_c_338_n 0.0179762f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_99 VPB N_A3_c_339_n 0.0170611f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.4
cc_100 VPB N_A3_c_340_n 0.0210531f $X=-0.19 $Y=1.66 $X2=1.78 $Y2=1.26
cc_101 VPB N_A3_c_334_n 0.0159625f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.365
cc_102 VPB N_A2_M1013_g 0.0264878f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_103 VPB N_A2_M1016_g 0.0205309f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.4
cc_104 VPB N_A2_M1019_g 0.0205309f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.185
cc_105 VPB N_A2_M1022_g 0.0211645f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=1.367
cc_106 VPB N_A1_M1025_g 0.0217357f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_107 VPB N_A1_M1026_g 0.0219153f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_108 VPB N_A1_M1035_g 0.0219153f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=0.74
cc_109 VPB N_A1_M1036_g 0.028082f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_110 VPB N_VPWR_c_609_n 0.0119967f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=2.4
cc_111 VPB N_VPWR_c_610_n 0.0553391f $X=-0.19 $Y=1.66 $X2=1.355 $Y2=1.185
cc_112 VPB N_VPWR_c_611_n 0.0139267f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=0.74
cc_113 VPB N_VPWR_c_612_n 0.00559929f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_613_n 0.00559929f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=1.385
cc_115 VPB N_VPWR_c_614_n 0.0183788f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.367
cc_116 VPB N_VPWR_c_615_n 0.154956f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.365
cc_117 VPB N_VPWR_c_616_n 0.0185924f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_617_n 0.0177062f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_608_n 0.105088f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_619_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_620_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_621_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_Y_c_716_n 0.00326394f $X=-0.19 $Y=1.66 $X2=1.78 $Y2=1.26
cc_124 VPB N_Y_c_717_n 0.0059192f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_125 VPB N_Y_c_718_n 0.0043231f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_Y_c_715_n 0.00201193f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=1.367
cc_127 VPB N_Y_c_720_n 0.00297633f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=1.385
cc_128 VPB N_Y_c_721_n 0.0101507f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=1.365
cc_129 VPB N_A_339_368#_c_795_n 0.00761891f $X=-0.19 $Y=1.66 $X2=1.78 $Y2=1.26
cc_130 VPB N_A_339_368#_c_796_n 0.00192243f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.185
cc_131 VPB N_A_339_368#_c_797_n 0.00413156f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=0.74
cc_132 VPB N_A_339_368#_c_798_n 0.00192243f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_339_368#_c_799_n 0.00245929f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.367
cc_134 VPB N_A_339_368#_c_800_n 0.0026766f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.385
cc_135 VPB N_A_339_368#_c_801_n 0.00605183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_339_368#_c_802_n 0.00759021f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.365
cc_137 VPB N_A_339_368#_c_803_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_339_368#_c_804_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_339_368#_c_805_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_791_368#_c_889_n 9.51563e-19 $X=-0.19 $Y=1.66 $X2=1.78 $Y2=1.26
cc_141 VPB N_A_791_368#_c_890_n 0.0188562f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_142 VPB N_A_791_368#_c_891_n 0.00535008f $X=-0.19 $Y=1.66 $X2=0.3 $Y2=1.385
cc_143 VPB N_A_791_368#_c_892_n 0.00186725f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.367
cc_144 VPB N_A_1191_368#_c_935_n 0.00749658f $X=-0.19 $Y=1.66 $X2=1.78 $Y2=1.26
cc_145 VPB N_A_1191_368#_c_936_n 0.00192524f $X=-0.19 $Y=1.66 $X2=1.855
+ $Y2=1.185
cc_146 VPB N_A_1191_368#_c_937_n 0.00426372f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=0.74
cc_147 VPB N_A_1191_368#_c_938_n 0.00467254f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_1191_368#_c_939_n 0.00443091f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.385
cc_149 VPB N_A_1191_368#_c_940_n 0.00234762f $X=-0.19 $Y=1.66 $X2=0.98 $Y2=1.385
cc_150 VPB N_A_1191_368#_c_941_n 0.00223845f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.365
cc_151 VPB N_A_1191_368#_c_942_n 0.0131052f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.365
cc_152 VPB N_A_1191_368#_c_943_n 0.0441882f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_1191_368#_c_944_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_1191_368#_c_945_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 N_B1_c_162_n N_A4_c_223_n 0.0177689f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_156 N_B1_c_160_n N_A4_c_227_n 0.00932861f $X=1.78 $Y=1.26 $X2=0 $Y2=0
cc_157 N_B1_c_162_n N_A4_c_229_n 0.00137652f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_158 N_B1_M1004_g N_VPWR_c_610_n 0.0205921f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_159 N_B1_M1008_g N_VPWR_c_610_n 5.94268e-19 $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_160 N_B1_c_161_n N_VPWR_c_610_n 0.00628686f $X=1.43 $Y=1.26 $X2=0 $Y2=0
cc_161 N_B1_c_163_n N_VPWR_c_610_n 0.019114f $X=0.98 $Y=1.385 $X2=0 $Y2=0
cc_162 N_B1_M1004_g N_VPWR_c_611_n 5.34972e-19 $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_163 N_B1_M1008_g N_VPWR_c_611_n 0.0203923f $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_164 N_B1_M1004_g N_VPWR_c_614_n 0.00460063f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_165 N_B1_M1008_g N_VPWR_c_614_n 0.00460063f $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_166 N_B1_M1004_g N_VPWR_c_608_n 0.00909486f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_167 N_B1_M1008_g N_VPWR_c_608_n 0.00909486f $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_168 N_B1_M1004_g N_Y_c_716_n 4.86047e-19 $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_169 N_B1_M1008_g N_Y_c_716_n 4.86047e-19 $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_170 N_B1_c_157_n N_Y_c_724_n 0.00955428f $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_171 N_B1_c_159_n N_Y_c_724_n 0.015868f $X=1.355 $Y=1.185 $X2=0 $Y2=0
cc_172 N_B1_c_161_n N_Y_c_724_n 0.00190994f $X=1.43 $Y=1.26 $X2=0 $Y2=0
cc_173 N_B1_c_163_n N_Y_c_724_n 0.0224794f $X=0.98 $Y=1.385 $X2=0 $Y2=0
cc_174 N_B1_M1008_g N_Y_c_717_n 0.017948f $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_175 N_B1_c_161_n N_Y_c_717_n 0.0106118f $X=1.43 $Y=1.26 $X2=0 $Y2=0
cc_176 N_B1_c_163_n N_Y_c_717_n 0.0144526f $X=0.98 $Y=1.385 $X2=0 $Y2=0
cc_177 N_B1_M1004_g N_Y_c_718_n 0.00365076f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_178 N_B1_c_161_n N_Y_c_718_n 0.00491508f $X=1.43 $Y=1.26 $X2=0 $Y2=0
cc_179 N_B1_c_163_n N_Y_c_718_n 0.0280525f $X=0.98 $Y=1.385 $X2=0 $Y2=0
cc_180 N_B1_c_162_n N_Y_c_734_n 0.0054601f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_181 N_B1_c_159_n N_Y_c_715_n 0.00255143f $X=1.355 $Y=1.185 $X2=0 $Y2=0
cc_182 N_B1_c_160_n N_Y_c_715_n 0.0205092f $X=1.78 $Y=1.26 $X2=0 $Y2=0
cc_183 N_B1_c_161_n N_Y_c_715_n 0.00682632f $X=1.43 $Y=1.26 $X2=0 $Y2=0
cc_184 N_B1_c_162_n N_Y_c_715_n 0.0048483f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_185 N_B1_c_163_n N_Y_c_715_n 0.0181698f $X=0.98 $Y=1.385 $X2=0 $Y2=0
cc_186 N_B1_c_160_n N_Y_c_720_n 0.00411697f $X=1.78 $Y=1.26 $X2=0 $Y2=0
cc_187 N_B1_c_161_n N_Y_c_741_n 7.43006e-19 $X=1.43 $Y=1.26 $X2=0 $Y2=0
cc_188 N_B1_c_163_n N_Y_c_741_n 0.0140705f $X=0.98 $Y=1.385 $X2=0 $Y2=0
cc_189 N_B1_M1008_g N_A_339_368#_c_795_n 0.00189033f $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_190 N_B1_M1008_g N_A_339_368#_c_797_n 6.08298e-19 $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_191 N_B1_c_156_n N_A_27_74#_c_1016_n 0.00796844f $X=0.495 $Y=1.185 $X2=0
+ $Y2=0
cc_192 N_B1_c_157_n N_A_27_74#_c_1016_n 5.73078e-19 $X=0.925 $Y=1.185 $X2=0
+ $Y2=0
cc_193 N_B1_c_161_n N_A_27_74#_c_1016_n 0.00205251f $X=1.43 $Y=1.26 $X2=0 $Y2=0
cc_194 N_B1_c_163_n N_A_27_74#_c_1016_n 0.0251377f $X=0.98 $Y=1.385 $X2=0 $Y2=0
cc_195 N_B1_c_156_n N_A_27_74#_c_1017_n 0.0100711f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_196 N_B1_c_157_n N_A_27_74#_c_1017_n 0.00789822f $X=0.925 $Y=1.185 $X2=0
+ $Y2=0
cc_197 N_B1_c_156_n N_A_27_74#_c_1018_n 0.00282152f $X=0.495 $Y=1.185 $X2=0
+ $Y2=0
cc_198 N_B1_c_159_n N_A_27_74#_c_1019_n 0.00829147f $X=1.355 $Y=1.185 $X2=0
+ $Y2=0
cc_199 N_B1_c_162_n N_A_27_74#_c_1019_n 0.0137299f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_200 N_B1_c_156_n N_A_27_74#_c_1032_n 6.04287e-19 $X=0.495 $Y=1.185 $X2=0
+ $Y2=0
cc_201 N_B1_c_157_n N_A_27_74#_c_1032_n 0.00642184f $X=0.925 $Y=1.185 $X2=0
+ $Y2=0
cc_202 N_B1_c_159_n N_A_27_74#_c_1032_n 0.00684618f $X=1.355 $Y=1.185 $X2=0
+ $Y2=0
cc_203 N_B1_c_162_n N_A_27_74#_c_1032_n 6.66855e-19 $X=1.855 $Y=1.185 $X2=0
+ $Y2=0
cc_204 N_B1_c_156_n N_VGND_c_1217_n 0.00278247f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_205 N_B1_c_157_n N_VGND_c_1217_n 0.00279469f $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_206 N_B1_c_159_n N_VGND_c_1217_n 0.00279469f $X=1.355 $Y=1.185 $X2=0 $Y2=0
cc_207 N_B1_c_162_n N_VGND_c_1217_n 0.00278271f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_208 N_B1_c_156_n N_VGND_c_1223_n 0.00357084f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_209 N_B1_c_157_n N_VGND_c_1223_n 0.00352518f $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_210 N_B1_c_159_n N_VGND_c_1223_n 0.00353176f $X=1.355 $Y=1.185 $X2=0 $Y2=0
cc_211 N_B1_c_162_n N_VGND_c_1223_n 0.00354798f $X=1.855 $Y=1.185 $X2=0 $Y2=0
cc_212 N_A4_c_233_n N_A3_c_335_n 0.0127977f $X=3.415 $Y=1.725 $X2=-0.19
+ $Y2=-0.245
cc_213 N_A4_c_226_n N_A3_c_328_n 0.0149207f $X=3.895 $Y=1.26 $X2=0 $Y2=0
cc_214 N_A4_c_227_n N_A3_c_328_n 0.0127977f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_215 N_A4_c_228_n N_A3_c_329_n 0.00804366f $X=3.97 $Y=1.185 $X2=0 $Y2=0
cc_216 N_A4_c_226_n N_A3_c_334_n 0.00804366f $X=3.895 $Y=1.26 $X2=0 $Y2=0
cc_217 N_A4_c_230_n N_VPWR_c_611_n 0.00284685f $X=2.065 $Y=1.725 $X2=0 $Y2=0
cc_218 N_A4_c_230_n N_VPWR_c_615_n 0.00333921f $X=2.065 $Y=1.725 $X2=0 $Y2=0
cc_219 N_A4_c_231_n N_VPWR_c_615_n 0.00333921f $X=2.515 $Y=1.725 $X2=0 $Y2=0
cc_220 N_A4_c_232_n N_VPWR_c_615_n 0.00333921f $X=2.965 $Y=1.725 $X2=0 $Y2=0
cc_221 N_A4_c_233_n N_VPWR_c_615_n 0.00333921f $X=3.415 $Y=1.725 $X2=0 $Y2=0
cc_222 N_A4_c_230_n N_VPWR_c_608_n 0.00424184f $X=2.065 $Y=1.725 $X2=0 $Y2=0
cc_223 N_A4_c_231_n N_VPWR_c_608_n 0.00419051f $X=2.515 $Y=1.725 $X2=0 $Y2=0
cc_224 N_A4_c_232_n N_VPWR_c_608_n 0.00419051f $X=2.965 $Y=1.725 $X2=0 $Y2=0
cc_225 N_A4_c_233_n N_VPWR_c_608_n 0.00419162f $X=3.415 $Y=1.725 $X2=0 $Y2=0
cc_226 N_A4_c_223_n N_Y_c_715_n 5.71389e-19 $X=2.355 $Y=1.185 $X2=0 $Y2=0
cc_227 N_A4_c_227_n N_Y_c_715_n 0.00868138f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_228 N_A4_c_229_n N_Y_c_715_n 0.0248693f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_229 N_A4_c_230_n N_Y_c_720_n 0.0141359f $X=2.065 $Y=1.725 $X2=0 $Y2=0
cc_230 N_A4_c_227_n N_Y_c_720_n 0.00368436f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_231 N_A4_c_229_n N_Y_c_720_n 0.00796928f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_232 N_A4_c_230_n N_Y_c_749_n 0.0213574f $X=2.065 $Y=1.725 $X2=0 $Y2=0
cc_233 N_A4_c_231_n N_Y_c_749_n 0.0126519f $X=2.515 $Y=1.725 $X2=0 $Y2=0
cc_234 N_A4_c_232_n N_Y_c_749_n 4.21044e-19 $X=2.965 $Y=1.725 $X2=0 $Y2=0
cc_235 N_A4_c_227_n N_Y_c_749_n 0.00644625f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_236 N_A4_c_229_n N_Y_c_749_n 0.0225374f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_237 N_A4_c_231_n Y 4.21044e-19 $X=2.515 $Y=1.725 $X2=0 $Y2=0
cc_238 N_A4_c_232_n Y 0.0126519f $X=2.965 $Y=1.725 $X2=0 $Y2=0
cc_239 N_A4_c_233_n Y 0.0179904f $X=3.415 $Y=1.725 $X2=0 $Y2=0
cc_240 N_A4_c_227_n Y 0.0126784f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_241 N_A4_c_229_n Y 0.00885397f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_242 N_A4_c_231_n N_Y_c_759_n 0.0201953f $X=2.515 $Y=1.725 $X2=0 $Y2=0
cc_243 N_A4_c_232_n N_Y_c_759_n 0.0201953f $X=2.965 $Y=1.725 $X2=0 $Y2=0
cc_244 N_A4_c_227_n N_Y_c_759_n 0.0109996f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_245 N_A4_c_229_n N_Y_c_759_n 0.0478219f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_246 N_A4_c_230_n N_A_339_368#_c_795_n 0.0166317f $X=2.065 $Y=1.725 $X2=0
+ $Y2=0
cc_247 N_A4_c_231_n N_A_339_368#_c_795_n 6.77408e-19 $X=2.515 $Y=1.725 $X2=0
+ $Y2=0
cc_248 N_A4_c_230_n N_A_339_368#_c_796_n 0.0130835f $X=2.065 $Y=1.725 $X2=0
+ $Y2=0
cc_249 N_A4_c_231_n N_A_339_368#_c_796_n 0.0130835f $X=2.515 $Y=1.725 $X2=0
+ $Y2=0
cc_250 N_A4_c_230_n N_A_339_368#_c_797_n 0.00239394f $X=2.065 $Y=1.725 $X2=0
+ $Y2=0
cc_251 N_A4_c_230_n N_A_339_368#_c_813_n 5.48759e-19 $X=2.065 $Y=1.725 $X2=0
+ $Y2=0
cc_252 N_A4_c_231_n N_A_339_368#_c_813_n 0.0086655f $X=2.515 $Y=1.725 $X2=0
+ $Y2=0
cc_253 N_A4_c_232_n N_A_339_368#_c_813_n 0.0086655f $X=2.965 $Y=1.725 $X2=0
+ $Y2=0
cc_254 N_A4_c_233_n N_A_339_368#_c_813_n 5.48759e-19 $X=3.415 $Y=1.725 $X2=0
+ $Y2=0
cc_255 N_A4_c_227_n N_A_339_368#_c_813_n 3.00056e-19 $X=3.615 $Y=1.26 $X2=0
+ $Y2=0
cc_256 N_A4_c_232_n N_A_339_368#_c_798_n 0.0130835f $X=2.965 $Y=1.725 $X2=0
+ $Y2=0
cc_257 N_A4_c_233_n N_A_339_368#_c_798_n 0.0130393f $X=3.415 $Y=1.725 $X2=0
+ $Y2=0
cc_258 N_A4_c_232_n N_A_339_368#_c_799_n 7.59096e-19 $X=2.965 $Y=1.725 $X2=0
+ $Y2=0
cc_259 N_A4_c_233_n N_A_339_368#_c_799_n 0.0171693f $X=3.415 $Y=1.725 $X2=0
+ $Y2=0
cc_260 N_A4_c_227_n N_A_339_368#_c_799_n 0.00152446f $X=3.615 $Y=1.26 $X2=0
+ $Y2=0
cc_261 N_A4_c_231_n N_A_339_368#_c_803_n 0.00141876f $X=2.515 $Y=1.725 $X2=0
+ $Y2=0
cc_262 N_A4_c_232_n N_A_339_368#_c_803_n 0.00141876f $X=2.965 $Y=1.725 $X2=0
+ $Y2=0
cc_263 N_A4_c_233_n N_A_339_368#_c_804_n 0.00139249f $X=3.415 $Y=1.725 $X2=0
+ $Y2=0
cc_264 N_A4_c_223_n N_A_27_74#_c_1019_n 0.00353966f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_265 N_A4_c_223_n N_A_27_74#_c_1047_n 0.0124539f $X=2.355 $Y=1.185 $X2=0 $Y2=0
cc_266 N_A4_c_223_n N_A_27_74#_c_1048_n 0.00979933f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_267 N_A4_c_224_n N_A_27_74#_c_1048_n 0.0111145f $X=3.085 $Y=1.185 $X2=0 $Y2=0
cc_268 N_A4_c_227_n N_A_27_74#_c_1048_n 0.00274914f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_269 N_A4_c_229_n N_A_27_74#_c_1048_n 0.0612456f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_270 N_A4_c_223_n N_A_27_74#_c_1052_n 7.32094e-19 $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_271 N_A4_c_227_n N_A_27_74#_c_1052_n 0.00304121f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_272 N_A4_c_229_n N_A_27_74#_c_1052_n 0.0199556f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_273 N_A4_c_224_n N_A_27_74#_c_1020_n 2.68164e-19 $X=3.085 $Y=1.185 $X2=0
+ $Y2=0
cc_274 N_A4_c_225_n N_A_27_74#_c_1020_n 0.00604445f $X=3.54 $Y=1.185 $X2=0 $Y2=0
cc_275 N_A4_c_224_n N_A_27_74#_c_1021_n 0.0032036f $X=3.085 $Y=1.185 $X2=0 $Y2=0
cc_276 N_A4_c_225_n N_A_27_74#_c_1021_n 0.00281435f $X=3.54 $Y=1.185 $X2=0 $Y2=0
cc_277 N_A4_c_227_n N_A_27_74#_c_1021_n 0.00726193f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_278 N_A4_c_229_n N_A_27_74#_c_1021_n 0.00900371f $X=2.995 $Y=1.385 $X2=0
+ $Y2=0
cc_279 N_A4_c_226_n N_A_27_74#_c_1022_n 0.018043f $X=3.895 $Y=1.26 $X2=0 $Y2=0
cc_280 N_A4_c_227_n N_A_27_74#_c_1022_n 0.0105089f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_281 N_A4_c_227_n N_A_27_74#_c_1063_n 0.0139f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_282 N_A4_c_229_n N_A_27_74#_c_1063_n 0.0143906f $X=2.995 $Y=1.385 $X2=0 $Y2=0
cc_283 N_A4_c_228_n N_A_27_74#_c_1023_n 0.00574886f $X=3.97 $Y=1.185 $X2=0 $Y2=0
cc_284 N_A4_c_226_n N_A_27_74#_c_1024_n 0.00388347f $X=3.895 $Y=1.26 $X2=0 $Y2=0
cc_285 N_A4_c_228_n N_A_27_74#_c_1024_n 0.00267912f $X=3.97 $Y=1.185 $X2=0 $Y2=0
cc_286 N_A4_c_225_n N_A_27_74#_c_1068_n 0.00184154f $X=3.54 $Y=1.185 $X2=0 $Y2=0
cc_287 N_A4_c_227_n N_A_27_74#_c_1068_n 0.00381215f $X=3.615 $Y=1.26 $X2=0 $Y2=0
cc_288 N_A4_c_228_n N_A_27_74#_c_1070_n 0.0017646f $X=3.97 $Y=1.185 $X2=0 $Y2=0
cc_289 N_A4_c_225_n N_VGND_c_1206_n 0.00313396f $X=3.54 $Y=1.185 $X2=0 $Y2=0
cc_290 N_A4_c_226_n N_VGND_c_1206_n 0.00230361f $X=3.895 $Y=1.26 $X2=0 $Y2=0
cc_291 N_A4_c_228_n N_VGND_c_1206_n 0.00313962f $X=3.97 $Y=1.185 $X2=0 $Y2=0
cc_292 N_A4_c_228_n N_VGND_c_1207_n 0.00434272f $X=3.97 $Y=1.185 $X2=0 $Y2=0
cc_293 N_A4_c_224_n N_VGND_c_1215_n 0.00461464f $X=3.085 $Y=1.185 $X2=0 $Y2=0
cc_294 N_A4_c_225_n N_VGND_c_1215_n 0.00422942f $X=3.54 $Y=1.185 $X2=0 $Y2=0
cc_295 N_A4_c_223_n N_VGND_c_1217_n 0.00789845f $X=2.355 $Y=1.185 $X2=0 $Y2=0
cc_296 N_A4_c_224_n N_VGND_c_1217_n 0.00590535f $X=3.085 $Y=1.185 $X2=0 $Y2=0
cc_297 N_A4_c_223_n N_VGND_c_1223_n 0.00447853f $X=2.355 $Y=1.185 $X2=0 $Y2=0
cc_298 N_A4_c_224_n N_VGND_c_1223_n 0.00465356f $X=3.085 $Y=1.185 $X2=0 $Y2=0
cc_299 N_A4_c_225_n N_VGND_c_1223_n 0.00783843f $X=3.54 $Y=1.185 $X2=0 $Y2=0
cc_300 N_A4_c_228_n N_VGND_c_1223_n 0.00820382f $X=3.97 $Y=1.185 $X2=0 $Y2=0
cc_301 N_A3_c_332_n N_A2_c_430_n 0.00936575f $X=5.83 $Y=1.22 $X2=-0.19
+ $Y2=-0.245
cc_302 A3 N_A2_c_430_n 0.0044767f $X=5.915 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_303 A3 A2 0.0247108f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_304 N_A3_c_334_n A2 2.21735e-19 $X=5.58 $Y=1.385 $X2=0 $Y2=0
cc_305 N_A3_c_334_n N_A2_c_439_n 0.0132359f $X=5.58 $Y=1.385 $X2=0 $Y2=0
cc_306 N_A3_c_335_n N_VPWR_c_615_n 0.00333896f $X=3.865 $Y=1.725 $X2=0 $Y2=0
cc_307 N_A3_c_338_n N_VPWR_c_615_n 0.00333896f $X=4.415 $Y=1.725 $X2=0 $Y2=0
cc_308 N_A3_c_339_n N_VPWR_c_615_n 0.00333896f $X=4.865 $Y=1.725 $X2=0 $Y2=0
cc_309 N_A3_c_340_n N_VPWR_c_615_n 0.00333896f $X=5.315 $Y=1.725 $X2=0 $Y2=0
cc_310 N_A3_c_335_n N_VPWR_c_608_n 0.00423728f $X=3.865 $Y=1.725 $X2=0 $Y2=0
cc_311 N_A3_c_338_n N_VPWR_c_608_n 0.00423617f $X=4.415 $Y=1.725 $X2=0 $Y2=0
cc_312 N_A3_c_339_n N_VPWR_c_608_n 0.00422685f $X=4.865 $Y=1.725 $X2=0 $Y2=0
cc_313 N_A3_c_340_n N_VPWR_c_608_n 0.00427818f $X=5.315 $Y=1.725 $X2=0 $Y2=0
cc_314 N_A3_c_328_n Y 2.28955e-19 $X=3.955 $Y=1.65 $X2=0 $Y2=0
cc_315 N_A3_c_335_n N_A_339_368#_c_799_n 0.0160548f $X=3.865 $Y=1.725 $X2=0
+ $Y2=0
cc_316 N_A3_c_338_n N_A_339_368#_c_799_n 6.74102e-19 $X=4.415 $Y=1.725 $X2=0
+ $Y2=0
cc_317 N_A3_c_335_n N_A_339_368#_c_800_n 0.0121897f $X=3.865 $Y=1.725 $X2=0
+ $Y2=0
cc_318 N_A3_c_338_n N_A_339_368#_c_800_n 0.0121897f $X=4.415 $Y=1.725 $X2=0
+ $Y2=0
cc_319 N_A3_c_335_n N_A_339_368#_c_830_n 5.96905e-19 $X=3.865 $Y=1.725 $X2=0
+ $Y2=0
cc_320 N_A3_c_338_n N_A_339_368#_c_830_n 0.015148f $X=4.415 $Y=1.725 $X2=0 $Y2=0
cc_321 N_A3_c_339_n N_A_339_368#_c_830_n 0.0146914f $X=4.865 $Y=1.725 $X2=0
+ $Y2=0
cc_322 N_A3_c_340_n N_A_339_368#_c_830_n 6.15772e-19 $X=5.315 $Y=1.725 $X2=0
+ $Y2=0
cc_323 N_A3_c_334_n N_A_339_368#_c_830_n 4.79751e-19 $X=5.58 $Y=1.385 $X2=0
+ $Y2=0
cc_324 N_A3_c_339_n N_A_339_368#_c_801_n 0.0116345f $X=4.865 $Y=1.725 $X2=0
+ $Y2=0
cc_325 N_A3_c_340_n N_A_339_368#_c_801_n 0.014552f $X=5.315 $Y=1.725 $X2=0 $Y2=0
cc_326 N_A3_c_339_n N_A_339_368#_c_802_n 6.15772e-19 $X=4.865 $Y=1.725 $X2=0
+ $Y2=0
cc_327 N_A3_c_340_n N_A_339_368#_c_802_n 0.017253f $X=5.315 $Y=1.725 $X2=0 $Y2=0
cc_328 N_A3_c_335_n N_A_339_368#_c_804_n 0.001916f $X=3.865 $Y=1.725 $X2=0 $Y2=0
cc_329 N_A3_c_338_n N_A_339_368#_c_805_n 0.00194226f $X=4.415 $Y=1.725 $X2=0
+ $Y2=0
cc_330 N_A3_c_339_n N_A_339_368#_c_805_n 0.00194226f $X=4.865 $Y=1.725 $X2=0
+ $Y2=0
cc_331 N_A3_c_327_n N_A_791_368#_c_893_n 6.90257e-19 $X=4.325 $Y=1.65 $X2=0
+ $Y2=0
cc_332 N_A3_c_338_n N_A_791_368#_c_893_n 0.0132979f $X=4.415 $Y=1.725 $X2=0
+ $Y2=0
cc_333 N_A3_c_339_n N_A_791_368#_c_893_n 0.0129823f $X=4.865 $Y=1.725 $X2=0
+ $Y2=0
cc_334 A3 N_A_791_368#_c_893_n 0.0417698f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_335 N_A3_c_334_n N_A_791_368#_c_893_n 0.0128552f $X=5.58 $Y=1.385 $X2=0 $Y2=0
cc_336 N_A3_c_335_n N_A_791_368#_c_889_n 0.00186623f $X=3.865 $Y=1.725 $X2=0
+ $Y2=0
cc_337 N_A3_c_327_n N_A_791_368#_c_889_n 0.0123144f $X=4.325 $Y=1.65 $X2=0 $Y2=0
cc_338 N_A3_c_340_n N_A_791_368#_c_890_n 0.0150422f $X=5.315 $Y=1.725 $X2=0
+ $Y2=0
cc_339 A3 N_A_791_368#_c_890_n 0.0697636f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_340 N_A3_c_334_n N_A_791_368#_c_890_n 0.0118396f $X=5.58 $Y=1.385 $X2=0 $Y2=0
cc_341 A3 N_A_791_368#_c_903_n 0.0185129f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_342 N_A3_c_334_n N_A_791_368#_c_903_n 0.0056879f $X=5.58 $Y=1.385 $X2=0 $Y2=0
cc_343 N_A3_c_340_n N_A_1191_368#_c_935_n 0.00211027f $X=5.315 $Y=1.725 $X2=0
+ $Y2=0
cc_344 N_A3_c_340_n N_A_1191_368#_c_937_n 6.38202e-19 $X=5.315 $Y=1.725 $X2=0
+ $Y2=0
cc_345 N_A3_c_327_n N_A_27_74#_c_1022_n 0.00358745f $X=4.325 $Y=1.65 $X2=0 $Y2=0
cc_346 N_A3_c_328_n N_A_27_74#_c_1022_n 0.00462373f $X=3.955 $Y=1.65 $X2=0 $Y2=0
cc_347 A3 N_A_27_74#_c_1022_n 0.013152f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_348 N_A3_c_334_n N_A_27_74#_c_1022_n 0.00422915f $X=5.58 $Y=1.385 $X2=0 $Y2=0
cc_349 N_A3_c_329_n N_A_27_74#_c_1023_n 0.00722697f $X=4.4 $Y=1.22 $X2=0 $Y2=0
cc_350 N_A3_c_330_n N_A_27_74#_c_1023_n 7.0998e-19 $X=4.9 $Y=1.22 $X2=0 $Y2=0
cc_351 N_A3_c_329_n N_A_27_74#_c_1024_n 0.00418933f $X=4.4 $Y=1.22 $X2=0 $Y2=0
cc_352 A3 N_A_27_74#_c_1024_n 0.00818182f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_353 N_A3_c_329_n N_A_27_74#_c_1079_n 0.010267f $X=4.4 $Y=1.22 $X2=0 $Y2=0
cc_354 N_A3_c_330_n N_A_27_74#_c_1079_n 0.0100105f $X=4.9 $Y=1.22 $X2=0 $Y2=0
cc_355 A3 N_A_27_74#_c_1079_n 0.0422704f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_356 N_A3_c_334_n N_A_27_74#_c_1079_n 0.00106284f $X=5.58 $Y=1.385 $X2=0 $Y2=0
cc_357 N_A3_c_330_n N_A_27_74#_c_1025_n 2.29136e-19 $X=4.9 $Y=1.22 $X2=0 $Y2=0
cc_358 N_A3_c_331_n N_A_27_74#_c_1025_n 0.00703259f $X=5.33 $Y=1.22 $X2=0 $Y2=0
cc_359 N_A3_c_332_n N_A_27_74#_c_1025_n 7.13338e-19 $X=5.83 $Y=1.22 $X2=0 $Y2=0
cc_360 N_A3_c_331_n N_A_27_74#_c_1086_n 0.00892313f $X=5.33 $Y=1.22 $X2=0 $Y2=0
cc_361 N_A3_c_332_n N_A_27_74#_c_1086_n 0.0100105f $X=5.83 $Y=1.22 $X2=0 $Y2=0
cc_362 A3 N_A_27_74#_c_1086_n 0.0454799f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_363 N_A3_c_334_n N_A_27_74#_c_1086_n 0.00107356f $X=5.58 $Y=1.385 $X2=0 $Y2=0
cc_364 N_A3_c_332_n N_A_27_74#_c_1026_n 2.29136e-19 $X=5.83 $Y=1.22 $X2=0 $Y2=0
cc_365 N_A3_c_327_n N_A_27_74#_c_1070_n 0.00315685f $X=4.325 $Y=1.65 $X2=0 $Y2=0
cc_366 N_A3_c_329_n N_A_27_74#_c_1070_n 0.00157416f $X=4.4 $Y=1.22 $X2=0 $Y2=0
cc_367 N_A3_c_331_n N_A_27_74#_c_1093_n 7.17169e-19 $X=5.33 $Y=1.22 $X2=0 $Y2=0
cc_368 A3 N_A_27_74#_c_1093_n 0.0189543f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_369 N_A3_c_334_n N_A_27_74#_c_1093_n 7.00387e-19 $X=5.58 $Y=1.385 $X2=0 $Y2=0
cc_370 A3 N_A_27_74#_c_1096_n 0.0134301f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_371 N_A3_c_329_n N_VGND_c_1207_n 0.00434272f $X=4.4 $Y=1.22 $X2=0 $Y2=0
cc_372 N_A3_c_329_n N_VGND_c_1208_n 0.00482414f $X=4.4 $Y=1.22 $X2=0 $Y2=0
cc_373 N_A3_c_330_n N_VGND_c_1208_n 0.00771106f $X=4.9 $Y=1.22 $X2=0 $Y2=0
cc_374 N_A3_c_331_n N_VGND_c_1208_n 4.39845e-19 $X=5.33 $Y=1.22 $X2=0 $Y2=0
cc_375 N_A3_c_330_n N_VGND_c_1209_n 0.00383152f $X=4.9 $Y=1.22 $X2=0 $Y2=0
cc_376 N_A3_c_331_n N_VGND_c_1209_n 0.00434272f $X=5.33 $Y=1.22 $X2=0 $Y2=0
cc_377 N_A3_c_331_n N_VGND_c_1210_n 0.00335277f $X=5.33 $Y=1.22 $X2=0 $Y2=0
cc_378 N_A3_c_332_n N_VGND_c_1210_n 0.00771106f $X=5.83 $Y=1.22 $X2=0 $Y2=0
cc_379 N_A3_c_332_n N_VGND_c_1218_n 0.00383152f $X=5.83 $Y=1.22 $X2=0 $Y2=0
cc_380 N_A3_c_329_n N_VGND_c_1223_n 0.00445593f $X=4.4 $Y=1.22 $X2=0 $Y2=0
cc_381 N_A3_c_330_n N_VGND_c_1223_n 0.00383967f $X=4.9 $Y=1.22 $X2=0 $Y2=0
cc_382 N_A3_c_331_n N_VGND_c_1223_n 0.00445496f $X=5.33 $Y=1.22 $X2=0 $Y2=0
cc_383 N_A3_c_332_n N_VGND_c_1223_n 0.00384065f $X=5.83 $Y=1.22 $X2=0 $Y2=0
cc_384 N_A2_c_436_n N_A1_c_528_n 0.00901198f $X=7.655 $Y=1.22 $X2=0 $Y2=0
cc_385 A2 N_A1_c_528_n 0.00453332f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_386 N_A2_M1022_g N_A1_c_533_n 0.0242466f $X=7.675 $Y=2.4 $X2=0 $Y2=0
cc_387 N_A2_c_439_n N_A1_c_533_n 0.0135263f $X=7.675 $Y=1.385 $X2=0 $Y2=0
cc_388 A2 A1 0.0247094f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_389 N_A2_c_439_n A1 2.11798e-19 $X=7.675 $Y=1.385 $X2=0 $Y2=0
cc_390 N_A2_M1022_g N_VPWR_c_612_n 4.4669e-19 $X=7.675 $Y=2.4 $X2=0 $Y2=0
cc_391 N_A2_M1013_g N_VPWR_c_615_n 0.00333896f $X=6.325 $Y=2.4 $X2=0 $Y2=0
cc_392 N_A2_M1016_g N_VPWR_c_615_n 0.00333896f $X=6.775 $Y=2.4 $X2=0 $Y2=0
cc_393 N_A2_M1019_g N_VPWR_c_615_n 0.00333896f $X=7.225 $Y=2.4 $X2=0 $Y2=0
cc_394 N_A2_M1022_g N_VPWR_c_615_n 0.00333896f $X=7.675 $Y=2.4 $X2=0 $Y2=0
cc_395 N_A2_M1013_g N_VPWR_c_608_n 0.00427818f $X=6.325 $Y=2.4 $X2=0 $Y2=0
cc_396 N_A2_M1016_g N_VPWR_c_608_n 0.00422685f $X=6.775 $Y=2.4 $X2=0 $Y2=0
cc_397 N_A2_M1019_g N_VPWR_c_608_n 0.00422685f $X=7.225 $Y=2.4 $X2=0 $Y2=0
cc_398 N_A2_M1022_g N_VPWR_c_608_n 0.00422796f $X=7.675 $Y=2.4 $X2=0 $Y2=0
cc_399 N_A2_M1013_g N_A_339_368#_c_801_n 6.06861e-19 $X=6.325 $Y=2.4 $X2=0 $Y2=0
cc_400 N_A2_M1013_g N_A_339_368#_c_802_n 0.00213642f $X=6.325 $Y=2.4 $X2=0 $Y2=0
cc_401 N_A2_M1013_g N_A_791_368#_c_890_n 0.0217401f $X=6.325 $Y=2.4 $X2=0 $Y2=0
cc_402 A2 N_A_791_368#_c_890_n 0.00508283f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_403 N_A2_c_439_n N_A_791_368#_c_890_n 0.00207531f $X=7.675 $Y=1.385 $X2=0
+ $Y2=0
cc_404 N_A2_M1016_g N_A_791_368#_c_891_n 0.0156079f $X=6.775 $Y=2.4 $X2=0 $Y2=0
cc_405 N_A2_M1019_g N_A_791_368#_c_891_n 0.0154829f $X=7.225 $Y=2.4 $X2=0 $Y2=0
cc_406 N_A2_M1022_g N_A_791_368#_c_891_n 0.00108804f $X=7.675 $Y=2.4 $X2=0 $Y2=0
cc_407 A2 N_A_791_368#_c_891_n 0.0689321f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_408 N_A2_c_439_n N_A_791_368#_c_891_n 0.00421298f $X=7.675 $Y=1.385 $X2=0
+ $Y2=0
cc_409 A2 N_A_791_368#_c_892_n 0.0195526f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_410 N_A2_c_439_n N_A_791_368#_c_892_n 0.00209661f $X=7.675 $Y=1.385 $X2=0
+ $Y2=0
cc_411 N_A2_M1013_g N_A_1191_368#_c_935_n 0.0170853f $X=6.325 $Y=2.4 $X2=0 $Y2=0
cc_412 N_A2_M1016_g N_A_1191_368#_c_935_n 6.11696e-19 $X=6.775 $Y=2.4 $X2=0
+ $Y2=0
cc_413 N_A2_M1013_g N_A_1191_368#_c_936_n 0.0120835f $X=6.325 $Y=2.4 $X2=0 $Y2=0
cc_414 N_A2_M1016_g N_A_1191_368#_c_936_n 0.0120835f $X=6.775 $Y=2.4 $X2=0 $Y2=0
cc_415 N_A2_M1013_g N_A_1191_368#_c_937_n 0.00295841f $X=6.325 $Y=2.4 $X2=0
+ $Y2=0
cc_416 N_A2_M1013_g N_A_1191_368#_c_953_n 6.11696e-19 $X=6.325 $Y=2.4 $X2=0
+ $Y2=0
cc_417 N_A2_M1016_g N_A_1191_368#_c_953_n 0.0145237f $X=6.775 $Y=2.4 $X2=0 $Y2=0
cc_418 N_A2_M1019_g N_A_1191_368#_c_953_n 0.0144041f $X=7.225 $Y=2.4 $X2=0 $Y2=0
cc_419 N_A2_M1022_g N_A_1191_368#_c_953_n 5.71937e-19 $X=7.675 $Y=2.4 $X2=0
+ $Y2=0
cc_420 N_A2_M1019_g N_A_1191_368#_c_938_n 0.0115958f $X=7.225 $Y=2.4 $X2=0 $Y2=0
cc_421 N_A2_M1022_g N_A_1191_368#_c_938_n 0.0133188f $X=7.675 $Y=2.4 $X2=0 $Y2=0
cc_422 N_A2_M1019_g N_A_1191_368#_c_959_n 6.63195e-19 $X=7.225 $Y=2.4 $X2=0
+ $Y2=0
cc_423 N_A2_M1022_g N_A_1191_368#_c_959_n 0.01352f $X=7.675 $Y=2.4 $X2=0 $Y2=0
cc_424 A2 N_A_1191_368#_c_939_n 0.00156259f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_425 N_A2_M1022_g N_A_1191_368#_c_940_n 0.00368403f $X=7.675 $Y=2.4 $X2=0
+ $Y2=0
cc_426 A2 N_A_1191_368#_c_940_n 0.0247125f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_427 N_A2_M1016_g N_A_1191_368#_c_944_n 0.00198322f $X=6.775 $Y=2.4 $X2=0
+ $Y2=0
cc_428 N_A2_M1019_g N_A_1191_368#_c_944_n 0.00223038f $X=7.225 $Y=2.4 $X2=0
+ $Y2=0
cc_429 N_A2_c_430_n N_A_27_74#_c_1026_n 0.00703259f $X=6.26 $Y=1.22 $X2=0 $Y2=0
cc_430 N_A2_c_432_n N_A_27_74#_c_1026_n 7.13338e-19 $X=6.76 $Y=1.22 $X2=0 $Y2=0
cc_431 N_A2_c_430_n N_A_27_74#_c_1099_n 0.0126582f $X=6.26 $Y=1.22 $X2=0 $Y2=0
cc_432 N_A2_c_432_n N_A_27_74#_c_1099_n 0.0100105f $X=6.76 $Y=1.22 $X2=0 $Y2=0
cc_433 A2 N_A_27_74#_c_1099_n 0.0352336f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_434 N_A2_c_439_n N_A_27_74#_c_1099_n 0.00106692f $X=7.675 $Y=1.385 $X2=0
+ $Y2=0
cc_435 N_A2_c_432_n N_A_27_74#_c_1027_n 2.23968e-19 $X=6.76 $Y=1.22 $X2=0 $Y2=0
cc_436 N_A2_c_434_n N_A_27_74#_c_1027_n 2.23968e-19 $X=7.19 $Y=1.22 $X2=0 $Y2=0
cc_437 N_A2_c_434_n N_A_27_74#_c_1105_n 0.00982315f $X=7.19 $Y=1.22 $X2=0 $Y2=0
cc_438 N_A2_c_436_n N_A_27_74#_c_1105_n 0.0100509f $X=7.655 $Y=1.22 $X2=0 $Y2=0
cc_439 A2 N_A_27_74#_c_1105_n 0.046858f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_440 N_A2_c_439_n N_A_27_74#_c_1105_n 8.48385e-19 $X=7.675 $Y=1.385 $X2=0
+ $Y2=0
cc_441 N_A2_c_436_n N_A_27_74#_c_1028_n 2.6818e-19 $X=7.655 $Y=1.22 $X2=0 $Y2=0
cc_442 N_A2_c_430_n N_A_27_74#_c_1096_n 0.00151008f $X=6.26 $Y=1.22 $X2=0 $Y2=0
cc_443 A2 N_A_27_74#_c_1111_n 0.0146489f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_444 N_A2_c_439_n N_A_27_74#_c_1111_n 7.03576e-19 $X=7.675 $Y=1.385 $X2=0
+ $Y2=0
cc_445 A2 N_A_27_74#_c_1113_n 0.0205097f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_446 N_A2_c_430_n N_VGND_c_1210_n 4.39845e-19 $X=6.26 $Y=1.22 $X2=0 $Y2=0
cc_447 N_A2_c_430_n N_VGND_c_1211_n 0.00335277f $X=6.26 $Y=1.22 $X2=0 $Y2=0
cc_448 N_A2_c_432_n N_VGND_c_1211_n 0.00759025f $X=6.76 $Y=1.22 $X2=0 $Y2=0
cc_449 N_A2_c_434_n N_VGND_c_1211_n 4.20905e-19 $X=7.19 $Y=1.22 $X2=0 $Y2=0
cc_450 N_A2_c_432_n N_VGND_c_1212_n 4.20905e-19 $X=6.76 $Y=1.22 $X2=0 $Y2=0
cc_451 N_A2_c_434_n N_VGND_c_1212_n 0.00749469f $X=7.19 $Y=1.22 $X2=0 $Y2=0
cc_452 N_A2_c_436_n N_VGND_c_1212_n 0.00192221f $X=7.655 $Y=1.22 $X2=0 $Y2=0
cc_453 N_A2_c_436_n N_VGND_c_1213_n 4.08135e-19 $X=7.655 $Y=1.22 $X2=0 $Y2=0
cc_454 N_A2_c_430_n N_VGND_c_1218_n 0.00434272f $X=6.26 $Y=1.22 $X2=0 $Y2=0
cc_455 N_A2_c_432_n N_VGND_c_1219_n 0.00383152f $X=6.76 $Y=1.22 $X2=0 $Y2=0
cc_456 N_A2_c_434_n N_VGND_c_1219_n 0.00383152f $X=7.19 $Y=1.22 $X2=0 $Y2=0
cc_457 N_A2_c_436_n N_VGND_c_1220_n 0.00461464f $X=7.655 $Y=1.22 $X2=0 $Y2=0
cc_458 N_A2_c_430_n N_VGND_c_1223_n 0.00445593f $X=6.26 $Y=1.22 $X2=0 $Y2=0
cc_459 N_A2_c_432_n N_VGND_c_1223_n 0.00383967f $X=6.76 $Y=1.22 $X2=0 $Y2=0
cc_460 N_A2_c_434_n N_VGND_c_1223_n 0.00383967f $X=7.19 $Y=1.22 $X2=0 $Y2=0
cc_461 N_A2_c_436_n N_VGND_c_1223_n 0.00463521f $X=7.655 $Y=1.22 $X2=0 $Y2=0
cc_462 N_A1_M1025_g N_VPWR_c_612_n 0.0163394f $X=8.125 $Y=2.4 $X2=0 $Y2=0
cc_463 N_A1_M1026_g N_VPWR_c_612_n 0.00283364f $X=8.625 $Y=2.4 $X2=0 $Y2=0
cc_464 N_A1_M1035_g N_VPWR_c_613_n 0.00283364f $X=9.075 $Y=2.4 $X2=0 $Y2=0
cc_465 N_A1_M1036_g N_VPWR_c_613_n 0.0195914f $X=9.575 $Y=2.4 $X2=0 $Y2=0
cc_466 N_A1_M1025_g N_VPWR_c_615_n 0.00460063f $X=8.125 $Y=2.4 $X2=0 $Y2=0
cc_467 N_A1_M1026_g N_VPWR_c_616_n 0.00520371f $X=8.625 $Y=2.4 $X2=0 $Y2=0
cc_468 N_A1_M1035_g N_VPWR_c_616_n 0.00520371f $X=9.075 $Y=2.4 $X2=0 $Y2=0
cc_469 N_A1_M1036_g N_VPWR_c_617_n 0.00460063f $X=9.575 $Y=2.4 $X2=0 $Y2=0
cc_470 N_A1_M1025_g N_VPWR_c_608_n 0.00908665f $X=8.125 $Y=2.4 $X2=0 $Y2=0
cc_471 N_A1_M1026_g N_VPWR_c_608_n 0.00981712f $X=8.625 $Y=2.4 $X2=0 $Y2=0
cc_472 N_A1_M1035_g N_VPWR_c_608_n 0.00981712f $X=9.075 $Y=2.4 $X2=0 $Y2=0
cc_473 N_A1_M1036_g N_VPWR_c_608_n 0.00912296f $X=9.575 $Y=2.4 $X2=0 $Y2=0
cc_474 N_A1_M1025_g N_A_1191_368#_c_938_n 0.00100119f $X=8.125 $Y=2.4 $X2=0
+ $Y2=0
cc_475 N_A1_M1025_g N_A_1191_368#_c_939_n 0.0212455f $X=8.125 $Y=2.4 $X2=0 $Y2=0
cc_476 N_A1_M1026_g N_A_1191_368#_c_939_n 0.0132272f $X=8.625 $Y=2.4 $X2=0 $Y2=0
cc_477 N_A1_c_533_n N_A_1191_368#_c_939_n 0.00313888f $X=9.575 $Y=1.55 $X2=0
+ $Y2=0
cc_478 A1 N_A_1191_368#_c_939_n 0.0297341f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_479 N_A1_M1025_g N_A_1191_368#_c_941_n 7.8029e-19 $X=8.125 $Y=2.4 $X2=0 $Y2=0
cc_480 N_A1_M1026_g N_A_1191_368#_c_941_n 0.0158898f $X=8.625 $Y=2.4 $X2=0 $Y2=0
cc_481 N_A1_M1035_g N_A_1191_368#_c_941_n 0.0158898f $X=9.075 $Y=2.4 $X2=0 $Y2=0
cc_482 N_A1_M1036_g N_A_1191_368#_c_941_n 7.8029e-19 $X=9.575 $Y=2.4 $X2=0 $Y2=0
cc_483 N_A1_M1035_g N_A_1191_368#_c_942_n 0.0132272f $X=9.075 $Y=2.4 $X2=0 $Y2=0
cc_484 N_A1_c_533_n N_A_1191_368#_c_942_n 0.00313888f $X=9.575 $Y=1.55 $X2=0
+ $Y2=0
cc_485 N_A1_M1036_g N_A_1191_368#_c_942_n 0.0169522f $X=9.575 $Y=2.4 $X2=0 $Y2=0
cc_486 A1 N_A_1191_368#_c_942_n 0.0736603f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_487 N_A1_M1036_g N_A_1191_368#_c_943_n 0.00282914f $X=9.575 $Y=2.4 $X2=0
+ $Y2=0
cc_488 N_A1_M1026_g N_A_1191_368#_c_945_n 0.00228751f $X=8.625 $Y=2.4 $X2=0
+ $Y2=0
cc_489 N_A1_M1035_g N_A_1191_368#_c_945_n 0.00228751f $X=9.075 $Y=2.4 $X2=0
+ $Y2=0
cc_490 N_A1_c_533_n N_A_1191_368#_c_945_n 0.00215577f $X=9.575 $Y=1.55 $X2=0
+ $Y2=0
cc_491 A1 N_A_1191_368#_c_945_n 0.0277828f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_492 N_A1_c_528_n N_A_27_74#_c_1028_n 2.68041e-19 $X=8.14 $Y=1.22 $X2=0 $Y2=0
cc_493 N_A1_c_528_n N_A_27_74#_c_1115_n 0.0147786f $X=8.14 $Y=1.22 $X2=0 $Y2=0
cc_494 N_A1_c_530_n N_A_27_74#_c_1115_n 0.00899821f $X=8.655 $Y=1.22 $X2=0 $Y2=0
cc_495 N_A1_c_533_n N_A_27_74#_c_1115_n 0.00116455f $X=9.575 $Y=1.55 $X2=0 $Y2=0
cc_496 A1 N_A_27_74#_c_1115_n 0.0301154f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_497 N_A1_c_528_n N_A_27_74#_c_1029_n 4.37256e-19 $X=8.14 $Y=1.22 $X2=0 $Y2=0
cc_498 N_A1_c_530_n N_A_27_74#_c_1029_n 0.0073734f $X=8.655 $Y=1.22 $X2=0 $Y2=0
cc_499 N_A1_c_532_n N_A_27_74#_c_1029_n 0.00723778f $X=9.085 $Y=1.22 $X2=0 $Y2=0
cc_500 N_A1_c_535_n N_A_27_74#_c_1029_n 7.0998e-19 $X=9.585 $Y=1.22 $X2=0 $Y2=0
cc_501 N_A1_c_532_n N_A_27_74#_c_1123_n 0.00892313f $X=9.085 $Y=1.22 $X2=0 $Y2=0
cc_502 N_A1_c_533_n N_A_27_74#_c_1123_n 0.00107107f $X=9.575 $Y=1.55 $X2=0 $Y2=0
cc_503 N_A1_c_535_n N_A_27_74#_c_1123_n 0.0100105f $X=9.585 $Y=1.22 $X2=0 $Y2=0
cc_504 A1 N_A_27_74#_c_1123_n 0.0454799f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_505 A1 N_A_27_74#_c_1030_n 0.0208616f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_506 N_A1_c_535_n N_A_27_74#_c_1031_n 8.26992e-19 $X=9.585 $Y=1.22 $X2=0 $Y2=0
cc_507 N_A1_c_530_n N_A_27_74#_c_1129_n 7.17169e-19 $X=8.655 $Y=1.22 $X2=0 $Y2=0
cc_508 N_A1_c_532_n N_A_27_74#_c_1129_n 7.17169e-19 $X=9.085 $Y=1.22 $X2=0 $Y2=0
cc_509 N_A1_c_533_n N_A_27_74#_c_1129_n 7.03992e-19 $X=9.575 $Y=1.55 $X2=0 $Y2=0
cc_510 A1 N_A_27_74#_c_1129_n 0.0232596f $X=9.755 $Y=1.21 $X2=0 $Y2=0
cc_511 N_A1_c_528_n N_VGND_c_1213_n 0.00685728f $X=8.14 $Y=1.22 $X2=0 $Y2=0
cc_512 N_A1_c_530_n N_VGND_c_1213_n 0.00352333f $X=8.655 $Y=1.22 $X2=0 $Y2=0
cc_513 N_A1_c_532_n N_VGND_c_1214_n 0.00344221f $X=9.085 $Y=1.22 $X2=0 $Y2=0
cc_514 N_A1_c_535_n N_VGND_c_1214_n 0.0105358f $X=9.585 $Y=1.22 $X2=0 $Y2=0
cc_515 N_A1_c_528_n N_VGND_c_1220_n 0.00429299f $X=8.14 $Y=1.22 $X2=0 $Y2=0
cc_516 N_A1_c_530_n N_VGND_c_1221_n 0.00434272f $X=8.655 $Y=1.22 $X2=0 $Y2=0
cc_517 N_A1_c_532_n N_VGND_c_1221_n 0.00434272f $X=9.085 $Y=1.22 $X2=0 $Y2=0
cc_518 N_A1_c_535_n N_VGND_c_1222_n 0.00383152f $X=9.585 $Y=1.22 $X2=0 $Y2=0
cc_519 N_A1_c_528_n N_VGND_c_1223_n 0.00430064f $X=8.14 $Y=1.22 $X2=0 $Y2=0
cc_520 N_A1_c_530_n N_VGND_c_1223_n 0.00445625f $X=8.655 $Y=1.22 $X2=0 $Y2=0
cc_521 N_A1_c_532_n N_VGND_c_1223_n 0.00445496f $X=9.085 $Y=1.22 $X2=0 $Y2=0
cc_522 N_A1_c_535_n N_VGND_c_1223_n 0.00387625f $X=9.585 $Y=1.22 $X2=0 $Y2=0
cc_523 N_VPWR_c_610_n N_Y_c_716_n 0.0416899f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_524 N_VPWR_c_611_n N_Y_c_716_n 0.0353111f $X=1.28 $Y=2.225 $X2=0 $Y2=0
cc_525 N_VPWR_c_614_n N_Y_c_716_n 0.0146357f $X=1.115 $Y=3.33 $X2=0 $Y2=0
cc_526 N_VPWR_c_608_n N_Y_c_716_n 0.0121141f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_527 N_VPWR_M1008_d N_Y_c_717_n 0.00264175f $X=1.145 $Y=1.84 $X2=0 $Y2=0
cc_528 N_VPWR_c_611_n N_Y_c_717_n 0.0219147f $X=1.28 $Y=2.225 $X2=0 $Y2=0
cc_529 N_VPWR_c_610_n N_Y_c_718_n 0.00352479f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_530 N_VPWR_c_611_n N_A_339_368#_c_795_n 0.0565977f $X=1.28 $Y=2.225 $X2=0
+ $Y2=0
cc_531 N_VPWR_c_615_n N_A_339_368#_c_796_n 0.038868f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_532 N_VPWR_c_608_n N_A_339_368#_c_796_n 0.021711f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_533 N_VPWR_c_611_n N_A_339_368#_c_797_n 0.0121616f $X=1.28 $Y=2.225 $X2=0
+ $Y2=0
cc_534 N_VPWR_c_615_n N_A_339_368#_c_797_n 0.0218469f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_535 N_VPWR_c_608_n N_A_339_368#_c_797_n 0.0118348f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_536 N_VPWR_c_615_n N_A_339_368#_c_798_n 0.038868f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_537 N_VPWR_c_608_n N_A_339_368#_c_798_n 0.021711f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_538 N_VPWR_c_615_n N_A_339_368#_c_800_n 0.0422345f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_539 N_VPWR_c_608_n N_A_339_368#_c_800_n 0.0238184f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_540 N_VPWR_c_615_n N_A_339_368#_c_801_n 0.0593439f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_541 N_VPWR_c_608_n N_A_339_368#_c_801_n 0.032751f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_542 N_VPWR_c_615_n N_A_339_368#_c_803_n 0.0200371f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_543 N_VPWR_c_608_n N_A_339_368#_c_803_n 0.01084f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_544 N_VPWR_c_615_n N_A_339_368#_c_804_n 0.0217415f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_545 N_VPWR_c_608_n N_A_339_368#_c_804_n 0.0116975f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_546 N_VPWR_c_615_n N_A_339_368#_c_805_n 0.0234458f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_547 N_VPWR_c_608_n N_A_339_368#_c_805_n 0.0125551f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_548 N_VPWR_c_615_n N_A_1191_368#_c_936_n 0.0359969f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_549 N_VPWR_c_608_n N_A_1191_368#_c_936_n 0.0200963f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_550 N_VPWR_c_615_n N_A_1191_368#_c_937_n 0.0235512f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_551 N_VPWR_c_608_n N_A_1191_368#_c_937_n 0.0126924f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_552 N_VPWR_c_612_n N_A_1191_368#_c_938_n 0.0117236f $X=8.35 $Y=2.225 $X2=0
+ $Y2=0
cc_553 N_VPWR_c_615_n N_A_1191_368#_c_938_n 0.0557595f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_554 N_VPWR_c_608_n N_A_1191_368#_c_938_n 0.0308071f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_555 N_VPWR_M1025_d N_A_1191_368#_c_939_n 0.00218982f $X=8.215 $Y=1.84 $X2=0
+ $Y2=0
cc_556 N_VPWR_c_612_n N_A_1191_368#_c_939_n 0.0189268f $X=8.35 $Y=2.225 $X2=0
+ $Y2=0
cc_557 N_VPWR_c_612_n N_A_1191_368#_c_941_n 0.0368936f $X=8.35 $Y=2.225 $X2=0
+ $Y2=0
cc_558 N_VPWR_c_613_n N_A_1191_368#_c_941_n 0.0368936f $X=9.35 $Y=2.225 $X2=0
+ $Y2=0
cc_559 N_VPWR_c_616_n N_A_1191_368#_c_941_n 0.0157306f $X=9.185 $Y=3.33 $X2=0
+ $Y2=0
cc_560 N_VPWR_c_608_n N_A_1191_368#_c_941_n 0.0119807f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_561 N_VPWR_M1035_d N_A_1191_368#_c_942_n 0.00218982f $X=9.165 $Y=1.84 $X2=0
+ $Y2=0
cc_562 N_VPWR_c_613_n N_A_1191_368#_c_942_n 0.0189268f $X=9.35 $Y=2.225 $X2=0
+ $Y2=0
cc_563 N_VPWR_c_613_n N_A_1191_368#_c_943_n 0.0368537f $X=9.35 $Y=2.225 $X2=0
+ $Y2=0
cc_564 N_VPWR_c_617_n N_A_1191_368#_c_943_n 0.0134846f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_565 N_VPWR_c_608_n N_A_1191_368#_c_943_n 0.0103893f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_566 N_VPWR_c_615_n N_A_1191_368#_c_944_n 0.0234458f $X=8.185 $Y=3.33 $X2=0
+ $Y2=0
cc_567 N_VPWR_c_608_n N_A_1191_368#_c_944_n 0.0125551f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_568 N_Y_c_720_n N_A_339_368#_M1015_s 0.00119058f $X=2.15 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_569 N_Y_c_721_n N_A_339_368#_M1015_s 0.00149404f $X=1.64 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_570 N_Y_c_759_n N_A_339_368#_M1018_s 0.00170631f $X=3.05 $Y=1.935 $X2=0 $Y2=0
cc_571 N_Y_c_720_n N_A_339_368#_c_795_n 0.00941962f $X=2.15 $Y=1.805 $X2=0 $Y2=0
cc_572 N_Y_c_721_n N_A_339_368#_c_795_n 0.011698f $X=1.64 $Y=1.805 $X2=0 $Y2=0
cc_573 N_Y_c_749_n N_A_339_368#_c_795_n 0.0501993f $X=2.29 $Y=1.965 $X2=0 $Y2=0
cc_574 N_Y_M1015_d N_A_339_368#_c_796_n 0.00165831f $X=2.155 $Y=1.84 $X2=0 $Y2=0
cc_575 N_Y_c_749_n N_A_339_368#_c_796_n 0.0123692f $X=2.29 $Y=1.965 $X2=0 $Y2=0
cc_576 N_Y_c_749_n N_A_339_368#_c_813_n 0.0303695f $X=2.29 $Y=1.965 $X2=0 $Y2=0
cc_577 Y N_A_339_368#_c_813_n 0.0303695f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_578 N_Y_c_759_n N_A_339_368#_c_813_n 0.0141053f $X=3.05 $Y=1.935 $X2=0 $Y2=0
cc_579 N_Y_M1020_d N_A_339_368#_c_798_n 0.00165831f $X=3.055 $Y=1.84 $X2=0 $Y2=0
cc_580 Y N_A_339_368#_c_798_n 0.0123692f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_581 Y N_A_339_368#_c_799_n 0.0708362f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_582 Y N_A_791_368#_c_889_n 0.0025132f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_583 N_Y_c_724_n N_A_27_74#_M1010_d 0.00433624f $X=1.475 $Y=0.925 $X2=0 $Y2=0
cc_584 N_Y_M1009_s N_A_27_74#_c_1017_n 0.00176461f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_585 N_Y_c_724_n N_A_27_74#_c_1017_n 0.0035136f $X=1.475 $Y=0.925 $X2=0 $Y2=0
cc_586 N_Y_c_741_n N_A_27_74#_c_1017_n 0.0121701f $X=0.71 $Y=0.8 $X2=0 $Y2=0
cc_587 N_Y_M1029_s N_A_27_74#_c_1019_n 0.00250873f $X=1.43 $Y=0.37 $X2=0 $Y2=0
cc_588 N_Y_c_724_n N_A_27_74#_c_1019_n 0.00352531f $X=1.475 $Y=0.925 $X2=0 $Y2=0
cc_589 N_Y_c_734_n N_A_27_74#_c_1019_n 0.019744f $X=1.64 $Y=1.01 $X2=0 $Y2=0
cc_590 N_Y_c_724_n N_A_27_74#_c_1032_n 0.0160355f $X=1.475 $Y=0.925 $X2=0 $Y2=0
cc_591 N_Y_c_724_n N_VGND_c_1223_n 0.00143802f $X=1.475 $Y=0.925 $X2=0 $Y2=0
cc_592 N_A_339_368#_c_800_n N_A_791_368#_M1003_s 0.00275122f $X=4.475 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_593 N_A_339_368#_c_801_n N_A_791_368#_M1024_s 0.00165831f $X=5.375 $Y=2.99
+ $X2=0 $Y2=0
cc_594 N_A_339_368#_c_800_n N_A_791_368#_c_918_n 0.0194849f $X=4.475 $Y=2.99
+ $X2=0 $Y2=0
cc_595 N_A_339_368#_M1021_d N_A_791_368#_c_893_n 0.00165831f $X=4.505 $Y=1.84
+ $X2=0 $Y2=0
cc_596 N_A_339_368#_c_830_n N_A_791_368#_c_893_n 0.0170258f $X=4.64 $Y=2.145
+ $X2=0 $Y2=0
cc_597 N_A_339_368#_c_799_n N_A_791_368#_c_889_n 0.00517049f $X=3.64 $Y=1.965
+ $X2=0 $Y2=0
cc_598 N_A_339_368#_c_801_n N_A_791_368#_c_922_n 0.0118736f $X=5.375 $Y=2.99
+ $X2=0 $Y2=0
cc_599 N_A_339_368#_M1028_d N_A_791_368#_c_890_n 0.00264175f $X=5.405 $Y=1.84
+ $X2=0 $Y2=0
cc_600 N_A_339_368#_c_802_n N_A_791_368#_c_890_n 0.0219146f $X=5.54 $Y=2.145
+ $X2=0 $Y2=0
cc_601 N_A_339_368#_c_802_n N_A_1191_368#_c_935_n 0.0559235f $X=5.54 $Y=2.145
+ $X2=0 $Y2=0
cc_602 N_A_339_368#_c_801_n N_A_1191_368#_c_937_n 0.0128664f $X=5.375 $Y=2.99
+ $X2=0 $Y2=0
cc_603 N_A_339_368#_c_802_n N_A_1191_368#_c_937_n 0.00103927f $X=5.54 $Y=2.145
+ $X2=0 $Y2=0
cc_604 N_A_339_368#_c_799_n N_A_27_74#_c_1022_n 0.0159621f $X=3.64 $Y=1.965
+ $X2=0 $Y2=0
cc_605 N_A_791_368#_c_890_n N_A_1191_368#_M1013_s 0.00264175f $X=6.435 $Y=1.805
+ $X2=-0.19 $Y2=1.66
cc_606 N_A_791_368#_c_891_n N_A_1191_368#_M1016_s 0.00165831f $X=7.335 $Y=1.805
+ $X2=0 $Y2=0
cc_607 N_A_791_368#_c_890_n N_A_1191_368#_c_935_n 0.0219147f $X=6.435 $Y=1.805
+ $X2=0 $Y2=0
cc_608 N_A_791_368#_M1013_d N_A_1191_368#_c_936_n 0.00166264f $X=6.415 $Y=1.84
+ $X2=0 $Y2=0
cc_609 N_A_791_368#_c_929_p N_A_1191_368#_c_936_n 0.0119845f $X=6.55 $Y=1.965
+ $X2=0 $Y2=0
cc_610 N_A_791_368#_c_891_n N_A_1191_368#_c_953_n 0.0170259f $X=7.335 $Y=1.805
+ $X2=0 $Y2=0
cc_611 N_A_791_368#_M1019_d N_A_1191_368#_c_938_n 0.00165831f $X=7.315 $Y=1.84
+ $X2=0 $Y2=0
cc_612 N_A_791_368#_c_932_p N_A_1191_368#_c_938_n 0.0118736f $X=7.45 $Y=2.045
+ $X2=0 $Y2=0
cc_613 N_A_791_368#_c_891_n N_A_1191_368#_c_940_n 0.0127663f $X=7.335 $Y=1.805
+ $X2=0 $Y2=0
cc_614 N_A_791_368#_c_889_n N_A_27_74#_c_1022_n 0.0139914f $X=4.305 $Y=1.805
+ $X2=0 $Y2=0
cc_615 N_A_27_74#_c_1048_n N_VGND_M1000_d 0.0117286f $X=3.16 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_616 N_A_27_74#_c_1079_n N_VGND_M1001_d 0.00462121f $X=5.03 $Y=0.925 $X2=0
+ $Y2=0
cc_617 N_A_27_74#_c_1086_n N_VGND_M1034_d 0.00462121f $X=5.96 $Y=0.925 $X2=0
+ $Y2=0
cc_618 N_A_27_74#_c_1099_n N_VGND_M1002_s 0.00462121f $X=6.89 $Y=0.925 $X2=0
+ $Y2=0
cc_619 N_A_27_74#_c_1105_n N_VGND_M1014_s 0.00395707f $X=7.785 $Y=0.925 $X2=0
+ $Y2=0
cc_620 N_A_27_74#_c_1115_n N_VGND_M1005_s 0.00530982f $X=8.705 $Y=0.925 $X2=0
+ $Y2=0
cc_621 N_A_27_74#_c_1123_n N_VGND_M1032_s 0.00462121f $X=9.715 $Y=0.925 $X2=0
+ $Y2=0
cc_622 N_A_27_74#_c_1020_n N_VGND_c_1206_n 0.0191473f $X=3.325 $Y=0.515 $X2=0
+ $Y2=0
cc_623 N_A_27_74#_c_1021_n N_VGND_c_1206_n 0.00474779f $X=3.415 $Y=1.3 $X2=0
+ $Y2=0
cc_624 N_A_27_74#_c_1022_n N_VGND_c_1206_n 0.013555f $X=4.02 $Y=1.385 $X2=0
+ $Y2=0
cc_625 N_A_27_74#_c_1023_n N_VGND_c_1206_n 0.018213f $X=4.185 $Y=0.515 $X2=0
+ $Y2=0
cc_626 N_A_27_74#_c_1024_n N_VGND_c_1206_n 0.00453882f $X=4.105 $Y=1.3 $X2=0
+ $Y2=0
cc_627 N_A_27_74#_c_1023_n N_VGND_c_1207_n 0.014477f $X=4.185 $Y=0.515 $X2=0
+ $Y2=0
cc_628 N_A_27_74#_c_1023_n N_VGND_c_1208_n 0.0127977f $X=4.185 $Y=0.515 $X2=0
+ $Y2=0
cc_629 N_A_27_74#_c_1079_n N_VGND_c_1208_n 0.0205261f $X=5.03 $Y=0.925 $X2=0
+ $Y2=0
cc_630 N_A_27_74#_c_1025_n N_VGND_c_1208_n 0.0121972f $X=5.115 $Y=0.515 $X2=0
+ $Y2=0
cc_631 N_A_27_74#_c_1025_n N_VGND_c_1209_n 0.0109704f $X=5.115 $Y=0.515 $X2=0
+ $Y2=0
cc_632 N_A_27_74#_c_1025_n N_VGND_c_1210_n 0.0122975f $X=5.115 $Y=0.515 $X2=0
+ $Y2=0
cc_633 N_A_27_74#_c_1086_n N_VGND_c_1210_n 0.0205261f $X=5.96 $Y=0.925 $X2=0
+ $Y2=0
cc_634 N_A_27_74#_c_1026_n N_VGND_c_1210_n 0.0121972f $X=6.045 $Y=0.515 $X2=0
+ $Y2=0
cc_635 N_A_27_74#_c_1026_n N_VGND_c_1211_n 0.0122975f $X=6.045 $Y=0.515 $X2=0
+ $Y2=0
cc_636 N_A_27_74#_c_1099_n N_VGND_c_1211_n 0.0205261f $X=6.89 $Y=0.925 $X2=0
+ $Y2=0
cc_637 N_A_27_74#_c_1027_n N_VGND_c_1211_n 0.0121558f $X=6.975 $Y=0.515 $X2=0
+ $Y2=0
cc_638 N_A_27_74#_c_1027_n N_VGND_c_1212_n 0.0121558f $X=6.975 $Y=0.515 $X2=0
+ $Y2=0
cc_639 N_A_27_74#_c_1105_n N_VGND_c_1212_n 0.0177409f $X=7.785 $Y=0.925 $X2=0
+ $Y2=0
cc_640 N_A_27_74#_c_1028_n N_VGND_c_1212_n 0.00131301f $X=7.87 $Y=0.515 $X2=0
+ $Y2=0
cc_641 N_A_27_74#_c_1028_n N_VGND_c_1213_n 0.0127651f $X=7.87 $Y=0.515 $X2=0
+ $Y2=0
cc_642 N_A_27_74#_c_1115_n N_VGND_c_1213_n 0.020602f $X=8.705 $Y=0.925 $X2=0
+ $Y2=0
cc_643 N_A_27_74#_c_1029_n N_VGND_c_1213_n 0.0127977f $X=8.87 $Y=0.515 $X2=0
+ $Y2=0
cc_644 N_A_27_74#_c_1029_n N_VGND_c_1214_n 0.0127977f $X=8.87 $Y=0.515 $X2=0
+ $Y2=0
cc_645 N_A_27_74#_c_1123_n N_VGND_c_1214_n 0.0205261f $X=9.715 $Y=0.925 $X2=0
+ $Y2=0
cc_646 N_A_27_74#_c_1031_n N_VGND_c_1214_n 0.0121972f $X=9.8 $Y=0.515 $X2=0
+ $Y2=0
cc_647 N_A_27_74#_c_1020_n N_VGND_c_1215_n 0.0149638f $X=3.325 $Y=0.515 $X2=0
+ $Y2=0
cc_648 N_A_27_74#_c_1017_n N_VGND_c_1217_n 0.0333877f $X=0.975 $Y=0.34 $X2=0
+ $Y2=0
cc_649 N_A_27_74#_c_1018_n N_VGND_c_1217_n 0.0235688f $X=0.445 $Y=0.34 $X2=0
+ $Y2=0
cc_650 N_A_27_74#_c_1019_n N_VGND_c_1217_n 0.0781546f $X=1.975 $Y=0.34 $X2=0
+ $Y2=0
cc_651 N_A_27_74#_c_1048_n N_VGND_c_1217_n 0.0278307f $X=3.16 $Y=0.925 $X2=0
+ $Y2=0
cc_652 N_A_27_74#_c_1020_n N_VGND_c_1217_n 0.0112517f $X=3.325 $Y=0.515 $X2=0
+ $Y2=0
cc_653 N_A_27_74#_c_1032_n N_VGND_c_1217_n 0.0225055f $X=1.14 $Y=0.34 $X2=0
+ $Y2=0
cc_654 N_A_27_74#_c_1026_n N_VGND_c_1218_n 0.0109704f $X=6.045 $Y=0.515 $X2=0
+ $Y2=0
cc_655 N_A_27_74#_c_1027_n N_VGND_c_1219_n 0.00747999f $X=6.975 $Y=0.515 $X2=0
+ $Y2=0
cc_656 N_A_27_74#_c_1028_n N_VGND_c_1220_n 0.0110419f $X=7.87 $Y=0.515 $X2=0
+ $Y2=0
cc_657 N_A_27_74#_c_1029_n N_VGND_c_1221_n 0.0144609f $X=8.87 $Y=0.515 $X2=0
+ $Y2=0
cc_658 N_A_27_74#_c_1031_n N_VGND_c_1222_n 0.0110419f $X=9.8 $Y=0.515 $X2=0
+ $Y2=0
cc_659 N_A_27_74#_c_1017_n N_VGND_c_1223_n 0.0187857f $X=0.975 $Y=0.34 $X2=0
+ $Y2=0
cc_660 N_A_27_74#_c_1018_n N_VGND_c_1223_n 0.0127152f $X=0.445 $Y=0.34 $X2=0
+ $Y2=0
cc_661 N_A_27_74#_c_1019_n N_VGND_c_1223_n 0.0366503f $X=1.975 $Y=0.34 $X2=0
+ $Y2=0
cc_662 N_A_27_74#_c_1048_n N_VGND_c_1223_n 0.0117436f $X=3.16 $Y=0.925 $X2=0
+ $Y2=0
cc_663 N_A_27_74#_c_1020_n N_VGND_c_1223_n 0.0123131f $X=3.325 $Y=0.515 $X2=0
+ $Y2=0
cc_664 N_A_27_74#_c_1023_n N_VGND_c_1223_n 0.0118767f $X=4.185 $Y=0.515 $X2=0
+ $Y2=0
cc_665 N_A_27_74#_c_1079_n N_VGND_c_1223_n 0.0113542f $X=5.03 $Y=0.925 $X2=0
+ $Y2=0
cc_666 N_A_27_74#_c_1025_n N_VGND_c_1223_n 0.00903439f $X=5.115 $Y=0.515 $X2=0
+ $Y2=0
cc_667 N_A_27_74#_c_1086_n N_VGND_c_1223_n 0.0113542f $X=5.96 $Y=0.925 $X2=0
+ $Y2=0
cc_668 N_A_27_74#_c_1026_n N_VGND_c_1223_n 0.00903439f $X=6.045 $Y=0.515 $X2=0
+ $Y2=0
cc_669 N_A_27_74#_c_1099_n N_VGND_c_1223_n 0.0113542f $X=6.89 $Y=0.925 $X2=0
+ $Y2=0
cc_670 N_A_27_74#_c_1027_n N_VGND_c_1223_n 0.00619848f $X=6.975 $Y=0.515 $X2=0
+ $Y2=0
cc_671 N_A_27_74#_c_1105_n N_VGND_c_1223_n 0.0126991f $X=7.785 $Y=0.925 $X2=0
+ $Y2=0
cc_672 N_A_27_74#_c_1028_n N_VGND_c_1223_n 0.00915013f $X=7.87 $Y=0.515 $X2=0
+ $Y2=0
cc_673 N_A_27_74#_c_1115_n N_VGND_c_1223_n 0.0109057f $X=8.705 $Y=0.925 $X2=0
+ $Y2=0
cc_674 N_A_27_74#_c_1029_n N_VGND_c_1223_n 0.0118703f $X=8.87 $Y=0.515 $X2=0
+ $Y2=0
cc_675 N_A_27_74#_c_1123_n N_VGND_c_1223_n 0.0113542f $X=9.715 $Y=0.925 $X2=0
+ $Y2=0
cc_676 N_A_27_74#_c_1031_n N_VGND_c_1223_n 0.00915013f $X=9.8 $Y=0.515 $X2=0
+ $Y2=0
cc_677 N_A_27_74#_c_1032_n N_VGND_c_1223_n 0.0123739f $X=1.14 $Y=0.34 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__a41oi_2.pxi.spice
* Created: Wed Sep  2 11:56:45 2020
* 
x_PM_SKY130_FD_SC_MS__A41OI_2%B1 N_B1_M1007_g N_B1_M1013_g N_B1_M1009_g B1 B1
+ N_B1_c_91_n N_B1_c_92_n PM_SKY130_FD_SC_MS__A41OI_2%B1
x_PM_SKY130_FD_SC_MS__A41OI_2%A1 N_A1_c_133_n N_A1_M1002_g N_A1_M1011_g
+ N_A1_M1018_g N_A1_c_134_n N_A1_M1006_g A1 N_A1_c_135_n N_A1_c_132_n
+ PM_SKY130_FD_SC_MS__A41OI_2%A1
x_PM_SKY130_FD_SC_MS__A41OI_2%A2 N_A2_c_195_n N_A2_M1010_g N_A2_M1001_g
+ N_A2_c_197_n N_A2_M1016_g N_A2_M1005_g A2 A2 N_A2_c_200_n
+ PM_SKY130_FD_SC_MS__A41OI_2%A2
x_PM_SKY130_FD_SC_MS__A41OI_2%A3 N_A3_M1000_g N_A3_M1004_g N_A3_M1003_g
+ N_A3_M1017_g A3 A3 N_A3_c_267_n PM_SKY130_FD_SC_MS__A41OI_2%A3
x_PM_SKY130_FD_SC_MS__A41OI_2%A4 N_A4_M1014_g N_A4_M1008_g N_A4_M1012_g
+ N_A4_M1015_g A4 A4 N_A4_c_324_n PM_SKY130_FD_SC_MS__A41OI_2%A4
x_PM_SKY130_FD_SC_MS__A41OI_2%A_27_368# N_A_27_368#_M1007_d N_A_27_368#_M1009_d
+ N_A_27_368#_M1006_d N_A_27_368#_M1005_d N_A_27_368#_M1003_d
+ N_A_27_368#_M1012_s N_A_27_368#_c_361_n N_A_27_368#_c_362_n
+ N_A_27_368#_c_363_n N_A_27_368#_c_377_n N_A_27_368#_c_378_n
+ N_A_27_368#_c_379_n N_A_27_368#_c_364_n N_A_27_368#_c_383_n
+ N_A_27_368#_c_365_n N_A_27_368#_c_392_n N_A_27_368#_c_366_n
+ N_A_27_368#_c_399_n N_A_27_368#_c_367_n N_A_27_368#_c_416_n
+ N_A_27_368#_c_368_n N_A_27_368#_c_369_n N_A_27_368#_c_385_n
+ N_A_27_368#_c_401_n N_A_27_368#_c_412_n PM_SKY130_FD_SC_MS__A41OI_2%A_27_368#
x_PM_SKY130_FD_SC_MS__A41OI_2%Y N_Y_M1013_d N_Y_M1011_d N_Y_M1007_s N_Y_c_457_n
+ N_Y_c_458_n N_Y_c_459_n N_Y_c_470_n N_Y_c_482_n N_Y_c_463_n N_Y_c_472_n
+ N_Y_c_460_n Y N_Y_c_461_n Y PM_SKY130_FD_SC_MS__A41OI_2%Y
x_PM_SKY130_FD_SC_MS__A41OI_2%VPWR N_VPWR_M1002_s N_VPWR_M1001_s N_VPWR_M1000_s
+ N_VPWR_M1008_d N_VPWR_c_525_n N_VPWR_c_526_n N_VPWR_c_527_n N_VPWR_c_528_n
+ N_VPWR_c_529_n N_VPWR_c_530_n N_VPWR_c_531_n N_VPWR_c_532_n VPWR
+ N_VPWR_c_533_n N_VPWR_c_534_n N_VPWR_c_535_n N_VPWR_c_524_n N_VPWR_c_537_n
+ N_VPWR_c_538_n PM_SKY130_FD_SC_MS__A41OI_2%VPWR
x_PM_SKY130_FD_SC_MS__A41OI_2%VGND N_VGND_M1013_s N_VGND_M1014_s N_VGND_c_598_n
+ N_VGND_c_599_n N_VGND_c_600_n VGND N_VGND_c_601_n N_VGND_c_602_n
+ N_VGND_c_603_n N_VGND_c_604_n PM_SKY130_FD_SC_MS__A41OI_2%VGND
x_PM_SKY130_FD_SC_MS__A41OI_2%A_239_74# N_A_239_74#_M1011_s N_A_239_74#_M1018_s
+ N_A_239_74#_M1016_d N_A_239_74#_c_651_n N_A_239_74#_c_652_n
+ N_A_239_74#_c_653_n N_A_239_74#_c_662_n N_A_239_74#_c_664_n
+ N_A_239_74#_c_654_n PM_SKY130_FD_SC_MS__A41OI_2%A_239_74#
x_PM_SKY130_FD_SC_MS__A41OI_2%A_512_74# N_A_512_74#_M1010_s N_A_512_74#_M1004_s
+ N_A_512_74#_c_695_n N_A_512_74#_c_696_n PM_SKY130_FD_SC_MS__A41OI_2%A_512_74#
x_PM_SKY130_FD_SC_MS__A41OI_2%A_709_74# N_A_709_74#_M1004_d N_A_709_74#_M1017_d
+ N_A_709_74#_M1015_d N_A_709_74#_c_716_n N_A_709_74#_c_717_n
+ N_A_709_74#_c_718_n N_A_709_74#_c_719_n N_A_709_74#_c_720_n
+ PM_SKY130_FD_SC_MS__A41OI_2%A_709_74#
cc_1 VNB N_B1_M1013_g 0.0324508f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.79
cc_2 VNB N_B1_c_91_n 0.0165437f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.515
cc_3 VNB N_B1_c_92_n 0.0527642f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.515
cc_4 VNB N_A1_M1011_g 0.0303832f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.79
cc_5 VNB N_A1_M1018_g 0.0222307f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_6 VNB N_A1_c_132_n 0.0490906f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.515
cc_7 VNB N_A2_c_195_n 0.0160246f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.68
cc_8 VNB N_A2_M1001_g 0.00169644f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.79
cc_9 VNB N_A2_c_197_n 0.0201419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A2_M1005_g 0.00141159f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_11 VNB A2 0.0100854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_c_200_n 0.0803198f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_13 VNB N_A3_M1000_g 0.00792799f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_14 VNB N_A3_M1004_g 0.0298132f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.79
cc_15 VNB N_A3_M1017_g 0.0239845f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB A3 0.00664811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A3_c_267_n 0.044085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A4_M1014_g 0.0237305f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_19 VNB N_A4_M1015_g 0.0333521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB A4 0.0171287f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A4_c_324_n 0.0393506f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_22 VNB N_Y_c_457_n 0.00935246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_458_n 0.022726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_459_n 0.00203445f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.515
cc_25 VNB N_Y_c_460_n 7.09812e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_461_n 0.007391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB Y 0.00225532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_524_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_598_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.79
cc_30 VNB N_VGND_c_599_n 0.0498697f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.68
cc_31 VNB N_VGND_c_600_n 0.00641104f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_32 VNB N_VGND_c_601_n 0.108993f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.515
cc_33 VNB N_VGND_c_602_n 0.0191315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_603_n 0.331124f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_35 VNB N_VGND_c_604_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_239_74#_c_651_n 0.00384069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_239_74#_c_652_n 0.00566166f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_38 VNB N_A_239_74#_c_653_n 0.00613558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_239_74#_c_654_n 0.00383032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_512_74#_c_695_n 0.0022973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_512_74#_c_696_n 0.0197244f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_42 VNB N_A_709_74#_c_716_n 0.00883436f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_43 VNB N_A_709_74#_c_717_n 0.00178889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_709_74#_c_718_n 0.0163059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_709_74#_c_719_n 0.0278949f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.515
cc_46 VNB N_A_709_74#_c_720_n 0.00213459f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_47 VPB N_B1_M1007_g 0.0258571f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_48 VPB N_B1_M1009_g 0.0214873f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_49 VPB N_B1_c_91_n 0.0115973f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.515
cc_50 VPB N_B1_c_92_n 0.00644459f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.515
cc_51 VPB N_A1_c_133_n 0.0212143f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.68
cc_52 VPB N_A1_c_134_n 0.0213575f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A1_c_135_n 0.00221857f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.515
cc_54 VPB N_A1_c_132_n 0.0195426f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.515
cc_55 VPB N_A2_M1001_g 0.0239547f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.79
cc_56 VPB N_A2_M1005_g 0.022916f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_57 VPB A2 0.00533426f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A3_M1000_g 0.0233287f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_59 VPB N_A3_M1003_g 0.0226891f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_60 VPB A3 0.00691685f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A3_c_267_n 0.00552972f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A4_M1008_g 0.0220427f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.79
cc_63 VPB N_A4_M1012_g 0.0262488f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_64 VPB A4 0.0110721f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A4_c_324_n 0.00487321f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_66 VPB N_A_27_368#_c_361_n 0.0366851f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.515
cc_67 VPB N_A_27_368#_c_362_n 0.00459762f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_68 VPB N_A_27_368#_c_363_n 0.00965867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_27_368#_c_364_n 0.0059777f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_27_368#_c_365_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_27_368#_c_366_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_27_368#_c_367_n 0.00321179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_27_368#_c_368_n 0.0075506f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_27_368#_c_369_n 0.0362086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_Y_c_463_n 0.00201719f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_76 VPB N_VPWR_c_525_n 0.0105945f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_526_n 0.0083004f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=1.515
cc_78 VPB N_VPWR_c_527_n 0.00891313f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.515
cc_79 VPB N_VPWR_c_528_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_529_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.565
cc_81 VPB N_VPWR_c_530_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_531_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_532_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_533_n 0.0405994f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_534_n 0.0192638f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_535_n 0.0182986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_524_n 0.067976f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_537_n 0.00997248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_538_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 N_B1_M1009_g N_A1_c_133_n 0.0206339f $X=1.005 $Y=2.4 $X2=-0.19 $Y2=-0.245
cc_91 N_B1_c_91_n N_A1_c_135_n 0.0164601f $X=0.92 $Y=1.515 $X2=0 $Y2=0
cc_92 N_B1_c_92_n N_A1_c_135_n 0.00152595f $X=1.005 $Y=1.515 $X2=0 $Y2=0
cc_93 N_B1_c_91_n N_A1_c_132_n 0.00209039f $X=0.92 $Y=1.515 $X2=0 $Y2=0
cc_94 N_B1_c_92_n N_A1_c_132_n 0.0206339f $X=1.005 $Y=1.515 $X2=0 $Y2=0
cc_95 N_B1_M1007_g N_A_27_368#_c_361_n 0.0128753f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_96 N_B1_M1009_g N_A_27_368#_c_361_n 5.96058e-19 $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_97 N_B1_c_91_n N_A_27_368#_c_361_n 0.0254127f $X=0.92 $Y=1.515 $X2=0 $Y2=0
cc_98 N_B1_M1007_g N_A_27_368#_c_362_n 0.0119307f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_99 N_B1_M1009_g N_A_27_368#_c_362_n 0.0144846f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_100 N_B1_M1007_g N_A_27_368#_c_363_n 0.00291744f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_101 N_B1_M1013_g N_Y_c_457_n 0.00835524f $X=0.565 $Y=0.79 $X2=0 $Y2=0
cc_102 N_B1_c_91_n N_Y_c_458_n 0.0107014f $X=0.92 $Y=1.515 $X2=0 $Y2=0
cc_103 N_B1_c_92_n N_Y_c_458_n 0.00410333f $X=1.005 $Y=1.515 $X2=0 $Y2=0
cc_104 N_B1_M1013_g N_Y_c_459_n 0.00264023f $X=0.565 $Y=0.79 $X2=0 $Y2=0
cc_105 N_B1_c_91_n N_Y_c_459_n 0.0282314f $X=0.92 $Y=1.515 $X2=0 $Y2=0
cc_106 N_B1_c_92_n N_Y_c_459_n 0.00775596f $X=1.005 $Y=1.515 $X2=0 $Y2=0
cc_107 N_B1_M1009_g N_Y_c_470_n 0.013466f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_108 N_B1_c_91_n N_Y_c_470_n 0.010181f $X=0.92 $Y=1.515 $X2=0 $Y2=0
cc_109 N_B1_M1009_g N_Y_c_472_n 0.0108419f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_110 N_B1_c_91_n N_Y_c_472_n 0.0246996f $X=0.92 $Y=1.515 $X2=0 $Y2=0
cc_111 N_B1_c_92_n N_Y_c_472_n 8.62986e-19 $X=1.005 $Y=1.515 $X2=0 $Y2=0
cc_112 N_B1_M1007_g N_VPWR_c_533_n 0.00333896f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_113 N_B1_M1009_g N_VPWR_c_533_n 0.00333926f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_114 N_B1_M1007_g N_VPWR_c_524_n 0.00426915f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_115 N_B1_M1009_g N_VPWR_c_524_n 0.00423742f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_116 N_B1_M1013_g N_VGND_c_599_n 0.0199087f $X=0.565 $Y=0.79 $X2=0 $Y2=0
cc_117 N_B1_c_91_n N_VGND_c_599_n 0.0286397f $X=0.92 $Y=1.515 $X2=0 $Y2=0
cc_118 N_B1_c_92_n N_VGND_c_599_n 7.89955e-19 $X=1.005 $Y=1.515 $X2=0 $Y2=0
cc_119 N_B1_M1013_g N_VGND_c_601_n 0.00517302f $X=0.565 $Y=0.79 $X2=0 $Y2=0
cc_120 N_B1_M1013_g N_VGND_c_603_n 0.00529924f $X=0.565 $Y=0.79 $X2=0 $Y2=0
cc_121 N_B1_M1013_g N_A_239_74#_c_651_n 8.49936e-19 $X=0.565 $Y=0.79 $X2=0 $Y2=0
cc_122 N_B1_M1013_g N_A_239_74#_c_653_n 0.00318346f $X=0.565 $Y=0.79 $X2=0 $Y2=0
cc_123 N_A1_M1018_g N_A2_c_195_n 0.0233638f $X=1.985 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_124 N_A1_c_134_n N_A2_M1001_g 0.0107448f $X=2.245 $Y=1.725 $X2=0 $Y2=0
cc_125 N_A1_M1018_g A2 2.3232e-19 $X=1.985 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A1_c_132_n A2 2.24269e-19 $X=1.985 $Y=1.537 $X2=0 $Y2=0
cc_127 N_A1_M1018_g N_A2_c_200_n 0.00420591f $X=1.985 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A1_c_132_n N_A2_c_200_n 0.0107448f $X=1.985 $Y=1.537 $X2=0 $Y2=0
cc_129 N_A1_c_133_n N_A_27_368#_c_362_n 0.00364476f $X=1.505 $Y=1.725 $X2=0
+ $Y2=0
cc_130 N_A1_c_133_n N_A_27_368#_c_377_n 8.84614e-19 $X=1.505 $Y=1.725 $X2=0
+ $Y2=0
cc_131 N_A1_c_133_n N_A_27_368#_c_378_n 0.0114943f $X=1.505 $Y=1.725 $X2=0 $Y2=0
cc_132 N_A1_c_133_n N_A_27_368#_c_379_n 0.0139713f $X=1.505 $Y=1.725 $X2=0 $Y2=0
cc_133 N_A1_c_134_n N_A_27_368#_c_379_n 0.0166137f $X=2.245 $Y=1.725 $X2=0 $Y2=0
cc_134 N_A1_c_132_n N_A_27_368#_c_379_n 5.03511e-19 $X=1.985 $Y=1.537 $X2=0
+ $Y2=0
cc_135 N_A1_c_134_n N_A_27_368#_c_364_n 0.00513936f $X=2.245 $Y=1.725 $X2=0
+ $Y2=0
cc_136 N_A1_c_134_n N_A_27_368#_c_383_n 0.0076999f $X=2.245 $Y=1.725 $X2=0 $Y2=0
cc_137 N_A1_c_134_n N_A_27_368#_c_365_n 0.013005f $X=2.245 $Y=1.725 $X2=0 $Y2=0
cc_138 N_A1_c_134_n N_A_27_368#_c_385_n 4.64231e-19 $X=2.245 $Y=1.725 $X2=0
+ $Y2=0
cc_139 N_A1_M1011_g N_Y_c_457_n 0.00489466f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A1_M1011_g N_Y_c_458_n 0.0146133f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_141 N_A1_c_135_n N_Y_c_458_n 0.0146656f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_142 N_A1_c_132_n N_Y_c_458_n 0.00178697f $X=1.985 $Y=1.537 $X2=0 $Y2=0
cc_143 N_A1_c_133_n N_Y_c_470_n 0.0129773f $X=1.505 $Y=1.725 $X2=0 $Y2=0
cc_144 N_A1_c_135_n N_Y_c_470_n 0.0264917f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_145 N_A1_c_132_n N_Y_c_470_n 0.007249f $X=1.985 $Y=1.537 $X2=0 $Y2=0
cc_146 N_A1_M1018_g N_Y_c_482_n 0.00579199f $X=1.985 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A1_c_133_n N_Y_c_463_n 0.00324782f $X=1.505 $Y=1.725 $X2=0 $Y2=0
cc_148 N_A1_c_134_n N_Y_c_463_n 0.00387175f $X=2.245 $Y=1.725 $X2=0 $Y2=0
cc_149 N_A1_c_132_n N_Y_c_463_n 0.00550079f $X=1.985 $Y=1.537 $X2=0 $Y2=0
cc_150 N_A1_c_133_n N_Y_c_472_n 7.34652e-19 $X=1.505 $Y=1.725 $X2=0 $Y2=0
cc_151 N_A1_c_132_n N_Y_c_460_n 0.0159795f $X=1.985 $Y=1.537 $X2=0 $Y2=0
cc_152 N_A1_M1011_g N_Y_c_461_n 0.00243405f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A1_M1018_g N_Y_c_461_n 0.0147903f $X=1.985 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A1_c_135_n N_Y_c_461_n 0.00925742f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_155 N_A1_c_132_n N_Y_c_461_n 0.0032074f $X=1.985 $Y=1.537 $X2=0 $Y2=0
cc_156 N_A1_M1011_g Y 4.94356e-19 $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A1_M1018_g Y 0.00302831f $X=1.985 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A1_c_135_n Y 0.0263674f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_159 N_A1_c_132_n Y 0.00773729f $X=1.985 $Y=1.537 $X2=0 $Y2=0
cc_160 N_A1_c_133_n N_VPWR_c_525_n 0.00448106f $X=1.505 $Y=1.725 $X2=0 $Y2=0
cc_161 N_A1_c_134_n N_VPWR_c_525_n 0.00507697f $X=2.245 $Y=1.725 $X2=0 $Y2=0
cc_162 N_A1_c_134_n N_VPWR_c_529_n 0.005209f $X=2.245 $Y=1.725 $X2=0 $Y2=0
cc_163 N_A1_c_133_n N_VPWR_c_533_n 0.00517089f $X=1.505 $Y=1.725 $X2=0 $Y2=0
cc_164 N_A1_c_133_n N_VPWR_c_524_n 0.00979649f $X=1.505 $Y=1.725 $X2=0 $Y2=0
cc_165 N_A1_c_134_n N_VPWR_c_524_n 0.00983982f $X=2.245 $Y=1.725 $X2=0 $Y2=0
cc_166 N_A1_M1011_g N_VGND_c_601_n 0.00278247f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A1_M1018_g N_VGND_c_601_n 0.00278271f $X=1.985 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A1_M1011_g N_VGND_c_603_n 0.00358425f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A1_M1018_g N_VGND_c_603_n 0.0035414f $X=1.985 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A1_M1011_g N_A_239_74#_c_651_n 0.00709316f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A1_M1018_g N_A_239_74#_c_651_n 4.4915e-19 $X=1.985 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A1_M1011_g N_A_239_74#_c_652_n 0.00792642f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A1_M1018_g N_A_239_74#_c_652_n 0.0110411f $X=1.985 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A1_M1011_g N_A_239_74#_c_653_n 0.00395315f $X=1.555 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A1_c_132_n N_A_239_74#_c_662_n 0.00224943f $X=1.985 $Y=1.537 $X2=0
+ $Y2=0
cc_176 N_A2_M1005_g N_A3_M1000_g 0.01694f $X=3.245 $Y=2.4 $X2=0 $Y2=0
cc_177 A2 N_A3_M1000_g 0.00990912f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_178 A2 N_A3_M1004_g 0.00154933f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_179 N_A2_c_200_n N_A3_M1004_g 0.00482007f $X=3.17 $Y=1.465 $X2=0 $Y2=0
cc_180 A2 A3 0.0279378f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_181 A2 N_A3_c_267_n 0.00776743f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_182 N_A2_c_200_n N_A3_c_267_n 0.01694f $X=3.17 $Y=1.465 $X2=0 $Y2=0
cc_183 N_A2_M1001_g N_A_27_368#_c_364_n 0.00492664f $X=2.695 $Y=2.4 $X2=0 $Y2=0
cc_184 N_A2_M1005_g N_A_27_368#_c_364_n 5.96661e-19 $X=3.245 $Y=2.4 $X2=0 $Y2=0
cc_185 N_A2_c_200_n N_A_27_368#_c_364_n 0.00677746f $X=3.17 $Y=1.465 $X2=0 $Y2=0
cc_186 N_A2_M1001_g N_A_27_368#_c_383_n 0.00384899f $X=2.695 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A2_M1005_g N_A_27_368#_c_383_n 3.46565e-19 $X=3.245 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A2_M1001_g N_A_27_368#_c_365_n 0.0066771f $X=2.695 $Y=2.4 $X2=0 $Y2=0
cc_189 N_A2_M1001_g N_A_27_368#_c_392_n 0.0150458f $X=2.695 $Y=2.4 $X2=0 $Y2=0
cc_190 N_A2_M1005_g N_A_27_368#_c_392_n 0.0134861f $X=3.245 $Y=2.4 $X2=0 $Y2=0
cc_191 A2 N_A_27_368#_c_392_n 0.0138359f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_192 A2 N_A_27_368#_c_392_n 0.0209965f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_193 N_A2_c_200_n N_A_27_368#_c_392_n 0.00331749f $X=3.17 $Y=1.465 $X2=0 $Y2=0
cc_194 N_A2_M1001_g N_A_27_368#_c_366_n 4.92941e-19 $X=2.695 $Y=2.4 $X2=0 $Y2=0
cc_195 N_A2_M1005_g N_A_27_368#_c_366_n 0.0119155f $X=3.245 $Y=2.4 $X2=0 $Y2=0
cc_196 A2 N_A_27_368#_c_399_n 0.00585617f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_197 N_A2_M1001_g N_A_27_368#_c_385_n 0.00193648f $X=2.695 $Y=2.4 $X2=0 $Y2=0
cc_198 N_A2_M1005_g N_A_27_368#_c_401_n 8.84614e-19 $X=3.245 $Y=2.4 $X2=0 $Y2=0
cc_199 A2 N_A_27_368#_c_401_n 0.0237863f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_200 N_A2_M1001_g N_Y_c_463_n 3.26833e-19 $X=2.695 $Y=2.4 $X2=0 $Y2=0
cc_201 N_A2_c_200_n N_Y_c_460_n 3.4212e-19 $X=3.17 $Y=1.465 $X2=0 $Y2=0
cc_202 N_A2_c_195_n N_Y_c_461_n 0.00538827f $X=2.485 $Y=1.185 $X2=0 $Y2=0
cc_203 A2 Y 0.0144379f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_204 N_A2_c_200_n Y 0.0039377f $X=3.17 $Y=1.465 $X2=0 $Y2=0
cc_205 N_A2_M1001_g N_VPWR_c_526_n 0.00212994f $X=2.695 $Y=2.4 $X2=0 $Y2=0
cc_206 N_A2_M1005_g N_VPWR_c_526_n 0.00212994f $X=3.245 $Y=2.4 $X2=0 $Y2=0
cc_207 N_A2_M1001_g N_VPWR_c_529_n 0.005209f $X=2.695 $Y=2.4 $X2=0 $Y2=0
cc_208 N_A2_M1005_g N_VPWR_c_531_n 0.005209f $X=3.245 $Y=2.4 $X2=0 $Y2=0
cc_209 N_A2_M1001_g N_VPWR_c_524_n 0.00982636f $X=2.695 $Y=2.4 $X2=0 $Y2=0
cc_210 N_A2_M1005_g N_VPWR_c_524_n 0.00982636f $X=3.245 $Y=2.4 $X2=0 $Y2=0
cc_211 N_A2_c_195_n N_VGND_c_601_n 0.00329872f $X=2.485 $Y=1.185 $X2=0 $Y2=0
cc_212 N_A2_c_197_n N_VGND_c_601_n 0.00288916f $X=2.915 $Y=1.185 $X2=0 $Y2=0
cc_213 N_A2_c_195_n N_VGND_c_603_n 0.0042865f $X=2.485 $Y=1.185 $X2=0 $Y2=0
cc_214 N_A2_c_197_n N_VGND_c_603_n 0.00361255f $X=2.915 $Y=1.185 $X2=0 $Y2=0
cc_215 N_A2_c_195_n N_A_239_74#_c_652_n 0.00282675f $X=2.485 $Y=1.185 $X2=0
+ $Y2=0
cc_216 N_A2_c_195_n N_A_239_74#_c_664_n 0.0139295f $X=2.485 $Y=1.185 $X2=0 $Y2=0
cc_217 N_A2_c_197_n N_A_239_74#_c_664_n 0.00887373f $X=2.915 $Y=1.185 $X2=0
+ $Y2=0
cc_218 A2 N_A_239_74#_c_664_n 0.0104844f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_219 N_A2_c_200_n N_A_239_74#_c_664_n 0.0027376f $X=3.17 $Y=1.465 $X2=0 $Y2=0
cc_220 N_A2_c_195_n N_A_239_74#_c_654_n 8.61657e-19 $X=2.485 $Y=1.185 $X2=0
+ $Y2=0
cc_221 N_A2_c_197_n N_A_239_74#_c_654_n 0.00450644f $X=2.915 $Y=1.185 $X2=0
+ $Y2=0
cc_222 A2 N_A_239_74#_c_654_n 0.0194992f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_223 N_A2_c_200_n N_A_239_74#_c_654_n 0.00860041f $X=3.17 $Y=1.465 $X2=0 $Y2=0
cc_224 N_A2_c_195_n N_A_512_74#_c_696_n 0.00360761f $X=2.485 $Y=1.185 $X2=0
+ $Y2=0
cc_225 N_A2_c_197_n N_A_512_74#_c_696_n 0.013308f $X=2.915 $Y=1.185 $X2=0 $Y2=0
cc_226 N_A2_c_200_n N_A_512_74#_c_696_n 0.00139415f $X=3.17 $Y=1.465 $X2=0 $Y2=0
cc_227 N_A2_c_197_n N_A_709_74#_c_716_n 0.00102896f $X=2.915 $Y=1.185 $X2=0
+ $Y2=0
cc_228 A2 N_A_709_74#_c_716_n 0.0160865f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_229 N_A3_M1017_g N_A4_M1014_g 0.01695f $X=4.335 $Y=0.74 $X2=0 $Y2=0
cc_230 N_A3_M1003_g N_A4_M1008_g 0.0255613f $X=4.245 $Y=2.4 $X2=0 $Y2=0
cc_231 A3 A4 0.0291763f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_232 N_A3_c_267_n A4 2.08437e-19 $X=4.245 $Y=1.515 $X2=0 $Y2=0
cc_233 A3 N_A4_c_324_n 0.00519974f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_234 N_A3_c_267_n N_A4_c_324_n 0.01695f $X=4.245 $Y=1.515 $X2=0 $Y2=0
cc_235 N_A3_M1000_g N_A_27_368#_c_366_n 0.0119155f $X=3.695 $Y=2.4 $X2=0 $Y2=0
cc_236 N_A3_M1003_g N_A_27_368#_c_366_n 4.92941e-19 $X=4.245 $Y=2.4 $X2=0 $Y2=0
cc_237 N_A3_M1000_g N_A_27_368#_c_399_n 0.0155005f $X=3.695 $Y=2.4 $X2=0 $Y2=0
cc_238 N_A3_M1003_g N_A_27_368#_c_399_n 0.0134861f $X=4.245 $Y=2.4 $X2=0 $Y2=0
cc_239 A3 N_A_27_368#_c_399_n 0.0239743f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_240 N_A3_c_267_n N_A_27_368#_c_399_n 0.0053207f $X=4.245 $Y=1.515 $X2=0 $Y2=0
cc_241 N_A3_M1000_g N_A_27_368#_c_367_n 4.96476e-19 $X=3.695 $Y=2.4 $X2=0 $Y2=0
cc_242 N_A3_M1003_g N_A_27_368#_c_367_n 0.012643f $X=4.245 $Y=2.4 $X2=0 $Y2=0
cc_243 N_A3_M1000_g N_A_27_368#_c_401_n 8.84614e-19 $X=3.695 $Y=2.4 $X2=0 $Y2=0
cc_244 N_A3_M1003_g N_A_27_368#_c_412_n 8.84614e-19 $X=4.245 $Y=2.4 $X2=0 $Y2=0
cc_245 A3 N_A_27_368#_c_412_n 0.0277936f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_246 N_A3_c_267_n N_A_27_368#_c_412_n 3.1404e-19 $X=4.245 $Y=1.515 $X2=0 $Y2=0
cc_247 N_A3_M1000_g N_VPWR_c_527_n 0.00212994f $X=3.695 $Y=2.4 $X2=0 $Y2=0
cc_248 N_A3_M1003_g N_VPWR_c_527_n 0.00312091f $X=4.245 $Y=2.4 $X2=0 $Y2=0
cc_249 N_A3_M1003_g N_VPWR_c_528_n 6.00394e-19 $X=4.245 $Y=2.4 $X2=0 $Y2=0
cc_250 N_A3_M1000_g N_VPWR_c_531_n 0.005209f $X=3.695 $Y=2.4 $X2=0 $Y2=0
cc_251 N_A3_M1003_g N_VPWR_c_534_n 0.00520371f $X=4.245 $Y=2.4 $X2=0 $Y2=0
cc_252 N_A3_M1000_g N_VPWR_c_524_n 0.00982636f $X=3.695 $Y=2.4 $X2=0 $Y2=0
cc_253 N_A3_M1003_g N_VPWR_c_524_n 0.00983018f $X=4.245 $Y=2.4 $X2=0 $Y2=0
cc_254 N_A3_M1017_g N_VGND_c_600_n 6.60052e-19 $X=4.335 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A3_M1004_g N_VGND_c_601_n 0.00288916f $X=3.905 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A3_M1017_g N_VGND_c_601_n 0.00432706f $X=4.335 $Y=0.74 $X2=0 $Y2=0
cc_257 N_A3_M1004_g N_VGND_c_603_n 0.00362189f $X=3.905 $Y=0.74 $X2=0 $Y2=0
cc_258 N_A3_M1017_g N_VGND_c_603_n 0.00448861f $X=4.335 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A3_M1004_g N_A_239_74#_c_654_n 0.00145088f $X=3.905 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A3_M1004_g N_A_512_74#_c_695_n 0.00588379f $X=3.905 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A3_M1017_g N_A_512_74#_c_695_n 0.00476696f $X=4.335 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A3_M1004_g N_A_512_74#_c_696_n 0.0121895f $X=3.905 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A3_M1004_g N_A_709_74#_c_716_n 0.0161611f $X=3.905 $Y=0.74 $X2=0 $Y2=0
cc_264 N_A3_M1017_g N_A_709_74#_c_716_n 0.0132419f $X=4.335 $Y=0.74 $X2=0 $Y2=0
cc_265 A3 N_A_709_74#_c_716_n 0.0323753f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_266 N_A3_c_267_n N_A_709_74#_c_716_n 0.00736176f $X=4.245 $Y=1.515 $X2=0
+ $Y2=0
cc_267 N_A3_M1017_g N_A_709_74#_c_717_n 3.92031e-19 $X=4.335 $Y=0.74 $X2=0 $Y2=0
cc_268 A3 N_A_709_74#_c_718_n 0.00320175f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_269 N_A3_M1017_g N_A_709_74#_c_720_n 0.00158218f $X=4.335 $Y=0.74 $X2=0 $Y2=0
cc_270 A3 N_A_709_74#_c_720_n 0.0153286f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_271 N_A4_M1008_g N_A_27_368#_c_367_n 0.00523548f $X=4.78 $Y=2.4 $X2=0 $Y2=0
cc_272 N_A4_M1008_g N_A_27_368#_c_416_n 0.0221979f $X=4.78 $Y=2.4 $X2=0 $Y2=0
cc_273 N_A4_M1012_g N_A_27_368#_c_416_n 0.0142562f $X=5.23 $Y=2.4 $X2=0 $Y2=0
cc_274 A4 N_A_27_368#_c_416_n 0.0289485f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_275 N_A4_c_324_n N_A_27_368#_c_416_n 4.90767e-19 $X=5.245 $Y=1.515 $X2=0
+ $Y2=0
cc_276 A4 N_A_27_368#_c_368_n 0.0244344f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_277 N_A4_M1012_g N_A_27_368#_c_369_n 0.00137891f $X=5.23 $Y=2.4 $X2=0 $Y2=0
cc_278 N_A4_M1008_g N_VPWR_c_528_n 0.0127956f $X=4.78 $Y=2.4 $X2=0 $Y2=0
cc_279 N_A4_M1012_g N_VPWR_c_528_n 0.0151142f $X=5.23 $Y=2.4 $X2=0 $Y2=0
cc_280 N_A4_M1008_g N_VPWR_c_534_n 0.00460063f $X=4.78 $Y=2.4 $X2=0 $Y2=0
cc_281 N_A4_M1012_g N_VPWR_c_535_n 0.00460063f $X=5.23 $Y=2.4 $X2=0 $Y2=0
cc_282 N_A4_M1008_g N_VPWR_c_524_n 0.00909416f $X=4.78 $Y=2.4 $X2=0 $Y2=0
cc_283 N_A4_M1012_g N_VPWR_c_524_n 0.0091238f $X=5.23 $Y=2.4 $X2=0 $Y2=0
cc_284 N_A4_M1014_g N_VGND_c_600_n 0.0107027f $X=4.765 $Y=0.74 $X2=0 $Y2=0
cc_285 N_A4_M1015_g N_VGND_c_600_n 0.00388319f $X=5.245 $Y=0.74 $X2=0 $Y2=0
cc_286 N_A4_M1014_g N_VGND_c_601_n 0.00383152f $X=4.765 $Y=0.74 $X2=0 $Y2=0
cc_287 N_A4_M1015_g N_VGND_c_602_n 0.00456932f $X=5.245 $Y=0.74 $X2=0 $Y2=0
cc_288 N_A4_M1014_g N_VGND_c_603_n 0.00757637f $X=4.765 $Y=0.74 $X2=0 $Y2=0
cc_289 N_A4_M1015_g N_VGND_c_603_n 0.00893404f $X=5.245 $Y=0.74 $X2=0 $Y2=0
cc_290 N_A4_M1014_g N_A_709_74#_c_717_n 3.92313e-19 $X=4.765 $Y=0.74 $X2=0 $Y2=0
cc_291 N_A4_M1014_g N_A_709_74#_c_718_n 0.0178155f $X=4.765 $Y=0.74 $X2=0 $Y2=0
cc_292 N_A4_M1015_g N_A_709_74#_c_718_n 0.0144542f $X=5.245 $Y=0.74 $X2=0 $Y2=0
cc_293 A4 N_A_709_74#_c_718_n 0.0581505f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_294 N_A4_c_324_n N_A_709_74#_c_718_n 0.00359948f $X=5.245 $Y=1.515 $X2=0
+ $Y2=0
cc_295 N_A4_M1014_g N_A_709_74#_c_719_n 8.86531e-19 $X=4.765 $Y=0.74 $X2=0 $Y2=0
cc_296 N_A4_M1015_g N_A_709_74#_c_719_n 0.00890364f $X=5.245 $Y=0.74 $X2=0 $Y2=0
cc_297 N_A_27_368#_c_362_n N_Y_M1007_s 0.00218982f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_298 N_A_27_368#_M1009_d N_Y_c_470_n 0.0100499f $X=1.095 $Y=1.84 $X2=0 $Y2=0
cc_299 N_A_27_368#_c_377_n N_Y_c_470_n 0.0189689f $X=1.28 $Y=2.46 $X2=0 $Y2=0
cc_300 N_A_27_368#_c_379_n N_Y_c_470_n 0.0436069f $X=2.305 $Y=2.375 $X2=0 $Y2=0
cc_301 N_A_27_368#_c_364_n N_Y_c_463_n 0.00562343f $X=2.47 $Y=2.12 $X2=0 $Y2=0
cc_302 N_A_27_368#_c_362_n N_Y_c_472_n 0.0177084f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_303 N_A_27_368#_c_379_n N_Y_c_460_n 0.00322071f $X=2.305 $Y=2.375 $X2=0 $Y2=0
cc_304 N_A_27_368#_c_379_n N_VPWR_M1002_s 0.0111892f $X=2.305 $Y=2.375 $X2=-0.19
+ $Y2=1.66
cc_305 N_A_27_368#_c_392_n N_VPWR_M1001_s 0.0056699f $X=3.305 $Y=2.035 $X2=0
+ $Y2=0
cc_306 N_A_27_368#_c_399_n N_VPWR_M1000_s 0.0058542f $X=4.305 $Y=2.035 $X2=0
+ $Y2=0
cc_307 N_A_27_368#_c_416_n N_VPWR_M1008_d 0.00314376f $X=5.34 $Y=2.035 $X2=0
+ $Y2=0
cc_308 N_A_27_368#_c_362_n N_VPWR_c_525_n 0.0122626f $X=1.115 $Y=2.99 $X2=0
+ $Y2=0
cc_309 N_A_27_368#_c_379_n N_VPWR_c_525_n 0.0333945f $X=2.305 $Y=2.375 $X2=0
+ $Y2=0
cc_310 N_A_27_368#_c_365_n N_VPWR_c_525_n 0.0132291f $X=2.47 $Y=2.815 $X2=0
+ $Y2=0
cc_311 N_A_27_368#_c_365_n N_VPWR_c_526_n 0.0202646f $X=2.47 $Y=2.815 $X2=0
+ $Y2=0
cc_312 N_A_27_368#_c_392_n N_VPWR_c_526_n 0.0208278f $X=3.305 $Y=2.035 $X2=0
+ $Y2=0
cc_313 N_A_27_368#_c_366_n N_VPWR_c_526_n 0.0266809f $X=3.47 $Y=2.815 $X2=0
+ $Y2=0
cc_314 N_A_27_368#_c_366_n N_VPWR_c_527_n 0.0266809f $X=3.47 $Y=2.815 $X2=0
+ $Y2=0
cc_315 N_A_27_368#_c_399_n N_VPWR_c_527_n 0.0208278f $X=4.305 $Y=2.035 $X2=0
+ $Y2=0
cc_316 N_A_27_368#_c_367_n N_VPWR_c_527_n 0.0286777f $X=4.485 $Y=2.44 $X2=0
+ $Y2=0
cc_317 N_A_27_368#_c_367_n N_VPWR_c_528_n 0.0282884f $X=4.485 $Y=2.44 $X2=0
+ $Y2=0
cc_318 N_A_27_368#_c_416_n N_VPWR_c_528_n 0.0170259f $X=5.34 $Y=2.035 $X2=0
+ $Y2=0
cc_319 N_A_27_368#_c_369_n N_VPWR_c_528_n 0.0282442f $X=5.465 $Y=2.44 $X2=0
+ $Y2=0
cc_320 N_A_27_368#_c_365_n N_VPWR_c_529_n 0.0144623f $X=2.47 $Y=2.815 $X2=0
+ $Y2=0
cc_321 N_A_27_368#_c_366_n N_VPWR_c_531_n 0.0144623f $X=3.47 $Y=2.815 $X2=0
+ $Y2=0
cc_322 N_A_27_368#_c_362_n N_VPWR_c_533_n 0.0656628f $X=1.115 $Y=2.99 $X2=0
+ $Y2=0
cc_323 N_A_27_368#_c_363_n N_VPWR_c_533_n 0.0235512f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_324 N_A_27_368#_c_367_n N_VPWR_c_534_n 0.0175179f $X=4.485 $Y=2.44 $X2=0
+ $Y2=0
cc_325 N_A_27_368#_c_369_n N_VPWR_c_535_n 0.0146972f $X=5.465 $Y=2.44 $X2=0
+ $Y2=0
cc_326 N_A_27_368#_c_362_n N_VPWR_c_524_n 0.036369f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_327 N_A_27_368#_c_363_n N_VPWR_c_524_n 0.0126924f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_328 N_A_27_368#_c_365_n N_VPWR_c_524_n 0.0118344f $X=2.47 $Y=2.815 $X2=0
+ $Y2=0
cc_329 N_A_27_368#_c_366_n N_VPWR_c_524_n 0.0118344f $X=3.47 $Y=2.815 $X2=0
+ $Y2=0
cc_330 N_A_27_368#_c_367_n N_VPWR_c_524_n 0.0134273f $X=4.485 $Y=2.44 $X2=0
+ $Y2=0
cc_331 N_A_27_368#_c_369_n N_VPWR_c_524_n 0.0113236f $X=5.465 $Y=2.44 $X2=0
+ $Y2=0
cc_332 N_Y_c_470_n N_VPWR_M1002_s 0.0110685f $X=1.965 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_333 N_Y_c_463_n N_VPWR_M1002_s 0.00181463f $X=2.05 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_334 N_Y_c_457_n N_VGND_c_599_n 0.0236416f $X=0.78 $Y=0.565 $X2=0 $Y2=0
cc_335 N_Y_c_459_n N_VGND_c_599_n 0.00795492f $X=0.945 $Y=1.095 $X2=0 $Y2=0
cc_336 N_Y_c_457_n N_VGND_c_601_n 0.0121139f $X=0.78 $Y=0.565 $X2=0 $Y2=0
cc_337 N_Y_c_457_n N_VGND_c_603_n 0.0117201f $X=0.78 $Y=0.565 $X2=0 $Y2=0
cc_338 N_Y_c_458_n N_A_239_74#_M1011_s 0.00299905f $X=1.685 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_339 N_Y_c_461_n N_A_239_74#_M1018_s 0.00201792f $X=2.12 $Y=1.26 $X2=0 $Y2=0
cc_340 N_Y_c_457_n N_A_239_74#_c_651_n 0.027945f $X=0.78 $Y=0.565 $X2=0 $Y2=0
cc_341 N_Y_c_458_n N_A_239_74#_c_651_n 0.021673f $X=1.685 $Y=1.095 $X2=0 $Y2=0
cc_342 N_Y_M1011_d N_A_239_74#_c_652_n 0.00176461f $X=1.63 $Y=0.37 $X2=0 $Y2=0
cc_343 N_Y_c_458_n N_A_239_74#_c_652_n 0.00304353f $X=1.685 $Y=1.095 $X2=0 $Y2=0
cc_344 N_Y_c_482_n N_A_239_74#_c_652_n 0.014283f $X=1.77 $Y=0.76 $X2=0 $Y2=0
cc_345 N_Y_c_461_n N_A_239_74#_c_652_n 0.00296068f $X=2.12 $Y=1.26 $X2=0 $Y2=0
cc_346 N_Y_c_457_n N_A_239_74#_c_653_n 0.00178848f $X=0.78 $Y=0.565 $X2=0 $Y2=0
cc_347 N_Y_c_461_n N_A_239_74#_c_662_n 0.0140442f $X=2.12 $Y=1.26 $X2=0 $Y2=0
cc_348 N_VGND_c_601_n N_A_239_74#_c_652_n 0.0556865f $X=4.815 $Y=0 $X2=0 $Y2=0
cc_349 N_VGND_c_603_n N_A_239_74#_c_652_n 0.0310135f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_350 N_VGND_c_601_n N_A_239_74#_c_653_n 0.0233048f $X=4.815 $Y=0 $X2=0 $Y2=0
cc_351 N_VGND_c_603_n N_A_239_74#_c_653_n 0.0126653f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_352 N_VGND_c_601_n N_A_239_74#_c_664_n 0.00197884f $X=4.815 $Y=0 $X2=0 $Y2=0
cc_353 N_VGND_c_603_n N_A_239_74#_c_664_n 0.00471412f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_354 N_VGND_c_600_n N_A_512_74#_c_695_n 5.95781e-19 $X=4.98 $Y=0.675 $X2=0
+ $Y2=0
cc_355 N_VGND_c_601_n N_A_512_74#_c_696_n 0.0780839f $X=4.815 $Y=0 $X2=0 $Y2=0
cc_356 N_VGND_c_603_n N_A_512_74#_c_696_n 0.0618436f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_357 N_VGND_c_603_n N_A_709_74#_c_716_n 0.00692405f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_358 N_VGND_c_600_n N_A_709_74#_c_717_n 0.0182488f $X=4.98 $Y=0.675 $X2=0
+ $Y2=0
cc_359 N_VGND_c_601_n N_A_709_74#_c_717_n 0.00749631f $X=4.815 $Y=0 $X2=0 $Y2=0
cc_360 N_VGND_c_603_n N_A_709_74#_c_717_n 0.0062048f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_361 N_VGND_M1014_s N_A_709_74#_c_718_n 0.00229612f $X=4.84 $Y=0.37 $X2=0
+ $Y2=0
cc_362 N_VGND_c_600_n N_A_709_74#_c_718_n 0.0193595f $X=4.98 $Y=0.675 $X2=0
+ $Y2=0
cc_363 N_VGND_c_600_n N_A_709_74#_c_719_n 0.0191764f $X=4.98 $Y=0.675 $X2=0
+ $Y2=0
cc_364 N_VGND_c_602_n N_A_709_74#_c_719_n 0.0146237f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_365 N_VGND_c_603_n N_A_709_74#_c_719_n 0.0120948f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_366 N_A_239_74#_c_664_n N_A_512_74#_M1010_s 0.0047246f $X=2.965 $Y=0.835
+ $X2=-0.19 $Y2=-0.245
cc_367 N_A_239_74#_M1016_d N_A_512_74#_c_696_n 0.00346043f $X=2.99 $Y=0.37 $X2=0
+ $Y2=0
cc_368 N_A_239_74#_c_652_n N_A_512_74#_c_696_n 0.00550602f $X=2.105 $Y=0.34
+ $X2=0 $Y2=0
cc_369 N_A_239_74#_c_664_n N_A_512_74#_c_696_n 0.0220487f $X=2.965 $Y=0.835
+ $X2=0 $Y2=0
cc_370 N_A_239_74#_c_654_n N_A_512_74#_c_696_n 0.02055f $X=3.13 $Y=0.835 $X2=0
+ $Y2=0
cc_371 N_A_239_74#_c_654_n N_A_709_74#_c_716_n 0.0163825f $X=3.13 $Y=0.835 $X2=0
+ $Y2=0
cc_372 N_A_512_74#_c_696_n N_A_709_74#_M1004_d 0.0042464f $X=3.955 $Y=0.505
+ $X2=-0.19 $Y2=-0.245
cc_373 N_A_512_74#_M1004_s N_A_709_74#_c_716_n 0.00177318f $X=3.98 $Y=0.37 $X2=0
+ $Y2=0
cc_374 N_A_512_74#_c_695_n N_A_709_74#_c_716_n 0.0164606f $X=4.12 $Y=0.515 $X2=0
+ $Y2=0
cc_375 N_A_512_74#_c_696_n N_A_709_74#_c_716_n 0.0184982f $X=3.955 $Y=0.505
+ $X2=0 $Y2=0
cc_376 N_A_512_74#_c_695_n N_A_709_74#_c_717_n 0.0135087f $X=4.12 $Y=0.515 $X2=0
+ $Y2=0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor4bb_1 A B C_N D_N VGND VNB VPB VPWR Y
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 VGND D_N a_611_244# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X2 a_400_368# a_27_112# a_533_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 Y a_611_244# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_27_112# C_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X6 a_533_368# a_611_244# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 VPWR A a_316_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 a_316_368# B a_400_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X9 VGND a_27_112# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 VPWR D_N a_611_244# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X11 a_27_112# C_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
.ends

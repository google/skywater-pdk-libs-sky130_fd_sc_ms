* File: sky130_fd_sc_ms__nor4b_4.pxi.spice
* Created: Wed Sep  2 12:17:10 2020
* 
x_PM_SKY130_FD_SC_MS__NOR4B_4%D_N N_D_N_c_149_n N_D_N_M1012_g N_D_N_M1013_g
+ N_D_N_c_150_n N_D_N_M1010_g D_N D_N N_D_N_c_151_n
+ PM_SKY130_FD_SC_MS__NOR4B_4%D_N
x_PM_SKY130_FD_SC_MS__NOR4B_4%A_47_88# N_A_47_88#_M1010_s N_A_47_88#_M1012_d
+ N_A_47_88#_M1002_g N_A_47_88#_M1003_g N_A_47_88#_c_193_n N_A_47_88#_M1022_g
+ N_A_47_88#_c_194_n N_A_47_88#_M1024_g N_A_47_88#_M1011_g N_A_47_88#_M1028_g
+ N_A_47_88#_c_195_n N_A_47_88#_M1026_g N_A_47_88#_c_188_n N_A_47_88#_c_189_n
+ N_A_47_88#_c_198_n N_A_47_88#_M1027_g N_A_47_88#_c_190_n N_A_47_88#_c_199_n
+ N_A_47_88#_c_293_p N_A_47_88#_c_191_n N_A_47_88#_c_192_n N_A_47_88#_c_200_n
+ N_A_47_88#_c_215_n PM_SKY130_FD_SC_MS__NOR4B_4%A_47_88#
x_PM_SKY130_FD_SC_MS__NOR4B_4%C N_C_c_304_n N_C_M1006_g N_C_c_305_n N_C_M1000_g
+ N_C_c_306_n N_C_M1025_g N_C_M1001_g N_C_M1031_g N_C_c_307_n N_C_M1030_g
+ N_C_c_308_n N_C_c_309_n N_C_M1034_g N_C_M1032_g N_C_c_311_n C C C N_C_c_313_n
+ N_C_c_314_n PM_SKY130_FD_SC_MS__NOR4B_4%C
x_PM_SKY130_FD_SC_MS__NOR4B_4%B N_B_M1004_g N_B_M1014_g N_B_M1008_g N_B_M1016_g
+ N_B_M1009_g N_B_M1017_g N_B_M1019_g N_B_M1018_g B B B B N_B_c_405_n
+ PM_SKY130_FD_SC_MS__NOR4B_4%B
x_PM_SKY130_FD_SC_MS__NOR4B_4%A N_A_M1020_g N_A_M1005_g N_A_M1007_g N_A_M1021_g
+ N_A_M1015_g N_A_M1023_g N_A_M1029_g N_A_M1033_g A A A A N_A_c_499_n
+ PM_SKY130_FD_SC_MS__NOR4B_4%A
x_PM_SKY130_FD_SC_MS__NOR4B_4%VPWR N_VPWR_M1012_s N_VPWR_M1013_s N_VPWR_M1020_d
+ N_VPWR_M1023_d N_VPWR_c_577_n N_VPWR_c_578_n N_VPWR_c_579_n N_VPWR_c_580_n
+ N_VPWR_c_581_n VPWR N_VPWR_c_582_n N_VPWR_c_583_n N_VPWR_c_584_n
+ N_VPWR_c_585_n N_VPWR_c_576_n N_VPWR_c_587_n N_VPWR_c_588_n N_VPWR_c_589_n
+ PM_SKY130_FD_SC_MS__NOR4B_4%VPWR
x_PM_SKY130_FD_SC_MS__NOR4B_4%A_319_368# N_A_319_368#_M1022_s
+ N_A_319_368#_M1024_s N_A_319_368#_M1027_s N_A_319_368#_M1001_s
+ N_A_319_368#_M1032_s N_A_319_368#_c_680_n N_A_319_368#_c_681_n
+ N_A_319_368#_c_682_n N_A_319_368#_c_721_p N_A_319_368#_c_683_n
+ N_A_319_368#_c_695_n N_A_319_368#_c_696_n N_A_319_368#_c_684_n
+ N_A_319_368#_c_698_n N_A_319_368#_c_700_n N_A_319_368#_c_685_n
+ N_A_319_368#_c_702_n PM_SKY130_FD_SC_MS__NOR4B_4%A_319_368#
x_PM_SKY130_FD_SC_MS__NOR4B_4%Y N_Y_M1002_d N_Y_M1011_d N_Y_M1006_s N_Y_M1030_s
+ N_Y_M1004_d N_Y_M1009_d N_Y_M1005_d N_Y_M1015_d N_Y_M1022_d N_Y_M1026_d
+ N_Y_c_745_n N_Y_c_746_n N_Y_c_747_n N_Y_c_767_n N_Y_c_784_n N_Y_c_768_n
+ N_Y_c_748_n N_Y_c_749_n N_Y_c_795_n N_Y_c_797_n N_Y_c_750_n N_Y_c_751_n
+ N_Y_c_752_n N_Y_c_753_n N_Y_c_754_n N_Y_c_755_n N_Y_c_756_n N_Y_c_757_n
+ N_Y_c_758_n N_Y_c_759_n N_Y_c_760_n N_Y_c_761_n N_Y_c_799_n N_Y_c_769_n
+ N_Y_c_762_n N_Y_c_763_n N_Y_c_764_n N_Y_c_765_n Y Y
+ PM_SKY130_FD_SC_MS__NOR4B_4%Y
x_PM_SKY130_FD_SC_MS__NOR4B_4%A_781_368# N_A_781_368#_M1000_d
+ N_A_781_368#_M1031_d N_A_781_368#_M1014_d N_A_781_368#_M1017_d
+ N_A_781_368#_c_946_n N_A_781_368#_c_947_n N_A_781_368#_c_962_n
+ N_A_781_368#_c_948_n N_A_781_368#_c_967_n N_A_781_368#_c_949_n
+ N_A_781_368#_c_950_n N_A_781_368#_c_951_n
+ PM_SKY130_FD_SC_MS__NOR4B_4%A_781_368#
x_PM_SKY130_FD_SC_MS__NOR4B_4%A_1191_368# N_A_1191_368#_M1014_s
+ N_A_1191_368#_M1016_s N_A_1191_368#_M1018_s N_A_1191_368#_M1021_s
+ N_A_1191_368#_M1033_s N_A_1191_368#_c_1013_n N_A_1191_368#_c_1017_n
+ N_A_1191_368#_c_1019_n N_A_1191_368#_c_1007_n N_A_1191_368#_c_1033_n
+ N_A_1191_368#_c_1008_n N_A_1191_368#_c_1041_n N_A_1191_368#_c_1009_n
+ N_A_1191_368#_c_1010_n N_A_1191_368#_c_1011_n N_A_1191_368#_c_1028_n
+ N_A_1191_368#_c_1047_n N_A_1191_368#_c_1048_n
+ PM_SKY130_FD_SC_MS__NOR4B_4%A_1191_368#
x_PM_SKY130_FD_SC_MS__NOR4B_4%VGND N_VGND_M1010_d N_VGND_M1003_s N_VGND_M1028_s
+ N_VGND_M1025_d N_VGND_M1034_d N_VGND_M1008_s N_VGND_M1019_s N_VGND_M1007_s
+ N_VGND_M1029_s N_VGND_c_1077_n N_VGND_c_1078_n N_VGND_c_1079_n N_VGND_c_1080_n
+ N_VGND_c_1081_n N_VGND_c_1082_n N_VGND_c_1083_n N_VGND_c_1084_n
+ N_VGND_c_1085_n VGND N_VGND_c_1086_n N_VGND_c_1087_n N_VGND_c_1088_n
+ N_VGND_c_1089_n N_VGND_c_1090_n N_VGND_c_1091_n N_VGND_c_1092_n
+ N_VGND_c_1093_n N_VGND_c_1094_n N_VGND_c_1095_n N_VGND_c_1096_n
+ N_VGND_c_1097_n N_VGND_c_1098_n N_VGND_c_1099_n N_VGND_c_1100_n
+ N_VGND_c_1101_n N_VGND_c_1102_n PM_SKY130_FD_SC_MS__NOR4B_4%VGND
cc_1 VNB N_D_N_c_149_n 0.101479f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.93
cc_2 VNB N_D_N_c_150_n 0.018845f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.185
cc_3 VNB N_D_N_c_151_n 0.0370874f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.085
cc_4 VNB N_A_47_88#_M1002_g 0.0230393f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.185
cc_5 VNB N_A_47_88#_M1003_g 0.0231678f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_6 VNB N_A_47_88#_M1011_g 0.0219865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_47_88#_M1028_g 0.0233014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_47_88#_c_188_n 0.016153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_47_88#_c_189_n 0.0877822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_47_88#_c_190_n 0.010652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_47_88#_c_191_n 0.00104905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_47_88#_c_192_n 0.00696627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_C_c_304_n 0.0162244f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.93
cc_14 VNB N_C_c_305_n 0.00881176f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.885
cc_15 VNB N_C_c_306_n 0.0172723f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_16 VNB N_C_c_307_n 0.01639f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.765
cc_17 VNB N_C_c_308_n 0.00902811f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.295
cc_18 VNB N_C_c_309_n 0.0162419f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.665
cc_19 VNB N_C_M1032_g 0.0215897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_C_c_311_n 0.00889195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB C 0.0042803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_C_c_313_n 0.0116767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_C_c_314_n 0.0924002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B_M1004_g 0.0280319f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_25 VNB N_B_M1008_g 0.024496f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_26 VNB N_B_M1009_g 0.0240482f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.765
cc_27 VNB N_B_M1019_g 0.0255763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB B 0.00547741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B_c_405_n 0.084315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_M1005_g 0.0255734f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.54
cc_31 VNB N_A_M1007_g 0.0224928f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_32 VNB N_A_M1015_g 0.0224928f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.765
cc_33 VNB N_A_M1029_g 0.0305461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB A 0.00266041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_c_499_n 0.0825172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_576_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_745_n 0.00253603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_Y_c_746_n 0.0034414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_Y_c_747_n 0.00223541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Y_c_748_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_Y_c_749_n 0.0105947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_Y_c_750_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_Y_c_751_n 0.00844257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_Y_c_752_n 0.0024006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_Y_c_753_n 0.0115474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_Y_c_754_n 0.00491298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_Y_c_755_n 0.00280455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_Y_c_756_n 0.00307912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_Y_c_757_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_Y_c_758_n 0.00408994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_Y_c_759_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_Y_c_760_n 0.0050343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_Y_c_761_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_Y_c_762_n 0.00324275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_Y_c_763_n 0.00231148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_Y_c_764_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_Y_c_765_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB Y 0.0122064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1077_n 0.00607168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1078_n 0.00509474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1079_n 0.0108774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1080_n 0.0119347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1081_n 0.00516528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1082_n 0.008436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1083_n 0.00269659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1084_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1085_n 0.0541576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1086_n 0.031535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1087_n 0.0170944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1088_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1089_n 0.0423352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1090_n 0.0187266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1091_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1092_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1093_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1094_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1095_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1096_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1097_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1098_n 0.0129835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1099_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1100_n 0.00682834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1101_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1102_n 0.528476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VPB N_D_N_c_149_n 0.0467396f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.93
cc_86 VPB N_D_N_M1012_g 0.028805f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_87 VPB N_D_N_M1013_g 0.0277343f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.54
cc_88 VPB N_D_N_c_151_n 0.0146866f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.085
cc_89 VPB N_A_47_88#_c_193_n 0.0229849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_47_88#_c_194_n 0.0183461f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.085
cc_91 VPB N_A_47_88#_c_195_n 0.0183461f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_47_88#_c_188_n 0.00630042f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_47_88#_c_189_n 0.0407083f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_47_88#_c_198_n 0.0181892f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_47_88#_c_199_n 0.00639286f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_47_88#_c_200_n 0.00184377f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_C_M1000_g 0.0217568f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_C_M1001_g 0.0210627f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_C_M1031_g 0.0207635f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.765
cc_100 VPB N_C_M1032_g 0.0250146f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB C 0.0102122f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_C_c_314_n 0.0119392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_B_M1014_g 0.0248261f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.54
cc_104 VPB N_B_M1016_g 0.0207967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_B_M1017_g 0.0202197f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_B_M1018_g 0.0208623f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB B 0.0139193f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_B_c_405_n 0.0181092f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_M1020_g 0.0202417f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_110 VPB N_A_M1021_g 0.020498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_M1023_g 0.0204973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_M1033_g 0.0285289f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB A 0.0110376f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_c_499_n 0.0123259f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_577_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_116 VPB N_VPWR_c_578_n 0.0462542f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_579_n 0.0206214f $X=-0.19 $Y=1.66 $X2=0.645 $Y2=1.765
cc_118 VPB N_VPWR_c_580_n 0.00554449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_581_n 0.00554449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_582_n 0.0199677f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_583_n 0.160986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_584_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_585_n 0.0180274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_576_n 0.104399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_587_n 0.00516749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_588_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_589_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_319_368#_c_680_n 0.0127902f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.085
cc_129 VPB N_A_319_368#_c_681_n 0.00240659f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.085
cc_130 VPB N_A_319_368#_c_682_n 0.00376758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_319_368#_c_683_n 0.00401291f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.765
cc_132 VPB N_A_319_368#_c_684_n 0.00203831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_319_368#_c_685_n 0.00316175f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_Y_c_767_n 0.00222771f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_Y_c_768_n 0.00265934f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_Y_c_769_n 0.00235306f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB Y 0.00430194f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_781_368#_c_946_n 0.00245644f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_139 VPB N_A_781_368#_c_947_n 0.016918f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_781_368#_c_948_n 0.00422885f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.765
cc_141 VPB N_A_781_368#_c_949_n 0.00328286f $X=-0.19 $Y=1.66 $X2=0.337 $Y2=1.765
cc_142 VPB N_A_781_368#_c_950_n 0.00213199f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_781_368#_c_951_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_1191_368#_c_1007_n 0.00232987f $X=-0.19 $Y=1.66 $X2=0.337
+ $Y2=1.765
cc_145 VPB N_A_1191_368#_c_1008_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_1191_368#_c_1009_n 0.0222704f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_1191_368#_c_1010_n 0.033959f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_1191_368#_c_1011_n 0.00966886f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 N_D_N_c_150_n N_A_47_88#_M1002_g 0.0178975f $X=0.995 $Y=1.185 $X2=0 $Y2=0
cc_150 N_D_N_c_149_n N_A_47_88#_c_189_n 0.0200161f $X=0.505 $Y=1.93 $X2=0 $Y2=0
cc_151 N_D_N_c_149_n N_A_47_88#_c_190_n 0.00519978f $X=0.505 $Y=1.93 $X2=0 $Y2=0
cc_152 N_D_N_c_151_n N_A_47_88#_c_190_n 0.0229928f $X=0.385 $Y=1.085 $X2=0 $Y2=0
cc_153 N_D_N_c_149_n N_A_47_88#_c_199_n 0.00160824f $X=0.505 $Y=1.93 $X2=0 $Y2=0
cc_154 N_D_N_M1012_g N_A_47_88#_c_199_n 0.0151088f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_155 N_D_N_M1013_g N_A_47_88#_c_199_n 0.0131455f $X=0.955 $Y=2.54 $X2=0 $Y2=0
cc_156 N_D_N_c_149_n N_A_47_88#_c_191_n 0.0108506f $X=0.505 $Y=1.93 $X2=0 $Y2=0
cc_157 N_D_N_c_150_n N_A_47_88#_c_191_n 0.005256f $X=0.995 $Y=1.185 $X2=0 $Y2=0
cc_158 N_D_N_c_151_n N_A_47_88#_c_191_n 0.0298646f $X=0.385 $Y=1.085 $X2=0 $Y2=0
cc_159 N_D_N_c_149_n N_A_47_88#_c_192_n 0.0247534f $X=0.505 $Y=1.93 $X2=0 $Y2=0
cc_160 N_D_N_c_149_n N_A_47_88#_c_200_n 0.0195581f $X=0.505 $Y=1.93 $X2=0 $Y2=0
cc_161 N_D_N_M1013_g N_A_47_88#_c_200_n 0.0101739f $X=0.955 $Y=2.54 $X2=0 $Y2=0
cc_162 N_D_N_c_151_n N_A_47_88#_c_200_n 0.0205445f $X=0.385 $Y=1.085 $X2=0 $Y2=0
cc_163 N_D_N_c_149_n N_A_47_88#_c_215_n 0.0100663f $X=0.505 $Y=1.93 $X2=0 $Y2=0
cc_164 N_D_N_c_151_n N_A_47_88#_c_215_n 0.0268332f $X=0.385 $Y=1.085 $X2=0 $Y2=0
cc_165 N_D_N_c_149_n N_VPWR_c_578_n 0.00112612f $X=0.505 $Y=1.93 $X2=0 $Y2=0
cc_166 N_D_N_M1012_g N_VPWR_c_578_n 0.00870081f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_167 N_D_N_c_151_n N_VPWR_c_578_n 0.0216458f $X=0.385 $Y=1.085 $X2=0 $Y2=0
cc_168 N_D_N_M1013_g N_VPWR_c_579_n 0.00841865f $X=0.955 $Y=2.54 $X2=0 $Y2=0
cc_169 N_D_N_M1012_g N_VPWR_c_582_n 0.005209f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_170 N_D_N_M1013_g N_VPWR_c_582_n 0.005209f $X=0.955 $Y=2.54 $X2=0 $Y2=0
cc_171 N_D_N_M1012_g N_VPWR_c_576_n 0.00986008f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_172 N_D_N_M1013_g N_VPWR_c_576_n 0.00986951f $X=0.955 $Y=2.54 $X2=0 $Y2=0
cc_173 N_D_N_c_149_n N_A_319_368#_c_680_n 0.00862776f $X=0.505 $Y=1.93 $X2=0
+ $Y2=0
cc_174 N_D_N_c_150_n N_VGND_c_1077_n 0.0170704f $X=0.995 $Y=1.185 $X2=0 $Y2=0
cc_175 N_D_N_c_150_n N_VGND_c_1086_n 0.00429299f $X=0.995 $Y=1.185 $X2=0 $Y2=0
cc_176 N_D_N_c_150_n N_VGND_c_1102_n 0.00852523f $X=0.995 $Y=1.185 $X2=0 $Y2=0
cc_177 N_A_47_88#_M1028_g N_C_c_304_n 0.011234f $X=2.88 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_178 N_A_47_88#_c_188_n N_C_c_305_n 0.00444043f $X=3.275 $Y=1.65 $X2=0 $Y2=0
cc_179 N_A_47_88#_c_189_n N_C_c_305_n 0.011234f $X=3.005 $Y=1.65 $X2=0 $Y2=0
cc_180 N_A_47_88#_c_198_n N_C_M1000_g 0.0213081f $X=3.365 $Y=1.725 $X2=0 $Y2=0
cc_181 N_A_47_88#_c_188_n C 5.33406e-19 $X=3.275 $Y=1.65 $X2=0 $Y2=0
cc_182 N_A_47_88#_c_188_n N_C_c_314_n 0.0213081f $X=3.275 $Y=1.65 $X2=0 $Y2=0
cc_183 N_A_47_88#_c_199_n N_VPWR_c_578_n 0.030311f $X=0.73 $Y=2.265 $X2=0 $Y2=0
cc_184 N_A_47_88#_c_193_n N_VPWR_c_579_n 8.7202e-19 $X=1.965 $Y=1.725 $X2=0
+ $Y2=0
cc_185 N_A_47_88#_c_189_n N_VPWR_c_579_n 5.29226e-19 $X=3.005 $Y=1.65 $X2=0
+ $Y2=0
cc_186 N_A_47_88#_c_199_n N_VPWR_c_579_n 0.0329775f $X=0.73 $Y=2.265 $X2=0 $Y2=0
cc_187 N_A_47_88#_c_192_n N_VPWR_c_579_n 0.0119664f $X=2.165 $Y=1.485 $X2=0
+ $Y2=0
cc_188 N_A_47_88#_c_199_n N_VPWR_c_582_n 0.0144623f $X=0.73 $Y=2.265 $X2=0 $Y2=0
cc_189 N_A_47_88#_c_193_n N_VPWR_c_583_n 0.00333926f $X=1.965 $Y=1.725 $X2=0
+ $Y2=0
cc_190 N_A_47_88#_c_194_n N_VPWR_c_583_n 0.00333926f $X=2.415 $Y=1.725 $X2=0
+ $Y2=0
cc_191 N_A_47_88#_c_195_n N_VPWR_c_583_n 0.00333926f $X=2.915 $Y=1.725 $X2=0
+ $Y2=0
cc_192 N_A_47_88#_c_198_n N_VPWR_c_583_n 0.00333926f $X=3.365 $Y=1.725 $X2=0
+ $Y2=0
cc_193 N_A_47_88#_c_193_n N_VPWR_c_576_n 0.0042782f $X=1.965 $Y=1.725 $X2=0
+ $Y2=0
cc_194 N_A_47_88#_c_194_n N_VPWR_c_576_n 0.00423176f $X=2.415 $Y=1.725 $X2=0
+ $Y2=0
cc_195 N_A_47_88#_c_195_n N_VPWR_c_576_n 0.00423176f $X=2.915 $Y=1.725 $X2=0
+ $Y2=0
cc_196 N_A_47_88#_c_198_n N_VPWR_c_576_n 0.00422798f $X=3.365 $Y=1.725 $X2=0
+ $Y2=0
cc_197 N_A_47_88#_c_199_n N_VPWR_c_576_n 0.0118344f $X=0.73 $Y=2.265 $X2=0 $Y2=0
cc_198 N_A_47_88#_c_193_n N_A_319_368#_c_680_n 0.00147281f $X=1.965 $Y=1.725
+ $X2=0 $Y2=0
cc_199 N_A_47_88#_c_189_n N_A_319_368#_c_680_n 0.00680866f $X=3.005 $Y=1.65
+ $X2=0 $Y2=0
cc_200 N_A_47_88#_c_192_n N_A_319_368#_c_680_n 0.0209125f $X=2.165 $Y=1.485
+ $X2=0 $Y2=0
cc_201 N_A_47_88#_c_193_n N_A_319_368#_c_681_n 0.0149445f $X=1.965 $Y=1.725
+ $X2=0 $Y2=0
cc_202 N_A_47_88#_c_194_n N_A_319_368#_c_681_n 0.0142213f $X=2.415 $Y=1.725
+ $X2=0 $Y2=0
cc_203 N_A_47_88#_c_195_n N_A_319_368#_c_683_n 0.0142213f $X=2.915 $Y=1.725
+ $X2=0 $Y2=0
cc_204 N_A_47_88#_c_198_n N_A_319_368#_c_683_n 0.0139961f $X=3.365 $Y=1.725
+ $X2=0 $Y2=0
cc_205 N_A_47_88#_M1002_g N_Y_c_745_n 0.00335659f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A_47_88#_M1003_g N_Y_c_745_n 4.79304e-19 $X=1.95 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A_47_88#_M1003_g N_Y_c_746_n 0.013154f $X=1.95 $Y=0.74 $X2=0 $Y2=0
cc_208 N_A_47_88#_M1011_g N_Y_c_746_n 0.0144352f $X=2.45 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A_47_88#_c_189_n N_Y_c_746_n 0.00421375f $X=3.005 $Y=1.65 $X2=0 $Y2=0
cc_210 N_A_47_88#_c_192_n N_Y_c_746_n 0.0377337f $X=2.165 $Y=1.485 $X2=0 $Y2=0
cc_211 N_A_47_88#_M1002_g N_Y_c_747_n 0.00151697f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A_47_88#_c_189_n N_Y_c_747_n 0.00436753f $X=3.005 $Y=1.65 $X2=0 $Y2=0
cc_213 N_A_47_88#_c_192_n N_Y_c_747_n 0.0210847f $X=2.165 $Y=1.485 $X2=0 $Y2=0
cc_214 N_A_47_88#_c_193_n N_Y_c_767_n 0.00279295f $X=1.965 $Y=1.725 $X2=0 $Y2=0
cc_215 N_A_47_88#_c_194_n N_Y_c_767_n 0.00146862f $X=2.415 $Y=1.725 $X2=0 $Y2=0
cc_216 N_A_47_88#_c_189_n N_Y_c_767_n 0.00239121f $X=3.005 $Y=1.65 $X2=0 $Y2=0
cc_217 N_A_47_88#_c_192_n N_Y_c_767_n 0.0255666f $X=2.165 $Y=1.485 $X2=0 $Y2=0
cc_218 N_A_47_88#_c_193_n N_Y_c_784_n 0.00971651f $X=1.965 $Y=1.725 $X2=0 $Y2=0
cc_219 N_A_47_88#_c_194_n N_Y_c_784_n 0.0102924f $X=2.415 $Y=1.725 $X2=0 $Y2=0
cc_220 N_A_47_88#_c_195_n N_Y_c_784_n 5.83379e-19 $X=2.915 $Y=1.725 $X2=0 $Y2=0
cc_221 N_A_47_88#_c_194_n N_Y_c_768_n 0.0152815f $X=2.415 $Y=1.725 $X2=0 $Y2=0
cc_222 N_A_47_88#_c_195_n N_Y_c_768_n 0.0148147f $X=2.915 $Y=1.725 $X2=0 $Y2=0
cc_223 N_A_47_88#_c_189_n N_Y_c_768_n 0.00402675f $X=3.005 $Y=1.65 $X2=0 $Y2=0
cc_224 N_A_47_88#_M1003_g N_Y_c_748_n 9.70813e-19 $X=1.95 $Y=0.74 $X2=0 $Y2=0
cc_225 N_A_47_88#_M1011_g N_Y_c_748_n 0.00933152f $X=2.45 $Y=0.74 $X2=0 $Y2=0
cc_226 N_A_47_88#_M1028_g N_Y_c_748_n 0.00767492f $X=2.88 $Y=0.74 $X2=0 $Y2=0
cc_227 N_A_47_88#_M1028_g N_Y_c_749_n 0.00612947f $X=2.88 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A_47_88#_c_189_n N_Y_c_749_n 0.0210533f $X=3.005 $Y=1.65 $X2=0 $Y2=0
cc_229 N_A_47_88#_c_195_n N_Y_c_795_n 0.00766694f $X=2.915 $Y=1.725 $X2=0 $Y2=0
cc_230 N_A_47_88#_c_198_n N_Y_c_795_n 0.00883449f $X=3.365 $Y=1.725 $X2=0 $Y2=0
cc_231 N_A_47_88#_c_198_n N_Y_c_797_n 0.0147998f $X=3.365 $Y=1.725 $X2=0 $Y2=0
cc_232 N_A_47_88#_M1028_g N_Y_c_750_n 6.91376e-19 $X=2.88 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A_47_88#_M1003_g N_Y_c_799_n 8.81603e-19 $X=1.95 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A_47_88#_M1011_g N_Y_c_799_n 0.00666364f $X=2.45 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A_47_88#_M1028_g N_Y_c_799_n 0.00762747f $X=2.88 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A_47_88#_c_189_n N_Y_c_799_n 0.0154748f $X=3.005 $Y=1.65 $X2=0 $Y2=0
cc_237 N_A_47_88#_c_192_n N_Y_c_799_n 0.0118939f $X=2.165 $Y=1.485 $X2=0 $Y2=0
cc_238 N_A_47_88#_c_194_n N_Y_c_769_n 6.60808e-19 $X=2.415 $Y=1.725 $X2=0 $Y2=0
cc_239 N_A_47_88#_c_195_n N_Y_c_769_n 0.00426294f $X=2.915 $Y=1.725 $X2=0 $Y2=0
cc_240 N_A_47_88#_c_188_n N_Y_c_769_n 0.00226086f $X=3.275 $Y=1.65 $X2=0 $Y2=0
cc_241 N_A_47_88#_c_198_n N_Y_c_769_n 0.00411963f $X=3.365 $Y=1.725 $X2=0 $Y2=0
cc_242 N_A_47_88#_c_189_n N_Y_c_762_n 2.78242e-19 $X=3.005 $Y=1.65 $X2=0 $Y2=0
cc_243 N_A_47_88#_M1002_g N_VGND_c_1077_n 0.0136496f $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A_47_88#_M1003_g N_VGND_c_1077_n 5.37974e-19 $X=1.95 $Y=0.74 $X2=0
+ $Y2=0
cc_245 N_A_47_88#_c_189_n N_VGND_c_1077_n 0.00108047f $X=3.005 $Y=1.65 $X2=0
+ $Y2=0
cc_246 N_A_47_88#_c_191_n N_VGND_c_1077_n 0.0149733f $X=0.805 $Y=1.32 $X2=0
+ $Y2=0
cc_247 N_A_47_88#_c_192_n N_VGND_c_1077_n 0.0263407f $X=2.165 $Y=1.485 $X2=0
+ $Y2=0
cc_248 N_A_47_88#_M1002_g N_VGND_c_1078_n 4.4638e-19 $X=1.44 $Y=0.74 $X2=0 $Y2=0
cc_249 N_A_47_88#_M1003_g N_VGND_c_1078_n 0.00983095f $X=1.95 $Y=0.74 $X2=0
+ $Y2=0
cc_250 N_A_47_88#_M1011_g N_VGND_c_1078_n 0.00406778f $X=2.45 $Y=0.74 $X2=0
+ $Y2=0
cc_251 N_A_47_88#_M1028_g N_VGND_c_1079_n 0.00666821f $X=2.88 $Y=0.74 $X2=0
+ $Y2=0
cc_252 N_A_47_88#_c_190_n N_VGND_c_1086_n 0.0145959f $X=0.72 $Y=0.585 $X2=0
+ $Y2=0
cc_253 N_A_47_88#_c_293_p N_VGND_c_1086_n 0.00530359f $X=0.805 $Y=0.75 $X2=0
+ $Y2=0
cc_254 N_A_47_88#_M1002_g N_VGND_c_1087_n 0.00383152f $X=1.44 $Y=0.74 $X2=0
+ $Y2=0
cc_255 N_A_47_88#_M1003_g N_VGND_c_1087_n 0.00383152f $X=1.95 $Y=0.74 $X2=0
+ $Y2=0
cc_256 N_A_47_88#_M1011_g N_VGND_c_1088_n 0.00434272f $X=2.45 $Y=0.74 $X2=0
+ $Y2=0
cc_257 N_A_47_88#_M1028_g N_VGND_c_1088_n 0.00434272f $X=2.88 $Y=0.74 $X2=0
+ $Y2=0
cc_258 N_A_47_88#_M1002_g N_VGND_c_1102_n 0.00758285f $X=1.44 $Y=0.74 $X2=0
+ $Y2=0
cc_259 N_A_47_88#_M1003_g N_VGND_c_1102_n 0.00758285f $X=1.95 $Y=0.74 $X2=0
+ $Y2=0
cc_260 N_A_47_88#_M1011_g N_VGND_c_1102_n 0.00820718f $X=2.45 $Y=0.74 $X2=0
+ $Y2=0
cc_261 N_A_47_88#_M1028_g N_VGND_c_1102_n 0.00821312f $X=2.88 $Y=0.74 $X2=0
+ $Y2=0
cc_262 N_A_47_88#_c_190_n N_VGND_c_1102_n 0.0152957f $X=0.72 $Y=0.585 $X2=0
+ $Y2=0
cc_263 N_A_47_88#_c_293_p N_VGND_c_1102_n 0.00600684f $X=0.805 $Y=0.75 $X2=0
+ $Y2=0
cc_264 N_C_c_311_n N_B_M1004_g 0.00222113f $X=5.307 $Y=1.26 $X2=0 $Y2=0
cc_265 N_C_M1032_g N_B_c_405_n 0.00222113f $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_266 N_C_M1000_g N_VPWR_c_583_n 0.00517089f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_267 N_C_M1001_g N_VPWR_c_583_n 0.00335119f $X=4.315 $Y=2.4 $X2=0 $Y2=0
cc_268 N_C_M1031_g N_VPWR_c_583_n 0.00335143f $X=4.84 $Y=2.4 $X2=0 $Y2=0
cc_269 N_C_M1032_g N_VPWR_c_583_n 0.00335119f $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_270 N_C_M1000_g N_VPWR_c_576_n 0.00534445f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_271 N_C_M1001_g N_VPWR_c_576_n 0.0042298f $X=4.315 $Y=2.4 $X2=0 $Y2=0
cc_272 N_C_M1031_g N_VPWR_c_576_n 0.00419108f $X=4.84 $Y=2.4 $X2=0 $Y2=0
cc_273 N_C_M1032_g N_VPWR_c_576_n 0.00427159f $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_274 N_C_M1000_g N_A_319_368#_c_683_n 0.00335819f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_275 N_C_M1000_g N_A_319_368#_c_695_n 9.22099e-19 $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_276 N_C_M1000_g N_A_319_368#_c_696_n 0.00628213f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_277 N_C_M1001_g N_A_319_368#_c_696_n 3.52569e-19 $X=4.315 $Y=2.4 $X2=0 $Y2=0
cc_278 N_C_M1000_g N_A_319_368#_c_698_n 0.0102593f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_279 N_C_M1001_g N_A_319_368#_c_698_n 0.0114298f $X=4.315 $Y=2.4 $X2=0 $Y2=0
cc_280 N_C_M1031_g N_A_319_368#_c_700_n 0.00494786f $X=4.84 $Y=2.4 $X2=0 $Y2=0
cc_281 N_C_M1032_g N_A_319_368#_c_700_n 6.4049e-19 $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_282 N_C_M1031_g N_A_319_368#_c_702_n 0.011157f $X=4.84 $Y=2.4 $X2=0 $Y2=0
cc_283 N_C_M1032_g N_A_319_368#_c_702_n 0.0112357f $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_284 N_C_c_304_n N_Y_c_748_n 4.05063e-19 $X=3.45 $Y=1.185 $X2=0 $Y2=0
cc_285 N_C_c_305_n N_Y_c_749_n 0.00783639f $X=3.525 $Y=1.26 $X2=0 $Y2=0
cc_286 N_C_c_314_n N_Y_c_749_n 5.43413e-19 $X=4.93 $Y=1.432 $X2=0 $Y2=0
cc_287 N_C_c_305_n N_Y_c_797_n 8.66207e-19 $X=3.525 $Y=1.26 $X2=0 $Y2=0
cc_288 N_C_M1000_g N_Y_c_797_n 0.0171336f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_289 N_C_M1001_g N_Y_c_797_n 0.0126077f $X=4.315 $Y=2.4 $X2=0 $Y2=0
cc_290 N_C_M1031_g N_Y_c_797_n 0.0121477f $X=4.84 $Y=2.4 $X2=0 $Y2=0
cc_291 N_C_M1032_g N_Y_c_797_n 0.0184794f $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_292 C N_Y_c_797_n 0.0861559f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_293 N_C_c_314_n N_Y_c_797_n 0.00165024f $X=4.93 $Y=1.432 $X2=0 $Y2=0
cc_294 N_C_c_304_n N_Y_c_750_n 0.00775604f $X=3.45 $Y=1.185 $X2=0 $Y2=0
cc_295 N_C_c_306_n N_Y_c_750_n 3.97481e-19 $X=3.88 $Y=1.185 $X2=0 $Y2=0
cc_296 N_C_c_306_n N_Y_c_751_n 0.0181545f $X=3.88 $Y=1.185 $X2=0 $Y2=0
cc_297 N_C_c_307_n N_Y_c_751_n 0.0131906f $X=4.855 $Y=1.185 $X2=0 $Y2=0
cc_298 C N_Y_c_751_n 0.0949583f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_299 N_C_c_314_n N_Y_c_751_n 0.0200647f $X=4.93 $Y=1.432 $X2=0 $Y2=0
cc_300 N_C_c_307_n N_Y_c_752_n 0.0138478f $X=4.855 $Y=1.185 $X2=0 $Y2=0
cc_301 N_C_c_309_n N_Y_c_752_n 0.0138478f $X=5.285 $Y=1.185 $X2=0 $Y2=0
cc_302 N_C_c_307_n N_Y_c_754_n 0.00161307f $X=4.855 $Y=1.185 $X2=0 $Y2=0
cc_303 N_C_c_308_n N_Y_c_754_n 0.00233369f $X=5.21 $Y=1.26 $X2=0 $Y2=0
cc_304 N_C_c_309_n N_Y_c_754_n 0.0195028f $X=5.285 $Y=1.185 $X2=0 $Y2=0
cc_305 N_C_c_311_n N_Y_c_754_n 0.00223761f $X=5.307 $Y=1.26 $X2=0 $Y2=0
cc_306 N_C_c_305_n N_Y_c_799_n 4.2021e-19 $X=3.525 $Y=1.26 $X2=0 $Y2=0
cc_307 N_C_M1000_g N_Y_c_769_n 0.00158489f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_308 N_C_c_304_n N_Y_c_762_n 0.00300516f $X=3.45 $Y=1.185 $X2=0 $Y2=0
cc_309 N_C_c_305_n N_Y_c_762_n 0.00296331f $X=3.525 $Y=1.26 $X2=0 $Y2=0
cc_310 N_C_c_306_n N_Y_c_762_n 2.86737e-19 $X=3.88 $Y=1.185 $X2=0 $Y2=0
cc_311 C N_Y_c_762_n 0.00931227f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_312 N_C_c_313_n N_Y_c_762_n 0.00857906f $X=3.725 $Y=1.432 $X2=0 $Y2=0
cc_313 N_C_c_314_n N_Y_c_762_n 0.0130569f $X=4.93 $Y=1.432 $X2=0 $Y2=0
cc_314 N_C_c_311_n Y 0.018562f $X=5.307 $Y=1.26 $X2=0 $Y2=0
cc_315 C Y 0.0281249f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_316 N_C_M1001_g N_A_781_368#_c_946_n 0.00934879f $X=4.315 $Y=2.4 $X2=0 $Y2=0
cc_317 N_C_M1031_g N_A_781_368#_c_946_n 0.0105329f $X=4.84 $Y=2.4 $X2=0 $Y2=0
cc_318 N_C_M1032_g N_A_781_368#_c_947_n 0.0111722f $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_319 N_C_M1000_g N_A_781_368#_c_949_n 0.00100515f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_320 N_C_M1001_g N_A_781_368#_c_949_n 0.00740307f $X=4.315 $Y=2.4 $X2=0 $Y2=0
cc_321 N_C_M1031_g N_A_781_368#_c_949_n 6.70462e-19 $X=4.84 $Y=2.4 $X2=0 $Y2=0
cc_322 N_C_M1001_g N_A_781_368#_c_950_n 6.397e-19 $X=4.315 $Y=2.4 $X2=0 $Y2=0
cc_323 N_C_M1031_g N_A_781_368#_c_950_n 0.00682065f $X=4.84 $Y=2.4 $X2=0 $Y2=0
cc_324 N_C_M1032_g N_A_781_368#_c_950_n 0.0151184f $X=5.315 $Y=2.4 $X2=0 $Y2=0
cc_325 N_C_M1032_g N_A_1191_368#_c_1011_n 0.00875054f $X=5.315 $Y=2.4 $X2=0
+ $Y2=0
cc_326 N_C_c_304_n N_VGND_c_1079_n 0.00657876f $X=3.45 $Y=1.185 $X2=0 $Y2=0
cc_327 N_C_c_309_n N_VGND_c_1080_n 0.0060502f $X=5.285 $Y=1.185 $X2=0 $Y2=0
cc_328 N_C_c_304_n N_VGND_c_1089_n 0.00485667f $X=3.45 $Y=1.185 $X2=0 $Y2=0
cc_329 N_C_c_306_n N_VGND_c_1089_n 0.0175569f $X=3.88 $Y=1.185 $X2=0 $Y2=0
cc_330 N_C_c_307_n N_VGND_c_1089_n 0.00607183f $X=4.855 $Y=1.185 $X2=0 $Y2=0
cc_331 N_C_c_307_n N_VGND_c_1090_n 0.00434272f $X=4.855 $Y=1.185 $X2=0 $Y2=0
cc_332 N_C_c_309_n N_VGND_c_1090_n 0.00434272f $X=5.285 $Y=1.185 $X2=0 $Y2=0
cc_333 N_C_c_304_n N_VGND_c_1102_n 0.00821312f $X=3.45 $Y=1.185 $X2=0 $Y2=0
cc_334 N_C_c_306_n N_VGND_c_1102_n 0.0075754f $X=3.88 $Y=1.185 $X2=0 $Y2=0
cc_335 N_C_c_307_n N_VGND_c_1102_n 0.00825059f $X=4.855 $Y=1.185 $X2=0 $Y2=0
cc_336 N_C_c_309_n N_VGND_c_1102_n 0.00825059f $X=5.285 $Y=1.185 $X2=0 $Y2=0
cc_337 N_B_M1018_g N_A_M1020_g 0.0113899f $X=7.775 $Y=2.4 $X2=0 $Y2=0
cc_338 N_B_M1019_g N_A_M1005_g 0.0242687f $X=7.63 $Y=0.74 $X2=0 $Y2=0
cc_339 N_B_M1018_g A 0.00345577f $X=7.775 $Y=2.4 $X2=0 $Y2=0
cc_340 B A 0.0269711f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_341 N_B_c_405_n A 0.0118953f $X=7.775 $Y=1.515 $X2=0 $Y2=0
cc_342 N_B_c_405_n N_A_c_499_n 0.0181186f $X=7.775 $Y=1.515 $X2=0 $Y2=0
cc_343 N_B_M1018_g N_VPWR_c_580_n 5.51283e-19 $X=7.775 $Y=2.4 $X2=0 $Y2=0
cc_344 N_B_M1014_g N_VPWR_c_583_n 0.00333926f $X=6.325 $Y=2.4 $X2=0 $Y2=0
cc_345 N_B_M1016_g N_VPWR_c_583_n 0.00333896f $X=6.825 $Y=2.4 $X2=0 $Y2=0
cc_346 N_B_M1017_g N_VPWR_c_583_n 0.00333926f $X=7.325 $Y=2.4 $X2=0 $Y2=0
cc_347 N_B_M1018_g N_VPWR_c_583_n 0.00517089f $X=7.775 $Y=2.4 $X2=0 $Y2=0
cc_348 N_B_M1014_g N_VPWR_c_576_n 0.00428309f $X=6.325 $Y=2.4 $X2=0 $Y2=0
cc_349 N_B_M1016_g N_VPWR_c_576_n 0.00423662f $X=6.825 $Y=2.4 $X2=0 $Y2=0
cc_350 N_B_M1017_g N_VPWR_c_576_n 0.00423176f $X=7.325 $Y=2.4 $X2=0 $Y2=0
cc_351 N_B_M1018_g N_VPWR_c_576_n 0.00978686f $X=7.775 $Y=2.4 $X2=0 $Y2=0
cc_352 N_B_M1014_g N_A_319_368#_c_685_n 6.69392e-19 $X=6.325 $Y=2.4 $X2=0 $Y2=0
cc_353 N_B_M1004_g N_Y_c_753_n 0.0131906f $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_354 B N_Y_c_753_n 0.0285229f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_355 N_B_M1004_g N_Y_c_755_n 0.0137366f $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_356 N_B_M1008_g N_Y_c_755_n 0.00350341f $X=6.7 $Y=0.74 $X2=0 $Y2=0
cc_357 N_B_M1008_g N_Y_c_756_n 0.0151601f $X=6.7 $Y=0.74 $X2=0 $Y2=0
cc_358 N_B_M1009_g N_Y_c_756_n 0.0115433f $X=7.2 $Y=0.74 $X2=0 $Y2=0
cc_359 B N_Y_c_756_n 0.0502964f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_360 N_B_c_405_n N_Y_c_756_n 0.00436308f $X=7.775 $Y=1.515 $X2=0 $Y2=0
cc_361 N_B_M1008_g N_Y_c_757_n 7.24002e-19 $X=6.7 $Y=0.74 $X2=0 $Y2=0
cc_362 N_B_M1009_g N_Y_c_757_n 0.00991175f $X=7.2 $Y=0.74 $X2=0 $Y2=0
cc_363 N_B_M1019_g N_Y_c_757_n 0.0101239f $X=7.63 $Y=0.74 $X2=0 $Y2=0
cc_364 N_B_M1019_g N_Y_c_758_n 0.0156506f $X=7.63 $Y=0.74 $X2=0 $Y2=0
cc_365 N_B_c_405_n N_Y_c_758_n 0.00573225f $X=7.775 $Y=1.515 $X2=0 $Y2=0
cc_366 N_B_M1019_g N_Y_c_759_n 0.00100994f $X=7.63 $Y=0.74 $X2=0 $Y2=0
cc_367 N_B_M1004_g N_Y_c_763_n 0.00173883f $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_368 B N_Y_c_763_n 0.0282341f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_369 N_B_c_405_n N_Y_c_763_n 0.00451245f $X=7.775 $Y=1.515 $X2=0 $Y2=0
cc_370 N_B_M1009_g N_Y_c_764_n 0.00157732f $X=7.2 $Y=0.74 $X2=0 $Y2=0
cc_371 N_B_M1019_g N_Y_c_764_n 0.00243516f $X=7.63 $Y=0.74 $X2=0 $Y2=0
cc_372 B N_Y_c_764_n 0.0260877f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_373 N_B_c_405_n N_Y_c_764_n 0.00272398f $X=7.775 $Y=1.515 $X2=0 $Y2=0
cc_374 N_B_M1004_g Y 0.00303248f $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_375 N_B_M1014_g Y 0.00305482f $X=6.325 $Y=2.4 $X2=0 $Y2=0
cc_376 B Y 0.0281718f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_377 N_B_c_405_n Y 8.72526e-19 $X=7.775 $Y=1.515 $X2=0 $Y2=0
cc_378 N_B_M1014_g N_A_781_368#_c_947_n 0.0163444f $X=6.325 $Y=2.4 $X2=0 $Y2=0
cc_379 N_B_M1016_g N_A_781_368#_c_962_n 0.00877172f $X=6.825 $Y=2.4 $X2=0 $Y2=0
cc_380 N_B_M1017_g N_A_781_368#_c_962_n 8.6734e-19 $X=7.325 $Y=2.4 $X2=0 $Y2=0
cc_381 N_B_M1016_g N_A_781_368#_c_948_n 0.0119307f $X=6.825 $Y=2.4 $X2=0 $Y2=0
cc_382 N_B_M1017_g N_A_781_368#_c_948_n 0.0143183f $X=7.325 $Y=2.4 $X2=0 $Y2=0
cc_383 N_B_M1018_g N_A_781_368#_c_948_n 0.00414503f $X=7.775 $Y=2.4 $X2=0 $Y2=0
cc_384 N_B_M1018_g N_A_781_368#_c_967_n 0.00727215f $X=7.775 $Y=2.4 $X2=0 $Y2=0
cc_385 N_B_M1016_g N_A_781_368#_c_951_n 0.00214324f $X=6.825 $Y=2.4 $X2=0 $Y2=0
cc_386 N_B_M1014_g N_A_1191_368#_c_1013_n 0.0132272f $X=6.325 $Y=2.4 $X2=0 $Y2=0
cc_387 N_B_M1016_g N_A_1191_368#_c_1013_n 0.0145524f $X=6.825 $Y=2.4 $X2=0 $Y2=0
cc_388 B N_A_1191_368#_c_1013_n 0.046225f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_389 N_B_c_405_n N_A_1191_368#_c_1013_n 7.55656e-19 $X=7.775 $Y=1.515 $X2=0
+ $Y2=0
cc_390 N_B_M1017_g N_A_1191_368#_c_1017_n 0.010699f $X=7.325 $Y=2.4 $X2=0 $Y2=0
cc_391 N_B_M1018_g N_A_1191_368#_c_1017_n 4.41999e-19 $X=7.775 $Y=2.4 $X2=0
+ $Y2=0
cc_392 N_B_M1017_g N_A_1191_368#_c_1019_n 0.012931f $X=7.325 $Y=2.4 $X2=0 $Y2=0
cc_393 N_B_M1018_g N_A_1191_368#_c_1019_n 0.0177447f $X=7.775 $Y=2.4 $X2=0 $Y2=0
cc_394 B N_A_1191_368#_c_1019_n 0.0199917f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_395 N_B_c_405_n N_A_1191_368#_c_1019_n 0.00176071f $X=7.775 $Y=1.515 $X2=0
+ $Y2=0
cc_396 N_B_M1018_g N_A_1191_368#_c_1007_n 2.20696e-19 $X=7.775 $Y=2.4 $X2=0
+ $Y2=0
cc_397 N_B_M1014_g N_A_1191_368#_c_1011_n 0.0127636f $X=6.325 $Y=2.4 $X2=0 $Y2=0
cc_398 N_B_M1016_g N_A_1191_368#_c_1011_n 4.54422e-19 $X=6.825 $Y=2.4 $X2=0
+ $Y2=0
cc_399 B N_A_1191_368#_c_1011_n 0.0263957f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_400 N_B_c_405_n N_A_1191_368#_c_1011_n 5.27311e-19 $X=7.775 $Y=1.515 $X2=0
+ $Y2=0
cc_401 N_B_M1017_g N_A_1191_368#_c_1028_n 8.84614e-19 $X=7.325 $Y=2.4 $X2=0
+ $Y2=0
cc_402 B N_A_1191_368#_c_1028_n 0.0246996f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_403 N_B_c_405_n N_A_1191_368#_c_1028_n 8.55208e-19 $X=7.775 $Y=1.515 $X2=0
+ $Y2=0
cc_404 N_B_M1004_g N_VGND_c_1080_n 0.0060502f $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_405 N_B_M1004_g N_VGND_c_1081_n 4.90868e-19 $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_406 N_B_M1008_g N_VGND_c_1081_n 0.0101619f $X=6.7 $Y=0.74 $X2=0 $Y2=0
cc_407 N_B_M1009_g N_VGND_c_1081_n 0.00414597f $X=7.2 $Y=0.74 $X2=0 $Y2=0
cc_408 N_B_M1019_g N_VGND_c_1082_n 0.00481771f $X=7.63 $Y=0.74 $X2=0 $Y2=0
cc_409 N_B_M1004_g N_VGND_c_1091_n 0.00434272f $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_410 N_B_M1008_g N_VGND_c_1091_n 0.00383152f $X=6.7 $Y=0.74 $X2=0 $Y2=0
cc_411 N_B_M1009_g N_VGND_c_1092_n 0.00434272f $X=7.2 $Y=0.74 $X2=0 $Y2=0
cc_412 N_B_M1019_g N_VGND_c_1092_n 0.00434272f $X=7.63 $Y=0.74 $X2=0 $Y2=0
cc_413 N_B_M1004_g N_VGND_c_1102_n 0.00825717f $X=6.2 $Y=0.74 $X2=0 $Y2=0
cc_414 N_B_M1008_g N_VGND_c_1102_n 0.00758198f $X=6.7 $Y=0.74 $X2=0 $Y2=0
cc_415 N_B_M1009_g N_VGND_c_1102_n 0.00820718f $X=7.2 $Y=0.74 $X2=0 $Y2=0
cc_416 N_B_M1019_g N_VGND_c_1102_n 0.00821489f $X=7.63 $Y=0.74 $X2=0 $Y2=0
cc_417 N_A_M1020_g N_VPWR_c_580_n 0.0119688f $X=8.225 $Y=2.4 $X2=0 $Y2=0
cc_418 N_A_M1021_g N_VPWR_c_580_n 0.002979f $X=8.675 $Y=2.4 $X2=0 $Y2=0
cc_419 N_A_M1023_g N_VPWR_c_581_n 0.002979f $X=9.125 $Y=2.4 $X2=0 $Y2=0
cc_420 N_A_M1033_g N_VPWR_c_581_n 0.0153844f $X=9.575 $Y=2.4 $X2=0 $Y2=0
cc_421 N_A_M1020_g N_VPWR_c_583_n 0.00460063f $X=8.225 $Y=2.4 $X2=0 $Y2=0
cc_422 N_A_M1021_g N_VPWR_c_584_n 0.005209f $X=8.675 $Y=2.4 $X2=0 $Y2=0
cc_423 N_A_M1023_g N_VPWR_c_584_n 0.005209f $X=9.125 $Y=2.4 $X2=0 $Y2=0
cc_424 N_A_M1033_g N_VPWR_c_585_n 0.00460063f $X=9.575 $Y=2.4 $X2=0 $Y2=0
cc_425 N_A_M1020_g N_VPWR_c_576_n 0.00908665f $X=8.225 $Y=2.4 $X2=0 $Y2=0
cc_426 N_A_M1021_g N_VPWR_c_576_n 0.00982266f $X=8.675 $Y=2.4 $X2=0 $Y2=0
cc_427 N_A_M1023_g N_VPWR_c_576_n 0.00982266f $X=9.125 $Y=2.4 $X2=0 $Y2=0
cc_428 N_A_M1033_g N_VPWR_c_576_n 0.00912296f $X=9.575 $Y=2.4 $X2=0 $Y2=0
cc_429 N_A_M1005_g N_Y_c_757_n 0.00100644f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_430 N_A_M1005_g N_Y_c_758_n 0.0118978f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_431 A N_Y_c_758_n 0.0367696f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_432 N_A_M1005_g N_Y_c_759_n 0.00977465f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_433 N_A_M1007_g N_Y_c_759_n 3.97481e-19 $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_434 N_A_M1007_g N_Y_c_760_n 0.0131257f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_435 N_A_M1015_g N_Y_c_760_n 0.0131257f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_436 N_A_M1029_g N_Y_c_760_n 0.00483035f $X=9.515 $Y=0.74 $X2=0 $Y2=0
cc_437 A N_Y_c_760_n 0.0730968f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_438 N_A_c_499_n N_Y_c_760_n 0.00492645f $X=9.515 $Y=1.515 $X2=0 $Y2=0
cc_439 N_A_M1015_g N_Y_c_761_n 3.97481e-19 $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_440 N_A_M1029_g N_Y_c_761_n 0.0079794f $X=9.515 $Y=0.74 $X2=0 $Y2=0
cc_441 N_A_M1005_g N_Y_c_765_n 0.00157732f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_442 A N_Y_c_765_n 0.0213626f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_443 N_A_c_499_n N_Y_c_765_n 0.00238873f $X=9.515 $Y=1.515 $X2=0 $Y2=0
cc_444 N_A_M1020_g N_A_781_368#_c_948_n 2.96504e-19 $X=8.225 $Y=2.4 $X2=0 $Y2=0
cc_445 A N_A_1191_368#_c_1019_n 0.00521059f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_446 N_A_M1020_g N_A_1191_368#_c_1007_n 2.21024e-19 $X=8.225 $Y=2.4 $X2=0
+ $Y2=0
cc_447 N_A_M1020_g N_A_1191_368#_c_1033_n 0.0142562f $X=8.225 $Y=2.4 $X2=0 $Y2=0
cc_448 N_A_M1021_g N_A_1191_368#_c_1033_n 0.012931f $X=8.675 $Y=2.4 $X2=0 $Y2=0
cc_449 A N_A_1191_368#_c_1033_n 0.0422425f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_450 N_A_c_499_n N_A_1191_368#_c_1033_n 4.90415e-19 $X=9.515 $Y=1.515 $X2=0
+ $Y2=0
cc_451 N_A_M1020_g N_A_1191_368#_c_1008_n 6.6858e-19 $X=8.225 $Y=2.4 $X2=0 $Y2=0
cc_452 N_A_M1021_g N_A_1191_368#_c_1008_n 0.0122399f $X=8.675 $Y=2.4 $X2=0 $Y2=0
cc_453 N_A_M1023_g N_A_1191_368#_c_1008_n 0.0123116f $X=9.125 $Y=2.4 $X2=0 $Y2=0
cc_454 N_A_M1033_g N_A_1191_368#_c_1008_n 6.74232e-19 $X=9.575 $Y=2.4 $X2=0
+ $Y2=0
cc_455 N_A_M1023_g N_A_1191_368#_c_1041_n 0.012931f $X=9.125 $Y=2.4 $X2=0 $Y2=0
cc_456 N_A_M1033_g N_A_1191_368#_c_1041_n 0.0195925f $X=9.575 $Y=2.4 $X2=0 $Y2=0
cc_457 A N_A_1191_368#_c_1041_n 0.0278429f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_458 N_A_c_499_n N_A_1191_368#_c_1041_n 4.87593e-19 $X=9.515 $Y=1.515 $X2=0
+ $Y2=0
cc_459 N_A_M1033_g N_A_1191_368#_c_1009_n 8.13654e-19 $X=9.575 $Y=2.4 $X2=0
+ $Y2=0
cc_460 N_A_M1033_g N_A_1191_368#_c_1010_n 0.00147311f $X=9.575 $Y=2.4 $X2=0
+ $Y2=0
cc_461 A N_A_1191_368#_c_1047_n 0.0170102f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_462 N_A_M1021_g N_A_1191_368#_c_1048_n 8.84614e-19 $X=8.675 $Y=2.4 $X2=0
+ $Y2=0
cc_463 N_A_M1023_g N_A_1191_368#_c_1048_n 8.84614e-19 $X=9.125 $Y=2.4 $X2=0
+ $Y2=0
cc_464 A N_A_1191_368#_c_1048_n 0.0235495f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_465 N_A_c_499_n N_A_1191_368#_c_1048_n 5.53009e-19 $X=9.515 $Y=1.515 $X2=0
+ $Y2=0
cc_466 N_A_M1005_g N_VGND_c_1082_n 0.00472678f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_467 N_A_M1005_g N_VGND_c_1083_n 5.07377e-19 $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_468 N_A_M1007_g N_VGND_c_1083_n 0.0100479f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_469 N_A_M1015_g N_VGND_c_1083_n 0.0100479f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_470 N_A_M1029_g N_VGND_c_1083_n 5.07377e-19 $X=9.515 $Y=0.74 $X2=0 $Y2=0
cc_471 N_A_M1029_g N_VGND_c_1085_n 0.018401f $X=9.515 $Y=0.74 $X2=0 $Y2=0
cc_472 N_A_c_499_n N_VGND_c_1085_n 0.00132967f $X=9.515 $Y=1.515 $X2=0 $Y2=0
cc_473 N_A_M1005_g N_VGND_c_1093_n 0.00434272f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_474 N_A_M1007_g N_VGND_c_1093_n 0.00383152f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_475 N_A_M1015_g N_VGND_c_1094_n 0.00383152f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_476 N_A_M1029_g N_VGND_c_1094_n 0.00434272f $X=9.515 $Y=0.74 $X2=0 $Y2=0
cc_477 N_A_M1005_g N_VGND_c_1102_n 0.00821489f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_478 N_A_M1007_g N_VGND_c_1102_n 0.0075754f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_479 N_A_M1015_g N_VGND_c_1102_n 0.0075754f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_480 N_A_M1029_g N_VGND_c_1102_n 0.00823934f $X=9.515 $Y=0.74 $X2=0 $Y2=0
cc_481 N_VPWR_c_579_n N_A_319_368#_c_680_n 0.0523105f $X=1.18 $Y=2.265 $X2=0
+ $Y2=0
cc_482 N_VPWR_c_583_n N_A_319_368#_c_681_n 0.0439866f $X=8.285 $Y=3.33 $X2=0
+ $Y2=0
cc_483 N_VPWR_c_576_n N_A_319_368#_c_681_n 0.0246722f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_484 N_VPWR_c_579_n N_A_319_368#_c_682_n 0.0119897f $X=1.18 $Y=2.265 $X2=0
+ $Y2=0
cc_485 N_VPWR_c_583_n N_A_319_368#_c_682_n 0.0179217f $X=8.285 $Y=3.33 $X2=0
+ $Y2=0
cc_486 N_VPWR_c_576_n N_A_319_368#_c_682_n 0.00971942f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_487 N_VPWR_c_583_n N_A_319_368#_c_683_n 0.0620209f $X=8.285 $Y=3.33 $X2=0
+ $Y2=0
cc_488 N_VPWR_c_576_n N_A_319_368#_c_683_n 0.0342927f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_489 N_VPWR_c_583_n N_A_319_368#_c_684_n 0.0200723f $X=8.285 $Y=3.33 $X2=0
+ $Y2=0
cc_490 N_VPWR_c_576_n N_A_319_368#_c_684_n 0.0108858f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_491 N_VPWR_c_576_n N_A_319_368#_c_698_n 0.00573193f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_492 N_VPWR_c_583_n N_A_781_368#_c_946_n 0.0422142f $X=8.285 $Y=3.33 $X2=0
+ $Y2=0
cc_493 N_VPWR_c_576_n N_A_781_368#_c_946_n 0.0237116f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_494 N_VPWR_c_583_n N_A_781_368#_c_947_n 0.0749947f $X=8.285 $Y=3.33 $X2=0
+ $Y2=0
cc_495 N_VPWR_c_576_n N_A_781_368#_c_947_n 0.0428557f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_496 N_VPWR_c_580_n N_A_781_368#_c_948_n 0.00273527f $X=8.45 $Y=2.455 $X2=0
+ $Y2=0
cc_497 N_VPWR_c_583_n N_A_781_368#_c_948_n 0.0618931f $X=8.285 $Y=3.33 $X2=0
+ $Y2=0
cc_498 N_VPWR_c_576_n N_A_781_368#_c_948_n 0.0343914f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_499 N_VPWR_c_583_n N_A_781_368#_c_949_n 0.0225681f $X=8.285 $Y=3.33 $X2=0
+ $Y2=0
cc_500 N_VPWR_c_576_n N_A_781_368#_c_949_n 0.0124607f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_501 N_VPWR_c_583_n N_A_781_368#_c_950_n 0.0226702f $X=8.285 $Y=3.33 $X2=0
+ $Y2=0
cc_502 N_VPWR_c_576_n N_A_781_368#_c_950_n 0.0124639f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_503 N_VPWR_c_583_n N_A_781_368#_c_951_n 0.0235512f $X=8.285 $Y=3.33 $X2=0
+ $Y2=0
cc_504 N_VPWR_c_576_n N_A_781_368#_c_951_n 0.0126924f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_505 N_VPWR_c_580_n N_A_1191_368#_c_1007_n 0.0255604f $X=8.45 $Y=2.455 $X2=0
+ $Y2=0
cc_506 N_VPWR_c_583_n N_A_1191_368#_c_1007_n 0.0101736f $X=8.285 $Y=3.33 $X2=0
+ $Y2=0
cc_507 N_VPWR_c_576_n N_A_1191_368#_c_1007_n 0.0084208f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_508 N_VPWR_M1020_d N_A_1191_368#_c_1033_n 0.00314376f $X=8.315 $Y=1.84 $X2=0
+ $Y2=0
cc_509 N_VPWR_c_580_n N_A_1191_368#_c_1033_n 0.0148589f $X=8.45 $Y=2.455 $X2=0
+ $Y2=0
cc_510 N_VPWR_c_580_n N_A_1191_368#_c_1008_n 0.0234083f $X=8.45 $Y=2.455 $X2=0
+ $Y2=0
cc_511 N_VPWR_c_581_n N_A_1191_368#_c_1008_n 0.0234083f $X=9.35 $Y=2.455 $X2=0
+ $Y2=0
cc_512 N_VPWR_c_584_n N_A_1191_368#_c_1008_n 0.0144623f $X=9.265 $Y=3.33 $X2=0
+ $Y2=0
cc_513 N_VPWR_c_576_n N_A_1191_368#_c_1008_n 0.0118344f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_514 N_VPWR_M1023_d N_A_1191_368#_c_1041_n 0.00314376f $X=9.215 $Y=1.84 $X2=0
+ $Y2=0
cc_515 N_VPWR_c_581_n N_A_1191_368#_c_1041_n 0.0148589f $X=9.35 $Y=2.455 $X2=0
+ $Y2=0
cc_516 N_VPWR_c_581_n N_A_1191_368#_c_1010_n 0.0224614f $X=9.35 $Y=2.455 $X2=0
+ $Y2=0
cc_517 N_VPWR_c_585_n N_A_1191_368#_c_1010_n 0.011066f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_518 N_VPWR_c_576_n N_A_1191_368#_c_1010_n 0.00915947f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_519 N_A_319_368#_c_681_n N_Y_M1022_d 0.00165831f $X=2.525 $Y=2.99 $X2=0 $Y2=0
cc_520 N_A_319_368#_c_683_n N_Y_M1026_d 0.00165831f $X=3.475 $Y=2.99 $X2=0 $Y2=0
cc_521 N_A_319_368#_c_680_n N_Y_c_767_n 0.00696138f $X=1.74 $Y=1.985 $X2=0 $Y2=0
cc_522 N_A_319_368#_c_681_n N_Y_c_784_n 0.0159318f $X=2.525 $Y=2.99 $X2=0 $Y2=0
cc_523 N_A_319_368#_M1024_s N_Y_c_768_n 0.00218982f $X=2.505 $Y=1.84 $X2=0 $Y2=0
cc_524 N_A_319_368#_c_721_p N_Y_c_768_n 0.0167599f $X=2.66 $Y=2.325 $X2=0 $Y2=0
cc_525 N_A_319_368#_c_683_n N_Y_c_795_n 0.0159318f $X=3.475 $Y=2.99 $X2=0 $Y2=0
cc_526 N_A_319_368#_M1027_s N_Y_c_797_n 0.00400506f $X=3.455 $Y=1.84 $X2=0 $Y2=0
cc_527 N_A_319_368#_M1001_s N_Y_c_797_n 0.0045988f $X=4.405 $Y=1.84 $X2=0 $Y2=0
cc_528 N_A_319_368#_M1032_s N_Y_c_797_n 0.00459125f $X=5.405 $Y=1.84 $X2=0 $Y2=0
cc_529 N_A_319_368#_c_695_n N_Y_c_797_n 0.0132121f $X=3.615 $Y=2.49 $X2=0 $Y2=0
cc_530 N_A_319_368#_c_698_n N_Y_c_797_n 0.0328444f $X=4.425 $Y=2.505 $X2=0 $Y2=0
cc_531 N_A_319_368#_c_700_n N_Y_c_797_n 0.0554982f $X=4.755 $Y=2.505 $X2=0 $Y2=0
cc_532 N_A_319_368#_c_685_n N_Y_c_797_n 0.0144054f $X=5.54 $Y=2.375 $X2=0 $Y2=0
cc_533 N_A_319_368#_M1032_s Y 0.00219719f $X=5.405 $Y=1.84 $X2=0 $Y2=0
cc_534 N_A_319_368#_c_698_n N_A_781_368#_M1000_d 0.00438523f $X=4.425 $Y=2.505
+ $X2=-0.19 $Y2=1.66
cc_535 N_A_319_368#_c_702_n N_A_781_368#_M1031_d 0.00385282f $X=5.44 $Y=2.415
+ $X2=0 $Y2=0
cc_536 N_A_319_368#_M1001_s N_A_781_368#_c_946_n 0.00255072f $X=4.405 $Y=1.84
+ $X2=0 $Y2=0
cc_537 N_A_319_368#_c_698_n N_A_781_368#_c_946_n 0.00421866f $X=4.425 $Y=2.505
+ $X2=0 $Y2=0
cc_538 N_A_319_368#_c_700_n N_A_781_368#_c_946_n 0.0160324f $X=4.755 $Y=2.505
+ $X2=0 $Y2=0
cc_539 N_A_319_368#_c_702_n N_A_781_368#_c_946_n 0.00527089f $X=5.44 $Y=2.415
+ $X2=0 $Y2=0
cc_540 N_A_319_368#_M1032_s N_A_781_368#_c_947_n 0.0037093f $X=5.405 $Y=1.84
+ $X2=0 $Y2=0
cc_541 N_A_319_368#_c_685_n N_A_781_368#_c_947_n 0.00899023f $X=5.54 $Y=2.375
+ $X2=0 $Y2=0
cc_542 N_A_319_368#_c_702_n N_A_781_368#_c_947_n 0.00464895f $X=5.44 $Y=2.415
+ $X2=0 $Y2=0
cc_543 N_A_319_368#_c_683_n N_A_781_368#_c_949_n 0.0119238f $X=3.475 $Y=2.99
+ $X2=0 $Y2=0
cc_544 N_A_319_368#_c_698_n N_A_781_368#_c_949_n 0.017773f $X=4.425 $Y=2.505
+ $X2=0 $Y2=0
cc_545 N_A_319_368#_c_700_n N_A_781_368#_c_950_n 0.0067138f $X=4.755 $Y=2.505
+ $X2=0 $Y2=0
cc_546 N_A_319_368#_c_702_n N_A_781_368#_c_950_n 0.0165787f $X=5.44 $Y=2.415
+ $X2=0 $Y2=0
cc_547 N_A_319_368#_c_685_n N_A_1191_368#_c_1011_n 0.0173479f $X=5.54 $Y=2.375
+ $X2=0 $Y2=0
cc_548 N_Y_c_797_n N_A_781_368#_M1000_d 0.0042731f $X=5.405 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_549 N_Y_c_797_n N_A_781_368#_M1031_d 0.00411427f $X=5.405 $Y=2.035 $X2=0
+ $Y2=0
cc_550 N_Y_c_797_n N_A_1191_368#_c_1011_n 0.0103789f $X=5.405 $Y=2.035 $X2=0
+ $Y2=0
cc_551 N_Y_c_746_n N_VGND_M1003_s 0.00263002f $X=2.5 $Y=1.065 $X2=0 $Y2=0
cc_552 N_Y_c_751_n N_VGND_M1025_d 0.0101061f $X=4.905 $Y=1.095 $X2=0 $Y2=0
cc_553 N_Y_c_753_n N_VGND_M1034_d 0.00628546f $X=6.25 $Y=1.095 $X2=0 $Y2=0
cc_554 N_Y_c_754_n N_VGND_M1034_d 0.00283795f $X=5.635 $Y=1.095 $X2=0 $Y2=0
cc_555 N_Y_c_756_n N_VGND_M1008_s 0.00271958f $X=7.25 $Y=1.095 $X2=0 $Y2=0
cc_556 N_Y_c_758_n N_VGND_M1019_s 0.0042801f $X=8.275 $Y=1.095 $X2=0 $Y2=0
cc_557 N_Y_c_760_n N_VGND_M1007_s 0.00191292f $X=9.215 $Y=1.095 $X2=0 $Y2=0
cc_558 N_Y_c_745_n N_VGND_c_1077_n 0.023308f $X=1.735 $Y=0.515 $X2=0 $Y2=0
cc_559 N_Y_c_747_n N_VGND_c_1077_n 0.00625076f $X=1.82 $Y=1.065 $X2=0 $Y2=0
cc_560 N_Y_c_745_n N_VGND_c_1078_n 0.0164981f $X=1.735 $Y=0.515 $X2=0 $Y2=0
cc_561 N_Y_c_746_n N_VGND_c_1078_n 0.0193036f $X=2.5 $Y=1.065 $X2=0 $Y2=0
cc_562 N_Y_c_748_n N_VGND_c_1078_n 0.0173003f $X=2.665 $Y=0.515 $X2=0 $Y2=0
cc_563 N_Y_c_748_n N_VGND_c_1079_n 0.0308109f $X=2.665 $Y=0.515 $X2=0 $Y2=0
cc_564 N_Y_c_749_n N_VGND_c_1079_n 0.0277025f $X=3.5 $Y=1.385 $X2=0 $Y2=0
cc_565 N_Y_c_750_n N_VGND_c_1079_n 0.0295934f $X=3.665 $Y=0.515 $X2=0 $Y2=0
cc_566 N_Y_c_752_n N_VGND_c_1080_n 0.0192667f $X=5.07 $Y=0.515 $X2=0 $Y2=0
cc_567 N_Y_c_754_n N_VGND_c_1080_n 0.0529279f $X=5.635 $Y=1.095 $X2=0 $Y2=0
cc_568 N_Y_c_755_n N_VGND_c_1080_n 0.0192667f $X=6.415 $Y=0.515 $X2=0 $Y2=0
cc_569 N_Y_c_755_n N_VGND_c_1081_n 0.0178632f $X=6.415 $Y=0.515 $X2=0 $Y2=0
cc_570 N_Y_c_756_n N_VGND_c_1081_n 0.0182382f $X=7.25 $Y=1.095 $X2=0 $Y2=0
cc_571 N_Y_c_757_n N_VGND_c_1081_n 0.0178632f $X=7.415 $Y=0.515 $X2=0 $Y2=0
cc_572 N_Y_c_757_n N_VGND_c_1082_n 0.017872f $X=7.415 $Y=0.515 $X2=0 $Y2=0
cc_573 N_Y_c_758_n N_VGND_c_1082_n 0.0234251f $X=8.275 $Y=1.095 $X2=0 $Y2=0
cc_574 N_Y_c_759_n N_VGND_c_1082_n 0.0171608f $X=8.44 $Y=0.515 $X2=0 $Y2=0
cc_575 N_Y_c_759_n N_VGND_c_1083_n 0.0170358f $X=8.44 $Y=0.515 $X2=0 $Y2=0
cc_576 N_Y_c_760_n N_VGND_c_1083_n 0.0148206f $X=9.215 $Y=1.095 $X2=0 $Y2=0
cc_577 N_Y_c_761_n N_VGND_c_1083_n 0.0170358f $X=9.3 $Y=0.515 $X2=0 $Y2=0
cc_578 N_Y_c_760_n N_VGND_c_1085_n 0.00584871f $X=9.215 $Y=1.095 $X2=0 $Y2=0
cc_579 N_Y_c_761_n N_VGND_c_1085_n 0.0244878f $X=9.3 $Y=0.515 $X2=0 $Y2=0
cc_580 N_Y_c_745_n N_VGND_c_1087_n 0.011066f $X=1.735 $Y=0.515 $X2=0 $Y2=0
cc_581 N_Y_c_748_n N_VGND_c_1088_n 0.0144922f $X=2.665 $Y=0.515 $X2=0 $Y2=0
cc_582 N_Y_c_750_n N_VGND_c_1089_n 0.0313451f $X=3.665 $Y=0.515 $X2=0 $Y2=0
cc_583 N_Y_c_751_n N_VGND_c_1089_n 0.0596318f $X=4.905 $Y=1.095 $X2=0 $Y2=0
cc_584 N_Y_c_752_n N_VGND_c_1089_n 0.019268f $X=5.07 $Y=0.515 $X2=0 $Y2=0
cc_585 N_Y_c_752_n N_VGND_c_1090_n 0.0144609f $X=5.07 $Y=0.515 $X2=0 $Y2=0
cc_586 N_Y_c_755_n N_VGND_c_1091_n 0.0145639f $X=6.415 $Y=0.515 $X2=0 $Y2=0
cc_587 N_Y_c_757_n N_VGND_c_1092_n 0.0144922f $X=7.415 $Y=0.515 $X2=0 $Y2=0
cc_588 N_Y_c_759_n N_VGND_c_1093_n 0.0109942f $X=8.44 $Y=0.515 $X2=0 $Y2=0
cc_589 N_Y_c_761_n N_VGND_c_1094_n 0.0109942f $X=9.3 $Y=0.515 $X2=0 $Y2=0
cc_590 N_Y_c_745_n N_VGND_c_1102_n 0.00915947f $X=1.735 $Y=0.515 $X2=0 $Y2=0
cc_591 N_Y_c_748_n N_VGND_c_1102_n 0.0118826f $X=2.665 $Y=0.515 $X2=0 $Y2=0
cc_592 N_Y_c_750_n N_VGND_c_1102_n 0.00904371f $X=3.665 $Y=0.515 $X2=0 $Y2=0
cc_593 N_Y_c_752_n N_VGND_c_1102_n 0.0118703f $X=5.07 $Y=0.515 $X2=0 $Y2=0
cc_594 N_Y_c_755_n N_VGND_c_1102_n 0.0119984f $X=6.415 $Y=0.515 $X2=0 $Y2=0
cc_595 N_Y_c_757_n N_VGND_c_1102_n 0.0118826f $X=7.415 $Y=0.515 $X2=0 $Y2=0
cc_596 N_Y_c_759_n N_VGND_c_1102_n 0.00904371f $X=8.44 $Y=0.515 $X2=0 $Y2=0
cc_597 N_Y_c_761_n N_VGND_c_1102_n 0.00904371f $X=9.3 $Y=0.515 $X2=0 $Y2=0
cc_598 N_A_781_368#_c_947_n N_A_1191_368#_M1014_s 0.00266942f $X=6.435 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_599 N_A_781_368#_c_948_n N_A_1191_368#_M1016_s 0.00218982f $X=7.465 $Y=2.99
+ $X2=0 $Y2=0
cc_600 N_A_781_368#_M1014_d N_A_1191_368#_c_1013_n 0.00410979f $X=6.415 $Y=1.84
+ $X2=0 $Y2=0
cc_601 N_A_781_368#_c_962_n N_A_1191_368#_c_1013_n 0.0189268f $X=6.6 $Y=2.455
+ $X2=0 $Y2=0
cc_602 N_A_781_368#_c_948_n N_A_1191_368#_c_1017_n 0.0177084f $X=7.465 $Y=2.99
+ $X2=0 $Y2=0
cc_603 N_A_781_368#_M1017_d N_A_1191_368#_c_1019_n 0.00420477f $X=7.415 $Y=1.84
+ $X2=0 $Y2=0
cc_604 N_A_781_368#_c_967_n N_A_1191_368#_c_1019_n 0.0148589f $X=7.55 $Y=2.455
+ $X2=0 $Y2=0
cc_605 N_A_781_368#_c_948_n N_A_1191_368#_c_1007_n 0.00391086f $X=7.465 $Y=2.99
+ $X2=0 $Y2=0
cc_606 N_A_781_368#_c_947_n N_A_1191_368#_c_1011_n 0.0205035f $X=6.435 $Y=2.99
+ $X2=0 $Y2=0

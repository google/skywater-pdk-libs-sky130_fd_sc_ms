* NGSPICE file created from sky130_fd_sc_ms__a31oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 a_200_74# A1 Y VNB nlowvt w=740000u l=150000u
+  ad=4.773e+11p pd=4.25e+06u as=7.548e+11p ps=5e+06u
M1001 Y B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=5.217e+11p ps=4.37e+06u
M1002 a_27_368# A3 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=1.6464e+12p pd=1.414e+07u as=9.744e+11p ps=8.46e+06u
M1003 VPWR A2 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A3 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y A1 a_200_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A3 a_114_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.662e+11p ps=4.22e+06u
M1007 a_114_74# A2 a_200_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_368# A2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1010 VPWR A1 a_27_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_114_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_200_74# A2 a_114_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_368# B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__nand4b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.985000 1.510000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.350000 2.590000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.350000 4.195000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.558000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.445000 1.350000 5.635000 1.780000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.573400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 0.800000 1.895000 1.010000 ;
        RECT 1.535000 1.010000 3.235000 1.180000 ;
        RECT 1.550000 1.850000 1.825000 1.950000 ;
        RECT 1.550000 1.950000 5.190000 2.120000 ;
        RECT 1.550000 2.120000 1.825000 2.980000 ;
        RECT 2.760000 1.820000 3.235000 1.950000 ;
        RECT 2.760000 2.120000 3.090000 2.980000 ;
        RECT 3.005000 1.180000 3.235000 1.820000 ;
        RECT 3.760000 2.120000 4.090000 2.980000 ;
        RECT 4.860000 2.120000 5.190000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  0.350000 0.365000 0.840000 ;
      RECT 0.115000  0.840000 1.325000 1.010000 ;
      RECT 0.505000  1.680000 1.325000 1.850000 ;
      RECT 0.505000  1.850000 0.835000 2.860000 ;
      RECT 0.545000  0.085000 0.875000 0.670000 ;
      RECT 1.040000  2.020000 1.370000 3.245000 ;
      RECT 1.105000  0.350000 2.325000 0.630000 ;
      RECT 1.155000  1.010000 1.325000 1.350000 ;
      RECT 1.155000  1.350000 1.720000 1.680000 ;
      RECT 1.995000  2.290000 2.590000 3.245000 ;
      RECT 2.075000  0.630000 2.325000 0.670000 ;
      RECT 2.075000  0.670000 3.345000 0.840000 ;
      RECT 2.505000  0.255000 4.335000 0.425000 ;
      RECT 2.505000  0.425000 2.835000 0.500000 ;
      RECT 3.015000  0.595000 3.345000 0.670000 ;
      RECT 3.260000  2.290000 3.590000 3.245000 ;
      RECT 3.575000  0.595000 3.825000 0.930000 ;
      RECT 3.575000  0.930000 5.645000 1.180000 ;
      RECT 4.005000  0.425000 4.335000 0.760000 ;
      RECT 4.320000  2.290000 4.650000 3.245000 ;
      RECT 4.505000  0.400000 4.695000 0.930000 ;
      RECT 4.865000  0.085000 5.195000 0.760000 ;
      RECT 5.360000  1.950000 5.645000 3.245000 ;
      RECT 5.395000  0.400000 5.645000 0.930000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_ms__nand4b_2
END LIBRARY

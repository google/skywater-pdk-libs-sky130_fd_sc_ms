* File: sky130_fd_sc_ms__or4_4.pex.spice
* Created: Fri Aug 28 18:09:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__OR4_4%A_83_264# 1 2 3 12 16 20 24 28 32 36 40 42 48
+ 49 50 53 55 59 61 63 66 69 70 71 77
c164 61 0 6.34286e-20 $X=6.465 $Y=1.11
r165 84 85 59.4247 $w=2.92e-07 $l=3.6e-07 $layer=POLY_cond $X=1.495 $Y=1.485
+ $X2=1.855 $Y2=1.485
r166 81 82 67.6781 $w=2.92e-07 $l=4.1e-07 $layer=POLY_cond $X=0.995 $Y=1.485
+ $X2=1.405 $Y2=1.485
r167 75 77 8.91885 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=5.46 $Y=2.07
+ $X2=5.625 $Y2=2.07
r168 71 72 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=4.935 $Y=0.875
+ $X2=4.935 $Y2=1.11
r169 69 87 14.8562 $w=2.92e-07 $l=9e-08 $layer=POLY_cond $X=2.16 $Y=1.485
+ $X2=2.25 $Y2=1.485
r170 69 85 50.3459 $w=2.92e-07 $l=3.05e-07 $layer=POLY_cond $X=2.16 $Y=1.485
+ $X2=1.855 $Y2=1.485
r171 68 69 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.16
+ $Y=1.485 $X2=2.16 $Y2=1.485
r172 65 66 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=6.55 $Y=1.195
+ $X2=6.55 $Y2=1.95
r173 63 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.465 $Y=2.035
+ $X2=6.55 $Y2=1.95
r174 63 77 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=6.465 $Y=2.035
+ $X2=5.625 $Y2=2.035
r175 62 72 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.1 $Y=1.11
+ $X2=4.935 $Y2=1.11
r176 61 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.465 $Y=1.11
+ $X2=6.55 $Y2=1.195
r177 61 62 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=6.465 $Y=1.11
+ $X2=5.1 $Y2=1.11
r178 57 71 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.935 $Y=0.79
+ $X2=4.935 $Y2=0.875
r179 57 59 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.935 $Y=0.79
+ $X2=4.935 $Y2=0.515
r180 56 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.25 $Y=0.875
+ $X2=3.085 $Y2=0.875
r181 55 71 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.77 $Y=0.875
+ $X2=4.935 $Y2=0.875
r182 55 56 99.1658 $w=1.68e-07 $l=1.52e-06 $layer=LI1_cond $X=4.77 $Y=0.875
+ $X2=3.25 $Y2=0.875
r183 51 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=0.79
+ $X2=3.085 $Y2=0.875
r184 51 53 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.085 $Y=0.79
+ $X2=3.085 $Y2=0.515
r185 49 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.92 $Y=0.875
+ $X2=3.085 $Y2=0.875
r186 49 50 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.92 $Y=0.875
+ $X2=2.325 $Y2=0.875
r187 48 68 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=1.32
+ $X2=2.24 $Y2=1.485
r188 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.24 $Y=0.96
+ $X2=2.325 $Y2=0.875
r189 47 48 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.24 $Y=0.96
+ $X2=2.24 $Y2=1.32
r190 45 84 2.47603 $w=2.92e-07 $l=1.5e-08 $layer=POLY_cond $X=1.48 $Y=1.485
+ $X2=1.495 $Y2=1.485
r191 45 82 12.3801 $w=2.92e-07 $l=7.5e-08 $layer=POLY_cond $X=1.48 $Y=1.485
+ $X2=1.405 $Y2=1.485
r192 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.48
+ $Y=1.485 $X2=1.48 $Y2=1.485
r193 42 68 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=1.485
+ $X2=2.24 $Y2=1.485
r194 42 44 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.155 $Y=1.485
+ $X2=1.48 $Y2=1.485
r195 38 87 18.3338 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.32
+ $X2=2.25 $Y2=1.485
r196 38 40 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.25 $Y=1.32
+ $X2=2.25 $Y2=0.74
r197 34 85 14.0951 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.65
+ $X2=1.855 $Y2=1.485
r198 34 36 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=1.855 $Y=1.65
+ $X2=1.855 $Y2=2.4
r199 30 84 18.3338 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.495 $Y=1.32
+ $X2=1.495 $Y2=1.485
r200 30 32 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.495 $Y=1.32
+ $X2=1.495 $Y2=0.74
r201 26 82 14.0951 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.65
+ $X2=1.405 $Y2=1.485
r202 26 28 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=1.405 $Y=1.65
+ $X2=1.405 $Y2=2.4
r203 22 81 18.3338 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.32
+ $X2=0.995 $Y2=1.485
r204 22 24 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.995 $Y=1.32
+ $X2=0.995 $Y2=0.74
r205 18 81 6.60274 $w=2.92e-07 $l=4e-08 $layer=POLY_cond $X=0.955 $Y=1.485
+ $X2=0.995 $Y2=1.485
r206 18 79 64.3767 $w=2.92e-07 $l=3.9e-07 $layer=POLY_cond $X=0.955 $Y=1.485
+ $X2=0.565 $Y2=1.485
r207 18 20 322.629 $w=1.8e-07 $l=8.3e-07 $layer=POLY_cond $X=0.955 $Y=1.57
+ $X2=0.955 $Y2=2.4
r208 14 79 18.3338 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=1.32
+ $X2=0.565 $Y2=1.485
r209 14 16 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.565 $Y=1.32
+ $X2=0.565 $Y2=0.74
r210 10 79 9.90411 $w=2.92e-07 $l=6e-08 $layer=POLY_cond $X=0.505 $Y=1.485
+ $X2=0.565 $Y2=1.485
r211 10 12 322.629 $w=1.8e-07 $l=8.3e-07 $layer=POLY_cond $X=0.505 $Y=1.57
+ $X2=0.505 $Y2=2.4
r212 3 75 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.325
+ $Y=1.96 $X2=5.46 $Y2=2.105
r213 2 59 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.795
+ $Y=0.37 $X2=4.935 $Y2=0.515
r214 1 53 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.945
+ $Y=0.37 $X2=3.085 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR4_4%B 1 3 5 7 10 12 13 14 18 20 21
c83 14 0 1.3894e-19 $X=4.23 $Y=1.215
c84 10 0 1.72297e-19 $X=4.235 $Y=2.46
r85 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.78
+ $Y=1.385 $X2=2.78 $Y2=1.385
r86 21 26 10.3184 $w=4.02e-07 $l=3.4e-07 $layer=LI1_cond $X=3.12 $Y=1.34
+ $X2=2.78 $Y2=1.34
r87 20 26 4.24876 $w=4.02e-07 $l=1.4e-07 $layer=LI1_cond $X=2.64 $Y=1.34
+ $X2=2.78 $Y2=1.34
r88 18 29 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.23 $Y=1.385
+ $X2=4.23 $Y2=1.55
r89 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.23
+ $Y=1.385 $X2=4.23 $Y2=1.385
r90 14 17 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.23 $Y=1.215
+ $X2=4.23 $Y2=1.385
r91 13 21 7.646 $w=4.02e-07 $l=1.73205e-07 $layer=LI1_cond $X=3.235 $Y=1.215
+ $X2=3.12 $Y2=1.34
r92 12 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.065 $Y=1.215
+ $X2=4.23 $Y2=1.215
r93 12 13 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.065 $Y=1.215
+ $X2=3.235 $Y2=1.215
r94 10 29 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=4.235 $Y=2.46
+ $X2=4.235 $Y2=1.55
r95 5 25 38.5662 $w=2.97e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.87 $Y=1.22
+ $X2=2.785 $Y2=1.385
r96 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.87 $Y=1.22 $X2=2.87
+ $Y2=0.74
r97 1 25 48.8089 $w=2.97e-07 $l=2.92276e-07 $layer=POLY_cond $X=2.865 $Y=1.64
+ $X2=2.785 $Y2=1.385
r98 1 3 318.742 $w=1.8e-07 $l=8.2e-07 $layer=POLY_cond $X=2.865 $Y=1.64
+ $X2=2.865 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__OR4_4%A 3 7 11 13 21
c47 7 0 1.55268e-19 $X=3.315 $Y=2.46
r48 19 21 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=3.57 $Y=1.635
+ $X2=3.765 $Y2=1.635
r49 17 19 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=3.315 $Y=1.635
+ $X2=3.57 $Y2=1.635
r50 15 17 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.3 $Y=1.635
+ $X2=3.315 $Y2=1.635
r51 13 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.635 $X2=3.57 $Y2=1.635
r52 9 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.765 $Y=1.8
+ $X2=3.765 $Y2=1.635
r53 9 11 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.765 $Y=1.8
+ $X2=3.765 $Y2=2.46
r54 5 17 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.315 $Y=1.8
+ $X2=3.315 $Y2=1.635
r55 5 7 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.315 $Y=1.8 $X2=3.315
+ $Y2=2.46
r56 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.3 $Y=1.47 $X2=3.3
+ $Y2=1.635
r57 1 3 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=3.3 $Y=1.47 $X2=3.3
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__OR4_4%C 3 7 11 13 14 15 20 25 26 29
c67 20 0 1.3894e-19 $X=4.77 $Y=1.605
c68 7 0 2.84905e-19 $X=4.735 $Y=2.46
c69 3 0 6.34286e-20 $X=4.72 $Y=0.74
r70 25 28 55.5535 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=6.15 $Y=1.53
+ $X2=6.15 $Y2=1.78
r71 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.15
+ $Y=1.53 $X2=6.15 $Y2=1.53
r72 20 23 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=1.605
+ $X2=4.77 $Y2=1.77
r73 20 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=1.605
+ $X2=4.77 $Y2=1.44
r74 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.77
+ $Y=1.605 $X2=4.77 $Y2=1.605
r75 15 26 4.16546 $w=4.13e-07 $l=1.5e-07 $layer=LI1_cond $X=6 $Y=1.572 $X2=6.15
+ $Y2=1.572
r76 14 15 13.3295 $w=4.13e-07 $l=4.8e-07 $layer=LI1_cond $X=5.52 $Y=1.572 $X2=6
+ $Y2=1.572
r77 14 29 4.99855 $w=4.13e-07 $l=1.8e-07 $layer=LI1_cond $X=5.52 $Y=1.572
+ $X2=5.34 $Y2=1.572
r78 13 29 8.81928 $w=4.15e-07 $l=3e-07 $layer=LI1_cond $X=5.04 $Y=1.572 $X2=5.34
+ $Y2=1.572
r79 13 21 8.03415 $w=4.1e-07 $l=2.7e-07 $layer=LI1_cond $X=5.04 $Y=1.572
+ $X2=4.77 $Y2=1.572
r80 11 28 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=6.135 $Y=2.46
+ $X2=6.135 $Y2=1.78
r81 7 23 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=4.735 $Y=2.46
+ $X2=4.735 $Y2=1.77
r82 3 22 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=4.72 $Y=0.74 $X2=4.72
+ $Y2=1.44
.ends

.subckt PM_SKY130_FD_SC_MS__OR4_4%D 1 3 6 10 13 14 15 20 23 26 27
c56 26 0 7.13014e-20 $X=6.45 $Y=0.42
r57 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.45
+ $Y=0.42 $X2=6.45 $Y2=0.42
r58 23 27 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=6.45 $Y=0.555
+ $X2=6.45 $Y2=0.42
r59 22 26 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=6.45 $Y=0.775
+ $X2=6.45 $Y2=0.42
r60 19 20 2.99935 $w=3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.685 $Y=1.335 $X2=5.7
+ $Y2=1.335
r61 18 19 89.9803 $w=3e-07 $l=4.5e-07 $layer=POLY_cond $X=5.235 $Y=1.335
+ $X2=5.685 $Y2=1.335
r62 16 18 2.99935 $w=3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.22 $Y=1.335
+ $X2=5.235 $Y2=1.335
r63 14 22 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=6.285 $Y=0.85
+ $X2=6.45 $Y2=0.775
r64 14 15 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=6.285 $Y=0.85
+ $X2=5.775 $Y2=0.85
r65 13 20 18.9685 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=5.7 $Y=1.185 $X2=5.7
+ $Y2=1.335
r66 12 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.7 $Y=0.925
+ $X2=5.775 $Y2=0.85
r67 12 13 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=5.7 $Y=0.925 $X2=5.7
+ $Y2=1.185
r68 8 19 14.7197 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.685 $Y=1.485
+ $X2=5.685 $Y2=1.335
r69 8 10 378.992 $w=1.8e-07 $l=9.75e-07 $layer=POLY_cond $X=5.685 $Y=1.485
+ $X2=5.685 $Y2=2.46
r70 4 18 14.7197 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.235 $Y=1.485
+ $X2=5.235 $Y2=1.335
r71 4 6 378.992 $w=1.8e-07 $l=9.75e-07 $layer=POLY_cond $X=5.235 $Y=1.485
+ $X2=5.235 $Y2=2.46
r72 1 16 18.9685 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=5.22 $Y=1.185
+ $X2=5.22 $Y2=1.335
r73 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.22 $Y=1.185
+ $X2=5.22 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__OR4_4%VPWR 1 2 3 4 13 15 19 23 27 29 31 36 41 51 52
+ 58 61 64
r86 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r87 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r88 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r89 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r90 51 52 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r91 49 52 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=6.48 $Y2=3.33
r92 49 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r93 48 51 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=6.48 $Y2=3.33
r94 48 49 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r95 46 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=3.54 $Y2=3.33
r96 46 48 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=4.08 $Y2=3.33
r97 45 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r98 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r99 42 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.08 $Y2=3.33
r100 42 44 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=3.12 $Y2=3.33
r101 41 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=3.33
+ $X2=3.54 $Y2=3.33
r102 41 44 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.375 $Y=3.33
+ $X2=3.12 $Y2=3.33
r103 40 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r104 40 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r105 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r106 37 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.18 $Y2=3.33
r107 37 39 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r108 36 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.915 $Y=3.33
+ $X2=2.08 $Y2=3.33
r109 36 39 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.915 $Y=3.33
+ $X2=1.68 $Y2=3.33
r110 35 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r111 35 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r112 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r113 32 55 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r114 32 34 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r115 31 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.18 $Y2=3.33
r116 31 34 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.72 $Y2=3.33
r117 29 65 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.6 $Y2=3.33
r118 29 45 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r119 25 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=3.245
+ $X2=3.54 $Y2=3.33
r120 25 27 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.54 $Y=3.245
+ $X2=3.54 $Y2=2.815
r121 21 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=3.245
+ $X2=2.08 $Y2=3.33
r122 21 23 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=2.08 $Y=3.245
+ $X2=2.08 $Y2=2.405
r123 17 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r124 17 19 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.405
r125 13 55 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r126 13 15 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.405
r127 4 27 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.96 $X2=3.54 $Y2=2.815
r128 3 23 300 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=2 $X=1.945
+ $Y=1.84 $X2=2.08 $Y2=2.405
r129 2 19 300 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=2 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.405
r130 1 15 300 $w=1.7e-07 $l=6.33364e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.405
.ends

.subckt PM_SKY130_FD_SC_MS__OR4_4%X 1 2 3 4 15 17 19 21 25 29 31 33 34 35 42
r69 43 53 5.02295 $w=3.3e-07 $l=4.1e-07 $layer=LI1_cond $X=0.945 $Y=1.985
+ $X2=0.535 $Y2=1.985
r70 34 42 3.78902 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=1.63 $Y=1.985
+ $X2=1.515 $Y2=1.985
r71 34 46 3.78902 $w=3.3e-07 $l=1.15e-07 $layer=LI1_cond $X=1.63 $Y=1.985
+ $X2=1.745 $Y2=1.985
r72 34 35 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=1.755 $Y=1.985
+ $X2=2.16 $Y2=1.985
r73 34 46 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=1.755 $Y=1.985
+ $X2=1.745 $Y2=1.985
r74 33 42 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.2 $Y=1.985
+ $X2=1.515 $Y2=1.985
r75 33 43 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.2 $Y=1.985
+ $X2=0.945 $Y2=1.985
r76 31 53 0.890511 $w=6.85e-07 $l=5e-08 $layer=LI1_cond $X=0.535 $Y=2.035
+ $X2=0.535 $Y2=1.985
r77 27 29 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.78 $Y=0.98
+ $X2=1.78 $Y2=0.515
r78 23 34 2.66947 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.63 $Y=2.15
+ $X2=1.63 $Y2=1.985
r79 23 25 11.775 $w=2.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.63 $Y=2.15
+ $X2=1.63 $Y2=2.385
r80 22 53 16.3854 $w=6.85e-07 $l=1.10616e-06 $layer=LI1_cond $X=0.945 $Y=1.065
+ $X2=0.535 $Y2=1.985
r81 21 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.615 $Y=1.065
+ $X2=1.78 $Y2=0.98
r82 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=1.065
+ $X2=0.945 $Y2=1.065
r83 17 31 7.81937 $w=6.85e-07 $l=2.45866e-07 $layer=LI1_cond $X=0.73 $Y=2.15
+ $X2=0.535 $Y2=2.035
r84 17 19 11.775 $w=2.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.73 $Y=2.15
+ $X2=0.73 $Y2=2.385
r85 13 22 4.8017 $w=6.85e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.78 $Y=0.98
+ $X2=0.945 $Y2=1.065
r86 13 15 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.78 $Y=0.98
+ $X2=0.78 $Y2=0.515
r87 4 34 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.84 $X2=1.63 $Y2=1.985
r88 4 25 300 $w=1.7e-07 $l=6.08769e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.84 $X2=1.63 $Y2=2.385
r89 3 53 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=1.985
r90 3 19 300 $w=1.7e-07 $l=6.08769e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.385
r91 2 29 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.57
+ $Y=0.37 $X2=1.78 $Y2=0.515
r92 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.64
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR4_4%A_499_392# 1 2 3 10 12 14 16 17 20 22 30 32
c70 20 0 1.72297e-19 $X=4.51 $Y=2.815
r71 23 30 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.675 $Y=2.445
+ $X2=4.51 $Y2=2.445
r72 22 32 4.85386 $w=1.7e-07 $l=1.81659e-07 $layer=LI1_cond $X=6.245 $Y=2.445
+ $X2=6.41 $Y2=2.41
r73 22 23 102.428 $w=1.68e-07 $l=1.57e-06 $layer=LI1_cond $X=6.245 $Y=2.445
+ $X2=4.675 $Y2=2.445
r74 18 30 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.51 $Y=2.53 $X2=4.51
+ $Y2=2.445
r75 18 20 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=4.51 $Y=2.53
+ $X2=4.51 $Y2=2.815
r76 17 30 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.51 $Y=2.36 $X2=4.51
+ $Y2=2.445
r77 16 29 2.77363 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=4.51 $Y=2.14 $X2=4.51
+ $Y2=2.04
r78 16 17 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=4.51 $Y=2.14
+ $X2=4.51 $Y2=2.36
r79 15 27 3.96311 $w=1.7e-07 $l=1.69926e-07 $layer=LI1_cond $X=2.805 $Y=2.055
+ $X2=2.64 $Y2=2.065
r80 14 29 4.99254 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=4.345 $Y=2.055
+ $X2=4.51 $Y2=2.04
r81 14 15 100.471 $w=1.68e-07 $l=1.54e-06 $layer=LI1_cond $X=4.345 $Y=2.055
+ $X2=2.805 $Y2=2.055
r82 10 27 3.39695 $w=2.8e-07 $l=1.36931e-07 $layer=LI1_cond $X=2.615 $Y=2.19
+ $X2=2.64 $Y2=2.065
r83 10 12 10.4955 $w=2.78e-07 $l=2.55e-07 $layer=LI1_cond $X=2.615 $Y=2.19
+ $X2=2.615 $Y2=2.445
r84 3 32 300 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_PDIFF $count=2 $X=6.225
+ $Y=1.96 $X2=6.41 $Y2=2.455
r85 2 29 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=4.325
+ $Y=1.96 $X2=4.51 $Y2=2.105
r86 2 20 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=4.325
+ $Y=1.96 $X2=4.51 $Y2=2.815
r87 1 27 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=1.96 $X2=2.64 $Y2=2.105
r88 1 12 300 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=2 $X=2.495
+ $Y=1.96 $X2=2.64 $Y2=2.445
.ends

.subckt PM_SKY130_FD_SC_MS__OR4_4%A_591_392# 1 2 7 9 11 13 15
c28 15 0 1.09092e-19 $X=4 $Y=2.815
c29 9 0 1.55268e-19 $X=3.09 $Y=2.815
r30 13 20 3.14031 $w=2.8e-07 $l=1.41421e-07 $layer=LI1_cond $X=4.035 $Y=2.56
+ $X2=4 $Y2=2.435
r31 13 15 10.4955 $w=2.78e-07 $l=2.55e-07 $layer=LI1_cond $X=4.035 $Y=2.56
+ $X2=4.035 $Y2=2.815
r32 12 18 4.12165 $w=2e-07 $l=1.4e-07 $layer=LI1_cond $X=3.205 $Y=2.46 $X2=3.065
+ $Y2=2.46
r33 11 20 3.92538 $w=2e-07 $l=1.87083e-07 $layer=LI1_cond $X=3.825 $Y=2.46 $X2=4
+ $Y2=2.435
r34 11 12 34.3818 $w=1.98e-07 $l=6.2e-07 $layer=LI1_cond $X=3.825 $Y=2.46
+ $X2=3.205 $Y2=2.46
r35 7 18 2.94404 $w=2.8e-07 $l=1e-07 $layer=LI1_cond $X=3.065 $Y=2.56 $X2=3.065
+ $Y2=2.46
r36 7 9 10.4955 $w=2.78e-07 $l=2.55e-07 $layer=LI1_cond $X=3.065 $Y=2.56
+ $X2=3.065 $Y2=2.815
r37 2 20 600 $w=1.7e-07 $l=5.02295e-07 $layer=licon1_PDIFF $count=1 $X=3.855
+ $Y=1.96 $X2=4 $Y2=2.395
r38 2 15 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.855
+ $Y=1.96 $X2=4 $Y2=2.815
r39 1 18 600 $w=1.7e-07 $l=5.63471e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=1.96 $X2=3.09 $Y2=2.46
r40 1 9 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=1.96 $X2=3.09 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__OR4_4%A_965_392# 1 2 11
c13 11 0 1.75814e-19 $X=5.91 $Y=2.8
r14 8 11 37.0428 $w=2.78e-07 $l=9e-07 $layer=LI1_cond $X=5.01 $Y=2.84 $X2=5.91
+ $Y2=2.84
r15 2 11 600 $w=1.7e-07 $l=9.04986e-07 $layer=licon1_PDIFF $count=1 $X=5.775
+ $Y=1.96 $X2=5.91 $Y2=2.8
r16 1 8 600 $w=1.7e-07 $l=9.27901e-07 $layer=licon1_PDIFF $count=1 $X=4.825
+ $Y=1.96 $X2=5.01 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_MS__OR4_4%VGND 1 2 3 4 5 16 18 22 26 28 30 35 52 53 59
+ 62 66 75 78 84
c77 53 0 7.13014e-20 $X=6.48 $Y=0
r78 82 84 10.4353 $w=7.63e-07 $l=1.15e-07 $layer=LI1_cond $X=6 $Y=0.297
+ $X2=6.115 $Y2=0.297
r79 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r80 80 82 0.781751 $w=7.63e-07 $l=5e-08 $layer=LI1_cond $X=5.95 $Y=0.297 $X2=6
+ $Y2=0.297
r81 77 80 8.05203 $w=7.63e-07 $l=5.15e-07 $layer=LI1_cond $X=5.435 $Y=0.297
+ $X2=5.95 $Y2=0.297
r82 77 78 11.2171 $w=7.63e-07 $l=1.65e-07 $layer=LI1_cond $X=5.435 $Y=0.297
+ $X2=5.27 $Y2=0.297
r83 74 75 10.8372 $w=7.03e-07 $l=1.65e-07 $layer=LI1_cond $X=4.425 $Y=0.267
+ $X2=4.59 $Y2=0.267
r84 71 74 5.85315 $w=7.03e-07 $l=3.45e-07 $layer=LI1_cond $X=4.08 $Y=0.267
+ $X2=4.425 $Y2=0.267
r85 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r86 69 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r87 68 71 8.14351 $w=7.03e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=0.267
+ $X2=4.08 $Y2=0.267
r88 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r89 65 68 0.0848283 $w=7.03e-07 $l=5e-09 $layer=LI1_cond $X=3.595 $Y=0.267
+ $X2=3.6 $Y2=0.267
r90 65 66 10.8372 $w=7.03e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=0.267
+ $X2=3.43 $Y2=0.267
r91 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r92 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r93 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r94 53 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r95 52 84 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.48 $Y=0 $X2=6.115
+ $Y2=0
r96 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r97 49 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r98 49 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.08
+ $Y2=0
r99 48 78 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=5.27
+ $Y2=0
r100 48 75 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=4.59
+ $Y2=0
r101 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r102 44 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r103 43 66 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=3.43
+ $Y2=0
r104 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r105 41 62 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.74 $Y=0 $X2=2.56
+ $Y2=0
r106 41 43 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.74 $Y=0 $X2=3.12
+ $Y2=0
r107 39 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r108 39 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r109 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r110 36 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=0 $X2=1.28
+ $Y2=0
r111 36 38 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.445 $Y=0
+ $X2=2.16 $Y2=0
r112 35 62 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.38 $Y=0 $X2=2.56
+ $Y2=0
r113 35 38 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.38 $Y=0 $X2=2.16
+ $Y2=0
r114 34 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r115 34 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r116 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r117 31 56 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r118 31 33 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r119 30 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.28
+ $Y2=0
r120 30 33 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=0
+ $X2=0.72 $Y2=0
r121 28 69 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=3.6
+ $Y2=0
r122 28 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0
+ $X2=3.12 $Y2=0
r123 24 62 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=0.085
+ $X2=2.56 $Y2=0
r124 24 26 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.56 $Y=0.085
+ $X2=2.56 $Y2=0.455
r125 20 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0
r126 20 22 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.28 $Y=0.085
+ $X2=1.28 $Y2=0.58
r127 16 56 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r128 16 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.515
r129 5 80 182 $w=1.7e-07 $l=7.23878e-07 $layer=licon1_NDIFF $count=1 $X=5.295
+ $Y=0.37 $X2=5.95 $Y2=0.515
r130 5 77 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.295
+ $Y=0.37 $X2=5.435 $Y2=0.515
r131 4 74 121.333 $w=1.7e-07 $l=1.09167e-06 $layer=licon1_NDIFF $count=1
+ $X=3.375 $Y=0.37 $X2=4.425 $Y2=0.455
r132 4 65 121.333 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1
+ $X=3.375 $Y=0.37 $X2=3.595 $Y2=0.455
r133 3 26 182 $w=1.7e-07 $l=2.74226e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.37 $X2=2.56 $Y2=0.455
r134 2 22 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.28 $Y2=0.58
r135 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends


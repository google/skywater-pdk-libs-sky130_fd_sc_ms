* File: sky130_fd_sc_ms__o221ai_2.pex.spice
* Created: Wed Sep  2 12:23:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O221AI_2%C1 3 7 11 15 17 21 24
r43 23 24 58.8939 $w=3.11e-07 $l=3.8e-07 $layer=POLY_cond $X=0.545 $Y=1.465
+ $X2=0.925 $Y2=1.465
r44 22 23 7.7492 $w=3.11e-07 $l=5e-08 $layer=POLY_cond $X=0.495 $Y=1.465
+ $X2=0.545 $Y2=1.465
r45 20 22 34.8714 $w=3.11e-07 $l=2.25e-07 $layer=POLY_cond $X=0.27 $Y=1.465
+ $X2=0.495 $Y2=1.465
r46 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r47 17 21 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.27 $Y=1.665 $X2=0.27
+ $Y2=1.465
r48 13 24 10.8489 $w=3.11e-07 $l=7e-08 $layer=POLY_cond $X=0.995 $Y=1.465
+ $X2=0.925 $Y2=1.465
r49 13 15 314.855 $w=1.8e-07 $l=8.1e-07 $layer=POLY_cond $X=0.995 $Y=1.59
+ $X2=0.995 $Y2=2.4
r50 9 24 19.8172 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.3
+ $X2=0.925 $Y2=1.465
r51 9 11 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.925 $Y=1.3
+ $X2=0.925 $Y2=0.74
r52 5 23 15.5536 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.63
+ $X2=0.545 $Y2=1.465
r53 5 7 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.545 $Y=1.63
+ $X2=0.545 $Y2=2.4
r54 1 22 19.8172 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.465
r55 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O221AI_2%B1 1 3 5 7 10 14 16 20 21 23 24 25 43
c91 14 0 1.19923e-19 $X=3.33 $Y=0.795
c92 10 0 8.04709e-20 $X=3.255 $Y=2.4
c93 3 0 7.71556e-20 $X=1.805 $Y=2.4
c94 1 0 1.93102e-19 $X=1.805 $Y=1.68
r95 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.795
+ $Y=1.515 $X2=1.795 $Y2=1.515
r96 25 43 10.4716 $w=7.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.16 $Y=1.735
+ $X2=2.275 $Y2=1.735
r97 25 31 5.66972 $w=7.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.16 $Y=1.735
+ $X2=1.795 $Y2=1.735
r98 24 31 1.78635 $w=7.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=1.735
+ $X2=1.795 $Y2=1.735
r99 23 24 7.45607 $w=7.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.735
+ $X2=1.68 $Y2=1.735
r100 21 34 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.24 $Y=1.515
+ $X2=3.24 $Y2=1.68
r101 21 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.24 $Y=1.515
+ $X2=3.24 $Y2=1.35
r102 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.24
+ $Y=1.515 $X2=3.24 $Y2=1.515
r103 18 20 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=3.24 $Y=1.95
+ $X2=3.24 $Y2=1.515
r104 16 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.075 $Y=2.035
+ $X2=3.24 $Y2=1.95
r105 16 43 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=3.075 $Y=2.035
+ $X2=2.275 $Y2=2.035
r106 14 33 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.33 $Y=0.795
+ $X2=3.33 $Y2=1.35
r107 10 34 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.255 $Y=2.4
+ $X2=3.255 $Y2=1.68
r108 5 30 47.1698 $w=3.41e-07 $l=2.72489e-07 $layer=POLY_cond $X=1.915 $Y=1.29
+ $X2=1.81 $Y2=1.515
r109 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.915 $Y=1.29
+ $X2=1.915 $Y2=0.795
r110 1 30 34.0112 $w=3.41e-07 $l=1.67481e-07 $layer=POLY_cond $X=1.805 $Y=1.68
+ $X2=1.81 $Y2=1.515
r111 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.805 $Y=1.68
+ $X2=1.805 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O221AI_2%B2 1 3 6 8 10 14 16 22
c52 22 0 1.93102e-19 $X=2.685 $Y=1.515
c53 8 0 5.73497e-20 $X=2.755 $Y=1.68
r54 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.685
+ $Y=1.515 $X2=2.685 $Y2=1.515
r55 19 21 49.9634 $w=3.28e-07 $l=3.4e-07 $layer=POLY_cond $X=2.345 $Y=1.56
+ $X2=2.685 $Y2=1.56
r56 18 19 8.08232 $w=3.28e-07 $l=5.5e-08 $layer=POLY_cond $X=2.29 $Y=1.56
+ $X2=2.345 $Y2=1.56
r57 16 22 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.685 $Y=1.665
+ $X2=2.685 $Y2=1.515
r58 12 24 21.0783 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.775 $Y=1.35
+ $X2=2.775 $Y2=1.56
r59 12 14 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.775 $Y=1.35
+ $X2=2.775 $Y2=0.795
r60 8 24 2.93902 $w=3.28e-07 $l=2e-08 $layer=POLY_cond $X=2.755 $Y=1.56
+ $X2=2.775 $Y2=1.56
r61 8 21 10.2866 $w=3.28e-07 $l=7e-08 $layer=POLY_cond $X=2.755 $Y=1.56
+ $X2=2.685 $Y2=1.56
r62 8 10 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.755 $Y=1.68
+ $X2=2.755 $Y2=2.4
r63 4 19 21.0783 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.345 $Y=1.35
+ $X2=2.345 $Y2=1.56
r64 4 6 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.345 $Y=1.35
+ $X2=2.345 $Y2=0.795
r65 1 18 16.7902 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=2.29 $Y=1.77 $X2=2.29
+ $Y2=1.56
r66 1 3 168.7 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=2.29 $Y=1.77 $X2=2.29
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O221AI_2%A1 3 7 11 15 19 20 22 23 24 32 33
c87 7 0 1.76091e-19 $X=3.805 $Y=2.4
c88 3 0 2.04231e-19 $X=3.76 $Y=0.795
r89 32 35 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.28 $Y=1.515
+ $X2=5.28 $Y2=1.68
r90 32 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.28 $Y=1.515
+ $X2=5.28 $Y2=1.35
r91 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.28
+ $Y=1.515 $X2=5.28 $Y2=1.515
r92 24 41 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=5.28 $Y=1.665
+ $X2=5.28 $Y2=2.035
r93 24 33 2.52693 $w=7.08e-07 $l=1.5e-07 $layer=LI1_cond $X=5.28 $Y=1.665
+ $X2=5.28 $Y2=1.515
r94 22 41 9.41505 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=4.925 $Y=2.035
+ $X2=5.28 $Y2=2.035
r95 22 23 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=4.925 $Y=2.035
+ $X2=3.975 $Y2=2.035
r96 20 30 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.81 $Y=1.515
+ $X2=3.81 $Y2=1.68
r97 20 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.81 $Y=1.515
+ $X2=3.81 $Y2=1.35
r98 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.81
+ $Y=1.515 $X2=3.81 $Y2=1.515
r99 17 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.81 $Y=1.95
+ $X2=3.975 $Y2=2.035
r100 17 19 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=3.81 $Y=1.95
+ $X2=3.81 $Y2=1.515
r101 15 34 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=5.26 $Y=0.795
+ $X2=5.26 $Y2=1.35
r102 11 35 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.205 $Y=2.4
+ $X2=5.205 $Y2=1.68
r103 7 30 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.805 $Y=2.4
+ $X2=3.805 $Y2=1.68
r104 3 29 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.76 $Y=0.795
+ $X2=3.76 $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__O221AI_2%A2 3 7 11 15 17 24 26
c52 24 0 9.55934e-20 $X=4.51 $Y=1.515
r53 25 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.755 $Y=1.515
+ $X2=4.77 $Y2=1.515
r54 23 25 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=4.51 $Y=1.515
+ $X2=4.755 $Y2=1.515
r55 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.51
+ $Y=1.515 $X2=4.51 $Y2=1.515
r56 21 23 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=4.305 $Y=1.515
+ $X2=4.51 $Y2=1.515
r57 19 21 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.29 $Y=1.515
+ $X2=4.305 $Y2=1.515
r58 17 24 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.51 $Y=1.665
+ $X2=4.51 $Y2=1.515
r59 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=1.35
+ $X2=4.77 $Y2=1.515
r60 13 15 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=4.77 $Y=1.35
+ $X2=4.77 $Y2=0.795
r61 9 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.755 $Y=1.68
+ $X2=4.755 $Y2=1.515
r62 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.755 $Y=1.68
+ $X2=4.755 $Y2=2.4
r63 5 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.305 $Y=1.68
+ $X2=4.305 $Y2=1.515
r64 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.305 $Y=1.68
+ $X2=4.305 $Y2=2.4
r65 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.29 $Y=1.35
+ $X2=4.29 $Y2=1.515
r66 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=4.29 $Y=1.35 $X2=4.29
+ $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_MS__O221AI_2%VPWR 1 2 3 4 13 15 21 23 25 27 29 34 39 51
+ 60 64
r71 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r72 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r73 55 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r74 54 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r75 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r76 51 54 9.99847 $w=6.38e-07 $l=5.35e-07 $layer=LI1_cond $X=1.375 $Y=2.795
+ $X2=1.375 $Y2=3.33
r77 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r78 46 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r79 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r80 43 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r81 43 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r82 42 45 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=3.33 $X2=5.04
+ $Y2=3.33
r83 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r84 40 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.695 $Y=3.33
+ $X2=3.53 $Y2=3.33
r85 40 42 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.695 $Y=3.33
+ $X2=4.08 $Y2=3.33
r86 39 63 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.537 $Y2=3.33
r87 39 45 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.315 $Y=3.33
+ $X2=5.04 $Y2=3.33
r88 38 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r89 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r90 35 54 8.73481 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=1.695 $Y=3.33
+ $X2=1.375 $Y2=3.33
r91 35 37 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=1.695 $Y=3.33
+ $X2=3.12 $Y2=3.33
r92 34 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=3.33
+ $X2=3.53 $Y2=3.33
r93 34 37 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.365 $Y=3.33
+ $X2=3.12 $Y2=3.33
r94 33 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r95 33 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r96 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r97 30 48 3.96192 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=3.33
+ $X2=0.202 $Y2=3.33
r98 30 32 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.405 $Y=3.33
+ $X2=0.72 $Y2=3.33
r99 29 54 8.73481 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.375 $Y2=3.33
r100 29 32 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.72 $Y2=3.33
r101 27 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r102 27 57 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=1.68 $Y2=3.33
r103 23 63 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.48 $Y=3.245
+ $X2=5.537 $Y2=3.33
r104 23 25 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=5.48 $Y=3.245
+ $X2=5.48 $Y2=2.455
r105 19 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.53 $Y=3.245
+ $X2=3.53 $Y2=3.33
r106 19 21 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.53 $Y=3.245
+ $X2=3.53 $Y2=2.805
r107 15 18 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=0.28 $Y=2.115
+ $X2=0.28 $Y2=2.815
r108 13 48 3.18124 $w=2.5e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.202 $Y2=3.33
r109 13 18 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r110 4 25 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=5.295
+ $Y=1.84 $X2=5.48 $Y2=2.455
r111 3 21 600 $w=1.7e-07 $l=1.05345e-06 $layer=licon1_PDIFF $count=1 $X=3.345
+ $Y=1.84 $X2=3.53 $Y2=2.805
r112 2 51 300 $w=1.7e-07 $l=1.17675e-06 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=1.84 $X2=1.58 $Y2=2.795
r113 1 18 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.84 $X2=0.32 $Y2=2.815
r114 1 15 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.84 $X2=0.32 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__O221AI_2%Y 1 2 3 4 15 17 22 23 24 25 26 27 28 29
r60 28 37 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=2.375
+ $X2=0.74 $Y2=2.29
r61 28 49 3.58051 $w=2.6e-07 $l=8.9861e-08 $layer=LI1_cond $X=0.74 $Y=2.375
+ $X2=0.73 $Y2=2.46
r62 28 29 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=0.73 $Y=2.475 $X2=0.73
+ $Y2=2.775
r63 28 49 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=0.73 $Y=2.475
+ $X2=0.73 $Y2=2.46
r64 27 37 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.74 $Y=1.985
+ $X2=0.74 $Y2=2.29
r65 26 27 13.6586 $w=2.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.74 $Y=1.665
+ $X2=0.74 $Y2=1.985
r66 25 26 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.74 $Y=1.295
+ $X2=0.74 $Y2=1.665
r67 24 25 18.5671 $w=2.68e-07 $l=4.35e-07 $layer=LI1_cond $X=0.74 $Y=0.86
+ $X2=0.74 $Y2=1.295
r68 21 23 8.86124 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=2.53 $Y=2.512
+ $X2=2.695 $Y2=2.512
r69 21 22 8.86124 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=2.53 $Y=2.512
+ $X2=2.365 $Y2=2.512
r70 17 19 2.44 $w=2.5e-07 $l=5e-08 $layer=LI1_cond $X=4.49 $Y=2.46 $X2=4.49
+ $Y2=2.51
r71 15 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.365 $Y=2.375
+ $X2=4.49 $Y2=2.46
r72 15 23 108.952 $w=1.68e-07 $l=1.67e-06 $layer=LI1_cond $X=4.365 $Y=2.375
+ $X2=2.695 $Y2=2.375
r73 14 28 2.90867 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.875 $Y=2.375
+ $X2=0.74 $Y2=2.375
r74 14 22 97.2086 $w=1.68e-07 $l=1.49e-06 $layer=LI1_cond $X=0.875 $Y=2.375
+ $X2=2.365 $Y2=2.375
r75 4 19 600 $w=1.7e-07 $l=7.34405e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.84 $X2=4.53 $Y2=2.51
r76 3 21 600 $w=1.7e-07 $l=7.41215e-07 $layer=licon1_PDIFF $count=1 $X=2.38
+ $Y=1.84 $X2=2.53 $Y2=2.51
r77 2 28 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=0.635
+ $Y=1.84 $X2=0.77 $Y2=2.4
r78 2 27 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.635
+ $Y=1.84 $X2=0.77 $Y2=1.985
r79 1 24 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__O221AI_2%A_379_368# 1 2 7 10 15
c28 7 0 1.57627e-19 $X=2.865 $Y=2.99
r29 15 17 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=3.03 $Y=2.805
+ $X2=3.03 $Y2=2.99
r30 10 12 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.03 $Y=2.805
+ $X2=2.03 $Y2=2.99
r31 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=2.99
+ $X2=2.03 $Y2=2.99
r32 7 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.865 $Y=2.99
+ $X2=3.03 $Y2=2.99
r33 7 8 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.865 $Y=2.99
+ $X2=2.195 $Y2=2.99
r34 2 15 600 $w=1.7e-07 $l=1.05345e-06 $layer=licon1_PDIFF $count=1 $X=2.845
+ $Y=1.84 $X2=3.03 $Y2=2.805
r35 1 10 600 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=1.895
+ $Y=1.84 $X2=2.03 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_MS__O221AI_2%A_779_368# 1 2 7 11 14
c28 7 0 8.04979e-20 $X=4.815 $Y=2.99
r29 14 16 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=4.03 $Y=2.805
+ $X2=4.03 $Y2=2.99
r30 9 11 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.98 $Y=2.905
+ $X2=4.98 $Y2=2.455
r31 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.195 $Y=2.99
+ $X2=4.03 $Y2=2.99
r32 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.815 $Y=2.99
+ $X2=4.98 $Y2=2.905
r33 7 8 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.815 $Y=2.99
+ $X2=4.195 $Y2=2.99
r34 2 11 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=4.845
+ $Y=1.84 $X2=4.98 $Y2=2.455
r35 1 14 600 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=3.895
+ $Y=1.84 $X2=4.03 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_MS__O221AI_2%A_27_74# 1 2 3 4 15 17 18 22 23 24 27 29 33
+ 35
c51 35 0 5.73497e-20 $X=2.13 $Y=1.095
c52 33 0 1.48041e-19 $X=3.085 $Y=0.68
c53 29 0 5.61893e-20 $X=2.895 $Y=1.095
r54 31 33 9.87808 $w=3.83e-07 $l=3.3e-07 $layer=LI1_cond $X=3.087 $Y=1.01
+ $X2=3.087 $Y2=0.68
r55 30 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.215 $Y=1.095
+ $X2=2.13 $Y2=1.095
r56 29 31 8.24022 $w=1.7e-07 $l=2.30617e-07 $layer=LI1_cond $X=2.895 $Y=1.095
+ $X2=3.087 $Y2=1.01
r57 29 30 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.895 $Y=1.095
+ $X2=2.215 $Y2=1.095
r58 25 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.13 $Y=1.01 $X2=2.13
+ $Y2=1.095
r59 25 27 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.13 $Y=1.01
+ $X2=2.13 $Y2=0.885
r60 23 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=1.095
+ $X2=2.13 $Y2=1.095
r61 23 24 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.045 $Y=1.095
+ $X2=1.305 $Y2=1.095
r62 20 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.18 $Y=1.01
+ $X2=1.305 $Y2=1.095
r63 20 22 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.18 $Y=1.01
+ $X2=1.18 $Y2=0.515
r64 19 22 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.18 $Y=0.425 $X2=1.18
+ $Y2=0.515
r65 17 19 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.055 $Y=0.34
+ $X2=1.18 $Y2=0.425
r66 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.055 $Y=0.34
+ $X2=0.365 $Y2=0.34
r67 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.425
+ $X2=0.365 $Y2=0.34
r68 13 15 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.24 $Y=0.425 $X2=0.24
+ $Y2=0.515
r69 4 33 91 $w=1.7e-07 $l=3.53483e-07 $layer=licon1_NDIFF $count=2 $X=2.85
+ $Y=0.425 $X2=3.085 $Y2=0.68
r70 3 27 182 $w=1.7e-07 $l=5.25357e-07 $layer=licon1_NDIFF $count=1 $X=1.99
+ $Y=0.425 $X2=2.13 $Y2=0.885
r71 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1 $Y=0.37
+ $X2=1.14 $Y2=0.515
r72 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O221AI_2%A_311_85# 1 2 3 4 5 18 20 21 24 26 31 32 33
+ 36 38 42 44 45
c79 33 0 1.19923e-19 $X=3.71 $Y=1.095
r80 40 42 19.8853 $w=2.53e-07 $l=4.4e-07 $layer=LI1_cond $X=5.517 $Y=1.01
+ $X2=5.517 $Y2=0.57
r81 39 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.71 $Y=1.095
+ $X2=4.545 $Y2=1.095
r82 38 40 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=5.39 $Y=1.095
+ $X2=5.517 $Y2=1.01
r83 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.39 $Y=1.095
+ $X2=4.71 $Y2=1.095
r84 34 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.545 $Y=1.01
+ $X2=4.545 $Y2=1.095
r85 34 36 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=4.545 $Y=1.01
+ $X2=4.545 $Y2=0.57
r86 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.38 $Y=1.095
+ $X2=4.545 $Y2=1.095
r87 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.38 $Y=1.095
+ $X2=3.71 $Y2=1.095
r88 29 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.585 $Y=1.01
+ $X2=3.71 $Y2=1.095
r89 29 31 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=3.585 $Y=1.01
+ $X2=3.585 $Y2=0.57
r90 28 31 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=3.585 $Y=0.425
+ $X2=3.585 $Y2=0.57
r91 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=0.34
+ $X2=2.56 $Y2=0.34
r92 26 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.46 $Y=0.34
+ $X2=3.585 $Y2=0.425
r93 26 27 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=3.46 $Y=0.34
+ $X2=2.725 $Y2=0.34
r94 22 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=0.425
+ $X2=2.56 $Y2=0.34
r95 22 24 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.56 $Y=0.425
+ $X2=2.56 $Y2=0.655
r96 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=0.34
+ $X2=2.56 $Y2=0.34
r97 20 21 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.395 $Y=0.34
+ $X2=1.865 $Y2=0.34
r98 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.7 $Y=0.425
+ $X2=1.865 $Y2=0.34
r99 16 18 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.7 $Y=0.425 $X2=1.7
+ $Y2=0.655
r100 5 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.335
+ $Y=0.425 $X2=5.475 $Y2=0.57
r101 4 36 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=4.365
+ $Y=0.425 $X2=4.545 $Y2=0.57
r102 3 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.405
+ $Y=0.425 $X2=3.545 $Y2=0.57
r103 2 24 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=2.42
+ $Y=0.425 $X2=2.56 $Y2=0.655
r104 1 18 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.425 $X2=1.7 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_MS__O221AI_2%VGND 1 2 9 13 15 17 25 32 33 36 39
r52 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r53 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r54 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r55 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r56 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.21 $Y=0 $X2=5.045
+ $Y2=0
r57 30 32 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.21 $Y=0 $X2=5.52
+ $Y2=0
r58 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r59 29 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r60 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r61 26 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.045
+ $Y2=0
r62 26 28 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.56
+ $Y2=0
r63 25 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.88 $Y=0 $X2=5.045
+ $Y2=0
r64 25 28 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.88 $Y=0 $X2=4.56
+ $Y2=0
r65 24 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r66 23 24 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r67 19 23 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=3.6
+ $Y2=0
r68 19 20 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r69 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.88 $Y=0 $X2=4.045
+ $Y2=0
r70 17 23 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.88 $Y=0 $X2=3.6
+ $Y2=0
r71 15 24 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.6
+ $Y2=0
r72 15 20 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=0.24
+ $Y2=0
r73 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=0.085
+ $X2=5.045 $Y2=0
r74 11 13 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=5.045 $Y=0.085
+ $X2=5.045 $Y2=0.655
r75 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.045 $Y=0.085
+ $X2=4.045 $Y2=0
r76 7 9 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=4.045 $Y=0.085
+ $X2=4.045 $Y2=0.655
r77 2 13 182 $w=1.7e-07 $l=3.14484e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.425 $X2=5.045 $Y2=0.655
r78 1 9 182 $w=1.7e-07 $l=3.18119e-07 $layer=licon1_NDIFF $count=1 $X=3.835
+ $Y=0.425 $X2=4.045 $Y2=0.655
.ends


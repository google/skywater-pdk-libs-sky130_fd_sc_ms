* File: sky130_fd_sc_ms__o32ai_4.pex.spice
* Created: Fri Aug 28 18:04:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O32AI_4%B2 3 7 11 15 19 23 27 31 33 34 35 36 58
r84 57 58 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.855 $Y=1.515
+ $X2=1.87 $Y2=1.515
r85 55 57 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=1.6 $Y=1.515
+ $X2=1.855 $Y2=1.515
r86 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=1.515 $X2=1.6 $Y2=1.515
r87 53 55 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=1.425 $Y=1.515
+ $X2=1.6 $Y2=1.515
r88 52 53 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.405 $Y=1.515
+ $X2=1.425 $Y2=1.515
r89 51 56 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=1.26 $Y=1.605
+ $X2=1.6 $Y2=1.605
r90 50 52 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=1.26 $Y=1.515
+ $X2=1.405 $Y2=1.515
r91 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.26
+ $Y=1.515 $X2=1.26 $Y2=1.515
r92 48 50 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=0.955 $Y=1.515
+ $X2=1.26 $Y2=1.515
r93 47 48 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=0.925 $Y=1.515
+ $X2=0.955 $Y2=1.515
r94 45 47 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=0.92 $Y=1.515
+ $X2=0.925 $Y2=1.515
r95 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.92
+ $Y=1.515 $X2=0.92 $Y2=1.515
r96 43 45 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=0.505 $Y=1.515
+ $X2=0.92 $Y2=1.515
r97 41 43 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.515
+ $X2=0.505 $Y2=1.515
r98 36 56 2.63416 $w=3.48e-07 $l=8e-08 $layer=LI1_cond $X=1.68 $Y=1.605 $X2=1.6
+ $Y2=1.605
r99 35 51 1.97562 $w=3.48e-07 $l=6e-08 $layer=LI1_cond $X=1.2 $Y=1.605 $X2=1.26
+ $Y2=1.605
r100 35 46 9.21954 $w=3.48e-07 $l=2.8e-07 $layer=LI1_cond $X=1.2 $Y=1.605
+ $X2=0.92 $Y2=1.605
r101 34 46 6.58539 $w=3.48e-07 $l=2e-07 $layer=LI1_cond $X=0.72 $Y=1.605
+ $X2=0.92 $Y2=1.605
r102 33 34 15.8049 $w=3.48e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.605
+ $X2=0.72 $Y2=1.605
r103 29 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.87 $Y=1.35
+ $X2=1.87 $Y2=1.515
r104 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.87 $Y=1.35
+ $X2=1.87 $Y2=0.74
r105 25 57 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.68
+ $X2=1.855 $Y2=1.515
r106 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.855 $Y=1.68
+ $X2=1.855 $Y2=2.4
r107 21 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=1.515
r108 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.425 $Y2=0.74
r109 17 52 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.68
+ $X2=1.405 $Y2=1.515
r110 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.405 $Y=1.68
+ $X2=1.405 $Y2=2.4
r111 13 48 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.68
+ $X2=0.955 $Y2=1.515
r112 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.955 $Y=1.68
+ $X2=0.955 $Y2=2.4
r113 9 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=1.515
r114 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=0.74
r115 5 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.515
r116 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
r117 1 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.68
+ $X2=0.505 $Y2=1.515
r118 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.505 $Y=1.68
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_4%B1 3 7 11 15 19 23 27 31 33 34 35 36 37 63
r97 61 63 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=3.74 $Y=1.515
+ $X2=3.855 $Y2=1.515
r98 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.74
+ $Y=1.515 $X2=3.74 $Y2=1.515
r99 59 61 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.665 $Y=1.515
+ $X2=3.74 $Y2=1.515
r100 57 59 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=3.4 $Y=1.515
+ $X2=3.665 $Y2=1.515
r101 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.4
+ $Y=1.515 $X2=3.4 $Y2=1.515
r102 55 57 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=3.355 $Y=1.515
+ $X2=3.4 $Y2=1.515
r103 54 55 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=3.205 $Y=1.515
+ $X2=3.355 $Y2=1.515
r104 52 54 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=3.06 $Y=1.515
+ $X2=3.205 $Y2=1.515
r105 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.06
+ $Y=1.515 $X2=3.06 $Y2=1.515
r106 50 52 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=2.855 $Y=1.515
+ $X2=3.06 $Y2=1.515
r107 49 50 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=2.755 $Y=1.515
+ $X2=2.855 $Y2=1.515
r108 48 53 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=2.72 $Y=1.605
+ $X2=3.06 $Y2=1.605
r109 47 49 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=2.72 $Y=1.515
+ $X2=2.755 $Y2=1.515
r110 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.72
+ $Y=1.515 $X2=2.72 $Y2=1.515
r111 45 47 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=2.355 $Y=1.515
+ $X2=2.72 $Y2=1.515
r112 43 45 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=2.305 $Y=1.515
+ $X2=2.355 $Y2=1.515
r113 37 62 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=4.08 $Y=1.605
+ $X2=3.74 $Y2=1.605
r114 36 62 4.60977 $w=3.48e-07 $l=1.4e-07 $layer=LI1_cond $X=3.6 $Y=1.605
+ $X2=3.74 $Y2=1.605
r115 36 58 6.58539 $w=3.48e-07 $l=2e-07 $layer=LI1_cond $X=3.6 $Y=1.605 $X2=3.4
+ $Y2=1.605
r116 35 58 9.21954 $w=3.48e-07 $l=2.8e-07 $layer=LI1_cond $X=3.12 $Y=1.605
+ $X2=3.4 $Y2=1.605
r117 35 53 1.97562 $w=3.48e-07 $l=6e-08 $layer=LI1_cond $X=3.12 $Y=1.605
+ $X2=3.06 $Y2=1.605
r118 34 48 2.63416 $w=3.48e-07 $l=8e-08 $layer=LI1_cond $X=2.64 $Y=1.605
+ $X2=2.72 $Y2=1.605
r119 33 34 15.8049 $w=3.48e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.605
+ $X2=2.64 $Y2=1.605
r120 29 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.855 $Y=1.35
+ $X2=3.855 $Y2=1.515
r121 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.855 $Y=1.35
+ $X2=3.855 $Y2=0.74
r122 25 59 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.665 $Y=1.68
+ $X2=3.665 $Y2=1.515
r123 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.665 $Y=1.68
+ $X2=3.665 $Y2=2.4
r124 21 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.355 $Y=1.35
+ $X2=3.355 $Y2=1.515
r125 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.355 $Y=1.35
+ $X2=3.355 $Y2=0.74
r126 17 54 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=1.68
+ $X2=3.205 $Y2=1.515
r127 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.205 $Y=1.68
+ $X2=3.205 $Y2=2.4
r128 13 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.855 $Y=1.35
+ $X2=2.855 $Y2=1.515
r129 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.855 $Y=1.35
+ $X2=2.855 $Y2=0.74
r130 9 49 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.755 $Y=1.68
+ $X2=2.755 $Y2=1.515
r131 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.755 $Y=1.68
+ $X2=2.755 $Y2=2.4
r132 5 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.355 $Y=1.35
+ $X2=2.355 $Y2=1.515
r133 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.355 $Y=1.35
+ $X2=2.355 $Y2=0.74
r134 1 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=1.68
+ $X2=2.305 $Y2=1.515
r135 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.305 $Y=1.68
+ $X2=2.305 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_4%A3 3 5 6 9 13 17 21 25 29 33 35 36 37 52
c96 9 0 1.72955e-19 $X=4.675 $Y=2.4
r97 51 52 46.6452 $w=3.1e-07 $l=3e-07 $layer=POLY_cond $X=5.575 $Y=1.515
+ $X2=5.875 $Y2=1.515
r98 50 51 20.9903 $w=3.1e-07 $l=1.35e-07 $layer=POLY_cond $X=5.44 $Y=1.515
+ $X2=5.575 $Y2=1.515
r99 48 50 1.55484 $w=3.1e-07 $l=1e-08 $layer=POLY_cond $X=5.43 $Y=1.515 $X2=5.44
+ $Y2=1.515
r100 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.43
+ $Y=1.515 $X2=5.43 $Y2=1.515
r101 46 48 47.4226 $w=3.1e-07 $l=3.05e-07 $layer=POLY_cond $X=5.125 $Y=1.515
+ $X2=5.43 $Y2=1.515
r102 45 49 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=5.09 $Y=1.605
+ $X2=5.43 $Y2=1.605
r103 44 46 5.44194 $w=3.1e-07 $l=3.5e-08 $layer=POLY_cond $X=5.09 $Y=1.515
+ $X2=5.125 $Y2=1.515
r104 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.09
+ $Y=1.515 $X2=5.09 $Y2=1.515
r105 42 44 22.5452 $w=3.1e-07 $l=1.45e-07 $layer=POLY_cond $X=4.945 $Y=1.515
+ $X2=5.09 $Y2=1.515
r106 41 42 41.9806 $w=3.1e-07 $l=2.7e-07 $layer=POLY_cond $X=4.675 $Y=1.515
+ $X2=4.945 $Y2=1.515
r107 37 49 2.96342 $w=3.48e-07 $l=9e-08 $layer=LI1_cond $X=5.52 $Y=1.605
+ $X2=5.43 $Y2=1.605
r108 36 45 1.64635 $w=3.48e-07 $l=5e-08 $layer=LI1_cond $X=5.04 $Y=1.605
+ $X2=5.09 $Y2=1.605
r109 35 36 15.8049 $w=3.48e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.605
+ $X2=5.04 $Y2=1.605
r110 31 52 23.3226 $w=3.1e-07 $l=2.2798e-07 $layer=POLY_cond $X=6.025 $Y=1.68
+ $X2=5.875 $Y2=1.515
r111 31 33 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.025 $Y=1.68
+ $X2=6.025 $Y2=2.4
r112 27 52 19.7411 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.875 $Y=1.35
+ $X2=5.875 $Y2=1.515
r113 27 29 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.875 $Y=1.35
+ $X2=5.875 $Y2=0.74
r114 23 51 15.4789 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.575 $Y=1.68
+ $X2=5.575 $Y2=1.515
r115 23 25 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.575 $Y=1.68
+ $X2=5.575 $Y2=2.4
r116 19 50 19.7411 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.44 $Y=1.35
+ $X2=5.44 $Y2=1.515
r117 19 21 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.44 $Y=1.35
+ $X2=5.44 $Y2=0.74
r118 15 46 15.4789 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.125 $Y=1.68
+ $X2=5.125 $Y2=1.515
r119 15 17 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.125 $Y=1.68
+ $X2=5.125 $Y2=2.4
r120 11 42 19.7411 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.945 $Y=1.35
+ $X2=4.945 $Y2=1.515
r121 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.945 $Y=1.35
+ $X2=4.945 $Y2=0.74
r122 7 41 15.4789 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.675 $Y=1.68
+ $X2=4.675 $Y2=1.515
r123 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.675 $Y=1.68
+ $X2=4.675 $Y2=2.4
r124 5 41 26.8705 $w=3.1e-07 $l=1.27279e-07 $layer=POLY_cond $X=4.585 $Y=1.425
+ $X2=4.675 $Y2=1.515
r125 5 6 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=4.585 $Y=1.425
+ $X2=4.43 $Y2=1.425
r126 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.355 $Y=1.35
+ $X2=4.43 $Y2=1.425
r127 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.355 $Y=1.35
+ $X2=4.355 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_4%A2 1 3 6 10 14 18 22 26 30 32 33 34 35 36 53
r97 53 55 36.1862 $w=3.33e-07 $l=2.5e-07 $layer=POLY_cond $X=8.04 $Y=1.56
+ $X2=8.29 $Y2=1.56
r98 53 54 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=8.04
+ $Y=1.515 $X2=8.04 $Y2=1.515
r99 44 46 5.78979 $w=3.33e-07 $l=4e-08 $layer=POLY_cond $X=6.68 $Y=1.56 $X2=6.72
+ $Y2=1.56
r100 44 45 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=6.68
+ $Y=1.515 $X2=6.68 $Y2=1.515
r101 42 44 15.1982 $w=3.33e-07 $l=1.05e-07 $layer=POLY_cond $X=6.575 $Y=1.56
+ $X2=6.68 $Y2=1.56
r102 36 54 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=8.4 $Y=1.565
+ $X2=8.04 $Y2=1.565
r103 35 54 3.21612 $w=4.28e-07 $l=1.2e-07 $layer=LI1_cond $X=7.92 $Y=1.565
+ $X2=8.04 $Y2=1.565
r104 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.92 $Y2=1.565
r105 33 34 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.44 $Y2=1.565
r106 33 45 7.50428 $w=4.28e-07 $l=2.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=6.68 $Y2=1.565
r107 32 45 5.3602 $w=4.28e-07 $l=2e-07 $layer=LI1_cond $X=6.48 $Y=1.565 $X2=6.68
+ $Y2=1.565
r108 28 55 21.4384 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=8.29 $Y=1.35
+ $X2=8.29 $Y2=1.56
r109 28 30 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.29 $Y=1.35
+ $X2=8.29 $Y2=0.74
r110 24 53 2.17117 $w=3.33e-07 $l=1.5e-08 $layer=POLY_cond $X=8.025 $Y=1.56
+ $X2=8.04 $Y2=1.56
r111 24 50 44.1471 $w=3.33e-07 $l=3.05e-07 $layer=POLY_cond $X=8.025 $Y=1.56
+ $X2=7.72 $Y2=1.56
r112 24 26 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.025 $Y=1.68
+ $X2=8.025 $Y2=2.4
r113 20 50 21.4384 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.72 $Y=1.35
+ $X2=7.72 $Y2=1.56
r114 20 22 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.72 $Y=1.35
+ $X2=7.72 $Y2=0.74
r115 16 50 28.2252 $w=3.33e-07 $l=1.95e-07 $layer=POLY_cond $X=7.525 $Y=1.56
+ $X2=7.72 $Y2=1.56
r116 16 48 34.015 $w=3.33e-07 $l=2.35e-07 $layer=POLY_cond $X=7.525 $Y=1.56
+ $X2=7.29 $Y2=1.56
r117 16 18 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.525 $Y=1.68
+ $X2=7.525 $Y2=2.4
r118 12 48 21.4384 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.29 $Y=1.35
+ $X2=7.29 $Y2=1.56
r119 12 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.29 $Y=1.35
+ $X2=7.29 $Y2=0.74
r120 8 48 38.3574 $w=3.33e-07 $l=2.65e-07 $layer=POLY_cond $X=7.025 $Y=1.56
+ $X2=7.29 $Y2=1.56
r121 8 46 44.1471 $w=3.33e-07 $l=3.05e-07 $layer=POLY_cond $X=7.025 $Y=1.56
+ $X2=6.72 $Y2=1.56
r122 8 10 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.025 $Y=1.68
+ $X2=7.025 $Y2=2.4
r123 4 46 21.4384 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.72 $Y=1.35
+ $X2=6.72 $Y2=1.56
r124 4 6 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.72 $Y=1.35 $X2=6.72
+ $Y2=0.74
r125 1 42 17.1428 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=6.575 $Y=1.77
+ $X2=6.575 $Y2=1.56
r126 1 3 168.7 $w=1.8e-07 $l=6.3e-07 $layer=POLY_cond $X=6.575 $Y=1.77 $X2=6.575
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_4%A1 3 7 11 15 19 23 27 31 33 34 35 36 37 55
r83 54 55 21.8356 $w=2.98e-07 $l=1.35e-07 $layer=POLY_cond $X=10.085 $Y=1.515
+ $X2=10.22 $Y2=1.515
r84 52 54 21.8356 $w=2.98e-07 $l=1.35e-07 $layer=POLY_cond $X=9.95 $Y=1.515
+ $X2=10.085 $Y2=1.515
r85 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.95
+ $Y=1.515 $X2=9.95 $Y2=1.515
r86 50 52 37.2013 $w=2.98e-07 $l=2.3e-07 $layer=POLY_cond $X=9.72 $Y=1.515
+ $X2=9.95 $Y2=1.515
r87 49 50 29.9228 $w=2.98e-07 $l=1.85e-07 $layer=POLY_cond $X=9.535 $Y=1.515
+ $X2=9.72 $Y2=1.515
r88 48 49 39.6275 $w=2.98e-07 $l=2.45e-07 $layer=POLY_cond $X=9.29 $Y=1.515
+ $X2=9.535 $Y2=1.515
r89 46 48 3.2349 $w=2.98e-07 $l=2e-08 $layer=POLY_cond $X=9.27 $Y=1.515 $X2=9.29
+ $Y2=1.515
r90 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.27
+ $Y=1.515 $X2=9.27 $Y2=1.515
r91 44 46 29.9228 $w=2.98e-07 $l=1.85e-07 $layer=POLY_cond $X=9.085 $Y=1.515
+ $X2=9.27 $Y2=1.515
r92 43 44 47.7148 $w=2.98e-07 $l=2.95e-07 $layer=POLY_cond $X=8.79 $Y=1.515
+ $X2=9.085 $Y2=1.515
r93 36 37 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=10.32 $Y=1.565
+ $X2=10.8 $Y2=1.565
r94 36 53 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.32 $Y=1.565
+ $X2=9.95 $Y2=1.565
r95 35 53 2.94811 $w=4.28e-07 $l=1.1e-07 $layer=LI1_cond $X=9.84 $Y=1.565
+ $X2=9.95 $Y2=1.565
r96 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=9.36 $Y=1.565
+ $X2=9.84 $Y2=1.565
r97 34 47 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=9.36 $Y=1.565 $X2=9.27
+ $Y2=1.565
r98 33 47 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=8.88 $Y=1.565
+ $X2=9.27 $Y2=1.565
r99 29 55 50.9497 $w=2.98e-07 $l=3.88844e-07 $layer=POLY_cond $X=10.535 $Y=1.68
+ $X2=10.22 $Y2=1.515
r100 29 31 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=10.535 $Y=1.68
+ $X2=10.535 $Y2=2.4
r101 25 55 18.8112 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.22 $Y=1.35
+ $X2=10.22 $Y2=1.515
r102 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=10.22 $Y=1.35
+ $X2=10.22 $Y2=0.74
r103 21 54 14.565 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.085 $Y=1.68
+ $X2=10.085 $Y2=1.515
r104 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=10.085 $Y=1.68
+ $X2=10.085 $Y2=2.4
r105 17 50 18.8112 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.72 $Y=1.35
+ $X2=9.72 $Y2=1.515
r106 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.72 $Y=1.35
+ $X2=9.72 $Y2=0.74
r107 13 49 14.565 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.535 $Y=1.68
+ $X2=9.535 $Y2=1.515
r108 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=9.535 $Y=1.68
+ $X2=9.535 $Y2=2.4
r109 9 48 18.8112 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.29 $Y=1.35
+ $X2=9.29 $Y2=1.515
r110 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.29 $Y=1.35
+ $X2=9.29 $Y2=0.74
r111 5 44 14.565 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.085 $Y=1.68
+ $X2=9.085 $Y2=1.515
r112 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=9.085 $Y=1.68
+ $X2=9.085 $Y2=2.4
r113 1 43 18.8112 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.79 $Y=1.35
+ $X2=8.79 $Y2=1.515
r114 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.79 $Y=1.35 $X2=8.79
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_4%A_27_368# 1 2 3 4 5 18 22 23 26 28 30 31 32
+ 36 40 44 46
c68 46 0 1.72955e-19 $X=3.89 $Y=2.455
r69 37 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.145 $Y=2.375
+ $X2=2.98 $Y2=2.375
r70 36 46 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.725 $Y=2.375
+ $X2=3.89 $Y2=2.375
r71 36 37 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.725 $Y=2.375
+ $X2=3.145 $Y2=2.375
r72 33 42 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.245 $Y=2.375
+ $X2=2.12 $Y2=2.375
r73 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=2.375
+ $X2=2.98 $Y2=2.375
r74 32 33 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.815 $Y=2.375
+ $X2=2.245 $Y2=2.375
r75 30 42 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=2.46 $X2=2.12
+ $Y2=2.375
r76 30 31 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=2.12 $Y=2.46
+ $X2=2.12 $Y2=2.905
r77 29 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.265 $Y=2.99
+ $X2=1.14 $Y2=2.99
r78 28 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.995 $Y=2.99
+ $X2=2.12 $Y2=2.905
r79 28 29 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.995 $Y=2.99
+ $X2=1.265 $Y2=2.99
r80 24 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=2.905
+ $X2=1.14 $Y2=2.99
r81 24 26 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=1.14 $Y=2.905
+ $X2=1.14 $Y2=2.455
r82 22 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.015 $Y=2.99
+ $X2=1.14 $Y2=2.99
r83 22 23 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.015 $Y=2.99
+ $X2=0.445 $Y2=2.99
r84 18 21 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.28 $Y=2.115 $X2=0.28
+ $Y2=2.815
r85 16 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.445 $Y2=2.99
r86 16 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=2.905 $X2=0.28
+ $Y2=2.815
r87 5 46 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=3.755
+ $Y=1.84 $X2=3.89 $Y2=2.455
r88 4 44 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=2.845
+ $Y=1.84 $X2=2.98 $Y2=2.455
r89 3 42 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.945
+ $Y=1.84 $X2=2.08 $Y2=2.455
r90 2 26 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.455
r91 1 21 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r92 1 18 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_4%Y 1 2 3 4 5 6 7 8 27 31 33 34 37 39 41 45 47
+ 51 53 57 62 64 67 68 69 70 72 74 75
r158 65 75 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.63 $Y=2.12
+ $X2=1.63 $Y2=2.405
r159 65 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=2.12
+ $X2=1.63 $Y2=2.035
r160 62 74 3.70735 $w=2.5e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.89 $Y=1.95
+ $X2=5.805 $Y2=2.035
r161 61 62 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.89 $Y=1.26
+ $X2=5.89 $Y2=1.95
r162 58 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.065 $Y=2.035
+ $X2=4.9 $Y2=2.035
r163 57 74 2.76166 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.635 $Y=2.035
+ $X2=5.805 $Y2=2.035
r164 57 58 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.635 $Y=2.035
+ $X2=5.065 $Y2=2.035
r165 54 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.805 $Y=1.175
+ $X2=3.64 $Y2=1.175
r166 53 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.805 $Y=1.175
+ $X2=5.89 $Y2=1.26
r167 53 54 130.481 $w=1.68e-07 $l=2e-06 $layer=LI1_cond $X=5.805 $Y=1.175
+ $X2=3.805 $Y2=1.175
r168 49 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=1.09
+ $X2=3.64 $Y2=1.175
r169 49 51 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=3.64 $Y=1.09
+ $X2=3.64 $Y2=0.86
r170 48 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=1.175
+ $X2=2.64 $Y2=1.175
r171 47 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.475 $Y=1.175
+ $X2=3.64 $Y2=1.175
r172 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.475 $Y=1.175
+ $X2=2.805 $Y2=1.175
r173 43 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=1.09
+ $X2=2.64 $Y2=1.175
r174 43 45 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.64 $Y=1.09
+ $X2=2.64 $Y2=0.86
r175 42 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.805 $Y=1.175
+ $X2=1.68 $Y2=1.175
r176 41 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=1.175
+ $X2=2.64 $Y2=1.175
r177 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.475 $Y=1.175
+ $X2=1.805 $Y2=1.175
r178 40 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=2.035
+ $X2=1.63 $Y2=2.035
r179 39 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.735 $Y=2.035
+ $X2=4.9 $Y2=2.035
r180 39 40 191.807 $w=1.68e-07 $l=2.94e-06 $layer=LI1_cond $X=4.735 $Y=2.035
+ $X2=1.795 $Y2=2.035
r181 35 68 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=1.09
+ $X2=1.68 $Y2=1.175
r182 35 37 10.6025 $w=2.48e-07 $l=2.3e-07 $layer=LI1_cond $X=1.68 $Y=1.09
+ $X2=1.68 $Y2=0.86
r183 33 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.555 $Y=1.175
+ $X2=1.68 $Y2=1.175
r184 33 34 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.555 $Y=1.175
+ $X2=0.875 $Y2=1.175
r185 32 64 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=2.035
+ $X2=0.73 $Y2=2.035
r186 31 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=2.035
+ $X2=1.63 $Y2=2.035
r187 31 32 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.465 $Y=2.035
+ $X2=0.815 $Y2=2.035
r188 25 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.71 $Y=1.09
+ $X2=0.875 $Y2=1.175
r189 25 27 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.71 $Y=1.09
+ $X2=0.71 $Y2=0.86
r190 8 74 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=5.665
+ $Y=1.84 $X2=5.8 $Y2=2.115
r191 7 72 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=4.765
+ $Y=1.84 $X2=4.9 $Y2=2.115
r192 6 67 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.84 $X2=1.63 $Y2=2.115
r193 5 64 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.115
r194 4 51 182 $w=1.7e-07 $l=5.85662e-07 $layer=licon1_NDIFF $count=1 $X=3.43
+ $Y=0.37 $X2=3.64 $Y2=0.86
r195 3 45 182 $w=1.7e-07 $l=5.85662e-07 $layer=licon1_NDIFF $count=1 $X=2.43
+ $Y=0.37 $X2=2.64 $Y2=0.86
r196 2 37 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.64 $Y2=0.86
r197 1 27 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_4%VPWR 1 2 3 4 5 18 22 26 30 32 34 39 40 42 43
+ 45 46 47 65 69 75 79
r119 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r120 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r121 73 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r122 73 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r123 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r124 70 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.975 $Y=3.33
+ $X2=9.81 $Y2=3.33
r125 70 72 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.975 $Y=3.33
+ $X2=10.32 $Y2=3.33
r126 69 78 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=10.675 $Y=3.33
+ $X2=10.857 $Y2=3.33
r127 69 72 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=10.675 $Y=3.33
+ $X2=10.32 $Y2=3.33
r128 68 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r129 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r130 65 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.645 $Y=3.33
+ $X2=9.81 $Y2=3.33
r131 65 67 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.645 $Y=3.33
+ $X2=9.36 $Y2=3.33
r132 64 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r133 63 64 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r134 60 63 313.155 $w=1.68e-07 $l=4.8e-06 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=8.4
+ $Y2=3.33
r135 60 61 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r136 58 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r137 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r138 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r139 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r140 51 55 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r141 50 54 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r142 50 51 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r143 47 64 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=8.4 $Y2=3.33
r144 47 61 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=3.6 $Y2=3.33
r145 45 63 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.695 $Y=3.33
+ $X2=8.4 $Y2=3.33
r146 45 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.695 $Y=3.33
+ $X2=8.82 $Y2=3.33
r147 44 67 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=8.945 $Y=3.33
+ $X2=9.36 $Y2=3.33
r148 44 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.945 $Y=3.33
+ $X2=8.82 $Y2=3.33
r149 42 57 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.345 $Y=3.33
+ $X2=3.12 $Y2=3.33
r150 42 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.345 $Y=3.33
+ $X2=3.43 $Y2=3.33
r151 41 60 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=3.33
+ $X2=3.6 $Y2=3.33
r152 41 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=3.33
+ $X2=3.43 $Y2=3.33
r153 39 54 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=2.16 $Y2=3.33
r154 39 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=2.53 $Y2=3.33
r155 38 57 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.615 $Y=3.33
+ $X2=3.12 $Y2=3.33
r156 38 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=3.33
+ $X2=2.53 $Y2=3.33
r157 34 37 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=10.8 $Y=2.115
+ $X2=10.8 $Y2=2.815
r158 32 78 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.8 $Y=3.245
+ $X2=10.857 $Y2=3.33
r159 32 37 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.8 $Y=3.245
+ $X2=10.8 $Y2=2.815
r160 28 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.81 $Y=3.245
+ $X2=9.81 $Y2=3.33
r161 28 30 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=9.81 $Y=3.245
+ $X2=9.81 $Y2=2.455
r162 24 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.82 $Y=3.245
+ $X2=8.82 $Y2=3.33
r163 24 26 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=8.82 $Y=3.245
+ $X2=8.82 $Y2=2.455
r164 20 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=3.245
+ $X2=3.43 $Y2=3.33
r165 20 22 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.43 $Y=3.245
+ $X2=3.43 $Y2=2.805
r166 16 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=3.245
+ $X2=2.53 $Y2=3.33
r167 16 18 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.53 $Y=3.245
+ $X2=2.53 $Y2=2.805
r168 5 37 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.625
+ $Y=1.84 $X2=10.76 $Y2=2.815
r169 5 34 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=10.625
+ $Y=1.84 $X2=10.76 $Y2=2.115
r170 4 30 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=9.625
+ $Y=1.84 $X2=9.81 $Y2=2.455
r171 3 26 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=8.715
+ $Y=1.84 $X2=8.86 $Y2=2.455
r172 2 22 600 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=3.295
+ $Y=1.84 $X2=3.43 $Y2=2.805
r173 1 18 600 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=2.395
+ $Y=1.84 $X2=2.53 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_4%A_861_368# 1 2 3 4 5 18 20 21 24 26 30 34 38
+ 40 44 46 47 48
r59 42 44 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=8.3 $Y=2.905 $X2=8.3
+ $Y2=2.455
r60 41 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.465 $Y=2.99
+ $X2=7.3 $Y2=2.99
r61 40 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.135 $Y=2.99
+ $X2=8.3 $Y2=2.905
r62 40 41 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.135 $Y=2.99
+ $X2=7.465 $Y2=2.99
r63 36 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.3 $Y=2.905 $X2=7.3
+ $Y2=2.99
r64 36 38 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=7.3 $Y=2.905 $X2=7.3
+ $Y2=2.455
r65 35 47 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=6.465 $Y=2.99
+ $X2=6.305 $Y2=2.99
r66 34 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.135 $Y=2.99
+ $X2=7.3 $Y2=2.99
r67 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.135 $Y=2.99
+ $X2=6.465 $Y2=2.99
r68 30 33 25.2097 $w=3.18e-07 $l=7e-07 $layer=LI1_cond $X=6.305 $Y=2.115
+ $X2=6.305 $Y2=2.815
r69 28 47 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=6.305 $Y=2.905
+ $X2=6.305 $Y2=2.99
r70 28 33 3.24125 $w=3.18e-07 $l=9e-08 $layer=LI1_cond $X=6.305 $Y=2.905
+ $X2=6.305 $Y2=2.815
r71 27 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.435 $Y=2.99
+ $X2=5.35 $Y2=2.99
r72 26 47 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=6.145 $Y=2.99
+ $X2=6.305 $Y2=2.99
r73 26 27 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=6.145 $Y=2.99
+ $X2=5.435 $Y2=2.99
r74 22 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.35 $Y=2.905
+ $X2=5.35 $Y2=2.99
r75 22 24 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=5.35 $Y=2.905
+ $X2=5.35 $Y2=2.455
r76 20 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.265 $Y=2.99
+ $X2=5.35 $Y2=2.99
r77 20 21 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.265 $Y=2.99
+ $X2=4.535 $Y2=2.99
r78 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.41 $Y=2.905
+ $X2=4.535 $Y2=2.99
r79 16 18 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=4.41 $Y=2.905
+ $X2=4.41 $Y2=2.455
r80 5 44 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=8.115
+ $Y=1.84 $X2=8.3 $Y2=2.455
r81 4 38 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=7.115
+ $Y=1.84 $X2=7.3 $Y2=2.455
r82 3 33 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=6.115
+ $Y=1.84 $X2=6.3 $Y2=2.815
r83 3 30 400 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=1 $X=6.115
+ $Y=1.84 $X2=6.3 $Y2=2.115
r84 2 24 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=5.215
+ $Y=1.84 $X2=5.35 $Y2=2.455
r85 1 18 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=4.305
+ $Y=1.84 $X2=4.45 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_4%A_1333_368# 1 2 3 4 15 19 23 25 27 29 32 34
+ 36
r59 27 38 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.31 $Y=2.12
+ $X2=10.31 $Y2=2.035
r60 27 29 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=10.31 $Y=2.12
+ $X2=10.31 $Y2=2.815
r61 26 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.475 $Y=2.035
+ $X2=9.31 $Y2=2.035
r62 25 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.145 $Y=2.035
+ $X2=10.31 $Y2=2.035
r63 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.145 $Y=2.035
+ $X2=9.475 $Y2=2.035
r64 21 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.31 $Y=2.12 $X2=9.31
+ $Y2=2.035
r65 21 23 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=9.31 $Y=2.12
+ $X2=9.31 $Y2=2.815
r66 20 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.965 $Y=2.035
+ $X2=7.8 $Y2=2.035
r67 19 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.145 $Y=2.035
+ $X2=9.31 $Y2=2.035
r68 19 20 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=9.145 $Y=2.035
+ $X2=7.965 $Y2=2.035
r69 16 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.965 $Y=2.035
+ $X2=6.8 $Y2=2.035
r70 15 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.635 $Y=2.035
+ $X2=7.8 $Y2=2.035
r71 15 16 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.635 $Y=2.035
+ $X2=6.965 $Y2=2.035
r72 4 38 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=10.175
+ $Y=1.84 $X2=10.31 $Y2=2.115
r73 4 29 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.175
+ $Y=1.84 $X2=10.31 $Y2=2.815
r74 3 36 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=9.175
+ $Y=1.84 $X2=9.31 $Y2=2.115
r75 3 23 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.175
+ $Y=1.84 $X2=9.31 $Y2=2.815
r76 2 34 300 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=2 $X=7.615
+ $Y=1.84 $X2=7.8 $Y2=2.115
r77 1 32 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=6.665
+ $Y=1.84 $X2=6.8 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_4%A_27_74# 1 2 3 4 5 6 7 8 9 10 11 36 38 39 42
+ 44 48 50 54 56 61 62 63 66 68 70 74 76 80 82 86 88 92 94 95 96 98 102 104 105
+ 106
r184 102 103 4.15909 $w=5.72e-07 $l=1.95e-07 $layer=LI1_cond $X=6.332 $Y=0.9
+ $X2=6.332 $Y2=1.095
r185 100 102 1.38636 $w=5.72e-07 $l=6.5e-08 $layer=LI1_cond $X=6.332 $Y=0.835
+ $X2=6.332 $Y2=0.9
r186 90 92 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.505 $Y=1.01
+ $X2=10.505 $Y2=0.515
r187 89 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.67 $Y=1.095
+ $X2=9.505 $Y2=1.095
r188 88 90 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.34 $Y=1.095
+ $X2=10.505 $Y2=1.01
r189 88 89 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.34 $Y=1.095
+ $X2=9.67 $Y2=1.095
r190 84 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.505 $Y=1.01
+ $X2=9.505 $Y2=1.095
r191 84 86 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=9.505 $Y=1.01
+ $X2=9.505 $Y2=0.515
r192 83 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.67 $Y=1.095
+ $X2=8.505 $Y2=1.095
r193 82 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.34 $Y=1.095
+ $X2=9.505 $Y2=1.095
r194 82 83 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.34 $Y=1.095
+ $X2=8.67 $Y2=1.095
r195 78 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.505 $Y=1.01
+ $X2=8.505 $Y2=1.095
r196 78 80 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=8.505 $Y=1.01
+ $X2=8.505 $Y2=0.515
r197 77 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.67 $Y=1.095
+ $X2=7.505 $Y2=1.095
r198 76 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.34 $Y=1.095
+ $X2=8.505 $Y2=1.095
r199 76 77 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.34 $Y=1.095
+ $X2=7.67 $Y2=1.095
r200 72 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.505 $Y=1.01
+ $X2=7.505 $Y2=1.095
r201 72 74 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=7.505 $Y=1.01
+ $X2=7.505 $Y2=0.515
r202 71 103 8.0097 $w=1.7e-07 $l=3.38e-07 $layer=LI1_cond $X=6.67 $Y=1.095
+ $X2=6.332 $Y2=1.095
r203 70 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.34 $Y=1.095
+ $X2=7.505 $Y2=1.095
r204 70 71 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.34 $Y=1.095
+ $X2=6.67 $Y2=1.095
r205 69 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.325 $Y=0.835
+ $X2=5.16 $Y2=0.835
r206 68 100 8.0097 $w=1.7e-07 $l=3.37e-07 $layer=LI1_cond $X=5.995 $Y=0.835
+ $X2=6.332 $Y2=0.835
r207 68 69 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.995 $Y=0.835
+ $X2=5.325 $Y2=0.835
r208 64 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.16 $Y=0.75
+ $X2=5.16 $Y2=0.835
r209 64 66 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.16 $Y=0.75
+ $X2=5.16 $Y2=0.495
r210 62 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.995 $Y=0.835
+ $X2=5.16 $Y2=0.835
r211 62 63 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.995 $Y=0.835
+ $X2=4.305 $Y2=0.835
r212 59 63 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.14 $Y=0.75
+ $X2=4.305 $Y2=0.835
r213 59 61 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=4.14 $Y=0.75
+ $X2=4.14 $Y2=0.635
r214 58 61 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=4.14 $Y=0.425
+ $X2=4.14 $Y2=0.635
r215 57 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.305 $Y=0.34
+ $X2=3.14 $Y2=0.34
r216 56 58 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.975 $Y=0.34
+ $X2=4.14 $Y2=0.425
r217 56 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.975 $Y=0.34
+ $X2=3.305 $Y2=0.34
r218 52 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=0.425
+ $X2=3.14 $Y2=0.34
r219 52 54 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=3.14 $Y=0.425
+ $X2=3.14 $Y2=0.635
r220 51 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=0.34
+ $X2=2.14 $Y2=0.34
r221 50 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=0.34
+ $X2=3.14 $Y2=0.34
r222 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.975 $Y=0.34
+ $X2=2.305 $Y2=0.34
r223 46 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.425
+ $X2=2.14 $Y2=0.34
r224 46 48 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.14 $Y=0.425
+ $X2=2.14 $Y2=0.635
r225 45 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0.34
+ $X2=1.21 $Y2=0.34
r226 44 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=0.34
+ $X2=2.14 $Y2=0.34
r227 44 45 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.975 $Y=0.34
+ $X2=1.375 $Y2=0.34
r228 40 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.425
+ $X2=1.21 $Y2=0.34
r229 40 42 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.21 $Y=0.425
+ $X2=1.21 $Y2=0.635
r230 38 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=1.21 $Y2=0.34
r231 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.045 $Y=0.34
+ $X2=0.365 $Y2=0.34
r232 34 39 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.425
+ $X2=0.365 $Y2=0.34
r233 34 36 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.24 $Y=0.425
+ $X2=0.24 $Y2=0.515
r234 11 92 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=10.295
+ $Y=0.37 $X2=10.505 $Y2=0.515
r235 10 86 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.365
+ $Y=0.37 $X2=9.505 $Y2=0.515
r236 9 80 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.365
+ $Y=0.37 $X2=8.505 $Y2=0.515
r237 8 74 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.365
+ $Y=0.37 $X2=7.505 $Y2=0.515
r238 7 102 121.333 $w=1.7e-07 $l=7.75999e-07 $layer=licon1_NDIFF $count=1
+ $X=5.95 $Y=0.37 $X2=6.505 $Y2=0.9
r239 7 100 121.333 $w=1.7e-07 $l=5.60245e-07 $layer=licon1_NDIFF $count=1
+ $X=5.95 $Y=0.37 $X2=6.16 $Y2=0.835
r240 6 98 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=5.02
+ $Y=0.37 $X2=5.16 $Y2=0.835
r241 6 66 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=5.02
+ $Y=0.37 $X2=5.16 $Y2=0.495
r242 5 61 182 $w=1.7e-07 $l=3.54789e-07 $layer=licon1_NDIFF $count=1 $X=3.93
+ $Y=0.37 $X2=4.14 $Y2=0.635
r243 4 54 182 $w=1.7e-07 $l=3.54789e-07 $layer=licon1_NDIFF $count=1 $X=2.93
+ $Y=0.37 $X2=3.14 $Y2=0.635
r244 3 48 182 $w=1.7e-07 $l=3.49142e-07 $layer=licon1_NDIFF $count=1 $X=1.945
+ $Y=0.37 $X2=2.14 $Y2=0.635
r245 2 42 182 $w=1.7e-07 $l=3.54789e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.37 $X2=1.21 $Y2=0.635
r246 1 36 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O32AI_4%VGND 1 2 3 4 5 6 21 23 27 31 33 37 39 43 45
+ 49 51 53 58 65 66 69 72 75 78 81 84
r134 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r135 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r136 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r137 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.88
+ $Y2=0
r138 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r139 76 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r140 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r141 69 70 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r142 66 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=0 $X2=9.84
+ $Y2=0
r143 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r144 63 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.17 $Y=0
+ $X2=10.005 $Y2=0
r145 63 65 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=10.17 $Y=0 $X2=10.8
+ $Y2=0
r146 62 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r147 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r148 59 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.825 $Y=0 $X2=5.66
+ $Y2=0
r149 59 61 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.825 $Y=0
+ $X2=6.48 $Y2=0
r150 58 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.84 $Y=0 $X2=7.005
+ $Y2=0
r151 58 61 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.84 $Y=0 $X2=6.48
+ $Y2=0
r152 56 70 1.20413 $w=4.9e-07 $l=4.32e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=4.56
+ $Y2=0
r153 55 56 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r154 53 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.485 $Y=0 $X2=4.65
+ $Y2=0
r155 53 55 276.947 $w=1.68e-07 $l=4.245e-06 $layer=LI1_cond $X=4.485 $Y=0
+ $X2=0.24 $Y2=0
r156 51 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r157 51 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r158 51 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r159 47 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.005 $Y=0.085
+ $X2=10.005 $Y2=0
r160 47 49 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=10.005 $Y=0.085
+ $X2=10.005 $Y2=0.595
r161 46 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.17 $Y=0 $X2=9.005
+ $Y2=0
r162 45 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.84 $Y=0
+ $X2=10.005 $Y2=0
r163 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.84 $Y=0 $X2=9.17
+ $Y2=0
r164 41 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.005 $Y=0.085
+ $X2=9.005 $Y2=0
r165 41 43 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=9.005 $Y=0.085
+ $X2=9.005 $Y2=0.595
r166 40 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.17 $Y=0 $X2=8.005
+ $Y2=0
r167 39 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.84 $Y=0 $X2=9.005
+ $Y2=0
r168 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.84 $Y=0 $X2=8.17
+ $Y2=0
r169 35 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.005 $Y=0.085
+ $X2=8.005 $Y2=0
r170 35 37 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=8.005 $Y=0.085
+ $X2=8.005 $Y2=0.595
r171 34 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.17 $Y=0 $X2=7.005
+ $Y2=0
r172 33 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.84 $Y=0 $X2=8.005
+ $Y2=0
r173 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.84 $Y=0 $X2=7.17
+ $Y2=0
r174 29 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.005 $Y=0.085
+ $X2=7.005 $Y2=0
r175 29 31 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=7.005 $Y=0.085
+ $X2=7.005 $Y2=0.595
r176 25 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.66 $Y=0.085
+ $X2=5.66 $Y2=0
r177 25 27 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=5.66 $Y=0.085
+ $X2=5.66 $Y2=0.495
r178 24 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.815 $Y=0 $X2=4.65
+ $Y2=0
r179 23 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.495 $Y=0 $X2=5.66
+ $Y2=0
r180 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.495 $Y=0
+ $X2=4.815 $Y2=0
r181 19 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.65 $Y=0.085
+ $X2=4.65 $Y2=0
r182 19 21 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=4.65 $Y=0.085
+ $X2=4.65 $Y2=0.415
r183 6 49 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=9.795
+ $Y=0.37 $X2=10.005 $Y2=0.595
r184 5 43 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=8.865
+ $Y=0.37 $X2=9.005 $Y2=0.595
r185 4 37 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=7.795
+ $Y=0.37 $X2=8.005 $Y2=0.595
r186 3 31 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=6.795
+ $Y=0.37 $X2=7.005 $Y2=0.595
r187 2 27 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=5.515
+ $Y=0.37 $X2=5.66 $Y2=0.495
r188 1 21 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.37 $X2=4.65 $Y2=0.415
.ends


* File: sky130_fd_sc_ms__sedfxtp_1.pex.spice
* Created: Fri Aug 28 18:16:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SEDFXTP_1%D 2 5 9 11 12 13 17 18
c41 17 0 4.24886e-20 $X=0.58 $Y=1.275
r42 17 19 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.575 $Y=1.275
+ $X2=0.575 $Y2=1.11
r43 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.58
+ $Y=1.275 $X2=0.58 $Y2=1.275
r44 12 13 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.615 $Y=1.295
+ $X2=0.615 $Y2=1.665
r45 12 18 0.606549 $w=3.78e-07 $l=2e-08 $layer=LI1_cond $X=0.615 $Y=1.295
+ $X2=0.615 $Y2=1.275
r46 9 19 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.64 $Y=0.58 $X2=0.64
+ $Y2=1.11
r47 5 11 334.29 $w=1.8e-07 $l=8.6e-07 $layer=POLY_cond $X=0.495 $Y=2.64
+ $X2=0.495 $Y2=1.78
r48 2 11 41.5618 $w=3.4e-07 $l=1.7e-07 $layer=POLY_cond $X=0.575 $Y=1.61
+ $X2=0.575 $Y2=1.78
r49 1 17 0.848592 $w=3.4e-07 $l=5e-09 $layer=POLY_cond $X=0.575 $Y=1.28
+ $X2=0.575 $Y2=1.275
r50 1 2 56.007 $w=3.4e-07 $l=3.3e-07 $layer=POLY_cond $X=0.575 $Y=1.28 $X2=0.575
+ $Y2=1.61
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_1%A_159_404# 1 2 7 9 13 21 22 23 24 25 26 29
+ 33 35 39 42 47
c116 42 0 9.40653e-20 $X=1.79 $Y=2.035
c117 24 0 4.24886e-20 $X=1.305 $Y=1.065
c118 22 0 1.72336e-19 $X=1.14 $Y=1.605
r119 40 47 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=2.22 $Y=1.685
+ $X2=2.45 $Y2=1.685
r120 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.22
+ $Y=1.685 $X2=2.22 $Y2=1.685
r121 37 39 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.22 $Y=1.95
+ $X2=2.22 $Y2=1.685
r122 36 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=2.035
+ $X2=1.79 $Y2=2.035
r123 35 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.055 $Y=2.035
+ $X2=2.22 $Y2=1.95
r124 35 36 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.055 $Y=2.035
+ $X2=1.875 $Y2=2.035
r125 31 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.79 $Y=2.12
+ $X2=1.79 $Y2=2.035
r126 31 33 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.79 $Y=2.12
+ $X2=1.79 $Y2=2.515
r127 27 29 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=1.765 $Y=0.98
+ $X2=1.765 $Y2=0.765
r128 25 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=2.035
+ $X2=1.79 $Y2=2.035
r129 25 26 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.705 $Y=2.035
+ $X2=1.305 $Y2=2.035
r130 23 27 14.8321 $w=1.01e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.64 $Y=1.065
+ $X2=1.765 $Y2=0.98
r131 23 24 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.64 $Y=1.065
+ $X2=1.305 $Y2=1.065
r132 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.14
+ $Y=1.605 $X2=1.14 $Y2=1.605
r133 19 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.14 $Y=1.95
+ $X2=1.305 $Y2=2.035
r134 19 21 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.14 $Y=1.95
+ $X2=1.14 $Y2=1.605
r135 18 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.14 $Y=1.15
+ $X2=1.305 $Y2=1.065
r136 18 21 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=1.14 $Y=1.15
+ $X2=1.14 $Y2=1.605
r137 17 22 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=1.14 $Y=2.02
+ $X2=1.14 $Y2=1.605
r138 11 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.45 $Y=1.52
+ $X2=2.45 $Y2=1.685
r139 11 13 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.45 $Y=1.52
+ $X2=2.45 $Y2=0.765
r140 7 17 96.0234 $w=1.28e-07 $l=2.55e-07 $layer=POLY_cond $X=0.885 $Y=2.095
+ $X2=1.14 $Y2=2.095
r141 7 9 182.694 $w=1.8e-07 $l=4.7e-07 $layer=POLY_cond $X=0.885 $Y=2.17
+ $X2=0.885 $Y2=2.64
r142 2 33 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=1.645
+ $Y=2.315 $X2=1.79 $Y2=2.515
r143 1 29 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.66
+ $Y=0.555 $X2=1.805 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_1%DE 3 5 6 10 11 13 14 16 17 18 19 21 23 28
+ 31 32 33
c90 33 0 9.40653e-20 $X=1.68 $Y=1.65
c91 32 0 1.3237e-19 $X=1.68 $Y=1.485
r92 31 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=1.485
+ $X2=1.68 $Y2=1.65
r93 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.485 $X2=1.68 $Y2=1.485
r94 28 32 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=1.68 $Y2=1.485
r95 19 21 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.695 $Y=2.24
+ $X2=2.695 $Y2=2.635
r96 17 19 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.605 $Y=2.165
+ $X2=2.695 $Y2=2.24
r97 17 18 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.605 $Y=2.165
+ $X2=2.105 $Y2=2.165
r98 14 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.02 $Y=1.05
+ $X2=2.02 $Y2=1.125
r99 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.02 $Y=1.05 $X2=2.02
+ $Y2=0.765
r100 11 18 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.015 $Y=2.165
+ $X2=2.105 $Y2=2.165
r101 11 25 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=2.015 $Y=2.165
+ $X2=1.74 $Y2=2.165
r102 11 13 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.015 $Y=2.24
+ $X2=2.015 $Y2=2.635
r103 10 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.74 $Y=2.09
+ $X2=1.74 $Y2=2.165
r104 10 33 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.74 $Y=2.09
+ $X2=1.74 $Y2=1.65
r105 7 23 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.68 $Y=1.125
+ $X2=2.02 $Y2=1.125
r106 7 31 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=1.68 $Y=1.2
+ $X2=1.68 $Y2=1.485
r107 5 7 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=1.125
+ $X2=1.68 $Y2=1.125
r108 5 6 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.515 $Y=1.125
+ $X2=1.105 $Y2=1.125
r109 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.03 $Y=1.05
+ $X2=1.105 $Y2=1.125
r110 1 3 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.03 $Y=1.05 $X2=1.03
+ $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_1%A_547_301# 1 2 9 13 15 17 18 19 22 26 29
+ 33 36 40 43 44 45 51 52 58 59 62 69
c234 52 0 8.71884e-20 $X=14.16 $Y=1.665
c235 44 0 7.68314e-20 $X=14.015 $Y=1.665
c236 13 0 1.92249e-19 $X=3.085 $Y=2.635
r237 57 59 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=2.9 $Y=1.67
+ $X2=3.085 $Y2=1.67
r238 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.9
+ $Y=1.67 $X2=2.9 $Y2=1.67
r239 54 57 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.84 $Y=1.67 $X2=2.9
+ $Y2=1.67
r240 52 69 6.51792 $w=2.38e-07 $l=1.15e-07 $layer=LI1_cond $X=14.165 $Y=1.665
+ $X2=14.165 $Y2=1.55
r241 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=1.665
+ $X2=14.16 $Y2=1.665
r242 48 58 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.64 $Y=1.67
+ $X2=2.9 $Y2=1.67
r243 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=1.665
r244 45 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=1.665
+ $X2=2.64 $Y2=1.665
r245 44 51 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.015 $Y=1.665
+ $X2=14.16 $Y2=1.665
r246 44 45 13.8985 $w=1.4e-07 $l=1.123e-05 $layer=MET1_cond $X=14.015 $Y=1.665
+ $X2=2.785 $Y2=1.665
r247 42 69 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=14.2 $Y=0.81
+ $X2=14.2 $Y2=1.55
r248 40 42 10.5918 $w=3.58e-07 $l=2.3e-07 $layer=LI1_cond $X=14.105 $Y=0.58
+ $X2=14.105 $Y2=0.81
r249 36 43 5.46396 $w=2.85e-07 $l=1.73043e-07 $layer=LI1_cond $X=14.165 $Y=2.075
+ $X2=14.12 $Y2=2.227
r250 35 52 0.240092 $w=2.38e-07 $l=5e-09 $layer=LI1_cond $X=14.165 $Y=1.67
+ $X2=14.165 $Y2=1.665
r251 35 36 19.4475 $w=2.38e-07 $l=4.05e-07 $layer=LI1_cond $X=14.165 $Y=1.67
+ $X2=14.165 $Y2=2.075
r252 31 43 5.46396 $w=2.85e-07 $l=1.53e-07 $layer=LI1_cond $X=14.12 $Y=2.38
+ $X2=14.12 $Y2=2.227
r253 31 33 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=14.12 $Y=2.38
+ $X2=14.12 $Y2=2.465
r254 29 63 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.23 $Y=2.215
+ $X2=13.23 $Y2=2.38
r255 29 62 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.23 $Y=2.215
+ $X2=13.23 $Y2=2.05
r256 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.23
+ $Y=2.215 $X2=13.23 $Y2=2.215
r257 26 43 1.09951 $w=3.05e-07 $l=1.65e-07 $layer=LI1_cond $X=13.955 $Y=2.227
+ $X2=14.12 $Y2=2.227
r258 26 28 27.3941 $w=3.03e-07 $l=7.25e-07 $layer=LI1_cond $X=13.955 $Y=2.227
+ $X2=13.23 $Y2=2.227
r259 24 62 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=13.29 $Y=1.015
+ $X2=13.29 $Y2=2.05
r260 22 63 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=13.185 $Y=2.75
+ $X2=13.185 $Y2=2.38
r261 18 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.215 $Y=0.94
+ $X2=13.29 $Y2=1.015
r262 18 19 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=13.215 $Y=0.94
+ $X2=12.825 $Y2=0.94
r263 15 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.75 $Y=0.865
+ $X2=12.825 $Y2=0.94
r264 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=12.75 $Y=0.865
+ $X2=12.75 $Y2=0.58
r265 11 59 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.085 $Y=1.835
+ $X2=3.085 $Y2=1.67
r266 11 13 310.968 $w=1.8e-07 $l=8e-07 $layer=POLY_cond $X=3.085 $Y=1.835
+ $X2=3.085 $Y2=2.635
r267 7 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=1.505
+ $X2=2.84 $Y2=1.67
r268 7 9 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.84 $Y=1.505
+ $X2=2.84 $Y2=0.765
r269 2 33 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=13.985
+ $Y=2.32 $X2=14.12 $Y2=2.465
r270 1 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=13.95
+ $Y=0.37 $X2=14.09 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_1%A_639_85# 1 2 7 9 10 11 14 18 20 23 24 29
+ 30 32 33 37 38 43 45 49
c110 43 0 1.30585e-19 $X=4.41 $Y=0.805
c111 38 0 1.64952e-19 $X=5.655 $Y=1.58
r112 46 49 4.60989 $w=4.78e-07 $l=1.85e-07 $layer=LI1_cond $X=4.1 $Y=2.495
+ $X2=4.285 $Y2=2.495
r113 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.655
+ $Y=1.58 $X2=5.655 $Y2=1.58
r114 35 37 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.655 $Y=1.915
+ $X2=5.655 $Y2=1.58
r115 34 45 2.36881 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.185 $Y=2 $X2=4.045
+ $Y2=2
r116 33 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.49 $Y=2
+ $X2=5.655 $Y2=1.915
r117 33 34 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=5.49 $Y=2
+ $X2=4.185 $Y2=2
r118 32 46 6.90116 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=4.1 $Y=2.255 $X2=4.1
+ $Y2=2.495
r119 31 45 4.06715 $w=2.25e-07 $l=1.09087e-07 $layer=LI1_cond $X=4.1 $Y=2.085
+ $X2=4.045 $Y2=2
r120 31 32 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.1 $Y=2.085
+ $X2=4.1 $Y2=2.255
r121 29 30 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.995
+ $Y=1.78 $X2=3.995 $Y2=1.78
r122 27 45 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=4.045 $Y=1.915
+ $X2=4.045 $Y2=2
r123 27 29 5.55642 $w=2.78e-07 $l=1.35e-07 $layer=LI1_cond $X=4.045 $Y=1.915
+ $X2=4.045 $Y2=1.78
r124 26 29 31.6922 $w=2.78e-07 $l=7.7e-07 $layer=LI1_cond $X=4.045 $Y=1.01
+ $X2=4.045 $Y2=1.78
r125 23 24 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.995
+ $Y=0.42 $X2=3.995 $Y2=0.42
r126 21 43 10.3862 $w=4.03e-07 $l=3.65e-07 $layer=LI1_cond $X=4.045 $Y=0.807
+ $X2=4.41 $Y2=0.807
r127 21 26 2.89865 $w=2.8e-07 $l=2.03e-07 $layer=LI1_cond $X=4.045 $Y=0.807
+ $X2=4.045 $Y2=1.01
r128 21 23 7.61436 $w=2.78e-07 $l=1.85e-07 $layer=LI1_cond $X=4.045 $Y=0.605
+ $X2=4.045 $Y2=0.42
r129 19 38 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.655 $Y=1.92
+ $X2=5.655 $Y2=1.58
r130 19 20 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.655 $Y=1.92
+ $X2=5.655 $Y2=2.085
r131 17 30 101.42 $w=3.3e-07 $l=5.8e-07 $layer=POLY_cond $X=3.995 $Y=1.2
+ $X2=3.995 $Y2=1.78
r132 17 18 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.995 $Y=1.2
+ $X2=3.995 $Y2=1.125
r133 16 24 110.163 $w=3.3e-07 $l=6.3e-07 $layer=POLY_cond $X=3.995 $Y=1.05
+ $X2=3.995 $Y2=0.42
r134 16 18 10.1687 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.995 $Y=1.05
+ $X2=3.995 $Y2=1.125
r135 14 20 198.242 $w=1.8e-07 $l=5.1e-07 $layer=POLY_cond $X=5.58 $Y=2.595
+ $X2=5.58 $Y2=2.085
r136 10 18 16.9349 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.83 $Y=1.125
+ $X2=3.995 $Y2=1.125
r137 10 11 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=3.83 $Y=1.125
+ $X2=3.345 $Y2=1.125
r138 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.27 $Y=1.05
+ $X2=3.345 $Y2=1.125
r139 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.27 $Y=1.05 $X2=3.27
+ $Y2=0.765
r140 2 49 600 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_PDIFF $count=1 $X=4.155
+ $Y=2.275 $X2=4.285 $Y2=2.495
r141 1 43 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=4.27
+ $Y=0.625 $X2=4.41 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_1%SCD 3 7 9 12
c41 12 0 1.14523e-19 $X=5.115 $Y=1.58
c42 3 0 1.30585e-19 $X=5.055 $Y=0.835
r43 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.115 $Y=1.58
+ $X2=5.115 $Y2=1.745
r44 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.115 $Y=1.58
+ $X2=5.115 $Y2=1.415
r45 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.115
+ $Y=1.58 $X2=5.115 $Y2=1.58
r46 9 13 9.25201 $w=3.53e-07 $l=2.85e-07 $layer=LI1_cond $X=5.102 $Y=1.295
+ $X2=5.102 $Y2=1.58
r47 7 15 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=5.19 $Y=2.595
+ $X2=5.19 $Y2=1.745
r48 3 14 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.055 $Y=0.835
+ $X2=5.055 $Y2=1.415
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_1%SCE 1 3 4 5 9 13 14 15 18 20 23
c77 23 0 5.07631e-20 $X=4.565 $Y=1.345
c78 20 0 1.14523e-19 $X=4.56 $Y=1.295
c79 1 0 1.43862e-19 $X=3.535 $Y=3.03
r80 23 26 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.565 $Y=1.345
+ $X2=4.565 $Y2=1.51
r81 23 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.565 $Y=1.345
+ $X2=4.565 $Y2=1.18
r82 20 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.565
+ $Y=1.345 $X2=4.565 $Y2=1.345
r83 16 18 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.415 $Y=0.255
+ $X2=5.415 $Y2=0.835
r84 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.34 $Y=0.18
+ $X2=5.415 $Y2=0.255
r85 14 15 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=5.34 $Y=0.18 $X2=4.7
+ $Y2=0.18
r86 13 25 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=4.625 $Y=0.835
+ $X2=4.625 $Y2=1.18
r87 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.625 $Y=0.255
+ $X2=4.7 $Y2=0.18
r88 10 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.625 $Y=0.255
+ $X2=4.625 $Y2=0.835
r89 9 26 421.75 $w=1.8e-07 $l=1.085e-06 $layer=POLY_cond $X=4.51 $Y=2.595
+ $X2=4.51 $Y2=1.51
r90 7 9 169.089 $w=1.8e-07 $l=4.35e-07 $layer=POLY_cond $X=4.51 $Y=3.03 $X2=4.51
+ $Y2=2.595
r91 4 7 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.42 $Y=3.105
+ $X2=4.51 $Y2=3.03
r92 4 5 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=4.42 $Y=3.105
+ $X2=3.625 $Y2=3.105
r93 1 5 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.535 $Y=3.03
+ $X2=3.625 $Y2=3.105
r94 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.535 $Y=3.03
+ $X2=3.535 $Y2=2.635
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_1%CLK 3 6 8 11 13
c39 11 0 1.38172e-19 $X=6.495 $Y=1.385
r40 11 14 40.6969 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=6.492 $Y=1.385
+ $X2=6.492 $Y2=1.55
r41 11 13 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=6.492 $Y=1.385
+ $X2=6.492 $Y2=1.22
r42 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.495
+ $Y=1.385 $X2=6.495 $Y2=1.385
r43 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.495 $Y=1.295
+ $X2=6.495 $Y2=1.385
r44 6 14 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=6.55 $Y=2.34 $X2=6.55
+ $Y2=1.55
r45 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.4 $Y=0.74 $X2=6.4
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_1%A_1492_74# 1 2 9 11 13 16 20 24 26 27 28
+ 33 34 37 40 41 43 46 47 48 50 51 52 53 55 56 58 60 64 65 68 72
c229 72 0 2.60684e-20 $X=12.84 $Y=1.39
c230 64 0 8.92139e-20 $X=8.575 $Y=2.17
c231 56 0 6.25838e-20 $X=11.76 $Y=1.635
c232 55 0 4.09651e-20 $X=11.76 $Y=1.635
c233 37 0 1.94394e-19 $X=9.17 $Y=0.85
c234 33 0 1.24564e-19 $X=8.49 $Y=1.82
c235 20 0 1.18952e-19 $X=12.765 $Y=2.75
r236 72 85 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.84 $Y=1.39
+ $X2=12.84 $Y2=1.555
r237 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.84
+ $Y=1.39 $X2=12.84 $Y2=1.39
r238 68 71 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=12.84 $Y=1.195
+ $X2=12.84 $Y2=1.39
r239 66 67 14.0135 $w=2.22e-07 $l=2.55e-07 $layer=LI1_cond $X=11.71 $Y=0.94
+ $X2=11.71 $Y2=1.195
r240 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.575
+ $Y=2.17 $X2=8.575 $Y2=2.17
r241 59 67 2.3025 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=11.86 $Y=1.195
+ $X2=11.71 $Y2=1.195
r242 58 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.675 $Y=1.195
+ $X2=12.84 $Y2=1.195
r243 58 59 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=12.675 $Y=1.195
+ $X2=11.86 $Y2=1.195
r244 56 81 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.76 $Y=1.635
+ $X2=11.76 $Y2=1.47
r245 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.76
+ $Y=1.635 $X2=11.76 $Y2=1.635
r246 53 67 4.30642 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.71 $Y=1.28
+ $X2=11.71 $Y2=1.195
r247 53 55 13.6372 $w=2.98e-07 $l=3.55e-07 $layer=LI1_cond $X=11.71 $Y=1.28
+ $X2=11.71 $Y2=1.635
r248 51 66 2.3025 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=11.56 $Y=0.94
+ $X2=11.71 $Y2=0.94
r249 51 52 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=11.56 $Y=0.94
+ $X2=11.02 $Y2=0.94
r250 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.935 $Y=0.855
+ $X2=11.02 $Y2=0.94
r251 49 50 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=10.935 $Y=0.425
+ $X2=10.935 $Y2=0.855
r252 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.85 $Y=0.34
+ $X2=10.935 $Y2=0.425
r253 47 48 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=10.85 $Y=0.34
+ $X2=10.34 $Y2=0.34
r254 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.255 $Y=0.425
+ $X2=10.34 $Y2=0.34
r255 45 46 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=10.255 $Y=0.425
+ $X2=10.255 $Y2=0.85
r256 44 65 2.15711 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=9.34 $Y=0.935
+ $X2=9.212 $Y2=0.935
r257 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.17 $Y=0.935
+ $X2=10.255 $Y2=0.85
r258 43 44 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=10.17 $Y=0.935
+ $X2=9.34 $Y2=0.935
r259 41 76 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=9.175 $Y=1.18
+ $X2=9.045 $Y2=1.18
r260 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.175
+ $Y=1.18 $X2=9.175 $Y2=1.18
r261 38 65 4.27425 $w=2.12e-07 $l=8.5e-08 $layer=LI1_cond $X=9.212 $Y=1.02
+ $X2=9.212 $Y2=0.935
r262 38 40 7.23101 $w=2.53e-07 $l=1.6e-07 $layer=LI1_cond $X=9.212 $Y=1.02
+ $X2=9.212 $Y2=1.18
r263 37 65 4.27425 $w=2.12e-07 $l=1.03899e-07 $layer=LI1_cond $X=9.17 $Y=0.85
+ $X2=9.212 $Y2=0.935
r264 36 37 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=9.17 $Y=0.425
+ $X2=9.17 $Y2=0.85
r265 35 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.575 $Y=0.34
+ $X2=8.49 $Y2=0.34
r266 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.085 $Y=0.34
+ $X2=9.17 $Y2=0.425
r267 34 35 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.085 $Y=0.34
+ $X2=8.575 $Y2=0.34
r268 32 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.49 $Y=0.425
+ $X2=8.49 $Y2=0.34
r269 32 33 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=8.49 $Y=0.425
+ $X2=8.49 $Y2=1.82
r270 28 63 9.54783 $w=2.3e-07 $l=1.8e-07 $layer=LI1_cond $X=8.535 $Y=1.99
+ $X2=8.535 $Y2=2.17
r271 28 33 9.87245 $w=2.3e-07 $l=1.91181e-07 $layer=LI1_cond $X=8.535 $Y=1.99
+ $X2=8.49 $Y2=1.82
r272 28 30 9.49071 $w=3.38e-07 $l=2.8e-07 $layer=LI1_cond $X=8.405 $Y=1.99
+ $X2=8.125 $Y2=1.99
r273 26 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.405 $Y=0.34
+ $X2=8.49 $Y2=0.34
r274 26 27 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=8.405 $Y=0.34
+ $X2=7.765 $Y2=0.34
r275 22 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.64 $Y=0.425
+ $X2=7.765 $Y2=0.34
r276 22 24 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=7.64 $Y=0.425
+ $X2=7.64 $Y2=0.515
r277 20 85 464.508 $w=1.8e-07 $l=1.195e-06 $layer=POLY_cond $X=12.765 $Y=2.75
+ $X2=12.765 $Y2=1.555
r278 16 81 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=11.85 $Y=0.69
+ $X2=11.85 $Y2=1.47
r279 11 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.045 $Y=1.015
+ $X2=9.045 $Y2=1.18
r280 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.045 $Y=1.015
+ $X2=9.045 $Y2=0.695
r281 7 64 56.2646 $w=2.57e-07 $l=3.73497e-07 $layer=POLY_cond $X=8.875 $Y=2.335
+ $X2=8.575 $Y2=2.17
r282 7 9 161.315 $w=1.8e-07 $l=4.15e-07 $layer=POLY_cond $X=8.875 $Y=2.335
+ $X2=8.875 $Y2=2.75
r283 2 30 600 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=1 $X=7.99
+ $Y=1.84 $X2=8.125 $Y2=1.99
r284 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.46
+ $Y=0.37 $X2=7.6 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_1%A_1295_74# 1 2 9 11 13 15 16 20 22 28 32
+ 36 39 40 41 44 47 50 51 53 56 59 60 61 63 66 72 76 77 82
c204 82 0 1.24564e-19 $X=9.34 $Y=1.925
c205 72 0 1.38172e-19 $X=7 $Y=1.96
c206 60 0 1.18952e-19 $X=12.03 $Y=2.475
c207 59 0 2.75377e-20 $X=9.57 $Y=2.39
c208 53 0 3.8828e-20 $X=9.485 $Y=2.09
c209 32 0 4.09651e-20 $X=12.23 $Y=2.46
c210 28 0 7.25971e-20 $X=9.375 $Y=2.75
c211 20 0 1.94394e-19 $X=8.365 $Y=0.695
r212 77 86 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.3 $Y=1.59
+ $X2=12.3 $Y2=1.755
r213 77 85 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.3 $Y=1.59
+ $X2=12.3 $Y2=1.425
r214 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.3
+ $Y=1.59 $X2=12.3 $Y2=1.59
r215 73 76 7.48077 $w=2.83e-07 $l=1.85e-07 $layer=LI1_cond $X=12.115 $Y=1.592
+ $X2=12.3 $Y2=1.592
r216 71 72 2.83598 $w=3.98e-07 $l=8.5e-08 $layer=LI1_cond $X=6.915 $Y=1.96 $X2=7
+ $Y2=1.96
r217 69 71 4.03355 $w=3.98e-07 $l=1.4e-07 $layer=LI1_cond $X=6.775 $Y=1.96
+ $X2=6.915 $Y2=1.96
r218 62 73 3.76007 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=12.115 $Y=1.735
+ $X2=12.115 $Y2=1.592
r219 62 63 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=12.115 $Y=1.735
+ $X2=12.115 $Y2=2.39
r220 60 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.03 $Y=2.475
+ $X2=12.115 $Y2=2.39
r221 60 61 154.947 $w=1.68e-07 $l=2.375e-06 $layer=LI1_cond $X=12.03 $Y=2.475
+ $X2=9.655 $Y2=2.475
r222 59 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.57 $Y=2.39
+ $X2=9.655 $Y2=2.475
r223 58 59 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=9.57 $Y=2.22
+ $X2=9.57 $Y2=2.39
r224 56 83 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.34 $Y=2.09
+ $X2=9.34 $Y2=2.255
r225 56 82 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.34 $Y=2.09
+ $X2=9.34 $Y2=1.925
r226 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.34
+ $Y=2.09 $X2=9.34 $Y2=2.09
r227 53 58 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=9.485 $Y=2.09
+ $X2=9.57 $Y2=2.22
r228 53 55 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=9.485 $Y=2.09
+ $X2=9.34 $Y2=2.09
r229 50 72 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=7.225 $Y=1.995
+ $X2=7 $Y2=1.995
r230 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.225
+ $Y=1.995 $X2=7.225 $Y2=1.995
r231 47 71 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=6.915 $Y=1.76
+ $X2=6.915 $Y2=1.96
r232 46 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.915 $Y=1.01
+ $X2=6.915 $Y2=0.925
r233 46 47 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=6.915 $Y=1.01
+ $X2=6.915 $Y2=1.76
r234 42 66 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.615 $Y=0.925
+ $X2=6.915 $Y2=0.925
r235 42 44 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=6.615 $Y=0.84
+ $X2=6.615 $Y2=0.515
r236 38 51 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=7.225 $Y=1.765
+ $X2=7.225 $Y2=1.995
r237 38 39 13.5877 $w=2.4e-07 $l=9.08295e-08 $layer=POLY_cond $X=7.225 $Y=1.765
+ $X2=7.26 $Y2=1.69
r238 36 85 433.287 $w=1.5e-07 $l=8.45e-07 $layer=POLY_cond $X=12.36 $Y=0.58
+ $X2=12.36 $Y2=1.425
r239 32 86 274.04 $w=1.8e-07 $l=7.05e-07 $layer=POLY_cond $X=12.23 $Y=2.46
+ $X2=12.23 $Y2=1.755
r240 28 83 192.411 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=9.375 $Y=2.75
+ $X2=9.375 $Y2=2.255
r241 24 82 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=9.25 $Y=1.765
+ $X2=9.25 $Y2=1.925
r242 23 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.44 $Y=1.69
+ $X2=8.365 $Y2=1.69
r243 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.175 $Y=1.69
+ $X2=9.25 $Y2=1.765
r244 22 23 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=9.175 $Y=1.69
+ $X2=8.44 $Y2=1.69
r245 18 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.365 $Y=1.615
+ $X2=8.365 $Y2=1.69
r246 18 20 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=8.365 $Y=1.615
+ $X2=8.365 $Y2=0.695
r247 17 40 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.99 $Y=1.69 $X2=7.9
+ $Y2=1.69
r248 16 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.29 $Y=1.69
+ $X2=8.365 $Y2=1.69
r249 16 17 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=8.29 $Y=1.69 $X2=7.99
+ $Y2=1.69
r250 13 40 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=7.9 $Y=1.765 $X2=7.9
+ $Y2=1.69
r251 13 15 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=7.9 $Y=1.765
+ $X2=7.9 $Y2=2.4
r252 12 39 12.1617 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=7.46 $Y=1.69 $X2=7.26
+ $Y2=1.69
r253 11 40 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=7.81 $Y=1.69 $X2=7.9
+ $Y2=1.69
r254 11 12 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=7.81 $Y=1.69
+ $X2=7.46 $Y2=1.69
r255 7 39 13.5877 $w=2.4e-07 $l=1.58114e-07 $layer=POLY_cond $X=7.385 $Y=1.615
+ $X2=7.26 $Y2=1.69
r256 7 9 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=7.385 $Y=1.615
+ $X2=7.385 $Y2=0.74
r257 2 69 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=6.64
+ $Y=1.78 $X2=6.775 $Y2=1.96
r258 1 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.475
+ $Y=0.37 $X2=6.615 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_1%A_1910_71# 1 2 9 13 19 21 23 24 28 31 32
+ 34 35 41 45 52 55
c113 34 0 6.25838e-20 $X=11.22 $Y=1.36
r114 47 48 5.82061 $w=2.62e-07 $l=1.25e-07 $layer=LI1_cond $X=10.595 $Y=1.36
+ $X2=10.72 $Y2=1.36
r115 43 45 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=10.55 $Y=2.095
+ $X2=10.72 $Y2=2.095
r116 39 52 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.73 $Y=1.32
+ $X2=9.805 $Y2=1.32
r117 39 49 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=9.73 $Y=1.32
+ $X2=9.625 $Y2=1.32
r118 38 41 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=9.73 $Y=1.32
+ $X2=9.895 $Y2=1.32
r119 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.73
+ $Y=1.32 $X2=9.73 $Y2=1.32
r120 35 55 12.8191 $w=2.82e-07 $l=7.5e-08 $layer=POLY_cond $X=11.22 $Y=1.317
+ $X2=11.295 $Y2=1.317
r121 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.22
+ $Y=1.36 $X2=11.22 $Y2=1.36
r122 32 48 3.69502 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.805 $Y=1.36
+ $X2=10.72 $Y2=1.36
r123 32 34 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=10.805 $Y=1.36
+ $X2=11.22 $Y2=1.36
r124 31 45 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.72 $Y=1.97
+ $X2=10.72 $Y2=2.095
r125 30 48 3.26844 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.72 $Y=1.525
+ $X2=10.72 $Y2=1.36
r126 30 31 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=10.72 $Y=1.525
+ $X2=10.72 $Y2=1.97
r127 26 47 3.26844 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.595 $Y=1.195
+ $X2=10.595 $Y2=1.36
r128 26 28 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.595 $Y=1.195
+ $X2=10.595 $Y2=0.81
r129 24 47 5.45986 $w=2.62e-07 $l=1.18427e-07 $layer=LI1_cond $X=10.51 $Y=1.28
+ $X2=10.595 $Y2=1.36
r130 24 41 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=10.51 $Y=1.28
+ $X2=9.895 $Y2=1.28
r131 21 55 33.3298 $w=2.82e-07 $l=2.88468e-07 $layer=POLY_cond $X=11.49 $Y=1.11
+ $X2=11.295 $Y2=1.317
r132 21 23 134.96 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=11.49 $Y=1.11
+ $X2=11.49 $Y2=0.69
r133 17 55 13.2911 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=11.295 $Y=1.525
+ $X2=11.295 $Y2=1.317
r134 17 19 363.444 $w=1.8e-07 $l=9.35e-07 $layer=POLY_cond $X=11.295 $Y=1.525
+ $X2=11.295 $Y2=2.46
r135 11 52 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.805 $Y=1.485
+ $X2=9.805 $Y2=1.32
r136 11 13 491.718 $w=1.8e-07 $l=1.265e-06 $layer=POLY_cond $X=9.805 $Y=1.485
+ $X2=9.805 $Y2=2.75
r137 7 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.625 $Y=1.155
+ $X2=9.625 $Y2=1.32
r138 7 9 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=9.625 $Y=1.155
+ $X2=9.625 $Y2=0.695
r139 2 43 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.415
+ $Y=1.99 $X2=10.55 $Y2=2.135
r140 1 28 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=10.455
+ $Y=0.37 $X2=10.595 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_1%A_1688_97# 1 2 9 13 17 23 27 28 29 31 32
+ 33
r104 32 37 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.3 $Y=1.665
+ $X2=10.3 $Y2=1.83
r105 32 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.3 $Y=1.665
+ $X2=10.3 $Y2=1.5
r106 31 33 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=10.3 $Y=1.665
+ $X2=10.135 $Y2=1.665
r107 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.3
+ $Y=1.665 $X2=10.3 $Y2=1.665
r108 28 29 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=9.075 $Y=2.39
+ $X2=9.075 $Y2=2.56
r109 26 27 1.34256 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.005 $Y=1.705
+ $X2=8.875 $Y2=1.705
r110 26 33 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=9.005 $Y=1.705
+ $X2=10.135 $Y2=1.705
r111 23 29 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=9.15 $Y=2.75
+ $X2=9.15 $Y2=2.56
r112 19 27 5.16603 $w=1.7e-07 $l=1.05119e-07 $layer=LI1_cond $X=8.92 $Y=1.79
+ $X2=8.875 $Y2=1.705
r113 19 28 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=8.92 $Y=1.79 $X2=8.92
+ $Y2=2.39
r114 15 27 5.16603 $w=1.7e-07 $l=1.05119e-07 $layer=LI1_cond $X=8.83 $Y=1.62
+ $X2=8.875 $Y2=1.705
r115 15 17 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=8.83 $Y=1.62
+ $X2=8.83 $Y2=0.76
r116 13 36 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=10.38 $Y=0.69
+ $X2=10.38 $Y2=1.5
r117 9 37 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=10.325 $Y=2.41
+ $X2=10.325 $Y2=1.83
r118 2 23 600 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_PDIFF $count=1 $X=8.965
+ $Y=2.54 $X2=9.15 $Y2=2.75
r119 1 17 182 $w=1.7e-07 $l=5.09264e-07 $layer=licon1_NDIFF $count=1 $X=8.44
+ $Y=0.485 $X2=8.83 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_1%A_2385_74# 1 2 9 13 15 16 19 21 23 24 25
+ 27 29 31 33 35 38 39 42 48 50
c137 25 0 1.37761e-19 $X=12.065 $Y=0.77
r138 55 56 2.23148 $w=4.32e-07 $l=2e-08 $layer=POLY_cond $X=13.875 $Y=1.335
+ $X2=13.895 $Y2=1.335
r139 51 55 10.5995 $w=4.32e-07 $l=9.5e-08 $layer=POLY_cond $X=13.78 $Y=1.335
+ $X2=13.875 $Y2=1.335
r140 50 53 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=13.78 $Y=1.215
+ $X2=13.78 $Y2=1.38
r141 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.78
+ $Y=1.215 $X2=13.78 $Y2=1.215
r142 42 53 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=13.7 $Y=1.735
+ $X2=13.7 $Y2=1.38
r143 40 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.345 $Y=1.82
+ $X2=13.26 $Y2=1.82
r144 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.615 $Y=1.82
+ $X2=13.7 $Y2=1.735
r145 39 40 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=13.615 $Y=1.82
+ $X2=13.345 $Y2=1.82
r146 38 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.26 $Y=1.735
+ $X2=13.26 $Y2=1.82
r147 37 38 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=13.26 $Y=0.94
+ $X2=13.26 $Y2=1.735
r148 36 47 11.3627 $w=3.06e-07 $l=3.78622e-07 $layer=LI1_cond $X=12.805 $Y=1.82
+ $X2=12.587 $Y2=2.105
r149 35 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.175 $Y=1.82
+ $X2=13.26 $Y2=1.82
r150 35 36 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=13.175 $Y=1.82
+ $X2=12.805 $Y2=1.82
r151 31 47 2.54614 $w=4.35e-07 $l=5.2e-08 $layer=LI1_cond $X=12.587 $Y=2.157
+ $X2=12.587 $Y2=2.105
r152 31 33 17.4324 $w=4.33e-07 $l=6.58e-07 $layer=LI1_cond $X=12.587 $Y=2.157
+ $X2=12.587 $Y2=2.815
r153 30 44 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.23 $Y=0.855
+ $X2=12.065 $Y2=0.855
r154 29 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.175 $Y=0.855
+ $X2=13.26 $Y2=0.94
r155 29 30 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=13.175 $Y=0.855
+ $X2=12.23 $Y2=0.855
r156 25 44 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.065 $Y=0.77
+ $X2=12.065 $Y2=0.855
r157 25 27 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=12.065 $Y=0.77
+ $X2=12.065 $Y2=0.515
r158 21 24 38.8775 $w=1.65e-07 $l=1.95e-07 $layer=POLY_cond $X=14.865 $Y=1.23
+ $X2=14.865 $Y2=1.425
r159 21 23 157.453 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=14.865 $Y=1.23
+ $X2=14.865 $Y2=0.74
r160 17 24 38.8775 $w=1.65e-07 $l=1.95e-07 $layer=POLY_cond $X=14.865 $Y=1.62
+ $X2=14.865 $Y2=1.425
r161 17 19 303.194 $w=1.8e-07 $l=7.8e-07 $layer=POLY_cond $X=14.865 $Y=1.62
+ $X2=14.865 $Y2=2.4
r162 16 56 10.5996 $w=4.32e-07 $l=1.27279e-07 $layer=POLY_cond $X=13.985
+ $Y=1.425 $X2=13.895 $Y2=1.335
r163 15 24 5.85142 $w=3.9e-07 $l=9e-08 $layer=POLY_cond $X=14.775 $Y=1.425
+ $X2=14.865 $Y2=1.425
r164 15 16 112.657 $w=3.9e-07 $l=7.9e-07 $layer=POLY_cond $X=14.775 $Y=1.425
+ $X2=13.985 $Y2=1.425
r165 11 56 23.3057 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=13.895 $Y=1.62
+ $X2=13.895 $Y2=1.335
r166 11 13 396.484 $w=1.8e-07 $l=1.02e-06 $layer=POLY_cond $X=13.895 $Y=1.62
+ $X2=13.895 $Y2=2.64
r167 7 55 27.7542 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=13.875 $Y=1.05
+ $X2=13.875 $Y2=1.335
r168 7 9 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=13.875 $Y=1.05 $X2=13.875
+ $Y2=0.58
r169 2 47 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=12.32
+ $Y=1.96 $X2=12.455 $Y2=2.105
r170 2 33 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=12.32
+ $Y=1.96 $X2=12.455 $Y2=2.815
r171 1 44 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=11.925
+ $Y=0.37 $X2=12.065 $Y2=0.855
r172 1 27 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=11.925
+ $Y=0.37 $X2=12.065 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_1%A_27_74# 1 2 3 4 14 17 19 22 23 24 26 27
+ 28 31 35 38 42 44 47 49
c118 35 0 1.43862e-19 $X=3.31 $Y=2.46
r119 39 42 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=0.17 $Y=0.645
+ $X2=0.35 $Y2=0.645
r120 38 49 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=3.31 $Y=2.29
+ $X2=3.27 $Y2=2.375
r121 37 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.31 $Y=1.335
+ $X2=3.31 $Y2=1.25
r122 37 38 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=3.31 $Y=1.335
+ $X2=3.31 $Y2=2.29
r123 35 49 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.27 $Y=2.46 $X2=3.27
+ $Y2=2.375
r124 29 47 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.055 $Y=1.25
+ $X2=3.31 $Y2=1.25
r125 29 31 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=3.055 $Y=1.165
+ $X2=3.055 $Y2=0.765
r126 27 49 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.145 $Y=2.375
+ $X2=3.27 $Y2=2.375
r127 27 28 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.145 $Y=2.375
+ $X2=2.215 $Y2=2.375
r128 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.13 $Y=2.46
+ $X2=2.215 $Y2=2.375
r129 25 26 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.13 $Y=2.46
+ $X2=2.13 $Y2=2.905
r130 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.045 $Y=2.99
+ $X2=2.13 $Y2=2.905
r131 23 24 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.045 $Y=2.99
+ $X2=1.535 $Y2=2.99
r132 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.45 $Y=2.905
+ $X2=1.535 $Y2=2.99
r133 21 22 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.45 $Y=2.46
+ $X2=1.45 $Y2=2.905
r134 20 44 2.90867 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.435 $Y=2.375
+ $X2=0.26 $Y2=2.375
r135 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.365 $Y=2.375
+ $X2=1.45 $Y2=2.46
r136 19 20 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=1.365 $Y=2.375
+ $X2=0.435 $Y2=2.375
r137 15 44 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.46
+ $X2=0.26 $Y2=2.375
r138 15 17 0.164635 $w=3.48e-07 $l=5e-09 $layer=LI1_cond $X=0.26 $Y=2.46
+ $X2=0.26 $Y2=2.465
r139 14 44 3.58051 $w=2.6e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.17 $Y=2.29
+ $X2=0.26 $Y2=2.375
r140 13 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=0.81
+ $X2=0.17 $Y2=0.645
r141 13 14 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=0.17 $Y=0.81
+ $X2=0.17 $Y2=2.29
r142 4 35 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.175
+ $Y=2.315 $X2=3.31 $Y2=2.46
r143 3 17 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.27 $Y2=2.465
r144 2 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.915
+ $Y=0.555 $X2=3.055 $Y2=0.765
r145 1 42 182 $w=1.7e-07 $l=3.67083e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.35 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_1%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50
+ 54 58 60 62 67 68 70 71 73 74 76 77 79 80 81 93 100 118 125 131 134 137 141
c162 3 0 9.48608e-20 $X=4.6 $Y=2.275
r163 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r164 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r165 134 135 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r166 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r167 129 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=15.12 $Y2=3.33
r168 129 138 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=13.68 $Y2=3.33
r169 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r170 126 137 10.6558 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=13.785 $Y=3.33
+ $X2=13.557 $Y2=3.33
r171 126 128 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=13.785 $Y=3.33
+ $X2=14.64 $Y2=3.33
r172 125 140 4.02656 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=15.005 $Y=3.33
+ $X2=15.182 $Y2=3.33
r173 125 128 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=15.005 $Y=3.33
+ $X2=14.64 $Y2=3.33
r174 124 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r175 123 124 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r176 121 124 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=13.2 $Y2=3.33
r177 120 123 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=11.28 $Y=3.33
+ $X2=13.2 $Y2=3.33
r178 120 121 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r179 118 137 10.6558 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=13.33 $Y=3.33
+ $X2=13.557 $Y2=3.33
r180 118 123 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=13.33 $Y=3.33
+ $X2=13.2 $Y2=3.33
r181 117 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r182 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r183 114 117 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.8 $Y2=3.33
r184 113 114 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r185 111 114 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=9.84 $Y2=3.33
r186 110 113 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=7.92 $Y=3.33
+ $X2=9.84 $Y2=3.33
r187 110 111 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r188 108 135 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r189 107 108 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r190 105 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.49 $Y=3.33
+ $X2=6.325 $Y2=3.33
r191 105 107 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=6.49 $Y=3.33
+ $X2=7.44 $Y2=3.33
r192 104 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r193 104 132 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r194 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r195 101 131 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.13 $Y=3.33
+ $X2=5.005 $Y2=3.33
r196 101 103 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=5.13 $Y=3.33
+ $X2=6 $Y2=3.33
r197 100 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.16 $Y=3.33
+ $X2=6.325 $Y2=3.33
r198 100 103 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=6.16 $Y=3.33
+ $X2=6 $Y2=3.33
r199 99 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r200 98 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r201 96 99 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.56 $Y2=3.33
r202 95 98 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.56 $Y2=3.33
r203 95 96 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r204 93 131 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.88 $Y=3.33
+ $X2=5.005 $Y2=3.33
r205 93 98 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.88 $Y=3.33
+ $X2=4.56 $Y2=3.33
r206 92 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r207 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r208 89 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r209 88 91 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r210 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r211 85 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r212 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r213 81 111 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.68 $Y=3.33
+ $X2=7.92 $Y2=3.33
r214 81 108 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.68 $Y=3.33
+ $X2=7.44 $Y2=3.33
r215 79 116 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=10.905 $Y=3.33
+ $X2=10.8 $Y2=3.33
r216 79 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.905 $Y=3.33
+ $X2=11.07 $Y2=3.33
r217 78 120 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=11.235 $Y=3.33
+ $X2=11.28 $Y2=3.33
r218 78 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.235 $Y=3.33
+ $X2=11.07 $Y2=3.33
r219 76 113 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=9.865 $Y=3.33
+ $X2=9.84 $Y2=3.33
r220 76 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.865 $Y=3.33
+ $X2=10.03 $Y2=3.33
r221 75 116 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=10.195 $Y=3.33
+ $X2=10.8 $Y2=3.33
r222 75 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.195 $Y=3.33
+ $X2=10.03 $Y2=3.33
r223 73 107 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=7.51 $Y=3.33
+ $X2=7.44 $Y2=3.33
r224 73 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.51 $Y=3.33
+ $X2=7.675 $Y2=3.33
r225 72 110 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=7.84 $Y=3.33
+ $X2=7.92 $Y2=3.33
r226 72 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.84 $Y=3.33
+ $X2=7.675 $Y2=3.33
r227 70 91 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.385 $Y=3.33
+ $X2=2.16 $Y2=3.33
r228 70 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.385 $Y=3.33
+ $X2=2.51 $Y2=3.33
r229 69 95 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.635 $Y=3.33
+ $X2=2.64 $Y2=3.33
r230 69 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.635 $Y=3.33
+ $X2=2.51 $Y2=3.33
r231 67 84 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.72 $Y2=3.33
r232 67 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.07 $Y2=3.33
r233 66 88 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.195 $Y=3.33
+ $X2=1.2 $Y2=3.33
r234 66 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.195 $Y=3.33
+ $X2=1.07 $Y2=3.33
r235 62 65 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=15.13 $Y=1.985
+ $X2=15.13 $Y2=2.815
r236 60 140 3.1166 $w=2.5e-07 $l=1.07912e-07 $layer=LI1_cond $X=15.13 $Y=3.245
+ $X2=15.182 $Y2=3.33
r237 60 65 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=15.13 $Y=3.245
+ $X2=15.13 $Y2=2.815
r238 56 137 1.82608 $w=4.55e-07 $l=8.5e-08 $layer=LI1_cond $X=13.557 $Y=3.245
+ $X2=13.557 $Y2=3.33
r239 56 58 11.3036 $w=4.53e-07 $l=4.3e-07 $layer=LI1_cond $X=13.557 $Y=3.245
+ $X2=13.557 $Y2=2.815
r240 52 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.07 $Y=3.245
+ $X2=11.07 $Y2=3.33
r241 52 54 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.07 $Y=3.245
+ $X2=11.07 $Y2=2.815
r242 48 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.03 $Y=3.245
+ $X2=10.03 $Y2=3.33
r243 48 50 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.03 $Y=3.245
+ $X2=10.03 $Y2=2.815
r244 44 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.675 $Y=3.245
+ $X2=7.675 $Y2=3.33
r245 44 46 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=7.675 $Y=3.245
+ $X2=7.675 $Y2=2.785
r246 40 134 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.325 $Y=3.245
+ $X2=6.325 $Y2=3.33
r247 40 42 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=6.325 $Y=3.245
+ $X2=6.325 $Y2=2.755
r248 36 131 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=3.245
+ $X2=5.005 $Y2=3.33
r249 36 38 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=5.005 $Y=3.245
+ $X2=5.005 $Y2=2.765
r250 32 71 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=3.245
+ $X2=2.51 $Y2=3.33
r251 32 34 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=2.51 $Y=3.245
+ $X2=2.51 $Y2=2.8
r252 28 68 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=3.245
+ $X2=1.07 $Y2=3.33
r253 28 30 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=1.07 $Y=3.245
+ $X2=1.07 $Y2=2.805
r254 9 65 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=14.955
+ $Y=1.84 $X2=15.09 $Y2=2.815
r255 9 62 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=14.955
+ $Y=1.84 $X2=15.09 $Y2=1.985
r256 8 58 600 $w=1.7e-07 $l=3.94208e-07 $layer=licon1_PDIFF $count=1 $X=13.275
+ $Y=2.54 $X2=13.555 $Y2=2.815
r257 7 54 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=10.945
+ $Y=1.96 $X2=11.07 $Y2=2.815
r258 6 50 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=9.895
+ $Y=2.54 $X2=10.03 $Y2=2.815
r259 5 46 600 $w=1.7e-07 $l=1.00556e-06 $layer=licon1_PDIFF $count=1 $X=7.55
+ $Y=1.84 $X2=7.675 $Y2=2.785
r260 4 42 600 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=6.2
+ $Y=1.78 $X2=6.325 $Y2=2.755
r261 3 38 600 $w=1.7e-07 $l=6.47263e-07 $layer=licon1_PDIFF $count=1 $X=4.6
+ $Y=2.275 $X2=4.965 $Y2=2.765
r262 2 34 600 $w=1.7e-07 $l=6.42067e-07 $layer=licon1_PDIFF $count=1 $X=2.105
+ $Y=2.315 $X2=2.47 $Y2=2.8
r263 1 30 600 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=1 $X=0.975
+ $Y=2.32 $X2=1.11 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_1%A_669_111# 1 2 3 4 5 6 21 24 25 26 28 30
+ 33 37 38 40 41 44 45 46 47 51 54 55 57 60 63 65 66 68 69
c189 63 0 1.92249e-19 $X=3.705 $Y=2.295
c190 57 0 7.25971e-20 $X=8.65 $Y=2.815
c191 47 0 2.28482e-20 $X=8.01 $Y=2.415
c192 37 0 1.64952e-19 $X=5.99 $Y=1.16
c193 25 0 9.48608e-20 $X=4.54 $Y=2.99
r194 65 66 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=5.805 $Y=2.377
+ $X2=5.64 $Y2=2.377
r195 62 63 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=3.65 $Y=0.995
+ $X2=3.65 $Y2=2.295
r196 60 62 10.6507 $w=3.43e-07 $l=2.3e-07 $layer=LI1_cond $X=3.562 $Y=0.765
+ $X2=3.562 $Y2=0.995
r197 55 57 21.6659 $w=2.48e-07 $l=4.7e-07 $layer=LI1_cond $X=8.18 $Y=2.855
+ $X2=8.65 $Y2=2.855
r198 54 55 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.095 $Y=2.73
+ $X2=8.18 $Y2=2.855
r199 53 54 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=8.095 $Y=2.5
+ $X2=8.095 $Y2=2.73
r200 49 51 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=8.11 $Y=1.48
+ $X2=8.11 $Y2=0.76
r201 48 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.79 $Y=2.415
+ $X2=7.705 $Y2=2.415
r202 47 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.01 $Y=2.415
+ $X2=8.095 $Y2=2.5
r203 47 48 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.01 $Y=2.415
+ $X2=7.79 $Y2=2.415
r204 45 49 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.985 $Y=1.565
+ $X2=8.11 $Y2=1.48
r205 45 46 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=7.985 $Y=1.565
+ $X2=7.79 $Y2=1.565
r206 44 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.705 $Y=2.33
+ $X2=7.705 $Y2=2.415
r207 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.705 $Y=1.65
+ $X2=7.79 $Y2=1.565
r208 43 44 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.705 $Y=1.65
+ $X2=7.705 $Y2=2.33
r209 41 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.62 $Y=2.415
+ $X2=7.705 $Y2=2.415
r210 41 68 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=7.62 $Y=2.415
+ $X2=6.16 $Y2=2.415
r211 40 68 5.08946 $w=2.43e-07 $l=8.5e-08 $layer=LI1_cond $X=6.075 $Y=2.377
+ $X2=6.16 $Y2=2.377
r212 40 65 12.7004 $w=2.43e-07 $l=2.7e-07 $layer=LI1_cond $X=6.075 $Y=2.377
+ $X2=5.805 $Y2=2.377
r213 39 40 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=6.075 $Y=1.245
+ $X2=6.075 $Y2=2.255
r214 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.99 $Y=1.16
+ $X2=6.075 $Y2=1.245
r215 37 38 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.99 $Y=1.16
+ $X2=5.795 $Y2=1.16
r216 31 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.63 $Y=1.075
+ $X2=5.795 $Y2=1.16
r217 31 33 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=5.63 $Y=1.075
+ $X2=5.63 $Y2=0.835
r218 30 66 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=4.71 $Y=2.34
+ $X2=5.64 $Y2=2.34
r219 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.625 $Y=2.425
+ $X2=4.71 $Y2=2.34
r220 27 28 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.625 $Y=2.425
+ $X2=4.625 $Y2=2.905
r221 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.54 $Y=2.99
+ $X2=4.625 $Y2=2.905
r222 25 26 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.54 $Y=2.99
+ $X2=3.845 $Y2=2.99
r223 22 26 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.705 $Y=2.905
+ $X2=3.845 $Y2=2.99
r224 22 24 18.3156 $w=2.78e-07 $l=4.45e-07 $layer=LI1_cond $X=3.705 $Y=2.905
+ $X2=3.705 $Y2=2.46
r225 21 63 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=3.705 $Y=2.435
+ $X2=3.705 $Y2=2.295
r226 21 24 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=3.705 $Y=2.435
+ $X2=3.705 $Y2=2.46
r227 6 57 600 $w=1.7e-07 $l=3.33729e-07 $layer=licon1_PDIFF $count=1 $X=8.52
+ $Y=2.54 $X2=8.65 $Y2=2.815
r228 5 65 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=5.67
+ $Y=2.275 $X2=5.805 $Y2=2.42
r229 4 24 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.625
+ $Y=2.315 $X2=3.76 $Y2=2.46
r230 3 51 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=8.01
+ $Y=0.485 $X2=8.15 $Y2=0.76
r231 2 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.49
+ $Y=0.625 $X2=5.63 $Y2=0.835
r232 1 60 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=3.345
+ $Y=0.555 $X2=3.555 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_1%Q 1 2 7 8 9 10 11 12 13
r18 12 13 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=14.645 $Y=2.405
+ $X2=14.645 $Y2=2.775
r19 11 12 14.2361 $w=3.38e-07 $l=4.2e-07 $layer=LI1_cond $X=14.645 $Y=1.985
+ $X2=14.645 $Y2=2.405
r20 10 11 10.8465 $w=3.38e-07 $l=3.2e-07 $layer=LI1_cond $X=14.645 $Y=1.665
+ $X2=14.645 $Y2=1.985
r21 9 10 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=14.645 $Y=1.295
+ $X2=14.645 $Y2=1.665
r22 8 9 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=14.645 $Y=0.925
+ $X2=14.645 $Y2=1.295
r23 7 8 13.8971 $w=3.38e-07 $l=4.1e-07 $layer=LI1_cond $X=14.645 $Y=0.515
+ $X2=14.645 $Y2=0.925
r24 2 13 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=14.515
+ $Y=1.84 $X2=14.64 $Y2=2.815
r25 2 11 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=14.515
+ $Y=1.84 $X2=14.64 $Y2=1.985
r26 1 7 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=14.505
+ $Y=0.37 $X2=14.65 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SEDFXTP_1%VGND 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50
+ 54 56 58 61 62 64 65 67 68 69 71 76 97 104 117 123 126 129 132 137 143 146
c173 30 0 1.72336e-19 $X=1.245 $Y=0.58
r174 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r175 141 143 9.13714 $w=6.83e-07 $l=7.5e-08 $layer=LI1_cond $X=13.68 $Y=0.257
+ $X2=13.755 $Y2=0.257
r176 141 142 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r177 139 141 1.57149 $w=6.83e-07 $l=9e-08 $layer=LI1_cond $X=13.59 $Y=0.257
+ $X2=13.68 $Y2=0.257
r178 136 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=13.68 $Y2=0
r179 135 139 6.80979 $w=6.83e-07 $l=3.9e-07 $layer=LI1_cond $X=13.2 $Y=0.257
+ $X2=13.59 $Y2=0.257
r180 135 137 14.812 $w=6.83e-07 $l=4e-07 $layer=LI1_cond $X=13.2 $Y=0.257
+ $X2=12.8 $Y2=0.257
r181 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r182 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r183 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r184 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r185 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r186 121 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=15.12 $Y2=0
r187 121 142 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=13.68 $Y2=0
r188 120 143 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=14.64 $Y=0
+ $X2=13.755 $Y2=0
r189 120 121 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r190 117 145 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=14.995 $Y=0
+ $X2=15.177 $Y2=0
r191 117 120 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=14.995 $Y=0
+ $X2=14.64 $Y2=0
r192 116 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r193 115 137 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=12.72 $Y=0 $X2=12.8
+ $Y2=0
r194 115 116 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r195 113 116 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.72 $Y2=0
r196 113 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r197 112 115 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=11.76 $Y=0
+ $X2=12.72 $Y2=0
r198 112 113 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r199 110 132 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.44 $Y=0
+ $X2=11.315 $Y2=0
r200 110 112 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=11.44 $Y=0
+ $X2=11.76 $Y2=0
r201 108 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r202 108 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=9.84 $Y2=0
r203 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r204 105 129 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10 $Y=0 $X2=9.875
+ $Y2=0
r205 105 107 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=10 $Y=0 $X2=10.8
+ $Y2=0
r206 104 132 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.19 $Y=0
+ $X2=11.315 $Y2=0
r207 104 107 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=11.19 $Y=0
+ $X2=10.8 $Y2=0
r208 103 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r209 102 103 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r210 99 102 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=7.44 $Y=0
+ $X2=9.36 $Y2=0
r211 99 100 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r212 97 129 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.75 $Y=0
+ $X2=9.875 $Y2=0
r213 97 102 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=9.75 $Y=0 $X2=9.36
+ $Y2=0
r214 96 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r215 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r216 93 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r217 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r218 90 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r219 89 92 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r220 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r221 87 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r222 86 87 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r223 84 87 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.56 $Y2=0
r224 84 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=2.16 $Y2=0
r225 83 86 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r226 83 84 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r227 81 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.235
+ $Y2=0
r228 81 83 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r229 80 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r230 80 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r231 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r232 77 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.41 $Y=0
+ $X2=1.245 $Y2=0
r233 77 79 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.68
+ $Y2=0
r234 76 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.07 $Y=0
+ $X2=2.235 $Y2=0
r235 76 79 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.68
+ $Y2=0
r236 74 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r237 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r238 71 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.08 $Y=0
+ $X2=1.245 $Y2=0
r239 71 73 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.08 $Y=0 $X2=0.72
+ $Y2=0
r240 69 103 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=7.68 $Y=0
+ $X2=9.36 $Y2=0
r241 69 100 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.68 $Y=0
+ $X2=7.44 $Y2=0
r242 67 95 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=7.005 $Y=0 $X2=6.96
+ $Y2=0
r243 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.005 $Y=0 $X2=7.17
+ $Y2=0
r244 66 99 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.335 $Y=0
+ $X2=7.44 $Y2=0
r245 66 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.335 $Y=0 $X2=7.17
+ $Y2=0
r246 64 92 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=6.02 $Y=0 $X2=6 $Y2=0
r247 64 65 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.02 $Y=0 $X2=6.15
+ $Y2=0
r248 63 95 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.28 $Y=0 $X2=6.96
+ $Y2=0
r249 63 65 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.28 $Y=0 $X2=6.15
+ $Y2=0
r250 61 86 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=4.755 $Y=0
+ $X2=4.56 $Y2=0
r251 61 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.755 $Y=0 $X2=4.88
+ $Y2=0
r252 60 89 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=5.005 $Y=0 $X2=5.04
+ $Y2=0
r253 60 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.005 $Y=0 $X2=4.88
+ $Y2=0
r254 56 145 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=15.12 $Y=0.085
+ $X2=15.177 $Y2=0
r255 56 58 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=15.12 $Y=0.085
+ $X2=15.12 $Y2=0.515
r256 52 132 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.315 $Y=0.085
+ $X2=11.315 $Y2=0
r257 52 54 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.315 $Y=0.085
+ $X2=11.315 $Y2=0.515
r258 48 129 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.875 $Y=0.085
+ $X2=9.875 $Y2=0
r259 48 50 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.875 $Y=0.085
+ $X2=9.875 $Y2=0.515
r260 44 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.17 $Y=0.085
+ $X2=7.17 $Y2=0
r261 44 46 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=7.17 $Y=0.085
+ $X2=7.17 $Y2=0.55
r262 40 65 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.15 $Y=0.085
+ $X2=6.15 $Y2=0
r263 40 42 25.7083 $w=2.58e-07 $l=5.8e-07 $layer=LI1_cond $X=6.15 $Y=0.085
+ $X2=6.15 $Y2=0.665
r264 36 62 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.88 $Y=0.085
+ $X2=4.88 $Y2=0
r265 36 38 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=4.88 $Y=0.085
+ $X2=4.88 $Y2=0.805
r266 32 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.235 $Y=0.085
+ $X2=2.235 $Y2=0
r267 32 34 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.235 $Y=0.085
+ $X2=2.235 $Y2=0.765
r268 28 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=0.085
+ $X2=1.245 $Y2=0
r269 28 30 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.245 $Y=0.085
+ $X2=1.245 $Y2=0.58
r270 9 58 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.94
+ $Y=0.37 $X2=15.08 $Y2=0.515
r271 8 139 91 $w=1.7e-07 $l=8.34356e-07 $layer=licon1_NDIFF $count=2 $X=12.825
+ $Y=0.37 $X2=13.59 $Y2=0.515
r272 7 54 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=11.13
+ $Y=0.37 $X2=11.275 $Y2=0.515
r273 6 50 182 $w=1.7e-07 $l=2.2951e-07 $layer=licon1_NDIFF $count=1 $X=9.7
+ $Y=0.485 $X2=9.915 $Y2=0.515
r274 5 46 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=7.025
+ $Y=0.37 $X2=7.17 $Y2=0.55
r275 4 42 182 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_NDIFF $count=1 $X=6.04
+ $Y=0.37 $X2=6.185 $Y2=0.665
r276 3 38 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=4.7 $Y=0.625
+ $X2=4.84 $Y2=0.805
r277 2 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.095
+ $Y=0.555 $X2=2.235 $Y2=0.765
r278 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.105
+ $Y=0.37 $X2=1.245 $Y2=0.58
.ends


* File: sky130_fd_sc_ms__dlrtp_1.pxi.spice
* Created: Wed Sep  2 12:05:43 2020
* 
x_PM_SKY130_FD_SC_MS__DLRTP_1%D N_D_M1008_g N_D_M1017_g D N_D_c_137_n
+ N_D_c_138_n PM_SKY130_FD_SC_MS__DLRTP_1%D
x_PM_SKY130_FD_SC_MS__DLRTP_1%GATE N_GATE_M1006_g N_GATE_M1007_g GATE
+ N_GATE_c_165_n PM_SKY130_FD_SC_MS__DLRTP_1%GATE
x_PM_SKY130_FD_SC_MS__DLRTP_1%A_219_424# N_A_219_424#_M1007_d
+ N_A_219_424#_M1006_d N_A_219_424#_c_200_n N_A_219_424#_M1001_g
+ N_A_219_424#_M1012_g N_A_219_424#_c_217_n N_A_219_424#_M1000_g
+ N_A_219_424#_c_218_n N_A_219_424#_c_219_n N_A_219_424#_M1010_g
+ N_A_219_424#_c_204_n N_A_219_424#_c_220_n N_A_219_424#_c_205_n
+ N_A_219_424#_c_221_n N_A_219_424#_c_206_n N_A_219_424#_c_207_n
+ N_A_219_424#_c_208_n N_A_219_424#_c_209_n N_A_219_424#_c_210_n
+ N_A_219_424#_c_211_n N_A_219_424#_c_212_n N_A_219_424#_c_213_n
+ N_A_219_424#_c_214_n N_A_219_424#_c_215_n
+ PM_SKY130_FD_SC_MS__DLRTP_1%A_219_424#
x_PM_SKY130_FD_SC_MS__DLRTP_1%A_27_424# N_A_27_424#_M1017_s N_A_27_424#_M1008_s
+ N_A_27_424#_M1018_g N_A_27_424#_M1016_g N_A_27_424#_c_348_n
+ N_A_27_424#_c_354_n N_A_27_424#_c_355_n N_A_27_424#_c_356_n
+ N_A_27_424#_c_357_n N_A_27_424#_c_349_n N_A_27_424#_c_350_n
+ N_A_27_424#_c_351_n PM_SKY130_FD_SC_MS__DLRTP_1%A_27_424#
x_PM_SKY130_FD_SC_MS__DLRTP_1%A_363_74# N_A_363_74#_M1012_s N_A_363_74#_M1001_s
+ N_A_363_74#_M1019_g N_A_363_74#_M1005_g N_A_363_74#_c_433_n
+ N_A_363_74#_c_434_n N_A_363_74#_c_435_n N_A_363_74#_c_535_p
+ N_A_363_74#_c_436_n N_A_363_74#_c_443_n N_A_363_74#_c_444_n
+ N_A_363_74#_c_445_n N_A_363_74#_c_446_n N_A_363_74#_c_447_n
+ N_A_363_74#_c_478_n N_A_363_74#_c_437_n N_A_363_74#_c_438_n
+ N_A_363_74#_c_439_n PM_SKY130_FD_SC_MS__DLRTP_1%A_363_74#
x_PM_SKY130_FD_SC_MS__DLRTP_1%A_817_48# N_A_817_48#_M1015_s N_A_817_48#_M1003_d
+ N_A_817_48#_c_542_n N_A_817_48#_M1011_g N_A_817_48#_c_553_n
+ N_A_817_48#_M1013_g N_A_817_48#_c_543_n N_A_817_48#_M1014_g
+ N_A_817_48#_M1004_g N_A_817_48#_c_545_n N_A_817_48#_c_557_n
+ N_A_817_48#_c_546_n N_A_817_48#_c_558_n N_A_817_48#_c_547_n
+ N_A_817_48#_c_548_n N_A_817_48#_c_549_n N_A_817_48#_c_550_n
+ N_A_817_48#_c_559_n N_A_817_48#_c_551_n N_A_817_48#_c_552_n
+ PM_SKY130_FD_SC_MS__DLRTP_1%A_817_48#
x_PM_SKY130_FD_SC_MS__DLRTP_1%A_643_74# N_A_643_74#_M1019_d N_A_643_74#_M1000_d
+ N_A_643_74#_M1003_g N_A_643_74#_M1015_g N_A_643_74#_c_659_n
+ N_A_643_74#_c_660_n N_A_643_74#_c_661_n N_A_643_74#_c_668_n
+ N_A_643_74#_c_669_n N_A_643_74#_c_662_n N_A_643_74#_c_684_n
+ N_A_643_74#_c_670_n N_A_643_74#_c_663_n PM_SKY130_FD_SC_MS__DLRTP_1%A_643_74#
x_PM_SKY130_FD_SC_MS__DLRTP_1%RESET_B N_RESET_B_M1009_g N_RESET_B_M1002_g
+ RESET_B N_RESET_B_c_740_n N_RESET_B_c_741_n
+ PM_SKY130_FD_SC_MS__DLRTP_1%RESET_B
x_PM_SKY130_FD_SC_MS__DLRTP_1%VPWR N_VPWR_M1008_d N_VPWR_M1001_d N_VPWR_M1013_d
+ N_VPWR_M1002_d N_VPWR_c_781_n N_VPWR_c_782_n N_VPWR_c_783_n N_VPWR_c_784_n
+ N_VPWR_c_785_n VPWR N_VPWR_c_786_n N_VPWR_c_787_n N_VPWR_c_788_n
+ N_VPWR_c_789_n N_VPWR_c_780_n N_VPWR_c_791_n N_VPWR_c_792_n N_VPWR_c_793_n
+ PM_SKY130_FD_SC_MS__DLRTP_1%VPWR
x_PM_SKY130_FD_SC_MS__DLRTP_1%Q N_Q_M1014_d N_Q_M1004_d N_Q_c_863_n N_Q_c_864_n
+ N_Q_c_861_n Q PM_SKY130_FD_SC_MS__DLRTP_1%Q
x_PM_SKY130_FD_SC_MS__DLRTP_1%VGND N_VGND_M1017_d N_VGND_M1012_d N_VGND_M1011_d
+ N_VGND_M1009_d N_VGND_c_884_n N_VGND_c_885_n N_VGND_c_886_n N_VGND_c_887_n
+ N_VGND_c_888_n N_VGND_c_889_n N_VGND_c_890_n N_VGND_c_891_n N_VGND_c_892_n
+ N_VGND_c_893_n VGND N_VGND_c_894_n N_VGND_c_895_n N_VGND_c_896_n
+ N_VGND_c_897_n PM_SKY130_FD_SC_MS__DLRTP_1%VGND
cc_1 VNB N_D_M1017_g 0.0302124f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.835
cc_2 VNB N_D_c_137_n 0.00715327f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_3 VNB N_D_c_138_n 0.0657379f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.54
cc_4 VNB N_GATE_M1007_g 0.0370084f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.835
cc_5 VNB GATE 0.00257351f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_6 VNB N_GATE_c_165_n 0.024421f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.465
cc_7 VNB N_A_219_424#_c_200_n 0.0178334f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.835
cc_8 VNB N_A_219_424#_M1001_g 0.00889432f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.54
cc_9 VNB N_A_219_424#_M1012_g 0.0363752f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.3
cc_10 VNB N_A_219_424#_M1010_g 0.0350581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_219_424#_c_204_n 0.0103791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_219_424#_c_205_n 0.0100621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_219_424#_c_206_n 0.00636311f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_219_424#_c_207_n 0.00612679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_219_424#_c_208_n 0.00201944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_219_424#_c_209_n 0.0114186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_219_424#_c_210_n 0.00449969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_219_424#_c_211_n 0.00669166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_219_424#_c_212_n 0.00498474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_219_424#_c_213_n 0.0454379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_219_424#_c_214_n 0.00422813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_219_424#_c_215_n 0.0277565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_424#_M1018_g 0.0349143f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_24 VNB N_A_27_424#_c_348_n 0.00520606f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.665
cc_25 VNB N_A_27_424#_c_349_n 0.0305779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_424#_c_350_n 0.0016951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_424#_c_351_n 0.028196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_363_74#_c_433_n 0.00268395f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.3
cc_29 VNB N_A_363_74#_c_434_n 0.0198185f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.465
cc_30 VNB N_A_363_74#_c_435_n 0.00250666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_363_74#_c_436_n 0.00315036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_363_74#_c_437_n 0.0062466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_363_74#_c_438_n 0.0315985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_363_74#_c_439_n 0.0176429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_817_48#_c_542_n 0.0174955f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=0.835
cc_36 VNB N_A_817_48#_c_543_n 0.0398073f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.3
cc_37 VNB N_A_817_48#_M1004_g 0.0069424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_817_48#_c_545_n 0.0294045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_817_48#_c_546_n 0.00937344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_817_48#_c_547_n 0.0147792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_817_48#_c_548_n 0.00368394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_817_48#_c_549_n 0.0351541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_817_48#_c_550_n 0.00566982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_817_48#_c_551_n 0.00351959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_817_48#_c_552_n 0.0223702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_643_74#_M1015_g 0.0329854f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_47 VNB N_A_643_74#_c_659_n 0.0213847f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.3
cc_48 VNB N_A_643_74#_c_660_n 0.00641007f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.465
cc_49 VNB N_A_643_74#_c_661_n 0.0126245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_643_74#_c_662_n 0.00108293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_643_74#_c_663_n 0.00575851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_RESET_B_M1009_g 0.0237015f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_53 VNB N_RESET_B_c_740_n 0.0268844f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_54 VNB N_RESET_B_c_741_n 0.00165846f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.465
cc_55 VNB N_VPWR_c_780_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_Q_c_861_n 0.0390747f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.3
cc_57 VNB Q 0.030012f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.465
cc_58 VNB N_VGND_c_884_n 0.0139492f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.3
cc_59 VNB N_VGND_c_885_n 0.00396956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_886_n 0.0167618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_887_n 0.00647919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_888_n 0.0276506f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_889_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_890_n 0.0371416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_891_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_892_n 0.0306291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_893_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_894_n 0.0362066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_895_n 0.0234371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_896_n 0.394164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_897_n 0.00702378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VPB N_D_M1008_g 0.0443176f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_73 VPB N_D_c_137_n 0.00850726f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_74 VPB N_D_c_138_n 0.00693093f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.54
cc_75 VPB N_GATE_M1006_g 0.0380224f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_76 VPB N_GATE_c_165_n 0.0104858f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.465
cc_77 VPB N_A_219_424#_M1001_g 0.0295039f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.54
cc_78 VPB N_A_219_424#_c_217_n 0.0185217f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_219_424#_c_218_n 0.0305493f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_219_424#_c_219_n 0.00720675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_219_424#_c_220_n 0.011982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_219_424#_c_221_n 0.00393595f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_219_424#_c_210_n 0.00312026f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_A_219_424#_c_213_n 0.00892495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_219_424#_c_215_n 0.00937713f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_27_424#_M1016_g 0.0229223f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_87 VPB N_A_27_424#_c_348_n 0.00409706f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.665
cc_88 VPB N_A_27_424#_c_354_n 0.00887864f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_27_424#_c_355_n 0.00128303f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_27_424#_c_356_n 0.0186185f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_27_424#_c_357_n 0.0223062f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_27_424#_c_351_n 0.00568252f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_363_74#_M1005_g 0.0228797f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_94 VPB N_A_363_74#_c_433_n 0.00227193f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.3
cc_95 VPB N_A_363_74#_c_436_n 0.00230695f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_A_363_74#_c_443_n 0.00559023f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_363_74#_c_444_n 0.00198863f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_363_74#_c_445_n 0.00175682f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_363_74#_c_446_n 0.0433702f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_363_74#_c_447_n 0.00202812f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_817_48#_c_553_n 0.0321853f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_817_48#_M1013_g 0.0261338f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_103 VPB N_A_817_48#_c_543_n 0.0272317f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.3
cc_104 VPB N_A_817_48#_M1004_g 0.0303432f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_817_48#_c_557_n 0.00407784f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_817_48#_c_558_n 0.00275675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_817_48#_c_559_n 0.00766741f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_817_48#_c_551_n 0.00252622f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_643_74#_M1003_g 0.0237183f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_110 VPB N_A_643_74#_c_659_n 0.0179659f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.3
cc_111 VPB N_A_643_74#_c_660_n 0.00466185f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.465
cc_112 VPB N_A_643_74#_c_661_n 5.50244e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_643_74#_c_668_n 0.0289584f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_643_74#_c_669_n 0.00442275f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_643_74#_c_670_n 0.00292634f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_643_74#_c_663_n 0.00315245f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_RESET_B_M1002_g 0.0304708f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=0.835
cc_118 VPB N_RESET_B_c_740_n 0.00571098f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_119 VPB N_RESET_B_c_741_n 0.00383181f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.465
cc_120 VPB N_VPWR_c_781_n 0.00635773f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.3
cc_121 VPB N_VPWR_c_782_n 0.013027f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_783_n 0.0137588f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_784_n 0.0185677f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_785_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_786_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_787_n 0.0438518f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_788_n 0.0436554f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_789_n 0.0198718f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_780_n 0.0892898f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_791_n 0.00612764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_792_n 0.00699324f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_793_n 0.0176638f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_Q_c_863_n 0.0415472f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_134 VPB N_Q_c_864_n 0.0136968f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.54
cc_135 VPB N_Q_c_861_n 0.00769959f $X=-0.19 $Y=1.66 $X2=0.6 $Y2=1.3
cc_136 N_D_M1008_g N_GATE_M1006_g 0.0188194f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_137 N_D_M1017_g N_GATE_M1007_g 0.0162965f $X=0.6 $Y=0.835 $X2=0 $Y2=0
cc_138 N_D_c_138_n GATE 3.32426e-19 $X=0.505 $Y=1.54 $X2=0 $Y2=0
cc_139 N_D_c_138_n N_GATE_c_165_n 0.0264925f $X=0.505 $Y=1.54 $X2=0 $Y2=0
cc_140 N_D_M1008_g N_A_27_424#_c_348_n 0.0162003f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_141 N_D_M1017_g N_A_27_424#_c_348_n 0.00990189f $X=0.6 $Y=0.835 $X2=0 $Y2=0
cc_142 N_D_c_137_n N_A_27_424#_c_348_n 0.0343288f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_143 N_D_c_138_n N_A_27_424#_c_348_n 0.0148836f $X=0.505 $Y=1.54 $X2=0 $Y2=0
cc_144 N_D_M1008_g N_A_27_424#_c_356_n 0.00816171f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_145 N_D_M1008_g N_A_27_424#_c_357_n 0.0249256f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_146 N_D_c_137_n N_A_27_424#_c_357_n 0.0147162f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_147 N_D_c_138_n N_A_27_424#_c_357_n 0.00275637f $X=0.505 $Y=1.54 $X2=0 $Y2=0
cc_148 N_D_M1017_g N_A_27_424#_c_349_n 0.0202375f $X=0.6 $Y=0.835 $X2=0 $Y2=0
cc_149 N_D_c_137_n N_A_27_424#_c_349_n 0.0131784f $X=0.27 $Y=1.465 $X2=0 $Y2=0
cc_150 N_D_c_138_n N_A_27_424#_c_349_n 0.00817656f $X=0.505 $Y=1.54 $X2=0 $Y2=0
cc_151 N_D_M1008_g N_VPWR_c_781_n 0.00334717f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_152 N_D_M1008_g N_VPWR_c_786_n 0.005209f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_153 N_D_M1008_g N_VPWR_c_780_n 0.00520594f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_154 N_D_M1017_g N_VGND_c_884_n 0.0042545f $X=0.6 $Y=0.835 $X2=0 $Y2=0
cc_155 N_D_M1017_g N_VGND_c_888_n 0.00340649f $X=0.6 $Y=0.835 $X2=0 $Y2=0
cc_156 N_D_M1017_g N_VGND_c_896_n 0.00487769f $X=0.6 $Y=0.835 $X2=0 $Y2=0
cc_157 N_GATE_M1006_g N_A_219_424#_c_220_n 0.00615836f $X=1.005 $Y=2.54 $X2=0
+ $Y2=0
cc_158 GATE N_A_219_424#_c_220_n 0.00971996f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_159 N_GATE_c_165_n N_A_219_424#_c_220_n 0.00288243f $X=1.185 $Y=1.615 $X2=0
+ $Y2=0
cc_160 N_GATE_M1007_g N_A_219_424#_c_205_n 0.00634199f $X=1.185 $Y=0.74 $X2=0
+ $Y2=0
cc_161 N_GATE_M1006_g N_A_219_424#_c_221_n 0.0053844f $X=1.005 $Y=2.54 $X2=0
+ $Y2=0
cc_162 N_GATE_M1007_g N_A_219_424#_c_209_n 0.00469117f $X=1.185 $Y=0.74 $X2=0
+ $Y2=0
cc_163 GATE N_A_219_424#_c_209_n 0.00257643f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_164 GATE N_A_219_424#_c_210_n 0.027849f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_165 N_GATE_c_165_n N_A_219_424#_c_210_n 0.00638325f $X=1.185 $Y=1.615 $X2=0
+ $Y2=0
cc_166 N_GATE_M1007_g N_A_219_424#_c_211_n 0.00531887f $X=1.185 $Y=0.74 $X2=0
+ $Y2=0
cc_167 GATE N_A_219_424#_c_215_n 0.00100641f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_168 N_GATE_c_165_n N_A_219_424#_c_215_n 0.0181923f $X=1.185 $Y=1.615 $X2=0
+ $Y2=0
cc_169 N_GATE_M1007_g N_A_27_424#_c_348_n 0.00541079f $X=1.185 $Y=0.74 $X2=0
+ $Y2=0
cc_170 GATE N_A_27_424#_c_348_n 0.0208665f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_171 N_GATE_c_165_n N_A_27_424#_c_348_n 0.00737175f $X=1.185 $Y=1.615 $X2=0
+ $Y2=0
cc_172 N_GATE_M1006_g N_A_27_424#_c_354_n 0.0179499f $X=1.005 $Y=2.54 $X2=0
+ $Y2=0
cc_173 GATE N_A_27_424#_c_354_n 0.00480558f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_174 N_GATE_c_165_n N_A_27_424#_c_354_n 9.11879e-19 $X=1.185 $Y=1.615 $X2=0
+ $Y2=0
cc_175 N_GATE_M1006_g N_A_27_424#_c_356_n 6.13347e-19 $X=1.005 $Y=2.54 $X2=0
+ $Y2=0
cc_176 N_GATE_M1006_g N_A_27_424#_c_357_n 0.0056636f $X=1.005 $Y=2.54 $X2=0
+ $Y2=0
cc_177 N_GATE_M1006_g N_VPWR_c_781_n 0.0182479f $X=1.005 $Y=2.54 $X2=0 $Y2=0
cc_178 N_GATE_M1006_g N_VPWR_c_787_n 0.00460063f $X=1.005 $Y=2.54 $X2=0 $Y2=0
cc_179 N_GATE_M1006_g N_VPWR_c_780_n 0.0044838f $X=1.005 $Y=2.54 $X2=0 $Y2=0
cc_180 N_GATE_M1007_g N_VGND_c_884_n 0.00522565f $X=1.185 $Y=0.74 $X2=0 $Y2=0
cc_181 GATE N_VGND_c_884_n 0.00653399f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_182 N_GATE_c_165_n N_VGND_c_884_n 0.00368039f $X=1.185 $Y=1.615 $X2=0 $Y2=0
cc_183 N_GATE_M1007_g N_VGND_c_894_n 0.00434272f $X=1.185 $Y=0.74 $X2=0 $Y2=0
cc_184 N_GATE_M1007_g N_VGND_c_896_n 0.00830282f $X=1.185 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A_219_424#_M1012_g N_A_27_424#_M1018_g 0.0310105f $X=2.24 $Y=0.74 $X2=0
+ $Y2=0
cc_186 N_A_219_424#_c_206_n N_A_27_424#_M1018_g 0.0111444f $X=2.85 $Y=0.855
+ $X2=0 $Y2=0
cc_187 N_A_219_424#_c_208_n N_A_27_424#_M1018_g 0.0011351f $X=3.02 $Y=0.34 $X2=0
+ $Y2=0
cc_188 N_A_219_424#_M1001_g N_A_27_424#_M1016_g 0.0253489f $X=2.185 $Y=2.38
+ $X2=0 $Y2=0
cc_189 N_A_219_424#_c_217_n N_A_27_424#_M1016_g 0.0330636f $X=3.185 $Y=1.84
+ $X2=0 $Y2=0
cc_190 N_A_219_424#_c_220_n N_A_27_424#_c_348_n 0.00548112f $X=1.455 $Y=2.095
+ $X2=0 $Y2=0
cc_191 N_A_219_424#_M1006_d N_A_27_424#_c_354_n 0.0139832f $X=1.095 $Y=2.12
+ $X2=0 $Y2=0
cc_192 N_A_219_424#_M1001_g N_A_27_424#_c_354_n 0.0188987f $X=2.185 $Y=2.38
+ $X2=0 $Y2=0
cc_193 N_A_219_424#_c_220_n N_A_27_424#_c_354_n 0.0367029f $X=1.455 $Y=2.095
+ $X2=0 $Y2=0
cc_194 N_A_219_424#_c_210_n N_A_27_424#_c_354_n 0.00485156f $X=1.665 $Y=1.615
+ $X2=0 $Y2=0
cc_195 N_A_219_424#_c_215_n N_A_27_424#_c_354_n 0.0012498f $X=1.665 $Y=1.525
+ $X2=0 $Y2=0
cc_196 N_A_219_424#_M1001_g N_A_27_424#_c_355_n 0.00665439f $X=2.185 $Y=2.38
+ $X2=0 $Y2=0
cc_197 N_A_219_424#_c_217_n N_A_27_424#_c_355_n 2.17497e-19 $X=3.185 $Y=1.84
+ $X2=0 $Y2=0
cc_198 N_A_219_424#_c_220_n N_A_27_424#_c_357_n 0.0030406f $X=1.455 $Y=2.095
+ $X2=0 $Y2=0
cc_199 N_A_219_424#_M1001_g N_A_27_424#_c_350_n 7.12265e-19 $X=2.185 $Y=2.38
+ $X2=0 $Y2=0
cc_200 N_A_219_424#_c_204_n N_A_27_424#_c_350_n 5.7423e-19 $X=2.205 $Y=1.525
+ $X2=0 $Y2=0
cc_201 N_A_219_424#_M1001_g N_A_27_424#_c_351_n 0.00962915f $X=2.185 $Y=2.38
+ $X2=0 $Y2=0
cc_202 N_A_219_424#_c_219_n N_A_27_424#_c_351_n 0.0330636f $X=3.275 $Y=1.765
+ $X2=0 $Y2=0
cc_203 N_A_219_424#_c_204_n N_A_27_424#_c_351_n 0.00863303f $X=2.205 $Y=1.525
+ $X2=0 $Y2=0
cc_204 N_A_219_424#_c_206_n N_A_363_74#_M1012_s 0.00989832f $X=2.85 $Y=0.855
+ $X2=-0.19 $Y2=-0.245
cc_205 N_A_219_424#_c_200_n N_A_363_74#_c_433_n 0.00704085f $X=2.095 $Y=1.525
+ $X2=0 $Y2=0
cc_206 N_A_219_424#_M1001_g N_A_363_74#_c_433_n 0.0119051f $X=2.185 $Y=2.38
+ $X2=0 $Y2=0
cc_207 N_A_219_424#_M1012_g N_A_363_74#_c_433_n 0.00581595f $X=2.24 $Y=0.74
+ $X2=0 $Y2=0
cc_208 N_A_219_424#_c_204_n N_A_363_74#_c_433_n 0.00421753f $X=2.205 $Y=1.525
+ $X2=0 $Y2=0
cc_209 N_A_219_424#_c_220_n N_A_363_74#_c_433_n 0.00229419f $X=1.455 $Y=2.095
+ $X2=0 $Y2=0
cc_210 N_A_219_424#_c_221_n N_A_363_74#_c_433_n 0.00822183f $X=1.54 $Y=1.97
+ $X2=0 $Y2=0
cc_211 N_A_219_424#_c_210_n N_A_363_74#_c_433_n 0.0244847f $X=1.665 $Y=1.615
+ $X2=0 $Y2=0
cc_212 N_A_219_424#_c_211_n N_A_363_74#_c_433_n 0.00729783f $X=1.642 $Y=1.45
+ $X2=0 $Y2=0
cc_213 N_A_219_424#_c_215_n N_A_363_74#_c_433_n 0.00107984f $X=1.665 $Y=1.525
+ $X2=0 $Y2=0
cc_214 N_A_219_424#_M1012_g N_A_363_74#_c_434_n 0.0128465f $X=2.24 $Y=0.74 $X2=0
+ $Y2=0
cc_215 N_A_219_424#_c_206_n N_A_363_74#_c_434_n 0.0120886f $X=2.85 $Y=0.855
+ $X2=0 $Y2=0
cc_216 N_A_219_424#_c_200_n N_A_363_74#_c_435_n 7.98076e-19 $X=2.095 $Y=1.525
+ $X2=0 $Y2=0
cc_217 N_A_219_424#_M1012_g N_A_363_74#_c_435_n 0.00369563f $X=2.24 $Y=0.74
+ $X2=0 $Y2=0
cc_218 N_A_219_424#_c_206_n N_A_363_74#_c_435_n 0.0686872f $X=2.85 $Y=0.855
+ $X2=0 $Y2=0
cc_219 N_A_219_424#_c_209_n N_A_363_74#_c_435_n 0.0142477f $X=1.43 $Y=0.855
+ $X2=0 $Y2=0
cc_220 N_A_219_424#_c_210_n N_A_363_74#_c_435_n 0.00254949f $X=1.665 $Y=1.615
+ $X2=0 $Y2=0
cc_221 N_A_219_424#_c_215_n N_A_363_74#_c_435_n 0.00611482f $X=1.665 $Y=1.525
+ $X2=0 $Y2=0
cc_222 N_A_219_424#_c_217_n N_A_363_74#_c_436_n 0.00298724f $X=3.185 $Y=1.84
+ $X2=0 $Y2=0
cc_223 N_A_219_424#_c_219_n N_A_363_74#_c_436_n 0.00526986f $X=3.275 $Y=1.765
+ $X2=0 $Y2=0
cc_224 N_A_219_424#_c_217_n N_A_363_74#_c_443_n 0.0144279f $X=3.185 $Y=1.84
+ $X2=0 $Y2=0
cc_225 N_A_219_424#_c_217_n N_A_363_74#_c_445_n 5.09058e-19 $X=3.185 $Y=1.84
+ $X2=0 $Y2=0
cc_226 N_A_219_424#_c_217_n N_A_363_74#_c_446_n 0.0246196f $X=3.185 $Y=1.84
+ $X2=0 $Y2=0
cc_227 N_A_219_424#_c_218_n N_A_363_74#_c_446_n 0.0140765f $X=3.695 $Y=1.765
+ $X2=0 $Y2=0
cc_228 N_A_219_424#_c_213_n N_A_363_74#_c_446_n 0.00367833f $X=3.93 $Y=1.39
+ $X2=0 $Y2=0
cc_229 N_A_219_424#_c_200_n N_A_363_74#_c_447_n 0.0048198f $X=2.095 $Y=1.525
+ $X2=0 $Y2=0
cc_230 N_A_219_424#_M1001_g N_A_363_74#_c_447_n 0.00495647f $X=2.185 $Y=2.38
+ $X2=0 $Y2=0
cc_231 N_A_219_424#_c_220_n N_A_363_74#_c_447_n 0.0172708f $X=1.455 $Y=2.095
+ $X2=0 $Y2=0
cc_232 N_A_219_424#_c_210_n N_A_363_74#_c_447_n 0.00198601f $X=1.665 $Y=1.615
+ $X2=0 $Y2=0
cc_233 N_A_219_424#_c_215_n N_A_363_74#_c_447_n 2.26279e-19 $X=1.665 $Y=1.525
+ $X2=0 $Y2=0
cc_234 N_A_219_424#_c_217_n N_A_363_74#_c_478_n 0.00867708f $X=3.185 $Y=1.84
+ $X2=0 $Y2=0
cc_235 N_A_219_424#_c_219_n N_A_363_74#_c_437_n 9.2239e-19 $X=3.275 $Y=1.765
+ $X2=0 $Y2=0
cc_236 N_A_219_424#_c_219_n N_A_363_74#_c_438_n 0.0167481f $X=3.275 $Y=1.765
+ $X2=0 $Y2=0
cc_237 N_A_219_424#_M1010_g N_A_363_74#_c_438_n 0.011696f $X=3.77 $Y=0.58 $X2=0
+ $Y2=0
cc_238 N_A_219_424#_M1010_g N_A_363_74#_c_439_n 0.0168057f $X=3.77 $Y=0.58 $X2=0
+ $Y2=0
cc_239 N_A_219_424#_c_207_n N_A_363_74#_c_439_n 0.0132006f $X=3.835 $Y=0.34
+ $X2=0 $Y2=0
cc_240 N_A_219_424#_c_214_n N_A_363_74#_c_439_n 9.76507e-19 $X=3.965 $Y=1.225
+ $X2=0 $Y2=0
cc_241 N_A_219_424#_M1010_g N_A_817_48#_c_542_n 0.0385805f $X=3.77 $Y=0.58 $X2=0
+ $Y2=0
cc_242 N_A_219_424#_c_207_n N_A_817_48#_c_542_n 0.00133249f $X=3.835 $Y=0.34
+ $X2=0 $Y2=0
cc_243 N_A_219_424#_c_214_n N_A_817_48#_c_542_n 0.00729255f $X=3.965 $Y=1.225
+ $X2=0 $Y2=0
cc_244 N_A_219_424#_M1010_g N_A_817_48#_c_543_n 0.00426541f $X=3.77 $Y=0.58
+ $X2=0 $Y2=0
cc_245 N_A_219_424#_c_212_n N_A_817_48#_c_543_n 0.00197074f $X=3.93 $Y=1.39
+ $X2=0 $Y2=0
cc_246 N_A_219_424#_c_213_n N_A_817_48#_c_543_n 0.0287556f $X=3.93 $Y=1.39 $X2=0
+ $Y2=0
cc_247 N_A_219_424#_c_214_n N_A_817_48#_c_543_n 0.00399793f $X=3.965 $Y=1.225
+ $X2=0 $Y2=0
cc_248 N_A_219_424#_c_213_n N_A_817_48#_c_545_n 6.79409e-19 $X=3.93 $Y=1.39
+ $X2=0 $Y2=0
cc_249 N_A_219_424#_c_207_n N_A_643_74#_M1019_d 0.00417255f $X=3.835 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_250 N_A_219_424#_c_218_n N_A_643_74#_c_661_n 0.00639741f $X=3.695 $Y=1.765
+ $X2=0 $Y2=0
cc_251 N_A_219_424#_M1010_g N_A_643_74#_c_661_n 0.0129937f $X=3.77 $Y=0.58 $X2=0
+ $Y2=0
cc_252 N_A_219_424#_c_214_n N_A_643_74#_c_661_n 0.0457738f $X=3.965 $Y=1.225
+ $X2=0 $Y2=0
cc_253 N_A_219_424#_c_218_n N_A_643_74#_c_668_n 0.00141716f $X=3.695 $Y=1.765
+ $X2=0 $Y2=0
cc_254 N_A_219_424#_c_212_n N_A_643_74#_c_668_n 0.020194f $X=3.93 $Y=1.39 $X2=0
+ $Y2=0
cc_255 N_A_219_424#_c_213_n N_A_643_74#_c_668_n 0.0114646f $X=3.93 $Y=1.39 $X2=0
+ $Y2=0
cc_256 N_A_219_424#_c_217_n N_A_643_74#_c_669_n 0.00121322f $X=3.185 $Y=1.84
+ $X2=0 $Y2=0
cc_257 N_A_219_424#_c_218_n N_A_643_74#_c_669_n 0.0135404f $X=3.695 $Y=1.765
+ $X2=0 $Y2=0
cc_258 N_A_219_424#_M1010_g N_A_643_74#_c_662_n 0.00278503f $X=3.77 $Y=0.58
+ $X2=0 $Y2=0
cc_259 N_A_219_424#_c_207_n N_A_643_74#_c_662_n 0.0279134f $X=3.835 $Y=0.34
+ $X2=0 $Y2=0
cc_260 N_A_219_424#_c_214_n N_A_643_74#_c_662_n 0.0170435f $X=3.965 $Y=1.225
+ $X2=0 $Y2=0
cc_261 N_A_219_424#_c_217_n N_A_643_74#_c_684_n 0.00539728f $X=3.185 $Y=1.84
+ $X2=0 $Y2=0
cc_262 N_A_219_424#_c_218_n N_A_643_74#_c_684_n 0.00144029f $X=3.695 $Y=1.765
+ $X2=0 $Y2=0
cc_263 N_A_219_424#_c_217_n N_A_643_74#_c_670_n 0.00635318f $X=3.185 $Y=1.84
+ $X2=0 $Y2=0
cc_264 N_A_219_424#_c_218_n N_A_643_74#_c_670_n 0.00151884f $X=3.695 $Y=1.765
+ $X2=0 $Y2=0
cc_265 N_A_219_424#_c_212_n N_A_643_74#_c_663_n 0.00226545f $X=3.93 $Y=1.39
+ $X2=0 $Y2=0
cc_266 N_A_219_424#_M1001_g N_VPWR_c_782_n 0.00423353f $X=2.185 $Y=2.38 $X2=0
+ $Y2=0
cc_267 N_A_219_424#_c_217_n N_VPWR_c_782_n 2.77478e-19 $X=3.185 $Y=1.84 $X2=0
+ $Y2=0
cc_268 N_A_219_424#_M1001_g N_VPWR_c_787_n 0.00562877f $X=2.185 $Y=2.38 $X2=0
+ $Y2=0
cc_269 N_A_219_424#_c_217_n N_VPWR_c_788_n 0.00333926f $X=3.185 $Y=1.84 $X2=0
+ $Y2=0
cc_270 N_A_219_424#_M1001_g N_VPWR_c_780_n 0.00595788f $X=2.185 $Y=2.38 $X2=0
+ $Y2=0
cc_271 N_A_219_424#_c_217_n N_VPWR_c_780_n 0.00423366f $X=3.185 $Y=1.84 $X2=0
+ $Y2=0
cc_272 N_A_219_424#_c_206_n N_VGND_M1012_d 0.00508382f $X=2.85 $Y=0.855 $X2=0
+ $Y2=0
cc_273 N_A_219_424#_c_205_n N_VGND_c_884_n 0.0300165f $X=1.4 $Y=0.515 $X2=0
+ $Y2=0
cc_274 N_A_219_424#_M1012_g N_VGND_c_885_n 0.0126864f $X=2.24 $Y=0.74 $X2=0
+ $Y2=0
cc_275 N_A_219_424#_c_205_n N_VGND_c_885_n 0.00713841f $X=1.4 $Y=0.515 $X2=0
+ $Y2=0
cc_276 N_A_219_424#_c_206_n N_VGND_c_885_n 0.0210746f $X=2.85 $Y=0.855 $X2=0
+ $Y2=0
cc_277 N_A_219_424#_c_208_n N_VGND_c_885_n 0.0118766f $X=3.02 $Y=0.34 $X2=0
+ $Y2=0
cc_278 N_A_219_424#_M1010_g N_VGND_c_886_n 5.44443e-19 $X=3.77 $Y=0.58 $X2=0
+ $Y2=0
cc_279 N_A_219_424#_c_207_n N_VGND_c_886_n 0.0123564f $X=3.835 $Y=0.34 $X2=0
+ $Y2=0
cc_280 N_A_219_424#_c_214_n N_VGND_c_886_n 0.0246024f $X=3.965 $Y=1.225 $X2=0
+ $Y2=0
cc_281 N_A_219_424#_M1010_g N_VGND_c_890_n 0.00278262f $X=3.77 $Y=0.58 $X2=0
+ $Y2=0
cc_282 N_A_219_424#_c_207_n N_VGND_c_890_n 0.063753f $X=3.835 $Y=0.34 $X2=0
+ $Y2=0
cc_283 N_A_219_424#_c_208_n N_VGND_c_890_n 0.0121935f $X=3.02 $Y=0.34 $X2=0
+ $Y2=0
cc_284 N_A_219_424#_M1012_g N_VGND_c_894_n 0.00398535f $X=2.24 $Y=0.74 $X2=0
+ $Y2=0
cc_285 N_A_219_424#_c_205_n N_VGND_c_894_n 0.0172412f $X=1.4 $Y=0.515 $X2=0
+ $Y2=0
cc_286 N_A_219_424#_M1012_g N_VGND_c_896_n 0.00388856f $X=2.24 $Y=0.74 $X2=0
+ $Y2=0
cc_287 N_A_219_424#_M1010_g N_VGND_c_896_n 0.00354801f $X=3.77 $Y=0.58 $X2=0
+ $Y2=0
cc_288 N_A_219_424#_c_205_n N_VGND_c_896_n 0.0142144f $X=1.4 $Y=0.515 $X2=0
+ $Y2=0
cc_289 N_A_219_424#_c_206_n N_VGND_c_896_n 0.0302804f $X=2.85 $Y=0.855 $X2=0
+ $Y2=0
cc_290 N_A_219_424#_c_207_n N_VGND_c_896_n 0.0358785f $X=3.835 $Y=0.34 $X2=0
+ $Y2=0
cc_291 N_A_219_424#_c_208_n N_VGND_c_896_n 0.00661049f $X=3.02 $Y=0.34 $X2=0
+ $Y2=0
cc_292 N_A_219_424#_c_206_n A_565_74# 0.00142466f $X=2.85 $Y=0.855 $X2=-0.19
+ $Y2=-0.245
cc_293 N_A_219_424#_c_207_n A_769_74# 5.0299e-19 $X=3.835 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_294 N_A_219_424#_c_214_n A_769_74# 0.003195f $X=3.965 $Y=1.225 $X2=-0.19
+ $Y2=-0.245
cc_295 N_A_27_424#_c_354_n N_A_363_74#_M1001_s 0.00750563f $X=2.525 $Y=2.475
+ $X2=0 $Y2=0
cc_296 N_A_27_424#_M1018_g N_A_363_74#_c_433_n 8.66064e-19 $X=2.75 $Y=0.69 $X2=0
+ $Y2=0
cc_297 N_A_27_424#_M1016_g N_A_363_74#_c_433_n 2.02362e-19 $X=2.765 $Y=2.46
+ $X2=0 $Y2=0
cc_298 N_A_27_424#_c_350_n N_A_363_74#_c_433_n 0.0220207f $X=2.69 $Y=1.635 $X2=0
+ $Y2=0
cc_299 N_A_27_424#_c_351_n N_A_363_74#_c_433_n 0.00100444f $X=2.69 $Y=1.635
+ $X2=0 $Y2=0
cc_300 N_A_27_424#_M1018_g N_A_363_74#_c_434_n 0.0101442f $X=2.75 $Y=0.69 $X2=0
+ $Y2=0
cc_301 N_A_27_424#_c_350_n N_A_363_74#_c_434_n 0.0228816f $X=2.69 $Y=1.635 $X2=0
+ $Y2=0
cc_302 N_A_27_424#_c_351_n N_A_363_74#_c_434_n 0.00122248f $X=2.69 $Y=1.635
+ $X2=0 $Y2=0
cc_303 N_A_27_424#_c_355_n N_A_363_74#_c_436_n 0.00738713f $X=2.61 $Y=2.39 $X2=0
+ $Y2=0
cc_304 N_A_27_424#_c_350_n N_A_363_74#_c_436_n 0.0248017f $X=2.69 $Y=1.635 $X2=0
+ $Y2=0
cc_305 N_A_27_424#_c_351_n N_A_363_74#_c_436_n 0.00674601f $X=2.69 $Y=1.635
+ $X2=0 $Y2=0
cc_306 N_A_27_424#_M1016_g N_A_363_74#_c_444_n 0.0011745f $X=2.765 $Y=2.46 $X2=0
+ $Y2=0
cc_307 N_A_27_424#_c_354_n N_A_363_74#_c_447_n 0.0230002f $X=2.525 $Y=2.475
+ $X2=0 $Y2=0
cc_308 N_A_27_424#_c_355_n N_A_363_74#_c_447_n 0.0084011f $X=2.61 $Y=2.39 $X2=0
+ $Y2=0
cc_309 N_A_27_424#_M1018_g N_A_363_74#_c_437_n 0.0044995f $X=2.75 $Y=0.69 $X2=0
+ $Y2=0
cc_310 N_A_27_424#_M1018_g N_A_363_74#_c_439_n 0.0597211f $X=2.75 $Y=0.69 $X2=0
+ $Y2=0
cc_311 N_A_27_424#_c_354_n N_VPWR_M1008_d 0.0068978f $X=2.525 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_312 N_A_27_424#_c_357_n N_VPWR_M1008_d 0.00432546f $X=0.715 $Y=2.33 $X2=-0.19
+ $Y2=-0.245
cc_313 N_A_27_424#_c_354_n N_VPWR_M1001_d 0.0106965f $X=2.525 $Y=2.475 $X2=0
+ $Y2=0
cc_314 N_A_27_424#_c_355_n N_VPWR_M1001_d 0.00511383f $X=2.61 $Y=2.39 $X2=0
+ $Y2=0
cc_315 N_A_27_424#_c_356_n N_VPWR_c_781_n 0.0101711f $X=0.28 $Y=2.265 $X2=0
+ $Y2=0
cc_316 N_A_27_424#_c_357_n N_VPWR_c_781_n 0.0187086f $X=0.715 $Y=2.33 $X2=0
+ $Y2=0
cc_317 N_A_27_424#_M1016_g N_VPWR_c_782_n 0.00838194f $X=2.765 $Y=2.46 $X2=0
+ $Y2=0
cc_318 N_A_27_424#_c_354_n N_VPWR_c_782_n 0.0249123f $X=2.525 $Y=2.475 $X2=0
+ $Y2=0
cc_319 N_A_27_424#_c_356_n N_VPWR_c_786_n 0.0140571f $X=0.28 $Y=2.265 $X2=0
+ $Y2=0
cc_320 N_A_27_424#_M1016_g N_VPWR_c_788_n 0.00460063f $X=2.765 $Y=2.46 $X2=0
+ $Y2=0
cc_321 N_A_27_424#_M1016_g N_VPWR_c_780_n 0.00908371f $X=2.765 $Y=2.46 $X2=0
+ $Y2=0
cc_322 N_A_27_424#_c_354_n N_VPWR_c_780_n 0.0506441f $X=2.525 $Y=2.475 $X2=0
+ $Y2=0
cc_323 N_A_27_424#_c_356_n N_VPWR_c_780_n 0.011784f $X=0.28 $Y=2.265 $X2=0 $Y2=0
cc_324 N_A_27_424#_c_357_n N_VPWR_c_780_n 0.00701323f $X=0.715 $Y=2.33 $X2=0
+ $Y2=0
cc_325 N_A_27_424#_c_349_n N_VGND_c_884_n 0.0230738f $X=0.63 $Y=0.835 $X2=0
+ $Y2=0
cc_326 N_A_27_424#_M1018_g N_VGND_c_885_n 0.00507404f $X=2.75 $Y=0.69 $X2=0
+ $Y2=0
cc_327 N_A_27_424#_c_349_n N_VGND_c_888_n 0.0118661f $X=0.63 $Y=0.835 $X2=0
+ $Y2=0
cc_328 N_A_27_424#_M1018_g N_VGND_c_890_n 0.00444681f $X=2.75 $Y=0.69 $X2=0
+ $Y2=0
cc_329 N_A_27_424#_M1018_g N_VGND_c_896_n 0.00427328f $X=2.75 $Y=0.69 $X2=0
+ $Y2=0
cc_330 N_A_27_424#_c_349_n N_VGND_c_896_n 0.0158184f $X=0.63 $Y=0.835 $X2=0
+ $Y2=0
cc_331 N_A_363_74#_c_445_n N_A_817_48#_c_553_n 7.79074e-19 $X=3.88 $Y=2.215
+ $X2=0 $Y2=0
cc_332 N_A_363_74#_c_446_n N_A_817_48#_c_553_n 0.0170379f $X=3.88 $Y=2.215 $X2=0
+ $Y2=0
cc_333 N_A_363_74#_M1005_g N_A_817_48#_M1013_g 0.013785f $X=3.72 $Y=2.75 $X2=0
+ $Y2=0
cc_334 N_A_363_74#_c_443_n N_A_817_48#_M1013_g 0.00177596f $X=3.715 $Y=2.99
+ $X2=0 $Y2=0
cc_335 N_A_363_74#_c_445_n N_A_817_48#_M1013_g 0.00877775f $X=3.88 $Y=2.215
+ $X2=0 $Y2=0
cc_336 N_A_363_74#_c_445_n N_A_817_48#_c_557_n 0.0177637f $X=3.88 $Y=2.215 $X2=0
+ $Y2=0
cc_337 N_A_363_74#_c_446_n N_A_817_48#_c_557_n 0.00120301f $X=3.88 $Y=2.215
+ $X2=0 $Y2=0
cc_338 N_A_363_74#_c_443_n N_A_643_74#_M1000_d 0.00363537f $X=3.715 $Y=2.99
+ $X2=0 $Y2=0
cc_339 N_A_363_74#_c_436_n N_A_643_74#_c_661_n 0.0136696f $X=3.11 $Y=1.97 $X2=0
+ $Y2=0
cc_340 N_A_363_74#_c_437_n N_A_643_74#_c_661_n 0.0254068f $X=3.175 $Y=1.195
+ $X2=0 $Y2=0
cc_341 N_A_363_74#_c_438_n N_A_643_74#_c_661_n 0.00244597f $X=3.23 $Y=1.285
+ $X2=0 $Y2=0
cc_342 N_A_363_74#_c_439_n N_A_643_74#_c_661_n 0.00351644f $X=3.23 $Y=1.12 $X2=0
+ $Y2=0
cc_343 N_A_363_74#_c_445_n N_A_643_74#_c_668_n 0.0262119f $X=3.88 $Y=2.215 $X2=0
+ $Y2=0
cc_344 N_A_363_74#_c_436_n N_A_643_74#_c_669_n 0.0130064f $X=3.11 $Y=1.97 $X2=0
+ $Y2=0
cc_345 N_A_363_74#_c_446_n N_A_643_74#_c_669_n 0.00437073f $X=3.88 $Y=2.215
+ $X2=0 $Y2=0
cc_346 N_A_363_74#_c_437_n N_A_643_74#_c_662_n 0.00806711f $X=3.175 $Y=1.195
+ $X2=0 $Y2=0
cc_347 N_A_363_74#_c_438_n N_A_643_74#_c_662_n 0.00341895f $X=3.23 $Y=1.285
+ $X2=0 $Y2=0
cc_348 N_A_363_74#_c_439_n N_A_643_74#_c_662_n 0.00935059f $X=3.23 $Y=1.12 $X2=0
+ $Y2=0
cc_349 N_A_363_74#_M1005_g N_A_643_74#_c_684_n 0.00297227f $X=3.72 $Y=2.75 $X2=0
+ $Y2=0
cc_350 N_A_363_74#_c_443_n N_A_643_74#_c_684_n 0.0171624f $X=3.715 $Y=2.99 $X2=0
+ $Y2=0
cc_351 N_A_363_74#_c_436_n N_A_643_74#_c_670_n 0.00535063f $X=3.11 $Y=1.97 $X2=0
+ $Y2=0
cc_352 N_A_363_74#_c_445_n N_A_643_74#_c_670_n 0.0482167f $X=3.88 $Y=2.215 $X2=0
+ $Y2=0
cc_353 N_A_363_74#_c_446_n N_A_643_74#_c_670_n 0.00297227f $X=3.88 $Y=2.215
+ $X2=0 $Y2=0
cc_354 N_A_363_74#_c_478_n N_A_643_74#_c_670_n 0.0123438f $X=3.11 $Y=2.055 $X2=0
+ $Y2=0
cc_355 N_A_363_74#_c_444_n N_VPWR_c_782_n 0.0104713f $X=3.075 $Y=2.99 $X2=0
+ $Y2=0
cc_356 N_A_363_74#_M1005_g N_VPWR_c_788_n 0.00333833f $X=3.72 $Y=2.75 $X2=0
+ $Y2=0
cc_357 N_A_363_74#_c_443_n N_VPWR_c_788_n 0.063691f $X=3.715 $Y=2.99 $X2=0 $Y2=0
cc_358 N_A_363_74#_c_444_n N_VPWR_c_788_n 0.0121867f $X=3.075 $Y=2.99 $X2=0
+ $Y2=0
cc_359 N_A_363_74#_M1005_g N_VPWR_c_780_n 0.00425285f $X=3.72 $Y=2.75 $X2=0
+ $Y2=0
cc_360 N_A_363_74#_c_443_n N_VPWR_c_780_n 0.0352395f $X=3.715 $Y=2.99 $X2=0
+ $Y2=0
cc_361 N_A_363_74#_c_444_n N_VPWR_c_780_n 0.00660921f $X=3.075 $Y=2.99 $X2=0
+ $Y2=0
cc_362 N_A_363_74#_M1005_g N_VPWR_c_793_n 4.05858e-19 $X=3.72 $Y=2.75 $X2=0
+ $Y2=0
cc_363 N_A_363_74#_c_443_n N_VPWR_c_793_n 0.00796896f $X=3.715 $Y=2.99 $X2=0
+ $Y2=0
cc_364 N_A_363_74#_c_445_n N_VPWR_c_793_n 0.0109521f $X=3.88 $Y=2.215 $X2=0
+ $Y2=0
cc_365 N_A_363_74#_c_535_p A_571_392# 0.00327032f $X=2.99 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_366 N_A_363_74#_c_478_n A_571_392# 0.00478419f $X=3.11 $Y=2.055 $X2=-0.19
+ $Y2=-0.245
cc_367 N_A_363_74#_c_443_n A_762_508# 8.66307e-19 $X=3.715 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_368 N_A_363_74#_c_445_n A_762_508# 0.00564058f $X=3.88 $Y=2.215 $X2=-0.19
+ $Y2=-0.245
cc_369 N_A_363_74#_c_439_n N_VGND_c_885_n 2.63324e-19 $X=3.23 $Y=1.12 $X2=0
+ $Y2=0
cc_370 N_A_363_74#_c_439_n N_VGND_c_890_n 0.00278271f $X=3.23 $Y=1.12 $X2=0
+ $Y2=0
cc_371 N_A_363_74#_c_439_n N_VGND_c_896_n 0.00354802f $X=3.23 $Y=1.12 $X2=0
+ $Y2=0
cc_372 N_A_817_48#_c_553_n N_A_643_74#_M1003_g 0.00893844f $X=4.375 $Y=2.38
+ $X2=0 $Y2=0
cc_373 N_A_817_48#_M1013_g N_A_643_74#_M1003_g 0.0136165f $X=4.375 $Y=2.75 $X2=0
+ $Y2=0
cc_374 N_A_817_48#_c_543_n N_A_643_74#_M1003_g 0.00448135f $X=4.38 $Y=2.05 $X2=0
+ $Y2=0
cc_375 N_A_817_48#_c_557_n N_A_643_74#_M1003_g 0.0111402f $X=5.095 $Y=2.222
+ $X2=0 $Y2=0
cc_376 N_A_817_48#_c_559_n N_A_643_74#_M1003_g 0.0151752f $X=5.41 $Y=2.115 $X2=0
+ $Y2=0
cc_377 N_A_817_48#_c_551_n N_A_643_74#_M1003_g 0.00408593f $X=5.335 $Y=1.95
+ $X2=0 $Y2=0
cc_378 N_A_817_48#_c_545_n N_A_643_74#_M1015_g 0.00808109f $X=4.38 $Y=0.94 $X2=0
+ $Y2=0
cc_379 N_A_817_48#_c_546_n N_A_643_74#_M1015_g 0.012954f $X=4.935 $Y=0.515 $X2=0
+ $Y2=0
cc_380 N_A_817_48#_c_550_n N_A_643_74#_M1015_g 0.0127642f $X=5.017 $Y=1.095
+ $X2=0 $Y2=0
cc_381 N_A_817_48#_c_551_n N_A_643_74#_M1015_g 0.009378f $X=5.335 $Y=1.95 $X2=0
+ $Y2=0
cc_382 N_A_817_48#_c_543_n N_A_643_74#_c_659_n 0.0217577f $X=4.38 $Y=2.05 $X2=0
+ $Y2=0
cc_383 N_A_817_48#_c_557_n N_A_643_74#_c_659_n 0.00483936f $X=5.095 $Y=2.222
+ $X2=0 $Y2=0
cc_384 N_A_817_48#_c_550_n N_A_643_74#_c_659_n 0.00713037f $X=5.017 $Y=1.095
+ $X2=0 $Y2=0
cc_385 N_A_817_48#_c_551_n N_A_643_74#_c_660_n 0.0095273f $X=5.335 $Y=1.95 $X2=0
+ $Y2=0
cc_386 N_A_817_48#_c_553_n N_A_643_74#_c_668_n 0.00484368f $X=4.375 $Y=2.38
+ $X2=0 $Y2=0
cc_387 N_A_817_48#_c_543_n N_A_643_74#_c_668_n 0.0162584f $X=4.38 $Y=2.05 $X2=0
+ $Y2=0
cc_388 N_A_817_48#_c_557_n N_A_643_74#_c_668_n 0.0265217f $X=5.095 $Y=2.222
+ $X2=0 $Y2=0
cc_389 N_A_817_48#_c_543_n N_A_643_74#_c_663_n 0.00167264f $X=4.38 $Y=2.05 $X2=0
+ $Y2=0
cc_390 N_A_817_48#_c_557_n N_A_643_74#_c_663_n 0.0217299f $X=5.095 $Y=2.222
+ $X2=0 $Y2=0
cc_391 N_A_817_48#_c_550_n N_A_643_74#_c_663_n 0.00890275f $X=5.017 $Y=1.095
+ $X2=0 $Y2=0
cc_392 N_A_817_48#_c_551_n N_A_643_74#_c_663_n 0.0301206f $X=5.335 $Y=1.95 $X2=0
+ $Y2=0
cc_393 N_A_817_48#_c_546_n N_RESET_B_M1009_g 0.00222669f $X=4.935 $Y=0.515 $X2=0
+ $Y2=0
cc_394 N_A_817_48#_c_547_n N_RESET_B_M1009_g 0.0144185f $X=5.975 $Y=1.095 $X2=0
+ $Y2=0
cc_395 N_A_817_48#_c_548_n N_RESET_B_M1009_g 9.9568e-19 $X=6.14 $Y=1.385 $X2=0
+ $Y2=0
cc_396 N_A_817_48#_c_551_n N_RESET_B_M1009_g 0.00330038f $X=5.335 $Y=1.95 $X2=0
+ $Y2=0
cc_397 N_A_817_48#_c_552_n N_RESET_B_M1009_g 0.0290173f $X=6.14 $Y=1.22 $X2=0
+ $Y2=0
cc_398 N_A_817_48#_M1004_g N_RESET_B_M1002_g 0.0219072f $X=6.215 $Y=2.4 $X2=0
+ $Y2=0
cc_399 N_A_817_48#_c_558_n N_RESET_B_M1002_g 0.00732239f $X=5.41 $Y=2.465 $X2=0
+ $Y2=0
cc_400 N_A_817_48#_c_559_n N_RESET_B_M1002_g 0.00543339f $X=5.41 $Y=2.115 $X2=0
+ $Y2=0
cc_401 N_A_817_48#_c_551_n N_RESET_B_M1002_g 0.00339594f $X=5.335 $Y=1.95 $X2=0
+ $Y2=0
cc_402 N_A_817_48#_M1004_g N_RESET_B_c_740_n 0.0048174f $X=6.215 $Y=2.4 $X2=0
+ $Y2=0
cc_403 N_A_817_48#_c_547_n N_RESET_B_c_740_n 0.00124445f $X=5.975 $Y=1.095 $X2=0
+ $Y2=0
cc_404 N_A_817_48#_c_548_n N_RESET_B_c_740_n 6.9668e-19 $X=6.14 $Y=1.385 $X2=0
+ $Y2=0
cc_405 N_A_817_48#_c_549_n N_RESET_B_c_740_n 0.0121881f $X=6.14 $Y=1.385 $X2=0
+ $Y2=0
cc_406 N_A_817_48#_c_559_n N_RESET_B_c_740_n 6.64736e-19 $X=5.41 $Y=2.115 $X2=0
+ $Y2=0
cc_407 N_A_817_48#_c_551_n N_RESET_B_c_740_n 0.00174016f $X=5.335 $Y=1.95 $X2=0
+ $Y2=0
cc_408 N_A_817_48#_M1004_g N_RESET_B_c_741_n 0.00276707f $X=6.215 $Y=2.4 $X2=0
+ $Y2=0
cc_409 N_A_817_48#_c_547_n N_RESET_B_c_741_n 0.0247205f $X=5.975 $Y=1.095 $X2=0
+ $Y2=0
cc_410 N_A_817_48#_c_548_n N_RESET_B_c_741_n 0.0126449f $X=6.14 $Y=1.385 $X2=0
+ $Y2=0
cc_411 N_A_817_48#_c_549_n N_RESET_B_c_741_n 6.96581e-19 $X=6.14 $Y=1.385 $X2=0
+ $Y2=0
cc_412 N_A_817_48#_c_559_n N_RESET_B_c_741_n 0.0122442f $X=5.41 $Y=2.115 $X2=0
+ $Y2=0
cc_413 N_A_817_48#_c_551_n N_RESET_B_c_741_n 0.0327282f $X=5.335 $Y=1.95 $X2=0
+ $Y2=0
cc_414 N_A_817_48#_c_557_n N_VPWR_M1013_d 0.00544476f $X=5.095 $Y=2.222 $X2=0
+ $Y2=0
cc_415 N_A_817_48#_M1004_g N_VPWR_c_783_n 0.00943875f $X=6.215 $Y=2.4 $X2=0
+ $Y2=0
cc_416 N_A_817_48#_c_548_n N_VPWR_c_783_n 0.00419693f $X=6.14 $Y=1.385 $X2=0
+ $Y2=0
cc_417 N_A_817_48#_c_549_n N_VPWR_c_783_n 6.59514e-19 $X=6.14 $Y=1.385 $X2=0
+ $Y2=0
cc_418 N_A_817_48#_c_559_n N_VPWR_c_783_n 0.0407271f $X=5.41 $Y=2.115 $X2=0
+ $Y2=0
cc_419 N_A_817_48#_c_558_n N_VPWR_c_784_n 0.014549f $X=5.41 $Y=2.465 $X2=0 $Y2=0
cc_420 N_A_817_48#_M1013_g N_VPWR_c_788_n 0.00461464f $X=4.375 $Y=2.75 $X2=0
+ $Y2=0
cc_421 N_A_817_48#_M1004_g N_VPWR_c_789_n 0.005209f $X=6.215 $Y=2.4 $X2=0 $Y2=0
cc_422 N_A_817_48#_M1013_g N_VPWR_c_780_n 0.00910297f $X=4.375 $Y=2.75 $X2=0
+ $Y2=0
cc_423 N_A_817_48#_M1004_g N_VPWR_c_780_n 0.00987222f $X=6.215 $Y=2.4 $X2=0
+ $Y2=0
cc_424 N_A_817_48#_c_558_n N_VPWR_c_780_n 0.0119743f $X=5.41 $Y=2.465 $X2=0
+ $Y2=0
cc_425 N_A_817_48#_c_553_n N_VPWR_c_793_n 0.00352628f $X=4.375 $Y=2.38 $X2=0
+ $Y2=0
cc_426 N_A_817_48#_M1013_g N_VPWR_c_793_n 0.0169705f $X=4.375 $Y=2.75 $X2=0
+ $Y2=0
cc_427 N_A_817_48#_c_557_n N_VPWR_c_793_n 0.0327169f $X=5.095 $Y=2.222 $X2=0
+ $Y2=0
cc_428 N_A_817_48#_c_558_n N_VPWR_c_793_n 0.0144922f $X=5.41 $Y=2.465 $X2=0
+ $Y2=0
cc_429 N_A_817_48#_c_547_n N_Q_M1014_d 0.00234008f $X=5.975 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_430 N_A_817_48#_M1004_g N_Q_c_863_n 0.013562f $X=6.215 $Y=2.4 $X2=0 $Y2=0
cc_431 N_A_817_48#_M1004_g N_Q_c_864_n 0.00463751f $X=6.215 $Y=2.4 $X2=0 $Y2=0
cc_432 N_A_817_48#_c_548_n N_Q_c_864_n 0.00103105f $X=6.14 $Y=1.385 $X2=0 $Y2=0
cc_433 N_A_817_48#_c_547_n N_Q_c_861_n 0.0141806f $X=5.975 $Y=1.095 $X2=0 $Y2=0
cc_434 N_A_817_48#_c_548_n N_Q_c_861_n 0.0278652f $X=6.14 $Y=1.385 $X2=0 $Y2=0
cc_435 N_A_817_48#_c_549_n N_Q_c_861_n 0.0152417f $X=6.14 $Y=1.385 $X2=0 $Y2=0
cc_436 N_A_817_48#_c_552_n N_Q_c_861_n 0.00443182f $X=6.14 $Y=1.22 $X2=0 $Y2=0
cc_437 N_A_817_48#_c_547_n Q 0.0116838f $X=5.975 $Y=1.095 $X2=0 $Y2=0
cc_438 N_A_817_48#_c_549_n Q 0.00107479f $X=6.14 $Y=1.385 $X2=0 $Y2=0
cc_439 N_A_817_48#_c_552_n Q 0.00864397f $X=6.14 $Y=1.22 $X2=0 $Y2=0
cc_440 N_A_817_48#_c_547_n N_VGND_M1009_d 0.00261503f $X=5.975 $Y=1.095 $X2=0
+ $Y2=0
cc_441 N_A_817_48#_c_542_n N_VGND_c_886_n 0.0115327f $X=4.16 $Y=0.865 $X2=0
+ $Y2=0
cc_442 N_A_817_48#_c_545_n N_VGND_c_886_n 0.01149f $X=4.38 $Y=0.94 $X2=0 $Y2=0
cc_443 N_A_817_48#_c_546_n N_VGND_c_886_n 0.0310125f $X=4.935 $Y=0.515 $X2=0
+ $Y2=0
cc_444 N_A_817_48#_c_546_n N_VGND_c_887_n 0.0155235f $X=4.935 $Y=0.515 $X2=0
+ $Y2=0
cc_445 N_A_817_48#_c_547_n N_VGND_c_887_n 0.0218003f $X=5.975 $Y=1.095 $X2=0
+ $Y2=0
cc_446 N_A_817_48#_c_552_n N_VGND_c_887_n 0.00569497f $X=6.14 $Y=1.22 $X2=0
+ $Y2=0
cc_447 N_A_817_48#_c_542_n N_VGND_c_890_n 0.00383152f $X=4.16 $Y=0.865 $X2=0
+ $Y2=0
cc_448 N_A_817_48#_c_546_n N_VGND_c_892_n 0.0145639f $X=4.935 $Y=0.515 $X2=0
+ $Y2=0
cc_449 N_A_817_48#_c_552_n N_VGND_c_895_n 0.00434272f $X=6.14 $Y=1.22 $X2=0
+ $Y2=0
cc_450 N_A_817_48#_c_542_n N_VGND_c_896_n 0.0075725f $X=4.16 $Y=0.865 $X2=0
+ $Y2=0
cc_451 N_A_817_48#_c_546_n N_VGND_c_896_n 0.0119984f $X=4.935 $Y=0.515 $X2=0
+ $Y2=0
cc_452 N_A_817_48#_c_552_n N_VGND_c_896_n 0.00825201f $X=6.14 $Y=1.22 $X2=0
+ $Y2=0
cc_453 N_A_817_48#_c_547_n A_1045_74# 0.0048076f $X=5.975 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_454 N_A_643_74#_M1015_g N_RESET_B_M1009_g 0.0564763f $X=5.15 $Y=0.74 $X2=0
+ $Y2=0
cc_455 N_A_643_74#_c_660_n N_RESET_B_M1002_g 0.0148633f $X=5.135 $Y=1.635 $X2=0
+ $Y2=0
cc_456 N_A_643_74#_M1015_g N_RESET_B_c_740_n 0.020603f $X=5.15 $Y=0.74 $X2=0
+ $Y2=0
cc_457 N_A_643_74#_M1015_g N_RESET_B_c_741_n 3.79805e-19 $X=5.15 $Y=0.74 $X2=0
+ $Y2=0
cc_458 N_A_643_74#_c_660_n N_RESET_B_c_741_n 3.27182e-19 $X=5.135 $Y=1.635 $X2=0
+ $Y2=0
cc_459 N_A_643_74#_M1003_g N_VPWR_c_784_n 0.00461464f $X=5.135 $Y=2.46 $X2=0
+ $Y2=0
cc_460 N_A_643_74#_M1003_g N_VPWR_c_780_n 0.00909121f $X=5.135 $Y=2.46 $X2=0
+ $Y2=0
cc_461 N_A_643_74#_M1003_g N_VPWR_c_793_n 0.0155569f $X=5.135 $Y=2.46 $X2=0
+ $Y2=0
cc_462 N_A_643_74#_M1015_g N_VGND_c_886_n 0.00370782f $X=5.15 $Y=0.74 $X2=0
+ $Y2=0
cc_463 N_A_643_74#_M1015_g N_VGND_c_887_n 0.00194806f $X=5.15 $Y=0.74 $X2=0
+ $Y2=0
cc_464 N_A_643_74#_M1015_g N_VGND_c_892_n 0.00434272f $X=5.15 $Y=0.74 $X2=0
+ $Y2=0
cc_465 N_A_643_74#_M1015_g N_VGND_c_896_n 0.00825979f $X=5.15 $Y=0.74 $X2=0
+ $Y2=0
cc_466 N_RESET_B_M1002_g N_VPWR_c_783_n 0.00218742f $X=5.635 $Y=2.46 $X2=0 $Y2=0
cc_467 N_RESET_B_c_741_n N_VPWR_c_783_n 0.00163024f $X=5.6 $Y=1.515 $X2=0 $Y2=0
cc_468 N_RESET_B_M1002_g N_VPWR_c_784_n 0.005209f $X=5.635 $Y=2.46 $X2=0 $Y2=0
cc_469 N_RESET_B_M1002_g N_VPWR_c_780_n 0.00983375f $X=5.635 $Y=2.46 $X2=0 $Y2=0
cc_470 N_RESET_B_M1002_g N_VPWR_c_793_n 4.25103e-19 $X=5.635 $Y=2.46 $X2=0 $Y2=0
cc_471 N_RESET_B_M1002_g N_Q_c_864_n 8.22245e-19 $X=5.635 $Y=2.46 $X2=0 $Y2=0
cc_472 N_RESET_B_M1009_g N_VGND_c_887_n 0.0138667f $X=5.54 $Y=0.74 $X2=0 $Y2=0
cc_473 N_RESET_B_M1009_g N_VGND_c_892_n 0.00383152f $X=5.54 $Y=0.74 $X2=0 $Y2=0
cc_474 N_RESET_B_M1009_g N_VGND_c_896_n 0.0075725f $X=5.54 $Y=0.74 $X2=0 $Y2=0
cc_475 N_VPWR_c_789_n N_Q_c_863_n 0.0158876f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_476 N_VPWR_c_780_n N_Q_c_863_n 0.0130823f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_477 N_VPWR_c_783_n N_Q_c_864_n 0.0350603f $X=5.91 $Y=2.115 $X2=0 $Y2=0
cc_478 Q N_VGND_c_887_n 0.0196681f $X=6.395 $Y=0.47 $X2=0 $Y2=0
cc_479 Q N_VGND_c_895_n 0.0233346f $X=6.395 $Y=0.47 $X2=0 $Y2=0
cc_480 Q N_VGND_c_896_n 0.0194239f $X=6.395 $Y=0.47 $X2=0 $Y2=0

* NGSPICE file created from sky130_fd_sc_ms__or2_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__or2_1 A B VGND VNB VPB VPWR X
M1000 X a_63_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=5.7345e+11p ps=4.42e+06u
M1001 a_155_368# B a_63_368# VPB pshort w=840000u l=180000u
+  ad=2.016e+11p pd=2.16e+06u as=2.352e+11p ps=2.24e+06u
M1002 VGND A a_63_368# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=2.6125e+11p ps=2.05e+06u
M1003 a_63_368# B VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_63_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=6.398e+11p ps=3.46e+06u
M1005 VPWR A a_155_368# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


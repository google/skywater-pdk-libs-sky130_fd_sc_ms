* File: sky130_fd_sc_ms__nor2_4.spice
* Created: Fri Aug 28 17:46:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nor2_4.pex.spice"
.subckt sky130_fd_sc_ms__nor2_4  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_M1002_g N_Y_M1002_s VNB NLOWVT L=0.15 W=0.74 AD=0.2294
+ AS=0.4218 PD=2.1 PS=1.88 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2 SB=75003.5
+ A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g N_Y_M1002_s VNB NLOWVT L=0.15 W=0.74 AD=0.1221
+ AS=0.4218 PD=1.07 PS=1.88 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5 SB=75002.2
+ A=0.111 P=1.78 MULT=1
MM1005 N_Y_M1005_d N_B_M1005_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.74 AD=0.111
+ AS=0.1221 PD=1.04 PS=1.07 NRD=3.24 NRS=8.1 M=1 R=4.93333 SA=75002 SB=75001.7
+ A=0.111 P=1.78 MULT=1
MM1011 N_Y_M1005_d N_B_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.74 AD=0.111
+ AS=1.0138 PD=1.04 PS=4.22 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.5 SB=75001.3
+ A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_27_368#_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003.5 A=0.2016 P=2.6 MULT=1
MM1001 N_VPWR_M1000_d N_A_M1001_g N_A_27_368#_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90003 A=0.2016 P=2.6 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_A_27_368#_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90002.6 A=0.2016 P=2.6 MULT=1
MM1006 N_VPWR_M1003_d N_A_M1006_g N_A_27_368#_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90002.1 A=0.2016 P=2.6 MULT=1
MM1007 N_Y_M1007_d N_B_M1007_g N_A_27_368#_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1008 N_Y_M1007_d N_B_M1008_g N_A_27_368#_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.4
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1009 N_Y_M1009_d N_B_M1009_g N_A_27_368#_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90002.9
+ SB=90000.8 A=0.2016 P=2.6 MULT=1
MM1010 N_Y_M1009_d N_B_M1010_g N_A_27_368#_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.3808 PD=1.44 PS=2.92 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.4
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__nor2_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__mux2_2.pxi.spice
* Created: Wed Sep  2 12:11:46 2020
* 
x_PM_SKY130_FD_SC_MS__MUX2_2%A0 N_A0_M1000_g N_A0_c_96_n N_A0_M1002_g A0
+ N_A0_c_98_n PM_SKY130_FD_SC_MS__MUX2_2%A0
x_PM_SKY130_FD_SC_MS__MUX2_2%A1 N_A1_M1001_g N_A1_c_122_n N_A1_M1006_g A1
+ N_A1_c_123_n N_A1_c_124_n PM_SKY130_FD_SC_MS__MUX2_2%A1
x_PM_SKY130_FD_SC_MS__MUX2_2%S N_S_M1009_g N_S_M1007_g N_S_M1008_g N_S_M1012_g
+ N_S_c_158_n N_S_c_159_n N_S_c_160_n N_S_c_161_n N_S_c_162_n N_S_c_163_n S
+ N_S_c_164_n N_S_c_165_n S PM_SKY130_FD_SC_MS__MUX2_2%S
x_PM_SKY130_FD_SC_MS__MUX2_2%A_459_48# N_A_459_48#_M1012_s N_A_459_48#_M1008_s
+ N_A_459_48#_M1004_g N_A_459_48#_M1005_g N_A_459_48#_c_251_n
+ N_A_459_48#_c_252_n N_A_459_48#_c_253_n N_A_459_48#_c_254_n
+ N_A_459_48#_c_255_n N_A_459_48#_c_256_n N_A_459_48#_c_257_n
+ PM_SKY130_FD_SC_MS__MUX2_2%A_459_48#
x_PM_SKY130_FD_SC_MS__MUX2_2%A_119_368# N_A_119_368#_M1002_d
+ N_A_119_368#_M1000_d N_A_119_368#_M1010_g N_A_119_368#_M1003_g
+ N_A_119_368#_M1011_g N_A_119_368#_M1013_g N_A_119_368#_c_329_n
+ N_A_119_368#_c_335_n N_A_119_368#_c_385_p N_A_119_368#_c_346_n
+ N_A_119_368#_c_336_n N_A_119_368#_c_330_n N_A_119_368#_c_338_n
+ N_A_119_368#_c_339_n N_A_119_368#_c_340_n N_A_119_368#_c_341_n
+ N_A_119_368#_c_331_n N_A_119_368#_c_332_n N_A_119_368#_c_343_n
+ PM_SKY130_FD_SC_MS__MUX2_2%A_119_368#
x_PM_SKY130_FD_SC_MS__MUX2_2%A_27_368# N_A_27_368#_M1000_s N_A_27_368#_M1007_s
+ N_A_27_368#_c_431_n N_A_27_368#_c_432_n N_A_27_368#_c_433_n
+ N_A_27_368#_c_434_n PM_SKY130_FD_SC_MS__MUX2_2%A_27_368#
x_PM_SKY130_FD_SC_MS__MUX2_2%A_209_368# N_A_209_368#_M1001_d
+ N_A_209_368#_M1005_d N_A_209_368#_c_461_n N_A_209_368#_c_462_n
+ N_A_209_368#_c_463_n PM_SKY130_FD_SC_MS__MUX2_2%A_209_368#
x_PM_SKY130_FD_SC_MS__MUX2_2%VPWR N_VPWR_M1007_d N_VPWR_M1008_d N_VPWR_M1011_s
+ N_VPWR_c_491_n N_VPWR_c_492_n N_VPWR_c_493_n N_VPWR_c_494_n VPWR
+ N_VPWR_c_495_n N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_498_n N_VPWR_c_499_n
+ N_VPWR_c_490_n PM_SKY130_FD_SC_MS__MUX2_2%VPWR
x_PM_SKY130_FD_SC_MS__MUX2_2%X N_X_M1003_d N_X_M1010_d X X X
+ PM_SKY130_FD_SC_MS__MUX2_2%X
x_PM_SKY130_FD_SC_MS__MUX2_2%A_38_74# N_A_38_74#_M1002_s N_A_38_74#_M1004_d
+ N_A_38_74#_c_560_n N_A_38_74#_c_561_n N_A_38_74#_c_562_n N_A_38_74#_c_563_n
+ PM_SKY130_FD_SC_MS__MUX2_2%A_38_74#
x_PM_SKY130_FD_SC_MS__MUX2_2%VGND N_VGND_M1009_d N_VGND_M1012_d N_VGND_M1013_s
+ N_VGND_c_592_n N_VGND_c_593_n N_VGND_c_594_n N_VGND_c_595_n N_VGND_c_596_n
+ N_VGND_c_597_n N_VGND_c_598_n N_VGND_c_599_n VGND N_VGND_c_600_n
+ N_VGND_c_601_n N_VGND_c_602_n N_VGND_c_603_n PM_SKY130_FD_SC_MS__MUX2_2%VGND
cc_1 VNB N_A0_M1000_g 0.00936933f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.34
cc_2 VNB N_A0_c_96_n 0.0235456f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.22
cc_3 VNB A0 0.0103228f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A0_c_98_n 0.0604963f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.385
cc_5 VNB N_A1_M1001_g 0.00711076f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.34
cc_6 VNB N_A1_c_122_n 0.0187368f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.22
cc_7 VNB N_A1_c_123_n 0.0094737f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.385
cc_8 VNB N_A1_c_124_n 0.0444529f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.385
cc_9 VNB N_S_M1009_g 0.0325126f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.34
cc_10 VNB N_S_M1008_g 0.0137951f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_11 VNB N_S_M1012_g 0.0278673f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.385
cc_12 VNB N_S_c_158_n 0.0545147f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_13 VNB N_S_c_159_n 0.0155165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_S_c_160_n 0.00209218f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_15 VNB N_S_c_161_n 0.0140564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_S_c_162_n 0.0032759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_S_c_163_n 0.0109028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_S_c_164_n 0.0266077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_S_c_165_n 0.00231439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_459_48#_M1004_g 0.0375502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_459_48#_c_251_n 0.0043718f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.385
cc_22 VNB N_A_459_48#_c_252_n 0.00686707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_459_48#_c_253_n 0.00304223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_459_48#_c_254_n 0.00275007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_459_48#_c_255_n 0.00893193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_459_48#_c_256_n 0.00444253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_459_48#_c_257_n 0.0395517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_119_368#_M1010_g 0.00334301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_119_368#_M1003_g 0.0203836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_119_368#_M1011_g 0.00155254f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_31 VNB N_A_119_368#_M1013_g 0.0261234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_119_368#_c_329_n 0.0324906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_119_368#_c_330_n 0.01098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_119_368#_c_331_n 0.00436702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_119_368#_c_332_n 0.0514256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_490_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB X 0.00406431f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.74
cc_38 VNB N_A_38_74#_c_560_n 0.0209651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_38_74#_c_561_n 0.011561f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_40 VNB N_A_38_74#_c_562_n 0.00971514f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_41 VNB N_A_38_74#_c_563_n 0.00639207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_592_n 0.0117029f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_43 VNB N_VGND_c_593_n 0.0177565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_594_n 0.00577157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_595_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_596_n 0.0436438f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_47 VNB N_VGND_c_597_n 0.00279755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_598_n 0.07498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_599_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_600_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_601_n 0.0190307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_602_n 0.00729102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_603_n 0.305923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VPB N_A0_M1000_g 0.0284706f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.34
cc_55 VPB N_A1_M1001_g 0.0248477f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.34
cc_56 VPB N_S_M1007_g 0.0273367f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=0.74
cc_57 VPB N_S_M1008_g 0.0297276f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_58 VPB N_S_c_160_n 0.00236019f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_59 VPB N_S_c_164_n 0.0184547f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_S_c_165_n 0.00153509f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_A_459_48#_M1005_g 0.0314275f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_459_48#_c_251_n 0.00673795f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=1.385
cc_63 VPB N_A_459_48#_c_253_n 0.00258775f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_A_459_48#_c_254_n 0.0096756f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_459_48#_c_257_n 0.02195f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_119_368#_M1010_g 0.0229649f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_119_368#_M1011_g 0.0239122f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_68 VPB N_A_119_368#_c_335_n 0.00262435f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_119_368#_c_336_n 0.00452416f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_119_368#_c_330_n 0.00382251f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_119_368#_c_338_n 0.0119692f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_A_119_368#_c_339_n 0.00508827f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_119_368#_c_340_n 0.0143097f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_119_368#_c_341_n 0.00562225f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_119_368#_c_331_n 0.0259151f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_119_368#_c_343_n 0.00555493f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_27_368#_c_431_n 0.043538f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_27_368#_c_432_n 0.0202059f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_27_368#_c_433_n 0.0100805f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.385
cc_80 VPB N_A_27_368#_c_434_n 0.0066409f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_209_368#_c_461_n 0.0071967f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=0.74
cc_82 VPB N_A_209_368#_c_462_n 0.00415706f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_83 VPB N_A_209_368#_c_463_n 0.00262741f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_84 VPB N_VPWR_c_491_n 0.00928913f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_85 VPB N_VPWR_c_492_n 0.0164699f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_493_n 0.0130546f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_494_n 0.0221025f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_88 VPB N_VPWR_c_495_n 0.0512348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_496_n 0.0445926f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_497_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_498_n 0.00631825f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_499_n 0.00631974f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_490_n 0.0857431f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB X 0.00127169f $X=-0.19 $Y=1.66 $X2=0.55 $Y2=0.74
cc_95 N_A0_M1000_g N_A1_M1001_g 0.0314411f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_96 N_A0_c_96_n N_A1_c_122_n 0.0189176f $X=0.55 $Y=1.22 $X2=0 $Y2=0
cc_97 N_A0_c_96_n N_A1_c_123_n 0.00206978f $X=0.55 $Y=1.22 $X2=0 $Y2=0
cc_98 A0 N_A1_c_123_n 0.029162f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_99 N_A0_c_98_n N_A1_c_123_n 0.00941047f $X=0.55 $Y=1.385 $X2=0 $Y2=0
cc_100 A0 N_A1_c_124_n 2.04426e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_101 N_A0_c_98_n N_A1_c_124_n 0.0182447f $X=0.55 $Y=1.385 $X2=0 $Y2=0
cc_102 N_A0_M1000_g N_A_119_368#_c_335_n 2.91588e-19 $X=0.505 $Y=2.34 $X2=0
+ $Y2=0
cc_103 N_A0_M1000_g N_A_27_368#_c_431_n 0.0159776f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_104 A0 N_A_27_368#_c_431_n 0.0188569f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_105 N_A0_c_98_n N_A_27_368#_c_431_n 0.00223195f $X=0.55 $Y=1.385 $X2=0 $Y2=0
cc_106 N_A0_M1000_g N_A_27_368#_c_432_n 0.0106481f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_107 N_A0_M1000_g N_A_27_368#_c_433_n 0.00198263f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_108 N_A0_M1000_g N_VPWR_c_495_n 8.89343e-19 $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_109 N_A0_c_96_n N_A_38_74#_c_560_n 0.0142246f $X=0.55 $Y=1.22 $X2=0 $Y2=0
cc_110 A0 N_A_38_74#_c_560_n 0.022507f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_111 N_A0_c_98_n N_A_38_74#_c_560_n 0.00182108f $X=0.55 $Y=1.385 $X2=0 $Y2=0
cc_112 N_A0_c_96_n N_A_38_74#_c_561_n 0.0114763f $X=0.55 $Y=1.22 $X2=0 $Y2=0
cc_113 N_A0_c_96_n N_A_38_74#_c_562_n 0.00215133f $X=0.55 $Y=1.22 $X2=0 $Y2=0
cc_114 N_A0_c_96_n N_VGND_c_598_n 0.00283294f $X=0.55 $Y=1.22 $X2=0 $Y2=0
cc_115 N_A0_c_96_n N_VGND_c_603_n 0.00360528f $X=0.55 $Y=1.22 $X2=0 $Y2=0
cc_116 N_A1_c_122_n N_S_M1009_g 0.0331815f $X=1.275 $Y=1.22 $X2=0 $Y2=0
cc_117 N_A1_M1001_g N_S_c_164_n 0.00339876f $X=0.955 $Y=2.34 $X2=0 $Y2=0
cc_118 N_A1_c_124_n N_S_c_164_n 0.0331815f $X=1.275 $Y=1.385 $X2=0 $Y2=0
cc_119 N_A1_c_123_n N_A_119_368#_c_335_n 0.0141814f $X=1.03 $Y=1.385 $X2=0 $Y2=0
cc_120 N_A1_c_122_n N_A_119_368#_c_346_n 0.0221735f $X=1.275 $Y=1.22 $X2=0 $Y2=0
cc_121 N_A1_c_123_n N_A_119_368#_c_346_n 0.040728f $X=1.03 $Y=1.385 $X2=0 $Y2=0
cc_122 N_A1_c_124_n N_A_119_368#_c_346_n 0.00205655f $X=1.275 $Y=1.385 $X2=0
+ $Y2=0
cc_123 N_A1_M1001_g N_A_119_368#_c_336_n 0.023718f $X=0.955 $Y=2.34 $X2=0 $Y2=0
cc_124 N_A1_c_123_n N_A_119_368#_c_336_n 0.0193447f $X=1.03 $Y=1.385 $X2=0 $Y2=0
cc_125 N_A1_c_124_n N_A_119_368#_c_336_n 0.0093449f $X=1.275 $Y=1.385 $X2=0
+ $Y2=0
cc_126 N_A1_M1001_g N_A_119_368#_c_330_n 0.00564738f $X=0.955 $Y=2.34 $X2=0
+ $Y2=0
cc_127 N_A1_c_122_n N_A_119_368#_c_330_n 0.00512335f $X=1.275 $Y=1.22 $X2=0
+ $Y2=0
cc_128 N_A1_c_123_n N_A_119_368#_c_330_n 0.0292455f $X=1.03 $Y=1.385 $X2=0 $Y2=0
cc_129 N_A1_M1001_g N_A_27_368#_c_431_n 0.00102926f $X=0.955 $Y=2.34 $X2=0 $Y2=0
cc_130 N_A1_M1001_g N_A_27_368#_c_432_n 0.013283f $X=0.955 $Y=2.34 $X2=0 $Y2=0
cc_131 N_A1_M1001_g N_A_27_368#_c_434_n 0.00477191f $X=0.955 $Y=2.34 $X2=0 $Y2=0
cc_132 N_A1_M1001_g N_A_209_368#_c_462_n 0.00638486f $X=0.955 $Y=2.34 $X2=0
+ $Y2=0
cc_133 N_A1_M1001_g N_VPWR_c_495_n 8.71493e-19 $X=0.955 $Y=2.34 $X2=0 $Y2=0
cc_134 N_A1_c_122_n N_A_38_74#_c_561_n 0.010644f $X=1.275 $Y=1.22 $X2=0 $Y2=0
cc_135 N_A1_c_122_n N_VGND_c_597_n 2.11353e-19 $X=1.275 $Y=1.22 $X2=0 $Y2=0
cc_136 N_A1_c_122_n N_VGND_c_598_n 0.00283318f $X=1.275 $Y=1.22 $X2=0 $Y2=0
cc_137 N_A1_c_122_n N_VGND_c_603_n 0.00356414f $X=1.275 $Y=1.22 $X2=0 $Y2=0
cc_138 N_S_M1009_g N_A_459_48#_M1004_g 0.019636f $X=1.665 $Y=0.74 $X2=0 $Y2=0
cc_139 N_S_c_158_n N_A_459_48#_M1004_g 0.00509439f $X=3.635 $Y=1.295 $X2=0 $Y2=0
cc_140 N_S_c_160_n N_A_459_48#_M1004_g 0.00944274f $X=2.3 $Y=1.45 $X2=0 $Y2=0
cc_141 N_S_c_161_n N_A_459_48#_M1004_g 0.00666396f $X=3.125 $Y=1.215 $X2=0 $Y2=0
cc_142 N_S_c_162_n N_A_459_48#_M1004_g 0.00452171f $X=2.385 $Y=1.215 $X2=0 $Y2=0
cc_143 N_S_c_163_n N_A_459_48#_M1004_g 8.44761e-19 $X=3.29 $Y=1.215 $X2=0 $Y2=0
cc_144 N_S_c_164_n N_A_459_48#_M1004_g 0.00936723f $X=1.965 $Y=1.615 $X2=0 $Y2=0
cc_145 N_S_M1007_g N_A_459_48#_M1005_g 0.0189686f $X=1.965 $Y=2.46 $X2=0 $Y2=0
cc_146 N_S_M1008_g N_A_459_48#_c_251_n 5.82299e-19 $X=3.725 $Y=2.26 $X2=0 $Y2=0
cc_147 N_S_c_158_n N_A_459_48#_c_251_n 0.00147334f $X=3.635 $Y=1.295 $X2=0 $Y2=0
cc_148 N_S_c_161_n N_A_459_48#_c_251_n 0.0114196f $X=3.125 $Y=1.215 $X2=0 $Y2=0
cc_149 N_S_c_163_n N_A_459_48#_c_251_n 0.0157852f $X=3.29 $Y=1.215 $X2=0 $Y2=0
cc_150 N_S_M1012_g N_A_459_48#_c_252_n 0.00826909f $X=3.72 $Y=0.645 $X2=0 $Y2=0
cc_151 N_S_c_160_n N_A_459_48#_c_253_n 0.0254342f $X=2.3 $Y=1.45 $X2=0 $Y2=0
cc_152 N_S_c_161_n N_A_459_48#_c_253_n 0.0247729f $X=3.125 $Y=1.215 $X2=0 $Y2=0
cc_153 N_S_c_164_n N_A_459_48#_c_253_n 2.79763e-19 $X=1.965 $Y=1.615 $X2=0 $Y2=0
cc_154 N_S_M1008_g N_A_459_48#_c_254_n 0.0166639f $X=3.725 $Y=2.26 $X2=0 $Y2=0
cc_155 N_S_c_158_n N_A_459_48#_c_254_n 0.00819338f $X=3.635 $Y=1.295 $X2=0 $Y2=0
cc_156 N_S_c_163_n N_A_459_48#_c_254_n 0.00976597f $X=3.29 $Y=1.215 $X2=0 $Y2=0
cc_157 N_S_M1008_g N_A_459_48#_c_255_n 0.006214f $X=3.725 $Y=2.26 $X2=0 $Y2=0
cc_158 N_S_M1012_g N_A_459_48#_c_255_n 0.00663605f $X=3.72 $Y=0.645 $X2=0 $Y2=0
cc_159 N_S_c_158_n N_A_459_48#_c_255_n 0.00513851f $X=3.635 $Y=1.295 $X2=0 $Y2=0
cc_160 N_S_c_159_n N_A_459_48#_c_255_n 0.00687432f $X=3.725 $Y=1.295 $X2=0 $Y2=0
cc_161 N_S_c_163_n N_A_459_48#_c_255_n 0.0235661f $X=3.29 $Y=1.215 $X2=0 $Y2=0
cc_162 N_S_M1012_g N_A_459_48#_c_256_n 0.00826577f $X=3.72 $Y=0.645 $X2=0 $Y2=0
cc_163 N_S_c_158_n N_A_459_48#_c_256_n 0.00812293f $X=3.635 $Y=1.295 $X2=0 $Y2=0
cc_164 N_S_c_163_n N_A_459_48#_c_256_n 0.00870045f $X=3.29 $Y=1.215 $X2=0 $Y2=0
cc_165 N_S_c_160_n N_A_459_48#_c_257_n 0.00835613f $X=2.3 $Y=1.45 $X2=0 $Y2=0
cc_166 N_S_c_161_n N_A_459_48#_c_257_n 0.00578023f $X=3.125 $Y=1.215 $X2=0 $Y2=0
cc_167 N_S_c_164_n N_A_459_48#_c_257_n 0.0189686f $X=1.965 $Y=1.615 $X2=0 $Y2=0
cc_168 N_S_M1008_g N_A_119_368#_M1010_g 0.0201474f $X=3.725 $Y=2.26 $X2=0 $Y2=0
cc_169 N_S_M1012_g N_A_119_368#_M1003_g 0.0173258f $X=3.72 $Y=0.645 $X2=0 $Y2=0
cc_170 N_S_c_159_n N_A_119_368#_M1003_g 0.00887935f $X=3.725 $Y=1.295 $X2=0
+ $Y2=0
cc_171 N_S_c_159_n N_A_119_368#_c_329_n 0.0201474f $X=3.725 $Y=1.295 $X2=0 $Y2=0
cc_172 N_S_M1009_g N_A_119_368#_c_330_n 0.0116106f $X=1.665 $Y=0.74 $X2=0 $Y2=0
cc_173 N_S_M1007_g N_A_119_368#_c_330_n 0.00113754f $X=1.965 $Y=2.46 $X2=0 $Y2=0
cc_174 N_S_c_165_n N_A_119_368#_c_330_n 0.0250633f $X=2.215 $Y=1.615 $X2=0 $Y2=0
cc_175 N_S_M1007_g N_A_119_368#_c_338_n 0.0144312f $X=1.965 $Y=2.46 $X2=0 $Y2=0
cc_176 N_S_c_160_n N_A_119_368#_c_338_n 0.0124173f $X=2.3 $Y=1.45 $X2=0 $Y2=0
cc_177 N_S_c_161_n N_A_119_368#_c_338_n 0.00365018f $X=3.125 $Y=1.215 $X2=0
+ $Y2=0
cc_178 N_S_c_164_n N_A_119_368#_c_338_n 0.00858175f $X=1.965 $Y=1.615 $X2=0
+ $Y2=0
cc_179 N_S_c_165_n N_A_119_368#_c_338_n 0.0302603f $X=2.215 $Y=1.615 $X2=0 $Y2=0
cc_180 N_S_M1008_g N_A_119_368#_c_339_n 0.0033455f $X=3.725 $Y=2.26 $X2=0 $Y2=0
cc_181 N_S_M1008_g N_A_119_368#_c_340_n 0.016296f $X=3.725 $Y=2.26 $X2=0 $Y2=0
cc_182 N_S_M1007_g N_A_119_368#_c_343_n 0.00523517f $X=1.965 $Y=2.46 $X2=0 $Y2=0
cc_183 N_S_M1007_g N_A_27_368#_c_432_n 3.96096e-19 $X=1.965 $Y=2.46 $X2=0 $Y2=0
cc_184 N_S_M1007_g N_A_27_368#_c_434_n 0.00764577f $X=1.965 $Y=2.46 $X2=0 $Y2=0
cc_185 N_S_M1007_g N_A_209_368#_c_461_n 0.0154966f $X=1.965 $Y=2.46 $X2=0 $Y2=0
cc_186 N_S_M1007_g N_A_209_368#_c_462_n 0.00444581f $X=1.965 $Y=2.46 $X2=0 $Y2=0
cc_187 N_S_M1007_g N_A_209_368#_c_463_n 7.78134e-19 $X=1.965 $Y=2.46 $X2=0 $Y2=0
cc_188 N_S_M1007_g N_VPWR_c_491_n 0.00150765f $X=1.965 $Y=2.46 $X2=0 $Y2=0
cc_189 N_S_M1008_g N_VPWR_c_492_n 0.00385696f $X=3.725 $Y=2.26 $X2=0 $Y2=0
cc_190 N_S_M1007_g N_VPWR_c_495_n 0.00518311f $X=1.965 $Y=2.46 $X2=0 $Y2=0
cc_191 N_S_M1008_g N_VPWR_c_496_n 0.00482866f $X=3.725 $Y=2.26 $X2=0 $Y2=0
cc_192 N_S_M1007_g N_VPWR_c_490_n 0.00541438f $X=1.965 $Y=2.46 $X2=0 $Y2=0
cc_193 N_S_M1008_g N_VPWR_c_490_n 0.00555093f $X=3.725 $Y=2.26 $X2=0 $Y2=0
cc_194 N_S_M1012_g X 0.00278223f $X=3.72 $Y=0.645 $X2=0 $Y2=0
cc_195 N_S_c_159_n X 0.00848135f $X=3.725 $Y=1.295 $X2=0 $Y2=0
cc_196 N_S_M1009_g N_A_38_74#_c_561_n 0.0142791f $X=1.665 $Y=0.74 $X2=0 $Y2=0
cc_197 N_S_M1009_g N_A_38_74#_c_563_n 7.54552e-19 $X=1.665 $Y=0.74 $X2=0 $Y2=0
cc_198 N_S_M1012_g N_VGND_c_592_n 9.12408e-19 $X=3.72 $Y=0.645 $X2=0 $Y2=0
cc_199 N_S_c_158_n N_VGND_c_592_n 3.48248e-19 $X=3.635 $Y=1.295 $X2=0 $Y2=0
cc_200 N_S_c_161_n N_VGND_c_592_n 0.0538813f $X=3.125 $Y=1.215 $X2=0 $Y2=0
cc_201 N_S_c_162_n N_VGND_c_592_n 0.0113758f $X=2.385 $Y=1.215 $X2=0 $Y2=0
cc_202 N_S_c_163_n N_VGND_c_592_n 0.00372877f $X=3.29 $Y=1.215 $X2=0 $Y2=0
cc_203 N_S_c_164_n N_VGND_c_592_n 2.04362e-19 $X=1.965 $Y=1.615 $X2=0 $Y2=0
cc_204 N_S_c_165_n N_VGND_c_592_n 0.0061623f $X=2.215 $Y=1.615 $X2=0 $Y2=0
cc_205 N_S_M1012_g N_VGND_c_593_n 0.00257181f $X=3.72 $Y=0.645 $X2=0 $Y2=0
cc_206 N_S_M1012_g N_VGND_c_594_n 0.00341131f $X=3.72 $Y=0.645 $X2=0 $Y2=0
cc_207 N_S_M1009_g N_VGND_c_597_n 0.00470661f $X=1.665 $Y=0.74 $X2=0 $Y2=0
cc_208 N_S_c_164_n N_VGND_c_597_n 0.00685793f $X=1.965 $Y=1.615 $X2=0 $Y2=0
cc_209 N_S_c_165_n N_VGND_c_597_n 0.0162068f $X=2.215 $Y=1.615 $X2=0 $Y2=0
cc_210 N_S_M1009_g N_VGND_c_598_n 0.00283318f $X=1.665 $Y=0.74 $X2=0 $Y2=0
cc_211 N_S_M1012_g N_VGND_c_600_n 0.00434272f $X=3.72 $Y=0.645 $X2=0 $Y2=0
cc_212 N_S_M1009_g N_VGND_c_603_n 0.00356303f $X=1.665 $Y=0.74 $X2=0 $Y2=0
cc_213 N_S_M1012_g N_VGND_c_603_n 0.00434731f $X=3.72 $Y=0.645 $X2=0 $Y2=0
cc_214 N_A_459_48#_c_254_n N_A_119_368#_M1010_g 3.09569e-19 $X=3.565 $Y=1.715
+ $X2=0 $Y2=0
cc_215 N_A_459_48#_c_252_n N_A_119_368#_M1003_g 5.66031e-19 $X=3.505 $Y=0.645
+ $X2=0 $Y2=0
cc_216 N_A_459_48#_c_256_n N_A_119_368#_M1003_g 3.01611e-19 $X=3.567 $Y=0.94
+ $X2=0 $Y2=0
cc_217 N_A_459_48#_c_255_n N_A_119_368#_c_329_n 6.11181e-19 $X=3.565 $Y=1.63
+ $X2=0 $Y2=0
cc_218 N_A_459_48#_M1005_g N_A_119_368#_c_338_n 0.0157388f $X=2.515 $Y=2.46
+ $X2=0 $Y2=0
cc_219 N_A_459_48#_c_251_n N_A_119_368#_c_338_n 0.022268f $X=3.335 $Y=1.715
+ $X2=0 $Y2=0
cc_220 N_A_459_48#_c_253_n N_A_119_368#_c_338_n 0.0221432f $X=2.72 $Y=1.635
+ $X2=0 $Y2=0
cc_221 N_A_459_48#_c_254_n N_A_119_368#_c_338_n 0.0154042f $X=3.565 $Y=1.715
+ $X2=0 $Y2=0
cc_222 N_A_459_48#_c_257_n N_A_119_368#_c_338_n 0.00223579f $X=2.515 $Y=1.635
+ $X2=0 $Y2=0
cc_223 N_A_459_48#_M1005_g N_A_119_368#_c_339_n 0.00426053f $X=2.515 $Y=2.46
+ $X2=0 $Y2=0
cc_224 N_A_459_48#_M1008_s N_A_119_368#_c_340_n 0.00782185f $X=3.355 $Y=1.84
+ $X2=0 $Y2=0
cc_225 N_A_459_48#_c_251_n N_A_119_368#_c_340_n 0.00596701f $X=3.335 $Y=1.715
+ $X2=0 $Y2=0
cc_226 N_A_459_48#_c_254_n N_A_119_368#_c_340_n 0.0313619f $X=3.565 $Y=1.715
+ $X2=0 $Y2=0
cc_227 N_A_459_48#_M1005_g N_A_209_368#_c_461_n 0.0103147f $X=2.515 $Y=2.46
+ $X2=0 $Y2=0
cc_228 N_A_459_48#_M1005_g N_A_209_368#_c_463_n 0.00864019f $X=2.515 $Y=2.46
+ $X2=0 $Y2=0
cc_229 N_A_459_48#_M1005_g N_VPWR_c_491_n 0.00343717f $X=2.515 $Y=2.46 $X2=0
+ $Y2=0
cc_230 N_A_459_48#_M1005_g N_VPWR_c_496_n 0.005209f $X=2.515 $Y=2.46 $X2=0 $Y2=0
cc_231 N_A_459_48#_M1005_g N_VPWR_c_490_n 0.00540854f $X=2.515 $Y=2.46 $X2=0
+ $Y2=0
cc_232 N_A_459_48#_c_256_n X 0.11361f $X=3.567 $Y=0.94 $X2=0 $Y2=0
cc_233 N_A_459_48#_M1004_g N_A_38_74#_c_561_n 0.00894316f $X=2.37 $Y=0.74 $X2=0
+ $Y2=0
cc_234 N_A_459_48#_M1004_g N_A_38_74#_c_563_n 0.00658239f $X=2.37 $Y=0.74 $X2=0
+ $Y2=0
cc_235 N_A_459_48#_M1004_g N_VGND_c_592_n 0.0136534f $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A_459_48#_c_256_n N_VGND_c_592_n 0.013581f $X=3.567 $Y=0.94 $X2=0 $Y2=0
cc_237 N_A_459_48#_M1004_g N_VGND_c_593_n 0.0048753f $X=2.37 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A_459_48#_c_252_n N_VGND_c_593_n 0.0348474f $X=3.505 $Y=0.645 $X2=0
+ $Y2=0
cc_239 N_A_459_48#_c_252_n N_VGND_c_594_n 0.0101913f $X=3.505 $Y=0.645 $X2=0
+ $Y2=0
cc_240 N_A_459_48#_M1004_g N_VGND_c_597_n 0.00427381f $X=2.37 $Y=0.74 $X2=0
+ $Y2=0
cc_241 N_A_459_48#_M1004_g N_VGND_c_598_n 0.00284483f $X=2.37 $Y=0.74 $X2=0
+ $Y2=0
cc_242 N_A_459_48#_c_252_n N_VGND_c_600_n 0.0144337f $X=3.505 $Y=0.645 $X2=0
+ $Y2=0
cc_243 N_A_459_48#_M1004_g N_VGND_c_603_n 0.00360668f $X=2.37 $Y=0.74 $X2=0
+ $Y2=0
cc_244 N_A_459_48#_c_252_n N_VGND_c_603_n 0.0119481f $X=3.505 $Y=0.645 $X2=0
+ $Y2=0
cc_245 N_A_459_48#_c_256_n N_VGND_c_603_n 0.00423403f $X=3.567 $Y=0.94 $X2=0
+ $Y2=0
cc_246 N_A_119_368#_c_338_n N_A_27_368#_M1007_s 0.00562297f $X=2.995 $Y=2.055
+ $X2=0 $Y2=0
cc_247 N_A_119_368#_c_335_n N_A_27_368#_c_431_n 0.0122403f $X=0.73 $Y=2.14 $X2=0
+ $Y2=0
cc_248 N_A_119_368#_c_385_p N_A_27_368#_c_432_n 0.0137665f $X=0.73 $Y=2.56 $X2=0
+ $Y2=0
cc_249 N_A_119_368#_c_336_n N_A_209_368#_M1001_d 0.00407211f $X=1.365 $Y=1.98
+ $X2=-0.19 $Y2=-0.245
cc_250 N_A_119_368#_c_338_n N_A_209_368#_M1005_d 0.00675599f $X=2.995 $Y=2.055
+ $X2=0 $Y2=0
cc_251 N_A_119_368#_c_336_n N_A_209_368#_c_461_n 0.0015404f $X=1.365 $Y=1.98
+ $X2=0 $Y2=0
cc_252 N_A_119_368#_c_338_n N_A_209_368#_c_461_n 0.0616054f $X=2.995 $Y=2.055
+ $X2=0 $Y2=0
cc_253 N_A_119_368#_c_343_n N_A_209_368#_c_461_n 0.014265f $X=1.45 $Y=1.98 $X2=0
+ $Y2=0
cc_254 N_A_119_368#_c_336_n N_A_209_368#_c_462_n 0.0221185f $X=1.365 $Y=1.98
+ $X2=0 $Y2=0
cc_255 N_A_119_368#_c_338_n N_A_209_368#_c_463_n 0.015486f $X=2.995 $Y=2.055
+ $X2=0 $Y2=0
cc_256 N_A_119_368#_c_341_n N_A_209_368#_c_463_n 0.0156276f $X=3.165 $Y=2.395
+ $X2=0 $Y2=0
cc_257 N_A_119_368#_c_338_n N_VPWR_M1007_d 0.00554554f $X=2.995 $Y=2.055
+ $X2=-0.19 $Y2=-0.245
cc_258 N_A_119_368#_c_340_n N_VPWR_M1008_d 0.00793599f $X=4.835 $Y=2.395 $X2=0
+ $Y2=0
cc_259 N_A_119_368#_c_340_n N_VPWR_M1011_s 0.00449534f $X=4.835 $Y=2.395 $X2=0
+ $Y2=0
cc_260 N_A_119_368#_c_331_n N_VPWR_M1011_s 0.00600484f $X=5 $Y=1.465 $X2=0 $Y2=0
cc_261 N_A_119_368#_M1010_g N_VPWR_c_492_n 0.0120324f $X=4.27 $Y=2.4 $X2=0 $Y2=0
cc_262 N_A_119_368#_M1011_g N_VPWR_c_492_n 0.00128716f $X=4.72 $Y=2.4 $X2=0
+ $Y2=0
cc_263 N_A_119_368#_c_340_n N_VPWR_c_492_n 0.0221109f $X=4.835 $Y=2.395 $X2=0
+ $Y2=0
cc_264 N_A_119_368#_M1010_g N_VPWR_c_494_n 0.00128618f $X=4.27 $Y=2.4 $X2=0
+ $Y2=0
cc_265 N_A_119_368#_M1011_g N_VPWR_c_494_n 0.0121155f $X=4.72 $Y=2.4 $X2=0 $Y2=0
cc_266 N_A_119_368#_c_340_n N_VPWR_c_494_n 0.0283433f $X=4.835 $Y=2.395 $X2=0
+ $Y2=0
cc_267 N_A_119_368#_M1010_g N_VPWR_c_497_n 0.00460063f $X=4.27 $Y=2.4 $X2=0
+ $Y2=0
cc_268 N_A_119_368#_M1011_g N_VPWR_c_497_n 0.00460063f $X=4.72 $Y=2.4 $X2=0
+ $Y2=0
cc_269 N_A_119_368#_M1010_g N_VPWR_c_490_n 0.00463365f $X=4.27 $Y=2.4 $X2=0
+ $Y2=0
cc_270 N_A_119_368#_M1011_g N_VPWR_c_490_n 0.00463365f $X=4.72 $Y=2.4 $X2=0
+ $Y2=0
cc_271 N_A_119_368#_c_340_n N_VPWR_c_490_n 0.0433812f $X=4.835 $Y=2.395 $X2=0
+ $Y2=0
cc_272 N_A_119_368#_c_341_n N_VPWR_c_490_n 0.00645828f $X=3.165 $Y=2.395 $X2=0
+ $Y2=0
cc_273 N_A_119_368#_c_340_n N_X_M1010_d 0.00482128f $X=4.835 $Y=2.395 $X2=0
+ $Y2=0
cc_274 N_A_119_368#_M1010_g X 0.0206049f $X=4.27 $Y=2.4 $X2=0 $Y2=0
cc_275 N_A_119_368#_M1003_g X 0.0196086f $X=4.285 $Y=0.74 $X2=0 $Y2=0
cc_276 N_A_119_368#_M1011_g X 0.00901246f $X=4.72 $Y=2.4 $X2=0 $Y2=0
cc_277 N_A_119_368#_M1013_g X 0.0145881f $X=4.715 $Y=0.74 $X2=0 $Y2=0
cc_278 N_A_119_368#_c_329_n X 0.0265088f $X=4.81 $Y=1.465 $X2=0 $Y2=0
cc_279 N_A_119_368#_c_340_n X 0.0416825f $X=4.835 $Y=2.395 $X2=0 $Y2=0
cc_280 N_A_119_368#_c_331_n X 0.056393f $X=5 $Y=1.465 $X2=0 $Y2=0
cc_281 N_A_119_368#_M1002_d N_A_38_74#_c_561_n 0.00655559f $X=0.625 $Y=0.37
+ $X2=0 $Y2=0
cc_282 N_A_119_368#_c_346_n N_A_38_74#_c_561_n 0.0425349f $X=1.365 $Y=0.845
+ $X2=0 $Y2=0
cc_283 N_A_119_368#_c_346_n A_270_74# 0.00156414f $X=1.365 $Y=0.845 $X2=-0.19
+ $Y2=-0.245
cc_284 N_A_119_368#_M1003_g N_VGND_c_594_n 0.00905011f $X=4.285 $Y=0.74 $X2=0
+ $Y2=0
cc_285 N_A_119_368#_M1013_g N_VGND_c_594_n 0.00108248f $X=4.715 $Y=0.74 $X2=0
+ $Y2=0
cc_286 N_A_119_368#_M1013_g N_VGND_c_596_n 0.0185296f $X=4.715 $Y=0.74 $X2=0
+ $Y2=0
cc_287 N_A_119_368#_c_331_n N_VGND_c_596_n 0.0292427f $X=5 $Y=1.465 $X2=0 $Y2=0
cc_288 N_A_119_368#_c_332_n N_VGND_c_596_n 0.00259603f $X=5 $Y=1.465 $X2=0 $Y2=0
cc_289 N_A_119_368#_c_330_n N_VGND_c_597_n 0.00498752f $X=1.45 $Y=1.82 $X2=0
+ $Y2=0
cc_290 N_A_119_368#_M1003_g N_VGND_c_601_n 0.00398535f $X=4.285 $Y=0.74 $X2=0
+ $Y2=0
cc_291 N_A_119_368#_M1013_g N_VGND_c_601_n 0.00461464f $X=4.715 $Y=0.74 $X2=0
+ $Y2=0
cc_292 N_A_119_368#_M1003_g N_VGND_c_603_n 0.00383639f $X=4.285 $Y=0.74 $X2=0
+ $Y2=0
cc_293 N_A_119_368#_M1013_g N_VGND_c_603_n 0.00837987f $X=4.715 $Y=0.74 $X2=0
+ $Y2=0
cc_294 N_A_27_368#_M1007_s N_A_209_368#_c_461_n 0.00540141f $X=1.595 $Y=1.96
+ $X2=0 $Y2=0
cc_295 N_A_27_368#_c_432_n N_A_209_368#_c_461_n 0.00784501f $X=1.575 $Y=2.99
+ $X2=0 $Y2=0
cc_296 N_A_27_368#_c_434_n N_A_209_368#_c_461_n 0.020636f $X=1.74 $Y=2.815 $X2=0
+ $Y2=0
cc_297 N_A_27_368#_c_431_n N_A_209_368#_c_462_n 2.76983e-19 $X=0.28 $Y=1.99
+ $X2=0 $Y2=0
cc_298 N_A_27_368#_c_432_n N_A_209_368#_c_462_n 0.0222695f $X=1.575 $Y=2.99
+ $X2=0 $Y2=0
cc_299 N_A_27_368#_c_434_n N_A_209_368#_c_462_n 0.00573056f $X=1.74 $Y=2.815
+ $X2=0 $Y2=0
cc_300 N_A_27_368#_c_434_n N_VPWR_c_491_n 0.0206899f $X=1.74 $Y=2.815 $X2=0
+ $Y2=0
cc_301 N_A_27_368#_c_432_n N_VPWR_c_495_n 0.0727635f $X=1.575 $Y=2.99 $X2=0
+ $Y2=0
cc_302 N_A_27_368#_c_433_n N_VPWR_c_495_n 0.0236566f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_303 N_A_27_368#_c_434_n N_VPWR_c_495_n 0.0226073f $X=1.74 $Y=2.815 $X2=0
+ $Y2=0
cc_304 N_A_27_368#_c_432_n N_VPWR_c_490_n 0.0424815f $X=1.575 $Y=2.99 $X2=0
+ $Y2=0
cc_305 N_A_27_368#_c_433_n N_VPWR_c_490_n 0.0128296f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_306 N_A_27_368#_c_434_n N_VPWR_c_490_n 0.012468f $X=1.74 $Y=2.815 $X2=0 $Y2=0
cc_307 N_A_209_368#_c_461_n N_VPWR_M1007_d 0.00545544f $X=2.575 $Y=2.395
+ $X2=-0.19 $Y2=1.66
cc_308 N_A_209_368#_c_461_n N_VPWR_c_491_n 0.0203886f $X=2.575 $Y=2.395 $X2=0
+ $Y2=0
cc_309 N_A_209_368#_c_463_n N_VPWR_c_491_n 0.0126571f $X=2.74 $Y=2.475 $X2=0
+ $Y2=0
cc_310 N_A_209_368#_c_463_n N_VPWR_c_496_n 0.0109675f $X=2.74 $Y=2.475 $X2=0
+ $Y2=0
cc_311 N_A_209_368#_c_461_n N_VPWR_c_490_n 0.0118427f $X=2.575 $Y=2.395 $X2=0
+ $Y2=0
cc_312 N_A_209_368#_c_463_n N_VPWR_c_490_n 0.00901496f $X=2.74 $Y=2.475 $X2=0
+ $Y2=0
cc_313 N_VPWR_M1008_d X 0.00476832f $X=3.815 $Y=1.84 $X2=0 $Y2=0
cc_314 X N_VGND_M1012_d 0.00605429f $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_315 X N_VGND_c_594_n 0.0178564f $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_316 X N_VGND_c_596_n 0.0159437f $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_317 X N_VGND_c_603_n 0.0180187f $X=3.995 $Y=0.84 $X2=0 $Y2=0
cc_318 N_A_38_74#_c_561_n A_270_74# 0.00149916f $X=2.42 $Y=0.375 $X2=-0.19
+ $Y2=-0.245
cc_319 N_A_38_74#_c_561_n N_VGND_M1009_d 0.0073435f $X=2.42 $Y=0.375 $X2=-0.19
+ $Y2=-0.245
cc_320 N_A_38_74#_M1004_d N_VGND_c_592_n 0.0058155f $X=2.445 $Y=0.37 $X2=0 $Y2=0
cc_321 N_A_38_74#_c_561_n N_VGND_c_592_n 0.0120082f $X=2.42 $Y=0.375 $X2=0 $Y2=0
cc_322 N_A_38_74#_c_563_n N_VGND_c_592_n 0.0200984f $X=2.585 $Y=0.375 $X2=0
+ $Y2=0
cc_323 N_A_38_74#_c_563_n N_VGND_c_593_n 0.0199996f $X=2.585 $Y=0.375 $X2=0
+ $Y2=0
cc_324 N_A_38_74#_c_561_n N_VGND_c_597_n 0.0110999f $X=2.42 $Y=0.375 $X2=0 $Y2=0
cc_325 N_A_38_74#_c_561_n N_VGND_c_598_n 0.0999537f $X=2.42 $Y=0.375 $X2=0 $Y2=0
cc_326 N_A_38_74#_c_562_n N_VGND_c_598_n 0.0193579f $X=0.5 $Y=0.375 $X2=0 $Y2=0
cc_327 N_A_38_74#_c_563_n N_VGND_c_598_n 0.0181829f $X=2.585 $Y=0.375 $X2=0
+ $Y2=0
cc_328 N_A_38_74#_c_561_n N_VGND_c_603_n 0.0680944f $X=2.42 $Y=0.375 $X2=0 $Y2=0
cc_329 N_A_38_74#_c_562_n N_VGND_c_603_n 0.0125128f $X=0.5 $Y=0.375 $X2=0 $Y2=0
cc_330 N_A_38_74#_c_563_n N_VGND_c_603_n 0.0121696f $X=2.585 $Y=0.375 $X2=0
+ $Y2=0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
M1000 a_230_94# A3 VGND VNB nlowvt w=640000u l=150000u
+  ad=4.48e+11p pd=3.96e+06u as=6.755e+11p ps=4.76e+06u
M1001 a_84_48# B1 a_230_94# VNB nlowvt w=640000u l=150000u
+  ad=2.272e+11p pd=1.99e+06u as=0p ps=0u
M1002 a_84_48# A3 a_343_368# VPB pshort w=1e+06u l=180000u
+  ad=3.472e+11p pd=2.72e+06u as=3.3e+11p ps=2.66e+06u
M1003 VGND A2 a_230_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_259_368# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=9.36e+11p ps=5.86e+06u
M1005 VPWR B1 a_84_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR a_84_48# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1007 a_230_94# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_84_48# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1009 a_343_368# A2 a_259_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_ms__nand2b_2.spice
* Created: Wed Sep  2 12:13:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nand2b_2.pex.spice"
.subckt sky130_fd_sc_ms__nand2b_2  VNB VPB A_N B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_N_M1008_g N_A_27_74#_M1008_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.16675 AS=0.1824 PD=1.81 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1006 N_Y_M1006_d N_A_27_74#_M1006_g N_A_242_74#_M1006_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.20635 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1009 N_Y_M1006_d N_A_27_74#_M1009_g N_A_242_74#_M1009_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_B_M1002_g N_A_242_74#_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10545 AS=0.1036 PD=1.025 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1002_d N_B_M1007_g N_A_242_74#_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10545 AS=0.2109 PD=1.025 PS=2.05 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_VPWR_M1003_d N_A_N_M1003_g N_A_27_74#_M1003_s VPB PSHORT L=0.18 W=1
+ AD=0.420189 AS=0.28 PD=1.83019 PS=2.56 NRD=39.3803 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1000 N_Y_M1000_d N_A_27_74#_M1000_g N_VPWR_M1003_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.470611 PD=1.39 PS=2.04981 NRD=0 NRS=60.2426 M=1 R=6.22222
+ SA=90001.1 SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1001 N_Y_M1000_d N_A_27_74#_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.6
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1004_d N_B_M1004_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002 SB=90000.6
+ A=0.2016 P=2.6 MULT=1
MM1005 N_Y_M1004_d N_B_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.5 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
c_68 VPB 0 1.91337e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__nand2b_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__dlrbp_1.spice
* Created: Fri Aug 28 17:27:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dlrbp_1.pex.spice"
.subckt sky130_fd_sc_ms__dlrbp_1  VNB VPB D GATE RESET_B VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_D_M1002_g N_A_27_142#_M1002_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.123281 AS=0.15675 PD=0.98062 PS=1.67 NRD=18 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1016 N_A_226_104#_M1016_d N_GATE_M1016_g N_VGND_M1002_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2701 AS=0.165869 PD=2.21 PS=1.31938 NRD=12.972 NRS=8.1 M=1
+ R=4.93333 SA=75000.6 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A_226_104#_M1003_g N_A_353_98#_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.207066 AS=0.259 PD=1.59797 PS=2.18 NRD=36.456 NRS=5.664 M=1
+ R=4.93333 SA=75000.3 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1007 A_571_80# N_A_27_142#_M1007_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0672 AS=0.179084 PD=0.85 PS=1.38203 NRD=9.372 NRS=15.936 M=1 R=4.26667
+ SA=75000.8 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1008 N_A_643_80#_M1008_d N_A_353_98#_M1008_g A_571_80# VNB NLOWVT L=0.15
+ W=0.64 AD=0.162536 AS=0.0672 PD=1.38868 PS=0.85 NRD=21.552 NRS=9.372 M=1
+ R=4.26667 SA=75001.1 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1015 A_775_124# N_A_226_104#_M1015_g N_A_643_80#_M1008_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.106664 PD=0.66 PS=0.911321 NRD=18.564 NRS=32.856 M=1
+ R=2.8 SA=75001.9 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_823_98#_M1006_g A_775_124# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1020 A_1051_74# N_A_643_80#_M1020_g N_A_823_98#_M1020_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_RESET_B_M1017_g A_1051_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1332 AS=0.0888 PD=1.1 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75000.6
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1000 N_Q_M1000_d N_A_823_98#_M1000_g N_VGND_M1017_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1332 PD=2.05 PS=1.1 NRD=0 NRS=12.972 M=1 R=4.93333 SA=75001.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A_823_98#_M1010_g N_A_1342_74#_M1010_s VNB NLOWVT L=0.15
+ W=0.55 AD=0.105886 AS=0.15675 PD=0.937984 PS=1.67 NRD=18 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1022 N_Q_N_M1022_d N_A_1342_74#_M1022_g N_VGND_M1010_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2738 AS=0.142464 PD=2.22 PS=1.26202 NRD=12.972 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1023 N_VPWR_M1023_d N_D_M1023_g N_A_27_142#_M1023_s VPB PSHORT L=0.18 W=0.84
+ AD=0.21525 AS=0.2352 PD=1.49 PS=2.24 NRD=47.1815 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90000.9 A=0.1512 P=2.04 MULT=1
MM1012 N_A_226_104#_M1012_d N_GATE_M1012_g N_VPWR_M1023_d VPB PSHORT L=0.18
+ W=0.84 AD=0.294 AS=0.21525 PD=2.38 PS=1.49 NRD=0 NRS=47.1815 M=1 R=4.66667
+ SA=90000.8 SB=90000.3 A=0.1512 P=2.04 MULT=1
MM1011 N_VPWR_M1011_d N_A_226_104#_M1011_g N_A_353_98#_M1011_s VPB PSHORT L=0.18
+ W=0.84 AD=0.15887 AS=0.2352 PD=1.24174 PS=2.24 NRD=19.9167 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90002.1 A=0.1512 P=2.04 MULT=1
MM1021 A_567_392# N_A_27_142#_M1021_g N_VPWR_M1011_d VPB PSHORT L=0.18 W=1
+ AD=0.105 AS=0.18913 PD=1.21 PS=1.47826 NRD=9.8303 NRS=0 M=1 R=5.55556
+ SA=90000.6 SB=90001.9 A=0.18 P=2.36 MULT=1
MM1001 N_A_643_80#_M1001_d N_A_226_104#_M1001_g A_567_392# VPB PSHORT L=0.18 W=1
+ AD=0.233451 AS=0.105 PD=1.93662 PS=1.21 NRD=0.9653 NRS=9.8303 M=1 R=5.55556
+ SA=90001 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1019 A_756_508# N_A_353_98#_M1019_g N_A_643_80#_M1001_d VPB PSHORT L=0.18
+ W=0.42 AD=0.09975 AS=0.0980493 PD=0.895 PS=0.81338 NRD=85.5965 NRS=44.5417 M=1
+ R=2.33333 SA=90001.5 SB=90002.6 A=0.0756 P=1.2 MULT=1
MM1005 N_VPWR_M1005_d N_A_823_98#_M1005_g A_756_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.121036 AS=0.09975 PD=0.96 PS=0.895 NRD=0 NRS=85.5965 M=1 R=2.33333
+ SA=90002.1 SB=90002 A=0.0756 P=1.2 MULT=1
MM1009 N_A_823_98#_M1009_d N_A_643_80#_M1009_g N_VPWR_M1005_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1652 AS=0.322764 PD=1.415 PS=2.56 NRD=3.5066 NRS=3.5066 M=1
+ R=6.22222 SA=90001.2 SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1013 N_VPWR_M1013_d N_RESET_B_M1013_g N_A_823_98#_M1009_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1792 AS=0.1652 PD=1.44 PS=1.415 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.7 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1014 N_Q_M1014_d N_A_823_98#_M1014_g N_VPWR_M1013_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1792 PD=2.8 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1004 N_VPWR_M1004_d N_A_823_98#_M1004_g N_A_1342_74#_M1004_s VPB PSHORT L=0.18
+ W=0.84 AD=0.147 AS=0.2352 PD=1.23857 PS=2.24 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1018 N_Q_N_M1018_d N_A_1342_74#_M1018_g N_VPWR_M1004_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.196 PD=2.8 PS=1.65143 NRD=0 NRS=8.7862 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX24_noxref VNB VPB NWDIODE A=15.8844 P=20.8
c_90 VNB 0 6.46507e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__dlrbp_1.pxi.spice"
*
.ends
*
*

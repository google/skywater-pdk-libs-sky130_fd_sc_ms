* File: sky130_fd_sc_ms__o2111ai_2.pex.spice
* Created: Fri Aug 28 17:52:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O2111AI_2%D1 3 5 7 10 12 14 15 19 21
c48 12 0 2.41312e-19 $X=0.99 $Y=1.22
r49 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r50 21 25 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.385
r51 18 19 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=0.99 $Y=1.385
+ $X2=0.995 $Y2=1.385
r52 17 18 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.56 $Y=1.385
+ $X2=0.99 $Y2=1.385
r53 16 17 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.545 $Y=1.385
+ $X2=0.56 $Y2=1.385
r54 15 24 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=0.455 $Y=1.385
+ $X2=0.27 $Y2=1.385
r55 15 16 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.455 $Y=1.385
+ $X2=0.545 $Y2=1.385
r56 12 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=1.22
+ $X2=0.99 $Y2=1.385
r57 12 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.99 $Y=1.22 $X2=0.99
+ $Y2=0.74
r58 8 19 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.55
+ $X2=0.995 $Y2=1.385
r59 8 10 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.995 $Y=1.55
+ $X2=0.995 $Y2=2.4
r60 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.56 $Y=1.22
+ $X2=0.56 $Y2=1.385
r61 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.56 $Y=1.22 $X2=0.56
+ $Y2=0.74
r62 1 16 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.55
+ $X2=0.545 $Y2=1.385
r63 1 3 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.545 $Y=1.55
+ $X2=0.545 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_2%C1 3 7 11 15 17 26
c61 26 0 4.60698e-20 $X=1.945 $Y=1.465
c62 15 0 2.35345e-20 $X=1.945 $Y=2.4
c63 3 0 8.60869e-20 $X=1.42 $Y=0.74
r64 25 26 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.92 $Y=1.465
+ $X2=1.945 $Y2=1.465
r65 23 25 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=1.85 $Y=1.465 $X2=1.92
+ $Y2=1.465
r66 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.85
+ $Y=1.465 $X2=1.85 $Y2=1.465
r67 21 23 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.495 $Y=1.465
+ $X2=1.85 $Y2=1.465
r68 19 21 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.42 $Y=1.465
+ $X2=1.495 $Y2=1.465
r69 17 24 3.75725 $w=5.52e-07 $l=1.7e-07 $layer=LI1_cond $X=1.68 $Y=1.295
+ $X2=1.68 $Y2=1.465
r70 13 26 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.945 $Y=1.63
+ $X2=1.945 $Y2=1.465
r71 13 15 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.945 $Y=1.63
+ $X2=1.945 $Y2=2.4
r72 9 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.92 $Y=1.3 $X2=1.92
+ $Y2=1.465
r73 9 11 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.92 $Y=1.3 $X2=1.92
+ $Y2=0.74
r74 5 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.495 $Y=1.63
+ $X2=1.495 $Y2=1.465
r75 5 7 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.495 $Y=1.63
+ $X2=1.495 $Y2=2.4
r76 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=1.3 $X2=1.42
+ $Y2=1.465
r77 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.42 $Y=1.3 $X2=1.42
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_2%B1 3 5 6 9 13 17 20 21 22 23 24
r63 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.29
+ $Y=1.515 $X2=3.29 $Y2=1.515
r64 24 30 8.30831 $w=4.28e-07 $l=3.1e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.29 $Y2=1.565
r65 23 30 4.55617 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.29 $Y2=1.565
r66 22 23 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.12 $Y2=1.565
r67 21 29 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=3.335 $Y=1.515
+ $X2=3.29 $Y2=1.515
r68 19 29 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=2.985 $Y=1.515
+ $X2=3.29 $Y2=1.515
r69 19 20 7.86782 $w=3.3e-07 $l=2.37382e-07 $layer=POLY_cond $X=2.985 $Y=1.515
+ $X2=2.755 $Y2=1.53
r70 15 21 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.41 $Y=1.35
+ $X2=3.335 $Y2=1.515
r71 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.41 $Y=1.35
+ $X2=3.41 $Y2=0.74
r72 11 20 16.8416 $w=1.5e-07 $l=2.45561e-07 $layer=POLY_cond $X=2.91 $Y=1.35
+ $X2=2.755 $Y2=1.53
r73 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.91 $Y=1.35
+ $X2=2.91 $Y2=0.74
r74 7 20 16.8416 $w=1.8e-07 $l=1.89737e-07 $layer=POLY_cond $X=2.845 $Y=1.68
+ $X2=2.755 $Y2=1.53
r75 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.845 $Y=1.68
+ $X2=2.845 $Y2=2.4
r76 5 20 7.86782 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.755 $Y=1.605
+ $X2=2.755 $Y2=1.53
r77 5 6 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.755 $Y=1.605
+ $X2=2.485 $Y2=1.605
r78 1 6 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.395 $Y=1.68
+ $X2=2.485 $Y2=1.605
r79 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.395 $Y=1.68
+ $X2=2.395 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_2%A2 3 7 11 15 17 18 28
c48 28 0 1.8469e-19 $X=4.305 $Y=1.515
c49 18 0 7.17692e-20 $X=4.56 $Y=1.665
c50 15 0 1.88192e-19 $X=4.305 $Y=2.4
r51 27 28 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.29 $Y=1.515
+ $X2=4.305 $Y2=1.515
r52 25 27 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=4.13 $Y=1.515
+ $X2=4.29 $Y2=1.515
r53 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.13
+ $Y=1.515 $X2=4.13 $Y2=1.515
r54 23 25 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=3.855 $Y=1.515
+ $X2=4.13 $Y2=1.515
r55 21 23 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.84 $Y=1.515
+ $X2=3.855 $Y2=1.515
r56 18 26 11.5244 $w=4.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.13 $Y2=1.565
r57 17 26 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=4.08 $Y=1.565 $X2=4.13
+ $Y2=1.565
r58 13 28 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.305 $Y=1.68
+ $X2=4.305 $Y2=1.515
r59 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.305 $Y=1.68
+ $X2=4.305 $Y2=2.4
r60 9 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.29 $Y=1.35
+ $X2=4.29 $Y2=1.515
r61 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.29 $Y=1.35 $X2=4.29
+ $Y2=0.74
r62 5 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.855 $Y=1.68
+ $X2=3.855 $Y2=1.515
r63 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.855 $Y=1.68
+ $X2=3.855 $Y2=2.4
r64 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.84 $Y=1.35
+ $X2=3.84 $Y2=1.515
r65 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.84 $Y=1.35 $X2=3.84
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_2%A1 3 7 11 15 17 18 25
c45 18 0 1.8469e-19 $X=5.52 $Y=1.665
c46 15 0 7.17692e-20 $X=5.255 $Y=2.4
r47 25 27 0.760252 $w=3.17e-07 $l=5e-09 $layer=POLY_cond $X=5.25 $Y=1.515
+ $X2=5.255 $Y2=1.515
r48 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.25
+ $Y=1.515 $X2=5.25 $Y2=1.515
r49 23 25 4.56151 $w=3.17e-07 $l=3e-08 $layer=POLY_cond $X=5.22 $Y=1.515
+ $X2=5.25 $Y2=1.515
r50 18 26 7.23627 $w=4.28e-07 $l=2.7e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.25 $Y2=1.565
r51 17 26 5.62821 $w=4.28e-07 $l=2.1e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.25 $Y2=1.565
r52 13 27 15.9969 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.255 $Y=1.68
+ $X2=5.255 $Y2=1.515
r53 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.255 $Y=1.68
+ $X2=5.255 $Y2=2.4
r54 9 23 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.22 $Y=1.35 $X2=5.22
+ $Y2=1.515
r55 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.22 $Y=1.35 $X2=5.22
+ $Y2=0.74
r56 5 23 70.7035 $w=3.17e-07 $l=4.65e-07 $layer=POLY_cond $X=4.755 $Y=1.515
+ $X2=5.22 $Y2=1.515
r57 5 21 5.32177 $w=3.17e-07 $l=3.5e-08 $layer=POLY_cond $X=4.755 $Y=1.515
+ $X2=4.72 $Y2=1.515
r58 5 7 285.702 $w=1.8e-07 $l=7.35e-07 $layer=POLY_cond $X=4.755 $Y=1.665
+ $X2=4.755 $Y2=2.4
r59 1 21 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.72 $Y=1.35 $X2=4.72
+ $Y2=1.515
r60 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.72 $Y=1.35 $X2=4.72
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_2%VPWR 1 2 3 4 5 16 18 24 26 30 34 38 40 42
+ 47 52 62 63 69 72 75 78
c79 38 0 1.88192e-19 $X=4.98 $Y=2.455
r80 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r81 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r82 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r83 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r84 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r85 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r86 63 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r87 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r88 60 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.145 $Y=3.33
+ $X2=4.98 $Y2=3.33
r89 60 62 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.145 $Y=3.33
+ $X2=5.52 $Y2=3.33
r90 59 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r91 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r92 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r93 56 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r94 55 58 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r95 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r96 53 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.235 $Y=3.33
+ $X2=3.11 $Y2=3.33
r97 53 55 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.235 $Y=3.33
+ $X2=3.6 $Y2=3.33
r98 52 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.815 $Y=3.33
+ $X2=4.98 $Y2=3.33
r99 52 58 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.815 $Y=3.33
+ $X2=4.56 $Y2=3.33
r100 51 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r101 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r102 48 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.255 $Y=3.33
+ $X2=2.17 $Y2=3.33
r103 48 50 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.255 $Y=3.33
+ $X2=2.64 $Y2=3.33
r104 47 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.985 $Y=3.33
+ $X2=3.11 $Y2=3.33
r105 47 50 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.985 $Y=3.33
+ $X2=2.64 $Y2=3.33
r106 46 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r107 46 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r108 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r109 43 66 3.96192 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=3.33
+ $X2=0.202 $Y2=3.33
r110 43 45 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.405 $Y=3.33
+ $X2=0.72 $Y2=3.33
r111 42 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.105 $Y=3.33
+ $X2=1.23 $Y2=3.33
r112 42 45 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.105 $Y=3.33
+ $X2=0.72 $Y2=3.33
r113 40 76 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r114 40 51 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r115 36 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=3.245
+ $X2=4.98 $Y2=3.33
r116 36 38 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=4.98 $Y=3.245
+ $X2=4.98 $Y2=2.455
r117 32 75 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.11 $Y=3.245
+ $X2=3.11 $Y2=3.33
r118 32 34 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=3.11 $Y=3.245
+ $X2=3.11 $Y2=2.455
r119 28 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=3.33
r120 28 30 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=2.455
r121 27 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.355 $Y=3.33
+ $X2=1.23 $Y2=3.33
r122 26 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=2.17 $Y2=3.33
r123 26 27 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=1.355 $Y2=3.33
r124 22 69 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=3.33
r125 22 24 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=2.305
r126 18 21 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r127 16 66 3.18124 $w=2.5e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.202 $Y2=3.33
r128 16 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r129 5 38 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=4.845
+ $Y=1.84 $X2=4.98 $Y2=2.455
r130 4 34 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.84 $X2=3.07 $Y2=2.455
r131 3 30 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=2.035
+ $Y=1.84 $X2=2.17 $Y2=2.455
r132 2 24 300 $w=1.7e-07 $l=5.49773e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=1.84 $X2=1.27 $Y2=2.305
r133 1 21 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.84 $X2=0.32 $Y2=2.815
r134 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.84 $X2=0.32 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_2%Y 1 2 3 4 5 18 20 24 26 30 32 36 42 44 45
+ 46 47 48 49 57 65 75
c83 57 0 4.60698e-20 $X=0.77 $Y=1.345
c84 20 0 2.35345e-20 $X=1.555 $Y=1.885
r85 62 65 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.77 $Y=1.97
+ $X2=0.77 $Y2=1.985
r86 57 75 2.07824 $w=3.3e-07 $l=5.09902e-08 $layer=LI1_cond $X=0.77 $Y=1.345
+ $X2=0.772 $Y2=1.295
r87 48 49 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.77 $Y=2.405
+ $X2=0.77 $Y2=2.775
r88 47 58 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=1.885
+ $X2=0.77 $Y2=1.8
r89 47 62 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=1.885
+ $X2=0.77 $Y2=1.97
r90 47 48 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.77 $Y=2.045
+ $X2=0.77 $Y2=2.405
r91 47 65 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=0.77 $Y=2.045 $X2=0.77
+ $Y2=1.985
r92 46 58 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.77 $Y=1.665
+ $X2=0.77 $Y2=1.8
r93 45 75 0.7625 $w=2.88e-07 $l=1.8e-08 $layer=LI1_cond $X=0.772 $Y=1.277
+ $X2=0.772 $Y2=1.295
r94 45 46 10.5815 $w=3.28e-07 $l=3.03e-07 $layer=LI1_cond $X=0.77 $Y=1.362
+ $X2=0.77 $Y2=1.665
r95 45 57 0.593683 $w=3.28e-07 $l=1.7e-08 $layer=LI1_cond $X=0.77 $Y=1.362
+ $X2=0.77 $Y2=1.345
r96 39 40 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=1.72 $Y=1.985 $X2=1.72
+ $Y2=2.035
r97 36 39 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.72 $Y=1.885 $X2=1.72
+ $Y2=1.985
r98 33 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.785 $Y=2.035
+ $X2=2.62 $Y2=2.035
r99 32 44 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.915 $Y=2.035
+ $X2=4.08 $Y2=2.035
r100 32 33 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=3.915 $Y=2.035
+ $X2=2.785 $Y2=2.035
r101 28 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=2.12
+ $X2=2.62 $Y2=2.035
r102 28 30 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.62 $Y=2.12
+ $X2=2.62 $Y2=2.815
r103 27 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.885 $Y=2.035
+ $X2=1.72 $Y2=2.035
r104 26 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.455 $Y=2.035
+ $X2=2.62 $Y2=2.035
r105 26 27 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.455 $Y=2.035
+ $X2=1.885 $Y2=2.035
r106 22 40 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=2.12
+ $X2=1.72 $Y2=2.035
r107 22 24 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.72 $Y=2.12
+ $X2=1.72 $Y2=2.815
r108 21 47 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=1.885
+ $X2=0.77 $Y2=1.885
r109 20 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=1.885
+ $X2=1.72 $Y2=1.885
r110 20 21 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.555 $Y=1.885
+ $X2=0.935 $Y2=1.885
r111 16 45 11.7675 $w=2.88e-07 $l=2.92711e-07 $layer=LI1_cond $X=0.815 $Y=1.005
+ $X2=0.772 $Y2=1.277
r112 16 18 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=0.815 $Y=1.005
+ $X2=0.815 $Y2=0.86
r113 5 44 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=3.945
+ $Y=1.84 $X2=4.08 $Y2=2.115
r114 4 42 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.485
+ $Y=1.84 $X2=2.62 $Y2=2.115
r115 4 30 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.485
+ $Y=1.84 $X2=2.62 $Y2=2.815
r116 3 39 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.585
+ $Y=1.84 $X2=1.72 $Y2=1.985
r117 3 24 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.585
+ $Y=1.84 $X2=1.72 $Y2=2.815
r118 2 49 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.635
+ $Y=1.84 $X2=0.77 $Y2=2.815
r119 2 65 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.635
+ $Y=1.84 $X2=0.77 $Y2=1.985
r120 1 18 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=0.635
+ $Y=0.37 $X2=0.775 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_2%A_697_368# 1 2 3 12 14 15 16 20 22 24
r35 22 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=2.12 $X2=5.48
+ $Y2=2.035
r36 22 24 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.48 $Y=2.12
+ $X2=5.48 $Y2=2.815
r37 21 27 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.615 $Y=2.035
+ $X2=4.53 $Y2=2.035
r38 20 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.315 $Y=2.035
+ $X2=5.48 $Y2=2.035
r39 20 21 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.315 $Y=2.035
+ $X2=4.615 $Y2=2.035
r40 17 19 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.53 $Y=2.905 $X2=4.53
+ $Y2=2.815
r41 16 27 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.53 $Y=2.12 $X2=4.53
+ $Y2=2.035
r42 16 19 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.53 $Y=2.12
+ $X2=4.53 $Y2=2.815
r43 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.445 $Y=2.99
+ $X2=4.53 $Y2=2.905
r44 14 15 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.445 $Y=2.99
+ $X2=3.715 $Y2=2.99
r45 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.59 $Y=2.905
+ $X2=3.715 $Y2=2.99
r46 10 12 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=3.59 $Y=2.905
+ $X2=3.59 $Y2=2.455
r47 3 29 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=5.345
+ $Y=1.84 $X2=5.48 $Y2=2.115
r48 3 24 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.345
+ $Y=1.84 $X2=5.48 $Y2=2.815
r49 2 27 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.84 $X2=4.53 $Y2=2.115
r50 2 19 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.84 $X2=4.53 $Y2=2.815
r51 1 12 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=3.485
+ $Y=1.84 $X2=3.63 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_2%A_40_74# 1 2 3 12 14 15 17 25 26
c40 17 0 1.39672e-19 $X=1.205 $Y=0.84
r41 25 26 9.7361 $w=5.33e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=0.862
+ $X2=1.97 $Y2=0.862
r42 21 23 3.40825 $w=1.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=1.29 $Y=0.925
+ $X2=1.205 $Y2=0.985
r43 21 26 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.29 $Y=0.925
+ $X2=1.97 $Y2=0.925
r44 17 23 3.40825 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.205 $Y=0.84
+ $X2=1.205 $Y2=0.985
r45 17 19 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.205 $Y=0.84
+ $X2=1.205 $Y2=0.515
r46 16 19 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.205 $Y=0.425
+ $X2=1.205 $Y2=0.515
r47 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.12 $Y=0.34
+ $X2=1.205 $Y2=0.425
r48 14 15 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.12 $Y=0.34
+ $X2=0.51 $Y2=0.34
r49 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.345 $Y=0.425
+ $X2=0.51 $Y2=0.34
r50 10 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.345 $Y=0.425
+ $X2=0.345 $Y2=0.515
r51 3 25 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=1.995
+ $Y=0.37 $X2=2.135 $Y2=0.86
r52 2 23 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.37 $X2=1.205 $Y2=0.965
r53 2 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.37 $X2=1.205 $Y2=0.515
r54 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.2
+ $Y=0.37 $X2=0.345 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_2%A_299_74# 1 2 7 11 13
c26 13 0 1.01641e-19 $X=1.635 $Y=0.34
c27 7 0 8.60869e-20 $X=3.03 $Y=0.34
r28 13 16 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.635 $Y=0.34
+ $X2=1.635 $Y2=0.55
r29 9 11 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=3.195 $Y=0.425
+ $X2=3.195 $Y2=0.635
r30 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.8 $Y=0.34 $X2=1.635
+ $Y2=0.34
r31 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.03 $Y=0.34
+ $X2=3.195 $Y2=0.425
r32 7 8 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=3.03 $Y=0.34 $X2=1.8
+ $Y2=0.34
r33 2 11 182 $w=1.7e-07 $l=3.54789e-07 $layer=licon1_NDIFF $count=1 $X=2.985
+ $Y=0.37 $X2=3.195 $Y2=0.635
r34 1 16 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.495 $Y=0.37
+ $X2=1.635 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_2%A_510_74# 1 2 3 4 15 17 18 21 23 27 29 33
+ 35 36
r63 31 33 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=5.475 $Y=1.01
+ $X2=5.475 $Y2=0.515
r64 30 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.67 $Y=1.095
+ $X2=4.545 $Y2=1.095
r65 29 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.35 $Y=1.095
+ $X2=5.475 $Y2=1.01
r66 29 30 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.35 $Y=1.095
+ $X2=4.67 $Y2=1.095
r67 25 36 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.545 $Y=1.01
+ $X2=4.545 $Y2=1.095
r68 25 27 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=4.545 $Y=1.01
+ $X2=4.545 $Y2=0.515
r69 24 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.71 $Y=1.095
+ $X2=3.625 $Y2=1.095
r70 23 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.42 $Y=1.095
+ $X2=4.545 $Y2=1.095
r71 23 24 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.42 $Y=1.095
+ $X2=3.71 $Y2=1.095
r72 19 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=1.01
+ $X2=3.625 $Y2=1.095
r73 19 21 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.625 $Y=1.01
+ $X2=3.625 $Y2=0.515
r74 17 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=1.095
+ $X2=3.625 $Y2=1.095
r75 17 18 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.54 $Y=1.095
+ $X2=2.86 $Y2=1.095
r76 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.695 $Y=1.01
+ $X2=2.86 $Y2=1.095
r77 13 15 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.695 $Y=1.01
+ $X2=2.695 $Y2=0.86
r78 4 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.295
+ $Y=0.37 $X2=5.435 $Y2=0.515
r79 3 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.365
+ $Y=0.37 $X2=4.505 $Y2=0.515
r80 2 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.485
+ $Y=0.37 $X2=3.625 $Y2=0.515
r81 1 15 182 $w=1.7e-07 $l=5.57808e-07 $layer=licon1_NDIFF $count=1 $X=2.55
+ $Y=0.37 $X2=2.695 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_2%VGND 1 2 9 13 15 17 25 32 33 36 39
r58 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r59 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r60 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r61 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r62 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.17 $Y=0 $X2=5.005
+ $Y2=0
r63 30 32 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5.17 $Y=0 $X2=5.52
+ $Y2=0
r64 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r65 29 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r66 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r67 26 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.22 $Y=0 $X2=4.055
+ $Y2=0
r68 26 28 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.22 $Y=0 $X2=4.56
+ $Y2=0
r69 25 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.84 $Y=0 $X2=5.005
+ $Y2=0
r70 25 28 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.84 $Y=0 $X2=4.56
+ $Y2=0
r71 24 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r72 23 24 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r73 19 23 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=3.6
+ $Y2=0
r74 19 20 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r75 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.89 $Y=0 $X2=4.055
+ $Y2=0
r76 17 23 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.89 $Y=0 $X2=3.6
+ $Y2=0
r77 15 24 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.6
+ $Y2=0
r78 15 20 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=0.24
+ $Y2=0
r79 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=0.085
+ $X2=5.005 $Y2=0
r80 11 13 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=5.005 $Y=0.085
+ $X2=5.005 $Y2=0.595
r81 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.055 $Y=0.085
+ $X2=4.055 $Y2=0
r82 7 9 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=4.055 $Y=0.085
+ $X2=4.055 $Y2=0.595
r83 2 13 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=4.795
+ $Y=0.37 $X2=5.005 $Y2=0.595
r84 1 9 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=3.915
+ $Y=0.37 $X2=4.055 $Y2=0.595
.ends


* File: sky130_fd_sc_ms__a222o_2.pex.spice
* Created: Wed Sep  2 11:52:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A222O_2%C1 3 5 8 10 11 15 18
c32 15 0 1.32914e-19 $X=0.27 $Y=1.465
r33 17 18 0.524584 $w=3.3e-07 $l=3e-09 $layer=POLY_cond $X=0.492 $Y=1.465
+ $X2=0.495 $Y2=1.465
r34 14 17 38.8192 $w=3.3e-07 $l=2.22e-07 $layer=POLY_cond $X=0.27 $Y=1.465
+ $X2=0.492 $Y2=1.465
r35 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r36 11 15 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.27 $Y=1.665 $X2=0.27
+ $Y2=1.465
r37 6 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.465
r38 6 8 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.73
r39 3 10 36.5274 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.92 $X2=0.505
+ $Y2=1.83
r40 3 5 144.6 $w=1.8e-07 $l=5.4e-07 $layer=POLY_cond $X=0.505 $Y=1.92 $X2=0.505
+ $Y2=2.46
r41 1 17 20.5173 $w=1.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.492 $Y=1.63
+ $X2=0.492 $Y2=1.465
r42 1 10 95.6824 $w=1.55e-07 $l=2e-07 $layer=POLY_cond $X=0.492 $Y=1.63
+ $X2=0.492 $Y2=1.83
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_2%C2 3 7 9 12 13
c35 7 0 1.32914e-19 $X=0.955 $Y=2.46
r36 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.425
+ $X2=0.975 $Y2=1.59
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.425
+ $X2=0.975 $Y2=1.26
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.425 $X2=0.975 $Y2=1.425
r39 9 13 5.86538 $w=5.18e-07 $l=2.55e-07 $layer=LI1_cond $X=0.72 $Y=1.52
+ $X2=0.975 $Y2=1.52
r40 7 15 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=0.955 $Y=2.46
+ $X2=0.955 $Y2=1.59
r41 3 14 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.885 $Y=0.73
+ $X2=0.885 $Y2=1.26
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_2%A_27_82# 1 2 3 4 13 15 16 17 20 22 24 27 31
+ 33 35 37 38 39 44 46 47 48 50 53 54 56 60 61 63
c131 56 0 1.07056e-19 $X=3.265 $Y=1.095
r132 57 61 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=1.095
+ $X2=2.395 $Y2=1.095
r133 56 63 5.67212 $w=4.83e-07 $l=2.3e-07 $layer=LI1_cond $X=3.507 $Y=1.095
+ $X2=3.507 $Y2=0.865
r134 56 57 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=3.265 $Y=1.095
+ $X2=2.56 $Y2=1.095
r135 54 70 14.8853 $w=3.4e-07 $l=1.05e-07 $layer=POLY_cond $X=2.395 $Y=1.47
+ $X2=2.5 $Y2=1.47
r136 54 68 45.3647 $w=3.4e-07 $l=3.2e-07 $layer=POLY_cond $X=2.395 $Y=1.47
+ $X2=2.075 $Y2=1.47
r137 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.395
+ $Y=1.425 $X2=2.395 $Y2=1.425
r138 51 61 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.395 $Y=1.18
+ $X2=2.395 $Y2=1.095
r139 51 53 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.395 $Y=1.18
+ $X2=2.395 $Y2=1.425
r140 50 61 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.315 $Y=1.01
+ $X2=2.395 $Y2=1.095
r141 49 50 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.315 $Y=0.75
+ $X2=2.315 $Y2=1.01
r142 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.23 $Y=0.665
+ $X2=2.315 $Y2=0.75
r143 47 48 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.23 $Y=0.665
+ $X2=1.525 $Y2=0.665
r144 45 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.44 $Y=1.09
+ $X2=1.44 $Y2=1.005
r145 45 46 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=1.44 $Y=1.09
+ $X2=1.44 $Y2=1.95
r146 44 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.44 $Y=0.92
+ $X2=1.44 $Y2=1.005
r147 43 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.44 $Y=0.75
+ $X2=1.525 $Y2=0.665
r148 43 44 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.44 $Y=0.75
+ $X2=1.44 $Y2=0.92
r149 40 59 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=2.075
+ $X2=0.24 $Y2=2.075
r150 40 42 37.5696 $w=2.48e-07 $l=8.15e-07 $layer=LI1_cond $X=0.365 $Y=2.075
+ $X2=1.18 $Y2=2.075
r151 39 46 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.355 $Y=2.075
+ $X2=1.44 $Y2=1.95
r152 39 42 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=1.355 $Y=2.075
+ $X2=1.18 $Y2=2.075
r153 37 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.355 $Y=1.005
+ $X2=1.44 $Y2=1.005
r154 37 38 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=1.355 $Y=1.005
+ $X2=0.365 $Y2=1.005
r155 33 59 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=2.2
+ $X2=0.24 $Y2=2.075
r156 33 35 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=0.24 $Y=2.2
+ $X2=0.24 $Y2=2.465
r157 29 38 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=0.92
+ $X2=0.365 $Y2=1.005
r158 29 31 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=0.24 $Y=0.92
+ $X2=0.24 $Y2=0.555
r159 25 70 17.6285 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=2.5 $Y=1.68 $X2=2.5
+ $Y2=1.47
r160 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.5 $Y=1.68 $X2=2.5
+ $Y2=2.4
r161 22 68 21.9347 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.075 $Y=1.26
+ $X2=2.075 $Y2=1.47
r162 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.075 $Y=1.26
+ $X2=2.075 $Y2=0.78
r163 18 68 3.54412 $w=3.4e-07 $l=2.5e-08 $layer=POLY_cond $X=2.05 $Y=1.47
+ $X2=2.075 $Y2=1.47
r164 18 20 314.855 $w=1.8e-07 $l=8.1e-07 $layer=POLY_cond $X=2.05 $Y=1.59
+ $X2=2.05 $Y2=2.4
r165 16 18 28.0472 $w=3.4e-07 $l=1.74284e-07 $layer=POLY_cond $X=1.96 $Y=1.335
+ $X2=2.05 $Y2=1.47
r166 16 17 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.96 $Y=1.335
+ $X2=1.72 $Y2=1.335
r167 13 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.645 $Y=1.26
+ $X2=1.72 $Y2=1.335
r168 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.645 $Y=1.26
+ $X2=1.645 $Y2=0.78
r169 4 42 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.96 $X2=1.18 $Y2=2.115
r170 3 59 600 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.115
r171 3 35 300 $w=1.7e-07 $l=5.72931e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.465
r172 2 63 182 $w=1.7e-07 $l=6.07268e-07 $layer=licon1_NDIFF $count=1 $X=3.255
+ $Y=0.37 $X2=3.505 $Y2=0.865
r173 1 31 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.41 $X2=0.28 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_2%A1 3 7 9 10 14 15
r42 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=1.515
+ $X2=3.09 $Y2=1.68
r43 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.09 $Y=1.515
+ $X2=3.09 $Y2=1.35
r44 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.515 $X2=3.09 $Y2=1.515
r45 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.09 $Y=1.665
+ $X2=3.09 $Y2=2.035
r46 9 15 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.09 $Y=1.665
+ $X2=3.09 $Y2=1.515
r47 7 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.18 $Y=0.69 $X2=3.18
+ $Y2=1.35
r48 3 17 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.12 $Y=2.34 $X2=3.12
+ $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_2%B1 3 7 9 12 13
c36 13 0 8.45074e-20 $X=3.63 $Y=1.515
c37 7 0 1.07056e-19 $X=3.8 $Y=0.69
r38 12 15 40.172 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.515
+ $X2=3.67 $Y2=1.68
r39 12 14 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.515
+ $X2=3.67 $Y2=1.35
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.63
+ $Y=1.515 $X2=3.63 $Y2=1.515
r41 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.63 $Y=1.665
+ $X2=3.63 $Y2=1.515
r42 7 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.8 $Y=0.69 $X2=3.8
+ $Y2=1.35
r43 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.775 $Y=2.34
+ $X2=3.775 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_2%B2 3 7 9 12 13
c39 7 0 1.88727e-19 $X=4.225 $Y=2.34
r40 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.28 $Y=1.515
+ $X2=4.28 $Y2=1.68
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.28 $Y=1.515
+ $X2=4.28 $Y2=1.35
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.28
+ $Y=1.515 $X2=4.28 $Y2=1.515
r43 9 13 5.3602 $w=4.28e-07 $l=2e-07 $layer=LI1_cond $X=4.08 $Y=1.565 $X2=4.28
+ $Y2=1.565
r44 7 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=4.225 $Y=2.34
+ $X2=4.225 $Y2=1.68
r45 3 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.19 $Y=0.69 $X2=4.19
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_2%A2 3 7 9 12
c27 9 0 1.0422e-19 $X=5.04 $Y=1.665
r28 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.85 $Y=1.515
+ $X2=4.85 $Y2=1.68
r29 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.85 $Y=1.515
+ $X2=4.85 $Y2=1.35
r30 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.85
+ $Y=1.515 $X2=4.85 $Y2=1.515
r31 9 13 5.09219 $w=4.28e-07 $l=1.9e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=4.85 $Y2=1.565
r32 7 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=4.775 $Y=2.34
+ $X2=4.775 $Y2=1.68
r33 3 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.76 $Y=0.69 $X2=4.76
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_2%A_119_392# 1 2 9 13 16
r35 11 13 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=4 $Y=2.37 $X2=4
+ $Y2=2.115
r36 10 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=2.455
+ $X2=0.73 $Y2=2.455
r37 9 11 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.835 $Y=2.455
+ $X2=4 $Y2=2.37
r38 9 10 191.807 $w=1.68e-07 $l=2.94e-06 $layer=LI1_cond $X=3.835 $Y=2.455
+ $X2=0.895 $Y2=2.455
r39 2 13 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=3.865
+ $Y=1.84 $X2=4 $Y2=2.115
r40 1 16 300 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.96 $X2=0.73 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_2%VPWR 1 2 3 12 16 18 20 23 24 25 27 39 47 51
r51 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r52 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 45 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r54 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r55 42 45 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r56 41 44 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r57 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r58 39 50 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=4.835 $Y=3.33
+ $X2=5.057 $Y2=3.33
r59 39 44 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.835 $Y=3.33
+ $X2=4.56 $Y2=3.33
r60 35 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=1.74 $Y2=3.33
r61 35 37 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=2.64 $Y2=3.33
r62 34 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r64 30 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r65 29 33 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r66 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r67 27 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.74 $Y2=3.33
r68 27 33 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.2 $Y2=3.33
r69 25 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r70 25 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.68 $Y2=3.33
r71 25 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r72 23 37 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.645 $Y=3.33
+ $X2=2.64 $Y2=3.33
r73 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.645 $Y=3.33
+ $X2=2.81 $Y2=3.33
r74 22 41 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.975 $Y=3.33
+ $X2=3.12 $Y2=3.33
r75 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=3.33
+ $X2=2.81 $Y2=3.33
r76 18 50 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5 $Y=3.245
+ $X2=5.057 $Y2=3.33
r77 18 20 39.4624 $w=3.28e-07 $l=1.13e-06 $layer=LI1_cond $X=5 $Y=3.245 $X2=5
+ $Y2=2.115
r78 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=3.245
+ $X2=2.81 $Y2=3.33
r79 14 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.81 $Y=3.245
+ $X2=2.81 $Y2=2.875
r80 10 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=3.245
+ $X2=1.74 $Y2=3.33
r81 10 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.74 $Y=3.245
+ $X2=1.74 $Y2=2.875
r82 3 20 300 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=2 $X=4.865
+ $Y=1.84 $X2=5 $Y2=2.115
r83 2 16 600 $w=1.7e-07 $l=1.1397e-06 $layer=licon1_PDIFF $count=1 $X=2.59
+ $Y=1.84 $X2=2.81 $Y2=2.875
r84 1 12 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=2.73 $X2=1.74 $Y2=2.875
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_2%X 1 2 9 11 18
r28 11 18 3.48766 $w=3.78e-07 $l=1.15e-07 $layer=LI1_cond $X=2.16 $Y=2.01
+ $X2=2.275 $Y2=2.01
r29 11 13 9.09823 $w=3.78e-07 $l=3e-07 $layer=LI1_cond $X=2.16 $Y=2.01 $X2=1.86
+ $Y2=2.01
r30 7 13 1.56319 $w=3.3e-07 $l=1.9e-07 $layer=LI1_cond $X=1.86 $Y=1.82 $X2=1.86
+ $Y2=2.01
r31 7 9 28.4618 $w=3.28e-07 $l=8.15e-07 $layer=LI1_cond $X=1.86 $Y=1.82 $X2=1.86
+ $Y2=1.005
r32 2 18 600 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=2.14
+ $Y=1.84 $X2=2.275 $Y2=2.01
r33 1 9 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.72
+ $Y=0.41 $X2=1.86 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_2%A_642_368# 1 2 7 11 16
r22 16 18 3.63098 $w=3.63e-07 $l=1.15e-07 $layer=LI1_cond $X=3.447 $Y=2.875
+ $X2=3.447 $Y2=2.99
r23 11 14 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.5 $Y=2.035 $X2=4.5
+ $Y2=2.715
r24 9 14 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.5 $Y=2.905 $X2=4.5
+ $Y2=2.715
r25 8 18 5.2253 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=3.63 $Y=2.99 $X2=3.447
+ $Y2=2.99
r26 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.335 $Y=2.99
+ $X2=4.5 $Y2=2.905
r27 7 8 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=4.335 $Y=2.99
+ $X2=3.63 $Y2=2.99
r28 2 14 400 $w=1.7e-07 $l=9.63068e-07 $layer=licon1_PDIFF $count=1 $X=4.315
+ $Y=1.84 $X2=4.5 $Y2=2.715
r29 2 11 400 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_PDIFF $count=1 $X=4.315
+ $Y=1.84 $X2=4.5 $Y2=2.035
r30 1 16 600 $w=1.7e-07 $l=1.14649e-06 $layer=licon1_PDIFF $count=1 $X=3.21
+ $Y=1.84 $X2=3.445 $Y2=2.875
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_2%VGND 1 2 3 12 16 19 20 21 22 29 30 31 50 51
r63 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r64 48 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r65 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r66 44 47 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.08
+ $Y2=0
r67 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r68 39 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r69 38 41 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r70 38 39 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r71 35 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r72 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r73 31 48 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=4.08
+ $Y2=0
r74 31 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r75 31 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r76 29 47 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.26 $Y=0 $X2=4.08
+ $Y2=0
r77 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.26 $Y=0 $X2=4.425
+ $Y2=0
r78 28 50 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.59 $Y=0 $X2=5.04
+ $Y2=0
r79 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.59 $Y=0 $X2=4.425
+ $Y2=0
r80 24 44 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.535 $Y=0 $X2=2.64
+ $Y2=0
r81 22 41 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.16
+ $Y2=0
r82 21 26 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.37 $Y=0 $X2=2.37
+ $Y2=0.325
r83 21 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.37 $Y=0 $X2=2.535
+ $Y2=0
r84 21 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.37 $Y=0 $X2=2.205
+ $Y2=0
r85 19 34 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.72
+ $Y2=0
r86 19 20 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.06
+ $Y2=0
r87 18 38 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.2
+ $Y2=0
r88 18 20 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.06
+ $Y2=0
r89 14 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.425 $Y=0.085
+ $X2=4.425 $Y2=0
r90 14 16 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=4.425 $Y=0.085
+ $X2=4.425 $Y2=0.635
r91 10 20 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.06 $Y=0.085
+ $X2=1.06 $Y2=0
r92 10 12 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=1.06 $Y=0.085
+ $X2=1.06 $Y2=0.57
r93 3 16 182 $w=1.7e-07 $l=3.35596e-07 $layer=licon1_NDIFF $count=1 $X=4.265
+ $Y=0.37 $X2=4.425 $Y2=0.635
r94 2 26 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=2.15
+ $Y=0.41 $X2=2.37 $Y2=0.325
r95 1 12 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=0.96
+ $Y=0.41 $X2=1.1 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_MS__A222O_2%A_557_74# 1 2 7 10 11 12 15 17
c38 7 0 2.49076e-20 $X=3.92 $Y=0.435
r39 17 20 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.93 $Y=0.435 $X2=2.93
+ $Y2=0.635
r40 13 15 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.975 $Y=1.01
+ $X2=4.975 $Y2=0.515
r41 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.81 $Y=1.095
+ $X2=4.975 $Y2=1.01
r42 11 12 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=4.81 $Y=1.095
+ $X2=4.09 $Y2=1.095
r43 10 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.005 $Y=1.01
+ $X2=4.09 $Y2=1.095
r44 9 10 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=4.005 $Y=0.52
+ $X2=4.005 $Y2=1.01
r45 8 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.095 $Y=0.435
+ $X2=2.93 $Y2=0.435
r46 7 9 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.92 $Y=0.435
+ $X2=4.005 $Y2=0.52
r47 7 8 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=3.92 $Y=0.435
+ $X2=3.095 $Y2=0.435
r48 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.835
+ $Y=0.37 $X2=4.975 $Y2=0.515
r49 1 20 182 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_NDIFF $count=1 $X=2.785
+ $Y=0.37 $X2=2.93 $Y2=0.635
.ends


* File: sky130_fd_sc_ms__nand4bb_1.pex.spice
* Created: Fri Aug 28 17:45:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NAND4BB_1%A_N 1 3 8 10 14 16
r28 13 16 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.315 $Y=0.42
+ $X2=0.52 $Y2=0.42
r29 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.315
+ $Y=0.42 $X2=0.315 $Y2=0.42
r30 10 14 4.38253 $w=3.53e-07 $l=1.35e-07 $layer=LI1_cond $X=0.302 $Y=0.555
+ $X2=0.302 $Y2=0.42
r31 8 9 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=0.52 $Y=0.97 $X2=0.52
+ $Y2=1.375
r32 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=0.585
+ $X2=0.52 $Y2=0.42
r33 5 8 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.52 $Y=0.585
+ $X2=0.52 $Y2=0.97
r34 1 9 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.505 $Y=1.465 $X2=0.505
+ $Y2=1.375
r35 1 3 367.331 $w=1.8e-07 $l=9.45e-07 $layer=POLY_cond $X=0.505 $Y=1.465
+ $X2=0.505 $Y2=2.41
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4BB_1%B_N 3 7 9 10 14
c34 14 0 8.08011e-20 $X=1.01 $Y=1.635
r35 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.01 $Y=1.635
+ $X2=1.01 $Y2=1.8
r36 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.01 $Y=1.635
+ $X2=1.01 $Y2=1.47
r37 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.01
+ $Y=1.635 $X2=1.01 $Y2=1.635
r38 10 15 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=1.2 $Y=1.635
+ $X2=1.01 $Y2=1.635
r39 9 15 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=0.72 $Y=1.635
+ $X2=1.01 $Y2=1.635
r40 7 16 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.1 $Y=0.925 $X2=1.1
+ $Y2=1.47
r41 3 17 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=1.055 $Y=2.41
+ $X2=1.055 $Y2=1.8
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4BB_1%A_27_398# 1 2 9 11 13 18 20 26 27 28 37
c64 28 0 8.08011e-20 $X=1.85 $Y=1.215
c65 9 0 4.10042e-20 $X=2.065 $Y=2.4
r66 36 37 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=2.065 $Y=1.385
+ $X2=2.1 $Y2=1.385
r67 32 36 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.85 $Y=1.385
+ $X2=2.065 $Y2=1.385
r68 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.85
+ $Y=1.385 $X2=1.85 $Y2=1.385
r69 28 31 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.85 $Y=1.215
+ $X2=1.85 $Y2=1.385
r70 25 26 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.305 $Y=1.07
+ $X2=0.47 $Y2=1.07
r71 22 25 2.73018 $w=4.58e-07 $l=1.05e-07 $layer=LI1_cond $X=0.2 $Y=1.07
+ $X2=0.305 $Y2=1.07
r72 20 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.215
+ $X2=1.85 $Y2=1.215
r73 20 26 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=1.685 $Y=1.215
+ $X2=0.47 $Y2=1.215
r74 18 27 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=2.135
+ $X2=0.28 $Y2=1.97
r75 14 22 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.2 $Y=1.3 $X2=0.2
+ $Y2=1.07
r76 14 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.2 $Y=1.3 $X2=0.2
+ $Y2=1.97
r77 11 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.1 $Y=1.22 $X2=2.1
+ $Y2=1.385
r78 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.1 $Y=1.22 $X2=2.1
+ $Y2=0.74
r79 7 36 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.065 $Y=1.55
+ $X2=2.065 $Y2=1.385
r80 7 9 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.065 $Y=1.55
+ $X2=2.065 $Y2=2.4
r81 2 18 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.99 $X2=0.28 $Y2=2.135
r82 1 25 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.86 $X2=0.305 $Y2=1.05
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4BB_1%A_229_398# 1 2 9 12 16 18 21 23 25 29 33
+ 34 37
r77 34 38 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.58 $Y=1.385
+ $X2=2.58 $Y2=1.55
r78 34 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.58 $Y=1.385
+ $X2=2.58 $Y2=1.22
r79 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.58
+ $Y=1.385 $X2=2.58 $Y2=1.385
r80 30 33 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=2.27 $Y=1.385
+ $X2=2.58 $Y2=1.385
r81 27 29 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.32 $Y=0.795
+ $X2=1.49 $Y2=0.795
r82 22 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.27 $Y=1.55
+ $X2=2.27 $Y2=1.385
r83 22 23 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.27 $Y=1.55
+ $X2=2.27 $Y2=1.97
r84 21 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.27 $Y=1.22
+ $X2=2.27 $Y2=1.385
r85 20 21 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.27 $Y=0.96
+ $X2=2.27 $Y2=1.22
r86 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.185 $Y=0.875
+ $X2=2.27 $Y2=0.96
r87 18 29 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.185 $Y=0.875
+ $X2=1.49 $Y2=0.875
r88 17 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=2.055
+ $X2=1.28 $Y2=2.055
r89 16 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.185 $Y=2.055
+ $X2=2.27 $Y2=1.97
r90 16 17 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.185 $Y=2.055
+ $X2=1.445 $Y2=2.055
r91 12 38 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.655 $Y=2.4
+ $X2=2.655 $Y2=1.55
r92 9 37 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.49 $Y=0.74 $X2=2.49
+ $Y2=1.22
r93 2 25 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.145
+ $Y=1.99 $X2=1.28 $Y2=2.135
r94 1 27 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=1.175
+ $Y=0.65 $X2=1.32 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4BB_1%C 3 6 8 9 13 15
r45 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=1.385
+ $X2=3.15 $Y2=1.55
r46 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=1.385
+ $X2=3.15 $Y2=1.22
r47 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.15
+ $Y=1.385 $X2=3.15 $Y2=1.385
r48 9 14 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.15 $Y=1.295 $X2=3.15
+ $Y2=1.385
r49 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.15 $Y=0.925 $X2=3.15
+ $Y2=1.295
r50 6 16 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.155 $Y=2.4
+ $X2=3.155 $Y2=1.55
r51 3 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.06 $Y=0.74 $X2=3.06
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4BB_1%D 3 7 9 12 13
r40 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.72 $Y=1.515
+ $X2=3.72 $Y2=1.68
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.72 $Y=1.515
+ $X2=3.72 $Y2=1.35
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.72
+ $Y=1.515 $X2=3.72 $Y2=1.515
r43 9 13 4.32166 $w=3.98e-07 $l=1.5e-07 $layer=LI1_cond $X=3.685 $Y=1.665
+ $X2=3.685 $Y2=1.515
r44 7 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.705 $Y=2.4
+ $X2=3.705 $Y2=1.68
r45 3 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.63 $Y=0.74 $X2=3.63
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4BB_1%VPWR 1 2 3 12 16 20 23 24 26 27 28 30 46
+ 47 50
r58 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r60 44 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r61 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r62 38 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r63 37 40 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r64 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r65 35 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r66 35 37 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r67 33 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r68 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r69 30 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r70 30 32 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r71 28 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r72 28 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r73 28 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r74 26 43 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.265 $Y=3.33
+ $X2=3.12 $Y2=3.33
r75 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.265 $Y=3.33
+ $X2=3.43 $Y2=3.33
r76 25 46 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.595 $Y=3.33
+ $X2=4.08 $Y2=3.33
r77 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=3.33
+ $X2=3.43 $Y2=3.33
r78 23 40 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.175 $Y=3.33
+ $X2=2.16 $Y2=3.33
r79 23 24 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.175 $Y=3.33
+ $X2=2.385 $Y2=3.33
r80 22 43 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.595 $Y=3.33
+ $X2=3.12 $Y2=3.33
r81 22 24 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.595 $Y=3.33
+ $X2=2.385 $Y2=3.33
r82 18 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=3.245
+ $X2=3.43 $Y2=3.33
r83 18 20 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=3.43 $Y=3.245
+ $X2=3.43 $Y2=2.455
r84 14 24 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=3.245
+ $X2=2.385 $Y2=3.33
r85 14 16 11.7988 $w=4.18e-07 $l=4.3e-07 $layer=LI1_cond $X=2.385 $Y=3.245
+ $X2=2.385 $Y2=2.815
r86 10 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r87 10 12 38.764 $w=3.28e-07 $l=1.11e-06 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.135
r88 3 20 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=3.245
+ $Y=1.84 $X2=3.43 $Y2=2.455
r89 2 16 600 $w=1.7e-07 $l=1.08392e-06 $layer=licon1_PDIFF $count=1 $X=2.155
+ $Y=1.84 $X2=2.385 $Y2=2.815
r90 1 12 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.99 $X2=0.78 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4BB_1%Y 1 2 3 4 15 19 23 25 28 29 30 33 36 38 40
+ 41 44
c92 44 0 4.10042e-20 $X=2.93 $Y=1.985
r93 48 49 3.88629 $w=5.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=2.395
+ $X2=2.81 $Y2=2.48
r94 41 48 7.55418 $w=5.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.81 $Y=2.035
+ $X2=2.81 $Y2=2.395
r95 41 44 1.04919 $w=5.68e-07 $l=5e-08 $layer=LI1_cond $X=2.81 $Y=2.035 $X2=2.81
+ $Y2=1.985
r96 36 40 3.01263 $w=3.15e-07 $l=1.8262e-07 $layer=LI1_cond $X=4.14 $Y=1.95
+ $X2=3.995 $Y2=2.035
r97 35 36 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.14 $Y=1.18
+ $X2=4.14 $Y2=1.95
r98 31 40 3.01263 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.995 $Y=2.12
+ $X2=3.995 $Y2=2.035
r99 31 33 18.0712 $w=4.58e-07 $l=6.95e-07 $layer=LI1_cond $X=3.995 $Y=2.12
+ $X2=3.995 $Y2=2.815
r100 29 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.055 $Y=1.095
+ $X2=4.14 $Y2=1.18
r101 29 30 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=4.055 $Y=1.095
+ $X2=3.655 $Y2=1.095
r102 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.57 $Y=1.01
+ $X2=3.655 $Y2=1.095
r103 27 28 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.57 $Y=0.62
+ $X2=3.57 $Y2=1.01
r104 26 41 7.98728 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=3.095 $Y=2.035
+ $X2=2.81 $Y2=2.035
r105 25 40 3.63293 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.765 $Y=2.035
+ $X2=3.995 $Y2=2.035
r106 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.765 $Y=2.035
+ $X2=3.095 $Y2=2.035
r107 23 49 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.93 $Y=2.815
+ $X2=2.93 $Y2=2.48
r108 20 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=2.395
+ $X2=1.84 $Y2=2.395
r109 19 48 7.98728 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=2.525 $Y=2.395
+ $X2=2.81 $Y2=2.395
r110 19 20 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.525 $Y=2.395
+ $X2=2.005 $Y2=2.395
r111 15 27 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=3.485 $Y=0.485
+ $X2=3.57 $Y2=0.62
r112 15 17 68.2929 $w=2.68e-07 $l=1.6e-06 $layer=LI1_cond $X=3.485 $Y=0.485
+ $X2=1.885 $Y2=0.485
r113 4 40 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=3.795
+ $Y=1.84 $X2=3.93 $Y2=2.115
r114 4 33 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.795
+ $Y=1.84 $X2=3.93 $Y2=2.815
r115 3 44 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=2.745
+ $Y=1.84 $X2=2.93 $Y2=1.985
r116 3 23 600 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=1.84 $X2=2.93 $Y2=2.815
r117 2 38 300 $w=1.7e-07 $l=7.03776e-07 $layer=licon1_PDIFF $count=2 $X=1.695
+ $Y=1.84 $X2=1.84 $Y2=2.475
r118 1 17 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=1.74
+ $Y=0.37 $X2=1.885 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_MS__NAND4BB_1%VGND 1 2 11 13 15 17 19 28 32
r37 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r38 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r39 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r40 25 26 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r41 23 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r42 22 25 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r43 22 23 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r44 20 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=0.815
+ $Y2=0
r45 20 22 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.2
+ $Y2=0
r46 19 31 4.63344 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=3.825 $Y=0 $X2=4.072
+ $Y2=0
r47 19 25 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.825 $Y=0 $X2=3.6
+ $Y2=0
r48 17 26 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r49 17 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r50 13 31 3.13273 $w=3.3e-07 $l=1.19143e-07 $layer=LI1_cond $X=3.99 $Y=0.085
+ $X2=4.072 $Y2=0
r51 13 15 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=3.99 $Y=0.085
+ $X2=3.99 $Y2=0.595
r52 9 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0
r53 9 11 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0.795
r54 2 15 182 $w=1.7e-07 $l=3.81248e-07 $layer=licon1_NDIFF $count=1 $X=3.705
+ $Y=0.37 $X2=3.99 $Y2=0.595
r55 1 11 182 $w=1.7e-07 $l=2.6533e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.695 $X2=0.815 $Y2=0.795
.ends


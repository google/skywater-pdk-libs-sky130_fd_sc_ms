* File: sky130_fd_sc_ms__o211a_4.pex.spice
* Created: Wed Sep  2 12:20:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O211A_4%A_91_48# 1 2 3 4 15 19 23 27 31 35 39 43 45
+ 54 55 56 59 61 66 67 72 74 79 81 90
c173 90 0 1.89035e-19 $X=1.89 $Y=1.465
c174 81 0 5.47072e-20 $X=5.49 $Y=2.115
c175 61 0 8.88359e-21 $X=3.95 $Y=1.195
c176 39 0 1.6164e-19 $X=1.89 $Y=0.74
r177 90 91 16.8994 $w=3.28e-07 $l=1.15e-07 $layer=POLY_cond $X=1.89 $Y=1.465
+ $X2=2.005 $Y2=1.465
r178 87 88 13.9604 $w=3.28e-07 $l=9.5e-08 $layer=POLY_cond $X=1.46 $Y=1.465
+ $X2=1.555 $Y2=1.465
r179 86 87 66.8628 $w=3.28e-07 $l=4.55e-07 $layer=POLY_cond $X=1.005 $Y=1.465
+ $X2=1.46 $Y2=1.465
r180 85 86 6.6128 $w=3.28e-07 $l=4.5e-08 $layer=POLY_cond $X=0.96 $Y=1.465
+ $X2=1.005 $Y2=1.465
r181 82 83 3.67378 $w=3.28e-07 $l=2.5e-08 $layer=POLY_cond $X=0.53 $Y=1.465
+ $X2=0.555 $Y2=1.465
r182 74 76 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.555 $Y=1.105
+ $X2=3.555 $Y2=1.195
r183 68 79 4.30018 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.12 $Y=2.035
+ $X2=3.955 $Y2=2.035
r184 67 81 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.325 $Y=2.035
+ $X2=5.49 $Y2=2.035
r185 67 68 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=5.325 $Y=2.035
+ $X2=4.12 $Y2=2.035
r186 66 79 1.96316 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.035 $Y=1.95
+ $X2=3.955 $Y2=2.035
r187 65 66 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.035 $Y=1.28
+ $X2=4.035 $Y2=1.95
r188 62 76 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.72 $Y=1.195
+ $X2=3.555 $Y2=1.195
r189 61 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.95 $Y=1.195
+ $X2=4.035 $Y2=1.28
r190 61 62 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.95 $Y=1.195
+ $X2=3.72 $Y2=1.195
r191 60 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=2.035
+ $X2=2.94 $Y2=2.035
r192 59 79 4.30018 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.79 $Y=2.035
+ $X2=3.955 $Y2=2.035
r193 59 60 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.79 $Y=2.035
+ $X2=3.105 $Y2=2.035
r194 55 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=2.035
+ $X2=2.94 $Y2=2.035
r195 55 56 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.775 $Y=2.035
+ $X2=2.285 $Y2=2.035
r196 54 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.2 $Y=1.95
+ $X2=2.285 $Y2=2.035
r197 53 54 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.2 $Y=1.63 $X2=2.2
+ $Y2=1.95
r198 52 90 13.2256 $w=3.28e-07 $l=9e-08 $layer=POLY_cond $X=1.8 $Y=1.465
+ $X2=1.89 $Y2=1.465
r199 52 88 36.003 $w=3.28e-07 $l=2.45e-07 $layer=POLY_cond $X=1.8 $Y=1.465
+ $X2=1.555 $Y2=1.465
r200 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.8
+ $Y=1.465 $X2=1.8 $Y2=1.465
r201 48 85 26.4512 $w=3.28e-07 $l=1.8e-07 $layer=POLY_cond $X=0.78 $Y=1.465
+ $X2=0.96 $Y2=1.465
r202 48 83 33.064 $w=3.28e-07 $l=2.25e-07 $layer=POLY_cond $X=0.78 $Y=1.465
+ $X2=0.555 $Y2=1.465
r203 47 51 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=0.78 $Y=1.465
+ $X2=1.8 $Y2=1.465
r204 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.78
+ $Y=1.465 $X2=0.78 $Y2=1.465
r205 45 53 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.115 $Y=1.465
+ $X2=2.2 $Y2=1.63
r206 45 51 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.115 $Y=1.465
+ $X2=1.8 $Y2=1.465
r207 41 91 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.005 $Y=1.63
+ $X2=2.005 $Y2=1.465
r208 41 43 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=2.005 $Y=1.63
+ $X2=2.005 $Y2=2.4
r209 37 90 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=1.3
+ $X2=1.89 $Y2=1.465
r210 37 39 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.89 $Y=1.3
+ $X2=1.89 $Y2=0.74
r211 33 88 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.555 $Y=1.63
+ $X2=1.555 $Y2=1.465
r212 33 35 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.555 $Y=1.63
+ $X2=1.555 $Y2=2.4
r213 29 87 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.46 $Y=1.3
+ $X2=1.46 $Y2=1.465
r214 29 31 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.46 $Y=1.3
+ $X2=1.46 $Y2=0.74
r215 25 86 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.63
+ $X2=1.005 $Y2=1.465
r216 25 27 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.005 $Y=1.63
+ $X2=1.005 $Y2=2.4
r217 21 85 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.3
+ $X2=0.96 $Y2=1.465
r218 21 23 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.96 $Y=1.3
+ $X2=0.96 $Y2=0.74
r219 17 83 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.63
+ $X2=0.555 $Y2=1.465
r220 17 19 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.555 $Y=1.63
+ $X2=0.555 $Y2=2.4
r221 13 82 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.3
+ $X2=0.53 $Y2=1.465
r222 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.53 $Y=1.3
+ $X2=0.53 $Y2=0.74
r223 4 81 300 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_PDIFF $count=2 $X=5.305
+ $Y=1.955 $X2=5.49 $Y2=2.115
r224 3 79 300 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=2 $X=3.82
+ $Y=1.955 $X2=3.955 $Y2=2.115
r225 2 72 300 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=2 $X=2.805
+ $Y=1.955 $X2=2.94 $Y2=2.115
r226 1 74 182 $w=1.7e-07 $l=5.45527e-07 $layer=licon1_NDIFF $count=1 $X=3.415
+ $Y=0.625 $X2=3.555 $Y2=1.105
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_4%C1 1 3 6 8 10 13 15 22
c52 15 0 1.10453e-20 $X=3.6 $Y=1.665
c53 6 0 8.88359e-21 $X=3.34 $Y=0.945
r54 22 23 5.35556 $w=3.6e-07 $l=4e-08 $layer=POLY_cond $X=3.73 $Y=1.665 $X2=3.77
+ $Y2=1.665
r55 20 22 15.3972 $w=3.6e-07 $l=1.15e-07 $layer=POLY_cond $X=3.615 $Y=1.665
+ $X2=3.73 $Y2=1.665
r56 18 20 36.8194 $w=3.6e-07 $l=2.75e-07 $layer=POLY_cond $X=3.34 $Y=1.665
+ $X2=3.615 $Y2=1.665
r57 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.615
+ $Y=1.615 $X2=3.615 $Y2=1.615
r58 11 23 23.3057 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=3.77 $Y=1.45
+ $X2=3.77 $Y2=1.665
r59 11 13 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.77 $Y=1.45
+ $X2=3.77 $Y2=0.945
r60 8 22 18.9685 $w=1.8e-07 $l=2.15e-07 $layer=POLY_cond $X=3.73 $Y=1.88
+ $X2=3.73 $Y2=1.665
r61 8 10 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=3.73 $Y=1.88 $X2=3.73
+ $Y2=2.375
r62 4 18 23.3057 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=3.34 $Y=1.45
+ $X2=3.34 $Y2=1.665
r63 4 6 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.34 $Y=1.45 $X2=3.34
+ $Y2=0.945
r64 1 18 23.4306 $w=3.6e-07 $l=2.89569e-07 $layer=POLY_cond $X=3.165 $Y=1.88
+ $X2=3.34 $Y2=1.665
r65 1 3 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=3.165 $Y=1.88
+ $X2=3.165 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_4%B1 2 3 4 7 9 11 14 19 21 22 28
c81 22 0 1.89035e-19 $X=2.64 $Y=1.665
c82 19 0 2.18884e-20 $X=4.27 $Y=0.945
c83 7 0 4.59574e-20 $X=2.715 $Y=2.375
r84 26 28 5.99171 $w=3.62e-07 $l=4.5e-08 $layer=POLY_cond $X=2.67 $Y=1.552
+ $X2=2.715 $Y2=1.552
r85 24 26 35.9503 $w=3.62e-07 $l=2.7e-07 $layer=POLY_cond $X=2.4 $Y=1.552
+ $X2=2.67 $Y2=1.552
r86 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.67
+ $Y=1.6 $X2=2.67 $Y2=1.6
r87 20 21 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=4.217 $Y=1.34
+ $X2=4.217 $Y2=1.49
r88 19 20 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.27 $Y=0.945
+ $X2=4.27 $Y2=1.34
r89 16 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.27 $Y=0.255
+ $X2=4.27 $Y2=0.945
r90 14 21 344.008 $w=1.8e-07 $l=8.85e-07 $layer=POLY_cond $X=4.18 $Y=2.375
+ $X2=4.18 $Y2=1.49
r91 9 28 25.9641 $w=3.62e-07 $l=2.93741e-07 $layer=POLY_cond $X=2.91 $Y=1.34
+ $X2=2.715 $Y2=1.552
r92 9 11 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.91 $Y=1.34
+ $X2=2.91 $Y2=0.945
r93 5 28 19.0988 $w=1.8e-07 $l=2.13e-07 $layer=POLY_cond $X=2.715 $Y=1.765
+ $X2=2.715 $Y2=1.552
r94 5 7 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=2.715 $Y=1.765
+ $X2=2.715 $Y2=2.375
r95 3 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.195 $Y=0.18
+ $X2=4.27 $Y2=0.255
r96 3 4 881.957 $w=1.5e-07 $l=1.72e-06 $layer=POLY_cond $X=4.195 $Y=0.18
+ $X2=2.475 $Y2=0.18
r97 2 24 23.4391 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=2.4 $Y=1.34 $X2=2.4
+ $Y2=1.552
r98 1 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.4 $Y=0.255
+ $X2=2.475 $Y2=0.18
r99 1 2 556.351 $w=1.5e-07 $l=1.085e-06 $layer=POLY_cond $X=2.4 $Y=0.255 $X2=2.4
+ $Y2=1.34
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_4%A2 3 7 11 15 17 18 25 26
c48 26 0 1.81351e-19 $X=5.715 $Y=1.615
c49 15 0 1.59181e-19 $X=5.725 $Y=0.945
c50 11 0 3.56328e-20 $X=5.715 $Y=2.455
c51 7 0 1.64451e-19 $X=5.24 $Y=0.945
r52 26 27 1.51097 $w=3.19e-07 $l=1e-08 $layer=POLY_cond $X=5.715 $Y=1.615
+ $X2=5.725 $Y2=1.615
r53 24 26 6.79937 $w=3.19e-07 $l=4.5e-08 $layer=POLY_cond $X=5.67 $Y=1.615
+ $X2=5.715 $Y2=1.615
r54 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.67
+ $Y=1.615 $X2=5.67 $Y2=1.615
r55 22 24 64.9718 $w=3.19e-07 $l=4.3e-07 $layer=POLY_cond $X=5.24 $Y=1.615
+ $X2=5.67 $Y2=1.615
r56 21 22 3.77743 $w=3.19e-07 $l=2.5e-08 $layer=POLY_cond $X=5.215 $Y=1.615
+ $X2=5.24 $Y2=1.615
r57 18 25 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=5.52 $Y=1.615
+ $X2=5.67 $Y2=1.615
r58 17 18 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.615
+ $X2=5.52 $Y2=1.615
r59 13 27 20.418 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.725 $Y=1.45
+ $X2=5.725 $Y2=1.615
r60 13 15 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.725 $Y=1.45
+ $X2=5.725 $Y2=0.945
r61 9 26 16.143 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.715 $Y=1.78
+ $X2=5.715 $Y2=1.615
r62 9 11 262.379 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=5.715 $Y=1.78
+ $X2=5.715 $Y2=2.455
r63 5 22 20.418 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.24 $Y=1.45 $X2=5.24
+ $Y2=1.615
r64 5 7 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.24 $Y=1.45 $X2=5.24
+ $Y2=0.945
r65 1 21 16.143 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.215 $Y=1.78
+ $X2=5.215 $Y2=1.615
r66 1 3 262.379 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=5.215 $Y=1.78
+ $X2=5.215 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_4%A1 1 3 8 9 10 13 18 20 23
c63 13 0 5.47072e-20 $X=6.165 $Y=2.455
c64 8 0 1.33941e-19 $X=4.78 $Y=0.945
r65 23 26 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.24 $Y=1.615
+ $X2=6.24 $Y2=1.78
r66 23 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.24 $Y=1.615
+ $X2=6.24 $Y2=1.45
r67 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.24
+ $Y=1.615 $X2=6.24 $Y2=1.615
r68 20 24 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=6.48 $Y=1.615
+ $X2=6.24 $Y2=1.615
r69 18 25 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.225 $Y=0.945
+ $X2=6.225 $Y2=1.45
r70 15 18 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.225 $Y=0.255
+ $X2=6.225 $Y2=0.945
r71 13 26 262.379 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=6.165 $Y=2.455
+ $X2=6.165 $Y2=1.78
r72 9 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.15 $Y=0.18
+ $X2=6.225 $Y2=0.255
r73 9 10 664.032 $w=1.5e-07 $l=1.295e-06 $layer=POLY_cond $X=6.15 $Y=0.18
+ $X2=4.855 $Y2=0.18
r74 8 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.78 $Y=0.945
+ $X2=4.78 $Y2=1.34
r75 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.78 $Y=0.255
+ $X2=4.855 $Y2=0.18
r76 5 8 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.78 $Y=0.255 $X2=4.78
+ $Y2=0.945
r77 1 19 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.765 $Y=1.43 $X2=4.765
+ $Y2=1.34
r78 1 3 398.427 $w=1.8e-07 $l=1.025e-06 $layer=POLY_cond $X=4.765 $Y=1.43
+ $X2=4.765 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_4%VPWR 1 2 3 4 5 6 19 21 25 27 31 37 41 45 47
+ 52 53 54 56 65 69 81 84 87 91
r94 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r95 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r96 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r97 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r98 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r99 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r100 76 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r101 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r102 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r103 73 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r104 72 75 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r105 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r106 70 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.655 $Y=3.33
+ $X2=4.49 $Y2=3.33
r107 70 72 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.655 $Y=3.33
+ $X2=5.04 $Y2=3.33
r108 69 90 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6.497 $Y2=3.33
r109 69 75 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6 $Y2=3.33
r110 68 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r111 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r112 65 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.325 $Y=3.33
+ $X2=4.49 $Y2=3.33
r113 65 67 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.325 $Y=3.33
+ $X2=4.08 $Y2=3.33
r114 64 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r115 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r116 61 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=2.28 $Y2=3.33
r117 61 63 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.445 $Y=3.33
+ $X2=3.12 $Y2=3.33
r118 60 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r119 60 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r120 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r121 57 78 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r122 57 59 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r123 56 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=1.28 $Y2=3.33
r124 56 59 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=0.72 $Y2=3.33
r125 54 68 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.08 $Y2=3.33
r126 54 64 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r127 52 63 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.275 $Y=3.33
+ $X2=3.12 $Y2=3.33
r128 52 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.275 $Y=3.33
+ $X2=3.44 $Y2=3.33
r129 51 67 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.605 $Y=3.33
+ $X2=4.08 $Y2=3.33
r130 51 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.605 $Y=3.33
+ $X2=3.44 $Y2=3.33
r131 47 50 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=6.44 $Y=2.115
+ $X2=6.44 $Y2=2.81
r132 45 90 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=6.44 $Y=3.245
+ $X2=6.497 $Y2=3.33
r133 45 50 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=6.44 $Y=3.245
+ $X2=6.44 $Y2=2.81
r134 41 44 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=4.49 $Y=2.41 $X2=4.49
+ $Y2=2.81
r135 39 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=3.245
+ $X2=4.49 $Y2=3.33
r136 39 44 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=4.49 $Y=3.245
+ $X2=4.49 $Y2=2.81
r137 35 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=3.245
+ $X2=3.44 $Y2=3.33
r138 35 37 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=3.44 $Y=3.245
+ $X2=3.44 $Y2=2.455
r139 31 34 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.28 $Y=2.405
+ $X2=2.28 $Y2=2.815
r140 29 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=3.245
+ $X2=2.28 $Y2=3.33
r141 29 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.28 $Y=3.245
+ $X2=2.28 $Y2=2.815
r142 28 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=3.33
+ $X2=1.28 $Y2=3.33
r143 27 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=3.33
+ $X2=2.28 $Y2=3.33
r144 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.115 $Y=3.33
+ $X2=1.445 $Y2=3.33
r145 23 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=3.245
+ $X2=1.28 $Y2=3.33
r146 23 25 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=1.28 $Y=3.245
+ $X2=1.28 $Y2=2.305
r147 19 78 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r148 19 21 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.305
r149 6 50 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=6.255
+ $Y=1.955 $X2=6.44 $Y2=2.81
r150 6 47 400 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_PDIFF $count=1 $X=6.255
+ $Y=1.955 $X2=6.44 $Y2=2.115
r151 5 44 600 $w=1.7e-07 $l=9.5871e-07 $layer=licon1_PDIFF $count=1 $X=4.27
+ $Y=1.955 $X2=4.49 $Y2=2.81
r152 5 41 600 $w=1.7e-07 $l=5.54189e-07 $layer=licon1_PDIFF $count=1 $X=4.27
+ $Y=1.955 $X2=4.49 $Y2=2.41
r153 4 37 600 $w=1.7e-07 $l=5.85235e-07 $layer=licon1_PDIFF $count=1 $X=3.255
+ $Y=1.955 $X2=3.44 $Y2=2.455
r154 3 34 600 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=2.095
+ $Y=1.84 $X2=2.28 $Y2=2.815
r155 3 31 600 $w=1.7e-07 $l=6.50961e-07 $layer=licon1_PDIFF $count=1 $X=2.095
+ $Y=1.84 $X2=2.28 $Y2=2.405
r156 2 25 300 $w=1.7e-07 $l=5.49773e-07 $layer=licon1_PDIFF $count=2 $X=1.095
+ $Y=1.84 $X2=1.28 $Y2=2.305
r157 1 21 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.305
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_4%X 1 2 3 4 13 14 15 16 19 23 27 29 33 37 43
+ 44 45 46
c78 29 0 3.49122e-20 $X=1.615 $Y=1.885
c79 27 0 1.6164e-19 $X=1.51 $Y=1.045
r80 45 46 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r81 42 46 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.24 $Y=1.8
+ $X2=0.24 $Y2=1.665
r82 41 45 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.13
+ $X2=0.24 $Y2=1.295
r83 37 39 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.78 $Y=1.985
+ $X2=1.78 $Y2=2.815
r84 35 37 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.78 $Y=1.97
+ $X2=1.78 $Y2=1.985
r85 31 33 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=1.635 $Y=0.96
+ $X2=1.635 $Y2=0.515
r86 30 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=1.885
+ $X2=0.78 $Y2=1.885
r87 29 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.615 $Y=1.885
+ $X2=1.78 $Y2=1.97
r88 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=1.885
+ $X2=0.945 $Y2=1.885
r89 28 43 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.83 $Y=1.045
+ $X2=0.705 $Y2=1.045
r90 27 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.51 $Y=1.045
+ $X2=1.635 $Y2=0.96
r91 27 28 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.51 $Y=1.045
+ $X2=0.83 $Y2=1.045
r92 23 25 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.78 $Y=1.985
+ $X2=0.78 $Y2=2.815
r93 21 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=1.97 $X2=0.78
+ $Y2=1.885
r94 21 23 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.78 $Y=1.97
+ $X2=0.78 $Y2=1.985
r95 17 43 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.96
+ $X2=0.705 $Y2=1.045
r96 17 19 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.705 $Y=0.96
+ $X2=0.705 $Y2=0.515
r97 16 42 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.885
+ $X2=0.24 $Y2=1.8
r98 15 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=1.885
+ $X2=0.78 $Y2=1.885
r99 15 16 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.615 $Y=1.885
+ $X2=0.355 $Y2=1.885
r100 14 41 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.045
+ $X2=0.24 $Y2=1.13
r101 13 43 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.58 $Y=1.045
+ $X2=0.705 $Y2=1.045
r102 13 14 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.58 $Y=1.045
+ $X2=0.355 $Y2=1.045
r103 4 39 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.645
+ $Y=1.84 $X2=1.78 $Y2=2.815
r104 4 37 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.645
+ $Y=1.84 $X2=1.78 $Y2=1.985
r105 3 25 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.645
+ $Y=1.84 $X2=0.78 $Y2=2.815
r106 3 23 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.645
+ $Y=1.84 $X2=0.78 $Y2=1.985
r107 2 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.535
+ $Y=0.37 $X2=1.675 $Y2=0.515
r108 1 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.605
+ $Y=0.37 $X2=0.745 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_4%A_971_391# 1 2 9 11 12 15
c26 15 0 3.56328e-20 $X=5.94 $Y=2.115
r27 15 18 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=5.98 $Y=2.115
+ $X2=5.98 $Y2=2.81
r28 13 18 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=5.98 $Y=2.905
+ $X2=5.98 $Y2=2.81
r29 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.855 $Y=2.99
+ $X2=5.98 $Y2=2.905
r30 11 12 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.855 $Y=2.99
+ $X2=5.155 $Y2=2.99
r31 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.99 $Y=2.905
+ $X2=5.155 $Y2=2.99
r32 7 9 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.99 $Y=2.905
+ $X2=4.99 $Y2=2.41
r33 2 18 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.955 $X2=5.94 $Y2=2.81
r34 2 15 400 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.955 $X2=5.94 $Y2=2.115
r35 1 9 300 $w=1.7e-07 $l=5.18122e-07 $layer=licon1_PDIFF $count=2 $X=4.855
+ $Y=1.955 $X2=4.99 $Y2=2.41
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_4%VGND 1 2 3 4 5 16 18 22 26 30 34 36 38 43 48
+ 56 63 64 70 73 76 79
r88 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r89 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r90 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r91 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r92 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r93 64 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r94 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r95 61 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.105 $Y=0 $X2=5.94
+ $Y2=0
r96 61 63 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.105 $Y=0 $X2=6.48
+ $Y2=0
r97 60 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r98 60 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r99 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r100 57 76 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=5.175 $Y=0
+ $X2=5.002 $Y2=0
r101 57 59 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.175 $Y=0 $X2=5.52
+ $Y2=0
r102 56 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.775 $Y=0 $X2=5.94
+ $Y2=0
r103 56 59 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.775 $Y=0
+ $X2=5.52 $Y2=0
r104 55 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r105 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r106 52 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r107 51 54 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r108 51 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r109 49 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.105
+ $Y2=0
r110 49 51 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.64
+ $Y2=0
r111 48 76 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=5.002
+ $Y2=0
r112 48 54 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=4.56
+ $Y2=0
r113 47 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r114 47 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r115 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r116 44 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.34 $Y=0 $X2=1.175
+ $Y2=0
r117 44 46 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.34 $Y=0 $X2=1.68
+ $Y2=0
r118 43 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=2.105
+ $Y2=0
r119 43 46 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=1.68
+ $Y2=0
r120 42 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r121 42 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r122 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r123 39 67 3.96842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.4 $Y=0 $X2=0.2 $Y2=0
r124 39 41 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.4 $Y=0 $X2=0.72
+ $Y2=0
r125 38 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=1.175
+ $Y2=0
r126 38 41 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=0.72
+ $Y2=0
r127 36 55 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.56
+ $Y2=0
r128 36 52 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=2.64
+ $Y2=0
r129 32 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.94 $Y=0.085
+ $X2=5.94 $Y2=0
r130 32 34 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=5.94 $Y=0.085
+ $X2=5.94 $Y2=0.77
r131 28 76 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=5.002 $Y=0.085
+ $X2=5.002 $Y2=0
r132 28 30 22.8818 $w=3.43e-07 $l=6.85e-07 $layer=LI1_cond $X=5.002 $Y=0.085
+ $X2=5.002 $Y2=0.77
r133 24 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0
r134 24 26 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0.515
r135 20 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=0.085
+ $X2=1.175 $Y2=0
r136 20 22 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=1.175 $Y=0.085
+ $X2=1.175 $Y2=0.57
r137 16 67 3.17474 $w=2.5e-07 $l=1.16619e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.2 $Y2=0
r138 16 18 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.57
r139 5 34 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.8
+ $Y=0.625 $X2=5.94 $Y2=0.77
r140 4 30 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=4.855
+ $Y=0.625 $X2=5 $Y2=0.77
r141 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.965
+ $Y=0.37 $X2=2.105 $Y2=0.515
r142 2 22 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.37 $X2=1.175 $Y2=0.57
r143 1 18 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=0.17
+ $Y=0.37 $X2=0.315 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_4%A_510_125# 1 2 3 4 15 17 18 22 23 24 27 29
+ 33 35
c72 27 0 3.23633e-19 $X=5.51 $Y=0.77
c73 24 0 1.33941e-19 $X=4.65 $Y=1.195
c74 23 0 1.81351e-19 $X=5.345 $Y=1.195
r75 31 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=6.44 $Y=1.11
+ $X2=6.44 $Y2=0.77
r76 30 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.595 $Y=1.195
+ $X2=5.47 $Y2=1.195
r77 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.275 $Y=1.195
+ $X2=6.44 $Y2=1.11
r78 29 30 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.275 $Y=1.195
+ $X2=5.595 $Y2=1.195
r79 25 35 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.47 $Y=1.11
+ $X2=5.47 $Y2=1.195
r80 25 27 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=5.47 $Y=1.11
+ $X2=5.47 $Y2=0.77
r81 23 35 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.345 $Y=1.195
+ $X2=5.47 $Y2=1.195
r82 23 24 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=5.345 $Y=1.195
+ $X2=4.65 $Y2=1.195
r83 20 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.525 $Y=1.11
+ $X2=4.65 $Y2=1.195
r84 20 22 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=4.525 $Y=1.11
+ $X2=4.525 $Y2=0.77
r85 19 22 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=4.525 $Y=0.425
+ $X2=4.525 $Y2=0.77
r86 17 19 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.4 $Y=0.34
+ $X2=4.525 $Y2=0.425
r87 17 18 105.69 $w=1.68e-07 $l=1.62e-06 $layer=LI1_cond $X=4.4 $Y=0.34 $X2=2.78
+ $Y2=0.34
r88 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.655 $Y=0.425
+ $X2=2.78 $Y2=0.34
r89 13 15 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.655 $Y=0.425
+ $X2=2.655 $Y2=0.76
r90 4 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.3
+ $Y=0.625 $X2=6.44 $Y2=0.77
r91 3 27 91 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=2 $X=5.315
+ $Y=0.625 $X2=5.51 $Y2=0.77
r92 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.345
+ $Y=0.625 $X2=4.485 $Y2=0.77
r93 1 15 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.55
+ $Y=0.625 $X2=2.695 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_4%A_597_125# 1 2 9 11 12 13
c26 11 0 2.18884e-20 $X=3.89 $Y=0.68
r27 13 16 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.055 $Y=0.68
+ $X2=4.055 $Y2=0.77
r28 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.89 $Y=0.68
+ $X2=4.055 $Y2=0.68
r29 11 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.89 $Y=0.68
+ $X2=3.21 $Y2=0.68
r30 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.125 $Y=0.765
+ $X2=3.21 $Y2=0.68
r31 7 9 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.125 $Y=0.765
+ $X2=3.125 $Y2=0.77
r32 2 16 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.845
+ $Y=0.625 $X2=4.055 $Y2=0.77
r33 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.985
+ $Y=0.625 $X2=3.125 $Y2=0.77
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
M1000 a_1278_74# a_612_74# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.6502e+12p ps=1.426e+07u
M1001 a_1356_74# a_398_74# a_1278_74# VNB nlowvt w=640000u l=150000u
+  ad=2.713e+11p pd=2.31e+06u as=0p ps=0u
M1002 a_1057_118# a_612_74# a_767_384# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1003 a_1356_74# a_225_74# a_1269_341# VPB pshort w=1e+06u l=180000u
+  ad=5.278e+11p pd=4.58e+06u as=3.69625e+11p ps=3.16e+06u
M1004 VGND SET_B a_1596_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.764e+11p ps=1.68e+06u
M1005 VGND a_2022_94# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1006 VPWR a_1356_74# a_2022_94# VPB pshort w=1e+06u l=180000u
+  ad=2.34017e+12p pd=1.968e+07u as=2.8e+11p ps=2.56e+06u
M1007 a_1356_74# SET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_1489_118# a_225_74# a_1356_74# VNB nlowvt w=420000u l=150000u
+  ad=1.617e+11p pd=1.61e+06u as=0p ps=0u
M1009 a_767_384# a_612_74# VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1010 a_1524_508# a_398_74# a_1356_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1011 a_1269_341# a_612_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_781_74# a_398_74# a_612_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.919e+11p ps=2.23e+06u
M1013 VGND a_1356_74# a_2022_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1014 VPWR CLK a_225_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1015 a_398_74# a_225_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1016 VPWR SET_B a_767_384# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_398_74# a_225_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1018 a_612_74# a_225_74# a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=3.0635e+11p ps=3.21e+06u
M1019 a_1566_92# a_1356_74# VPWR VPB pshort w=420000u l=180000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1020 VPWR D a_27_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.8e+06u
M1021 a_719_456# a_225_74# a_612_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=1.344e+11p ps=1.48e+06u
M1022 VGND SET_B a_1057_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_612_74# a_398_74# a_27_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_767_384# a_781_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Q a_2022_94# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Q a_2022_94# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1027 a_1566_92# a_1356_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1028 VPWR a_1566_92# a_1524_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_2022_94# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1596_118# a_1566_92# a_1489_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND D a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR a_767_384# a_719_456# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND CLK a_225_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
.ends

* File: sky130_fd_sc_ms__o21ba_1.spice
* Created: Wed Sep  2 12:22:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o21ba_1.pex.spice"
.subckt sky130_fd_sc_ms__o21ba_1  VNB VPB A1 A2 B1_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1_N	B1_N
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A1_M1008_g N_A_27_74#_M1008_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1344 AS=0.1824 PD=1.06 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.3 A=0.096 P=1.58 MULT=1
MM1009 N_A_27_74#_M1009_d N_A2_M1009_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0944 AS=0.1344 PD=0.935 PS=1.06 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75000.8
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1005 N_A_203_392#_M1005_d N_A_281_244#_M1005_g N_A_27_74#_M1009_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.2176 AS=0.0944 PD=1.96 PS=0.935 NRD=10.308 NRS=2.808 M=1
+ R=4.26667 SA=75001.2 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1006_d N_B1_N_M1006_g N_A_281_244#_M1006_s VNB NLOWVT L=0.15
+ W=0.55 AD=0.123601 AS=0.275 PD=0.989147 PS=2.1 NRD=23.448 NRS=0 M=1 R=3.66667
+ SA=75000.4 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1001 N_X_M1001_d N_A_203_392#_M1001_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.166299 PD=2.05 PS=1.33085 NRD=0 NRS=5.664 M=1 R=4.93333
+ SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 A_119_392# N_A1_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.28 PD=1.24 PS=2.56 NRD=12.7853 NRS=0 M=1 R=5.55556 SA=90000.2 SB=90001.2
+ A=0.18 P=2.36 MULT=1
MM1003 N_A_203_392#_M1003_d N_A2_M1003_g A_119_392# VPB PSHORT L=0.18 W=1
+ AD=0.195 AS=0.12 PD=1.39 PS=1.24 NRD=12.7853 NRS=12.7853 M=1 R=5.55556
+ SA=90000.6 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_A_281_244#_M1004_g N_A_203_392#_M1003_d VPB PSHORT
+ L=0.18 W=1 AD=0.28 AS=0.195 PD=2.56 PS=1.39 NRD=0 NRS=8.8453 M=1 R=5.55556
+ SA=90001.2 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_B1_N_M1007_g N_A_281_244#_M1007_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1854 AS=0.2982 PD=1.30714 PS=2.39 NRD=38.8484 NRS=0 M=1 R=4.66667
+ SA=90000.3 SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1000 N_X_M1000_d N_A_203_392#_M1000_g N_VPWR_M1007_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.2472 PD=2.8 PS=1.74286 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90000.7 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ms__o21ba_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__o41ai_1.pxi.spice
* Created: Fri Aug 28 18:05:24 2020
* 
x_PM_SKY130_FD_SC_MS__O41AI_1%B1 N_B1_c_62_n N_B1_M1009_g N_B1_M1006_g
+ N_B1_c_64_n N_B1_c_65_n B1 PM_SKY130_FD_SC_MS__O41AI_1%B1
x_PM_SKY130_FD_SC_MS__O41AI_1%A4 N_A4_M1005_g N_A4_M1008_g A4 N_A4_c_100_n
+ N_A4_c_101_n PM_SKY130_FD_SC_MS__O41AI_1%A4
x_PM_SKY130_FD_SC_MS__O41AI_1%A3 N_A3_M1002_g N_A3_M1003_g A3 A3 A3 A3
+ N_A3_c_146_n N_A3_c_147_n PM_SKY130_FD_SC_MS__O41AI_1%A3
x_PM_SKY130_FD_SC_MS__O41AI_1%A2 N_A2_M1007_g N_A2_M1001_g N_A2_c_192_n
+ N_A2_c_193_n A2 A2 A2 N_A2_c_197_n A2 PM_SKY130_FD_SC_MS__O41AI_1%A2
x_PM_SKY130_FD_SC_MS__O41AI_1%A1 N_A1_M1000_g N_A1_M1004_g A1 N_A1_c_235_n
+ N_A1_c_236_n PM_SKY130_FD_SC_MS__O41AI_1%A1
x_PM_SKY130_FD_SC_MS__O41AI_1%VPWR N_VPWR_M1006_s N_VPWR_M1004_d N_VPWR_c_263_n
+ N_VPWR_c_264_n N_VPWR_c_265_n N_VPWR_c_266_n N_VPWR_c_267_n VPWR
+ N_VPWR_c_268_n N_VPWR_c_262_n PM_SKY130_FD_SC_MS__O41AI_1%VPWR
x_PM_SKY130_FD_SC_MS__O41AI_1%Y N_Y_M1009_s N_Y_M1006_d N_Y_c_297_n N_Y_c_301_n
+ N_Y_c_298_n N_Y_c_310_n N_Y_c_299_n Y N_Y_c_300_n
+ PM_SKY130_FD_SC_MS__O41AI_1%Y
x_PM_SKY130_FD_SC_MS__O41AI_1%A_157_74# N_A_157_74#_M1009_d N_A_157_74#_M1003_d
+ N_A_157_74#_M1000_d N_A_157_74#_c_342_n N_A_157_74#_c_343_n
+ N_A_157_74#_c_344_n N_A_157_74#_c_345_n N_A_157_74#_c_346_n
+ N_A_157_74#_c_347_n N_A_157_74#_c_348_n PM_SKY130_FD_SC_MS__O41AI_1%A_157_74#
x_PM_SKY130_FD_SC_MS__O41AI_1%VGND N_VGND_M1008_d N_VGND_M1007_d N_VGND_c_395_n
+ N_VGND_c_396_n N_VGND_c_397_n N_VGND_c_398_n N_VGND_c_399_n N_VGND_c_400_n
+ VGND N_VGND_c_401_n N_VGND_c_402_n PM_SKY130_FD_SC_MS__O41AI_1%VGND
cc_1 VNB N_B1_c_62_n 0.0231039f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.22
cc_2 VNB N_B1_M1006_g 0.00857766f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.4
cc_3 VNB N_B1_c_64_n 0.0679577f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.385
cc_4 VNB N_B1_c_65_n 0.013281f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.385
cc_5 VNB B1 0.00924172f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_A4_M1008_g 0.0272905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A4_c_100_n 0.0269258f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_8 VNB N_A4_c_101_n 0.00165618f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_9 VNB N_A3_M1003_g 0.0259452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A3_c_146_n 0.0226552f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_11 VNB N_A3_c_147_n 0.00442043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_M1007_g 0.0257812f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.74
cc_13 VNB N_A2_c_192_n 0.00484184f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_14 VNB N_A2_c_193_n 0.0224352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A1_M1000_g 0.0348798f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.74
cc_16 VNB N_A1_c_235_n 0.0331631f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_17 VNB N_A1_c_236_n 0.015292f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_18 VNB N_VPWR_c_262_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_297_n 0.00273786f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.385
cc_20 VNB N_Y_c_298_n 0.0036177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_299_n 0.0010381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_300_n 0.0380313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_157_74#_c_342_n 0.00207713f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_24 VNB N_A_157_74#_c_343_n 0.00809218f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_25 VNB N_A_157_74#_c_344_n 0.00541064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_157_74#_c_345_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_157_74#_c_346_n 0.0188655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_157_74#_c_347_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_157_74#_c_348_n 0.00781721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_395_n 0.00977876f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.385
cc_31 VNB N_VGND_c_396_n 0.00970653f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_32 VNB N_VGND_c_397_n 0.0388991f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_33 VNB N_VGND_c_398_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_399_n 0.0191721f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_35 VNB N_VGND_c_400_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_401_n 0.0199471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_402_n 0.215861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_B1_M1006_g 0.028912f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=2.4
cc_39 VPB N_A4_M1005_g 0.0221556f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=0.74
cc_40 VPB N_A4_c_100_n 0.00562503f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_41 VPB N_A4_c_101_n 0.00466172f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_42 VPB N_A3_M1002_g 0.0231826f $X=-0.19 $Y=1.66 $X2=0.71 $Y2=0.74
cc_43 VPB A3 0.00144367f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.385
cc_44 VPB N_A3_c_146_n 0.00926256f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_45 VPB N_A3_c_147_n 4.05978e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A2_M1001_g 0.0240144f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A2_c_192_n 4.54806e-19 $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_48 VPB N_A2_c_193_n 0.00879672f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A2_c_197_n 0.00150467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A1_M1004_g 0.0268938f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A1_c_235_n 0.00728271f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_52 VPB N_A1_c_236_n 0.00879038f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_53 VPB N_VPWR_c_263_n 0.0366597f $X=-0.19 $Y=1.66 $X2=0.725 $Y2=1.385
cc_54 VPB N_VPWR_c_264_n 0.0301664f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_55 VPB N_VPWR_c_265_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_56 VPB N_VPWR_c_266_n 0.0499543f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_267_n 0.0111029f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_268_n 0.0682324f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_262_n 0.0872524f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_Y_c_301_n 0.00275675f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_61 VPB N_Y_c_299_n 0.00135795f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 N_B1_M1006_g N_A4_M1005_g 0.013876f $X=0.725 $Y=2.4 $X2=0 $Y2=0
cc_63 N_B1_c_62_n N_A4_M1008_g 0.015975f $X=0.71 $Y=1.22 $X2=0 $Y2=0
cc_64 N_B1_c_65_n N_A4_M1008_g 0.00510291f $X=0.725 $Y=1.385 $X2=0 $Y2=0
cc_65 N_B1_c_65_n N_A4_c_100_n 0.0174074f $X=0.725 $Y=1.385 $X2=0 $Y2=0
cc_66 N_B1_M1006_g N_A4_c_101_n 3.06787e-19 $X=0.725 $Y=2.4 $X2=0 $Y2=0
cc_67 N_B1_c_65_n N_A4_c_101_n 3.60864e-19 $X=0.725 $Y=1.385 $X2=0 $Y2=0
cc_68 N_B1_M1006_g N_VPWR_c_263_n 0.00503518f $X=0.725 $Y=2.4 $X2=0 $Y2=0
cc_69 N_B1_c_64_n N_VPWR_c_263_n 0.00677105f $X=0.635 $Y=1.385 $X2=0 $Y2=0
cc_70 B1 N_VPWR_c_263_n 0.0192059f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_71 N_B1_M1006_g N_VPWR_c_264_n 0.00644626f $X=0.725 $Y=2.4 $X2=0 $Y2=0
cc_72 N_B1_M1006_g N_VPWR_c_267_n 0.00455257f $X=0.725 $Y=2.4 $X2=0 $Y2=0
cc_73 N_B1_M1006_g N_VPWR_c_268_n 0.00460063f $X=0.725 $Y=2.4 $X2=0 $Y2=0
cc_74 N_B1_M1006_g N_VPWR_c_262_n 0.00909121f $X=0.725 $Y=2.4 $X2=0 $Y2=0
cc_75 N_B1_c_62_n N_Y_c_297_n 0.00627667f $X=0.71 $Y=1.22 $X2=0 $Y2=0
cc_76 N_B1_c_64_n N_Y_c_297_n 0.00298425f $X=0.635 $Y=1.385 $X2=0 $Y2=0
cc_77 N_B1_c_65_n N_Y_c_297_n 0.00402065f $X=0.725 $Y=1.385 $X2=0 $Y2=0
cc_78 B1 N_Y_c_297_n 0.0124545f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_79 N_B1_c_64_n N_Y_c_298_n 0.00392281f $X=0.635 $Y=1.385 $X2=0 $Y2=0
cc_80 N_B1_c_65_n N_Y_c_298_n 0.00952428f $X=0.725 $Y=1.385 $X2=0 $Y2=0
cc_81 B1 N_Y_c_298_n 0.0125167f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_82 N_B1_M1006_g N_Y_c_310_n 0.00782039f $X=0.725 $Y=2.4 $X2=0 $Y2=0
cc_83 N_B1_M1006_g N_Y_c_299_n 0.0167424f $X=0.725 $Y=2.4 $X2=0 $Y2=0
cc_84 N_B1_c_65_n N_Y_c_299_n 0.00134511f $X=0.725 $Y=1.385 $X2=0 $Y2=0
cc_85 B1 N_Y_c_299_n 0.00143785f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_86 N_B1_c_62_n N_Y_c_300_n 0.013685f $X=0.71 $Y=1.22 $X2=0 $Y2=0
cc_87 N_B1_c_64_n N_Y_c_300_n 0.00875781f $X=0.635 $Y=1.385 $X2=0 $Y2=0
cc_88 B1 N_Y_c_300_n 0.0273814f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_89 N_B1_c_62_n N_A_157_74#_c_342_n 0.00464354f $X=0.71 $Y=1.22 $X2=0 $Y2=0
cc_90 N_B1_c_62_n N_A_157_74#_c_344_n 0.00131473f $X=0.71 $Y=1.22 $X2=0 $Y2=0
cc_91 N_B1_c_62_n N_VGND_c_397_n 0.00303976f $X=0.71 $Y=1.22 $X2=0 $Y2=0
cc_92 N_B1_c_62_n N_VGND_c_402_n 0.00404638f $X=0.71 $Y=1.22 $X2=0 $Y2=0
cc_93 N_A4_M1005_g N_A3_M1002_g 0.0534653f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_94 N_A4_c_101_n N_A3_M1002_g 3.15742e-19 $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_95 N_A4_M1008_g N_A3_M1003_g 0.0248295f $X=1.255 $Y=0.74 $X2=0 $Y2=0
cc_96 N_A4_M1005_g A3 0.0108981f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_97 N_A4_c_101_n A3 0.00778316f $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_98 N_A4_c_100_n N_A3_c_146_n 0.0174403f $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_99 N_A4_c_101_n N_A3_c_146_n 3.70595e-19 $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_100 N_A4_c_100_n N_A3_c_147_n 0.00201946f $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_101 N_A4_c_101_n N_A3_c_147_n 0.0253181f $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_102 N_A4_M1005_g N_VPWR_c_264_n 5.24148e-19 $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_103 N_A4_M1005_g N_VPWR_c_268_n 0.005209f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_104 N_A4_M1005_g N_VPWR_c_262_n 0.00984408f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_105 N_A4_M1008_g N_Y_c_297_n 9.38286e-19 $X=1.255 $Y=0.74 $X2=0 $Y2=0
cc_106 N_A4_M1005_g N_Y_c_301_n 0.014833f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_107 N_A4_c_100_n N_Y_c_298_n 9.98351e-19 $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_108 N_A4_c_101_n N_Y_c_298_n 0.0131895f $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_109 N_A4_M1005_g N_Y_c_310_n 0.00318117f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_110 N_A4_c_100_n N_Y_c_310_n 3.43696e-19 $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_111 N_A4_c_101_n N_Y_c_310_n 0.00677624f $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_112 N_A4_M1005_g N_Y_c_299_n 0.0034284f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_113 N_A4_c_100_n N_Y_c_299_n 9.07691e-19 $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_114 N_A4_c_101_n N_Y_c_299_n 0.0199516f $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_115 N_A4_M1008_g N_Y_c_300_n 3.37387e-19 $X=1.255 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A4_M1008_g N_A_157_74#_c_342_n 0.00959047f $X=1.255 $Y=0.74 $X2=0 $Y2=0
cc_117 N_A4_M1008_g N_A_157_74#_c_343_n 0.0118537f $X=1.255 $Y=0.74 $X2=0 $Y2=0
cc_118 N_A4_c_100_n N_A_157_74#_c_343_n 3.80672e-19 $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_119 N_A4_c_101_n N_A_157_74#_c_343_n 0.0132954f $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_120 N_A4_M1008_g N_A_157_74#_c_344_n 0.00154351f $X=1.255 $Y=0.74 $X2=0 $Y2=0
cc_121 N_A4_c_100_n N_A_157_74#_c_344_n 9.77176e-19 $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_122 N_A4_c_101_n N_A_157_74#_c_344_n 0.0127466f $X=1.22 $Y=1.515 $X2=0 $Y2=0
cc_123 N_A4_M1008_g N_A_157_74#_c_345_n 8.69432e-19 $X=1.255 $Y=0.74 $X2=0 $Y2=0
cc_124 N_A4_M1008_g N_VGND_c_395_n 0.00633237f $X=1.255 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A4_M1008_g N_VGND_c_397_n 0.00434272f $X=1.255 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A4_M1008_g N_VGND_c_402_n 0.00822486f $X=1.255 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A3_M1003_g N_A2_M1007_g 0.0199862f $X=1.84 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A3_M1002_g N_A2_M1001_g 0.0396048f $X=1.715 $Y=2.4 $X2=0 $Y2=0
cc_129 A3 N_A2_M1001_g 0.00127861f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_130 N_A3_c_146_n N_A2_c_192_n 0.00114507f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_131 N_A3_c_147_n N_A2_c_192_n 0.0269386f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_132 N_A3_c_146_n N_A2_c_193_n 0.0181729f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_133 N_A3_c_147_n N_A2_c_193_n 3.62017e-19 $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_134 N_A3_M1002_g A2 0.00683904f $X=1.715 $Y=2.4 $X2=0 $Y2=0
cc_135 A3 A2 0.0533612f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_136 N_A3_M1002_g N_A2_c_197_n 0.00156129f $X=1.715 $Y=2.4 $X2=0 $Y2=0
cc_137 A3 N_A2_c_197_n 0.0105527f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_138 N_A3_M1002_g N_VPWR_c_268_n 0.00375551f $X=1.715 $Y=2.4 $X2=0 $Y2=0
cc_139 A3 N_VPWR_c_268_n 0.00607813f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_140 N_A3_M1002_g N_VPWR_c_262_n 0.00485634f $X=1.715 $Y=2.4 $X2=0 $Y2=0
cc_141 A3 N_VPWR_c_262_n 0.0070933f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_142 N_A3_M1002_g N_Y_c_301_n 4.22454e-19 $X=1.715 $Y=2.4 $X2=0 $Y2=0
cc_143 N_A3_M1002_g N_Y_c_310_n 9.05389e-19 $X=1.715 $Y=2.4 $X2=0 $Y2=0
cc_144 A3 N_Y_c_310_n 0.0368493f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_145 A3 A_263_368# 0.0131286f $X=1.595 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_146 N_A3_M1003_g N_A_157_74#_c_342_n 8.64759e-19 $X=1.84 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A3_M1003_g N_A_157_74#_c_343_n 0.0118588f $X=1.84 $Y=0.74 $X2=0 $Y2=0
cc_148 N_A3_c_146_n N_A_157_74#_c_343_n 0.00369047f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_149 N_A3_c_147_n N_A_157_74#_c_343_n 0.0241717f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_150 N_A3_M1003_g N_A_157_74#_c_345_n 0.00988375f $X=1.84 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A3_M1003_g N_A_157_74#_c_348_n 0.00155819f $X=1.84 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A3_c_146_n N_A_157_74#_c_348_n 9.31826e-19 $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_153 N_A3_c_147_n N_A_157_74#_c_348_n 0.00536895f $X=1.79 $Y=1.515 $X2=0 $Y2=0
cc_154 N_A3_M1003_g N_VGND_c_395_n 0.00781129f $X=1.84 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A3_M1003_g N_VGND_c_399_n 0.00434272f $X=1.84 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A3_M1003_g N_VGND_c_402_n 0.00821853f $X=1.84 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A2_M1007_g N_A1_M1000_g 0.0260254f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A2_M1001_g N_A1_M1004_g 0.0419562f $X=2.285 $Y=2.4 $X2=0 $Y2=0
cc_159 N_A2_c_197_n N_A1_M1004_g 0.00603112f $X=2.17 $Y=1.92 $X2=0 $Y2=0
cc_160 N_A2_c_192_n N_A1_c_235_n 0.00127309f $X=2.36 $Y=1.515 $X2=0 $Y2=0
cc_161 N_A2_c_193_n N_A1_c_235_n 0.0178053f $X=2.36 $Y=1.515 $X2=0 $Y2=0
cc_162 N_A2_M1001_g N_A1_c_236_n 3.54703e-19 $X=2.285 $Y=2.4 $X2=0 $Y2=0
cc_163 N_A2_c_192_n N_A1_c_236_n 0.0169052f $X=2.36 $Y=1.515 $X2=0 $Y2=0
cc_164 N_A2_c_193_n N_A1_c_236_n 3.89752e-19 $X=2.36 $Y=1.515 $X2=0 $Y2=0
cc_165 N_A2_c_197_n N_A1_c_236_n 0.00291709f $X=2.17 $Y=1.92 $X2=0 $Y2=0
cc_166 N_A2_M1001_g N_VPWR_c_268_n 0.00449364f $X=2.285 $Y=2.4 $X2=0 $Y2=0
cc_167 A2 N_VPWR_c_268_n 0.00684978f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_168 N_A2_M1001_g N_VPWR_c_262_n 0.00737192f $X=2.285 $Y=2.4 $X2=0 $Y2=0
cc_169 A2 N_VPWR_c_262_n 0.00815361f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_170 A2 A_361_368# 0.0146718f $X=2.075 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_171 N_A2_c_197_n A_361_368# 9.2419e-19 $X=2.17 $Y=1.92 $X2=-0.19 $Y2=-0.245
cc_172 N_A2_M1007_g N_A_157_74#_c_345_n 0.00966073f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A2_M1007_g N_A_157_74#_c_346_n 0.0117984f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A2_c_192_n N_A_157_74#_c_346_n 0.0224209f $X=2.36 $Y=1.515 $X2=0 $Y2=0
cc_175 N_A2_c_193_n N_A_157_74#_c_346_n 0.0041539f $X=2.36 $Y=1.515 $X2=0 $Y2=0
cc_176 N_A2_M1007_g N_A_157_74#_c_347_n 6.28869e-19 $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A2_M1007_g N_A_157_74#_c_348_n 0.00155819f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A2_c_192_n N_A_157_74#_c_348_n 0.00818793f $X=2.36 $Y=1.515 $X2=0 $Y2=0
cc_179 N_A2_M1007_g N_VGND_c_396_n 0.00622602f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_180 N_A2_M1007_g N_VGND_c_399_n 0.00434272f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_181 N_A2_M1007_g N_VGND_c_402_n 0.0082141f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A1_M1004_g N_VPWR_c_266_n 0.00536186f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_183 N_A1_c_235_n N_VPWR_c_266_n 8.7069e-19 $X=2.975 $Y=1.515 $X2=0 $Y2=0
cc_184 N_A1_c_236_n N_VPWR_c_266_n 0.0208821f $X=2.975 $Y=1.515 $X2=0 $Y2=0
cc_185 N_A1_M1004_g N_VPWR_c_268_n 0.00553757f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_186 N_A1_M1004_g N_VPWR_c_262_n 0.0109354f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A1_M1000_g N_A_157_74#_c_345_n 6.28869e-19 $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_188 N_A1_M1000_g N_A_157_74#_c_346_n 0.0153462f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A1_c_235_n N_A_157_74#_c_346_n 0.00177798f $X=2.975 $Y=1.515 $X2=0
+ $Y2=0
cc_190 N_A1_c_236_n N_A_157_74#_c_346_n 0.0344691f $X=2.975 $Y=1.515 $X2=0 $Y2=0
cc_191 N_A1_M1000_g N_A_157_74#_c_347_n 0.0103339f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A1_M1000_g N_VGND_c_396_n 0.00622602f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_193 N_A1_M1000_g N_VGND_c_401_n 0.00434272f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A1_M1000_g N_VGND_c_402_n 0.00825053f $X=2.84 $Y=0.74 $X2=0 $Y2=0
cc_195 N_VPWR_c_267_n N_Y_c_301_n 0.0141382f $X=0.495 $Y=2.815 $X2=0 $Y2=0
cc_196 N_VPWR_c_268_n N_Y_c_301_n 0.014549f $X=2.995 $Y=3.33 $X2=0 $Y2=0
cc_197 N_VPWR_c_262_n N_Y_c_301_n 0.0119743f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_198 N_VPWR_c_263_n N_Y_c_299_n 0.0236074f $X=0.455 $Y=1.985 $X2=0 $Y2=0
cc_199 N_Y_c_300_n N_A_157_74#_c_342_n 0.0505664f $X=0.495 $Y=0.515 $X2=0 $Y2=0
cc_200 N_Y_c_297_n N_A_157_74#_c_344_n 0.0129299f $X=0.69 $Y=1.35 $X2=0 $Y2=0
cc_201 N_Y_c_300_n N_VGND_c_397_n 0.0284523f $X=0.495 $Y=0.515 $X2=0 $Y2=0
cc_202 N_Y_c_300_n N_VGND_c_402_n 0.0232443f $X=0.495 $Y=0.515 $X2=0 $Y2=0
cc_203 N_A_157_74#_c_343_n N_VGND_M1008_d 0.00378075f $X=1.89 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_204 N_A_157_74#_c_346_n N_VGND_M1007_d 0.00358162f $X=2.89 $Y=1.095 $X2=0
+ $Y2=0
cc_205 N_A_157_74#_c_342_n N_VGND_c_395_n 0.0184106f $X=1.04 $Y=0.515 $X2=0
+ $Y2=0
cc_206 N_A_157_74#_c_343_n N_VGND_c_395_n 0.0257907f $X=1.89 $Y=1.095 $X2=0
+ $Y2=0
cc_207 N_A_157_74#_c_345_n N_VGND_c_395_n 0.0356652f $X=2.055 $Y=0.515 $X2=0
+ $Y2=0
cc_208 N_A_157_74#_c_345_n N_VGND_c_396_n 0.0191765f $X=2.055 $Y=0.515 $X2=0
+ $Y2=0
cc_209 N_A_157_74#_c_346_n N_VGND_c_396_n 0.0248957f $X=2.89 $Y=1.095 $X2=0
+ $Y2=0
cc_210 N_A_157_74#_c_347_n N_VGND_c_396_n 0.0191765f $X=3.055 $Y=0.515 $X2=0
+ $Y2=0
cc_211 N_A_157_74#_c_342_n N_VGND_c_397_n 0.0109942f $X=1.04 $Y=0.515 $X2=0
+ $Y2=0
cc_212 N_A_157_74#_c_345_n N_VGND_c_399_n 0.0144922f $X=2.055 $Y=0.515 $X2=0
+ $Y2=0
cc_213 N_A_157_74#_c_347_n N_VGND_c_401_n 0.0145639f $X=3.055 $Y=0.515 $X2=0
+ $Y2=0
cc_214 N_A_157_74#_c_342_n N_VGND_c_402_n 0.00904371f $X=1.04 $Y=0.515 $X2=0
+ $Y2=0
cc_215 N_A_157_74#_c_345_n N_VGND_c_402_n 0.0118826f $X=2.055 $Y=0.515 $X2=0
+ $Y2=0
cc_216 N_A_157_74#_c_347_n N_VGND_c_402_n 0.0119984f $X=3.055 $Y=0.515 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__o2bb2ai_4.spice
* Created: Wed Sep  2 12:24:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o2bb2ai_4.pex.spice"
.subckt sky130_fd_sc_ms__o2bb2ai_4  VNB VPB A1_N A2_N B2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1012 N_A_27_74#_M1012_d N_A1_N_M1012_g N_VGND_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1032 N_A_27_74#_M1032_d N_A1_N_M1032_g N_VGND_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1073 AS=0.1036 PD=1.03 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1033 N_A_27_74#_M1032_d N_A1_N_M1033_g N_VGND_M1033_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1073 AS=0.1036 PD=1.03 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1034 N_A_27_74#_M1034_d N_A1_N_M1034_g N_VGND_M1033_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1008 N_A_27_74#_M1034_d N_A2_N_M1008_g N_A_117_368#_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.9 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1017 N_A_27_74#_M1017_d N_A2_N_M1017_g N_A_117_368#_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.13875 AS=0.1036 PD=1.115 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1022 N_A_27_74#_M1017_d N_A2_N_M1022_g N_A_117_368#_M1022_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.13875 AS=0.12025 PD=1.115 PS=1.065 NRD=4.044 NRS=7.296 M=1
+ R=4.93333 SA=75002.9 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1039 N_A_27_74#_M1039_d N_A2_N_M1039_g N_A_117_368#_M1022_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.12025 PD=2.05 PS=1.065 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.4 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_A_857_74#_M1009_d N_A_117_368#_M1009_g N_Y_M1009_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75005.1 A=0.111 P=1.78 MULT=1
MM1018 N_A_857_74#_M1018_d N_A_117_368#_M1018_g N_Y_M1009_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75004.7 A=0.111 P=1.78 MULT=1
MM1023 N_A_857_74#_M1018_d N_A_117_368#_M1023_g N_Y_M1023_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75004.3 A=0.111 P=1.78 MULT=1
MM1029 N_A_857_74#_M1029_d N_A_117_368#_M1029_g N_Y_M1023_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75003.9 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_B2_M1002_g N_A_857_74#_M1029_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75003.4 A=0.111 P=1.78 MULT=1
MM1024 N_VGND_M1002_d N_B2_M1024_g N_A_857_74#_M1024_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.4
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1025 N_VGND_M1025_d N_B2_M1025_g N_A_857_74#_M1024_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.9
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1038 N_VGND_M1025_d N_B2_M1038_g N_A_857_74#_M1038_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75003.4
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1006 N_A_857_74#_M1038_s N_B1_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.8
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1013 N_A_857_74#_M1013_d N_B1_M1013_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.2
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1016 N_A_857_74#_M1013_d N_B1_M1016_g N_VGND_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75004.6
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1035 N_A_857_74#_M1035_d N_B1_M1035_g N_VGND_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1026 N_A_117_368#_M1026_d N_A1_N_M1026_g N_VPWR_M1026_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3024 PD=1.39 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90005.1 A=0.2016 P=2.6 MULT=1
MM1027 N_A_117_368#_M1026_d N_A1_N_M1027_g N_VPWR_M1027_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90004.7 A=0.2016 P=2.6 MULT=1
MM1030 N_A_117_368#_M1030_d N_A1_N_M1030_g N_VPWR_M1027_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.1 SB=90004.2 A=0.2016 P=2.6 MULT=1
MM1036 N_A_117_368#_M1030_d N_A1_N_M1036_g N_VPWR_M1036_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.5 SB=90003.8 A=0.2016 P=2.6 MULT=1
MM1000 N_A_117_368#_M1000_d N_A2_N_M1000_g N_VPWR_M1036_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90003.3 A=0.2016 P=2.6 MULT=1
MM1003 N_A_117_368#_M1000_d N_A2_N_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90002.4 SB=90002.9 A=0.2016 P=2.6 MULT=1
MM1005 N_A_117_368#_M1005_d N_A2_N_M1005_g N_VPWR_M1003_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90002.9 SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1010 N_A_117_368#_M1005_d N_A2_N_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90003.3 SB=90002 A=0.2016 P=2.6 MULT=1
MM1014 N_Y_M1014_d N_A_117_368#_M1014_g N_VPWR_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.8
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1019 N_Y_M1014_d N_A_117_368#_M1019_g N_VPWR_M1019_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.2
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1021 N_Y_M1021_d N_A_117_368#_M1021_g N_VPWR_M1019_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.7
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1028 N_Y_M1021_d N_A_117_368#_M1028_g N_VPWR_M1028_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3024 PD=1.39 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222 SA=90005.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1001 N_Y_M1001_d N_B2_M1001_g N_A_1215_368#_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3024 PD=1.39 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003.3 A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1001_d N_B2_M1004_g N_A_1215_368#_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90002.9 A=0.2016 P=2.6 MULT=1
MM1031 N_Y_M1031_d N_B2_M1031_g N_A_1215_368#_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1037 N_Y_M1031_d N_B2_M1037_g N_A_1215_368#_M1037_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90002 A=0.2016 P=2.6 MULT=1
MM1007 N_VPWR_M1007_d N_B1_M1007_g N_A_1215_368#_M1037_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1011 N_VPWR_M1007_d N_B1_M1011_g N_A_1215_368#_M1011_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90002.4 SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1015 N_VPWR_M1015_d N_B1_M1015_g N_A_1215_368#_M1011_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90002.9 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1020 N_VPWR_M1015_d N_B1_M1020_g N_A_1215_368#_M1020_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3024 PD=1.39 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90003.3 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX40_noxref VNB VPB NWDIODE A=19.4556 P=24.64
c_94 VNB 0 1.74044e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__o2bb2ai_4.pxi.spice"
*
.ends
*
*

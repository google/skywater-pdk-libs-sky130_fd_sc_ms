* NGSPICE file created from sky130_fd_sc_ms__decap_4.ext - technology: sky130A

.subckt sky130_fd_sc_ms__decap_4 VGND VNB VPB VPWR
M1000 VPWR VGND VPWR VPB pshort w=1e+06u l=1e+06u
+  ad=5.6e+11p pd=5.12e+06u as=0p ps=0u
M1001 VGND VPWR VGND VNB nlowvt w=420000u l=1e+06u
+  ad=2.31e+11p pd=2.78e+06u as=0p ps=0u
.ends


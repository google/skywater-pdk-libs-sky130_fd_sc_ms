* NGSPICE file created from sky130_fd_sc_ms__and4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__and4b_1 A_N B C D VGND VNB VPB VPWR X
M1000 VGND D a_526_139# VNB nlowvt w=640000u l=150000u
+  ad=4.5645e+11p pd=3.97e+06u as=3.418e+11p ps=2.55e+06u
M1001 a_448_139# B a_353_124# VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=2.21125e+11p ps=2.08e+06u
M1002 a_229_424# a_27_74# VPWR VPB pshort w=840000u l=180000u
+  ad=5.628e+11p pd=4.7e+06u as=1.5316e+12p ps=9.08e+06u
M1003 a_353_124# a_27_74# a_229_424# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1004 VPWR A_N a_27_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1005 X a_229_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1006 VPWR B a_229_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A_N a_27_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1008 VPWR D a_229_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_229_424# C VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_229_424# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1011 a_526_139# C a_448_139# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__clkbuf_1.pex.spice
* Created: Wed Sep  2 12:00:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__CLKBUF_1%A 3 7 9 10 18
c35 7 0 1.37764e-19 $X=0.735 $Y=2.4
r36 16 18 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.66 $Y=1.465
+ $X2=0.735 $Y2=1.465
r37 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.66
+ $Y=1.465 $X2=0.66 $Y2=1.465
r38 13 16 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.465
+ $X2=0.66 $Y2=1.465
r39 10 17 1.4951 $w=4.78e-07 $l=6e-08 $layer=LI1_cond $X=0.72 $Y=1.54 $X2=0.66
+ $Y2=1.54
r40 9 17 10.4657 $w=4.78e-07 $l=4.2e-07 $layer=LI1_cond $X=0.24 $Y=1.54 $X2=0.66
+ $Y2=1.54
r41 5 18 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.735 $Y=1.63
+ $X2=0.735 $Y2=1.465
r42 5 7 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.735 $Y=1.63
+ $X2=0.735 $Y2=2.4
r43 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.465
r44 1 3 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__CLKBUF_1%A_27_74# 1 2 8 11 15 17 20 22 24 26 27 28
+ 30 31 33 38 39
r69 38 41 46.536 $w=4.35e-07 $l=1.65e-07 $layer=POLY_cond $X=1.282 $Y=1.125
+ $X2=1.282 $Y2=0.96
r70 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.23
+ $Y=1.125 $X2=1.23 $Y2=1.125
r71 33 39 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.09 $Y=1.95 $X2=1.09
+ $Y2=1.63
r72 31 39 9.49412 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=1.2 $Y=1.435
+ $X2=1.2 $Y2=1.63
r73 30 37 2.51472 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=1.13 $X2=1.2
+ $Y2=1.045
r74 30 31 9.0127 $w=3.88e-07 $l=3.05e-07 $layer=LI1_cond $X=1.2 $Y=1.13 $X2=1.2
+ $Y2=1.435
r75 29 35 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.675 $Y=2.035
+ $X2=0.51 $Y2=2.035
r76 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.005 $Y=2.035
+ $X2=1.09 $Y2=1.95
r77 28 29 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.005 $Y=2.035
+ $X2=0.675 $Y2=2.035
r78 26 37 5.76906 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.005 $Y=1.045
+ $X2=1.2 $Y2=1.045
r79 26 27 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.005 $Y=1.045
+ $X2=0.445 $Y2=1.045
r80 22 35 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.51 $Y=2.12 $X2=0.51
+ $Y2=2.035
r81 22 24 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.51 $Y=2.12
+ $X2=0.51 $Y2=2.815
r82 18 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.96
+ $X2=0.445 $Y2=1.045
r83 18 20 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=0.28 $Y=0.96
+ $X2=0.28 $Y2=0.58
r84 15 41 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=1.425 $Y=0.58
+ $X2=1.425 $Y2=0.96
r85 11 17 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.285 $Y=2.4
+ $X2=1.285 $Y2=1.63
r86 8 17 37.6912 $w=4.35e-07 $l=2.17e-07 $layer=POLY_cond $X=1.282 $Y=1.413
+ $X2=1.282 $Y2=1.63
r87 7 38 6.64828 $w=4.35e-07 $l=5.2e-08 $layer=POLY_cond $X=1.282 $Y=1.177
+ $X2=1.282 $Y2=1.125
r88 7 8 30.1729 $w=4.35e-07 $l=2.36e-07 $layer=POLY_cond $X=1.282 $Y=1.177
+ $X2=1.282 $Y2=1.413
r89 2 35 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.365
+ $Y=1.84 $X2=0.51 $Y2=2.115
r90 2 24 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.365
+ $Y=1.84 $X2=0.51 $Y2=2.815
r91 1 20 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__CLKBUF_1%VPWR 1 6 9 10 11 18 19
r22 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r23 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r24 11 19 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r25 11 15 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r26 9 14 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.845 $Y=3.33
+ $X2=0.72 $Y2=3.33
r27 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=3.33
+ $X2=1.01 $Y2=3.33
r28 8 18 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=1.175 $Y=3.33
+ $X2=1.68 $Y2=3.33
r29 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.175 $Y=3.33
+ $X2=1.01 $Y2=3.33
r30 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.01 $Y=3.245 $X2=1.01
+ $Y2=3.33
r31 4 6 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.01 $Y=3.245 $X2=1.01
+ $Y2=2.455
r32 1 6 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=0.825
+ $Y=1.84 $X2=1.01 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__CLKBUF_1%X 1 2 7 8 9 10 11 12 13 45 49
c24 45 0 1.37764e-19 $X=1.51 $Y=1.985
r25 45 46 7.01411 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=1.985
+ $X2=1.575 $Y2=1.82
r26 30 49 0.390026 $w=4.58e-07 $l=1.5e-08 $layer=LI1_cond $X=1.575 $Y=2.05
+ $X2=1.575 $Y2=2.035
r27 13 37 1.04007 $w=4.58e-07 $l=4e-08 $layer=LI1_cond $X=1.575 $Y=2.775
+ $X2=1.575 $Y2=2.815
r28 12 13 9.62063 $w=4.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.575 $Y=2.405
+ $X2=1.575 $Y2=2.775
r29 11 49 0.91006 $w=4.58e-07 $l=3.5e-08 $layer=LI1_cond $X=1.575 $Y=2 $X2=1.575
+ $Y2=2.035
r30 11 45 0.390026 $w=4.58e-07 $l=1.5e-08 $layer=LI1_cond $X=1.575 $Y=2
+ $X2=1.575 $Y2=1.985
r31 11 12 8.32055 $w=4.58e-07 $l=3.2e-07 $layer=LI1_cond $X=1.575 $Y=2.085
+ $X2=1.575 $Y2=2.405
r32 11 30 0.91006 $w=4.58e-07 $l=3.5e-08 $layer=LI1_cond $X=1.575 $Y=2.085
+ $X2=1.575 $Y2=2.05
r33 10 46 7.44286 $w=2.38e-07 $l=1.55e-07 $layer=LI1_cond $X=1.685 $Y=1.665
+ $X2=1.685 $Y2=1.82
r34 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.685 $Y=1.295
+ $X2=1.685 $Y2=1.665
r35 8 9 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.685 $Y=0.925
+ $X2=1.685 $Y2=1.295
r36 8 43 6.48249 $w=2.38e-07 $l=1.35e-07 $layer=LI1_cond $X=1.685 $Y=0.925
+ $X2=1.685 $Y2=0.79
r37 7 43 9.08452 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.64 $Y=0.555
+ $X2=1.64 $Y2=0.79
r38 2 45 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.375
+ $Y=1.84 $X2=1.51 $Y2=1.985
r39 2 37 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.375
+ $Y=1.84 $X2=1.51 $Y2=2.815
r40 1 7 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.64 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_MS__CLKBUF_1%VGND 1 4 13 14 19 25
r19 23 25 10.279 $w=7.63e-07 $l=1.05e-07 $layer=LI1_cond $X=1.2 $Y=0.297
+ $X2=1.305 $Y2=0.297
r20 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r21 21 23 0.938101 $w=7.63e-07 $l=6e-08 $layer=LI1_cond $X=1.14 $Y=0.297 $X2=1.2
+ $Y2=0.297
r22 17 21 6.5667 $w=7.63e-07 $l=4.2e-07 $layer=LI1_cond $X=0.72 $Y=0.297
+ $X2=1.14 $Y2=0.297
r23 17 19 10.279 $w=7.63e-07 $l=1.05e-07 $layer=LI1_cond $X=0.72 $Y=0.297
+ $X2=0.615 $Y2=0.297
r24 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r25 14 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r26 13 25 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=1.305
+ $Y2=0
r27 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r28 9 18 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r29 8 19 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=0.615
+ $Y2=0
r30 8 9 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r31 4 24 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r32 4 18 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r33 1 21 91 $w=1.7e-07 $l=6.38396e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=1.14 $Y2=0.515
.ends


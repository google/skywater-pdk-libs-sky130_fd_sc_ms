* File: sky130_fd_sc_ms__o2111ai_1.pex.spice
* Created: Fri Aug 28 17:51:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O2111AI_1%D1 3 7 8 11 13
c29 8 0 4.41642e-20 $X=0.72 $Y=1.295
r30 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.745 $Y=1.385
+ $X2=0.745 $Y2=1.55
r31 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.745 $Y=1.385
+ $X2=0.745 $Y2=1.22
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.745
+ $Y=1.385 $X2=0.745 $Y2=1.385
r33 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.745 $Y=1.295
+ $X2=0.745 $Y2=1.385
r34 7 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.835 $Y=0.74
+ $X2=0.835 $Y2=1.22
r35 3 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.82 $Y=2.4 $X2=0.82
+ $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_1%C1 3 6 8 9 10 15 17
c40 17 0 3.10838e-19 $X=1.285 $Y=1.22
r41 15 18 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.285 $Y=1.385
+ $X2=1.285 $Y2=1.55
r42 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.285 $Y=1.385
+ $X2=1.285 $Y2=1.22
r43 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.285
+ $Y=1.385 $X2=1.285 $Y2=1.385
r44 10 16 3.05058 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=1.255 $Y=1.295
+ $X2=1.255 $Y2=1.385
r45 9 10 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.255 $Y=0.925
+ $X2=1.255 $Y2=1.295
r46 8 9 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.255 $Y=0.555
+ $X2=1.255 $Y2=0.925
r47 6 18 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.27 $Y=2.4 $X2=1.27
+ $Y2=1.55
r48 3 17 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.225 $Y=0.74
+ $X2=1.225 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_1%B1 3 6 8 11 12 13
c33 13 0 3.90916e-20 $X=1.825 $Y=1.22
c34 12 0 2.68987e-19 $X=1.825 $Y=1.385
r35 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=1.385
+ $X2=1.825 $Y2=1.55
r36 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=1.385
+ $X2=1.825 $Y2=1.22
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.825
+ $Y=1.385 $X2=1.825 $Y2=1.385
r38 8 12 4.51633 $w=3.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=1.825 $Y2=1.365
r39 6 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.9 $Y=2.4 $X2=1.9
+ $Y2=1.55
r40 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.765 $Y=0.74
+ $X2=1.765 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_1%A2 3 6 8 11 13
c34 13 0 1.79793e-19 $X=2.365 $Y=1.22
c35 8 0 3.90916e-20 $X=2.64 $Y=1.295
r36 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.365 $Y=1.385
+ $X2=2.365 $Y2=1.55
r37 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.365 $Y=1.385
+ $X2=2.365 $Y2=1.22
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.365
+ $Y=1.385 $X2=2.365 $Y2=1.385
r39 8 12 8.56545 $w=3.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.64 $Y=1.365
+ $X2=2.365 $Y2=1.365
r40 6 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.375 $Y=2.4
+ $X2=2.375 $Y2=1.55
r41 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.275 $Y=0.74
+ $X2=2.275 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_1%A1 3 5 7 8 14
c26 8 0 2.40942e-20 $X=3.12 $Y=1.295
r27 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.385 $X2=3.09 $Y2=1.385
r28 12 14 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=2.865 $Y=1.385
+ $X2=3.09 $Y2=1.385
r29 10 12 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=2.83 $Y=1.385
+ $X2=2.865 $Y2=1.385
r30 8 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.09 $Y=1.295 $X2=3.09
+ $Y2=1.385
r31 5 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.22
+ $X2=2.865 $Y2=1.385
r32 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.865 $Y=1.22 $X2=2.865
+ $Y2=0.74
r33 1 10 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.83 $Y=1.55
+ $X2=2.83 $Y2=1.385
r34 1 3 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=2.83 $Y=1.55 $X2=2.83
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_1%VPWR 1 2 3 12 18 22 24 29 30 31 37 41 47
+ 51
r42 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 45 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 42 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=1.65 $Y2=3.33
r46 42 44 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 41 50 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=2.89 $Y=3.33
+ $X2=3.125 $Y2=3.33
r48 41 44 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.89 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r50 37 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.65 $Y2=3.33
r51 37 39 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 35 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r54 31 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r55 31 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 31 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 29 34 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=0.38 $Y=3.33
+ $X2=0.24 $Y2=3.33
r58 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.38 $Y=3.33
+ $X2=0.545 $Y2=3.33
r59 28 39 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=0.71 $Y=3.33 $X2=1.2
+ $Y2=3.33
r60 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.71 $Y=3.33
+ $X2=0.545 $Y2=3.33
r61 24 27 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=3.055 $Y=1.985
+ $X2=3.055 $Y2=2.815
r62 22 50 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=3.055 $Y=3.245
+ $X2=3.125 $Y2=3.33
r63 22 27 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.055 $Y=3.245
+ $X2=3.055 $Y2=2.815
r64 18 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.65 $Y=2.145
+ $X2=1.65 $Y2=2.825
r65 16 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.65 $Y=3.245
+ $X2=1.65 $Y2=3.33
r66 16 21 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.65 $Y=3.245
+ $X2=1.65 $Y2=2.825
r67 12 15 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.545 $Y=2.145
+ $X2=0.545 $Y2=2.825
r68 10 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.545 $Y=3.245
+ $X2=0.545 $Y2=3.33
r69 10 15 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=0.545 $Y=3.245
+ $X2=0.545 $Y2=2.825
r70 3 27 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.92
+ $Y=1.84 $X2=3.055 $Y2=2.815
r71 3 24 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.92
+ $Y=1.84 $X2=3.055 $Y2=1.985
r72 2 21 400 $w=1.7e-07 $l=1.12066e-06 $layer=licon1_PDIFF $count=1 $X=1.36
+ $Y=1.84 $X2=1.65 $Y2=2.825
r73 2 18 400 $w=1.7e-07 $l=4.25999e-07 $layer=licon1_PDIFF $count=1 $X=1.36
+ $Y=1.84 $X2=1.65 $Y2=2.145
r74 1 15 400 $w=1.7e-07 $l=1.05501e-06 $layer=licon1_PDIFF $count=1 $X=0.4
+ $Y=1.84 $X2=0.545 $Y2=2.825
r75 1 12 400 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_PDIFF $count=1 $X=0.4
+ $Y=1.84 $X2=0.545 $Y2=2.145
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_1%Y 1 2 3 11 12 13 14 18 25 28 29 30 31 36
r58 31 44 1.05972 $w=4.33e-07 $l=4e-08 $layer=LI1_cond $X=1.097 $Y=2.775
+ $X2=1.097 $Y2=2.815
r59 30 31 9.80239 $w=4.33e-07 $l=3.7e-07 $layer=LI1_cond $X=1.097 $Y=2.405
+ $X2=1.097 $Y2=2.775
r60 29 30 9.80239 $w=4.33e-07 $l=3.7e-07 $layer=LI1_cond $X=1.097 $Y=2.035
+ $X2=1.097 $Y2=2.405
r61 29 36 1.32465 $w=4.33e-07 $l=5e-08 $layer=LI1_cond $X=1.097 $Y=2.035
+ $X2=1.097 $Y2=1.985
r62 27 36 2.51683 $w=4.33e-07 $l=9.5e-08 $layer=LI1_cond $X=1.097 $Y=1.89
+ $X2=1.097 $Y2=1.985
r63 27 28 1.70358 $w=4.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.097 $Y=1.89
+ $X2=1.097 $Y2=1.805
r64 22 25 7.61141 $w=6.58e-07 $l=4.2e-07 $layer=LI1_cond $X=0.2 $Y=0.68 $X2=0.62
+ $Y2=0.68
r65 18 20 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.15 $Y=1.985
+ $X2=2.15 $Y2=2.815
r66 16 18 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.15 $Y=1.89
+ $X2=2.15 $Y2=1.985
r67 15 28 10.3577 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=1.315 $Y=1.805
+ $X2=1.097 $Y2=1.805
r68 14 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.985 $Y=1.805
+ $X2=2.15 $Y2=1.89
r69 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.985 $Y=1.805
+ $X2=1.315 $Y2=1.805
r70 12 28 10.3577 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=0.88 $Y=1.805
+ $X2=1.097 $Y2=1.805
r71 12 13 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=0.88 $Y=1.805
+ $X2=0.285 $Y2=1.805
r72 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.2 $Y=1.72
+ $X2=0.285 $Y2=1.805
r73 10 22 8.93547 $w=1.7e-07 $l=3.3e-07 $layer=LI1_cond $X=0.2 $Y=1.01 $X2=0.2
+ $Y2=0.68
r74 10 11 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.2 $Y=1.01 $X2=0.2
+ $Y2=1.72
r75 3 20 400 $w=1.7e-07 $l=1.05196e-06 $layer=licon1_PDIFF $count=1 $X=1.99
+ $Y=1.84 $X2=2.15 $Y2=2.815
r76 3 18 400 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=1.99
+ $Y=1.84 $X2=2.15 $Y2=1.985
r77 2 44 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=1.84 $X2=1.045 $Y2=2.815
r78 2 36 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=1.84 $X2=1.045 $Y2=1.985
r79 1 25 45.5 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_NDIFF $count=4 $X=0.135
+ $Y=0.37 $X2=0.62 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_1%A_368_74# 1 2 7 9 11 15
c28 7 0 1.53386e-19 $X=1.99 $Y=0.84
r29 13 15 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.08 $Y=0.84
+ $X2=3.08 $Y2=0.515
r30 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.155 $Y=0.925
+ $X2=1.99 $Y2=0.925
r31 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.915 $Y=0.925
+ $X2=3.08 $Y2=0.84
r32 11 12 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.915 $Y=0.925
+ $X2=2.155 $Y2=0.925
r33 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=0.84 $X2=1.99
+ $Y2=0.925
r34 7 9 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.99 $Y=0.84 $X2=1.99
+ $Y2=0.515
r35 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.94
+ $Y=0.37 $X2=3.08 $Y2=0.515
r36 1 18 182 $w=1.7e-07 $l=6.2552e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.37 $X2=1.99 $Y2=0.925
r37 1 9 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.37 $X2=1.99 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_1%VGND 1 6 8 10 20 21 24
r31 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r32 21 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r33 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r34 18 24 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.535
+ $Y2=0
r35 18 20 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=3.12
+ $Y2=0
r36 17 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r37 16 17 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r38 12 16 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r39 12 13 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r40 10 24 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.325 $Y=0 $X2=2.535
+ $Y2=0
r41 10 16 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=0 $X2=2.16
+ $Y2=0
r42 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r43 8 13 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r44 4 24 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.535 $Y=0.085
+ $X2=2.535 $Y2=0
r45 4 6 11.7988 $w=4.18e-07 $l=4.3e-07 $layer=LI1_cond $X=2.535 $Y=0.085
+ $X2=2.535 $Y2=0.515
r46 1 6 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=2.35
+ $Y=0.37 $X2=2.535 $Y2=0.515
.ends


* NGSPICE file created from sky130_fd_sc_ms__clkdlyinv3sd1_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__clkdlyinv3sd1_1 A VGND VNB VPB VPWR Y
M1000 Y a_288_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=1.0312e+12p ps=6.42e+06u
M1001 a_288_74# a_28_74# VPWR VPB pshort w=1e+06u l=150000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1002 VPWR A a_28_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=2.968e+11p ps=2.77e+06u
M1003 VGND A a_28_74# VNB nlowvt w=420000u l=150000u
+  ad=4.2e+11p pd=3.68e+06u as=1.113e+11p ps=1.37e+06u
M1004 a_288_74# a_28_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1005 Y a_288_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
.ends


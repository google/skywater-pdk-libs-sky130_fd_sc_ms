* File: sky130_fd_sc_ms__bufbuf_16.pex.spice
* Created: Wed Sep  2 11:59:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__BUFBUF_16%A 3 7 9 13 16
c34 3 0 5.52684e-20 $X=0.505 $Y=2.4
r35 15 16 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=0.505 $Y=1.465
+ $X2=0.51 $Y2=1.465
r36 12 15 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.34 $Y=1.465
+ $X2=0.505 $Y2=1.465
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.34
+ $Y=1.465 $X2=0.34 $Y2=1.465
r38 9 13 6.06549 $w=3.78e-07 $l=2e-07 $layer=LI1_cond $X=0.315 $Y=1.665
+ $X2=0.315 $Y2=1.465
r39 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.3 $X2=0.51
+ $Y2=1.465
r40 5 7 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.51 $Y=1.3 $X2=0.51
+ $Y2=0.74
r41 1 15 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=1.465
r42 1 3 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__BUFBUF_16%A_27_368# 1 2 9 13 17 21 25 29 31 33 37 39
+ 40 41 44 46 52 57 66
c111 9 0 1.78628e-19 $X=0.94 $Y=0.74
r112 65 66 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=1.805 $Y=1.465
+ $X2=1.855 $Y2=1.465
r113 62 63 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=1.37 $Y=1.465
+ $X2=1.405 $Y2=1.465
r114 58 60 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.94 $Y=1.465
+ $X2=0.955 $Y2=1.465
r115 53 65 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=1.71 $Y=1.465
+ $X2=1.805 $Y2=1.465
r116 53 63 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=1.71 $Y=1.465
+ $X2=1.405 $Y2=1.465
r117 52 53 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.465 $X2=1.71 $Y2=1.465
r118 50 62 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.03 $Y=1.465
+ $X2=1.37 $Y2=1.465
r119 50 60 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.03 $Y=1.465
+ $X2=0.955 $Y2=1.465
r120 49 52 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.03 $Y=1.465
+ $X2=1.71 $Y2=1.465
r121 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.03
+ $Y=1.465 $X2=1.03 $Y2=1.465
r122 47 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.845 $Y=1.465
+ $X2=0.76 $Y2=1.465
r123 47 49 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.845 $Y=1.465
+ $X2=1.03 $Y2=1.465
r124 45 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.76 $Y=1.63
+ $X2=0.76 $Y2=1.465
r125 45 46 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.76 $Y=1.63
+ $X2=0.76 $Y2=1.95
r126 44 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.76 $Y=1.3
+ $X2=0.76 $Y2=1.465
r127 43 44 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.76 $Y=1.13
+ $X2=0.76 $Y2=1.3
r128 42 56 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.035
+ $X2=0.28 $Y2=2.035
r129 41 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.675 $Y=2.035
+ $X2=0.76 $Y2=1.95
r130 41 42 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.675 $Y=2.035
+ $X2=0.445 $Y2=2.035
r131 39 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.675 $Y=1.045
+ $X2=0.76 $Y2=1.13
r132 39 40 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.675 $Y=1.045
+ $X2=0.38 $Y2=1.045
r133 35 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.255 $Y=0.96
+ $X2=0.38 $Y2=1.045
r134 35 37 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.255 $Y=0.96
+ $X2=0.255 $Y2=0.515
r135 31 56 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.12 $X2=0.28
+ $Y2=2.035
r136 31 33 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.28 $Y=2.12
+ $X2=0.28 $Y2=2.815
r137 27 66 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.63
+ $X2=1.855 $Y2=1.465
r138 27 29 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.855 $Y=1.63
+ $X2=1.855 $Y2=2.4
r139 23 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.805 $Y=1.3
+ $X2=1.805 $Y2=1.465
r140 23 25 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.805 $Y=1.3
+ $X2=1.805 $Y2=0.74
r141 19 63 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.63
+ $X2=1.405 $Y2=1.465
r142 19 21 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.405 $Y=1.63
+ $X2=1.405 $Y2=2.4
r143 15 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.37 $Y=1.3
+ $X2=1.37 $Y2=1.465
r144 15 17 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.37 $Y=1.3
+ $X2=1.37 $Y2=0.74
r145 11 60 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.63
+ $X2=0.955 $Y2=1.465
r146 11 13 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.955 $Y=1.63
+ $X2=0.955 $Y2=2.4
r147 7 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.94 $Y=1.3
+ $X2=0.94 $Y2=1.465
r148 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.94 $Y=1.3 $X2=0.94
+ $Y2=0.74
r149 2 56 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
r150 2 33 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r151 1 37 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.37 $X2=0.295 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__BUFBUF_16%A_203_74# 1 2 3 4 15 19 23 27 31 35 39 43
+ 47 51 55 59 63 69 71 72 73 74 77 81 86 88 94 97 98 99 114
c196 74 0 5.52684e-20 $X=1.345 $Y=1.885
c197 72 0 1.78628e-19 $X=1.24 $Y=1.045
c198 55 0 6.44981e-20 $X=5.14 $Y=2.4
r199 113 114 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.14 $Y=1.485
+ $X2=5.155 $Y2=1.485
r200 112 113 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=4.725 $Y=1.485
+ $X2=5.14 $Y2=1.485
r201 111 112 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=4.69 $Y=1.485
+ $X2=4.725 $Y2=1.485
r202 108 109 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=4.225 $Y=1.485
+ $X2=4.23 $Y2=1.485
r203 107 108 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.795 $Y=1.485
+ $X2=4.225 $Y2=1.485
r204 106 107 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.78 $Y=1.485
+ $X2=3.795 $Y2=1.485
r205 105 106 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=3.33 $Y=1.485
+ $X2=3.78 $Y2=1.485
r206 104 105 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=3.295 $Y=1.485
+ $X2=3.33 $Y2=1.485
r207 100 102 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.865 $Y=1.485
+ $X2=2.88 $Y2=1.485
r208 95 111 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=4.315 $Y=1.485
+ $X2=4.69 $Y2=1.485
r209 95 109 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=4.315 $Y=1.485
+ $X2=4.23 $Y2=1.485
r210 94 95 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.315
+ $Y=1.485 $X2=4.315 $Y2=1.485
r211 92 104 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.955 $Y=1.485
+ $X2=3.295 $Y2=1.485
r212 92 102 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.955 $Y=1.485
+ $X2=2.88 $Y2=1.485
r213 91 94 47.4946 $w=3.28e-07 $l=1.36e-06 $layer=LI1_cond $X=2.955 $Y=1.485
+ $X2=4.315 $Y2=1.485
r214 91 92 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.955
+ $Y=1.485 $X2=2.955 $Y2=1.485
r215 89 99 0.63164 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=2.245 $Y=1.485
+ $X2=2.145 $Y2=1.485
r216 89 91 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.245 $Y=1.485
+ $X2=2.955 $Y2=1.485
r217 88 98 3.52026 $w=2.65e-07 $l=1.12916e-07 $layer=LI1_cond $X=2.145 $Y=1.8
+ $X2=2.08 $Y2=1.885
r218 87 99 8.10876 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=1.65
+ $X2=2.145 $Y2=1.485
r219 87 88 8.31818 $w=1.98e-07 $l=1.5e-07 $layer=LI1_cond $X=2.145 $Y=1.65
+ $X2=2.145 $Y2=1.8
r220 86 99 8.10876 $w=1.85e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.13 $Y=1.32
+ $X2=2.145 $Y2=1.485
r221 85 97 3.52026 $w=2.65e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.13 $Y=1.13
+ $X2=2.035 $Y2=1.045
r222 85 86 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.13 $Y=1.13
+ $X2=2.13 $Y2=1.32
r223 81 83 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.08 $Y=1.985
+ $X2=2.08 $Y2=2.815
r224 79 98 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=1.97
+ $X2=2.08 $Y2=1.885
r225 79 81 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.08 $Y=1.97
+ $X2=2.08 $Y2=1.985
r226 75 97 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.035 $Y=0.96
+ $X2=2.035 $Y2=1.045
r227 75 77 14.2455 $w=3.58e-07 $l=4.45e-07 $layer=LI1_cond $X=2.035 $Y=0.96
+ $X2=2.035 $Y2=0.515
r228 73 98 2.98021 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.915 $Y=1.885
+ $X2=2.08 $Y2=1.885
r229 73 74 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.915 $Y=1.885
+ $X2=1.345 $Y2=1.885
r230 71 97 2.98021 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.855 $Y=1.045
+ $X2=2.035 $Y2=1.045
r231 71 72 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.855 $Y=1.045
+ $X2=1.24 $Y2=1.045
r232 67 72 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.155 $Y=0.96
+ $X2=1.24 $Y2=1.045
r233 67 69 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.155 $Y=0.96
+ $X2=1.155 $Y2=0.515
r234 63 65 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.18 $Y=1.985
+ $X2=1.18 $Y2=2.815
r235 61 74 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.18 $Y=1.97
+ $X2=1.345 $Y2=1.885
r236 61 63 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.18 $Y=1.97
+ $X2=1.18 $Y2=1.985
r237 57 114 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.155 $Y=1.32
+ $X2=5.155 $Y2=1.485
r238 57 59 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.155 $Y=1.32
+ $X2=5.155 $Y2=0.74
r239 53 113 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.14 $Y=1.65
+ $X2=5.14 $Y2=1.485
r240 53 55 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=5.14 $Y=1.65
+ $X2=5.14 $Y2=2.4
r241 49 112 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.725 $Y=1.32
+ $X2=4.725 $Y2=1.485
r242 49 51 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.725 $Y=1.32
+ $X2=4.725 $Y2=0.74
r243 45 111 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.69 $Y=1.65
+ $X2=4.69 $Y2=1.485
r244 45 47 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=4.69 $Y=1.65
+ $X2=4.69 $Y2=2.4
r245 41 108 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.225 $Y=1.32
+ $X2=4.225 $Y2=1.485
r246 41 43 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.225 $Y=1.32
+ $X2=4.225 $Y2=0.74
r247 37 109 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.23 $Y=1.65
+ $X2=4.23 $Y2=1.485
r248 37 39 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=4.23 $Y=1.65
+ $X2=4.23 $Y2=2.4
r249 33 107 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.795 $Y=1.32
+ $X2=3.795 $Y2=1.485
r250 33 35 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.795 $Y=1.32
+ $X2=3.795 $Y2=0.74
r251 29 106 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.78 $Y=1.65
+ $X2=3.78 $Y2=1.485
r252 29 31 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=3.78 $Y=1.65
+ $X2=3.78 $Y2=2.4
r253 25 105 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.33 $Y=1.65
+ $X2=3.33 $Y2=1.485
r254 25 27 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=3.33 $Y=1.65
+ $X2=3.33 $Y2=2.4
r255 21 104 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.295 $Y=1.32
+ $X2=3.295 $Y2=1.485
r256 21 23 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.295 $Y=1.32
+ $X2=3.295 $Y2=0.74
r257 17 102 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.88 $Y=1.65
+ $X2=2.88 $Y2=1.485
r258 17 19 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=2.88 $Y=1.65
+ $X2=2.88 $Y2=2.4
r259 13 100 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.32
+ $X2=2.865 $Y2=1.485
r260 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.865 $Y=1.32
+ $X2=2.865 $Y2=0.74
r261 4 83 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.945
+ $Y=1.84 $X2=2.08 $Y2=2.815
r262 4 81 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.945
+ $Y=1.84 $X2=2.08 $Y2=1.985
r263 3 65 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.815
r264 3 63 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=1.985
r265 2 77 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.88
+ $Y=0.37 $X2=2.02 $Y2=0.515
r266 1 69 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.015
+ $Y=0.37 $X2=1.155 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__BUFBUF_16%A_588_74# 1 2 3 4 5 6 21 25 29 33 37 41 45
+ 49 53 57 61 65 69 73 77 81 85 89 93 97 101 105 109 113 117 121 125 129 133 137
+ 141 145 149 151 153 155 156 157 161 165 167 169 171 173 177 180 184 185 186
+ 210 220 227 234 241 248 255 262 266
c490 171 0 1.38532e-19 $X=4.915 $Y=1.99
c491 125 0 9.40629e-20 $X=11.455 $Y=0.74
c492 41 0 1.04236e-19 $X=6.55 $Y=2.4
r493 297 299 2.0766 $w=4.7e-07 $l=8e-08 $layer=LI1_cond $X=5.077 $Y=1.905
+ $X2=5.077 $Y2=1.985
r494 265 266 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=12.395 $Y=1.485
+ $X2=12.45 $Y2=1.485
r495 264 265 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=11.965 $Y=1.485
+ $X2=12.395 $Y2=1.485
r496 263 264 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=11.95 $Y=1.485
+ $X2=11.965 $Y2=1.485
r497 261 263 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=11.685 $Y=1.485
+ $X2=11.95 $Y2=1.485
r498 261 262 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.685
+ $Y=1.485 $X2=11.685 $Y2=1.485
r499 259 261 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=11.5 $Y=1.485
+ $X2=11.685 $Y2=1.485
r500 258 259 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=11.455 $Y=1.485
+ $X2=11.5 $Y2=1.485
r501 257 258 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=11.05 $Y=1.485
+ $X2=11.455 $Y2=1.485
r502 256 257 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=11.025 $Y=1.485
+ $X2=11.05 $Y2=1.485
r503 254 256 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=10.76 $Y=1.485
+ $X2=11.025 $Y2=1.485
r504 254 255 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.76
+ $Y=1.485 $X2=10.76 $Y2=1.485
r505 252 254 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=10.6 $Y=1.485
+ $X2=10.76 $Y2=1.485
r506 251 252 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=10.525 $Y=1.485
+ $X2=10.6 $Y2=1.485
r507 250 251 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=10.15 $Y=1.485
+ $X2=10.525 $Y2=1.485
r508 249 250 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=10.095 $Y=1.485
+ $X2=10.15 $Y2=1.485
r509 247 249 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=9.815 $Y=1.485
+ $X2=10.095 $Y2=1.485
r510 247 248 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.815
+ $Y=1.485 $X2=9.815 $Y2=1.485
r511 245 247 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=9.7 $Y=1.485
+ $X2=9.815 $Y2=1.485
r512 244 245 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=9.595 $Y=1.485
+ $X2=9.7 $Y2=1.485
r513 243 244 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=9.25 $Y=1.485
+ $X2=9.595 $Y2=1.485
r514 242 243 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=9.165 $Y=1.485
+ $X2=9.25 $Y2=1.485
r515 240 242 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=8.905 $Y=1.485
+ $X2=9.165 $Y2=1.485
r516 240 241 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.905
+ $Y=1.485 $X2=8.905 $Y2=1.485
r517 238 240 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=8.8 $Y=1.485
+ $X2=8.905 $Y2=1.485
r518 237 238 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=8.665 $Y=1.485
+ $X2=8.8 $Y2=1.485
r519 236 237 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=8.35 $Y=1.485
+ $X2=8.665 $Y2=1.485
r520 235 236 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=8.235 $Y=1.485
+ $X2=8.35 $Y2=1.485
r521 233 235 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=7.985 $Y=1.485
+ $X2=8.235 $Y2=1.485
r522 233 234 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.985
+ $Y=1.485 $X2=7.985 $Y2=1.485
r523 231 233 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=7.9 $Y=1.485
+ $X2=7.985 $Y2=1.485
r524 230 231 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.735 $Y=1.485
+ $X2=7.9 $Y2=1.485
r525 229 230 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=7.45 $Y=1.485
+ $X2=7.735 $Y2=1.485
r526 228 229 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=7.305 $Y=1.485
+ $X2=7.45 $Y2=1.485
r527 226 228 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=7.085 $Y=1.485
+ $X2=7.305 $Y2=1.485
r528 226 227 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.085
+ $Y=1.485 $X2=7.085 $Y2=1.485
r529 224 226 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=7 $Y=1.485
+ $X2=7.085 $Y2=1.485
r530 223 224 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=6.875 $Y=1.485
+ $X2=7 $Y2=1.485
r531 222 223 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=6.55 $Y=1.485
+ $X2=6.875 $Y2=1.485
r532 221 222 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=6.445 $Y=1.485
+ $X2=6.55 $Y2=1.485
r533 219 221 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=6.21 $Y=1.485
+ $X2=6.445 $Y2=1.485
r534 219 220 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.21
+ $Y=1.485 $X2=6.21 $Y2=1.485
r535 217 219 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=6.05 $Y=1.485
+ $X2=6.21 $Y2=1.485
r536 216 217 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=6.015 $Y=1.485
+ $X2=6.05 $Y2=1.485
r537 215 216 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=5.6 $Y=1.485
+ $X2=6.015 $Y2=1.485
r538 213 215 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.585 $Y=1.485
+ $X2=5.6 $Y2=1.485
r539 211 262 5.25164 $w=3.93e-07 $l=1.8e-07 $layer=LI1_cond $X=11.692 $Y=1.665
+ $X2=11.692 $Y2=1.485
r540 210 211 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.685 $Y=1.665
+ $X2=11.685 $Y2=1.665
r541 208 255 5.53173 $w=3.73e-07 $l=1.8e-07 $layer=LI1_cond $X=10.752 $Y=1.665
+ $X2=10.752 $Y2=1.485
r542 207 210 0.593484 $w=2.3e-07 $l=9.25e-07 $layer=MET1_cond $X=10.76 $Y=1.665
+ $X2=11.685 $Y2=1.665
r543 207 208 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.76 $Y=1.665
+ $X2=10.76 $Y2=1.665
r544 205 248 6.38276 $w=3.23e-07 $l=1.8e-07 $layer=LI1_cond $X=9.812 $Y=1.665
+ $X2=9.812 $Y2=1.485
r545 204 207 0.606316 $w=2.3e-07 $l=9.45e-07 $layer=MET1_cond $X=9.815 $Y=1.665
+ $X2=10.76 $Y2=1.665
r546 204 205 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.815 $Y=1.665
+ $X2=9.815 $Y2=1.665
r547 202 241 7.03186 $w=2.93e-07 $l=1.8e-07 $layer=LI1_cond $X=8.897 $Y=1.665
+ $X2=8.897 $Y2=1.485
r548 201 204 0.58386 $w=2.3e-07 $l=9.1e-07 $layer=MET1_cond $X=8.905 $Y=1.665
+ $X2=9.815 $Y2=1.665
r549 201 202 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.905 $Y=1.665
+ $X2=8.905 $Y2=1.665
r550 199 234 7.82791 $w=2.63e-07 $l=1.8e-07 $layer=LI1_cond $X=7.982 $Y=1.665
+ $X2=7.982 $Y2=1.485
r551 198 201 0.590276 $w=2.3e-07 $l=9.2e-07 $layer=MET1_cond $X=7.985 $Y=1.665
+ $X2=8.905 $Y2=1.665
r552 198 199 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.985 $Y=1.665
+ $X2=7.985 $Y2=1.665
r553 196 227 7.82791 $w=2.63e-07 $l=1.8e-07 $layer=LI1_cond $X=7.082 $Y=1.665
+ $X2=7.082 $Y2=1.485
r554 195 198 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=7.085 $Y=1.665
+ $X2=7.985 $Y2=1.665
r555 195 196 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.085 $Y=1.665
+ $X2=7.085 $Y2=1.665
r556 193 220 6.6916 $w=3.08e-07 $l=1.8e-07 $layer=LI1_cond $X=6.21 $Y=1.665
+ $X2=6.21 $Y2=1.485
r557 192 195 0.561404 $w=2.3e-07 $l=8.75e-07 $layer=MET1_cond $X=6.21 $Y=1.665
+ $X2=7.085 $Y2=1.665
r558 192 193 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=1.665
+ $X2=6.21 $Y2=1.665
r559 189 297 6.22979 $w=4.7e-07 $l=2.4e-07 $layer=LI1_cond $X=5.077 $Y=1.665
+ $X2=5.077 $Y2=1.905
r560 188 192 0.606316 $w=2.3e-07 $l=9.45e-07 $layer=MET1_cond $X=5.265 $Y=1.665
+ $X2=6.21 $Y2=1.665
r561 188 189 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.265 $Y=1.665
+ $X2=5.265 $Y2=1.665
r562 180 189 11.3723 $w=4.7e-07 $l=3.92702e-07 $layer=LI1_cond $X=4.975 $Y=1.32
+ $X2=5.077 $Y2=1.665
r563 179 186 3.64284 $w=2.55e-07 $l=1.00995e-07 $layer=LI1_cond $X=4.975 $Y=1.15
+ $X2=4.94 $Y2=1.065
r564 179 180 7.5352 $w=2.58e-07 $l=1.7e-07 $layer=LI1_cond $X=4.975 $Y=1.15
+ $X2=4.975 $Y2=1.32
r565 175 186 3.64284 $w=2.55e-07 $l=1.03078e-07 $layer=LI1_cond $X=4.9 $Y=0.98
+ $X2=4.94 $Y2=1.065
r566 175 177 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=4.9 $Y=0.98
+ $X2=4.9 $Y2=0.515
r567 171 299 1.22671 $w=4.7e-07 $l=1.64481e-07 $layer=LI1_cond $X=4.915 $Y=1.99
+ $X2=5.077 $Y2=1.985
r568 171 173 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=4.915 $Y=1.99
+ $X2=4.915 $Y2=2.815
r569 170 184 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.17 $Y=1.905
+ $X2=4.005 $Y2=1.905
r570 169 297 6.76998 $w=1.7e-07 $l=3.27e-07 $layer=LI1_cond $X=4.75 $Y=1.905
+ $X2=5.077 $Y2=1.905
r571 169 170 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.75 $Y=1.905
+ $X2=4.17 $Y2=1.905
r572 168 185 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.095 $Y=1.065
+ $X2=3.97 $Y2=1.065
r573 167 186 2.83584 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.775 $Y=1.065
+ $X2=4.94 $Y2=1.065
r574 167 168 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.775 $Y=1.065
+ $X2=4.095 $Y2=1.065
r575 163 185 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.97 $Y=0.98
+ $X2=3.97 $Y2=1.065
r576 163 165 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=3.97 $Y=0.98
+ $X2=3.97 $Y2=0.515
r577 159 184 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.005 $Y=1.99
+ $X2=4.005 $Y2=1.905
r578 159 161 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=4.005 $Y=1.99
+ $X2=4.005 $Y2=2.815
r579 158 182 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.27 $Y=1.905
+ $X2=3.105 $Y2=1.905
r580 157 184 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.84 $Y=1.905
+ $X2=4.005 $Y2=1.905
r581 157 158 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.84 $Y=1.905
+ $X2=3.27 $Y2=1.905
r582 155 185 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.845 $Y=1.065
+ $X2=3.97 $Y2=1.065
r583 155 156 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.845 $Y=1.065
+ $X2=3.165 $Y2=1.065
r584 151 182 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.105 $Y=1.99
+ $X2=3.105 $Y2=1.905
r585 151 153 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=3.105 $Y=1.99
+ $X2=3.105 $Y2=2.815
r586 147 156 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.04 $Y=0.98
+ $X2=3.165 $Y2=1.065
r587 147 149 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=3.04 $Y=0.98
+ $X2=3.04 $Y2=0.515
r588 143 266 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=12.45 $Y=1.65
+ $X2=12.45 $Y2=1.485
r589 143 145 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=12.45 $Y=1.65
+ $X2=12.45 $Y2=2.4
r590 139 265 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.395 $Y=1.32
+ $X2=12.395 $Y2=1.485
r591 139 141 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=12.395 $Y=1.32
+ $X2=12.395 $Y2=0.74
r592 135 264 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.965 $Y=1.32
+ $X2=11.965 $Y2=1.485
r593 135 137 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=11.965 $Y=1.32
+ $X2=11.965 $Y2=0.74
r594 131 263 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=11.95 $Y=1.65
+ $X2=11.95 $Y2=1.485
r595 131 133 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=11.95 $Y=1.65
+ $X2=11.95 $Y2=2.4
r596 127 259 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=11.5 $Y=1.65
+ $X2=11.5 $Y2=1.485
r597 127 129 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=11.5 $Y=1.65
+ $X2=11.5 $Y2=2.4
r598 123 258 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.455 $Y=1.32
+ $X2=11.455 $Y2=1.485
r599 123 125 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=11.455 $Y=1.32
+ $X2=11.455 $Y2=0.74
r600 119 257 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=11.05 $Y=1.65
+ $X2=11.05 $Y2=1.485
r601 119 121 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=11.05 $Y=1.65
+ $X2=11.05 $Y2=2.4
r602 115 256 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.025 $Y=1.32
+ $X2=11.025 $Y2=1.485
r603 115 117 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=11.025 $Y=1.32
+ $X2=11.025 $Y2=0.74
r604 111 252 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.6 $Y=1.65
+ $X2=10.6 $Y2=1.485
r605 111 113 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=10.6 $Y=1.65
+ $X2=10.6 $Y2=2.4
r606 107 251 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.525 $Y=1.32
+ $X2=10.525 $Y2=1.485
r607 107 109 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=10.525 $Y=1.32
+ $X2=10.525 $Y2=0.74
r608 103 250 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.15 $Y=1.65
+ $X2=10.15 $Y2=1.485
r609 103 105 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=10.15 $Y=1.65
+ $X2=10.15 $Y2=2.4
r610 99 249 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.095 $Y=1.32
+ $X2=10.095 $Y2=1.485
r611 99 101 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=10.095 $Y=1.32
+ $X2=10.095 $Y2=0.74
r612 95 245 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.7 $Y=1.65
+ $X2=9.7 $Y2=1.485
r613 95 97 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=9.7 $Y=1.65 $X2=9.7
+ $Y2=2.4
r614 91 244 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.595 $Y=1.32
+ $X2=9.595 $Y2=1.485
r615 91 93 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=9.595 $Y=1.32
+ $X2=9.595 $Y2=0.74
r616 87 243 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.25 $Y=1.65
+ $X2=9.25 $Y2=1.485
r617 87 89 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=9.25 $Y=1.65
+ $X2=9.25 $Y2=2.4
r618 83 242 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.165 $Y=1.32
+ $X2=9.165 $Y2=1.485
r619 83 85 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=9.165 $Y=1.32
+ $X2=9.165 $Y2=0.74
r620 79 238 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.8 $Y=1.65
+ $X2=8.8 $Y2=1.485
r621 79 81 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=8.8 $Y=1.65 $X2=8.8
+ $Y2=2.4
r622 75 237 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.665 $Y=1.32
+ $X2=8.665 $Y2=1.485
r623 75 77 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.665 $Y=1.32
+ $X2=8.665 $Y2=0.74
r624 71 236 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.35 $Y=1.65
+ $X2=8.35 $Y2=1.485
r625 71 73 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=8.35 $Y=1.65
+ $X2=8.35 $Y2=2.4
r626 67 235 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.235 $Y=1.32
+ $X2=8.235 $Y2=1.485
r627 67 69 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.235 $Y=1.32
+ $X2=8.235 $Y2=0.74
r628 63 231 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.9 $Y=1.65
+ $X2=7.9 $Y2=1.485
r629 63 65 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=7.9 $Y=1.65 $X2=7.9
+ $Y2=2.4
r630 59 230 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.735 $Y=1.32
+ $X2=7.735 $Y2=1.485
r631 59 61 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.735 $Y=1.32
+ $X2=7.735 $Y2=0.74
r632 55 229 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.45 $Y=1.65
+ $X2=7.45 $Y2=1.485
r633 55 57 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=7.45 $Y=1.65
+ $X2=7.45 $Y2=2.4
r634 51 228 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.305 $Y=1.32
+ $X2=7.305 $Y2=1.485
r635 51 53 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.305 $Y=1.32
+ $X2=7.305 $Y2=0.74
r636 47 224 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7 $Y=1.65 $X2=7
+ $Y2=1.485
r637 47 49 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=7 $Y=1.65 $X2=7
+ $Y2=2.4
r638 43 223 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.875 $Y=1.32
+ $X2=6.875 $Y2=1.485
r639 43 45 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.875 $Y=1.32
+ $X2=6.875 $Y2=0.74
r640 39 222 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.55 $Y=1.65
+ $X2=6.55 $Y2=1.485
r641 39 41 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=6.55 $Y=1.65
+ $X2=6.55 $Y2=2.4
r642 35 221 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.445 $Y=1.32
+ $X2=6.445 $Y2=1.485
r643 35 37 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.445 $Y=1.32
+ $X2=6.445 $Y2=0.74
r644 31 217 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.05 $Y=1.65
+ $X2=6.05 $Y2=1.485
r645 31 33 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=6.05 $Y=1.65
+ $X2=6.05 $Y2=2.4
r646 27 216 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.015 $Y=1.32
+ $X2=6.015 $Y2=1.485
r647 27 29 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.015 $Y=1.32
+ $X2=6.015 $Y2=0.74
r648 23 215 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.6 $Y=1.65
+ $X2=5.6 $Y2=1.485
r649 23 25 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=5.6 $Y=1.65 $X2=5.6
+ $Y2=2.4
r650 19 213 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.585 $Y=1.32
+ $X2=5.585 $Y2=1.485
r651 19 21 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.585 $Y=1.32
+ $X2=5.585 $Y2=0.74
r652 6 299 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.78
+ $Y=1.84 $X2=4.915 $Y2=1.985
r653 6 173 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.78
+ $Y=1.84 $X2=4.915 $Y2=2.815
r654 5 184 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.87
+ $Y=1.84 $X2=4.005 $Y2=1.985
r655 5 161 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.87
+ $Y=1.84 $X2=4.005 $Y2=2.815
r656 4 182 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.97
+ $Y=1.84 $X2=3.105 $Y2=1.985
r657 4 153 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.97
+ $Y=1.84 $X2=3.105 $Y2=2.815
r658 3 177 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.8
+ $Y=0.37 $X2=4.94 $Y2=0.515
r659 2 165 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.87
+ $Y=0.37 $X2=4.01 $Y2=0.515
r660 1 149 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.94
+ $Y=0.37 $X2=3.08 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__BUFBUF_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 14 47
+ 51 55 61 65 69 75 79 83 89 93 97 101 105 111 115 117 122 123 125 126 128 129
+ 131 132 134 135 137 138 140 141 142 143 144 150 176 181 187 190 193 196 199
+ 203
r232 202 203 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r233 199 200 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r234 196 197 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r235 194 197 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.8 $Y2=3.33
r236 193 194 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r237 190 191 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r238 187 188 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r239 185 203 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r240 185 200 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r241 184 185 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r242 182 199 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.89 $Y=3.33
+ $X2=11.765 $Y2=3.33
r243 182 184 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=11.89 $Y=3.33
+ $X2=12.24 $Y2=3.33
r244 181 202 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=12.59 $Y=3.33
+ $X2=12.775 $Y2=3.33
r245 181 184 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=12.59 $Y=3.33
+ $X2=12.24 $Y2=3.33
r246 180 200 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r247 180 197 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r248 179 180 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r249 177 196 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.91 $Y=3.33
+ $X2=10.825 $Y2=3.33
r250 177 179 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=10.91 $Y=3.33
+ $X2=11.28 $Y2=3.33
r251 176 199 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.64 $Y=3.33
+ $X2=11.765 $Y2=3.33
r252 176 179 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=11.64 $Y=3.33
+ $X2=11.28 $Y2=3.33
r253 175 194 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.84 $Y2=3.33
r254 174 175 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r255 172 175 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r256 171 172 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r257 169 172 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r258 168 169 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r259 165 166 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r260 163 166 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6 $Y2=3.33
r261 162 163 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r262 160 163 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r263 159 160 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r264 157 160 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r265 157 191 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r266 156 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r267 154 190 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.74 $Y=3.33
+ $X2=2.615 $Y2=3.33
r268 154 156 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.74 $Y=3.33
+ $X2=3.12 $Y2=3.33
r269 153 191 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r270 152 153 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r271 150 190 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.49 $Y=3.33
+ $X2=2.615 $Y2=3.33
r272 150 152 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.49 $Y=3.33
+ $X2=2.16 $Y2=3.33
r273 149 153 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r274 149 188 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r275 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r276 146 187 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.73 $Y2=3.33
r277 146 148 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=1.2 $Y2=3.33
r278 144 169 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r279 144 166 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r280 142 174 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=8.94 $Y=3.33
+ $X2=8.88 $Y2=3.33
r281 142 143 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.94 $Y=3.33
+ $X2=9.025 $Y2=3.33
r282 140 171 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=8.04 $Y=3.33
+ $X2=7.92 $Y2=3.33
r283 140 141 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.04 $Y=3.33
+ $X2=8.125 $Y2=3.33
r284 139 174 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.21 $Y=3.33
+ $X2=8.88 $Y2=3.33
r285 139 141 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.21 $Y=3.33
+ $X2=8.125 $Y2=3.33
r286 137 168 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.14 $Y=3.33
+ $X2=6.96 $Y2=3.33
r287 137 138 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.14 $Y=3.33
+ $X2=7.225 $Y2=3.33
r288 136 171 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.31 $Y=3.33
+ $X2=7.92 $Y2=3.33
r289 136 138 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.31 $Y=3.33
+ $X2=7.225 $Y2=3.33
r290 134 165 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=6.16 $Y=3.33
+ $X2=6 $Y2=3.33
r291 134 135 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.16 $Y=3.33
+ $X2=6.285 $Y2=3.33
r292 133 168 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=6.41 $Y=3.33
+ $X2=6.96 $Y2=3.33
r293 133 135 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.41 $Y=3.33
+ $X2=6.285 $Y2=3.33
r294 131 162 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.28 $Y=3.33
+ $X2=5.04 $Y2=3.33
r295 131 132 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.28 $Y=3.33
+ $X2=5.365 $Y2=3.33
r296 130 165 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.45 $Y=3.33
+ $X2=6 $Y2=3.33
r297 130 132 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.45 $Y=3.33
+ $X2=5.365 $Y2=3.33
r298 128 159 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.37 $Y=3.33
+ $X2=4.08 $Y2=3.33
r299 128 129 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.37 $Y=3.33
+ $X2=4.455 $Y2=3.33
r300 127 162 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=4.54 $Y=3.33
+ $X2=5.04 $Y2=3.33
r301 127 129 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=3.33
+ $X2=4.455 $Y2=3.33
r302 125 156 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.47 $Y=3.33
+ $X2=3.12 $Y2=3.33
r303 125 126 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.47 $Y=3.33
+ $X2=3.555 $Y2=3.33
r304 124 159 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r305 124 126 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=3.33
+ $X2=3.555 $Y2=3.33
r306 122 148 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.2 $Y2=3.33
r307 122 123 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.63 $Y2=3.33
r308 121 152 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=2.16 $Y2=3.33
r309 121 123 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=1.63 $Y2=3.33
r310 117 120 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=12.715 $Y=1.985
+ $X2=12.715 $Y2=2.815
r311 115 202 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=12.715
+ $Y=3.245 $X2=12.775 $Y2=3.33
r312 115 120 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=12.715 $Y=3.245
+ $X2=12.715 $Y2=2.815
r313 111 114 33.4208 $w=2.48e-07 $l=7.25e-07 $layer=LI1_cond $X=11.765 $Y=2.09
+ $X2=11.765 $Y2=2.815
r314 109 199 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.765 $Y=3.245
+ $X2=11.765 $Y2=3.33
r315 109 114 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.765 $Y=3.245
+ $X2=11.765 $Y2=2.815
r316 105 108 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=10.825 $Y=2.09
+ $X2=10.825 $Y2=2.815
r317 103 196 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.825 $Y=3.245
+ $X2=10.825 $Y2=3.33
r318 103 108 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=10.825 $Y=3.245
+ $X2=10.825 $Y2=2.815
r319 102 193 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.01 $Y=3.33
+ $X2=9.925 $Y2=3.33
r320 101 196 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.74 $Y=3.33
+ $X2=10.825 $Y2=3.33
r321 101 102 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=10.74 $Y=3.33
+ $X2=10.01 $Y2=3.33
r322 97 100 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=9.925 $Y=2.09
+ $X2=9.925 $Y2=2.815
r323 95 193 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.925 $Y=3.245
+ $X2=9.925 $Y2=3.33
r324 95 100 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=9.925 $Y=3.245
+ $X2=9.925 $Y2=2.815
r325 94 143 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.11 $Y=3.33
+ $X2=9.025 $Y2=3.33
r326 93 193 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.84 $Y=3.33
+ $X2=9.925 $Y2=3.33
r327 93 94 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=9.84 $Y=3.33
+ $X2=9.11 $Y2=3.33
r328 89 92 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=9.025 $Y=2.09
+ $X2=9.025 $Y2=2.815
r329 87 143 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.025 $Y=3.245
+ $X2=9.025 $Y2=3.33
r330 87 92 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=9.025 $Y=3.245
+ $X2=9.025 $Y2=2.815
r331 83 86 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=8.125 $Y=2.09
+ $X2=8.125 $Y2=2.815
r332 81 141 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.125 $Y=3.245
+ $X2=8.125 $Y2=3.33
r333 81 86 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.125 $Y=3.245
+ $X2=8.125 $Y2=2.815
r334 77 138 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.225 $Y=3.245
+ $X2=7.225 $Y2=3.33
r335 77 79 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=7.225 $Y=3.245
+ $X2=7.225 $Y2=2.325
r336 73 135 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.285 $Y=3.245
+ $X2=6.285 $Y2=3.33
r337 73 75 42.4099 $w=2.48e-07 $l=9.2e-07 $layer=LI1_cond $X=6.285 $Y=3.245
+ $X2=6.285 $Y2=2.325
r338 69 72 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=5.365 $Y=2.09
+ $X2=5.365 $Y2=2.815
r339 67 132 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.365 $Y=3.245
+ $X2=5.365 $Y2=3.33
r340 67 72 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=5.365 $Y=3.245
+ $X2=5.365 $Y2=2.815
r341 63 129 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=3.245
+ $X2=4.455 $Y2=3.33
r342 63 65 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.455 $Y=3.245
+ $X2=4.455 $Y2=2.325
r343 59 126 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.555 $Y=3.245
+ $X2=3.555 $Y2=3.33
r344 59 61 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.555 $Y=3.245
+ $X2=3.555 $Y2=2.325
r345 55 58 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=2.615 $Y=1.985
+ $X2=2.615 $Y2=2.815
r346 53 190 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.615 $Y=3.245
+ $X2=2.615 $Y2=3.33
r347 53 58 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.615 $Y=3.245
+ $X2=2.615 $Y2=2.815
r348 49 123 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=3.33
r349 49 51 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=2.305
r350 45 187 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r351 45 47 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.455
r352 14 120 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=12.54
+ $Y=1.84 $X2=12.675 $Y2=2.815
r353 14 117 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=12.54
+ $Y=1.84 $X2=12.675 $Y2=1.985
r354 13 114 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=11.59
+ $Y=1.84 $X2=11.725 $Y2=2.815
r355 13 111 400 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_PDIFF $count=1 $X=11.59
+ $Y=1.84 $X2=11.725 $Y2=2.09
r356 12 108 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.69
+ $Y=1.84 $X2=10.825 $Y2=2.815
r357 12 105 400 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_PDIFF $count=1 $X=10.69
+ $Y=1.84 $X2=10.825 $Y2=2.09
r358 11 100 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.79
+ $Y=1.84 $X2=9.925 $Y2=2.815
r359 11 97 400 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_PDIFF $count=1 $X=9.79
+ $Y=1.84 $X2=9.925 $Y2=2.09
r360 10 92 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.89
+ $Y=1.84 $X2=9.025 $Y2=2.815
r361 10 89 400 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_PDIFF $count=1 $X=8.89
+ $Y=1.84 $X2=9.025 $Y2=2.09
r362 9 86 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.99
+ $Y=1.84 $X2=8.125 $Y2=2.815
r363 9 83 400 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_PDIFF $count=1 $X=7.99
+ $Y=1.84 $X2=8.125 $Y2=2.09
r364 8 79 300 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=2 $X=7.09
+ $Y=1.84 $X2=7.225 $Y2=2.325
r365 7 75 300 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_PDIFF $count=2 $X=6.14
+ $Y=1.84 $X2=6.325 $Y2=2.325
r366 6 72 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.23
+ $Y=1.84 $X2=5.365 $Y2=2.815
r367 6 69 400 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_PDIFF $count=1 $X=5.23
+ $Y=1.84 $X2=5.365 $Y2=2.09
r368 5 65 300 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=2 $X=4.32
+ $Y=1.84 $X2=4.455 $Y2=2.325
r369 4 61 300 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=2 $X=3.42
+ $Y=1.84 $X2=3.555 $Y2=2.325
r370 3 58 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=2.51
+ $Y=1.84 $X2=2.655 $Y2=2.815
r371 3 55 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.51
+ $Y=1.84 $X2=2.655 $Y2=1.985
r372 2 51 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.84 $X2=1.63 $Y2=2.305
r373 1 47 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__BUFBUF_16%X 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 51 53 55 59 65 69 75 79 85 89 95 99 105 109 113 117 122 125 127 128 129 130
+ 131 132 133 140 141 145 146 150 151 155 156 160 161 165 170 171
c277 171 0 1.38532e-19 $X=12.2 $Y=2.035
c278 161 0 3.07445e-20 $X=10.375 $Y=1.92
c279 156 0 3.07333e-20 $X=9.475 $Y=1.92
c280 151 0 3.07333e-20 $X=8.575 $Y=1.92
c281 146 0 3.07333e-20 $X=7.675 $Y=1.92
c282 141 0 3.07333e-20 $X=6.775 $Y=1.92
c283 132 0 9.40629e-20 $X=12.18 $Y=1.15
c284 53 0 1.04236e-19 $X=5.825 $Y=2.085
c285 51 0 6.44981e-20 $X=5.8 $Y=0.515
r286 170 172 0.769762 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=12.225 $Y=2.035
+ $X2=12.225 $Y2=2.02
r287 170 171 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.2 $Y=2.035
+ $X2=12.2 $Y2=2.035
r288 168 171 0.590276 $w=2.3e-07 $l=9.2e-07 $layer=MET1_cond $X=11.28 $Y=2.035
+ $X2=12.2 $Y2=2.035
r289 165 168 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=2.035
+ $X2=11.28 $Y2=2.035
r290 165 166 4.36643 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=11.275 $Y=2.005
+ $X2=11.275 $Y2=1.92
r291 163 168 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=10.38 $Y=2.035
+ $X2=11.28 $Y2=2.035
r292 160 163 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.38 $Y=2.035
+ $X2=10.38 $Y2=2.035
r293 160 161 5.17556 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=10.375 $Y=2.005
+ $X2=10.375 $Y2=1.92
r294 158 163 0.571028 $w=2.3e-07 $l=8.9e-07 $layer=MET1_cond $X=9.49 $Y=2.035
+ $X2=10.38 $Y2=2.035
r295 155 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.49 $Y=2.035
+ $X2=9.49 $Y2=2.035
r296 155 156 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=9.475 $Y=2.005
+ $X2=9.475 $Y2=1.92
r297 150 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.57 $Y=2.035
+ $X2=8.57 $Y2=2.035
r298 150 151 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.575 $Y=2.005
+ $X2=8.575 $Y2=1.92
r299 148 153 0.571028 $w=2.3e-07 $l=8.9e-07 $layer=MET1_cond $X=7.68 $Y=2.035
+ $X2=8.57 $Y2=2.035
r300 145 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.68 $Y=2.035
+ $X2=7.68 $Y2=2.035
r301 145 146 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=7.675 $Y=2.005
+ $X2=7.675 $Y2=1.92
r302 143 148 0.590276 $w=2.3e-07 $l=9.2e-07 $layer=MET1_cond $X=6.76 $Y=2.035
+ $X2=7.68 $Y2=2.035
r303 140 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.76 $Y=2.035
+ $X2=6.76 $Y2=2.035
r304 140 141 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=6.775 $Y=2.005
+ $X2=6.775 $Y2=1.92
r305 138 143 0.587068 $w=2.3e-07 $l=9.15e-07 $layer=MET1_cond $X=5.845 $Y=2.035
+ $X2=6.76 $Y2=2.035
r306 136 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.845 $Y=2.035
+ $X2=5.845 $Y2=2.035
r307 133 158 0.288722 $w=2.3e-07 $l=4.5e-07 $layer=MET1_cond $X=9.04 $Y=2.035
+ $X2=9.49 $Y2=2.035
r308 133 153 0.301554 $w=2.3e-07 $l=4.7e-07 $layer=MET1_cond $X=9.04 $Y=2.035
+ $X2=8.57 $Y2=2.035
r309 131 161 16.1867 $w=1.83e-07 $l=2.7e-07 $layer=LI1_cond $X=10.302 $Y=1.65
+ $X2=10.302 $Y2=1.92
r310 130 156 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.395 $Y=1.65
+ $X2=9.395 $Y2=1.92
r311 129 151 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.495 $Y=1.65
+ $X2=8.495 $Y2=1.92
r312 128 146 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.595 $Y=1.65
+ $X2=7.595 $Y2=1.92
r313 127 141 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.695 $Y=1.65
+ $X2=6.695 $Y2=1.92
r314 123 170 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=12.225 $Y=2.185
+ $X2=12.225 $Y2=2.035
r315 123 125 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=12.225 $Y=2.185
+ $X2=12.225 $Y2=2.4
r316 122 172 1.41528 $w=2.83e-07 $l=3.5e-08 $layer=LI1_cond $X=12.202 $Y=1.985
+ $X2=12.202 $Y2=2.02
r317 122 132 33.7646 $w=2.83e-07 $l=8.35e-07 $layer=LI1_cond $X=12.202 $Y=1.985
+ $X2=12.202 $Y2=1.15
r318 115 132 6.00814 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.18 $Y=0.985
+ $X2=12.18 $Y2=1.15
r319 115 117 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=12.18 $Y=0.985
+ $X2=12.18 $Y2=0.515
r320 111 165 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=11.275 $Y=2.085
+ $X2=11.275 $Y2=2.005
r321 111 113 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=11.275 $Y=2.085
+ $X2=11.275 $Y2=2.815
r322 109 166 75.3108 $w=2.13e-07 $l=1.405e-06 $layer=LI1_cond $X=11.217 $Y=0.515
+ $X2=11.217 $Y2=1.92
r323 103 160 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=10.375 $Y=2.085
+ $X2=10.375 $Y2=2.005
r324 103 105 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=10.375 $Y=2.085
+ $X2=10.375 $Y2=2.815
r325 97 131 6.56491 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=10.27 $Y=1.525
+ $X2=10.27 $Y2=1.65
r326 97 99 46.5587 $w=2.48e-07 $l=1.01e-06 $layer=LI1_cond $X=10.27 $Y=1.525
+ $X2=10.27 $Y2=0.515
r327 93 155 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=9.475 $Y=2.085
+ $X2=9.475 $Y2=2.005
r328 93 95 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=9.475 $Y=2.085
+ $X2=9.475 $Y2=2.815
r329 87 130 7.21712 $w=2.63e-07 $l=1.32e-07 $layer=LI1_cond $X=9.347 $Y=1.518
+ $X2=9.347 $Y2=1.65
r330 87 89 43.6189 $w=2.63e-07 $l=1.003e-06 $layer=LI1_cond $X=9.347 $Y=1.518
+ $X2=9.347 $Y2=0.515
r331 83 150 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=8.575 $Y=2.085
+ $X2=8.575 $Y2=2.005
r332 83 85 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=8.575 $Y=2.085
+ $X2=8.575 $Y2=2.815
r333 77 129 7.79447 $w=2.93e-07 $l=1.47e-07 $layer=LI1_cond $X=8.432 $Y=1.503
+ $X2=8.432 $Y2=1.65
r334 77 79 38.5971 $w=2.93e-07 $l=9.88e-07 $layer=LI1_cond $X=8.432 $Y=1.503
+ $X2=8.432 $Y2=0.515
r335 73 145 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.675 $Y=2.085
+ $X2=7.675 $Y2=2.005
r336 73 75 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=7.675 $Y=2.085
+ $X2=7.675 $Y2=2.815
r337 67 128 7.79447 $w=2.93e-07 $l=1.47e-07 $layer=LI1_cond $X=7.532 $Y=1.503
+ $X2=7.532 $Y2=1.65
r338 67 69 38.5971 $w=2.93e-07 $l=9.88e-07 $layer=LI1_cond $X=7.532 $Y=1.503
+ $X2=7.532 $Y2=0.515
r339 63 140 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=6.775 $Y=2.085
+ $X2=6.775 $Y2=2.005
r340 63 65 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=6.775 $Y=2.085
+ $X2=6.775 $Y2=2.815
r341 57 127 6.82988 $w=2.43e-07 $l=1.22e-07 $layer=LI1_cond $X=6.657 $Y=1.528
+ $X2=6.657 $Y2=1.65
r342 57 59 47.65 $w=2.43e-07 $l=1.013e-06 $layer=LI1_cond $X=6.657 $Y=1.528
+ $X2=6.657 $Y2=0.515
r343 53 136 2.98307 $w=3.3e-07 $l=8.12404e-08 $layer=LI1_cond $X=5.825 $Y=2.085
+ $X2=5.812 $Y2=2.01
r344 53 55 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=5.825 $Y=2.085
+ $X2=5.825 $Y2=2.815
r345 49 136 10.152 $w=2.9e-07 $l=2.59702e-07 $layer=LI1_cond $X=5.76 $Y=1.775
+ $X2=5.812 $Y2=2.01
r346 49 51 58.0831 $w=2.48e-07 $l=1.26e-06 $layer=LI1_cond $X=5.76 $Y=1.775
+ $X2=5.76 $Y2=0.515
r347 16 125 300 $w=1.7e-07 $l=6.4591e-07 $layer=licon1_PDIFF $count=2 $X=12.04
+ $Y=1.84 $X2=12.225 $Y2=2.4
r348 16 122 600 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=12.04
+ $Y=1.84 $X2=12.225 $Y2=1.985
r349 15 165 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=11.14
+ $Y=1.84 $X2=11.275 $Y2=2.005
r350 15 113 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=11.14
+ $Y=1.84 $X2=11.275 $Y2=2.815
r351 14 160 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=10.24
+ $Y=1.84 $X2=10.375 $Y2=2.005
r352 14 105 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.24
+ $Y=1.84 $X2=10.375 $Y2=2.815
r353 13 155 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=9.34
+ $Y=1.84 $X2=9.475 $Y2=2.005
r354 13 95 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.34
+ $Y=1.84 $X2=9.475 $Y2=2.815
r355 12 150 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=8.44
+ $Y=1.84 $X2=8.575 $Y2=2.005
r356 12 85 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.44
+ $Y=1.84 $X2=8.575 $Y2=2.815
r357 11 145 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=7.54
+ $Y=1.84 $X2=7.675 $Y2=2.005
r358 11 75 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.54
+ $Y=1.84 $X2=7.675 $Y2=2.815
r359 10 140 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=6.64
+ $Y=1.84 $X2=6.775 $Y2=2.005
r360 10 65 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.64
+ $Y=1.84 $X2=6.775 $Y2=2.815
r361 9 136 400 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=5.69
+ $Y=1.84 $X2=5.825 $Y2=2.01
r362 9 55 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.69
+ $Y=1.84 $X2=5.825 $Y2=2.815
r363 8 117 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.04
+ $Y=0.37 $X2=12.18 $Y2=0.515
r364 7 109 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.1
+ $Y=0.37 $X2=11.24 $Y2=0.515
r365 6 99 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.17
+ $Y=0.37 $X2=10.31 $Y2=0.515
r366 5 89 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.24
+ $Y=0.37 $X2=9.38 $Y2=0.515
r367 4 79 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.31
+ $Y=0.37 $X2=8.45 $Y2=0.515
r368 3 69 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.38
+ $Y=0.37 $X2=7.52 $Y2=0.515
r369 2 59 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.52
+ $Y=0.37 $X2=6.66 $Y2=0.515
r370 1 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.66
+ $Y=0.37 $X2=5.8 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__BUFBUF_16%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 14 45
+ 49 53 57 61 65 69 71 75 77 81 85 89 93 97 99 101 104 105 107 108 110 111 113
+ 114 115 116 118 119 120 122 131 148 153 158 167 172 175 178 181 184 187 190
+ 194
r222 193 194 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r223 190 191 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r224 187 188 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r225 184 185 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r226 181 182 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r227 179 182 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.92 $Y2=0
r228 178 179 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r229 175 176 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r230 172 173 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r231 170 194 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r232 169 170 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r233 167 193 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=12.515 $Y=0
+ $X2=12.737 $Y2=0
r234 167 169 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=12.515 $Y=0
+ $X2=12.24 $Y2=0
r235 166 170 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=12.24 $Y2=0
r236 166 191 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r237 165 166 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r238 163 190 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.905 $Y=0
+ $X2=10.74 $Y2=0
r239 163 165 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=10.905 $Y=0
+ $X2=11.28 $Y2=0
r240 162 191 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r241 162 188 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r242 161 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r243 159 187 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=9.975 $Y=0
+ $X2=9.82 $Y2=0
r244 159 161 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.975 $Y=0
+ $X2=10.32 $Y2=0
r245 158 190 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.575 $Y=0
+ $X2=10.74 $Y2=0
r246 158 161 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=10.575 $Y=0
+ $X2=10.32 $Y2=0
r247 157 188 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r248 157 185 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r249 156 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r250 154 184 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=9.045 $Y=0
+ $X2=8.897 $Y2=0
r251 154 156 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.045 $Y=0
+ $X2=9.36 $Y2=0
r252 153 187 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=9.665 $Y=0
+ $X2=9.82 $Y2=0
r253 153 156 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.665 $Y=0
+ $X2=9.36 $Y2=0
r254 152 185 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=8.88 $Y2=0
r255 152 182 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=7.92 $Y2=0
r256 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r257 149 181 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=8.115 $Y=0
+ $X2=7.982 $Y2=0
r258 149 151 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.115 $Y=0
+ $X2=8.4 $Y2=0
r259 148 184 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=8.75 $Y=0
+ $X2=8.897 $Y2=0
r260 148 151 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=8.75 $Y=0 $X2=8.4
+ $Y2=0
r261 146 147 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r262 144 147 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r263 143 144 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r264 141 144 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=5.04 $Y2=0
r265 140 141 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r266 138 141 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=4.08 $Y2=0
r267 138 176 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=2.64 $Y2=0
r268 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r269 135 175 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=0
+ $X2=2.58 $Y2=0
r270 135 137 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.745 $Y=0
+ $X2=3.12 $Y2=0
r271 134 176 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=2.64 $Y2=0
r272 133 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r273 131 175 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=0
+ $X2=2.58 $Y2=0
r274 131 133 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.415 $Y=0
+ $X2=2.16 $Y2=0
r275 130 134 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0
+ $X2=2.16 $Y2=0
r276 130 173 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0
+ $X2=0.72 $Y2=0
r277 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r278 127 172 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=0
+ $X2=0.725 $Y2=0
r279 127 129 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.89 $Y=0 $X2=1.2
+ $Y2=0
r280 125 173 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r281 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r282 122 172 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.56 $Y=0
+ $X2=0.725 $Y2=0
r283 122 124 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.24
+ $Y2=0
r284 120 179 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r285 120 147 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r286 118 165 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=11.505 $Y=0
+ $X2=11.28 $Y2=0
r287 118 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.505 $Y=0
+ $X2=11.67 $Y2=0
r288 117 169 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=11.835 $Y=0
+ $X2=12.24 $Y2=0
r289 117 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.835 $Y=0
+ $X2=11.67 $Y2=0
r290 115 146 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.065 $Y=0 $X2=6
+ $Y2=0
r291 115 116 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.065 $Y=0
+ $X2=6.19 $Y2=0
r292 113 143 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.275 $Y=0
+ $X2=5.04 $Y2=0
r293 113 114 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=5.275 $Y=0 $X2=5.365
+ $Y2=0
r294 112 146 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=5.455 $Y=0 $X2=6
+ $Y2=0
r295 112 114 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=5.455 $Y=0 $X2=5.365
+ $Y2=0
r296 110 140 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=4.275 $Y=0
+ $X2=4.08 $Y2=0
r297 110 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.275 $Y=0
+ $X2=4.44 $Y2=0
r298 109 143 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.605 $Y=0
+ $X2=5.04 $Y2=0
r299 109 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.605 $Y=0
+ $X2=4.44 $Y2=0
r300 107 137 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.345 $Y=0
+ $X2=3.12 $Y2=0
r301 107 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.345 $Y=0
+ $X2=3.51 $Y2=0
r302 106 140 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.675 $Y=0
+ $X2=4.08 $Y2=0
r303 106 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.675 $Y=0
+ $X2=3.51 $Y2=0
r304 104 129 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.42 $Y=0 $X2=1.2
+ $Y2=0
r305 104 105 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.42 $Y=0
+ $X2=1.545 $Y2=0
r306 103 133 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.67 $Y=0
+ $X2=2.16 $Y2=0
r307 103 105 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.67 $Y=0
+ $X2=1.545 $Y2=0
r308 99 193 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=12.68 $Y=0.085
+ $X2=12.737 $Y2=0
r309 99 101 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=12.68 $Y=0.085
+ $X2=12.68 $Y2=0.515
r310 95 119 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.67 $Y=0.085
+ $X2=11.67 $Y2=0
r311 95 97 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.67 $Y=0.085
+ $X2=11.67 $Y2=0.515
r312 91 190 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.74 $Y=0.085
+ $X2=10.74 $Y2=0
r313 91 93 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.74 $Y=0.085
+ $X2=10.74 $Y2=0.515
r314 87 187 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=9.82 $Y=0.085
+ $X2=9.82 $Y2=0
r315 87 89 15.9855 $w=3.08e-07 $l=4.3e-07 $layer=LI1_cond $X=9.82 $Y=0.085
+ $X2=9.82 $Y2=0.515
r316 83 184 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=8.897 $Y=0.085
+ $X2=8.897 $Y2=0
r317 83 85 16.7983 $w=2.93e-07 $l=4.3e-07 $layer=LI1_cond $X=8.897 $Y=0.085
+ $X2=8.897 $Y2=0.515
r318 79 181 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=7.982 $Y=0.085
+ $X2=7.982 $Y2=0
r319 79 81 18.7 $w=2.63e-07 $l=4.3e-07 $layer=LI1_cond $X=7.982 $Y=0.085
+ $X2=7.982 $Y2=0.515
r320 78 178 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=7.175 $Y=0
+ $X2=7.067 $Y2=0
r321 77 181 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=7.85 $Y=0
+ $X2=7.982 $Y2=0
r322 77 78 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=7.85 $Y=0
+ $X2=7.175 $Y2=0
r323 73 178 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=7.067 $Y=0.085
+ $X2=7.067 $Y2=0
r324 73 75 23.0489 $w=2.13e-07 $l=4.3e-07 $layer=LI1_cond $X=7.067 $Y=0.085
+ $X2=7.067 $Y2=0.515
r325 72 116 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.315 $Y=0
+ $X2=6.19 $Y2=0
r326 71 178 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=6.96 $Y=0
+ $X2=7.067 $Y2=0
r327 71 72 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=6.96 $Y=0
+ $X2=6.315 $Y2=0
r328 67 116 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.19 $Y=0.085
+ $X2=6.19 $Y2=0
r329 67 69 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6.19 $Y=0.085
+ $X2=6.19 $Y2=0.515
r330 63 114 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.365 $Y=0.085
+ $X2=5.365 $Y2=0
r331 63 65 30.5 $w=1.78e-07 $l=4.95e-07 $layer=LI1_cond $X=5.365 $Y=0.085
+ $X2=5.365 $Y2=0.58
r332 59 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.44 $Y=0.085
+ $X2=4.44 $Y2=0
r333 59 61 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=4.44 $Y=0.085
+ $X2=4.44 $Y2=0.645
r334 55 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.51 $Y=0.085
+ $X2=3.51 $Y2=0
r335 55 57 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=3.51 $Y=0.085
+ $X2=3.51 $Y2=0.645
r336 51 175 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=0.085
+ $X2=2.58 $Y2=0
r337 51 53 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.58 $Y=0.085
+ $X2=2.58 $Y2=0.515
r338 47 105 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.545 $Y=0.085
+ $X2=1.545 $Y2=0
r339 47 49 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=1.545 $Y=0.085
+ $X2=1.545 $Y2=0.625
r340 43 172 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=0.085
+ $X2=0.725 $Y2=0
r341 43 45 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=0.725 $Y=0.085
+ $X2=0.725 $Y2=0.625
r342 14 101 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=12.47
+ $Y=0.37 $X2=12.68 $Y2=0.515
r343 13 97 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.53
+ $Y=0.37 $X2=11.67 $Y2=0.515
r344 12 93 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.6
+ $Y=0.37 $X2=10.74 $Y2=0.515
r345 11 89 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.67
+ $Y=0.37 $X2=9.81 $Y2=0.515
r346 10 85 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.74
+ $Y=0.37 $X2=8.88 $Y2=0.515
r347 9 81 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.81
+ $Y=0.37 $X2=7.95 $Y2=0.515
r348 8 75 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.95
+ $Y=0.37 $X2=7.09 $Y2=0.515
r349 7 69 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.09
+ $Y=0.37 $X2=6.23 $Y2=0.515
r350 6 65 91 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=2 $X=5.23
+ $Y=0.37 $X2=5.37 $Y2=0.58
r351 5 61 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=4.3
+ $Y=0.37 $X2=4.44 $Y2=0.645
r352 4 57 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.37
+ $Y=0.37 $X2=3.51 $Y2=0.645
r353 3 53 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=2.435
+ $Y=0.37 $X2=2.58 $Y2=0.515
r354 2 49 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.37 $X2=1.585 $Y2=0.625
r355 1 45 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=0.585
+ $Y=0.37 $X2=0.725 $Y2=0.625
.ends


* File: sky130_fd_sc_ms__and4b_1.pxi.spice
* Created: Fri Aug 28 17:13:58 2020
* 
x_PM_SKY130_FD_SC_MS__AND4B_1%A_N N_A_N_M1004_g N_A_N_M1007_g N_A_N_c_86_n
+ N_A_N_c_91_n A_N N_A_N_c_87_n N_A_N_c_88_n PM_SKY130_FD_SC_MS__AND4B_1%A_N
x_PM_SKY130_FD_SC_MS__AND4B_1%A_27_74# N_A_27_74#_M1007_s N_A_27_74#_M1004_s
+ N_A_27_74#_M1002_g N_A_27_74#_c_124_n N_A_27_74#_c_125_n N_A_27_74#_c_126_n
+ N_A_27_74#_M1003_g N_A_27_74#_c_127_n N_A_27_74#_c_135_n N_A_27_74#_c_128_n
+ N_A_27_74#_c_129_n N_A_27_74#_c_136_n N_A_27_74#_c_137_n N_A_27_74#_c_130_n
+ N_A_27_74#_c_138_n N_A_27_74#_c_131_n N_A_27_74#_c_132_n N_A_27_74#_c_133_n
+ PM_SKY130_FD_SC_MS__AND4B_1%A_27_74#
x_PM_SKY130_FD_SC_MS__AND4B_1%B N_B_M1006_g N_B_M1001_g N_B_c_209_n N_B_c_210_n
+ B B PM_SKY130_FD_SC_MS__AND4B_1%B
x_PM_SKY130_FD_SC_MS__AND4B_1%C N_C_M1011_g N_C_M1009_g N_C_c_247_n C C
+ N_C_c_248_n N_C_c_249_n PM_SKY130_FD_SC_MS__AND4B_1%C
x_PM_SKY130_FD_SC_MS__AND4B_1%D N_D_M1008_g N_D_M1000_g D N_D_c_291_n
+ PM_SKY130_FD_SC_MS__AND4B_1%D
x_PM_SKY130_FD_SC_MS__AND4B_1%A_229_424# N_A_229_424#_M1003_s
+ N_A_229_424#_M1002_d N_A_229_424#_M1009_d N_A_229_424#_M1010_g
+ N_A_229_424#_M1005_g N_A_229_424#_c_328_n N_A_229_424#_c_329_n
+ N_A_229_424#_c_330_n N_A_229_424#_c_331_n N_A_229_424#_c_332_n
+ N_A_229_424#_c_338_n N_A_229_424#_c_341_n N_A_229_424#_c_375_n
+ N_A_229_424#_c_363_n N_A_229_424#_c_339_n N_A_229_424#_c_333_n
+ N_A_229_424#_c_334_n PM_SKY130_FD_SC_MS__AND4B_1%A_229_424#
x_PM_SKY130_FD_SC_MS__AND4B_1%VPWR N_VPWR_M1004_d N_VPWR_M1006_d N_VPWR_M1008_d
+ N_VPWR_c_432_n N_VPWR_c_433_n N_VPWR_c_434_n N_VPWR_c_435_n VPWR
+ N_VPWR_c_436_n N_VPWR_c_437_n N_VPWR_c_431_n N_VPWR_c_439_n N_VPWR_c_440_n
+ N_VPWR_c_441_n PM_SKY130_FD_SC_MS__AND4B_1%VPWR
x_PM_SKY130_FD_SC_MS__AND4B_1%X N_X_M1005_d N_X_M1010_d N_X_c_479_n N_X_c_480_n
+ X X X X N_X_c_481_n PM_SKY130_FD_SC_MS__AND4B_1%X
x_PM_SKY130_FD_SC_MS__AND4B_1%VGND N_VGND_M1007_d N_VGND_M1000_d N_VGND_c_503_n
+ N_VGND_c_504_n VGND N_VGND_c_505_n N_VGND_c_506_n N_VGND_c_507_n
+ N_VGND_c_508_n N_VGND_c_509_n N_VGND_c_510_n PM_SKY130_FD_SC_MS__AND4B_1%VGND
cc_1 VNB N_A_N_M1007_g 0.0371391f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_2 VNB N_A_N_c_86_n 0.0249613f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.695
cc_3 VNB N_A_N_c_87_n 0.0184956f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.355
cc_4 VNB N_A_N_c_88_n 0.0229758f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.355
cc_5 VNB N_A_27_74#_c_124_n 0.0305639f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_6 VNB N_A_27_74#_c_125_n 0.0108824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_74#_c_126_n 0.0132493f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.355
cc_8 VNB N_A_27_74#_c_127_n 0.0214334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_74#_c_128_n 0.0105312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_74#_c_129_n 0.00992961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_74#_c_130_n 0.0108784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_c_131_n 0.00226763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_132_n 0.0174747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_74#_c_133_n 0.0668854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_M1001_g 0.0301282f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_16 VNB N_B_c_209_n 0.0158757f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.355
cc_17 VNB N_B_c_210_n 0.0334807f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.19
cc_18 VNB B 0.00854044f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.86
cc_19 VNB N_C_M1011_g 0.00933542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_C_M1009_g 0.0196984f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_21 VNB N_C_c_247_n 0.0158127f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.19
cc_22 VNB N_C_c_248_n 0.0412509f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.355
cc_23 VNB N_C_c_249_n 0.025844f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.355
cc_24 VNB N_D_M1008_g 0.00218404f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_25 VNB N_D_M1000_g 0.0298855f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.645
cc_26 VNB D 0.00251027f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.355
cc_27 VNB N_D_c_291_n 0.0247607f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.86
cc_28 VNB N_A_229_424#_c_328_n 0.00846748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_229_424#_c_329_n 0.00939658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_229_424#_c_330_n 0.0105635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_229_424#_c_331_n 0.00482938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_229_424#_c_332_n 0.0214217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_229_424#_c_333_n 0.0279422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_229_424#_c_334_n 0.0215792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VPWR_c_431_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_X_c_479_n 0.0240518f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.355
cc_37 VNB N_X_c_480_n 0.00694384f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_38 VNB N_X_c_481_n 0.0219872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_503_n 0.0175884f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.355
cc_40 VNB N_VGND_c_504_n 0.0190854f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_41 VNB N_VGND_c_505_n 0.0181399f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=1.355
cc_42 VNB N_VGND_c_506_n 0.0705391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_507_n 0.019578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_508_n 0.293095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_509_n 0.00577043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_510_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VPB N_A_N_M1004_g 0.0379135f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_48 VPB N_A_N_c_86_n 0.00268144f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.695
cc_49 VPB N_A_N_c_91_n 0.0168639f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.86
cc_50 VPB N_A_N_c_88_n 0.0103985f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.355
cc_51 VPB N_A_27_74#_M1002_g 0.0292502f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.355
cc_52 VPB N_A_27_74#_c_135_n 0.0322185f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_27_74#_c_136_n 0.00746154f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_27_74#_c_137_n 0.00998527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_27_74#_c_138_n 0.0032226f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_27_74#_c_131_n 0.00358177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_27_74#_c_132_n 0.018232f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_B_M1006_g 0.029067f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_59 VPB N_B_c_209_n 8.35876e-19 $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.355
cc_60 VPB N_B_c_210_n 0.0153875f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.19
cc_61 VPB B 4.81172e-19 $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.86
cc_62 VPB N_C_M1009_g 0.0289389f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.645
cc_63 VPB N_D_M1008_g 0.0277097f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_64 VPB D 0.00257344f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.355
cc_65 VPB N_D_c_291_n 0.00982008f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.86
cc_66 VPB N_A_229_424#_M1010_g 0.0289595f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.86
cc_67 VPB N_A_229_424#_c_331_n 0.00176042f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A_229_424#_c_332_n 0.00422694f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A_229_424#_c_338_n 0.00275226f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_229_424#_c_339_n 0.00858131f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_229_424#_c_333_n 0.00616292f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_432_n 0.00983032f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.86
cc_73 VPB N_VPWR_c_433_n 0.0157671f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.525
cc_74 VPB N_VPWR_c_434_n 0.0207378f $X=-0.19 $Y=1.66 $X2=0.43 $Y2=1.525
cc_75 VPB N_VPWR_c_435_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_436_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_437_n 0.0202291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_431_n 0.0743094f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_439_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_440_n 0.0220529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_441_n 0.0274499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB X 0.00694384f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB X 0.040201f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_X_c_481_n 0.00904998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 N_A_N_M1004_g N_A_27_74#_M1002_g 0.0132466f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_86 N_A_N_M1007_g N_A_27_74#_c_125_n 0.0114901f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_87 N_A_N_M1007_g N_A_27_74#_c_127_n 0.00226722f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_88 N_A_N_M1004_g N_A_27_74#_c_135_n 0.0144049f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_89 N_A_N_M1007_g N_A_27_74#_c_128_n 0.0140234f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_90 N_A_N_c_87_n N_A_27_74#_c_128_n 0.00104829f $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_91 N_A_N_c_88_n N_A_27_74#_c_128_n 0.0144955f $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_92 N_A_N_c_87_n N_A_27_74#_c_129_n 0.00375152f $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_93 N_A_N_c_88_n N_A_27_74#_c_129_n 0.0254263f $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_94 N_A_N_M1004_g N_A_27_74#_c_136_n 0.0131848f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_95 N_A_N_c_88_n N_A_27_74#_c_136_n 0.0113214f $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_96 N_A_N_M1004_g N_A_27_74#_c_137_n 0.00269884f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_97 N_A_N_c_91_n N_A_27_74#_c_137_n 0.00402688f $X=0.43 $Y=1.86 $X2=0 $Y2=0
cc_98 N_A_N_c_88_n N_A_27_74#_c_137_n 0.0288658f $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_99 N_A_N_M1007_g N_A_27_74#_c_130_n 0.00374114f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_100 N_A_N_c_87_n N_A_27_74#_c_130_n 0.0013621f $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_101 N_A_N_c_88_n N_A_27_74#_c_130_n 0.0266416f $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_102 N_A_N_M1004_g N_A_27_74#_c_138_n 0.00321029f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_103 N_A_N_c_86_n N_A_27_74#_c_131_n 0.00120873f $X=0.43 $Y=1.695 $X2=0 $Y2=0
cc_104 N_A_N_c_91_n N_A_27_74#_c_131_n 5.12143e-19 $X=0.43 $Y=1.86 $X2=0 $Y2=0
cc_105 N_A_N_c_88_n N_A_27_74#_c_131_n 0.0248669f $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_106 N_A_N_c_86_n N_A_27_74#_c_132_n 0.0120054f $X=0.43 $Y=1.695 $X2=0 $Y2=0
cc_107 N_A_N_c_88_n N_A_27_74#_c_132_n 3.08399e-19 $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_108 N_A_N_c_87_n N_A_27_74#_c_133_n 0.00596009f $X=0.43 $Y=1.355 $X2=0 $Y2=0
cc_109 N_A_N_M1004_g N_A_229_424#_c_341_n 3.27875e-19 $X=0.505 $Y=2.54 $X2=0
+ $Y2=0
cc_110 N_A_N_M1004_g N_VPWR_c_432_n 0.00343717f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_111 N_A_N_M1004_g N_VPWR_c_436_n 0.005209f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_112 N_A_N_M1004_g N_VPWR_c_431_n 0.00986318f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_113 N_A_N_M1007_g N_VGND_c_503_n 0.00527104f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_114 N_A_N_M1007_g N_VGND_c_505_n 0.00461464f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_115 N_A_N_M1007_g N_VGND_c_508_n 0.00473629f $X=0.495 $Y=0.645 $X2=0 $Y2=0
cc_116 N_A_27_74#_c_126_n N_B_M1001_g 0.0314813f $X=1.69 $Y=0.545 $X2=0 $Y2=0
cc_117 N_A_27_74#_M1002_g N_B_c_209_n 0.0346297f $X=1.055 $Y=2.54 $X2=0 $Y2=0
cc_118 N_A_27_74#_c_126_n N_B_c_209_n 0.00834734f $X=1.69 $Y=0.545 $X2=0 $Y2=0
cc_119 N_A_27_74#_c_131_n N_B_c_209_n 0.00110467f $X=1.09 $Y=1.715 $X2=0 $Y2=0
cc_120 N_A_27_74#_c_132_n N_B_c_209_n 0.0141668f $X=1.09 $Y=1.715 $X2=0 $Y2=0
cc_121 N_A_27_74#_M1002_g B 2.76265e-19 $X=1.055 $Y=2.54 $X2=0 $Y2=0
cc_122 N_A_27_74#_c_126_n B 0.00104663f $X=1.69 $Y=0.545 $X2=0 $Y2=0
cc_123 N_A_27_74#_c_138_n B 0.00232826f $X=0.86 $Y=2.03 $X2=0 $Y2=0
cc_124 N_A_27_74#_c_131_n B 0.0170835f $X=1.09 $Y=1.715 $X2=0 $Y2=0
cc_125 N_A_27_74#_c_132_n B 8.62975e-19 $X=1.09 $Y=1.715 $X2=0 $Y2=0
cc_126 N_A_27_74#_c_124_n N_C_c_248_n 0.00170036f $X=1.615 $Y=0.47 $X2=0 $Y2=0
cc_127 N_A_27_74#_c_124_n N_C_c_249_n 0.00647686f $X=1.615 $Y=0.47 $X2=0 $Y2=0
cc_128 N_A_27_74#_c_124_n N_A_229_424#_c_328_n 0.0052648f $X=1.615 $Y=0.47 $X2=0
+ $Y2=0
cc_129 N_A_27_74#_c_126_n N_A_229_424#_c_328_n 0.0119422f $X=1.69 $Y=0.545 $X2=0
+ $Y2=0
cc_130 N_A_27_74#_c_128_n N_A_229_424#_c_328_n 0.0088137f $X=0.775 $Y=0.935
+ $X2=0 $Y2=0
cc_131 N_A_27_74#_c_130_n N_A_229_424#_c_328_n 0.00880168f $X=0.86 $Y=1.55 $X2=0
+ $Y2=0
cc_132 N_A_27_74#_c_133_n N_A_229_424#_c_328_n 0.0099514f $X=1.09 $Y=1.55 $X2=0
+ $Y2=0
cc_133 N_A_27_74#_c_126_n N_A_229_424#_c_329_n 0.0102279f $X=1.69 $Y=0.545 $X2=0
+ $Y2=0
cc_134 N_A_27_74#_c_126_n N_A_229_424#_c_330_n 0.00196337f $X=1.69 $Y=0.545
+ $X2=0 $Y2=0
cc_135 N_A_27_74#_c_130_n N_A_229_424#_c_330_n 0.00841426f $X=0.86 $Y=1.55 $X2=0
+ $Y2=0
cc_136 N_A_27_74#_c_133_n N_A_229_424#_c_330_n 0.00218369f $X=1.09 $Y=1.55 $X2=0
+ $Y2=0
cc_137 N_A_27_74#_M1002_g N_A_229_424#_c_341_n 0.0072371f $X=1.055 $Y=2.54 $X2=0
+ $Y2=0
cc_138 N_A_27_74#_c_135_n N_A_229_424#_c_341_n 0.00425729f $X=0.28 $Y=2.265
+ $X2=0 $Y2=0
cc_139 N_A_27_74#_c_131_n N_A_229_424#_c_341_n 0.00625929f $X=1.09 $Y=1.715
+ $X2=0 $Y2=0
cc_140 N_A_27_74#_c_132_n N_A_229_424#_c_341_n 0.0026046f $X=1.09 $Y=1.715 $X2=0
+ $Y2=0
cc_141 N_A_27_74#_c_136_n N_VPWR_M1004_d 0.00331335f $X=0.775 $Y=2.115 $X2=-0.19
+ $Y2=-0.245
cc_142 N_A_27_74#_M1002_g N_VPWR_c_432_n 0.00382308f $X=1.055 $Y=2.54 $X2=0
+ $Y2=0
cc_143 N_A_27_74#_c_135_n N_VPWR_c_432_n 0.0236791f $X=0.28 $Y=2.265 $X2=0 $Y2=0
cc_144 N_A_27_74#_c_136_n N_VPWR_c_432_n 0.0213327f $X=0.775 $Y=2.115 $X2=0
+ $Y2=0
cc_145 N_A_27_74#_c_135_n N_VPWR_c_436_n 0.014549f $X=0.28 $Y=2.265 $X2=0 $Y2=0
cc_146 N_A_27_74#_M1002_g N_VPWR_c_431_n 0.0108979f $X=1.055 $Y=2.54 $X2=0 $Y2=0
cc_147 N_A_27_74#_c_135_n N_VPWR_c_431_n 0.0119743f $X=0.28 $Y=2.265 $X2=0 $Y2=0
cc_148 N_A_27_74#_M1002_g N_VPWR_c_440_n 0.00553757f $X=1.055 $Y=2.54 $X2=0
+ $Y2=0
cc_149 N_A_27_74#_M1002_g N_VPWR_c_441_n 0.00255256f $X=1.055 $Y=2.54 $X2=0
+ $Y2=0
cc_150 N_A_27_74#_c_128_n N_VGND_M1007_d 0.0025118f $X=0.775 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_151 N_A_27_74#_c_125_n N_VGND_c_503_n 0.0059979f $X=1.255 $Y=0.47 $X2=0 $Y2=0
cc_152 N_A_27_74#_c_127_n N_VGND_c_503_n 0.00155433f $X=0.28 $Y=0.645 $X2=0
+ $Y2=0
cc_153 N_A_27_74#_c_128_n N_VGND_c_503_n 0.0206247f $X=0.775 $Y=0.935 $X2=0
+ $Y2=0
cc_154 N_A_27_74#_c_127_n N_VGND_c_505_n 0.0128369f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_155 N_A_27_74#_c_125_n N_VGND_c_506_n 0.017157f $X=1.255 $Y=0.47 $X2=0 $Y2=0
cc_156 N_A_27_74#_c_125_n N_VGND_c_508_n 0.0206598f $X=1.255 $Y=0.47 $X2=0 $Y2=0
cc_157 N_A_27_74#_c_127_n N_VGND_c_508_n 0.0106314f $X=0.28 $Y=0.645 $X2=0 $Y2=0
cc_158 N_A_27_74#_c_128_n N_VGND_c_508_n 0.00853677f $X=0.775 $Y=0.935 $X2=0
+ $Y2=0
cc_159 N_B_M1001_g N_C_M1009_g 0.013881f $X=2.165 $Y=1.015 $X2=0 $Y2=0
cc_160 B N_C_M1009_g 0.00297631f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_161 N_B_M1001_g N_C_c_248_n 0.0564627f $X=2.165 $Y=1.015 $X2=0 $Y2=0
cc_162 N_B_M1001_g N_C_c_249_n 0.0101643f $X=2.165 $Y=1.015 $X2=0 $Y2=0
cc_163 N_B_M1001_g N_A_229_424#_c_328_n 0.00265403f $X=2.165 $Y=1.015 $X2=0
+ $Y2=0
cc_164 N_B_M1001_g N_A_229_424#_c_329_n 0.0122201f $X=2.165 $Y=1.015 $X2=0 $Y2=0
cc_165 N_B_c_210_n N_A_229_424#_c_329_n 0.00185324f $X=2.09 $Y=1.795 $X2=0 $Y2=0
cc_166 B N_A_229_424#_c_329_n 0.0495197f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_167 N_B_c_209_n N_A_229_424#_c_330_n 0.00345348f $X=1.675 $Y=1.795 $X2=0
+ $Y2=0
cc_168 B N_A_229_424#_c_330_n 0.00662497f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_169 N_B_M1001_g N_A_229_424#_c_331_n 0.00134042f $X=2.165 $Y=1.015 $X2=0
+ $Y2=0
cc_170 B N_A_229_424#_c_331_n 0.0206597f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_171 N_B_M1006_g N_A_229_424#_c_363_n 0.0238183f $X=1.585 $Y=2.54 $X2=0 $Y2=0
cc_172 N_B_c_210_n N_A_229_424#_c_363_n 0.0131613f $X=2.09 $Y=1.795 $X2=0 $Y2=0
cc_173 B N_A_229_424#_c_363_n 0.0519859f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_174 N_B_M1006_g N_VPWR_c_431_n 0.00904737f $X=1.585 $Y=2.54 $X2=0 $Y2=0
cc_175 N_B_M1006_g N_VPWR_c_440_n 0.00460063f $X=1.585 $Y=2.54 $X2=0 $Y2=0
cc_176 N_B_M1006_g N_VPWR_c_441_n 0.0183038f $X=1.585 $Y=2.54 $X2=0 $Y2=0
cc_177 N_B_M1001_g N_VGND_c_506_n 4.64175e-19 $X=2.165 $Y=1.015 $X2=0 $Y2=0
cc_178 N_C_M1009_g N_D_M1008_g 0.0186986f $X=2.655 $Y=2.54 $X2=0 $Y2=0
cc_179 N_C_M1011_g N_D_M1000_g 0.0197345f $X=2.555 $Y=1.015 $X2=0 $Y2=0
cc_180 N_C_c_247_n N_D_M1000_g 0.00334362f $X=2.612 $Y=1.56 $X2=0 $Y2=0
cc_181 N_C_c_248_n N_D_M1000_g 0.0034753f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_182 N_C_c_249_n N_D_M1000_g 0.00131309f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_183 N_C_c_247_n D 4.09211e-19 $X=2.612 $Y=1.56 $X2=0 $Y2=0
cc_184 N_C_c_247_n N_D_c_291_n 0.017484f $X=2.612 $Y=1.56 $X2=0 $Y2=0
cc_185 N_C_c_249_n N_A_229_424#_c_328_n 0.0030474f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_186 N_C_M1011_g N_A_229_424#_c_329_n 0.0110338f $X=2.555 $Y=1.015 $X2=0 $Y2=0
cc_187 N_C_c_249_n N_A_229_424#_c_329_n 0.0149142f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_188 N_C_M1011_g N_A_229_424#_c_331_n 8.15891e-19 $X=2.555 $Y=1.015 $X2=0
+ $Y2=0
cc_189 N_C_M1009_g N_A_229_424#_c_331_n 0.0184715f $X=2.655 $Y=2.54 $X2=0 $Y2=0
cc_190 N_C_c_247_n N_A_229_424#_c_331_n 0.00724776f $X=2.612 $Y=1.56 $X2=0 $Y2=0
cc_191 N_C_c_248_n N_A_229_424#_c_332_n 2.05086e-19 $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_192 N_C_c_249_n N_A_229_424#_c_332_n 0.00154757f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_193 N_C_M1009_g N_A_229_424#_c_338_n 0.00102005f $X=2.655 $Y=2.54 $X2=0 $Y2=0
cc_194 N_C_M1011_g N_A_229_424#_c_375_n 0.00463728f $X=2.555 $Y=1.015 $X2=0
+ $Y2=0
cc_195 N_C_c_248_n N_A_229_424#_c_375_n 5.51222e-19 $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_196 N_C_c_249_n N_A_229_424#_c_375_n 0.00519212f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_197 N_C_M1009_g N_A_229_424#_c_363_n 0.00761391f $X=2.655 $Y=2.54 $X2=0 $Y2=0
cc_198 N_C_c_247_n N_A_229_424#_c_363_n 0.00169415f $X=2.612 $Y=1.56 $X2=0 $Y2=0
cc_199 N_C_M1009_g N_A_229_424#_c_339_n 0.0122449f $X=2.655 $Y=2.54 $X2=0 $Y2=0
cc_200 N_C_M1009_g N_VPWR_c_434_n 0.00460063f $X=2.655 $Y=2.54 $X2=0 $Y2=0
cc_201 N_C_M1009_g N_VPWR_c_431_n 0.00904483f $X=2.655 $Y=2.54 $X2=0 $Y2=0
cc_202 N_C_M1009_g N_VPWR_c_441_n 0.0135446f $X=2.655 $Y=2.54 $X2=0 $Y2=0
cc_203 N_C_c_248_n N_VGND_c_504_n 0.00126694f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_204 N_C_c_249_n N_VGND_c_504_n 0.0130106f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_205 N_C_c_248_n N_VGND_c_506_n 0.00783549f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_206 N_C_c_249_n N_VGND_c_506_n 0.0514254f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_207 N_C_c_248_n N_VGND_c_508_n 0.011167f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_208 N_C_c_249_n N_VGND_c_508_n 0.0291589f $X=2.645 $Y=0.42 $X2=0 $Y2=0
cc_209 N_D_M1008_g N_A_229_424#_M1010_g 0.0217089f $X=3.155 $Y=2.54 $X2=0 $Y2=0
cc_210 D N_A_229_424#_M1010_g 0.00109992f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_211 N_D_c_291_n N_A_229_424#_M1010_g 0.00642675f $X=3.15 $Y=1.715 $X2=0 $Y2=0
cc_212 N_D_M1008_g N_A_229_424#_c_331_n 0.00399192f $X=3.155 $Y=2.54 $X2=0 $Y2=0
cc_213 N_D_M1000_g N_A_229_424#_c_331_n 0.00283662f $X=3.245 $Y=0.92 $X2=0 $Y2=0
cc_214 D N_A_229_424#_c_331_n 0.0204438f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_215 N_D_c_291_n N_A_229_424#_c_331_n 0.00187683f $X=3.15 $Y=1.715 $X2=0 $Y2=0
cc_216 N_D_M1000_g N_A_229_424#_c_332_n 0.021225f $X=3.245 $Y=0.92 $X2=0 $Y2=0
cc_217 D N_A_229_424#_c_332_n 0.032803f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_218 N_D_c_291_n N_A_229_424#_c_332_n 0.00128722f $X=3.15 $Y=1.715 $X2=0 $Y2=0
cc_219 N_D_M1008_g N_A_229_424#_c_338_n 0.0107197f $X=3.155 $Y=2.54 $X2=0 $Y2=0
cc_220 N_D_M1008_g N_A_229_424#_c_339_n 0.00408353f $X=3.155 $Y=2.54 $X2=0 $Y2=0
cc_221 D N_A_229_424#_c_339_n 0.00686439f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_222 N_D_c_291_n N_A_229_424#_c_339_n 5.45701e-19 $X=3.15 $Y=1.715 $X2=0 $Y2=0
cc_223 N_D_M1000_g N_A_229_424#_c_333_n 0.0170787f $X=3.245 $Y=0.92 $X2=0 $Y2=0
cc_224 N_D_M1000_g N_A_229_424#_c_334_n 0.0185769f $X=3.245 $Y=0.92 $X2=0 $Y2=0
cc_225 N_D_M1008_g N_VPWR_c_433_n 0.0124353f $X=3.155 $Y=2.54 $X2=0 $Y2=0
cc_226 N_D_M1008_g N_VPWR_c_434_n 0.005209f $X=3.155 $Y=2.54 $X2=0 $Y2=0
cc_227 N_D_M1008_g N_VPWR_c_431_n 0.00985504f $X=3.155 $Y=2.54 $X2=0 $Y2=0
cc_228 N_D_M1008_g N_VPWR_c_441_n 6.72762e-19 $X=3.155 $Y=2.54 $X2=0 $Y2=0
cc_229 N_D_M1000_g N_X_c_479_n 7.43364e-19 $X=3.245 $Y=0.92 $X2=0 $Y2=0
cc_230 N_D_M1008_g X 0.00112687f $X=3.155 $Y=2.54 $X2=0 $Y2=0
cc_231 D X 8.49268e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_232 N_D_M1000_g N_VGND_c_504_n 0.00462414f $X=3.245 $Y=0.92 $X2=0 $Y2=0
cc_233 N_D_M1000_g N_VGND_c_506_n 0.00428744f $X=3.245 $Y=0.92 $X2=0 $Y2=0
cc_234 N_D_M1000_g N_VGND_c_508_n 0.00476395f $X=3.245 $Y=0.92 $X2=0 $Y2=0
cc_235 N_A_229_424#_c_363_n N_VPWR_M1006_d 0.0280016f $X=2.595 $Y=2.225 $X2=0
+ $Y2=0
cc_236 N_A_229_424#_M1010_g N_VPWR_c_433_n 0.0126713f $X=3.815 $Y=2.4 $X2=0
+ $Y2=0
cc_237 N_A_229_424#_c_332_n N_VPWR_c_433_n 0.00555466f $X=3.535 $Y=1.295 $X2=0
+ $Y2=0
cc_238 N_A_229_424#_c_338_n N_VPWR_c_433_n 0.0375645f $X=2.93 $Y=2.815 $X2=0
+ $Y2=0
cc_239 N_A_229_424#_c_339_n N_VPWR_c_433_n 0.0156416f $X=2.93 $Y=2.265 $X2=0
+ $Y2=0
cc_240 N_A_229_424#_c_333_n N_VPWR_c_433_n 7.25558e-19 $X=3.725 $Y=1.515 $X2=0
+ $Y2=0
cc_241 N_A_229_424#_c_338_n N_VPWR_c_434_n 0.0144686f $X=2.93 $Y=2.815 $X2=0
+ $Y2=0
cc_242 N_A_229_424#_M1010_g N_VPWR_c_437_n 0.005209f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_243 N_A_229_424#_M1010_g N_VPWR_c_431_n 0.00988007f $X=3.815 $Y=2.4 $X2=0
+ $Y2=0
cc_244 N_A_229_424#_c_338_n N_VPWR_c_431_n 0.0119429f $X=2.93 $Y=2.815 $X2=0
+ $Y2=0
cc_245 N_A_229_424#_c_338_n N_VPWR_c_441_n 0.0194969f $X=2.93 $Y=2.815 $X2=0
+ $Y2=0
cc_246 N_A_229_424#_c_363_n N_VPWR_c_441_n 0.0642899f $X=2.595 $Y=2.225 $X2=0
+ $Y2=0
cc_247 N_A_229_424#_c_334_n N_X_c_479_n 0.00609418f $X=3.732 $Y=1.35 $X2=0 $Y2=0
cc_248 N_A_229_424#_c_332_n N_X_c_480_n 0.001126f $X=3.535 $Y=1.295 $X2=0 $Y2=0
cc_249 N_A_229_424#_c_334_n N_X_c_480_n 0.00373327f $X=3.732 $Y=1.35 $X2=0 $Y2=0
cc_250 N_A_229_424#_M1010_g X 0.0043734f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_251 N_A_229_424#_c_332_n X 0.00112338f $X=3.535 $Y=1.295 $X2=0 $Y2=0
cc_252 N_A_229_424#_M1010_g X 0.0136647f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_253 N_A_229_424#_c_332_n N_X_c_481_n 0.0309163f $X=3.535 $Y=1.295 $X2=0 $Y2=0
cc_254 N_A_229_424#_c_333_n N_X_c_481_n 0.0118404f $X=3.725 $Y=1.515 $X2=0 $Y2=0
cc_255 N_A_229_424#_c_334_n N_X_c_481_n 0.00255066f $X=3.732 $Y=1.35 $X2=0 $Y2=0
cc_256 N_A_229_424#_c_332_n N_VGND_M1000_d 0.00339782f $X=3.535 $Y=1.295 $X2=0
+ $Y2=0
cc_257 N_A_229_424#_c_328_n N_VGND_c_503_n 0.00343679f $X=1.475 $Y=0.765 $X2=0
+ $Y2=0
cc_258 N_A_229_424#_c_332_n N_VGND_c_504_n 0.026684f $X=3.535 $Y=1.295 $X2=0
+ $Y2=0
cc_259 N_A_229_424#_c_333_n N_VGND_c_504_n 7.86248e-19 $X=3.725 $Y=1.515 $X2=0
+ $Y2=0
cc_260 N_A_229_424#_c_334_n N_VGND_c_504_n 0.00807563f $X=3.732 $Y=1.35 $X2=0
+ $Y2=0
cc_261 N_A_229_424#_c_328_n N_VGND_c_506_n 0.00707634f $X=1.475 $Y=0.765 $X2=0
+ $Y2=0
cc_262 N_A_229_424#_c_334_n N_VGND_c_507_n 0.00467453f $X=3.732 $Y=1.35 $X2=0
+ $Y2=0
cc_263 N_A_229_424#_c_328_n N_VGND_c_508_n 0.0101843f $X=1.475 $Y=0.765 $X2=0
+ $Y2=0
cc_264 N_A_229_424#_c_334_n N_VGND_c_508_n 0.00505379f $X=3.732 $Y=1.35 $X2=0
+ $Y2=0
cc_265 N_A_229_424#_c_329_n A_353_124# 0.00805082f $X=2.595 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_266 N_A_229_424#_c_329_n A_448_139# 0.00237138f $X=2.595 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_267 N_A_229_424#_c_332_n A_526_139# 0.0125125f $X=3.535 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_268 N_A_229_424#_c_375_n A_526_139# 0.00134898f $X=2.68 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_269 N_VPWR_c_433_n X 0.0584079f $X=3.5 $Y=2.265 $X2=0 $Y2=0
cc_270 N_VPWR_c_437_n X 0.0156645f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_271 N_VPWR_c_431_n X 0.0128976f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_272 N_X_c_479_n N_VGND_c_504_n 0.0220013f $X=4.04 $Y=0.645 $X2=0 $Y2=0
cc_273 N_X_c_479_n N_VGND_c_507_n 0.0102463f $X=4.04 $Y=0.645 $X2=0 $Y2=0
cc_274 N_X_c_479_n N_VGND_c_508_n 0.0119585f $X=4.04 $Y=0.645 $X2=0 $Y2=0

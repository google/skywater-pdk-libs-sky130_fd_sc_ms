* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 VPWR a_110_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 a_762_368# A2 a_1216_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X2 VPWR a_110_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 a_110_48# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X4 VGND A3 a_523_124# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 a_854_368# A4 a_110_48# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X6 VGND a_110_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_523_124# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_523_124# A4 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 VGND A2 a_523_124# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X10 a_110_48# A4 a_854_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X11 VGND A1 a_523_124# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X12 a_523_124# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 a_854_368# A3 a_762_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X14 X a_110_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 X a_110_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 X a_110_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X17 VPWR B1 a_110_48# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X18 a_1216_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X19 X a_110_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X20 VPWR A1 a_1216_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X21 a_762_368# A3 a_854_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X22 a_523_124# B1 a_110_48# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X23 a_110_48# B1 a_523_124# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X24 VGND A4 a_523_124# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X25 a_523_124# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X26 a_1216_368# A2 a_762_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X27 VGND a_110_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

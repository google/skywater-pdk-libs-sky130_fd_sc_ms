# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__dfbbp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__dfbbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.96000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.960000 1.825000 2.290000 2.155000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.502200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.525000 0.350000 12.860000 2.980000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.502100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.065000 0.350000 11.460000 1.130000 ;
        RECT 11.120000 1.820000 11.460000 2.980000 ;
        RECT 11.290000 1.130000 11.460000 1.820000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.235000 0.980000 10.580000 1.650000 ;
    END
  END RESET_B
  PIN SET_B
    ANTENNAGATEAREA  0.524700 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.230000 1.410000 4.560000 1.655000 ;
        RECT 4.360000 1.655000 4.530000 2.905000 ;
        RECT 4.360000 2.905000 5.330000 3.075000 ;
        RECT 5.160000 2.165000 6.210000 2.335000 ;
        RECT 5.160000 2.335000 5.330000 2.905000 ;
        RECT 6.040000 2.335000 6.210000 2.905000 ;
        RECT 6.040000 2.905000 7.450000 3.075000 ;
        RECT 7.280000 1.740000 8.570000 1.800000 ;
        RECT 7.280000 1.800000 8.515000 1.910000 ;
        RECT 7.280000 1.910000 7.450000 2.905000 ;
        RECT 8.240000 1.470000 8.570000 1.740000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.180000 0.805000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.960000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.960000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.960000 0.085000 ;
      RECT  0.000000  3.245000 12.960000 3.415000 ;
      RECT  0.085000  0.350000  0.445000 1.010000 ;
      RECT  0.085000  1.010000  0.255000 1.720000 ;
      RECT  0.085000  1.720000  1.145000 1.890000 ;
      RECT  0.085000  1.890000  0.535000 2.980000 ;
      RECT  0.615000  0.085000  0.945000 1.010000 ;
      RECT  0.705000  2.060000  1.035000 3.245000 ;
      RECT  0.975000  1.300000  1.145000 1.720000 ;
      RECT  1.125000  0.350000  1.485000 1.130000 ;
      RECT  1.315000  1.130000  1.485000 1.255000 ;
      RECT  1.315000  1.255000  2.615000 1.585000 ;
      RECT  1.315000  1.585000  1.565000 2.980000 ;
      RECT  1.655000  0.085000  1.905000 1.065000 ;
      RECT  1.805000  2.425000  2.410000 3.245000 ;
      RECT  2.085000  0.605000  2.335000 0.915000 ;
      RECT  2.085000  0.915000  2.955000 1.085000 ;
      RECT  2.575000  0.415000  3.295000 0.745000 ;
      RECT  2.580000  2.295000  2.955000 2.755000 ;
      RECT  2.785000  1.085000  2.955000 2.295000 ;
      RECT  3.125000  0.745000  3.295000 1.625000 ;
      RECT  3.125000  1.625000  4.060000 1.795000 ;
      RECT  3.125000  1.795000  3.430000 2.335000 ;
      RECT  3.465000  0.730000  5.335000 0.840000 ;
      RECT  3.465000  0.840000  6.020000 0.900000 ;
      RECT  3.465000  0.900000  3.720000 1.455000 ;
      RECT  3.560000  0.085000  4.155000 0.560000 ;
      RECT  3.890000  1.070000  4.915000 1.240000 ;
      RECT  3.890000  1.240000  4.060000 1.625000 ;
      RECT  3.940000  1.965000  4.190000 3.245000 ;
      RECT  4.415000  0.255000  5.840000 0.425000 ;
      RECT  4.415000  0.425000  4.825000 0.560000 ;
      RECT  4.700000  1.825000  6.020000 1.995000 ;
      RECT  4.700000  1.995000  4.950000 2.735000 ;
      RECT  4.745000  1.240000  4.915000 1.255000 ;
      RECT  4.745000  1.255000  5.100000 1.585000 ;
      RECT  5.015000  0.595000  5.335000 0.730000 ;
      RECT  5.085000  0.900000  6.020000 1.010000 ;
      RECT  5.310000  1.180000  5.640000 1.585000 ;
      RECT  5.500000  2.505000  5.870000 3.245000 ;
      RECT  5.510000  0.425000  5.840000 0.670000 ;
      RECT  5.850000  1.010000  6.020000 1.255000 ;
      RECT  5.850000  1.255000  6.180000 1.585000 ;
      RECT  5.850000  1.585000  6.020000 1.825000 ;
      RECT  6.060000  0.085000  6.430000 0.670000 ;
      RECT  6.190000  0.670000  6.430000 1.085000 ;
      RECT  6.440000  1.610000  6.770000 1.940000 ;
      RECT  6.540000  2.110000  7.110000 2.280000 ;
      RECT  6.540000  2.280000  6.870000 2.735000 ;
      RECT  6.600000  0.255000  7.670000 0.425000 ;
      RECT  6.600000  0.425000  6.770000 1.610000 ;
      RECT  6.940000  0.595000  7.175000 1.400000 ;
      RECT  6.940000  1.400000  8.070000 1.570000 ;
      RECT  6.940000  1.570000  7.110000 2.110000 ;
      RECT  7.345000  0.425000  7.670000 1.230000 ;
      RECT  7.620000  2.080000  9.385000 2.240000 ;
      RECT  7.620000  2.240000 10.950000 2.380000 ;
      RECT  7.620000  2.650000  8.420000 3.245000 ;
      RECT  7.900000  1.130000  9.045000 1.300000 ;
      RECT  7.900000  1.300000  8.070000 1.400000 ;
      RECT  8.085000  0.085000  8.415000 0.960000 ;
      RECT  8.585000  0.255000  9.725000 0.425000 ;
      RECT  8.585000  0.425000  8.915000 0.960000 ;
      RECT  8.685000  1.970000  9.385000 2.080000 ;
      RECT  8.685000  2.380000 10.950000 2.410000 ;
      RECT  8.685000  2.410000  8.935000 2.980000 ;
      RECT  8.780000  1.300000  9.045000 1.550000 ;
      RECT  9.085000  0.595000  9.385000 0.960000 ;
      RECT  9.215000  0.960000  9.385000 1.970000 ;
      RECT  9.470000  2.580000  9.800000 3.245000 ;
      RECT  9.555000  0.425000  9.725000 1.020000 ;
      RECT  9.710000  1.190000 10.065000 1.820000 ;
      RECT  9.710000  1.820000 10.405000 2.070000 ;
      RECT  9.895000  0.350000 10.385000 0.810000 ;
      RECT  9.895000  0.810000 10.065000 1.190000 ;
      RECT 10.565000  0.085000 10.895000 0.810000 ;
      RECT 10.590000  2.580000 10.920000 3.245000 ;
      RECT 10.780000  1.320000 11.120000 1.650000 ;
      RECT 10.780000  1.650000 10.950000 2.240000 ;
      RECT 11.640000  0.350000 11.875000 1.255000 ;
      RECT 11.640000  1.255000 12.355000 1.585000 ;
      RECT 11.640000  1.585000 11.810000 2.030000 ;
      RECT 11.640000  2.030000 11.890000 2.910000 ;
      RECT 12.055000  0.085000 12.305000 0.810000 ;
      RECT 12.075000  1.820000 12.325000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.210000  5.605000 1.380000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  1.210000  9.925000 1.380000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
    LAYER met1 ;
      RECT 5.375000 1.180000 5.665000 1.225000 ;
      RECT 5.375000 1.225000 9.985000 1.365000 ;
      RECT 5.375000 1.365000 5.665000 1.410000 ;
      RECT 9.695000 1.180000 9.985000 1.225000 ;
      RECT 9.695000 1.365000 9.985000 1.410000 ;
  END
END sky130_fd_sc_ms__dfbbp_1
END LIBRARY

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfstp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
X0 a_1804_424# a_795_74# a_2144_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X1 a_293_464# a_27_74# a_419_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X2 VGND a_2611_98# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_209_464# D a_293_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X4 a_608_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 a_239_74# D a_293_464# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X6 a_1804_424# a_608_74# a_2141_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X7 a_419_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X8 VGND a_608_74# a_795_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 VPWR a_2611_98# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X10 a_1185_55# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X11 a_1587_379# a_608_74# a_1804_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X12 a_27_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X13 VPWR SET_B a_1804_424# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X14 a_1641_74# a_795_74# a_1804_424# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 a_2219_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X16 a_293_464# SCE a_403_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X17 a_608_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 a_1641_74# a_991_81# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X19 a_293_464# a_608_74# a_991_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X20 a_2141_74# a_2186_367# a_2219_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X21 VGND a_27_74# a_239_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X22 a_1587_379# a_991_81# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X23 a_2186_367# a_1804_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X24 a_2611_98# a_1804_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X25 a_293_464# a_795_74# a_991_81# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X26 a_403_74# SCD VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X27 a_1804_424# a_795_74# a_1641_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X28 VPWR a_608_74# a_795_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X29 a_1804_424# a_608_74# a_1587_379# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X30 Q a_2611_98# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X31 a_1429_74# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X32 a_2144_508# a_2186_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X33 VGND a_991_81# a_1641_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X34 VPWR a_991_81# a_1185_55# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X35 a_1185_55# a_991_81# a_1429_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X36 a_1120_483# a_1185_55# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X37 VGND a_1804_424# a_2186_367# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X38 a_991_81# a_608_74# a_1120_483# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X39 a_991_81# a_795_74# a_1143_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X40 a_27_74# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X41 VPWR a_991_81# a_1587_379# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X42 a_2611_98# a_1804_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X43 VPWR SCE a_209_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X44 a_1143_81# a_1185_55# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X45 Q a_2611_98# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

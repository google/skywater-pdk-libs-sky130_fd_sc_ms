* File: sky130_fd_sc_ms__or4_1.pxi.spice
* Created: Fri Aug 28 18:08:47 2020
* 
x_PM_SKY130_FD_SC_MS__OR4_1%D N_D_M1003_g N_D_c_63_n N_D_M1001_g D N_D_c_64_n
+ PM_SKY130_FD_SC_MS__OR4_1%D
x_PM_SKY130_FD_SC_MS__OR4_1%C N_C_M1002_g N_C_M1008_g C N_C_c_91_n
+ PM_SKY130_FD_SC_MS__OR4_1%C
x_PM_SKY130_FD_SC_MS__OR4_1%B N_B_M1005_g N_B_M1006_g B N_B_c_124_n
+ PM_SKY130_FD_SC_MS__OR4_1%B
x_PM_SKY130_FD_SC_MS__OR4_1%A N_A_M1009_g N_A_M1004_g A N_A_c_156_n N_A_c_157_n
+ PM_SKY130_FD_SC_MS__OR4_1%A
x_PM_SKY130_FD_SC_MS__OR4_1%A_44_392# N_A_44_392#_M1003_d N_A_44_392#_M1006_d
+ N_A_44_392#_M1001_s N_A_44_392#_M1000_g N_A_44_392#_M1007_g
+ N_A_44_392#_c_207_n N_A_44_392#_c_208_n N_A_44_392#_c_209_n
+ N_A_44_392#_c_197_n N_A_44_392#_c_198_n N_A_44_392#_c_199_n
+ N_A_44_392#_c_200_n N_A_44_392#_c_201_n N_A_44_392#_c_202_n
+ N_A_44_392#_c_203_n N_A_44_392#_c_204_n N_A_44_392#_c_205_n
+ PM_SKY130_FD_SC_MS__OR4_1%A_44_392#
x_PM_SKY130_FD_SC_MS__OR4_1%VPWR N_VPWR_M1009_d N_VPWR_c_301_n VPWR
+ N_VPWR_c_302_n N_VPWR_c_303_n N_VPWR_c_300_n N_VPWR_c_305_n
+ PM_SKY130_FD_SC_MS__OR4_1%VPWR
x_PM_SKY130_FD_SC_MS__OR4_1%X N_X_M1007_d N_X_M1000_d N_X_c_327_n N_X_c_328_n X
+ X X X N_X_c_329_n PM_SKY130_FD_SC_MS__OR4_1%X
x_PM_SKY130_FD_SC_MS__OR4_1%VGND N_VGND_M1003_s N_VGND_M1002_d N_VGND_M1004_d
+ N_VGND_c_351_n N_VGND_c_352_n N_VGND_c_353_n N_VGND_c_354_n N_VGND_c_355_n
+ VGND N_VGND_c_356_n N_VGND_c_357_n N_VGND_c_358_n N_VGND_c_359_n
+ N_VGND_c_360_n PM_SKY130_FD_SC_MS__OR4_1%VGND
cc_1 VNB N_D_M1003_g 0.0360698f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.835
cc_2 VNB N_D_c_63_n 0.0241911f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.84
cc_3 VNB N_D_c_64_n 0.0135797f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.585
cc_4 VNB N_C_M1002_g 0.0312133f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.835
cc_5 VNB C 0.00378948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_C_c_91_n 0.0188753f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.585
cc_7 VNB N_B_M1006_g 0.0332829f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.46
cc_8 VNB B 0.00187616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B_c_124_n 0.0220243f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.585
cc_10 VNB N_A_M1004_g 0.0262449f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.46
cc_11 VNB N_A_c_156_n 0.00426371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_c_157_n 0.0252457f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.6
cc_13 VNB N_A_44_392#_M1000_g 0.00183668f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.585
cc_14 VNB N_A_44_392#_M1007_g 0.0287893f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.6
cc_15 VNB N_A_44_392#_c_197_n 0.00325236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_44_392#_c_198_n 0.0116367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_44_392#_c_199_n 0.0102551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_44_392#_c_200_n 0.00430793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_44_392#_c_201_n 0.00595784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_44_392#_c_202_n 0.0103286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_44_392#_c_203_n 3.93303e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_44_392#_c_204_n 0.00857761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_44_392#_c_205_n 0.0337537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_300_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_X_c_327_n 0.0279492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_X_c_328_n 0.012405f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.6
cc_27 VNB N_X_c_329_n 0.0247746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_351_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.585
cc_29 VNB N_VGND_c_352_n 0.0551753f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.585
cc_30 VNB N_VGND_c_353_n 0.0198125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_354_n 0.0288416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_355_n 0.0135712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_356_n 0.0252222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_357_n 0.0179969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_358_n 0.222079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_359_n 0.00913651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_360_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_D_c_63_n 0.0465435f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.84
cc_39 VPB N_D_c_64_n 0.0110488f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=1.585
cc_40 VPB N_C_M1008_g 0.0259174f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=2.46
cc_41 VPB C 0.00345409f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_C_c_91_n 0.00964655f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=1.585
cc_43 VPB N_B_M1005_g 0.0279229f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.835
cc_44 VPB B 0.00159046f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_B_c_124_n 0.0106136f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=1.585
cc_46 VPB N_A_M1009_g 0.0311121f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.835
cc_47 VPB N_A_c_156_n 0.00302988f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_c_157_n 0.00580281f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=1.6
cc_49 VPB N_A_44_392#_M1000_g 0.0311419f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=1.585
cc_50 VPB N_A_44_392#_c_207_n 0.00933413f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A_44_392#_c_208_n 0.0352562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_A_44_392#_c_209_n 0.0297607f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_44_392#_c_203_n 0.00298265f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_301_n 0.00684033f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=2.46
cc_55 VPB N_VPWR_c_302_n 0.0678403f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=1.585
cc_56 VPB N_VPWR_c_303_n 0.0245279f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_300_n 0.101532f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_305_n 0.00766803f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB X 0.0145515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB X 0.0421222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_X_c_329_n 0.00758261f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 N_D_M1003_g N_C_M1002_g 0.027997f $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_63 N_D_c_63_n N_C_M1008_g 0.075055f $X=0.59 $Y=1.84 $X2=0 $Y2=0
cc_64 N_D_c_63_n C 5.19548e-19 $X=0.59 $Y=1.84 $X2=0 $Y2=0
cc_65 N_D_c_64_n C 0.0195329f $X=0.485 $Y=1.585 $X2=0 $Y2=0
cc_66 N_D_c_63_n N_C_c_91_n 0.0156908f $X=0.59 $Y=1.84 $X2=0 $Y2=0
cc_67 N_D_c_64_n N_C_c_91_n 4.21003e-19 $X=0.485 $Y=1.585 $X2=0 $Y2=0
cc_68 N_D_c_63_n N_A_44_392#_c_207_n 0.00239488f $X=0.59 $Y=1.84 $X2=0 $Y2=0
cc_69 N_D_c_64_n N_A_44_392#_c_207_n 0.0291116f $X=0.485 $Y=1.585 $X2=0 $Y2=0
cc_70 N_D_c_63_n N_A_44_392#_c_208_n 0.0166884f $X=0.59 $Y=1.84 $X2=0 $Y2=0
cc_71 N_D_c_63_n N_A_44_392#_c_209_n 0.0134609f $X=0.59 $Y=1.84 $X2=0 $Y2=0
cc_72 N_D_c_64_n N_A_44_392#_c_209_n 0.00859598f $X=0.485 $Y=1.585 $X2=0 $Y2=0
cc_73 N_D_M1003_g N_A_44_392#_c_197_n 0.0065178f $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_74 N_D_M1003_g N_A_44_392#_c_199_n 0.00581878f $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_75 N_D_c_63_n N_A_44_392#_c_199_n 0.00120428f $X=0.59 $Y=1.84 $X2=0 $Y2=0
cc_76 N_D_c_64_n N_A_44_392#_c_199_n 0.00216782f $X=0.485 $Y=1.585 $X2=0 $Y2=0
cc_77 N_D_c_63_n N_VPWR_c_302_n 0.005209f $X=0.59 $Y=1.84 $X2=0 $Y2=0
cc_78 N_D_c_63_n N_VPWR_c_300_n 0.00987183f $X=0.59 $Y=1.84 $X2=0 $Y2=0
cc_79 N_D_M1003_g N_VGND_c_352_n 0.00867578f $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_80 N_D_c_63_n N_VGND_c_352_n 0.0026975f $X=0.59 $Y=1.84 $X2=0 $Y2=0
cc_81 N_D_c_64_n N_VGND_c_352_n 0.0190298f $X=0.485 $Y=1.585 $X2=0 $Y2=0
cc_82 N_D_M1003_g N_VGND_c_353_n 0.0043356f $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_83 N_D_M1003_g N_VGND_c_358_n 0.00487769f $X=0.565 $Y=0.835 $X2=0 $Y2=0
cc_84 N_C_M1008_g N_B_M1005_g 0.0497644f $X=1.01 $Y=2.46 $X2=0 $Y2=0
cc_85 N_C_M1002_g N_B_M1006_g 0.0175401f $X=0.995 $Y=0.835 $X2=0 $Y2=0
cc_86 C B 0.0259046f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_87 N_C_c_91_n B 3.84189e-19 $X=1.085 $Y=1.585 $X2=0 $Y2=0
cc_88 C N_B_c_124_n 0.0022324f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_89 N_C_c_91_n N_B_c_124_n 0.0174741f $X=1.085 $Y=1.585 $X2=0 $Y2=0
cc_90 N_C_M1008_g N_A_44_392#_c_208_n 0.00412931f $X=1.01 $Y=2.46 $X2=0 $Y2=0
cc_91 N_C_M1008_g N_A_44_392#_c_209_n 0.0175218f $X=1.01 $Y=2.46 $X2=0 $Y2=0
cc_92 C N_A_44_392#_c_209_n 0.028511f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_93 N_C_c_91_n N_A_44_392#_c_209_n 9.72837e-19 $X=1.085 $Y=1.585 $X2=0 $Y2=0
cc_94 N_C_M1002_g N_A_44_392#_c_197_n 0.0121196f $X=0.995 $Y=0.835 $X2=0 $Y2=0
cc_95 N_C_M1002_g N_A_44_392#_c_198_n 0.0124559f $X=0.995 $Y=0.835 $X2=0 $Y2=0
cc_96 C N_A_44_392#_c_198_n 0.0201443f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_97 N_C_c_91_n N_A_44_392#_c_198_n 0.00395915f $X=1.085 $Y=1.585 $X2=0 $Y2=0
cc_98 N_C_M1002_g N_A_44_392#_c_199_n 0.00256575f $X=0.995 $Y=0.835 $X2=0 $Y2=0
cc_99 C N_A_44_392#_c_199_n 0.00151542f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_100 N_C_M1008_g N_VPWR_c_302_n 0.00553757f $X=1.01 $Y=2.46 $X2=0 $Y2=0
cc_101 N_C_M1008_g N_VPWR_c_300_n 0.0109071f $X=1.01 $Y=2.46 $X2=0 $Y2=0
cc_102 N_C_M1002_g N_VGND_c_353_n 0.0043356f $X=0.995 $Y=0.835 $X2=0 $Y2=0
cc_103 N_C_M1002_g N_VGND_c_354_n 0.00598528f $X=0.995 $Y=0.835 $X2=0 $Y2=0
cc_104 N_C_M1002_g N_VGND_c_358_n 0.00487769f $X=0.995 $Y=0.835 $X2=0 $Y2=0
cc_105 N_B_M1005_g N_A_M1009_g 0.0454169f $X=1.58 $Y=2.46 $X2=0 $Y2=0
cc_106 N_B_M1006_g N_A_M1004_g 0.0208052f $X=1.73 $Y=0.835 $X2=0 $Y2=0
cc_107 N_B_M1006_g N_A_c_156_n 0.00151003f $X=1.73 $Y=0.835 $X2=0 $Y2=0
cc_108 B N_A_c_156_n 0.0233207f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_109 N_B_c_124_n N_A_c_156_n 0.00202099f $X=1.655 $Y=1.585 $X2=0 $Y2=0
cc_110 N_B_M1006_g N_A_c_157_n 0.00324793f $X=1.73 $Y=0.835 $X2=0 $Y2=0
cc_111 B N_A_c_157_n 4.10732e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_112 N_B_c_124_n N_A_c_157_n 0.0175264f $X=1.655 $Y=1.585 $X2=0 $Y2=0
cc_113 N_B_M1005_g N_A_44_392#_c_209_n 0.0182755f $X=1.58 $Y=2.46 $X2=0 $Y2=0
cc_114 B N_A_44_392#_c_209_n 0.0248886f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_115 N_B_c_124_n N_A_44_392#_c_209_n 9.53139e-19 $X=1.655 $Y=1.585 $X2=0 $Y2=0
cc_116 N_B_M1006_g N_A_44_392#_c_198_n 0.0171248f $X=1.73 $Y=0.835 $X2=0 $Y2=0
cc_117 B N_A_44_392#_c_198_n 0.0186612f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_118 N_B_c_124_n N_A_44_392#_c_198_n 0.00115436f $X=1.655 $Y=1.585 $X2=0 $Y2=0
cc_119 N_B_M1006_g N_A_44_392#_c_200_n 0.00299671f $X=1.73 $Y=0.835 $X2=0 $Y2=0
cc_120 N_B_M1005_g N_VPWR_c_301_n 0.00402353f $X=1.58 $Y=2.46 $X2=0 $Y2=0
cc_121 N_B_M1005_g N_VPWR_c_302_n 0.00553757f $X=1.58 $Y=2.46 $X2=0 $Y2=0
cc_122 N_B_M1005_g N_VPWR_c_300_n 0.0109203f $X=1.58 $Y=2.46 $X2=0 $Y2=0
cc_123 N_B_M1006_g N_VGND_c_354_n 0.00601282f $X=1.73 $Y=0.835 $X2=0 $Y2=0
cc_124 N_B_M1006_g N_VGND_c_356_n 0.00451272f $X=1.73 $Y=0.835 $X2=0 $Y2=0
cc_125 N_B_M1006_g N_VGND_c_358_n 0.00487769f $X=1.73 $Y=0.835 $X2=0 $Y2=0
cc_126 N_A_M1009_g N_A_44_392#_M1000_g 0.0183184f $X=2.15 $Y=2.46 $X2=0 $Y2=0
cc_127 N_A_c_157_n N_A_44_392#_M1000_g 0.00133909f $X=2.32 $Y=1.515 $X2=0 $Y2=0
cc_128 N_A_M1004_g N_A_44_392#_M1007_g 0.0183187f $X=2.32 $Y=0.835 $X2=0 $Y2=0
cc_129 N_A_M1009_g N_A_44_392#_c_209_n 0.0159386f $X=2.15 $Y=2.46 $X2=0 $Y2=0
cc_130 N_A_c_156_n N_A_44_392#_c_209_n 0.0264603f $X=2.225 $Y=1.515 $X2=0 $Y2=0
cc_131 N_A_c_157_n N_A_44_392#_c_209_n 0.0010246f $X=2.32 $Y=1.515 $X2=0 $Y2=0
cc_132 N_A_M1004_g N_A_44_392#_c_200_n 0.00299671f $X=2.32 $Y=0.835 $X2=0 $Y2=0
cc_133 N_A_M1004_g N_A_44_392#_c_201_n 0.0158031f $X=2.32 $Y=0.835 $X2=0 $Y2=0
cc_134 N_A_c_156_n N_A_44_392#_c_201_n 0.0147621f $X=2.225 $Y=1.515 $X2=0 $Y2=0
cc_135 N_A_c_157_n N_A_44_392#_c_201_n 3.80832e-19 $X=2.32 $Y=1.515 $X2=0 $Y2=0
cc_136 N_A_M1004_g N_A_44_392#_c_202_n 0.00539948f $X=2.32 $Y=0.835 $X2=0 $Y2=0
cc_137 N_A_c_156_n N_A_44_392#_c_202_n 0.0225675f $X=2.225 $Y=1.515 $X2=0 $Y2=0
cc_138 N_A_M1009_g N_A_44_392#_c_203_n 0.00351106f $X=2.15 $Y=2.46 $X2=0 $Y2=0
cc_139 N_A_c_156_n N_A_44_392#_c_203_n 0.0116888f $X=2.225 $Y=1.515 $X2=0 $Y2=0
cc_140 N_A_c_157_n N_A_44_392#_c_203_n 3.58193e-19 $X=2.32 $Y=1.515 $X2=0 $Y2=0
cc_141 N_A_c_156_n N_A_44_392#_c_204_n 0.0124267f $X=2.225 $Y=1.515 $X2=0 $Y2=0
cc_142 N_A_c_157_n N_A_44_392#_c_204_n 0.00100627f $X=2.32 $Y=1.515 $X2=0 $Y2=0
cc_143 N_A_M1004_g N_A_44_392#_c_205_n 0.0204349f $X=2.32 $Y=0.835 $X2=0 $Y2=0
cc_144 N_A_c_156_n N_A_44_392#_c_205_n 3.1599e-19 $X=2.225 $Y=1.515 $X2=0 $Y2=0
cc_145 N_A_M1009_g N_VPWR_c_301_n 0.0256718f $X=2.15 $Y=2.46 $X2=0 $Y2=0
cc_146 N_A_M1009_g N_VPWR_c_302_n 0.00275477f $X=2.15 $Y=2.46 $X2=0 $Y2=0
cc_147 N_A_M1009_g N_VPWR_c_300_n 0.00548615f $X=2.15 $Y=2.46 $X2=0 $Y2=0
cc_148 N_A_M1009_g X 8.59913e-19 $X=2.15 $Y=2.46 $X2=0 $Y2=0
cc_149 N_A_M1004_g N_VGND_c_355_n 0.00475377f $X=2.32 $Y=0.835 $X2=0 $Y2=0
cc_150 N_A_M1004_g N_VGND_c_356_n 0.00451272f $X=2.32 $Y=0.835 $X2=0 $Y2=0
cc_151 N_A_M1004_g N_VGND_c_358_n 0.00487769f $X=2.32 $Y=0.835 $X2=0 $Y2=0
cc_152 N_A_44_392#_c_209_n A_136_392# 0.0048076f $X=2.56 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_153 N_A_44_392#_c_209_n A_220_392# 0.010795f $X=2.56 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_154 N_A_44_392#_c_209_n A_334_392# 0.010795f $X=2.56 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_155 N_A_44_392#_c_209_n N_VPWR_M1009_d 0.013495f $X=2.56 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_156 N_A_44_392#_c_203_n N_VPWR_M1009_d 0.00221445f $X=2.645 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_157 N_A_44_392#_M1000_g N_VPWR_c_301_n 0.0101173f $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_158 N_A_44_392#_c_209_n N_VPWR_c_301_n 0.0280983f $X=2.56 $Y=2.035 $X2=0
+ $Y2=0
cc_159 N_A_44_392#_c_208_n N_VPWR_c_302_n 0.014549f $X=0.365 $Y=2.815 $X2=0
+ $Y2=0
cc_160 N_A_44_392#_M1000_g N_VPWR_c_303_n 0.005209f $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_161 N_A_44_392#_M1000_g N_VPWR_c_300_n 0.00989122f $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_162 N_A_44_392#_c_208_n N_VPWR_c_300_n 0.0119743f $X=0.365 $Y=2.815 $X2=0
+ $Y2=0
cc_163 N_A_44_392#_M1007_g N_X_c_327_n 0.00205928f $X=2.83 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A_44_392#_c_202_n N_X_c_328_n 0.00135284f $X=2.645 $Y=1.63 $X2=0 $Y2=0
cc_165 N_A_44_392#_M1000_g X 0.00298246f $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_166 N_A_44_392#_c_202_n X 0.00251595f $X=2.645 $Y=1.63 $X2=0 $Y2=0
cc_167 N_A_44_392#_c_203_n X 0.00568911f $X=2.645 $Y=1.95 $X2=0 $Y2=0
cc_168 N_A_44_392#_M1000_g X 0.0175931f $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_169 N_A_44_392#_M1000_g N_X_c_329_n 0.00305218f $X=2.84 $Y=2.4 $X2=0 $Y2=0
cc_170 N_A_44_392#_M1007_g N_X_c_329_n 0.00244983f $X=2.83 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A_44_392#_c_202_n N_X_c_329_n 0.0303927f $X=2.645 $Y=1.63 $X2=0 $Y2=0
cc_172 N_A_44_392#_c_203_n N_X_c_329_n 0.0060551f $X=2.645 $Y=1.95 $X2=0 $Y2=0
cc_173 N_A_44_392#_c_205_n N_X_c_329_n 0.00232633f $X=2.77 $Y=1.465 $X2=0 $Y2=0
cc_174 N_A_44_392#_c_198_n N_VGND_M1002_d 0.00623975f $X=1.86 $Y=1.095 $X2=0
+ $Y2=0
cc_175 N_A_44_392#_c_201_n N_VGND_M1004_d 0.00113743f $X=2.56 $Y=1.095 $X2=0
+ $Y2=0
cc_176 N_A_44_392#_c_202_n N_VGND_M1004_d 0.00214042f $X=2.645 $Y=1.63 $X2=0
+ $Y2=0
cc_177 N_A_44_392#_c_197_n N_VGND_c_352_n 0.0183885f $X=0.78 $Y=0.835 $X2=0
+ $Y2=0
cc_178 N_A_44_392#_c_199_n N_VGND_c_352_n 0.00584871f $X=0.945 $Y=1.095 $X2=0
+ $Y2=0
cc_179 N_A_44_392#_c_197_n N_VGND_c_353_n 0.00805448f $X=0.78 $Y=0.835 $X2=0
+ $Y2=0
cc_180 N_A_44_392#_c_197_n N_VGND_c_354_n 0.0115546f $X=0.78 $Y=0.835 $X2=0
+ $Y2=0
cc_181 N_A_44_392#_c_198_n N_VGND_c_354_n 0.0383199f $X=1.86 $Y=1.095 $X2=0
+ $Y2=0
cc_182 N_A_44_392#_c_200_n N_VGND_c_354_n 0.00120817f $X=2.025 $Y=0.835 $X2=0
+ $Y2=0
cc_183 N_A_44_392#_M1007_g N_VGND_c_355_n 0.0155432f $X=2.83 $Y=0.74 $X2=0 $Y2=0
cc_184 N_A_44_392#_c_200_n N_VGND_c_355_n 0.00117493f $X=2.025 $Y=0.835 $X2=0
+ $Y2=0
cc_185 N_A_44_392#_c_201_n N_VGND_c_355_n 0.00875025f $X=2.56 $Y=1.095 $X2=0
+ $Y2=0
cc_186 N_A_44_392#_c_202_n N_VGND_c_355_n 0.0136978f $X=2.645 $Y=1.63 $X2=0
+ $Y2=0
cc_187 N_A_44_392#_c_205_n N_VGND_c_355_n 4.70665e-19 $X=2.77 $Y=1.465 $X2=0
+ $Y2=0
cc_188 N_A_44_392#_c_200_n N_VGND_c_356_n 0.00817062f $X=2.025 $Y=0.835 $X2=0
+ $Y2=0
cc_189 N_A_44_392#_M1007_g N_VGND_c_357_n 0.00383152f $X=2.83 $Y=0.74 $X2=0
+ $Y2=0
cc_190 N_A_44_392#_M1007_g N_VGND_c_358_n 0.00761312f $X=2.83 $Y=0.74 $X2=0
+ $Y2=0
cc_191 N_A_44_392#_c_197_n N_VGND_c_358_n 0.0105848f $X=0.78 $Y=0.835 $X2=0
+ $Y2=0
cc_192 N_A_44_392#_c_200_n N_VGND_c_358_n 0.010638f $X=2.025 $Y=0.835 $X2=0
+ $Y2=0
cc_193 N_VPWR_c_301_n X 0.0327485f $X=2.375 $Y=2.455 $X2=0 $Y2=0
cc_194 N_VPWR_c_303_n X 0.0165569f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_195 N_VPWR_c_300_n X 0.0136363f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_196 N_X_c_327_n N_VGND_c_355_n 0.0183161f $X=3.045 $Y=0.515 $X2=0 $Y2=0
cc_197 N_X_c_327_n N_VGND_c_357_n 0.0139663f $X=3.045 $Y=0.515 $X2=0 $Y2=0
cc_198 N_X_c_327_n N_VGND_c_358_n 0.0115601f $X=3.045 $Y=0.515 $X2=0 $Y2=0

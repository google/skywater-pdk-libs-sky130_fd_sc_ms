* File: sky130_fd_sc_ms__a21o_4.pex.spice
* Created: Fri Aug 28 16:59:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A21O_4%A_91_48# 1 2 3 12 16 20 24 28 32 36 40 42 52
+ 54 55 58 60 64 67 77
c131 77 0 1.33616e-19 $X=1.895 $Y=1.465
c132 64 0 1.83628e-19 $X=4.055 $Y=0.76
c133 60 0 1.66816e-20 $X=3.96 $Y=1.195
c134 58 0 5.66563e-20 $X=3.09 $Y=2.125
c135 52 0 1.44963e-19 $X=2.525 $Y=0.615
c136 36 0 1.61246e-19 $X=1.82 $Y=0.74
r137 74 75 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=1.39 $Y=1.465
+ $X2=1.445 $Y2=1.465
r138 73 74 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=0.995 $Y=1.465
+ $X2=1.39 $Y2=1.465
r139 72 73 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=0.96 $Y=1.465
+ $X2=0.995 $Y2=1.465
r140 68 70 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.53 $Y=1.465
+ $X2=0.545 $Y2=1.465
r141 62 64 15.5137 $w=2.58e-07 $l=3.5e-07 $layer=LI1_cond $X=4.09 $Y=1.11
+ $X2=4.09 $Y2=0.76
r142 61 67 8.61065 $w=1.7e-07 $l=1.68953e-07 $layer=LI1_cond $X=3.255 $Y=1.195
+ $X2=3.09 $Y2=1.187
r143 60 62 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.96 $Y=1.195
+ $X2=4.09 $Y2=1.11
r144 60 61 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=3.96 $Y=1.195
+ $X2=3.255 $Y2=1.195
r145 56 67 0.89609 $w=3.3e-07 $l=9.3e-08 $layer=LI1_cond $X=3.09 $Y=1.28
+ $X2=3.09 $Y2=1.187
r146 56 58 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=3.09 $Y=1.28
+ $X2=3.09 $Y2=2.125
r147 54 67 8.61065 $w=1.7e-07 $l=1.68464e-07 $layer=LI1_cond $X=2.925 $Y=1.18
+ $X2=3.09 $Y2=1.187
r148 54 55 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.925 $Y=1.18
+ $X2=2.61 $Y2=1.18
r149 50 55 7.50571 $w=3.35e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.485 $Y=1.095
+ $X2=2.61 $Y2=1.18
r150 50 52 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=2.485 $Y=1.095
+ $X2=2.485 $Y2=0.615
r151 49 77 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.82 $Y=1.465
+ $X2=1.895 $Y2=1.465
r152 49 75 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=1.82 $Y=1.465
+ $X2=1.445 $Y2=1.465
r153 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.82
+ $Y=1.465 $X2=1.82 $Y2=1.465
r154 45 72 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=0.8 $Y=1.465
+ $X2=0.96 $Y2=1.465
r155 45 70 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=0.8 $Y=1.465
+ $X2=0.545 $Y2=1.465
r156 44 48 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=0.8 $Y=1.465
+ $X2=1.82 $Y2=1.465
r157 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.8
+ $Y=1.465 $X2=0.8 $Y2=1.465
r158 42 50 22.397 $w=3.35e-07 $l=7.78315e-07 $layer=LI1_cond $X=1.87 $Y=1.465
+ $X2=2.485 $Y2=1.095
r159 42 48 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=1.87 $Y=1.465
+ $X2=1.82 $Y2=1.465
r160 38 77 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=1.63
+ $X2=1.895 $Y2=1.465
r161 38 40 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.895 $Y=1.63
+ $X2=1.895 $Y2=2.4
r162 34 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.82 $Y=1.3
+ $X2=1.82 $Y2=1.465
r163 34 36 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.82 $Y=1.3
+ $X2=1.82 $Y2=0.74
r164 30 75 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.445 $Y=1.63
+ $X2=1.445 $Y2=1.465
r165 30 32 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.445 $Y=1.63
+ $X2=1.445 $Y2=2.4
r166 26 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.39 $Y=1.3
+ $X2=1.39 $Y2=1.465
r167 26 28 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.39 $Y=1.3
+ $X2=1.39 $Y2=0.74
r168 22 73 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.63
+ $X2=0.995 $Y2=1.465
r169 22 24 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.995 $Y=1.63
+ $X2=0.995 $Y2=2.4
r170 18 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.3
+ $X2=0.96 $Y2=1.465
r171 18 20 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.96 $Y=1.3
+ $X2=0.96 $Y2=0.74
r172 14 70 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.63
+ $X2=0.545 $Y2=1.465
r173 14 16 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.545 $Y=1.63
+ $X2=0.545 $Y2=2.4
r174 10 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.3
+ $X2=0.53 $Y2=1.465
r175 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.53 $Y=1.3
+ $X2=0.53 $Y2=0.74
r176 3 58 300 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=2 $X=2.955
+ $Y=1.96 $X2=3.09 $Y2=2.125
r177 2 64 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=3.915
+ $Y=0.37 $X2=4.055 $Y2=0.76
r178 1 52 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.385
+ $Y=0.47 $X2=2.525 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__A21O_4%B1 3 7 11 15 17 26
c51 17 0 1.33616e-19 $X=2.64 $Y=1.665
c52 15 0 2.71749e-19 $X=3.315 $Y=2.46
c53 7 0 1.44963e-19 $X=2.74 $Y=0.79
r54 25 26 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=2.865 $Y=1.6
+ $X2=3.315 $Y2=1.6
r55 24 25 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=2.74 $Y=1.6
+ $X2=2.865 $Y2=1.6
r56 22 24 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.59 $Y=1.6 $X2=2.74
+ $Y2=1.6
r57 19 22 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=2.31 $Y=1.6 $X2=2.59
+ $Y2=1.6
r58 17 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.59
+ $Y=1.6 $X2=2.59 $Y2=1.6
r59 13 26 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.315 $Y=1.765
+ $X2=3.315 $Y2=1.6
r60 13 15 270.153 $w=1.8e-07 $l=6.95e-07 $layer=POLY_cond $X=3.315 $Y=1.765
+ $X2=3.315 $Y2=2.46
r61 9 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.765
+ $X2=2.865 $Y2=1.6
r62 9 11 270.153 $w=1.8e-07 $l=6.95e-07 $layer=POLY_cond $X=2.865 $Y=1.765
+ $X2=2.865 $Y2=2.46
r63 5 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=1.435
+ $X2=2.74 $Y2=1.6
r64 5 7 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.74 $Y=1.435
+ $X2=2.74 $Y2=0.79
r65 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.31 $Y=1.435
+ $X2=2.31 $Y2=1.6
r66 1 3 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.31 $Y=1.435
+ $X2=2.31 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_MS__A21O_4%A1 3 7 11 15 17 18 25
c57 15 0 1.9142e-19 $X=4.27 $Y=0.69
c58 3 0 5.66563e-20 $X=3.765 $Y=2.46
r59 25 26 8.31034 $w=3.19e-07 $l=5.5e-08 $layer=POLY_cond $X=4.215 $Y=1.615
+ $X2=4.27 $Y2=1.615
r60 23 25 56.6614 $w=3.19e-07 $l=3.75e-07 $layer=POLY_cond $X=3.84 $Y=1.615
+ $X2=4.215 $Y2=1.615
r61 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.84
+ $Y=1.615 $X2=3.84 $Y2=1.615
r62 21 23 11.3323 $w=3.19e-07 $l=7.5e-08 $layer=POLY_cond $X=3.765 $Y=1.615
+ $X2=3.84 $Y2=1.615
r63 18 24 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=4.08 $Y=1.615
+ $X2=3.84 $Y2=1.615
r64 17 24 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.6 $Y=1.615 $X2=3.84
+ $Y2=1.615
r65 13 26 20.418 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.27 $Y=1.45
+ $X2=4.27 $Y2=1.615
r66 13 15 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=4.27 $Y=1.45
+ $X2=4.27 $Y2=0.69
r67 9 25 16.143 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.215 $Y=1.78
+ $X2=4.215 $Y2=1.615
r68 9 11 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=4.215 $Y=1.78
+ $X2=4.215 $Y2=2.46
r69 5 23 20.418 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.84 $Y=1.45 $X2=3.84
+ $Y2=1.615
r70 5 7 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=3.84 $Y=1.45 $X2=3.84
+ $Y2=0.69
r71 1 21 16.143 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.765 $Y=1.78
+ $X2=3.765 $Y2=1.615
r72 1 3 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=3.765 $Y=1.78
+ $X2=3.765 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A21O_4%A2 3 7 11 15 17 24 26
c44 26 0 1.66816e-20 $X=5.13 $Y=1.425
c45 7 0 1.83628e-19 $X=4.7 $Y=0.69
c46 3 0 1.53462e-19 $X=4.665 $Y=2.46
r47 25 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.115 $Y=1.425
+ $X2=5.13 $Y2=1.425
r48 23 25 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=4.74 $Y=1.425
+ $X2=5.115 $Y2=1.425
r49 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.74
+ $Y=1.425 $X2=4.74 $Y2=1.425
r50 21 23 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=4.7 $Y=1.425 $X2=4.74
+ $Y2=1.425
r51 19 21 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=4.665 $Y=1.425
+ $X2=4.7 $Y2=1.425
r52 17 24 6.24041 $w=4.58e-07 $l=2.4e-07 $layer=LI1_cond $X=4.675 $Y=1.665
+ $X2=4.675 $Y2=1.425
r53 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.13 $Y=1.26
+ $X2=5.13 $Y2=1.425
r54 13 15 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=5.13 $Y=1.26
+ $X2=5.13 $Y2=0.69
r55 9 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.115 $Y=1.59
+ $X2=5.115 $Y2=1.425
r56 9 11 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=5.115 $Y=1.59
+ $X2=5.115 $Y2=2.46
r57 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.7 $Y=1.26 $X2=4.7
+ $Y2=1.425
r58 5 7 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=4.7 $Y=1.26 $X2=4.7
+ $Y2=0.69
r59 1 19 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.665 $Y=1.59
+ $X2=4.665 $Y2=1.425
r60 1 3 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=4.665 $Y=1.59
+ $X2=4.665 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A21O_4%VPWR 1 2 3 4 5 16 18 22 26 32 36 39 40 42 43
+ 44 46 51 67 68 74 77
c83 32 0 1.87992e-19 $X=3.99 $Y=2.455
r84 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r85 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r86 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r87 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r88 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r89 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r90 62 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r91 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r92 59 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r93 58 61 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r94 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r95 56 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.285 $Y=3.33
+ $X2=2.16 $Y2=3.33
r96 56 58 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.285 $Y=3.33
+ $X2=2.64 $Y2=3.33
r97 55 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r98 55 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r99 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r100 52 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.305 $Y=3.33
+ $X2=1.18 $Y2=3.33
r101 52 54 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.305 $Y=3.33
+ $X2=1.68 $Y2=3.33
r102 51 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=2.16 $Y2=3.33
r103 51 54 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=1.68 $Y2=3.33
r104 50 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r105 50 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r106 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r107 47 71 4.64823 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=0.485 $Y=3.33
+ $X2=0.242 $Y2=3.33
r108 47 49 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.485 $Y=3.33
+ $X2=0.72 $Y2=3.33
r109 46 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.18 $Y2=3.33
r110 46 49 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.72 $Y2=3.33
r111 44 62 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.6 $Y2=3.33
r112 44 59 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r113 42 64 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.725 $Y=3.33
+ $X2=4.56 $Y2=3.33
r114 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.725 $Y=3.33
+ $X2=4.89 $Y2=3.33
r115 41 67 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=5.055 $Y=3.33
+ $X2=5.52 $Y2=3.33
r116 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.055 $Y=3.33
+ $X2=4.89 $Y2=3.33
r117 39 61 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.825 $Y=3.33
+ $X2=3.6 $Y2=3.33
r118 39 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.825 $Y=3.33
+ $X2=3.95 $Y2=3.33
r119 38 64 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=4.075 $Y=3.33
+ $X2=4.56 $Y2=3.33
r120 38 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.075 $Y=3.33
+ $X2=3.95 $Y2=3.33
r121 34 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.89 $Y=3.245
+ $X2=4.89 $Y2=3.33
r122 34 36 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=4.89 $Y=3.245
+ $X2=4.89 $Y2=2.455
r123 30 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.95 $Y=3.245
+ $X2=3.95 $Y2=3.33
r124 30 32 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=3.95 $Y=3.245
+ $X2=3.95 $Y2=2.455
r125 26 29 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=2.16 $Y=2.115
+ $X2=2.16 $Y2=2.815
r126 24 77 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=3.245
+ $X2=2.16 $Y2=3.33
r127 24 29 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.16 $Y=3.245
+ $X2=2.16 $Y2=2.815
r128 20 74 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r129 20 22 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.305
r130 16 71 3.11795 $w=3.3e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.32 $Y=3.245
+ $X2=0.242 $Y2=3.33
r131 16 18 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=0.32 $Y=3.245
+ $X2=0.32 $Y2=2.225
r132 5 36 300 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=2 $X=4.755
+ $Y=1.96 $X2=4.89 $Y2=2.455
r133 4 32 300 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=2 $X=3.855
+ $Y=1.96 $X2=3.99 $Y2=2.455
r134 3 29 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.985
+ $Y=1.84 $X2=2.12 $Y2=2.815
r135 3 26 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.985
+ $Y=1.84 $X2=2.12 $Y2=2.115
r136 2 22 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=1.84 $X2=1.22 $Y2=2.305
r137 1 18 300 $w=1.7e-07 $l=4.43114e-07 $layer=licon1_PDIFF $count=2 $X=0.195
+ $Y=1.84 $X2=0.32 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_MS__A21O_4%X 1 2 3 4 13 14 15 16 19 23 27 29 33 37 43 44
+ 45 46
c72 27 0 1.61246e-19 $X=1.44 $Y=1.045
r73 45 46 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r74 42 46 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.24 $Y=1.8
+ $X2=0.24 $Y2=1.665
r75 41 45 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.13
+ $X2=0.24 $Y2=1.295
r76 37 39 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.67 $Y=1.985
+ $X2=1.67 $Y2=2.815
r77 35 37 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.67 $Y=1.97
+ $X2=1.67 $Y2=1.985
r78 31 33 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=1.565 $Y=0.96
+ $X2=1.565 $Y2=0.515
r79 30 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.855 $Y=1.885
+ $X2=0.77 $Y2=1.885
r80 29 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.505 $Y=1.885
+ $X2=1.67 $Y2=1.97
r81 29 30 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.505 $Y=1.885
+ $X2=0.855 $Y2=1.885
r82 28 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.83 $Y=1.045
+ $X2=0.745 $Y2=1.045
r83 27 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.44 $Y=1.045
+ $X2=1.565 $Y2=0.96
r84 27 28 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.44 $Y=1.045
+ $X2=0.83 $Y2=1.045
r85 23 25 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=0.77 $Y=1.985
+ $X2=0.77 $Y2=2.815
r86 21 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=1.97 $X2=0.77
+ $Y2=1.885
r87 21 23 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.77 $Y=1.97
+ $X2=0.77 $Y2=1.985
r88 17 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=0.96
+ $X2=0.745 $Y2=1.045
r89 17 19 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=0.745 $Y=0.96
+ $X2=0.745 $Y2=0.515
r90 16 42 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.885
+ $X2=0.24 $Y2=1.8
r91 15 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=1.885
+ $X2=0.77 $Y2=1.885
r92 15 16 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.685 $Y=1.885
+ $X2=0.355 $Y2=1.885
r93 14 41 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.045
+ $X2=0.24 $Y2=1.13
r94 13 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.66 $Y=1.045
+ $X2=0.745 $Y2=1.045
r95 13 14 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.66 $Y=1.045
+ $X2=0.355 $Y2=1.045
r96 4 39 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.535
+ $Y=1.84 $X2=1.67 $Y2=2.815
r97 4 37 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.535
+ $Y=1.84 $X2=1.67 $Y2=1.985
r98 3 25 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.635
+ $Y=1.84 $X2=0.77 $Y2=2.815
r99 3 23 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.635
+ $Y=1.84 $X2=0.77 $Y2=1.985
r100 2 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.465
+ $Y=0.37 $X2=1.605 $Y2=0.515
r101 1 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.605
+ $Y=0.37 $X2=0.745 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A21O_4%A_503_392# 1 2 3 4 15 19 20 21 25 29 31 33 35
+ 40
c56 29 0 1.53462e-19 $X=4.44 $Y=2.815
c57 21 0 8.37567e-20 $X=3.54 $Y=2.12
r58 33 42 2.9222 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=5.38 $Y=2.12 $X2=5.38
+ $Y2=2.03
r59 33 35 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=5.38 $Y=2.12
+ $X2=5.38 $Y2=2.815
r60 32 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.525 $Y=2.035
+ $X2=4.4 $Y2=2.035
r61 31 42 4.22096 $w=1.7e-07 $l=1.27475e-07 $layer=LI1_cond $X=5.255 $Y=2.035
+ $X2=5.38 $Y2=2.03
r62 31 32 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.255 $Y=2.035
+ $X2=4.525 $Y2=2.035
r63 27 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.4 $Y=2.12
+ $X2=4.4 $Y2=2.035
r64 27 29 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=4.4 $Y=2.12 $X2=4.4
+ $Y2=2.815
r65 26 38 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=2.035
+ $X2=3.54 $Y2=2.035
r66 25 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.275 $Y=2.035
+ $X2=4.4 $Y2=2.035
r67 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.275 $Y=2.035
+ $X2=3.625 $Y2=2.035
r68 22 24 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.54 $Y=2.905 $X2=3.54
+ $Y2=2.815
r69 21 38 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=2.12 $X2=3.54
+ $Y2=2.035
r70 21 24 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.54 $Y=2.12
+ $X2=3.54 $Y2=2.815
r71 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.455 $Y=2.99
+ $X2=3.54 $Y2=2.905
r72 19 20 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.455 $Y=2.99
+ $X2=2.725 $Y2=2.99
r73 15 18 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=2.6 $Y=2.115 $X2=2.6
+ $Y2=2.815
r74 13 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.6 $Y=2.905
+ $X2=2.725 $Y2=2.99
r75 13 18 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=2.6 $Y=2.905 $X2=2.6
+ $Y2=2.815
r76 4 42 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.205
+ $Y=1.96 $X2=5.34 $Y2=2.105
r77 4 35 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.205
+ $Y=1.96 $X2=5.34 $Y2=2.815
r78 3 40 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=4.305
+ $Y=1.96 $X2=4.44 $Y2=2.115
r79 3 29 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.305
+ $Y=1.96 $X2=4.44 $Y2=2.815
r80 2 38 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.96 $X2=3.54 $Y2=2.115
r81 2 24 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.96 $X2=3.54 $Y2=2.815
r82 1 18 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.515
+ $Y=1.96 $X2=2.64 $Y2=2.815
r83 1 15 400 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=2.515
+ $Y=1.96 $X2=2.64 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__A21O_4%VGND 1 2 3 4 5 16 18 22 26 30 34 37 38 40 41
+ 43 44 46 47 48 67 68
c87 34 0 1.9142e-19 $X=4.915 $Y=0.585
r88 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r89 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r90 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r91 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r92 62 65 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.56
+ $Y2=0
r93 61 64 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.56
+ $Y2=0
r94 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r95 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r96 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r97 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r98 53 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r99 53 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r100 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r101 50 71 4.65971 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=0.48 $Y=0 $X2=0.24
+ $Y2=0
r102 50 52 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.48 $Y=0 $X2=0.72
+ $Y2=0
r103 48 62 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=3.12 $Y2=0
r104 48 59 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=2.64 $Y2=0
r105 46 64 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.75 $Y=0 $X2=4.56
+ $Y2=0
r106 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.75 $Y=0 $X2=4.915
+ $Y2=0
r107 45 67 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=5.52
+ $Y2=0
r108 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.08 $Y=0 $X2=4.915
+ $Y2=0
r109 44 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.955 $Y=0 $X2=3.12
+ $Y2=0
r110 43 58 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.79 $Y=0 $X2=2.64
+ $Y2=0
r111 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.79 $Y=0 $X2=2.955
+ $Y2=0
r112 40 55 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.87 $Y=0 $X2=1.68
+ $Y2=0
r113 40 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.87 $Y=0 $X2=1.995
+ $Y2=0
r114 39 58 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.12 $Y=0 $X2=2.64
+ $Y2=0
r115 39 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.12 $Y=0 $X2=1.995
+ $Y2=0
r116 37 52 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=0.72
+ $Y2=0
r117 37 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.01 $Y=0 $X2=1.135
+ $Y2=0
r118 36 55 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.68
+ $Y2=0
r119 36 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.135
+ $Y2=0
r120 32 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.915 $Y=0.085
+ $X2=4.915 $Y2=0
r121 32 34 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=4.915 $Y=0.085
+ $X2=4.915 $Y2=0.585
r122 28 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.955 $Y=0.085
+ $X2=2.955 $Y2=0
r123 28 30 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.955 $Y=0.085
+ $X2=2.955 $Y2=0.76
r124 24 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.995 $Y=0.085
+ $X2=1.995 $Y2=0
r125 24 26 28.5806 $w=2.48e-07 $l=6.2e-07 $layer=LI1_cond $X=1.995 $Y=0.085
+ $X2=1.995 $Y2=0.705
r126 20 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0.085
+ $X2=1.135 $Y2=0
r127 20 22 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=1.135 $Y=0.085
+ $X2=1.135 $Y2=0.625
r128 16 71 3.10647 $w=3.3e-07 $l=1.16619e-07 $layer=LI1_cond $X=0.315 $Y=0.085
+ $X2=0.24 $Y2=0
r129 16 18 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=0.315 $Y=0.085
+ $X2=0.315 $Y2=0.625
r130 5 34 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=4.775
+ $Y=0.37 $X2=4.915 $Y2=0.585
r131 4 30 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=2.815
+ $Y=0.47 $X2=2.955 $Y2=0.76
r132 3 26 182 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.37 $X2=2.035 $Y2=0.705
r133 2 22 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.37 $X2=1.175 $Y2=0.625
r134 1 18 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=0.17
+ $Y=0.37 $X2=0.315 $Y2=0.625
.ends

.subckt PM_SKY130_FD_SC_MS__A21O_4%A_700_74# 1 2 3 12 14 15 20 21 24
r37 22 24 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=5.385 $Y=0.92
+ $X2=5.385 $Y2=0.515
r38 20 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.26 $Y=1.005
+ $X2=5.385 $Y2=0.92
r39 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.26 $Y=1.005
+ $X2=4.57 $Y2=1.005
r40 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.485 $Y=0.92
+ $X2=4.57 $Y2=1.005
r41 17 19 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.485 $Y=0.92
+ $X2=4.485 $Y2=0.515
r42 16 19 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.485 $Y=0.425
+ $X2=4.485 $Y2=0.515
r43 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.4 $Y=0.34
+ $X2=4.485 $Y2=0.425
r44 14 15 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.4 $Y=0.34 $X2=3.79
+ $Y2=0.34
r45 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.625 $Y=0.425
+ $X2=3.79 $Y2=0.34
r46 10 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.625 $Y=0.425
+ $X2=3.625 $Y2=0.515
r47 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.205
+ $Y=0.37 $X2=5.345 $Y2=0.515
r48 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.345
+ $Y=0.37 $X2=4.485 $Y2=0.515
r49 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=3.5
+ $Y=0.37 $X2=3.625 $Y2=0.515
.ends


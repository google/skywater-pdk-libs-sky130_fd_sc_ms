* File: sky130_fd_sc_ms__dlrbn_2.spice
* Created: Fri Aug 28 17:26:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dlrbn_2.pex.spice"
.subckt sky130_fd_sc_ms__dlrbn_2  VNB VPB D GATE_N RESET_B VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1016 N_VGND_M1016_d N_D_M1016_g N_A_27_112#_M1016_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.129591 AS=0.15675 PD=0.997674 PS=1.67 NRD=17.988 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1013 N_A_230_74#_M1013_d N_GATE_N_M1013_g N_VGND_M1016_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1022_d N_A_230_74#_M1022_g N_A_363_74#_M1022_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.205591 AS=0.2109 PD=1.3942 PS=2.05 NRD=28.368 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1006 A_592_74# N_A_27_112#_M1006_g N_VGND_M1022_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.177809 PD=0.88 PS=1.2058 NRD=12.18 NRS=19.68 M=1 R=4.26667
+ SA=75000.9 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1007 N_A_670_74#_M1007_d N_A_230_74#_M1007_g A_592_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.147321 AS=0.0768 PD=1.31623 PS=0.88 NRD=15.936 NRS=12.18 M=1
+ R=4.26667 SA=75001.3 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1017 A_790_74# N_A_363_74#_M1017_g N_A_670_74#_M1007_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0966792 PD=0.66 PS=0.863774 NRD=18.564 NRS=24.276 M=1
+ R=2.8 SA=75001.9 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_A_838_48#_M1023_g A_790_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 A_1066_74# N_A_670_74#_M1001_g N_A_838_48#_M1001_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_RESET_B_M1002_g A_1066_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1628 AS=0.0888 PD=1.18 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75000.6
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1003 N_Q_M1003_d N_A_838_48#_M1003_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1628 PD=1.02 PS=1.18 NRD=0 NRS=25.944 M=1 R=4.93333 SA=75001.2
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1019 N_Q_M1003_d N_A_838_48#_M1019_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.133522 PD=1.02 PS=1.16899 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1018 N_A_1448_74#_M1018_d N_A_838_48#_M1018_g N_VGND_M1019_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.115478 PD=1.85 PS=1.01101 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75002.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1020 N_VGND_M1020_d N_A_1448_74#_M1020_g N_Q_N_M1020_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1184 PD=2.05 PS=1.06 NRD=0 NRS=3.24 M=1 R=4.93333
+ SA=75000.2 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1027 N_VGND_M1027_d N_A_1448_74#_M1027_g N_Q_N_M1020_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1184 PD=2.05 PS=1.06 NRD=0 NRS=3.24 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1012 N_VPWR_M1012_d N_D_M1012_g N_A_27_112#_M1012_s VPB PSHORT L=0.18 W=0.84
+ AD=0.21 AS=0.2352 PD=1.34 PS=2.24 NRD=0 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.9 A=0.1512 P=2.04 MULT=1
MM1015 N_A_230_74#_M1015_d N_GATE_N_M1015_g N_VPWR_M1012_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.21 PD=2.24 PS=1.34 NRD=0 NRS=52.7566 M=1 R=4.66667
+ SA=90000.9 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1005 N_VPWR_M1005_d N_A_230_74#_M1005_g N_A_363_74#_M1005_s VPB PSHORT L=0.18
+ W=0.84 AD=0.217898 AS=0.3704 PD=1.47 PS=2.85 NRD=47.9301 NRS=19.9167 M=1
+ R=4.66667 SA=90000.3 SB=90002.4 A=0.1512 P=2.04 MULT=1
MM1009 A_598_392# N_A_27_112#_M1009_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=1
+ AD=0.105 AS=0.259402 PD=1.21 PS=1.75 NRD=9.8303 NRS=16.7253 M=1 R=5.55556
+ SA=90000.8 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1024 N_A_670_74#_M1024_d N_A_363_74#_M1024_g A_598_392# VPB PSHORT L=0.18 W=1
+ AD=0.22993 AS=0.105 PD=1.92958 PS=1.21 NRD=0 NRS=9.8303 M=1 R=5.55556
+ SA=90001.2 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1014 A_786_508# N_A_230_74#_M1014_g N_A_670_74#_M1024_d VPB PSHORT L=0.18
+ W=0.42 AD=0.09345 AS=0.0965704 PD=0.865 PS=0.810423 NRD=78.5636 NRS=44.5417
+ M=1 R=2.33333 SA=90001.6 SB=90003.4 A=0.0756 P=1.2 MULT=1
MM1004 N_VPWR_M1004_d N_A_838_48#_M1004_g A_786_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.115882 AS=0.09345 PD=0.935455 PS=0.865 NRD=63.3158 NRS=78.5636 M=1
+ R=2.33333 SA=90002.2 SB=90002.7 A=0.0756 P=1.2 MULT=1
MM1011 N_A_838_48#_M1011_d N_A_670_74#_M1011_g N_VPWR_M1004_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1568 AS=0.309018 PD=1.4 PS=2.49455 NRD=0.8668 NRS=31.6579 M=1
+ R=6.22222 SA=90001.2 SB=90002 A=0.2016 P=2.6 MULT=1
MM1026 N_VPWR_M1026_d N_RESET_B_M1026_g N_A_838_48#_M1011_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1792 AS=0.1568 PD=1.44 PS=1.4 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90001.7 SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1000 N_VPWR_M1026_d N_A_838_48#_M1000_g N_Q_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.2
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1025 N_VPWR_M1025_d N_A_838_48#_M1025_g N_Q_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.187547 AS=0.1512 PD=1.52679 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.6
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1021 N_A_1448_74#_M1021_d N_A_838_48#_M1021_g N_VPWR_M1025_d VPB PSHORT L=0.18
+ W=1 AD=0.28 AS=0.167453 PD=2.56 PS=1.36321 NRD=0 NRS=9.8303 M=1 R=5.55556
+ SA=90003 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1008 N_Q_N_M1008_d N_A_1448_74#_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1010 N_Q_N_M1008_d N_A_1448_74#_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX28_noxref VNB VPB NWDIODE A=17.754 P=22.92
c_96 VNB 0 1.25688e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__dlrbn_2.pxi.spice"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sedfxbp_2 CLK D DE SCD SCE VGND VNB VPB VPWR Q Q_N
X0 VPWR a_575_87# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 a_2591_74# a_575_87# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X2 VGND a_183_290# a_527_113# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 a_141_74# DE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X4 a_1091_125# SCE a_691_113# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X5 a_691_113# a_1377_368# a_1784_97# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X6 VPWR a_2489_74# a_575_87# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 VGND a_2489_74# a_575_87# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_32_74# SCE a_691_113# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X9 a_661_87# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X10 VGND a_2013_71# a_2417_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X11 a_691_113# a_1586_74# a_1784_97# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X12 a_2377_392# a_1377_368# a_2489_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X13 VPWR DE a_581_462# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X14 a_1947_508# a_2013_71# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X15 VPWR SCD a_1091_453# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X16 a_2489_74# a_1377_368# a_2591_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X17 Q a_2489_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X18 VGND a_2489_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 VGND a_1377_368# a_1586_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 Q_N a_575_87# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X21 a_1091_453# a_661_87# a_691_113# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X22 a_2675_508# a_575_87# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X23 a_661_87# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X24 VPWR CLK a_1377_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X25 a_1784_97# a_1586_74# a_1920_97# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X26 a_2417_74# a_1586_74# a_2489_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X27 a_135_464# a_183_290# VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X28 VGND a_575_87# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X29 a_581_462# a_575_87# a_32_74# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X30 a_527_113# a_575_87# a_32_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X31 VPWR a_1377_368# a_1586_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X32 VGND CLK a_1377_368# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X33 Q a_2489_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X34 a_183_290# DE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X35 VPWR a_1784_97# a_2013_71# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X36 a_32_74# D a_141_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X37 a_1784_97# a_1377_368# a_1947_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X38 VGND SCD a_1091_125# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X39 VPWR a_2013_71# a_2377_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X40 a_32_74# D a_135_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X41 a_183_290# DE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X42 VGND a_1784_97# a_2013_71# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X43 Q_N a_575_87# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X44 a_2489_74# a_1586_74# a_2675_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X45 a_1920_97# a_2013_71# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X46 a_32_74# a_661_87# a_691_113# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X47 VPWR a_2489_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
.ends

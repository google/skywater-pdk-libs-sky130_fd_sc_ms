# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__sdfstp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__sdfstp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.92000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.820000 1.580000 2.150000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.513300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.380000 0.350000 13.815000 1.050000 ;
        RECT 13.565000 1.050000 13.815000 2.980000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 1.140000 2.805000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.280000 0.680000 1.440000 ;
        RECT 0.425000 1.440000 2.045000 1.610000 ;
        RECT 0.425000 1.610000 0.835000 1.950000 ;
        RECT 1.790000 1.260000 2.045000 1.440000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.277200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  7.145000 1.540000  7.555000 1.800000 ;
        RECT 10.685000 1.380000 11.030000 2.050000 ;
      LAYER mcon ;
        RECT  7.355000 1.580000  7.525000 1.750000 ;
        RECT 10.715000 1.580000 10.885000 1.750000 ;
      LAYER met1 ;
        RECT  7.295000 1.550000  7.585000 1.595000 ;
        RECT  7.295000 1.595000 10.945000 1.735000 ;
        RECT  7.295000 1.735000  7.585000 1.780000 ;
        RECT 10.655000 1.550000 10.945000 1.595000 ;
        RECT 10.655000 1.735000 10.945000 1.780000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.315000 1.180000 3.715000 1.550000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 13.920000 0.085000 ;
        RECT  0.695000  0.085000  1.025000 0.770000 ;
        RECT  2.375000  0.085000  2.705000 0.750000 ;
        RECT  3.475000  0.085000  3.805000 1.010000 ;
        RECT  6.115000  0.085000  6.445000 0.690000 ;
        RECT  7.455000  0.085000  8.305000 0.940000 ;
        RECT 10.825000  0.085000 11.155000 0.810000 ;
        RECT 12.880000  0.085000 13.210000 1.050000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.920000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 13.920000 3.415000 ;
        RECT  0.560000 2.660000  0.890000 3.245000 ;
        RECT  2.565000 2.830000  2.895000 3.245000 ;
        RECT  3.575000 2.580000  3.905000 3.245000 ;
        RECT  6.225000 2.685000  6.475000 3.245000 ;
        RECT  7.665000 2.310000  7.915000 3.245000 ;
        RECT 10.630000 2.560000 10.800000 3.245000 ;
        RECT 12.070000 2.560000 12.320000 3.245000 ;
        RECT 13.030000 1.995000 13.360000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 13.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.085000 0.350000  0.525000 0.940000 ;
      RECT  0.085000 0.940000  1.220000 1.110000 ;
      RECT  0.085000 1.110000  0.255000 2.300000 ;
      RECT  0.085000 2.300000  0.360000 2.320000 ;
      RECT  0.085000 2.320000  2.045000 2.490000 ;
      RECT  0.085000 2.490000  0.360000 2.980000 ;
      RECT  0.890000 1.110000  1.220000 1.270000 ;
      RECT  1.430000 2.660000  2.385000 2.910000 ;
      RECT  1.555000 0.350000  1.885000 0.920000 ;
      RECT  1.555000 0.920000  2.385000 1.090000 ;
      RECT  1.790000 1.830000  2.045000 2.320000 ;
      RECT  2.215000 1.090000  2.385000 2.490000 ;
      RECT  2.215000 2.490000  3.405000 2.660000 ;
      RECT  2.975000 0.350000  3.305000 1.010000 ;
      RECT  2.975000 1.010000  3.145000 1.820000 ;
      RECT  2.975000 1.820000  4.215000 2.070000 ;
      RECT  3.235000 2.240000  5.005000 2.410000 ;
      RECT  3.235000 2.410000  3.405000 2.490000 ;
      RECT  3.885000 1.350000  4.215000 1.820000 ;
      RECT  3.975000 0.255000  5.205000 0.425000 ;
      RECT  3.975000 0.425000  4.225000 1.130000 ;
      RECT  4.105000 2.580000  4.275000 2.895000 ;
      RECT  4.105000 2.895000  5.845000 3.065000 ;
      RECT  4.445000 0.595000  4.865000 0.765000 ;
      RECT  4.445000 0.765000  4.615000 2.240000 ;
      RECT  4.445000 2.410000  5.005000 2.725000 ;
      RECT  4.785000 0.935000  5.205000 1.105000 ;
      RECT  4.785000 1.105000  5.005000 2.070000 ;
      RECT  5.035000 0.425000  5.205000 0.935000 ;
      RECT  5.175000 1.275000  6.070000 1.435000 ;
      RECT  5.175000 1.435000  6.935000 1.445000 ;
      RECT  5.175000 1.445000  5.345000 2.265000 ;
      RECT  5.175000 2.265000  5.505000 2.725000 ;
      RECT  5.375000 0.385000  5.625000 1.275000 ;
      RECT  5.515000 1.615000  5.730000 1.775000 ;
      RECT  5.515000 1.775000  5.845000 1.945000 ;
      RECT  5.675000 1.945000  5.845000 2.345000 ;
      RECT  5.675000 2.345000  6.815000 2.515000 ;
      RECT  5.675000 2.515000  5.845000 2.895000 ;
      RECT  5.900000 1.445000  6.935000 1.605000 ;
      RECT  6.015000 1.795000  6.345000 2.005000 ;
      RECT  6.015000 2.005000  7.155000 2.175000 ;
      RECT  6.240000 0.860000  7.005000 1.030000 ;
      RECT  6.240000 1.030000  6.480000 1.265000 ;
      RECT  6.645000 2.515000  6.815000 2.895000 ;
      RECT  6.645000 2.895000  7.495000 3.065000 ;
      RECT  6.650000 1.200000  8.430000 1.370000 ;
      RECT  6.650000 1.370000  6.935000 1.435000 ;
      RECT  6.650000 1.605000  6.935000 1.835000 ;
      RECT  6.675000 0.570000  7.005000 0.860000 ;
      RECT  6.985000 2.175000  7.155000 2.725000 ;
      RECT  7.325000 1.970000  7.945000 2.140000 ;
      RECT  7.325000 2.140000  7.495000 2.895000 ;
      RECT  7.760000 1.120000  8.430000 1.200000 ;
      RECT  7.760000 1.370000  8.430000 1.410000 ;
      RECT  7.775000 1.580000  8.840000 1.750000 ;
      RECT  7.775000 1.750000  7.945000 1.970000 ;
      RECT  8.115000 1.920000  8.365000 2.350000 ;
      RECT  8.115000 2.350000  9.895000 2.520000 ;
      RECT  8.115000 2.520000  8.365000 2.725000 ;
      RECT  8.585000 2.690000  8.915000 2.905000 ;
      RECT  8.585000 2.905000 10.430000 3.075000 ;
      RECT  8.670000 1.120000  9.000000 1.450000 ;
      RECT  8.670000 1.450000  8.840000 1.580000 ;
      RECT  8.795000 0.350000  9.365000 0.940000 ;
      RECT  9.090000 1.620000 10.235000 1.790000 ;
      RECT  9.090000 1.790000  9.365000 2.180000 ;
      RECT  9.195000 0.940000  9.365000 1.620000 ;
      RECT  9.565000 1.960000  9.895000 2.350000 ;
      RECT  9.565000 2.520000  9.895000 2.735000 ;
      RECT  9.790000 0.980000 11.770000 1.040000 ;
      RECT  9.790000 1.040000 11.940000 1.210000 ;
      RECT  9.790000 1.210000 10.460000 1.310000 ;
      RECT 10.065000 1.790000 10.235000 2.220000 ;
      RECT 10.065000 2.220000 11.370000 2.390000 ;
      RECT 10.100000 2.560000 10.430000 2.905000 ;
      RECT 11.000000 2.390000 11.370000 2.980000 ;
      RECT 11.200000 1.380000 11.600000 2.050000 ;
      RECT 11.200000 2.050000 11.370000 2.220000 ;
      RECT 11.395000 0.350000 11.770000 0.980000 ;
      RECT 11.540000 2.220000 11.940000 2.390000 ;
      RECT 11.540000 2.390000 11.870000 2.980000 ;
      RECT 11.770000 1.210000 11.940000 2.220000 ;
      RECT 11.955000 0.540000 12.700000 0.870000 ;
      RECT 12.370000 0.870000 12.700000 1.005000 ;
      RECT 12.530000 1.005000 12.700000 1.220000 ;
      RECT 12.530000 1.220000 13.395000 1.550000 ;
      RECT 12.530000 1.550000 12.700000 1.995000 ;
      RECT 12.530000 1.995000 12.860000 2.875000 ;
  END
END sky130_fd_sc_ms__sdfstp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 VPWR B1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=9.184e+11p pd=8.36e+06u as=1.232e+12p ps=1.116e+07u
M1001 a_310_368# A2 a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=6.832e+11p pd=5.7e+06u as=9.744e+11p ps=8.46e+06u
M1002 a_28_368# A2 a_310_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_27_74# A1 VGND VNB nlowvt w=740000u l=150000u
+  ad=1.1174e+12p pd=1.042e+07u as=6.956e+11p ps=6.32e+06u
M1004 a_670_74# C1 Y VNB nlowvt w=740000u l=150000u
+  ad=5.18e+11p pd=4.36e+06u as=4.218e+11p ps=4.1e+06u
M1005 VPWR A1 a_28_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR C1 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_670_74# B1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A3 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y C1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y C1 a_670_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A2 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_74# A2 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_28_368# A1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_27_74# B1 a_670_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_74# A3 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_310_368# A3 Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A1 a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Y A3 a_310_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

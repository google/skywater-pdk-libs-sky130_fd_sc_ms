* File: sky130_fd_sc_ms__sdfxbp_1.pex.spice
* Created: Wed Sep  2 12:31:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SDFXBP_1%A_31_74# 1 2 9 13 15 17 20 22 23 25 34 35
c88 23 0 1.68868e-19 $X=0.915 $Y=2.04
r89 35 43 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.005 $Y=1.96
+ $X2=2.005 $Y2=2.125
r90 34 37 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.005 $Y=1.96 $X2=2.005
+ $Y2=2.04
r91 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.005
+ $Y=1.96 $X2=2.005 $Y2=1.96
r92 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.69 $X2=0.75 $Y2=1.69
r93 25 27 10.2392 $w=3.78e-07 $l=2.2e-07 $layer=LI1_cond $X=0.275 $Y=0.565
+ $X2=0.275 $Y2=0.785
r94 23 31 9.09243 $w=3.85e-07 $l=2.85832e-07 $layer=LI1_cond $X=0.915 $Y=2.04
+ $X2=0.75 $Y2=1.825
r95 22 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.84 $Y=2.04
+ $X2=2.005 $Y2=2.04
r96 22 23 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=1.84 $Y=2.04
+ $X2=0.915 $Y2=2.04
r97 18 31 14.0379 $w=3.85e-07 $l=4.43e-07 $layer=LI1_cond $X=0.307 $Y=1.825
+ $X2=0.75 $Y2=1.825
r98 18 28 4.3413 $w=3.85e-07 $l=1.37e-07 $layer=LI1_cond $X=0.307 $Y=1.825
+ $X2=0.17 $Y2=1.825
r99 18 20 15.7975 $w=4.43e-07 $l=6.1e-07 $layer=LI1_cond $X=0.307 $Y=1.855
+ $X2=0.307 $Y2=2.465
r100 17 28 5.54671 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=0.17 $Y=1.525 $X2=0.17
+ $Y2=1.825
r101 17 27 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=0.17 $Y=1.525
+ $X2=0.17 $Y2=0.785
r102 15 32 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.94 $Y=1.69
+ $X2=0.75 $Y2=1.69
r103 13 43 200.185 $w=1.8e-07 $l=5.15e-07 $layer=POLY_cond $X=1.96 $Y=2.64
+ $X2=1.96 $Y2=2.125
r104 7 15 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.015 $Y=1.525
+ $X2=0.94 $Y2=1.69
r105 7 9 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=1.015 $Y=1.525
+ $X2=1.015 $Y2=0.58
r106 2 20 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.22
+ $Y=2.32 $X2=0.365 $Y2=2.465
r107 1 25 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=0.155
+ $Y=0.37 $X2=0.3 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_1%SCE 2 3 4 7 9 11 12 14 16 17 19 20 26 29 33
+ 35 38
r79 32 35 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.885 $Y=1.065
+ $X2=2.095 $Y2=1.065
r80 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.885
+ $Y=1.065 $X2=1.885 $Y2=1.065
r81 26 33 5.16202 $w=4.73e-07 $l=2.05e-07 $layer=LI1_cond $X=1.68 $Y=1.047
+ $X2=1.885 $Y2=1.047
r82 26 38 4.02225 $w=4.73e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=1.047
+ $X2=1.565 $Y2=1.047
r83 24 29 9.23372 $w=2.61e-07 $l=5e-08 $layer=POLY_cond $X=0.565 $Y=1.12
+ $X2=0.515 $Y2=1.12
r84 23 38 34.9225 $w=3.28e-07 $l=1e-06 $layer=LI1_cond $X=0.565 $Y=1.12
+ $X2=1.565 $Y2=1.12
r85 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.565
+ $Y=1.12 $X2=0.565 $Y2=1.12
r86 17 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.095 $Y=0.9
+ $X2=2.095 $Y2=1.065
r87 17 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.095 $Y=0.9
+ $X2=2.095 $Y2=0.58
r88 14 16 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.09 $Y=2.245
+ $X2=1.09 $Y2=2.64
r89 13 20 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.68 $Y=2.17 $X2=0.59
+ $Y2=2.17
r90 12 14 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1 $Y=2.17
+ $X2=1.09 $Y2=2.245
r91 12 13 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1 $Y=2.17 $X2=0.68
+ $Y2=2.17
r92 9 20 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=0.59 $Y=2.245 $X2=0.59
+ $Y2=2.17
r93 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.59 $Y=2.245
+ $X2=0.59 $Y2=2.64
r94 5 29 15.717 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=0.955
+ $X2=0.515 $Y2=1.12
r95 5 7 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=0.515 $Y=0.955
+ $X2=0.515 $Y2=0.58
r96 3 20 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.5 $Y=2.17 $X2=0.59
+ $Y2=2.17
r97 3 4 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=0.5 $Y=2.17 $X2=0.345
+ $Y2=2.17
r98 2 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.27 $Y=2.095
+ $X2=0.345 $Y2=2.17
r99 1 29 45.2452 $w=2.61e-07 $l=3.16938e-07 $layer=POLY_cond $X=0.27 $Y=1.285
+ $X2=0.515 $Y2=1.12
r100 1 2 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.27 $Y=1.285 $X2=0.27
+ $Y2=2.095
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_1%D 3 7 9 12 13
c35 12 0 1.68868e-19 $X=1.465 $Y=1.62
r36 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.62
+ $X2=1.465 $Y2=1.785
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.62
+ $X2=1.465 $Y2=1.455
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.465
+ $Y=1.62 $X2=1.465 $Y2=1.62
r39 9 13 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=1.2 $Y=1.62
+ $X2=1.465 $Y2=1.62
r40 7 15 332.347 $w=1.8e-07 $l=8.55e-07 $layer=POLY_cond $X=1.51 $Y=2.64
+ $X2=1.51 $Y2=1.785
r41 3 14 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=1.405 $Y=0.58
+ $X2=1.405 $Y2=1.455
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_1%SCD 3 7 9 10 14
c41 14 0 6.03804e-20 $X=2.545 $Y=1.775
c42 3 0 8.79478e-20 $X=2.485 $Y=0.58
r43 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.545 $Y=1.775
+ $X2=2.545 $Y2=1.94
r44 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.545 $Y=1.775
+ $X2=2.545 $Y2=1.61
r45 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.545
+ $Y=1.775 $X2=2.545 $Y2=1.775
r46 10 15 8.68508 $w=3.43e-07 $l=2.6e-07 $layer=LI1_cond $X=2.552 $Y=2.035
+ $X2=2.552 $Y2=1.775
r47 9 15 3.67446 $w=3.43e-07 $l=1.1e-07 $layer=LI1_cond $X=2.552 $Y=1.665
+ $X2=2.552 $Y2=1.775
r48 7 17 272.097 $w=1.8e-07 $l=7e-07 $layer=POLY_cond $X=2.5 $Y=2.64 $X2=2.5
+ $Y2=1.94
r49 3 16 528.149 $w=1.5e-07 $l=1.03e-06 $layer=POLY_cond $X=2.485 $Y=0.58
+ $X2=2.485 $Y2=1.61
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_1%CLK 1 3 6 8 11
c41 8 0 8.79478e-20 $X=3.6 $Y=1.295
c42 6 0 6.77941e-20 $X=3.21 $Y=2.4
r43 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.4
+ $Y=1.385 $X2=3.4 $Y2=1.385
r44 11 13 33.6691 $w=2.72e-07 $l=1.9e-07 $layer=POLY_cond $X=3.21 $Y=1.385
+ $X2=3.4 $Y2=1.385
r45 8 14 6.22942 $w=3.68e-07 $l=2e-07 $layer=LI1_cond $X=3.6 $Y=1.365 $X2=3.4
+ $Y2=1.365
r46 4 11 12.4592 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=1.55
+ $X2=3.21 $Y2=1.385
r47 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.21 $Y=1.55 $X2=3.21
+ $Y2=2.4
r48 1 11 39.8713 $w=2.72e-07 $l=2.96226e-07 $layer=POLY_cond $X=2.985 $Y=1.22
+ $X2=3.21 $Y2=1.385
r49 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.985 $Y=1.22 $X2=2.985
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_1%A_828_74# 1 2 9 11 13 16 20 24 25 28 30 31
+ 33 34 37 40 41 43 46 47 48 55 56 61 62 64 65 67 68 69 72 73
c198 68 0 1.71252e-20 $X=7.615 $Y=1.255
c199 62 0 2.55557e-20 $X=5.075 $Y=2.155
c200 56 0 1.07508e-19 $X=8.515 $Y=1.52
c201 55 0 8.08518e-20 $X=8.515 $Y=1.52
c202 37 0 1.67448e-19 $X=5.892 $Y=0.69
c203 25 0 1.8865e-19 $X=8.395 $Y=2.17
c204 24 0 1.40714e-19 $X=8.395 $Y=2.02
r205 72 73 8.96645 $w=2.53e-07 $l=1.7e-07 $layer=LI1_cond $X=8.05 $Y=1.43
+ $X2=8.22 $Y2=1.43
r206 68 81 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.615 $Y=1.255
+ $X2=7.615 $Y2=1.09
r207 67 70 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.695 $Y=1.255
+ $X2=7.695 $Y2=1.335
r208 67 69 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.695 $Y=1.255
+ $X2=7.695 $Y2=1.09
r209 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.615
+ $Y=1.255 $X2=7.615 $Y2=1.255
r210 61 63 2.28037 $w=4.28e-07 $l=8e-08 $layer=LI1_cond $X=5.075 $Y=2.05
+ $X2=5.155 $Y2=2.05
r211 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.075
+ $Y=2.155 $X2=5.075 $Y2=2.155
r212 59 61 12.9696 $w=4.28e-07 $l=4.55e-07 $layer=LI1_cond $X=4.62 $Y=2.05
+ $X2=5.075 $Y2=2.05
r213 56 85 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.515 $Y=1.52
+ $X2=8.515 $Y2=1.685
r214 55 73 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=8.515 $Y=1.482
+ $X2=8.22 $Y2=1.482
r215 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.515
+ $Y=1.52 $X2=8.515 $Y2=1.52
r216 52 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.86 $Y=1.335
+ $X2=7.695 $Y2=1.335
r217 52 72 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=7.86 $Y=1.335
+ $X2=8.05 $Y2=1.335
r218 49 69 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=7.775 $Y=0.425
+ $X2=7.775 $Y2=1.09
r219 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.69 $Y=0.34
+ $X2=7.775 $Y2=0.425
r220 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.69 $Y=0.34
+ $X2=7.02 $Y2=0.34
r221 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.935 $Y=0.425
+ $X2=7.02 $Y2=0.34
r222 45 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.935 $Y=0.425
+ $X2=6.935 $Y2=0.69
r223 44 65 3.25423 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=6.035 $Y=0.775
+ $X2=5.892 $Y2=0.775
r224 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.85 $Y=0.775
+ $X2=6.935 $Y2=0.69
r225 43 44 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=6.85 $Y=0.775
+ $X2=6.035 $Y2=0.775
r226 41 76 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=5.87 $Y=1.195
+ $X2=5.71 $Y2=1.195
r227 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.87
+ $Y=1.195 $X2=5.87 $Y2=1.195
r228 38 65 3.29812 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=5.892 $Y=0.86
+ $X2=5.892 $Y2=0.775
r229 38 40 13.5463 $w=2.83e-07 $l=3.35e-07 $layer=LI1_cond $X=5.892 $Y=0.86
+ $X2=5.892 $Y2=1.195
r230 37 65 3.29812 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=5.892 $Y=0.69
+ $X2=5.892 $Y2=0.775
r231 36 37 10.7157 $w=2.83e-07 $l=2.65e-07 $layer=LI1_cond $X=5.892 $Y=0.425
+ $X2=5.892 $Y2=0.69
r232 35 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.24 $Y=0.34
+ $X2=5.155 $Y2=0.34
r233 34 36 7.39867 $w=1.7e-07 $l=1.79538e-07 $layer=LI1_cond $X=5.75 $Y=0.34
+ $X2=5.892 $Y2=0.425
r234 34 35 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.75 $Y=0.34
+ $X2=5.24 $Y2=0.34
r235 33 63 6.19161 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=5.155 $Y=1.82
+ $X2=5.155 $Y2=2.05
r236 32 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.155 $Y=0.425
+ $X2=5.155 $Y2=0.34
r237 32 33 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=5.155 $Y=0.425
+ $X2=5.155 $Y2=1.82
r238 30 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.07 $Y=0.34
+ $X2=5.155 $Y2=0.34
r239 30 31 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=5.07 $Y=0.34
+ $X2=4.445 $Y2=0.34
r240 26 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.32 $Y=0.425
+ $X2=4.445 $Y2=0.34
r241 26 28 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.32 $Y=0.425
+ $X2=4.32 $Y2=0.515
r242 24 25 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=8.395 $Y=2.02
+ $X2=8.395 $Y2=2.17
r243 24 85 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=8.425 $Y=2.02
+ $X2=8.425 $Y2=1.685
r244 20 25 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=8.38 $Y=2.75
+ $X2=8.38 $Y2=2.17
r245 16 81 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=7.57 $Y=0.645
+ $X2=7.57 $Y2=1.09
r246 11 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.71 $Y=1.03
+ $X2=5.71 $Y2=1.195
r247 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.71 $Y=1.03
+ $X2=5.71 $Y2=0.71
r248 7 62 56.2646 $w=2.57e-07 $l=3.73497e-07 $layer=POLY_cond $X=5.375 $Y=2.32
+ $X2=5.075 $Y2=2.155
r249 7 9 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=5.375 $Y=2.32
+ $X2=5.375 $Y2=2.69
r250 2 59 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=4.485
+ $Y=1.84 $X2=4.62 $Y2=2.02
r251 1 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.14
+ $Y=0.37 $X2=4.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_1%A_612_74# 1 2 9 11 13 15 16 20 22 28 32 35
+ 38 40 41 44 48 50 51 52 57 58 60 61 62 64 65 72 74 77 86 88
c214 77 0 1.40714e-19 $X=7.72 $Y=1.795
c215 74 0 2.55557e-20 $X=6.02 $Y=2.035
c216 52 0 6.77941e-20 $X=3.855 $Y=1.905
c217 44 0 5.43913e-20 $X=8.33 $Y=1.04
c218 20 0 1.67448e-19 $X=5.03 $Y=0.71
r219 78 88 22.6504 $w=2.66e-07 $l=1.25e-07 $layer=POLY_cond $X=7.72 $Y=1.795
+ $X2=7.845 $Y2=1.795
r220 77 80 8.46257 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=7.722 $Y=1.795
+ $X2=7.722 $Y2=1.96
r221 77 78 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.72
+ $Y=1.795 $X2=7.72 $Y2=1.795
r222 72 86 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.84 $Y=2.035
+ $X2=5.84 $Y2=2.2
r223 71 74 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=5.84 $Y=2.035
+ $X2=6.02 $Y2=2.035
r224 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.84
+ $Y=2.035 $X2=5.84 $Y2=2.035
r225 65 68 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.435 $Y=1.905
+ $X2=3.435 $Y2=2.02
r226 64 80 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.65 $Y=2.52
+ $X2=7.65 $Y2=1.96
r227 61 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.565 $Y=2.605
+ $X2=7.65 $Y2=2.52
r228 61 62 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=7.565 $Y=2.605
+ $X2=6.105 $Y2=2.605
r229 60 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.02 $Y=2.52
+ $X2=6.105 $Y2=2.605
r230 59 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.02 $Y=2.2
+ $X2=6.02 $Y2=2.035
r231 59 60 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.02 $Y=2.2 $X2=6.02
+ $Y2=2.52
r232 58 83 25.295 $w=3.65e-07 $l=1.6e-07 $layer=POLY_cond $X=3.957 $Y=1.515
+ $X2=3.957 $Y2=1.675
r233 58 82 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=3.957 $Y=1.515
+ $X2=3.957 $Y2=1.35
r234 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.94
+ $Y=1.515 $X2=3.94 $Y2=1.515
r235 55 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.94 $Y=1.82
+ $X2=3.94 $Y2=1.515
r236 54 57 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=3.94 $Y=1.01
+ $X2=3.94 $Y2=1.515
r237 53 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.6 $Y=1.905
+ $X2=3.435 $Y2=1.905
r238 52 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.855 $Y=1.905
+ $X2=3.94 $Y2=1.82
r239 52 53 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.855 $Y=1.905
+ $X2=3.6 $Y2=1.905
r240 50 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.855 $Y=0.925
+ $X2=3.94 $Y2=1.01
r241 50 51 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.855 $Y=0.925
+ $X2=3.365 $Y2=0.925
r242 46 51 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.2 $Y=0.84
+ $X2=3.365 $Y2=0.925
r243 46 48 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.2 $Y=0.84
+ $X2=3.2 $Y2=0.515
r244 42 44 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=8.065 $Y=1.04
+ $X2=8.33 $Y2=1.04
r245 36 44 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.33 $Y=0.965
+ $X2=8.33 $Y2=1.04
r246 36 38 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=8.33 $Y=0.965
+ $X2=8.33 $Y2=0.58
r247 35 88 39.8647 $w=2.66e-07 $l=2.91033e-07 $layer=POLY_cond $X=8.065 $Y=1.63
+ $X2=7.845 $Y2=1.795
r248 34 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.065 $Y=1.115
+ $X2=8.065 $Y2=1.04
r249 34 35 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=8.065 $Y=1.115
+ $X2=8.065 $Y2=1.63
r250 30 88 11.9456 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.845 $Y=1.96
+ $X2=7.845 $Y2=1.795
r251 30 32 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=7.845 $Y=1.96
+ $X2=7.845 $Y2=2.54
r252 28 86 190.468 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=5.825 $Y=2.69
+ $X2=5.825 $Y2=2.2
r253 24 72 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=5.84 $Y=1.75
+ $X2=5.84 $Y2=2.035
r254 23 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.105 $Y=1.675
+ $X2=5.03 $Y2=1.675
r255 22 24 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.675 $Y=1.675
+ $X2=5.84 $Y2=1.75
r256 22 23 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=5.675 $Y=1.675
+ $X2=5.105 $Y2=1.675
r257 18 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.03 $Y=1.6
+ $X2=5.03 $Y2=1.675
r258 18 20 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=5.03 $Y=1.6
+ $X2=5.03 $Y2=0.71
r259 17 40 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.485 $Y=1.675
+ $X2=4.395 $Y2=1.675
r260 16 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.955 $Y=1.675
+ $X2=5.03 $Y2=1.675
r261 16 17 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=4.955 $Y=1.675
+ $X2=4.485 $Y2=1.675
r262 13 40 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.395 $Y=1.75
+ $X2=4.395 $Y2=1.675
r263 13 15 174.056 $w=1.8e-07 $l=6.5e-07 $layer=POLY_cond $X=4.395 $Y=1.75
+ $X2=4.395 $Y2=2.4
r264 12 83 23.6381 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=4.14 $Y=1.675
+ $X2=3.957 $Y2=1.675
r265 11 40 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.305 $Y=1.675
+ $X2=4.395 $Y2=1.675
r266 11 12 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.305 $Y=1.675
+ $X2=4.14 $Y2=1.675
r267 9 82 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.065 $Y=0.74
+ $X2=4.065 $Y2=1.35
r268 2 68 600 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=1.84 $X2=3.435 $Y2=2.02
r269 1 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.06
+ $Y=0.37 $X2=3.2 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_1%A_1243_398# 1 2 7 9 13 16 17 20 22 23 27 33
c76 16 0 1.47351e-19 $X=6.305 $Y=1.99
r77 25 27 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=7.19 $Y=2.225
+ $X2=7.275 $Y2=2.225
r78 23 27 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.275 $Y=2.1
+ $X2=7.275 $Y2=2.225
r79 22 23 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=7.275 $Y=1.36
+ $X2=7.275 $Y2=2.1
r80 20 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.41 $Y=1.195
+ $X2=6.41 $Y2=1.36
r81 20 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.41 $Y=1.195
+ $X2=6.41 $Y2=1.03
r82 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.41
+ $Y=1.195 $X2=6.41 $Y2=1.195
r83 17 22 9.48765 $w=2.37e-07 $l=2.0106e-07 $layer=LI1_cond $X=7.355 $Y=1.195
+ $X2=7.275 $Y2=1.36
r84 17 30 24.7089 $w=2.37e-07 $l=4.8e-07 $layer=LI1_cond $X=7.355 $Y=1.195
+ $X2=7.355 $Y2=0.715
r85 17 19 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=7.19 $Y=1.195
+ $X2=6.41 $Y2=1.195
r86 16 34 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=6.32 $Y=1.99
+ $X2=6.32 $Y2=1.36
r87 13 33 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.32 $Y=0.71
+ $X2=6.32 $Y2=1.03
r88 7 16 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.305 $Y=2.08 $X2=6.305
+ $Y2=1.99
r89 7 9 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=6.305 $Y=2.08
+ $X2=6.305 $Y2=2.69
r90 2 25 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=7.015
+ $Y=2.12 $X2=7.19 $Y2=2.265
r91 1 30 182 $w=1.7e-07 $l=4.11157e-07 $layer=licon1_NDIFF $count=1 $X=7.21
+ $Y=0.37 $X2=7.355 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_1%A_1021_100# 1 2 9 13 17 21 23 25 26 28 37
c85 26 0 1.47351e-19 $X=5.587 $Y=2.46
r86 36 37 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=6.925 $Y=1.765
+ $X2=7.135 $Y2=1.765
r87 32 36 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=6.855 $Y=1.765
+ $X2=6.925 $Y2=1.765
r88 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.855
+ $Y=1.765 $X2=6.855 $Y2=1.765
r89 28 31 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=6.855 $Y=1.615
+ $X2=6.855 $Y2=1.765
r90 25 26 10.6092 $w=3.53e-07 $l=2.3e-07 $layer=LI1_cond $X=5.587 $Y=2.69
+ $X2=5.587 $Y2=2.46
r91 22 23 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.58 $Y=1.615
+ $X2=5.495 $Y2=1.615
r92 21 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.69 $Y=1.615
+ $X2=6.855 $Y2=1.615
r93 21 22 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=6.69 $Y=1.615
+ $X2=5.58 $Y2=1.615
r94 19 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.495 $Y=1.7
+ $X2=5.495 $Y2=1.615
r95 19 26 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=5.495 $Y=1.7
+ $X2=5.495 $Y2=2.46
r96 15 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.495 $Y=1.53
+ $X2=5.495 $Y2=1.615
r97 15 17 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=5.495 $Y=1.53
+ $X2=5.495 $Y2=0.765
r98 11 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.135 $Y=1.6
+ $X2=7.135 $Y2=1.765
r99 11 13 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=7.135 $Y=1.6
+ $X2=7.135 $Y2=0.645
r100 7 36 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.925 $Y=1.93
+ $X2=6.925 $Y2=1.765
r101 7 9 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=6.925 $Y=1.93
+ $X2=6.925 $Y2=2.54
r102 2 25 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=5.465
+ $Y=2.48 $X2=5.6 $Y2=2.69
r103 1 17 182 $w=1.7e-07 $l=5.05421e-07 $layer=licon1_NDIFF $count=1 $X=5.105
+ $Y=0.5 $X2=5.495 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_1%A_1723_48# 1 2 9 13 21 25 27 31 37 40 42 43
+ 44 45 48 50 55 58 63 64 66 68 69 71 73
c139 69 0 1.65961e-19 $X=9.775 $Y=1.94
c140 45 0 1.8865e-19 $X=9.6 $Y=2.235
c141 40 0 8.08518e-20 $X=8.965 $Y=1.07
c142 9 0 3.89393e-20 $X=8.69 $Y=0.58
r143 68 70 4.2805 $w=3.48e-07 $l=1.3e-07 $layer=LI1_cond $X=9.775 $Y=2.105
+ $X2=9.775 $Y2=2.235
r144 68 69 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=9.775 $Y=2.105
+ $X2=9.775 $Y2=1.94
r145 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.41
+ $Y=1.485 $X2=10.41 $Y2=1.485
r146 61 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.95 $Y=1.485
+ $X2=9.865 $Y2=1.485
r147 61 63 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=9.95 $Y=1.485
+ $X2=10.41 $Y2=1.485
r148 59 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.865 $Y=1.65
+ $X2=9.865 $Y2=1.485
r149 59 69 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=9.865 $Y=1.65
+ $X2=9.865 $Y2=1.94
r150 58 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.865 $Y=1.32
+ $X2=9.865 $Y2=1.485
r151 58 66 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=9.865 $Y=1.32
+ $X2=9.865 $Y2=0.93
r152 53 70 3.7866 $w=3.48e-07 $l=1.15e-07 $layer=LI1_cond $X=9.775 $Y=2.35
+ $X2=9.775 $Y2=2.235
r153 53 55 15.311 $w=3.48e-07 $l=4.65e-07 $layer=LI1_cond $X=9.775 $Y=2.35
+ $X2=9.775 $Y2=2.815
r154 50 66 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=9.77 $Y=0.75
+ $X2=9.77 $Y2=0.93
r155 50 52 3.72778 $w=3.6e-07 $l=1.1e-07 $layer=LI1_cond $X=9.77 $Y=0.75
+ $X2=9.77 $Y2=0.64
r156 48 74 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.875 $Y=2.215
+ $X2=8.875 $Y2=2.38
r157 48 73 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.875 $Y=2.215
+ $X2=8.875 $Y2=2.05
r158 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.875
+ $Y=2.215 $X2=8.875 $Y2=2.215
r159 45 70 3.19443 $w=2.3e-07 $l=1.75e-07 $layer=LI1_cond $X=9.6 $Y=2.235
+ $X2=9.775 $Y2=2.235
r160 45 47 36.327 $w=2.28e-07 $l=7.25e-07 $layer=LI1_cond $X=9.6 $Y=2.235
+ $X2=8.875 $Y2=2.235
r161 43 44 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=11.467 $Y=1.79
+ $X2=11.467 $Y2=1.94
r162 38 40 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=8.69 $Y=1.07
+ $X2=8.965 $Y2=1.07
r163 37 44 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=11.48 $Y=2.435
+ $X2=11.48 $Y2=1.94
r164 33 42 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.44 $Y=1.59
+ $X2=11.44 $Y2=1.455
r165 33 43 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=11.44 $Y=1.59
+ $X2=11.44 $Y2=1.79
r166 29 42 32.2453 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.44 $Y=1.32
+ $X2=11.44 $Y2=1.455
r167 29 31 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=11.44 $Y=1.32
+ $X2=11.44 $Y2=0.835
r168 28 64 5.72191 $w=2.7e-07 $l=1.27118e-07 $layer=POLY_cond $X=10.6 $Y=1.455
+ $X2=10.487 $Y2=1.485
r169 27 42 2.60871 $w=2.7e-07 $l=7.5e-08 $layer=POLY_cond $X=11.365 $Y=1.455
+ $X2=11.44 $Y2=1.455
r170 27 28 169.963 $w=2.7e-07 $l=7.65e-07 $layer=POLY_cond $X=11.365 $Y=1.455
+ $X2=10.6 $Y2=1.455
r171 23 64 19.9095 $w=1.8e-07 $l=1.76125e-07 $layer=POLY_cond $X=10.51 $Y=1.65
+ $X2=10.487 $Y2=1.485
r172 23 25 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=10.51 $Y=1.65
+ $X2=10.51 $Y2=2.4
r173 19 64 19.9095 $w=1.5e-07 $l=1.82565e-07 $layer=POLY_cond $X=10.45 $Y=1.32
+ $X2=10.487 $Y2=1.485
r174 19 21 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=10.45 $Y=1.32
+ $X2=10.45 $Y2=0.74
r175 15 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.965 $Y=1.145
+ $X2=8.965 $Y2=1.07
r176 15 73 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=8.965 $Y=1.145
+ $X2=8.965 $Y2=2.05
r177 13 74 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=8.8 $Y=2.75 $X2=8.8
+ $Y2=2.38
r178 7 38 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.69 $Y=0.995
+ $X2=8.69 $Y2=1.07
r179 7 9 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=8.69 $Y=0.995
+ $X2=8.69 $Y2=0.58
r180 2 68 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.63
+ $Y=1.96 $X2=9.765 $Y2=2.105
r181 2 55 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=9.63
+ $Y=1.96 $X2=9.765 $Y2=2.815
r182 1 52 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=9.535
+ $Y=0.37 $X2=9.675 $Y2=0.64
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_1%A_1529_74# 1 2 8 11 15 17 20 22 26 27 29 30
+ 31 33 34 38 42 44 48 49
c120 44 0 9.33306e-20 $X=8.935 $Y=1.065
c121 42 0 1.07508e-19 $X=8.475 $Y=0.58
c122 31 0 1.71252e-20 $X=8.56 $Y=1.065
r123 49 51 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.455 $Y=1.265
+ $X2=9.455 $Y2=1.1
r124 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.445
+ $Y=1.265 $X2=9.445 $Y2=1.265
r125 44 46 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=8.935 $Y=1.065
+ $X2=8.935 $Y2=1.185
r126 40 42 9.36061 $w=4.58e-07 $l=3.6e-07 $layer=LI1_cond $X=8.115 $Y=0.58
+ $X2=8.475 $Y2=0.58
r127 35 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.02 $Y=1.185
+ $X2=8.935 $Y2=1.185
r128 34 48 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.28 $Y=1.185
+ $X2=9.445 $Y2=1.185
r129 34 35 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=9.28 $Y=1.185
+ $X2=9.02 $Y2=1.185
r130 32 46 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=8.935 $Y=1.27
+ $X2=8.935 $Y2=1.185
r131 32 33 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.935 $Y=1.27
+ $X2=8.935 $Y2=1.78
r132 30 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.85 $Y=1.065
+ $X2=8.935 $Y2=1.065
r133 30 31 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=8.85 $Y=1.065
+ $X2=8.56 $Y2=1.065
r134 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.475 $Y=0.98
+ $X2=8.56 $Y2=1.065
r135 28 42 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=8.475 $Y=0.81
+ $X2=8.475 $Y2=0.58
r136 28 29 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.475 $Y=0.81
+ $X2=8.475 $Y2=0.98
r137 26 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.85 $Y=1.865
+ $X2=8.935 $Y2=1.78
r138 26 27 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=8.85 $Y=1.865
+ $X2=8.235 $Y2=1.865
r139 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.15 $Y=1.95
+ $X2=8.235 $Y2=1.865
r140 24 38 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.15 $Y=1.95
+ $X2=8.15 $Y2=2.13
r141 20 38 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.07 $Y=2.295
+ $X2=8.07 $Y2=2.13
r142 20 22 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=8.07 $Y=2.295
+ $X2=8.07 $Y2=2.815
r143 15 17 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=9.54 $Y=2.46
+ $X2=9.54 $Y2=1.77
r144 11 51 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=9.46 $Y=0.645
+ $X2=9.46 $Y2=1.1
r145 8 17 42.4214 $w=3.5e-07 $l=1.75e-07 $layer=POLY_cond $X=9.455 $Y=1.595
+ $X2=9.455 $Y2=1.77
r146 7 49 1.64869 $w=3.5e-07 $l=1e-08 $layer=POLY_cond $X=9.455 $Y=1.275
+ $X2=9.455 $Y2=1.265
r147 7 8 52.7581 $w=3.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.455 $Y=1.275
+ $X2=9.455 $Y2=1.595
r148 2 22 600 $w=1.7e-07 $l=7.59506e-07 $layer=licon1_PDIFF $count=1 $X=7.935
+ $Y=2.12 $X2=8.07 $Y2=2.815
r149 2 20 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=7.935
+ $Y=2.12 $X2=8.07 $Y2=2.295
r150 1 40 182 $w=1.7e-07 $l=5.65332e-07 $layer=licon1_NDIFF $count=1 $X=7.645
+ $Y=0.37 $X2=8.115 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_1%A_2216_112# 1 2 7 9 11 13 16 20 24 27
r49 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.89
+ $Y=1.385 $X2=11.89 $Y2=1.385
r50 22 27 0.153733 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=11.34 $Y=1.385
+ $X2=11.215 $Y2=1.385
r51 22 24 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=11.34 $Y=1.385
+ $X2=11.89 $Y2=1.385
r52 18 27 6.7841 $w=2.35e-07 $l=1.65e-07 $layer=LI1_cond $X=11.215 $Y=1.55
+ $X2=11.215 $Y2=1.385
r53 18 20 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=11.215 $Y=1.55
+ $X2=11.215 $Y2=2.16
r54 14 27 6.7841 $w=2.35e-07 $l=1.72337e-07 $layer=LI1_cond $X=11.2 $Y=1.22
+ $X2=11.215 $Y2=1.385
r55 14 16 20.1678 $w=2.18e-07 $l=3.85e-07 $layer=LI1_cond $X=11.2 $Y=1.22
+ $X2=11.2 $Y2=0.835
r56 11 25 38.5481 $w=3.01e-07 $l=2.03101e-07 $layer=POLY_cond $X=11.985 $Y=1.22
+ $X2=11.9 $Y2=1.385
r57 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=11.985 $Y=1.22
+ $X2=11.985 $Y2=0.74
r58 7 25 48.5617 $w=3.01e-07 $l=2.94449e-07 $layer=POLY_cond $X=11.985 $Y=1.64
+ $X2=11.9 $Y2=1.385
r59 7 9 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=11.985 $Y=1.64
+ $X2=11.985 $Y2=2.4
r60 2 20 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=11.13
+ $Y=2.015 $X2=11.255 $Y2=2.16
r61 1 16 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=11.08
+ $Y=0.56 $X2=11.225 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_1%VPWR 1 2 3 4 5 6 7 26 30 34 38 42 48 50 52
+ 57 62 67 72 77 84 85 88 91 98 101 104 107 110
r141 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r142 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r143 104 105 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r144 101 102 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r145 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r146 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r147 91 94 10.4403 $w=5.88e-07 $l=5.15e-07 $layer=LI1_cond $X=2.855 $Y=2.815
+ $X2=2.855 $Y2=3.33
r148 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r149 85 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r150 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r151 82 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.87 $Y=3.33
+ $X2=11.705 $Y2=3.33
r152 82 84 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=11.87 $Y=3.33
+ $X2=12.24 $Y2=3.33
r153 81 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r154 81 108 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.32 $Y2=3.33
r155 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r156 78 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.45 $Y=3.33
+ $X2=10.285 $Y2=3.33
r157 78 80 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=10.45 $Y=3.33
+ $X2=11.28 $Y2=3.33
r158 77 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.54 $Y=3.33
+ $X2=11.705 $Y2=3.33
r159 77 80 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=11.54 $Y=3.33
+ $X2=11.28 $Y2=3.33
r160 76 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r161 76 105 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=8.88 $Y2=3.33
r162 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r163 73 104 12.1981 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=9.43 $Y=3.33
+ $X2=9.145 $Y2=3.33
r164 73 75 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=9.43 $Y=3.33
+ $X2=9.84 $Y2=3.33
r165 72 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.12 $Y=3.33
+ $X2=10.285 $Y2=3.33
r166 72 75 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.12 $Y=3.33
+ $X2=9.84 $Y2=3.33
r167 71 105 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.88 $Y2=3.33
r168 71 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r169 70 71 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r170 68 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.78 $Y=3.33
+ $X2=6.615 $Y2=3.33
r171 68 70 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.78 $Y=3.33
+ $X2=6.96 $Y2=3.33
r172 67 104 12.1981 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=8.86 $Y=3.33
+ $X2=9.145 $Y2=3.33
r173 67 70 123.957 $w=1.68e-07 $l=1.9e-06 $layer=LI1_cond $X=8.86 $Y=3.33
+ $X2=6.96 $Y2=3.33
r174 66 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r175 65 66 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r176 63 98 11.3601 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=4.335 $Y=3.33
+ $X2=4.082 $Y2=3.33
r177 63 65 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=4.335 $Y=3.33
+ $X2=4.56 $Y2=3.33
r178 62 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.45 $Y=3.33
+ $X2=6.615 $Y2=3.33
r179 62 65 123.305 $w=1.68e-07 $l=1.89e-06 $layer=LI1_cond $X=6.45 $Y=3.33
+ $X2=4.56 $Y2=3.33
r180 61 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r181 61 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r182 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r183 58 94 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=3.15 $Y=3.33
+ $X2=2.855 $Y2=3.33
r184 58 60 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.15 $Y=3.33
+ $X2=3.6 $Y2=3.33
r185 57 98 11.3601 $w=1.7e-07 $l=2.52e-07 $layer=LI1_cond $X=3.83 $Y=3.33
+ $X2=4.082 $Y2=3.33
r186 57 60 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.83 $Y=3.33
+ $X2=3.6 $Y2=3.33
r187 56 95 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r188 56 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r189 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r190 53 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.03 $Y=3.33
+ $X2=0.865 $Y2=3.33
r191 53 55 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.03 $Y=3.33
+ $X2=1.2 $Y2=3.33
r192 52 94 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=2.56 $Y=3.33
+ $X2=2.855 $Y2=3.33
r193 52 55 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.56 $Y=3.33
+ $X2=1.2 $Y2=3.33
r194 50 102 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.24 $Y=3.33
+ $X2=6.48 $Y2=3.33
r195 50 66 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.24 $Y=3.33
+ $X2=4.56 $Y2=3.33
r196 46 110 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.705 $Y=3.245
+ $X2=11.705 $Y2=3.33
r197 46 48 37.8909 $w=3.28e-07 $l=1.085e-06 $layer=LI1_cond $X=11.705 $Y=3.245
+ $X2=11.705 $Y2=2.16
r198 42 45 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=10.285 $Y=1.985
+ $X2=10.285 $Y2=2.815
r199 40 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.285 $Y=3.245
+ $X2=10.285 $Y2=3.33
r200 40 45 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.285 $Y=3.245
+ $X2=10.285 $Y2=2.815
r201 36 104 2.39972 $w=5.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.145 $Y=3.245
+ $X2=9.145 $Y2=3.33
r202 36 38 9.02305 $w=5.68e-07 $l=4.3e-07 $layer=LI1_cond $X=9.145 $Y=3.245
+ $X2=9.145 $Y2=2.815
r203 32 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.615 $Y=3.245
+ $X2=6.615 $Y2=3.33
r204 32 34 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=6.615 $Y=3.245
+ $X2=6.615 $Y2=3.025
r205 28 98 2.09999 $w=5.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.082 $Y=3.245
+ $X2=4.082 $Y2=3.33
r206 28 30 10.1844 $w=5.03e-07 $l=4.3e-07 $layer=LI1_cond $X=4.082 $Y=3.245
+ $X2=4.082 $Y2=2.815
r207 24 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.865 $Y=3.245
+ $X2=0.865 $Y2=3.33
r208 24 26 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=0.865 $Y=3.245
+ $X2=0.865 $Y2=2.465
r209 7 48 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=11.57
+ $Y=2.015 $X2=11.705 $Y2=2.16
r210 6 45 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=10.16
+ $Y=1.84 $X2=10.285 $Y2=2.815
r211 6 42 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=10.16
+ $Y=1.84 $X2=10.285 $Y2=1.985
r212 5 38 600 $w=1.7e-07 $l=3.87137e-07 $layer=licon1_PDIFF $count=1 $X=8.89
+ $Y=2.54 $X2=9.16 $Y2=2.815
r213 4 34 600 $w=1.7e-07 $l=6.45697e-07 $layer=licon1_PDIFF $count=1 $X=6.395
+ $Y=2.48 $X2=6.615 $Y2=3.025
r214 3 30 600 $w=1.7e-07 $l=1.08392e-06 $layer=licon1_PDIFF $count=1 $X=3.85
+ $Y=1.84 $X2=4.08 $Y2=2.815
r215 2 91 600 $w=1.7e-07 $l=6.13351e-07 $layer=licon1_PDIFF $count=1 $X=2.59
+ $Y=2.32 $X2=2.855 $Y2=2.815
r216 1 26 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=0.68
+ $Y=2.32 $X2=0.865 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_1%A_296_74# 1 2 3 4 13 19 22 23 24 26 27 30
+ 31 32 35 37 38 41 44 45
c128 24 0 6.03804e-20 $X=2.39 $Y=1.265
c129 22 0 2.47416e-20 $X=2.305 $Y=1.18
r130 39 41 2.76586 $w=2.48e-07 $l=6e-08 $layer=LI1_cond $X=5.11 $Y=2.63 $X2=5.11
+ $Y2=2.69
r131 38 46 25.0585 $w=1.94e-07 $l=4.12129e-07 $layer=LI1_cond $X=4.675 $Y=2.545
+ $X2=4.28 $Y2=2.51
r132 37 39 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.985 $Y=2.545
+ $X2=5.11 $Y2=2.63
r133 37 38 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.985 $Y=2.545
+ $X2=4.675 $Y2=2.545
r134 33 35 32.9599 $w=2.48e-07 $l=7.15e-07 $layer=LI1_cond $X=4.775 $Y=1.48
+ $X2=4.775 $Y2=0.765
r135 31 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.65 $Y=1.565
+ $X2=4.775 $Y2=1.48
r136 31 32 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.65 $Y=1.565
+ $X2=4.365 $Y2=1.565
r137 30 46 1.50975 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.28 $Y=2.39
+ $X2=4.28 $Y2=2.51
r138 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.28 $Y=1.65
+ $X2=4.365 $Y2=1.565
r139 29 30 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=4.28 $Y=1.65
+ $X2=4.28 $Y2=2.39
r140 28 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=2.475
+ $X2=2.98 $Y2=2.475
r141 27 46 5.56362 $w=1.94e-07 $l=1.00995e-07 $layer=LI1_cond $X=4.195 $Y=2.475
+ $X2=4.28 $Y2=2.51
r142 27 28 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=4.195 $Y=2.475
+ $X2=3.065 $Y2=2.475
r143 26 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=2.39
+ $X2=2.98 $Y2=2.475
r144 25 26 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=2.98 $Y=1.35
+ $X2=2.98 $Y2=2.39
r145 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.895 $Y=1.265
+ $X2=2.98 $Y2=1.35
r146 23 24 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.895 $Y=1.265
+ $X2=2.39 $Y2=1.265
r147 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.305 $Y=1.18
+ $X2=2.39 $Y2=1.265
r148 21 22 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.305 $Y=0.64
+ $X2=2.305 $Y2=1.18
r149 20 44 4.79676 $w=1.7e-07 $l=1.86145e-07 $layer=LI1_cond $X=1.9 $Y=2.475
+ $X2=1.735 $Y2=2.43
r150 19 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=2.475
+ $X2=2.98 $Y2=2.475
r151 19 20 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=2.895 $Y=2.475
+ $X2=1.9 $Y2=2.475
r152 13 21 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.22 $Y=0.515
+ $X2=2.305 $Y2=0.64
r153 13 15 21.6659 $w=2.48e-07 $l=4.7e-07 $layer=LI1_cond $X=2.22 $Y=0.515
+ $X2=1.75 $Y2=0.515
r154 4 41 600 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_PDIFF $count=1 $X=5.02
+ $Y=2.48 $X2=5.15 $Y2=2.69
r155 3 44 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.6
+ $Y=2.32 $X2=1.735 $Y2=2.465
r156 2 35 182 $w=1.7e-07 $l=3.25576e-07 $layer=licon1_NDIFF $count=1 $X=4.68
+ $Y=0.5 $X2=4.815 $Y2=0.765
r157 1 15 182 $w=1.7e-07 $l=3.505e-07 $layer=licon1_NDIFF $count=1 $X=1.48
+ $Y=0.37 $X2=1.75 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_1%Q 1 2 7 9 15 16 17 23 29
r30 21 29 0.0555394 $w=4.13e-07 $l=2e-09 $layer=LI1_cond $X=10.707 $Y=0.923
+ $X2=10.707 $Y2=0.925
r31 17 31 8.68557 $w=4.13e-07 $l=1.64e-07 $layer=LI1_cond $X=10.707 $Y=0.966
+ $X2=10.707 $Y2=1.13
r32 17 29 1.13856 $w=4.13e-07 $l=4.1e-08 $layer=LI1_cond $X=10.707 $Y=0.966
+ $X2=10.707 $Y2=0.925
r33 17 21 1.16633 $w=4.13e-07 $l=4.2e-08 $layer=LI1_cond $X=10.707 $Y=0.881
+ $X2=10.707 $Y2=0.923
r34 16 17 9.05293 $w=4.13e-07 $l=3.26e-07 $layer=LI1_cond $X=10.707 $Y=0.555
+ $X2=10.707 $Y2=0.881
r35 16 23 1.11079 $w=4.13e-07 $l=4e-08 $layer=LI1_cond $X=10.707 $Y=0.555
+ $X2=10.707 $Y2=0.515
r36 15 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=10.83 $Y=1.82
+ $X2=10.83 $Y2=1.13
r37 9 11 36.0954 $w=2.63e-07 $l=8.3e-07 $layer=LI1_cond $X=10.782 $Y=1.985
+ $X2=10.782 $Y2=2.815
r38 7 15 7.21712 $w=2.63e-07 $l=1.32e-07 $layer=LI1_cond $X=10.782 $Y=1.952
+ $X2=10.782 $Y2=1.82
r39 7 9 1.43512 $w=2.63e-07 $l=3.3e-08 $layer=LI1_cond $X=10.782 $Y=1.952
+ $X2=10.782 $Y2=1.985
r40 2 11 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.6
+ $Y=1.84 $X2=10.735 $Y2=2.815
r41 2 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.6
+ $Y=1.84 $X2=10.735 $Y2=1.985
r42 1 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.525
+ $Y=0.37 $X2=10.665 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_1%Q_N 1 2 7 8 9 10 11 12 13 38 47
r19 23 47 1.52529 $w=3.38e-07 $l=4.5e-08 $layer=LI1_cond $X=12.205 $Y=0.88
+ $X2=12.205 $Y2=0.925
r20 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.21 $Y=2.405
+ $X2=12.21 $Y2=2.775
r21 11 38 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=12.21 $Y=1.967
+ $X2=12.21 $Y2=1.985
r22 11 51 6.4171 $w=3.28e-07 $l=1.47e-07 $layer=LI1_cond $X=12.21 $Y=1.967
+ $X2=12.21 $Y2=1.82
r23 11 12 12.3276 $w=3.28e-07 $l=3.53e-07 $layer=LI1_cond $X=12.21 $Y=2.052
+ $X2=12.21 $Y2=2.405
r24 11 38 2.33981 $w=3.28e-07 $l=6.7e-08 $layer=LI1_cond $X=12.21 $Y=2.052
+ $X2=12.21 $Y2=1.985
r25 10 51 8.11948 $w=2.18e-07 $l=1.55e-07 $layer=LI1_cond $X=12.265 $Y=1.665
+ $X2=12.265 $Y2=1.82
r26 9 10 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=12.265 $Y=1.295
+ $X2=12.265 $Y2=1.665
r27 9 49 12.834 $w=2.18e-07 $l=2.45e-07 $layer=LI1_cond $X=12.265 $Y=1.295
+ $X2=12.265 $Y2=1.05
r28 8 49 4.99175 $w=3.38e-07 $l=1.05e-07 $layer=LI1_cond $X=12.205 $Y=0.945
+ $X2=12.205 $Y2=1.05
r29 8 47 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=12.205 $Y=0.945
+ $X2=12.205 $Y2=0.925
r30 8 23 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=12.205 $Y=0.86
+ $X2=12.205 $Y2=0.88
r31 7 8 11.6939 $w=3.38e-07 $l=3.45e-07 $layer=LI1_cond $X=12.205 $Y=0.515
+ $X2=12.205 $Y2=0.86
r32 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=12.075
+ $Y=1.84 $X2=12.21 $Y2=2.815
r33 2 38 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=12.075
+ $Y=1.84 $X2=12.21 $Y2=1.985
r34 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.06
+ $Y=0.37 $X2=12.2 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFXBP_1%VGND 1 2 3 4 5 6 7 24 28 30 34 38 42 46 50
+ 53 54 55 57 62 67 72 84 93 94 97 100 103 106 109 112
r143 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r144 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r145 106 107 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r146 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r147 101 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.6 $Y2=0
r148 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r149 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r150 94 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r151 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r152 91 112 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=11.865 $Y=0
+ $X2=11.677 $Y2=0
r153 91 93 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.865 $Y=0
+ $X2=12.24 $Y2=0
r154 90 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r155 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r156 87 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=11.28 $Y2=0
r157 86 89 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=10.32 $Y=0 $X2=11.28
+ $Y2=0
r158 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r159 84 112 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=11.49 $Y=0
+ $X2=11.677 $Y2=0
r160 84 89 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=11.49 $Y=0
+ $X2=11.28 $Y2=0
r161 83 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r162 83 110 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=8.88 $Y2=0
r163 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r164 80 109 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=9.41 $Y=0
+ $X2=9.075 $Y2=0
r165 80 82 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=9.41 $Y=0 $X2=9.84
+ $Y2=0
r166 79 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r167 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r168 76 79 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=0 $X2=8.4
+ $Y2=0
r169 76 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=6.48 $Y2=0
r170 75 78 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.96 $Y=0 $X2=8.4
+ $Y2=0
r171 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r172 73 106 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.68 $Y=0
+ $X2=6.555 $Y2=0
r173 73 75 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=6.68 $Y=0 $X2=6.96
+ $Y2=0
r174 72 109 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=8.74 $Y=0
+ $X2=9.075 $Y2=0
r175 72 78 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=8.74 $Y=0 $X2=8.4
+ $Y2=0
r176 71 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r177 70 71 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r178 68 103 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.935 $Y=0
+ $X2=3.765 $Y2=0
r179 68 70 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.935 $Y=0
+ $X2=4.08 $Y2=0
r180 67 106 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.43 $Y=0
+ $X2=6.555 $Y2=0
r181 67 70 153.316 $w=1.68e-07 $l=2.35e-06 $layer=LI1_cond $X=6.43 $Y=0 $X2=4.08
+ $Y2=0
r182 66 101 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0
+ $X2=2.64 $Y2=0
r183 66 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r184 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r185 63 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=0 $X2=0.8
+ $Y2=0
r186 63 65 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.965 $Y=0 $X2=1.2
+ $Y2=0
r187 62 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.615 $Y=0
+ $X2=2.74 $Y2=0
r188 62 65 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=2.615 $Y=0
+ $X2=1.2 $Y2=0
r189 60 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r190 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r191 57 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.635 $Y=0 $X2=0.8
+ $Y2=0
r192 57 59 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=0
+ $X2=0.24 $Y2=0
r193 55 107 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.24 $Y=0
+ $X2=6.48 $Y2=0
r194 55 71 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=6.24 $Y=0
+ $X2=4.08 $Y2=0
r195 54 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.235 $Y=0
+ $X2=10.32 $Y2=0
r196 53 82 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.15 $Y=0 $X2=9.84
+ $Y2=0
r197 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.15 $Y=0
+ $X2=10.235 $Y2=0
r198 48 112 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=11.677 $Y=0.085
+ $X2=11.677 $Y2=0
r199 48 50 13.2147 $w=3.73e-07 $l=4.3e-07 $layer=LI1_cond $X=11.677 $Y=0.085
+ $X2=11.677 $Y2=0.515
r200 44 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.235 $Y=0.085
+ $X2=10.235 $Y2=0
r201 44 46 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=10.235 $Y=0.085
+ $X2=10.235 $Y2=0.515
r202 40 109 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.075 $Y=0.085
+ $X2=9.075 $Y2=0
r203 40 42 8.8367 $w=6.68e-07 $l=4.95e-07 $layer=LI1_cond $X=9.075 $Y=0.085
+ $X2=9.075 $Y2=0.58
r204 36 106 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.555 $Y=0.085
+ $X2=6.555 $Y2=0
r205 36 38 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=6.555 $Y=0.085
+ $X2=6.555 $Y2=0.355
r206 32 103 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.765 $Y=0.085
+ $X2=3.765 $Y2=0
r207 32 34 14.2361 $w=3.38e-07 $l=4.2e-07 $layer=LI1_cond $X=3.765 $Y=0.085
+ $X2=3.765 $Y2=0.505
r208 31 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.865 $Y=0
+ $X2=2.74 $Y2=0
r209 30 103 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.595 $Y=0
+ $X2=3.765 $Y2=0
r210 30 31 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.595 $Y=0
+ $X2=2.865 $Y2=0
r211 26 100 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.74 $Y=0.085
+ $X2=2.74 $Y2=0
r212 26 28 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=2.74 $Y=0.085
+ $X2=2.74 $Y2=0.58
r213 22 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=0.085 $X2=0.8
+ $Y2=0
r214 22 24 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.8 $Y=0.085
+ $X2=0.8 $Y2=0.58
r215 7 50 91 $w=1.7e-07 $l=2.56515e-07 $layer=licon1_NDIFF $count=2 $X=11.515
+ $Y=0.56 $X2=11.75 $Y2=0.515
r216 6 46 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=10.09
+ $Y=0.37 $X2=10.235 $Y2=0.515
r217 5 42 91 $w=1.7e-07 $l=5.755e-07 $layer=licon1_NDIFF $count=2 $X=8.765
+ $Y=0.37 $X2=9.245 $Y2=0.58
r218 4 38 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=6.395
+ $Y=0.5 $X2=6.595 $Y2=0.355
r219 3 34 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=3.615
+ $Y=0.36 $X2=3.765 $Y2=0.505
r220 2 28 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=2.56
+ $Y=0.37 $X2=2.74 $Y2=0.58
r221 1 24 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=0.59
+ $Y=0.37 $X2=0.8 $Y2=0.58
.ends


* File: sky130_fd_sc_ms__fah_2.pex.spice
* Created: Fri Aug 28 17:35:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__FAH_2%A_81_260# 1 2 9 13 16 19 24 27 30 33
c60 30 0 1.98792e-19 $X=1.31 $Y=1.465
c61 16 0 1.11723e-19 $X=0.532 $Y=1.465
r62 33 35 16.3735 $w=4.78e-07 $l=4.45e-07 $layer=LI1_cond $X=1.465 $Y=0.675
+ $X2=1.465 $Y2=1.12
r63 29 30 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.215 $Y=1.465
+ $X2=1.31 $Y2=1.465
r64 26 29 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.985 $Y=1.465
+ $X2=1.215 $Y2=1.465
r65 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.985
+ $Y=1.465 $X2=0.985 $Y2=1.465
r66 24 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.31 $Y=1.3 $X2=1.31
+ $Y2=1.465
r67 24 35 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.31 $Y=1.3 $X2=1.31
+ $Y2=1.12
r68 19 21 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=1.215 $Y=2.105
+ $X2=1.215 $Y2=2.815
r69 17 29 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=1.215 $Y=1.63
+ $X2=1.215 $Y2=1.465
r70 17 19 21.8964 $w=2.48e-07 $l=4.75e-07 $layer=LI1_cond $X=1.215 $Y=1.63
+ $X2=1.215 $Y2=2.105
r71 15 27 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=0.66 $Y=1.465
+ $X2=0.985 $Y2=1.465
r72 15 16 3.90195 $w=3.3e-07 $l=1.28e-07 $layer=POLY_cond $X=0.66 $Y=1.465
+ $X2=0.532 $Y2=1.465
r73 11 16 34.7346 $w=1.65e-07 $l=1.89658e-07 $layer=POLY_cond $X=0.585 $Y=1.3
+ $X2=0.532 $Y2=1.465
r74 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.585 $Y=1.3
+ $X2=0.585 $Y2=0.74
r75 7 16 34.7346 $w=1.65e-07 $l=1.82565e-07 $layer=POLY_cond $X=0.495 $Y=1.63
+ $X2=0.532 $Y2=1.465
r76 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.495 $Y=1.63
+ $X2=0.495 $Y2=2.4
r77 2 21 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.96 $X2=1.255 $Y2=2.815
r78 2 19 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.96 $X2=1.255 $Y2=2.105
r79 1 33 91 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=2 $X=1.395
+ $Y=0.525 $X2=1.54 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_2%A 3 5 7 10 12 14 15 22 24
c60 10 0 2.05287e-19 $X=1.99 $Y=2.46
c61 5 0 2.24154e-20 $X=1.825 $Y=1.29
c62 3 0 8.42529e-20 $X=1.48 $Y=2.46
r63 23 24 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=1.99 $Y=1.455
+ $X2=2.255 $Y2=1.455
r64 21 23 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.915 $Y=1.455
+ $X2=1.99 $Y2=1.455
r65 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.915
+ $Y=1.455 $X2=1.915 $Y2=1.455
r66 19 21 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.825 $Y=1.455
+ $X2=1.915 $Y2=1.455
r67 17 19 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=1.48 $Y=1.455
+ $X2=1.825 $Y2=1.455
r68 15 22 5.73629 $w=4.88e-07 $l=2.35e-07 $layer=LI1_cond $X=1.68 $Y=1.535
+ $X2=1.915 $Y2=1.535
r69 12 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=1.29
+ $X2=2.255 $Y2=1.455
r70 12 14 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.255 $Y=1.29
+ $X2=2.255 $Y2=0.845
r71 8 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.99 $Y=1.62
+ $X2=1.99 $Y2=1.455
r72 8 10 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=1.99 $Y=1.62 $X2=1.99
+ $Y2=2.46
r73 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=1.29
+ $X2=1.825 $Y2=1.455
r74 5 7 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.825 $Y=1.29
+ $X2=1.825 $Y2=0.845
r75 1 17 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.48 $Y=1.62
+ $X2=1.48 $Y2=1.455
r76 1 3 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=1.48 $Y=1.62 $X2=1.48
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_2%B 3 7 11 14 16 18 19 20 23 27 28 31 35 36 38
+ 41 42 43 46 47 48 50 51 52 54 55 56 62 63 73
c214 62 0 4.67017e-20 $X=2.64 $Y=1.665
c215 55 0 1.90307e-19 $X=4.5 $Y=0.68
c216 51 0 1.75179e-20 $X=3.605 $Y=1.795
c217 43 0 1.42825e-19 $X=5.435 $Y=1.005
c218 42 0 5.25489e-20 $X=5.875 $Y=1.005
c219 35 0 3.17652e-19 $X=4.505 $Y=1.44
c220 23 0 9.95712e-20 $X=7.125 $Y=0.74
c221 20 0 1.6052e-19 $X=6.745 $Y=1.315
c222 19 0 1.97436e-19 $X=7.05 $Y=1.315
r223 62 63 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.725 $Y=1.665
+ $X2=2.725 $Y2=2.035
r224 60 77 56.0359 $w=5.29e-07 $l=6.15e-07 $layer=POLY_cond $X=6.04 $Y=1.387
+ $X2=6.655 $Y2=1.387
r225 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.04
+ $Y=1.085 $X2=6.04 $Y2=1.085
r226 56 59 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=6.04 $Y=1.005 $X2=6.04
+ $Y2=1.085
r227 51 71 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.605 $Y=1.795
+ $X2=3.605 $Y2=1.96
r228 50 52 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.605 $Y=1.795
+ $X2=3.605 $Y2=1.63
r229 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.605
+ $Y=1.795 $X2=3.605 $Y2=1.795
r230 47 67 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.52
+ $X2=2.705 $Y2=1.355
r231 46 48 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=1.52
+ $X2=2.725 $Y2=1.355
r232 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.705
+ $Y=1.52 $X2=2.705 $Y2=1.52
r233 44 62 4.74535 $w=3.38e-07 $l=1.4e-07 $layer=LI1_cond $X=2.725 $Y=1.525
+ $X2=2.725 $Y2=1.665
r234 44 46 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=2.725 $Y=1.525
+ $X2=2.725 $Y2=1.52
r235 42 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.875 $Y=1.005
+ $X2=6.04 $Y2=1.005
r236 42 43 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.875 $Y=1.005
+ $X2=5.435 $Y2=1.005
r237 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.35 $Y=0.92
+ $X2=5.435 $Y2=1.005
r238 40 41 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.35 $Y=0.765
+ $X2=5.35 $Y2=0.92
r239 39 55 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.595 $Y=0.68
+ $X2=4.5 $Y2=0.68
r240 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.265 $Y=0.68
+ $X2=5.35 $Y2=0.765
r241 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.265 $Y=0.68
+ $X2=4.595 $Y2=0.68
r242 36 73 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.505 $Y=1.44
+ $X2=4.505 $Y2=1.275
r243 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.505
+ $Y=1.44 $X2=4.505 $Y2=1.44
r244 33 55 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.5 $Y=0.765
+ $X2=4.5 $Y2=0.68
r245 33 35 39.4019 $w=1.88e-07 $l=6.75e-07 $layer=LI1_cond $X=4.5 $Y=0.765
+ $X2=4.5 $Y2=1.44
r246 32 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.735 $Y=0.68
+ $X2=3.65 $Y2=0.68
r247 31 55 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.405 $Y=0.68
+ $X2=4.5 $Y2=0.68
r248 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.405 $Y=0.68
+ $X2=3.735 $Y2=0.68
r249 29 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.65 $Y=0.765
+ $X2=3.65 $Y2=0.68
r250 29 52 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=3.65 $Y=0.765
+ $X2=3.65 $Y2=1.63
r251 27 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.565 $Y=0.68
+ $X2=3.65 $Y2=0.68
r252 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.565 $Y=0.68
+ $X2=2.895 $Y2=0.68
r253 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.81 $Y=0.765
+ $X2=2.895 $Y2=0.68
r254 25 48 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.81 $Y=0.765
+ $X2=2.81 $Y2=1.355
r255 21 23 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=7.125 $Y=1.24
+ $X2=7.125 $Y2=0.74
r256 20 77 35.8501 $w=5.29e-07 $l=1.20748e-07 $layer=POLY_cond $X=6.745 $Y=1.315
+ $X2=6.655 $Y2=1.387
r257 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.05 $Y=1.315
+ $X2=7.125 $Y2=1.24
r258 19 20 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=7.05 $Y=1.315
+ $X2=6.745 $Y2=1.315
r259 16 77 28.2554 $w=1.8e-07 $l=3.78e-07 $layer=POLY_cond $X=6.655 $Y=1.765
+ $X2=6.655 $Y2=1.387
r260 16 18 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=6.655 $Y=1.765
+ $X2=6.655 $Y2=2.4
r261 12 60 34.1682 $w=5.29e-07 $l=6.28111e-07 $layer=POLY_cond $X=5.665 $Y=1.855
+ $X2=6.04 $Y2=1.387
r262 12 14 266.266 $w=1.8e-07 $l=6.85e-07 $layer=POLY_cond $X=5.665 $Y=1.855
+ $X2=5.665 $Y2=2.54
r263 11 73 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.445 $Y=0.845
+ $X2=4.445 $Y2=1.275
r264 7 71 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=3.56 $Y=2.54
+ $X2=3.56 $Y2=1.96
r265 3 67 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.685 $Y=0.845
+ $X2=2.685 $Y2=1.355
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_2%A_481_379# 1 2 7 9 10 11 13 14 16 17 18 20 21
+ 23 24 28 32 33 34 36 39 40 42 45 46 54
c166 54 0 5.91111e-20 $X=6.88 $Y=1.845
c167 36 0 8.21497e-20 $X=6.715 $Y=1.845
c168 33 0 1.61089e-19 $X=5.2 $Y=1.42
c169 24 0 1.90025e-19 $X=5.035 $Y=1.92
c170 17 0 1.56563e-19 $X=3.98 $Y=1.315
r171 54 56 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=6.88 $Y=1.845
+ $X2=6.88 $Y2=1.985
r172 45 48 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=5.235 $Y=1.765
+ $X2=5.235 $Y2=1.845
r173 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.2
+ $Y=1.765 $X2=5.2 $Y2=1.765
r174 40 42 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=7.34 $Y=1.19
+ $X2=7.34 $Y2=0.795
r175 39 54 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=6.88 $Y=1.76
+ $X2=6.88 $Y2=1.845
r176 38 40 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=6.88 $Y=1.275
+ $X2=7.34 $Y2=1.275
r177 38 39 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=6.88 $Y=1.36 $X2=6.88
+ $Y2=1.76
r178 37 48 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.365 $Y=1.845
+ $X2=5.235 $Y2=1.845
r179 36 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.715 $Y=1.845
+ $X2=6.88 $Y2=1.845
r180 36 37 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=6.715 $Y=1.845
+ $X2=5.365 $Y2=1.845
r181 35 46 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=5.2 $Y=1.845 $X2=5.2
+ $Y2=1.765
r182 33 46 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=5.2 $Y=1.42
+ $X2=5.2 $Y2=1.765
r183 33 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.2 $Y=1.42
+ $X2=5.2 $Y2=1.255
r184 29 31 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.155 $Y=1.315
+ $X2=3.445 $Y2=1.315
r185 28 34 131.747 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=5.29 $Y=0.845
+ $X2=5.29 $Y2=1.255
r186 25 32 6.66866 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=4.26 $Y=1.92
+ $X2=4.12 $Y2=1.92
r187 24 35 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.035 $Y=1.92
+ $X2=5.2 $Y2=1.845
r188 24 25 397.394 $w=1.5e-07 $l=7.75e-07 $layer=POLY_cond $X=5.035 $Y=1.92
+ $X2=4.26 $Y2=1.92
r189 21 32 18.8402 $w=1.65e-07 $l=9.68246e-08 $layer=POLY_cond $X=4.17 $Y=1.995
+ $X2=4.12 $Y2=1.92
r190 21 23 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=4.17 $Y=1.995
+ $X2=4.17 $Y2=2.54
r191 20 32 18.8402 $w=1.65e-07 $l=1.0247e-07 $layer=POLY_cond $X=4.055 $Y=1.845
+ $X2=4.12 $Y2=1.92
r192 19 20 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.055 $Y=1.39
+ $X2=4.055 $Y2=1.845
r193 18 31 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.52 $Y=1.315
+ $X2=3.445 $Y2=1.315
r194 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.98 $Y=1.315
+ $X2=4.055 $Y2=1.39
r195 17 18 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=3.98 $Y=1.315
+ $X2=3.52 $Y2=1.315
r196 14 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.445 $Y=1.24
+ $X2=3.445 $Y2=1.315
r197 14 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.445 $Y=1.24
+ $X2=3.445 $Y2=0.845
r198 12 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.155 $Y=1.39
+ $X2=3.155 $Y2=1.315
r199 12 13 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.155 $Y=1.39
+ $X2=3.155 $Y2=1.895
r200 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.08 $Y=1.97
+ $X2=3.155 $Y2=1.895
r201 10 11 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.08 $Y=1.97
+ $X2=2.585 $Y2=1.97
r202 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.495 $Y=2.045
+ $X2=2.585 $Y2=1.97
r203 7 9 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=2.495 $Y=2.045
+ $X2=2.495 $Y2=2.54
r204 2 56 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.84 $X2=6.88 $Y2=1.985
r205 1 42 182 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_NDIFF $count=1 $X=7.2
+ $Y=0.37 $X2=7.34 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_2%A_517_424# 1 2 9 13 17 21 23 28 29 32 33 34 35
+ 38 40 41 42 45 46 48 53 54 55 57 59 65 66 71 72 75 76 78 79 80 85 86
c250 71 0 1.01409e-19 $X=7.34 $Y=1.795
c251 46 0 3.062e-19 $X=8.575 $Y=1.39
c252 23 0 1.53607e-19 $X=3.065 $Y=2.555
c253 21 0 1.00227e-19 $X=10.285 $Y=0.715
r254 86 99 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.375 $Y=1.52
+ $X2=10.375 $Y2=1.355
r255 85 86 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.375
+ $Y=1.52 $X2=10.375 $Y2=1.52
r256 82 85 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=10.17 $Y=1.52
+ $X2=10.375 $Y2=1.52
r257 79 97 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.475 $Y=1.795
+ $X2=9.475 $Y2=1.96
r258 78 81 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.41 $Y=1.795
+ $X2=9.41 $Y2=1.96
r259 78 80 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.41 $Y=1.795
+ $X2=9.41 $Y2=1.63
r260 78 79 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.475
+ $Y=1.795 $X2=9.475 $Y2=1.795
r261 72 88 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=7.34 $Y=1.795
+ $X2=7.18 $Y2=1.795
r262 71 74 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=7.36 $Y=1.795
+ $X2=7.36 $Y2=1.96
r263 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.34
+ $Y=1.795 $X2=7.34 $Y2=1.795
r264 66 68 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.31 $Y=2.185
+ $X2=6.31 $Y2=2.325
r265 64 65 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.285 $Y=2.555
+ $X2=3.45 $Y2=2.555
r266 62 64 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.15 $Y=2.555
+ $X2=3.285 $Y2=2.555
r267 59 61 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.23 $Y=1.02
+ $X2=3.23 $Y2=1.185
r268 57 82 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.17 $Y=1.355
+ $X2=10.17 $Y2=1.52
r269 56 57 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=10.17 $Y=0.765
+ $X2=10.17 $Y2=1.355
r270 54 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.085 $Y=0.68
+ $X2=10.17 $Y2=0.765
r271 54 55 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.085 $Y=0.68
+ $X2=9.415 $Y2=0.68
r272 53 81 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=9.49 $Y=2.905
+ $X2=9.49 $Y2=1.96
r273 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.33 $Y=0.765
+ $X2=9.415 $Y2=0.68
r274 50 80 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=9.33 $Y=0.765
+ $X2=9.33 $Y2=1.63
r275 49 76 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=8.735 $Y=2.99
+ $X2=8.607 $Y2=2.99
r276 48 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.405 $Y=2.99
+ $X2=9.49 $Y2=2.905
r277 48 49 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.405 $Y=2.99
+ $X2=8.735 $Y2=2.99
r278 46 93 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.575 $Y=1.39
+ $X2=8.575 $Y2=1.225
r279 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.575
+ $Y=1.39 $X2=8.575 $Y2=1.39
r280 43 76 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=8.607 $Y=2.905
+ $X2=8.607 $Y2=2.99
r281 43 45 68.4687 $w=2.53e-07 $l=1.515e-06 $layer=LI1_cond $X=8.607 $Y=2.905
+ $X2=8.607 $Y2=1.39
r282 41 76 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=8.48 $Y=2.99
+ $X2=8.607 $Y2=2.99
r283 41 42 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=8.48 $Y=2.99
+ $X2=7.385 $Y2=2.99
r284 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.3 $Y=2.905
+ $X2=7.385 $Y2=2.99
r285 39 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.3 $Y=2.41 $X2=7.3
+ $Y2=2.325
r286 39 40 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=7.3 $Y=2.41
+ $X2=7.3 $Y2=2.905
r287 38 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.3 $Y=2.24 $X2=7.3
+ $Y2=2.325
r288 38 74 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.3 $Y=2.24 $X2=7.3
+ $Y2=1.96
r289 36 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.395 $Y=2.325
+ $X2=6.31 $Y2=2.325
r290 35 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.215 $Y=2.325
+ $X2=7.3 $Y2=2.325
r291 35 36 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=7.215 $Y=2.325
+ $X2=6.395 $Y2=2.325
r292 33 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.225 $Y=2.185
+ $X2=6.31 $Y2=2.185
r293 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.225 $Y=2.185
+ $X2=5.555 $Y2=2.185
r294 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.47 $Y=2.27
+ $X2=5.555 $Y2=2.185
r295 31 32 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.47 $Y=2.27
+ $X2=5.47 $Y2=2.55
r296 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.385 $Y=2.635
+ $X2=5.47 $Y2=2.55
r297 29 65 126.241 $w=1.68e-07 $l=1.935e-06 $layer=LI1_cond $X=5.385 $Y=2.635
+ $X2=3.45 $Y2=2.635
r298 28 62 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.15 $Y=2.39
+ $X2=3.15 $Y2=2.555
r299 28 61 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=3.15 $Y=2.39
+ $X2=3.15 $Y2=1.185
r300 23 62 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=2.555
+ $X2=3.15 $Y2=2.555
r301 23 25 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.065 $Y=2.555
+ $X2=2.72 $Y2=2.555
r302 21 99 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=10.285 $Y=0.715
+ $X2=10.285 $Y2=1.355
r303 17 97 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=9.4 $Y=2.54 $X2=9.4
+ $Y2=1.96
r304 13 93 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=8.625 $Y=0.715
+ $X2=8.625 $Y2=1.225
r305 7 88 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.18 $Y=1.96
+ $X2=7.18 $Y2=1.795
r306 7 9 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=7.18 $Y=1.96 $X2=7.18
+ $Y2=2.54
r307 2 64 600 $w=1.7e-07 $l=8.91347e-07 $layer=licon1_PDIFF $count=1 $X=2.585
+ $Y=2.12 $X2=3.285 $Y2=2.555
r308 2 25 600 $w=1.7e-07 $l=4.97946e-07 $layer=licon1_PDIFF $count=1 $X=2.585
+ $Y=2.12 $X2=2.72 $Y2=2.555
r309 1 59 182 $w=1.7e-07 $l=6.9114e-07 $layer=licon1_NDIFF $count=1 $X=2.76
+ $Y=0.525 $X2=3.23 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_2%A_852_424# 1 2 7 9 10 11 14 16 19 20 21 24 26
+ 29 30 32 36 37 38 46 49 51 53 56 57 58 60 61 62 65 67 71 75 76 80
c200 80 0 2.97007e-19 $X=7.822 $Y=1.275
c201 71 0 1.90025e-19 $X=4.93 $Y=1.02
c202 53 0 2.83882e-20 $X=6.375 $Y=1.44
c203 24 0 1.66419e-19 $X=9.455 $Y=0.715
c204 7 0 1.77494e-19 $X=7.6 $Y=1.11
c205 1 0 1.90307e-19 $X=4.52 $Y=0.525
r206 76 78 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=5.62 $Y=1.345
+ $X2=5.62 $Y2=1.44
r207 73 74 5.66838 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.93 $Y=1.345
+ $X2=4.93 $Y2=1.43
r208 71 73 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.93 $Y=1.02
+ $X2=4.93 $Y2=1.345
r209 67 68 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.88
+ $Y=1.44 $X2=7.88 $Y2=1.44
r210 65 80 7.79447 $w=2.93e-07 $l=1.47e-07 $layer=LI1_cond $X=7.822 $Y=1.422
+ $X2=7.822 $Y2=1.275
r211 65 67 0.703186 $w=2.93e-07 $l=1.8e-08 $layer=LI1_cond $X=7.822 $Y=1.422
+ $X2=7.822 $Y2=1.44
r212 63 80 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=7.76 $Y=0.425
+ $X2=7.76 $Y2=1.275
r213 61 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.675 $Y=0.34
+ $X2=7.76 $Y2=0.425
r214 61 62 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.675 $Y=0.34
+ $X2=7.005 $Y2=0.34
r215 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.92 $Y=0.425
+ $X2=7.005 $Y2=0.34
r216 59 60 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=6.92 $Y=0.425
+ $X2=6.92 $Y2=0.85
r217 57 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.835 $Y=0.935
+ $X2=6.92 $Y2=0.85
r218 57 58 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.835 $Y=0.935
+ $X2=6.545 $Y2=0.935
r219 55 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.46 $Y=1.02
+ $X2=6.545 $Y2=0.935
r220 55 56 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.46 $Y=1.02
+ $X2=6.46 $Y2=1.355
r221 54 78 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.705 $Y=1.44
+ $X2=5.62 $Y2=1.44
r222 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.375 $Y=1.44
+ $X2=6.46 $Y2=1.355
r223 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.375 $Y=1.44
+ $X2=5.705 $Y2=1.44
r224 52 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.095 $Y=1.345
+ $X2=4.93 $Y2=1.345
r225 51 76 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.535 $Y=1.345
+ $X2=5.62 $Y2=1.345
r226 51 52 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.535 $Y=1.345
+ $X2=5.095 $Y2=1.345
r227 47 75 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.935 $Y=2.225
+ $X2=4.85 $Y2=2.225
r228 47 49 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=4.935 $Y=2.225
+ $X2=5.05 $Y2=2.225
r229 46 75 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.85 $Y=2.1
+ $X2=4.85 $Y2=2.225
r230 46 74 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.85 $Y=2.1
+ $X2=4.85 $Y2=1.43
r231 36 68 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=7.88 $Y=1.795
+ $X2=7.88 $Y2=1.44
r232 30 39 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=10.185 $Y=1.97
+ $X2=9.925 $Y2=1.97
r233 30 32 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=10.185 $Y=2.045
+ $X2=10.185 $Y2=2.54
r234 29 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.925 $Y=1.895
+ $X2=9.925 $Y2=1.97
r235 28 29 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=9.925 $Y=1.39
+ $X2=9.925 $Y2=1.895
r236 27 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.53 $Y=1.315
+ $X2=9.455 $Y2=1.315
r237 26 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.85 $Y=1.315
+ $X2=9.925 $Y2=1.39
r238 26 27 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.85 $Y=1.315
+ $X2=9.53 $Y2=1.315
r239 22 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.455 $Y=1.24
+ $X2=9.455 $Y2=1.315
r240 22 24 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=9.455 $Y=1.24
+ $X2=9.455 $Y2=0.715
r241 20 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.38 $Y=1.315
+ $X2=9.455 $Y2=1.315
r242 20 21 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=9.38 $Y=1.315
+ $X2=9.1 $Y2=1.315
r243 18 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.025 $Y=1.39
+ $X2=9.1 $Y2=1.315
r244 18 19 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=9.025 $Y=1.39
+ $X2=9.025 $Y2=1.795
r245 17 37 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.46 $Y=1.87 $X2=8.37
+ $Y2=1.87
r246 16 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.95 $Y=1.87
+ $X2=9.025 $Y2=1.795
r247 16 17 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=8.95 $Y=1.87
+ $X2=8.46 $Y2=1.87
r248 12 37 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=8.37 $Y=1.945
+ $X2=8.37 $Y2=1.87
r249 12 14 231.282 $w=1.8e-07 $l=5.95e-07 $layer=POLY_cond $X=8.37 $Y=1.945
+ $X2=8.37 $Y2=2.54
r250 11 36 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=8.045 $Y=1.87
+ $X2=7.88 $Y2=1.795
r251 10 37 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.28 $Y=1.87 $X2=8.37
+ $Y2=1.87
r252 10 11 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=8.28 $Y=1.87
+ $X2=8.045 $Y2=1.87
r253 7 68 65.1981 $w=2.07e-07 $l=3.52987e-07 $layer=POLY_cond $X=7.6 $Y=1.11
+ $X2=7.88 $Y2=1.275
r254 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=7.6 $Y=1.11 $X2=7.6
+ $Y2=0.715
r255 2 49 300 $w=1.7e-07 $l=8.59448e-07 $layer=licon1_PDIFF $count=2 $X=4.26
+ $Y=2.12 $X2=5.05 $Y2=2.265
r256 1 71 182 $w=1.7e-07 $l=6.69309e-07 $layer=licon1_NDIFF $count=1 $X=4.52
+ $Y=0.525 $X2=4.93 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_2%A_1692_424# 1 2 3 4 15 19 24 29 30 36 37 38 40
+ 42 44 45 47
c121 38 0 5.30342e-20 $X=11.24 $Y=2.075
r122 50 52 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=10.855 $Y=1.635
+ $X2=10.87 $Y2=1.635
r123 47 49 16.8178 $w=4.28e-07 $l=5.9e-07 $layer=LI1_cond $X=11.11 $Y=0.715
+ $X2=11.7 $Y2=0.715
r124 44 45 6.71605 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=9.07 $Y=2.245
+ $X2=9.07 $Y2=2.13
r125 42 45 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=8.99 $Y=1.055
+ $X2=8.99 $Y2=2.13
r126 38 40 24.2013 $w=2.48e-07 $l=5.25e-07 $layer=LI1_cond $X=11.24 $Y=2.075
+ $X2=11.765 $Y2=2.075
r127 37 52 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=11.075 $Y=1.635
+ $X2=10.87 $Y2=1.635
r128 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.075
+ $Y=1.635 $X2=11.075 $Y2=1.635
r129 34 38 6.8199 $w=2.5e-07 $l=1.82071e-07 $layer=LI1_cond $X=11.11 $Y=1.95
+ $X2=11.24 $Y2=2.075
r130 34 36 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=11.11 $Y=1.95
+ $X2=11.11 $Y2=1.635
r131 33 47 3.65327 $w=2.6e-07 $l=3.4e-07 $layer=LI1_cond $X=11.11 $Y=1.055
+ $X2=11.11 $Y2=0.715
r132 33 36 25.7083 $w=2.58e-07 $l=5.8e-07 $layer=LI1_cond $X=11.11 $Y=1.055
+ $X2=11.11 $Y2=1.635
r133 32 47 7.41121 $w=4.28e-07 $l=2.6e-07 $layer=LI1_cond $X=10.85 $Y=0.715
+ $X2=11.11 $Y2=0.715
r134 31 32 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=10.85 $Y=0.425
+ $X2=10.85 $Y2=0.675
r135 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.765 $Y=0.34
+ $X2=10.85 $Y2=0.425
r136 29 30 110.257 $w=1.68e-07 $l=1.69e-06 $layer=LI1_cond $X=10.765 $Y=0.34
+ $X2=9.075 $Y2=0.34
r137 22 42 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.91 $Y=0.89
+ $X2=8.91 $Y2=1.055
r138 22 24 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=8.91 $Y=0.89
+ $X2=8.91 $Y2=0.54
r139 21 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.91 $Y=0.425
+ $X2=9.075 $Y2=0.34
r140 21 24 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=8.91 $Y=0.425
+ $X2=8.91 $Y2=0.54
r141 17 52 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.87 $Y=1.8
+ $X2=10.87 $Y2=1.635
r142 17 19 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=10.87 $Y=1.8
+ $X2=10.87 $Y2=2.46
r143 13 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.855 $Y=1.47
+ $X2=10.855 $Y2=1.635
r144 13 15 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=10.855 $Y=1.47
+ $X2=10.855 $Y2=0.715
r145 4 40 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=11.63
+ $Y=1.96 $X2=11.765 $Y2=2.115
r146 3 44 300 $w=1.7e-07 $l=6.69589e-07 $layer=licon1_PDIFF $count=2 $X=8.46
+ $Y=2.12 $X2=9.07 $Y2=2.245
r147 2 49 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.56
+ $Y=0.395 $X2=11.7 $Y2=0.54
r148 1 24 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=8.7
+ $Y=0.395 $X2=8.91 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_2%CI 3 8 10 11 12 15 17
c46 15 0 1.08693e-19 $X=11.615 $Y=1.615
c47 10 0 2.46841e-20 $X=11.505 $Y=1.11
c48 8 0 1.35554e-19 $X=11.54 $Y=2.46
r49 15 18 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.615 $Y=1.615
+ $X2=11.615 $Y2=1.78
r50 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.615 $Y=1.615
+ $X2=11.615 $Y2=1.45
r51 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.615
+ $Y=1.615 $X2=11.615 $Y2=1.615
r52 12 16 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=11.76 $Y=1.615
+ $X2=11.615 $Y2=1.615
r53 11 17 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=11.525 $Y=1.26
+ $X2=11.525 $Y2=1.45
r54 10 11 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=11.505 $Y=1.11
+ $X2=11.505 $Y2=1.26
r55 8 18 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=11.54 $Y=2.46
+ $X2=11.54 $Y2=1.78
r56 3 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=11.485 $Y=0.715
+ $X2=11.485 $Y2=1.11
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_2%A_1454_424# 1 2 9 11 13 14 16 19 21 25 27 28
+ 34 35 41 42
c132 42 0 1.08693e-19 $X=12.24 $Y=0.925
c133 41 0 7.1893e-20 $X=12.24 $Y=0.925
c134 34 0 1.39782e-19 $X=12.095 $Y=0.925
c135 27 0 1.77494e-19 $X=8.225 $Y=1.04
c136 25 0 3.57146e-20 $X=12.98 $Y=1.385
c137 19 0 2.31759e-20 $X=12.98 $Y=2.4
c138 14 0 2.25411e-19 $X=12.965 $Y=1.22
r139 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.25
+ $Y=1.385 $X2=12.25 $Y2=1.385
r140 42 46 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=12.25 $Y=0.925
+ $X2=12.25 $Y2=1.385
r141 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0.925
+ $X2=12.24 $Y2=0.925
r142 38 53 10.6717 $w=4.63e-07 $l=4.05e-07 $layer=LI1_cond $X=8.285 $Y=0.925
+ $X2=8.285 $Y2=0.52
r143 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0.925
+ $X2=8.4 $Y2=0.925
r144 35 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.545 $Y=0.925
+ $X2=8.4 $Y2=0.925
r145 34 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.095 $Y=0.925
+ $X2=12.24 $Y2=0.925
r146 34 35 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=12.095 $Y=0.925
+ $X2=8.545 $Y2=0.925
r147 28 30 1.58159 $w=6.03e-07 $l=8e-08 $layer=LI1_cond $X=8.225 $Y=2.432
+ $X2=8.145 $Y2=2.432
r148 27 38 8.16564 $w=4.63e-07 $l=1.41863e-07 $layer=LI1_cond $X=8.225 $Y=1.04
+ $X2=8.285 $Y2=0.925
r149 27 28 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=8.225 $Y=1.04
+ $X2=8.225 $Y2=2.13
r150 24 25 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=12.965 $Y=1.385
+ $X2=12.98 $Y2=1.385
r151 23 24 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=12.535 $Y=1.385
+ $X2=12.965 $Y2=1.385
r152 22 23 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=12.53 $Y=1.385
+ $X2=12.535 $Y2=1.385
r153 21 45 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=12.44 $Y=1.385
+ $X2=12.25 $Y2=1.385
r154 21 22 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=12.44 $Y=1.385
+ $X2=12.53 $Y2=1.385
r155 17 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=12.98 $Y=1.55
+ $X2=12.98 $Y2=1.385
r156 17 19 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=12.98 $Y=1.55
+ $X2=12.98 $Y2=2.4
r157 14 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.965 $Y=1.22
+ $X2=12.965 $Y2=1.385
r158 14 16 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=12.965 $Y=1.22
+ $X2=12.965 $Y2=0.74
r159 11 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.535 $Y=1.22
+ $X2=12.535 $Y2=1.385
r160 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=12.535 $Y=1.22
+ $X2=12.535 $Y2=0.74
r161 7 22 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=12.53 $Y=1.55
+ $X2=12.53 $Y2=1.385
r162 7 9 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=12.53 $Y=1.55
+ $X2=12.53 $Y2=2.4
r163 2 30 150 $w=1.7e-07 $l=9.35414e-07 $layer=licon1_PDIFF $count=4 $X=7.27
+ $Y=2.12 $X2=8.145 $Y2=2.245
r164 1 53 91 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=2 $X=7.675
+ $Y=0.395 $X2=8.18 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_2%A_1898_424# 1 2 9 13 17 21 26 28 29 31 34 36
+ 39 40 44 51 59
c121 59 0 7.31945e-20 $X=13.905 $Y=1.465
c122 39 0 1.00227e-19 $X=9.91 $Y=2.1
r123 58 59 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=13.89 $Y=1.465
+ $X2=13.905 $Y2=1.465
r124 57 58 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=13.465 $Y=1.465
+ $X2=13.89 $Y2=1.465
r125 52 57 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=13.445 $Y=1.465
+ $X2=13.465 $Y2=1.465
r126 52 54 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=13.445 $Y=1.465
+ $X2=13.43 $Y2=1.465
r127 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.445
+ $Y=1.465 $X2=13.445 $Y2=1.465
r128 48 51 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=13.315 $Y=1.465
+ $X2=13.445 $Y2=1.465
r129 44 46 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=11.885 $Y=2.455
+ $X2=11.885 $Y2=2.685
r130 40 42 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=9.91 $Y=2.685
+ $X2=9.91 $Y2=2.815
r131 38 39 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=9.83 $Y=1.185
+ $X2=9.83 $Y2=2.1
r132 36 38 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.75 $Y=1.02
+ $X2=9.75 $Y2=1.185
r133 33 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.315 $Y=1.63
+ $X2=13.315 $Y2=1.465
r134 33 34 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=13.315 $Y=1.63
+ $X2=13.315 $Y2=2.37
r135 32 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.97 $Y=2.455
+ $X2=11.885 $Y2=2.455
r136 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.23 $Y=2.455
+ $X2=13.315 $Y2=2.37
r137 31 32 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=13.23 $Y=2.455
+ $X2=11.97 $Y2=2.455
r138 30 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.075 $Y=2.685
+ $X2=9.91 $Y2=2.685
r139 29 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.8 $Y=2.685
+ $X2=11.885 $Y2=2.685
r140 29 30 112.54 $w=1.68e-07 $l=1.725e-06 $layer=LI1_cond $X=11.8 $Y=2.685
+ $X2=10.075 $Y2=2.685
r141 28 39 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.91 $Y=2.265
+ $X2=9.91 $Y2=2.1
r142 26 40 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=9.91 $Y=2.6
+ $X2=9.91 $Y2=2.685
r143 26 28 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.91 $Y=2.6
+ $X2=9.91 $Y2=2.265
r144 19 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.905 $Y=1.3
+ $X2=13.905 $Y2=1.465
r145 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.905 $Y=1.3
+ $X2=13.905 $Y2=0.74
r146 15 58 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=13.89 $Y=1.63
+ $X2=13.89 $Y2=1.465
r147 15 17 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=13.89 $Y=1.63
+ $X2=13.89 $Y2=2.4
r148 11 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.465 $Y=1.3
+ $X2=13.465 $Y2=1.465
r149 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.465 $Y=1.3
+ $X2=13.465 $Y2=0.74
r150 7 54 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=13.43 $Y=1.63
+ $X2=13.43 $Y2=1.465
r151 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=13.43 $Y=1.63
+ $X2=13.43 $Y2=2.4
r152 2 42 600 $w=1.7e-07 $l=8.80298e-07 $layer=licon1_PDIFF $count=1 $X=9.49
+ $Y=2.12 $X2=9.91 $Y2=2.815
r153 2 28 600 $w=1.7e-07 $l=4.87134e-07 $layer=licon1_PDIFF $count=1 $X=9.49
+ $Y=2.12 $X2=9.91 $Y2=2.265
r154 1 36 182 $w=1.7e-07 $l=7.26722e-07 $layer=licon1_NDIFF $count=1 $X=9.53
+ $Y=0.395 $X2=9.75 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_2%VPWR 1 2 3 4 5 6 7 22 24 28 34 38 42 44 46 50
+ 52 57 65 73 78 83 92 95 98 105 108 112
c130 34 0 2.96008e-20 $X=6.43 $Y=2.745
r131 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r132 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r133 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r134 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r135 98 101 9.24987 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=11.205 $Y=3.025
+ $X2=11.205 $Y2=3.33
r136 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r137 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r138 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r139 87 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.16 $Y2=3.33
r140 87 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=13.2 $Y2=3.33
r141 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r142 84 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.37 $Y=3.33
+ $X2=13.205 $Y2=3.33
r143 84 86 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=13.37 $Y=3.33
+ $X2=13.68 $Y2=3.33
r144 83 111 4.02656 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=14.045 $Y=3.33
+ $X2=14.222 $Y2=3.33
r145 83 86 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=14.045 $Y=3.33
+ $X2=13.68 $Y2=3.33
r146 82 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r147 82 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=12.24 $Y2=3.33
r148 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r149 79 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.47 $Y=3.33
+ $X2=12.305 $Y2=3.33
r150 79 81 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=12.47 $Y=3.33
+ $X2=12.72 $Y2=3.33
r151 78 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.04 $Y=3.33
+ $X2=13.205 $Y2=3.33
r152 78 81 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=13.04 $Y=3.33
+ $X2=12.72 $Y2=3.33
r153 77 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r154 77 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=11.28 $Y2=3.33
r155 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r156 74 101 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.395 $Y=3.33
+ $X2=11.205 $Y2=3.33
r157 74 76 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=11.395 $Y=3.33
+ $X2=11.76 $Y2=3.33
r158 73 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.14 $Y=3.33
+ $X2=12.305 $Y2=3.33
r159 73 76 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=12.14 $Y=3.33
+ $X2=11.76 $Y2=3.33
r160 72 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r161 71 72 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r162 69 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r163 68 71 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=10.8 $Y2=3.33
r164 68 69 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r165 66 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.595 $Y=3.33
+ $X2=6.43 $Y2=3.33
r166 66 68 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.595 $Y=3.33
+ $X2=6.96 $Y2=3.33
r167 65 101 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.015 $Y=3.33
+ $X2=11.205 $Y2=3.33
r168 65 71 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=11.015 $Y=3.33
+ $X2=10.8 $Y2=3.33
r169 64 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r170 63 64 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6 $Y=3.33
+ $X2=6 $Y2=3.33
r171 61 64 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=2.16 $Y=3.33 $X2=6
+ $Y2=3.33
r172 61 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r173 60 63 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=6
+ $Y2=3.33
r174 60 61 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r175 58 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.87 $Y=3.33
+ $X2=1.705 $Y2=3.33
r176 58 60 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.87 $Y=3.33
+ $X2=2.16 $Y2=3.33
r177 57 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.265 $Y=3.33
+ $X2=6.43 $Y2=3.33
r178 57 63 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.265 $Y=3.33
+ $X2=6 $Y2=3.33
r179 56 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r180 56 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r181 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r182 53 89 4.0754 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.36 $Y=3.33 $X2=0.18
+ $Y2=3.33
r183 53 55 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=0.36 $Y=3.33
+ $X2=1.2 $Y2=3.33
r184 52 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=3.33
+ $X2=1.705 $Y2=3.33
r185 52 55 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.54 $Y=3.33
+ $X2=1.2 $Y2=3.33
r186 50 72 1.00344 $w=4.9e-07 $l=3.6e-06 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=10.8 $Y2=3.33
r187 50 69 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=6.96 $Y2=3.33
r188 46 49 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=14.17 $Y=1.985
+ $X2=14.17 $Y2=2.815
r189 44 111 3.1166 $w=2.5e-07 $l=1.07912e-07 $layer=LI1_cond $X=14.17 $Y=3.245
+ $X2=14.222 $Y2=3.33
r190 44 49 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=14.17 $Y=3.245
+ $X2=14.17 $Y2=2.815
r191 40 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.205 $Y=3.245
+ $X2=13.205 $Y2=3.33
r192 40 42 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=13.205 $Y=3.245
+ $X2=13.205 $Y2=2.805
r193 36 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.305 $Y=3.245
+ $X2=12.305 $Y2=3.33
r194 36 38 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=12.305 $Y=3.245
+ $X2=12.305 $Y2=2.805
r195 32 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.43 $Y=3.245
+ $X2=6.43 $Y2=3.33
r196 32 34 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=6.43 $Y=3.245
+ $X2=6.43 $Y2=2.745
r197 28 31 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=1.705 $Y=2.115
+ $X2=1.705 $Y2=2.815
r198 26 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=3.245
+ $X2=1.705 $Y2=3.33
r199 26 31 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.705 $Y=3.245
+ $X2=1.705 $Y2=2.815
r200 22 89 3.10183 $w=2.55e-07 $l=1.07912e-07 $layer=LI1_cond $X=0.232 $Y=3.245
+ $X2=0.18 $Y2=3.33
r201 22 24 41.5783 $w=2.53e-07 $l=9.2e-07 $layer=LI1_cond $X=0.232 $Y=3.245
+ $X2=0.232 $Y2=2.325
r202 7 49 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=13.98
+ $Y=1.84 $X2=14.13 $Y2=2.815
r203 7 46 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=13.98
+ $Y=1.84 $X2=14.13 $Y2=1.985
r204 6 42 600 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=13.07
+ $Y=1.84 $X2=13.205 $Y2=2.805
r205 5 38 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=12.17
+ $Y=2.65 $X2=12.305 $Y2=2.805
r206 4 98 600 $w=1.7e-07 $l=1.18116e-06 $layer=licon1_PDIFF $count=1 $X=10.96
+ $Y=1.96 $X2=11.205 $Y2=3.025
r207 3 34 600 $w=1.7e-07 $l=9.70155e-07 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=1.84 $X2=6.43 $Y2=2.745
r208 2 31 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=1.96 $X2=1.705 $Y2=2.815
r209 2 28 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=1.96 $X2=1.705 $Y2=2.115
r210 1 24 300 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.325
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_2%A_117_368# 1 2 3 4 14 17 21 23 27 28 32 34 35
+ 41 45
c105 35 0 1.93813e-19 $X=0.385 $Y=1.295
c106 34 0 1.29241e-19 $X=3.935 $Y=1.295
r107 42 48 10.7189 $w=3.13e-07 $l=2.75e-07 $layer=LI1_cond $X=4.07 $Y=1.295
+ $X2=4.07 $Y2=1.02
r108 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=1.295
+ $X2=4.08 $Y2=1.295
r109 38 45 10.6381 $w=2.89e-07 $l=2.52e-07 $layer=LI1_cond $X=0.24 $Y=1.215
+ $X2=0.492 $Y2=1.215
r110 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.295
r111 35 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.385 $Y=1.295
+ $X2=0.24 $Y2=1.295
r112 34 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.935 $Y=1.295
+ $X2=4.08 $Y2=1.295
r113 34 35 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=3.935 $Y=1.295
+ $X2=0.385 $Y2=1.295
r114 27 42 7.01145 $w=3.13e-07 $l=1.35647e-07 $layer=LI1_cond $X=4.025 $Y=1.41
+ $X2=4.07 $Y2=1.295
r115 27 28 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=4.025 $Y=1.41
+ $X2=4.025 $Y2=2.13
r116 23 28 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.94 $Y=2.255
+ $X2=4.025 $Y2=2.13
r117 23 25 3.45733 $w=2.48e-07 $l=7.5e-08 $layer=LI1_cond $X=3.94 $Y=2.255
+ $X2=3.865 $Y2=2.255
r118 19 45 14.4796 $w=2.89e-07 $l=4.52895e-07 $layer=LI1_cond $X=0.835 $Y=0.96
+ $X2=0.492 $Y2=1.215
r119 19 21 19.7245 $w=2.58e-07 $l=4.45e-07 $layer=LI1_cond $X=0.835 $Y=0.96
+ $X2=0.835 $Y2=0.515
r120 17 32 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=0.72 $Y=2.815
+ $X2=0.72 $Y2=1.99
r121 14 32 14.8749 $w=1.68e-07 $l=2.28e-07 $layer=LI1_cond $X=0.492 $Y=1.905
+ $X2=0.72 $Y2=1.905
r122 13 45 0.205252 $w=3.15e-07 $l=2.55e-07 $layer=LI1_cond $X=0.492 $Y=1.47
+ $X2=0.492 $Y2=1.215
r123 13 14 12.8049 $w=3.13e-07 $l=3.5e-07 $layer=LI1_cond $X=0.492 $Y=1.47
+ $X2=0.492 $Y2=1.82
r124 4 25 600 $w=1.7e-07 $l=2.89569e-07 $layer=licon1_PDIFF $count=1 $X=3.65
+ $Y=2.12 $X2=3.865 $Y2=2.295
r125 3 32 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.72 $Y2=1.985
r126 3 17 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.72 $Y2=2.815
r127 2 48 182 $w=1.7e-07 $l=7.58123e-07 $layer=licon1_NDIFF $count=1 $X=3.52
+ $Y=0.525 $X2=4.07 $Y2=1.02
r128 1 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.66
+ $Y=0.37 $X2=0.8 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_2%A_416_392# 1 2 3 4 13 16 22 23 24 25 26 29 31
+ 33 34
c87 34 0 2.83882e-20 $X=5.77 $Y=0.34
c88 26 0 2.24154e-20 $X=2.555 $Y=0.34
c89 24 0 8.42529e-20 $X=2.385 $Y=2.975
c90 2 0 1.42825e-19 $X=5.365 $Y=0.525
r91 34 37 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=5.77 $Y=0.34
+ $X2=5.77 $Y2=0.665
r92 32 33 9.02376 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=2.385 $Y=1.015
+ $X2=2.385 $Y2=1.185
r93 31 33 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.3 $Y=2.015 $X2=2.3
+ $Y2=1.185
r94 27 29 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=5.89 $Y=2.89
+ $X2=5.89 $Y2=2.605
r95 25 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.605 $Y=0.34
+ $X2=5.77 $Y2=0.34
r96 25 26 198.984 $w=1.68e-07 $l=3.05e-06 $layer=LI1_cond $X=5.605 $Y=0.34
+ $X2=2.555 $Y2=0.34
r97 23 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.725 $Y=2.975
+ $X2=5.89 $Y2=2.89
r98 23 24 217.904 $w=1.68e-07 $l=3.34e-06 $layer=LI1_cond $X=5.725 $Y=2.975
+ $X2=2.385 $Y2=2.975
r99 22 32 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=2.43 $Y=0.67
+ $X2=2.43 $Y2=1.015
r100 19 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.43 $Y=0.425
+ $X2=2.555 $Y2=0.34
r101 19 22 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=2.43 $Y=0.425
+ $X2=2.43 $Y2=0.67
r102 14 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.22 $Y=2.89
+ $X2=2.385 $Y2=2.975
r103 14 16 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=2.22 $Y=2.89
+ $X2=2.22 $Y2=2.245
r104 13 31 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=2.18
+ $X2=2.22 $Y2=2.015
r105 13 16 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=2.22 $Y=2.18
+ $X2=2.22 $Y2=2.245
r106 4 29 600 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=1 $X=5.755
+ $Y=2.12 $X2=5.89 $Y2=2.605
r107 3 16 300 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=2 $X=2.08
+ $Y=1.96 $X2=2.22 $Y2=2.245
r108 2 37 182 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_NDIFF $count=1 $X=5.365
+ $Y=0.525 $X2=5.77 $Y2=0.665
r109 1 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.33
+ $Y=0.525 $X2=2.47 $Y2=0.67
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_2%A_2055_424# 1 2 7 13 16 19
c39 19 0 2.46841e-20 $X=10.725 $Y=1.1
c40 16 0 1.35554e-19 $X=10.725 $Y=2.13
r41 17 19 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=10.51 $Y=1.1
+ $X2=10.725 $Y2=1.1
r42 15 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.725 $Y=1.185
+ $X2=10.725 $Y2=1.1
r43 15 16 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=10.725 $Y=1.185
+ $X2=10.725 $Y2=2.13
r44 11 17 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.51 $Y=1.015
+ $X2=10.51 $Y2=1.1
r45 11 13 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=10.51 $Y=1.015
+ $X2=10.51 $Y2=0.825
r46 7 16 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=10.64 $Y=2.28
+ $X2=10.725 $Y2=2.13
r47 7 9 5.57014 $w=2.98e-07 $l=1.45e-07 $layer=LI1_cond $X=10.64 $Y=2.28
+ $X2=10.495 $Y2=2.28
r48 2 9 600 $w=1.7e-07 $l=2.94788e-07 $layer=licon1_PDIFF $count=1 $X=10.275
+ $Y=2.12 $X2=10.495 $Y2=2.295
r49 1 13 182 $w=1.7e-07 $l=4.994e-07 $layer=licon1_NDIFF $count=1 $X=10.36
+ $Y=0.395 $X2=10.51 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_2%COUT 1 2 9 11 12 25
c22 11 0 7.31945e-20 $X=12.635 $Y=1.58
r23 16 25 1.78887 $w=3.33e-07 $l=5.2e-08 $layer=LI1_cond $X=12.752 $Y=1.717
+ $X2=12.752 $Y2=1.665
r24 11 25 0.584822 $w=3.33e-07 $l=1.7e-08 $layer=LI1_cond $X=12.752 $Y=1.648
+ $X2=12.752 $Y2=1.665
r25 11 23 4.13832 $w=3.33e-07 $l=9.8e-08 $layer=LI1_cond $X=12.752 $Y=1.648
+ $X2=12.752 $Y2=1.55
r26 11 12 9.52916 $w=3.33e-07 $l=2.77e-07 $layer=LI1_cond $X=12.752 $Y=1.733
+ $X2=12.752 $Y2=2.01
r27 11 16 0.550421 $w=3.33e-07 $l=1.6e-08 $layer=LI1_cond $X=12.752 $Y=1.733
+ $X2=12.752 $Y2=1.717
r28 9 23 47.7111 $w=2.48e-07 $l=1.035e-06 $layer=LI1_cond $X=12.71 $Y=0.515
+ $X2=12.71 $Y2=1.55
r29 2 12 600 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=12.62
+ $Y=1.84 $X2=12.755 $Y2=2.01
r30 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.61
+ $Y=0.37 $X2=12.75 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_2%SUM 1 2 9 11 13 19 20
c35 20 0 1.21085e-19 $X=14.16 $Y=1.295
c36 19 0 2.31759e-20 $X=13.722 $Y=1.82
c37 9 0 1.4004e-19 $X=13.685 $Y=0.52
r38 26 27 2.09656 $w=6.11e-07 $l=2.33675e-07 $layer=LI1_cond $X=13.685 $Y=0.965
+ $X2=13.79 $Y2=1.152
r39 20 27 7.38789 $w=6.11e-07 $l=3.7e-07 $layer=LI1_cond $X=14.16 $Y=1.152
+ $X2=13.79 $Y2=1.152
r40 17 27 8.43407 $w=1.7e-07 $l=3.53e-07 $layer=LI1_cond $X=13.79 $Y=1.505
+ $X2=13.79 $Y2=1.152
r41 17 19 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=13.79 $Y=1.505
+ $X2=13.79 $Y2=1.82
r42 13 15 31.3616 $w=3.03e-07 $l=8.3e-07 $layer=LI1_cond $X=13.722 $Y=1.985
+ $X2=13.722 $Y2=2.815
r43 11 19 7.98337 $w=3.03e-07 $l=1.52e-07 $layer=LI1_cond $X=13.722 $Y=1.972
+ $X2=13.722 $Y2=1.82
r44 11 13 0.491205 $w=3.03e-07 $l=1.3e-08 $layer=LI1_cond $X=13.722 $Y=1.972
+ $X2=13.722 $Y2=1.985
r45 7 26 0.698854 $w=6.11e-07 $l=1.81659e-07 $layer=LI1_cond $X=13.65 $Y=0.8
+ $X2=13.685 $Y2=0.965
r46 7 9 11.9513 $w=2.68e-07 $l=2.8e-07 $layer=LI1_cond $X=13.65 $Y=0.8 $X2=13.65
+ $Y2=0.52
r47 2 15 400 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=1 $X=13.52
+ $Y=1.84 $X2=13.66 $Y2=2.815
r48 2 13 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.52
+ $Y=1.84 $X2=13.66 $Y2=1.985
r49 1 26 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=13.54
+ $Y=0.37 $X2=13.685 $Y2=0.965
r50 1 9 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=13.54
+ $Y=0.37 $X2=13.685 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_MS__FAH_2%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44 46 48
+ 51 52 54 55 56 65 79 83 88 97 100 103 107
r136 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r137 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r138 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r139 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r140 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r141 92 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=14.16 $Y2=0
r142 92 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r143 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r144 89 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.345 $Y=0
+ $X2=13.18 $Y2=0
r145 89 91 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=13.345 $Y=0
+ $X2=13.68 $Y2=0
r146 88 106 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=13.955 $Y=0
+ $X2=14.177 $Y2=0
r147 88 91 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=13.955 $Y=0
+ $X2=13.68 $Y2=0
r148 87 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r149 87 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r150 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r151 84 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.405 $Y=0
+ $X2=12.24 $Y2=0
r152 84 86 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.405 $Y=0
+ $X2=12.72 $Y2=0
r153 83 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.015 $Y=0
+ $X2=13.18 $Y2=0
r154 83 86 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.015 $Y=0
+ $X2=12.72 $Y2=0
r155 82 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r156 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r157 79 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.075 $Y=0
+ $X2=12.24 $Y2=0
r158 79 81 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.075 $Y=0
+ $X2=11.76 $Y2=0
r159 78 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.76 $Y2=0
r160 77 78 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r161 75 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r162 74 77 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=6.96 $Y=0 $X2=10.8
+ $Y2=0
r163 74 75 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r164 72 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.665 $Y=0 $X2=6.5
+ $Y2=0
r165 72 74 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.665 $Y=0 $X2=6.96
+ $Y2=0
r166 71 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r167 70 71 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6 $Y=0 $X2=6
+ $Y2=0
r168 68 71 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=6
+ $Y2=0
r169 67 70 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=6
+ $Y2=0
r170 67 68 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r171 65 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.335 $Y=0 $X2=6.5
+ $Y2=0
r172 65 70 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.335 $Y=0 $X2=6
+ $Y2=0
r173 64 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r174 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r175 61 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r176 61 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r177 60 63 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r178 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r179 58 94 4.9356 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.267
+ $Y2=0
r180 58 60 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.535 $Y=0
+ $X2=0.72 $Y2=0
r181 56 78 1.00344 $w=4.9e-07 $l=3.6e-06 $layer=MET1_cond $X=7.2 $Y=0 $X2=10.8
+ $Y2=0
r182 56 75 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=0 $X2=6.96
+ $Y2=0
r183 54 77 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=11.105 $Y=0
+ $X2=10.8 $Y2=0
r184 54 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.105 $Y=0
+ $X2=11.23 $Y2=0
r185 53 81 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=11.355 $Y=0
+ $X2=11.76 $Y2=0
r186 53 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.355 $Y=0
+ $X2=11.23 $Y2=0
r187 51 63 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=1.68 $Y2=0
r188 51 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2
+ $Y2=0
r189 50 67 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.125 $Y=0 $X2=2.16
+ $Y2=0
r190 50 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=2
+ $Y2=0
r191 46 106 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=14.12 $Y=0.085
+ $X2=14.177 $Y2=0
r192 46 48 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=14.12 $Y=0.085
+ $X2=14.12 $Y2=0.53
r193 42 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.18 $Y=0.085
+ $X2=13.18 $Y2=0
r194 42 44 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.18 $Y=0.085
+ $X2=13.18 $Y2=0.515
r195 38 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.24 $Y=0.085
+ $X2=12.24 $Y2=0
r196 38 40 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=12.24 $Y=0.085
+ $X2=12.24 $Y2=0.475
r197 34 55 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.23 $Y=0.085
+ $X2=11.23 $Y2=0
r198 34 36 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=11.23 $Y=0.085
+ $X2=11.23 $Y2=0.34
r199 30 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.5 $Y=0.085 $X2=6.5
+ $Y2=0
r200 30 32 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.5 $Y=0.085
+ $X2=6.5 $Y2=0.515
r201 26 52 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2 $Y=0.085 $X2=2
+ $Y2=0
r202 26 28 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=2 $Y=0.085 $X2=2
+ $Y2=0.675
r203 22 94 3.13079 $w=3.65e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.352 $Y=0.085
+ $X2=0.267 $Y2=0
r204 22 24 18.1549 $w=3.63e-07 $l=5.75e-07 $layer=LI1_cond $X=0.352 $Y=0.085
+ $X2=0.352 $Y2=0.66
r205 7 48 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=13.98
+ $Y=0.37 $X2=14.12 $Y2=0.53
r206 6 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.04
+ $Y=0.37 $X2=13.18 $Y2=0.515
r207 5 40 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=12.105
+ $Y=0.33 $X2=12.24 $Y2=0.475
r208 4 36 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=10.93
+ $Y=0.395 $X2=11.19 $Y2=0.34
r209 3 32 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=6.355
+ $Y=0.37 $X2=6.5 $Y2=0.515
r210 2 28 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=1.9
+ $Y=0.525 $X2=2.04 $Y2=0.675
r211 1 24 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=0.21
+ $Y=0.37 $X2=0.37 $Y2=0.66
.ends


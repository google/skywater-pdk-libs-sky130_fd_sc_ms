* File: sky130_fd_sc_ms__sdlclkp_2.pxi.spice
* Created: Wed Sep  2 12:32:09 2020
* 
x_PM_SKY130_FD_SC_MS__SDLCLKP_2%SCE N_SCE_c_166_n N_SCE_M1022_g N_SCE_M1015_g
+ N_SCE_c_172_n SCE N_SCE_c_168_n N_SCE_c_169_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_2%SCE
x_PM_SKY130_FD_SC_MS__SDLCLKP_2%GATE N_GATE_M1008_g N_GATE_M1014_g GATE
+ N_GATE_c_199_n N_GATE_c_200_n PM_SKY130_FD_SC_MS__SDLCLKP_2%GATE
x_PM_SKY130_FD_SC_MS__SDLCLKP_2%A_318_74# N_A_318_74#_M1006_d
+ N_A_318_74#_M1012_d N_A_318_74#_M1005_g N_A_318_74#_M1018_g
+ N_A_318_74#_c_240_n N_A_318_74#_c_241_n N_A_318_74#_c_242_n
+ N_A_318_74#_c_243_n N_A_318_74#_c_244_n N_A_318_74#_c_245_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_2%A_318_74#
x_PM_SKY130_FD_SC_MS__SDLCLKP_2%A_288_48# N_A_288_48#_M1002_s
+ N_A_288_48#_M1010_s N_A_288_48#_c_319_n N_A_288_48#_M1006_g
+ N_A_288_48#_c_320_n N_A_288_48#_c_321_n N_A_288_48#_M1012_g
+ N_A_288_48#_c_339_n N_A_288_48#_c_340_n N_A_288_48#_c_323_n
+ N_A_288_48#_c_324_n N_A_288_48#_c_325_n N_A_288_48#_M1023_g
+ N_A_288_48#_M1013_g N_A_288_48#_c_326_n N_A_288_48#_c_327_n
+ N_A_288_48#_c_328_n N_A_288_48#_c_329_n N_A_288_48#_c_330_n
+ N_A_288_48#_c_331_n N_A_288_48#_c_380_p N_A_288_48#_c_332_n
+ N_A_288_48#_c_333_n N_A_288_48#_c_334_n N_A_288_48#_c_335_n
+ N_A_288_48#_c_336_n N_A_288_48#_c_342_n N_A_288_48#_c_337_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_2%A_288_48#
x_PM_SKY130_FD_SC_MS__SDLCLKP_2%A_706_317# N_A_706_317#_M1004_d
+ N_A_706_317#_M1000_d N_A_706_317#_M1019_g N_A_706_317#_M1007_g
+ N_A_706_317#_M1011_g N_A_706_317#_M1020_g N_A_706_317#_c_488_n
+ N_A_706_317#_c_489_n N_A_706_317#_c_490_n N_A_706_317#_c_477_n
+ N_A_706_317#_c_478_n N_A_706_317#_c_492_n N_A_706_317#_c_479_n
+ N_A_706_317#_c_480_n N_A_706_317#_c_481_n N_A_706_317#_c_482_n
+ N_A_706_317#_c_495_n N_A_706_317#_c_496_n N_A_706_317#_c_483_n
+ N_A_706_317#_c_484_n N_A_706_317#_c_485_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_2%A_706_317#
x_PM_SKY130_FD_SC_MS__SDLCLKP_2%A_580_74# N_A_580_74#_M1023_d
+ N_A_580_74#_M1005_d N_A_580_74#_M1000_g N_A_580_74#_M1004_g
+ N_A_580_74#_c_619_n N_A_580_74#_c_608_n N_A_580_74#_c_609_n
+ N_A_580_74#_c_615_n N_A_580_74#_c_610_n N_A_580_74#_c_631_n
+ N_A_580_74#_c_611_n N_A_580_74#_c_612_n N_A_580_74#_c_613_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_2%A_580_74#
x_PM_SKY130_FD_SC_MS__SDLCLKP_2%CLK N_CLK_M1010_g N_CLK_c_693_n N_CLK_M1002_g
+ N_CLK_M1021_g N_CLK_c_695_n N_CLK_M1016_g CLK N_CLK_c_697_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_2%CLK
x_PM_SKY130_FD_SC_MS__SDLCLKP_2%A_1198_374# N_A_1198_374#_M1011_d
+ N_A_1198_374#_M1021_d N_A_1198_374#_M1001_g N_A_1198_374#_M1009_g
+ N_A_1198_374#_M1003_g N_A_1198_374#_M1017_g N_A_1198_374#_c_758_n
+ N_A_1198_374#_c_749_n N_A_1198_374#_c_759_n N_A_1198_374#_c_760_n
+ N_A_1198_374#_c_750_n N_A_1198_374#_c_751_n N_A_1198_374#_c_752_n
+ N_A_1198_374#_c_753_n N_A_1198_374#_c_754_n N_A_1198_374#_c_755_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_2%A_1198_374#
x_PM_SKY130_FD_SC_MS__SDLCLKP_2%VPWR N_VPWR_M1022_s N_VPWR_M1012_s
+ N_VPWR_M1007_d N_VPWR_M1010_d N_VPWR_M1020_d N_VPWR_M1003_s N_VPWR_c_836_n
+ N_VPWR_c_837_n N_VPWR_c_838_n N_VPWR_c_839_n N_VPWR_c_840_n N_VPWR_c_841_n
+ N_VPWR_c_842_n N_VPWR_c_843_n N_VPWR_c_844_n N_VPWR_c_845_n VPWR
+ N_VPWR_c_846_n N_VPWR_c_847_n N_VPWR_c_848_n N_VPWR_c_849_n N_VPWR_c_850_n
+ N_VPWR_c_851_n N_VPWR_c_852_n N_VPWR_c_835_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_2%VPWR
x_PM_SKY130_FD_SC_MS__SDLCLKP_2%A_114_112# N_A_114_112#_M1015_d
+ N_A_114_112#_M1023_s N_A_114_112#_M1008_d N_A_114_112#_M1005_s
+ N_A_114_112#_c_927_n N_A_114_112#_c_942_n N_A_114_112#_c_928_n
+ N_A_114_112#_c_929_n N_A_114_112#_c_930_n N_A_114_112#_c_933_n
+ N_A_114_112#_c_931_n N_A_114_112#_c_935_n N_A_114_112#_c_936_n
+ N_A_114_112#_c_937_n N_A_114_112#_c_938_n N_A_114_112#_c_932_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_2%A_114_112#
x_PM_SKY130_FD_SC_MS__SDLCLKP_2%GCLK N_GCLK_M1009_d N_GCLK_M1001_d
+ N_GCLK_c_1025_n N_GCLK_c_1026_n GCLK GCLK GCLK GCLK N_GCLK_c_1027_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_2%GCLK
x_PM_SKY130_FD_SC_MS__SDLCLKP_2%VGND N_VGND_M1015_s N_VGND_M1014_d
+ N_VGND_M1019_d N_VGND_M1002_d N_VGND_M1009_s N_VGND_M1017_s N_VGND_c_1062_n
+ N_VGND_c_1063_n N_VGND_c_1064_n N_VGND_c_1065_n N_VGND_c_1066_n
+ N_VGND_c_1067_n N_VGND_c_1068_n N_VGND_c_1069_n N_VGND_c_1070_n
+ N_VGND_c_1071_n N_VGND_c_1072_n VGND N_VGND_c_1073_n N_VGND_c_1074_n
+ N_VGND_c_1075_n N_VGND_c_1076_n N_VGND_c_1077_n N_VGND_c_1078_n
+ PM_SKY130_FD_SC_MS__SDLCLKP_2%VGND
cc_1 VNB N_SCE_c_166_n 0.0160819f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.778
cc_2 VNB N_SCE_M1015_g 0.0259574f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_3 VNB N_SCE_c_168_n 0.0228767f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_4 VNB N_SCE_c_169_n 0.0150846f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_5 VNB N_GATE_M1014_g 0.0410235f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.29
cc_6 VNB N_GATE_c_199_n 0.00752165f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_GATE_c_200_n 0.0039698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_318_74#_M1018_g 0.0290535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_318_74#_c_240_n 0.00409123f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_10 VNB N_A_318_74#_c_241_n 0.00340601f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.29
cc_11 VNB N_A_318_74#_c_242_n 0.00392562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_318_74#_c_243_n 0.00407793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_318_74#_c_244_n 0.0039819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_318_74#_c_245_n 0.0624237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_288_48#_c_319_n 0.0222943f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.29
cc_16 VNB N_A_288_48#_c_320_n 0.0196979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_288_48#_c_321_n 0.00949141f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.96
cc_18 VNB N_A_288_48#_M1012_g 0.0197795f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_19 VNB N_A_288_48#_c_323_n 0.0286287f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.625
cc_20 VNB N_A_288_48#_c_324_n 0.0570203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_288_48#_c_325_n 0.018287f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_288_48#_c_326_n 0.0017689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_288_48#_c_327_n 0.00620923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_288_48#_c_328_n 0.0054008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_288_48#_c_329_n 4.56848e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_288_48#_c_330_n 0.0083234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_288_48#_c_331_n 0.00200416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_288_48#_c_332_n 0.0157841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_288_48#_c_333_n 0.00232637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_288_48#_c_334_n 0.00425067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_288_48#_c_335_n 0.0103992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_288_48#_c_336_n 0.001685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_288_48#_c_337_n 0.00971058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_706_317#_M1019_g 0.0516566f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_35 VNB N_A_706_317#_M1011_g 0.0244504f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.29
cc_36 VNB N_A_706_317#_M1020_g 0.00198024f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.625
cc_37 VNB N_A_706_317#_c_477_n 0.00340445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_706_317#_c_478_n 0.00882689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_706_317#_c_479_n 3.62031e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_706_317#_c_480_n 6.10912e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_706_317#_c_481_n 0.0137603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_706_317#_c_482_n 0.00147549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_706_317#_c_483_n 0.00121771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_706_317#_c_484_n 0.00835532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_706_317#_c_485_n 0.0398771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_580_74#_c_608_n 0.00278951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_580_74#_c_609_n 0.018075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_580_74#_c_610_n 0.0022609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_580_74#_c_611_n 0.00177044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_580_74#_c_612_n 0.0294365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_580_74#_c_613_n 0.019747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_CLK_M1010_g 5.51528e-19 $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.96
cc_53 VNB N_CLK_c_693_n 0.0198677f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.54
cc_54 VNB N_CLK_M1021_g 0.00279639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_CLK_c_695_n 0.0169383f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_56 VNB CLK 0.00534056f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.455
cc_57 VNB N_CLK_c_697_n 0.0485401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1198_374#_M1001_g 0.00170773f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=0.835
cc_59 VNB N_A_1198_374#_M1009_g 0.0224327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1198_374#_M1003_g 0.00231818f $X=-0.19 $Y=-0.245 $X2=0.402
+ $Y2=1.29
cc_61 VNB N_A_1198_374#_M1017_g 0.0266863f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.625
cc_62 VNB N_A_1198_374#_c_749_n 0.00882336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1198_374#_c_750_n 0.012386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1198_374#_c_751_n 0.0024413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1198_374#_c_752_n 5.02584e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1198_374#_c_753_n 0.00651904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1198_374#_c_754_n 0.00347217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1198_374#_c_755_n 0.0716999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VPWR_c_835_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_114_112#_c_927_n 0.011371f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.455
cc_71 VNB N_A_114_112#_c_928_n 0.00956352f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.29
cc_72 VNB N_A_114_112#_c_929_n 0.00325069f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.625
cc_73 VNB N_A_114_112#_c_930_n 0.0148174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_114_112#_c_931_n 0.00557558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_114_112#_c_932_n 0.00641776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_GCLK_c_1025_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_77 VNB N_GCLK_c_1026_n 0.00448002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_GCLK_c_1027_n 0.0030223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1062_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1063_n 0.0503665f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.625
cc_81 VNB N_VGND_c_1064_n 0.00858671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1065_n 0.006053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1066_n 0.0133405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1067_n 0.010359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1068_n 0.050871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1069_n 0.0621246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1070_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1071_n 0.0364191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1072_n 0.00615884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1073_n 0.0191861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1074_n 0.0291972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1075_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1076_n 0.017485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1077_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1078_n 0.469354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VPB N_SCE_c_166_n 0.00982416f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.778
cc_97 VPB N_SCE_M1022_g 0.0274725f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.54
cc_98 VPB N_SCE_c_172_n 0.0200571f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.96
cc_99 VPB N_SCE_c_169_n 0.0123922f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_100 VPB N_GATE_M1008_g 0.024602f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.96
cc_101 VPB N_GATE_c_199_n 0.0283399f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_102 VPB N_GATE_c_200_n 0.00419679f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_318_74#_M1005_g 0.0272096f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.835
cc_104 VPB N_A_318_74#_c_241_n 0.00494693f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.29
cc_105 VPB N_A_318_74#_c_243_n 0.00743775f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_318_74#_c_244_n 0.00290184f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_318_74#_c_245_n 0.0177902f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_288_48#_M1012_g 0.0428862f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_109 VPB N_A_288_48#_c_339_n 0.110986f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.455
cc_110 VPB N_A_288_48#_c_340_n 0.0140007f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.29
cc_111 VPB N_A_288_48#_M1013_g 0.0476078f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_288_48#_c_342_n 0.00707478f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_288_48#_c_337_n 0.0028341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_706_317#_M1007_g 0.0344967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_706_317#_M1020_g 0.0271145f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.625
cc_116 VPB N_A_706_317#_c_488_n 0.00518421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_706_317#_c_489_n 0.00409167f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_706_317#_c_490_n 0.0173867f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_706_317#_c_478_n 0.00382862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_706_317#_c_492_n 0.0134329f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_706_317#_c_479_n 0.00223394f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_706_317#_c_482_n 0.00836574f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_706_317#_c_495_n 0.00591409f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_706_317#_c_496_n 5.34456e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_706_317#_c_484_n 0.033672f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_580_74#_M1000_g 0.0285509f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.835
cc_127 VPB N_A_580_74#_c_615_n 0.00122269f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_580_74#_c_610_n 0.00731419f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_580_74#_c_611_n 0.00137316f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_580_74#_c_612_n 0.00657025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_CLK_M1010_g 0.0261983f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.96
cc_132 VPB N_CLK_M1021_g 0.0297633f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_1198_374#_M1001_g 0.0241244f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.835
cc_134 VPB N_A_1198_374#_M1003_g 0.0274024f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.29
cc_135 VPB N_A_1198_374#_c_758_n 0.00322246f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_1198_374#_c_759_n 0.00373308f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_1198_374#_c_760_n 0.0026267f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_1198_374#_c_752_n 0.00240894f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_836_n 0.0116777f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_837_n 0.0426189f $X=-0.19 $Y=1.66 $X2=0.385 $Y2=1.625
cc_141 VPB N_VPWR_c_838_n 0.0162732f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_839_n 0.0173157f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_840_n 0.0249044f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_841_n 0.0130501f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_842_n 0.0124065f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_843_n 0.0642794f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_844_n 0.0254743f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_845_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_846_n 0.0306291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_847_n 0.0663018f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_848_n 0.0376907f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_849_n 0.0194542f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_850_n 0.00626979f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_851_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_852_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_835_n 0.130581f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_A_114_112#_c_933_n 0.0105766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_A_114_112#_c_931_n 0.00849932f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_114_112#_c_935_n 0.0132079f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_114_112#_c_936_n 0.00684448f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_A_114_112#_c_937_n 0.00873239f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_114_112#_c_938_n 8.47548e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB GCLK 0.00441499f $X=-0.19 $Y=1.66 $X2=0.402 $Y2=1.455
cc_164 VPB GCLK 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_GCLK_c_1027_n 0.00122185f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 N_SCE_c_172_n N_GATE_M1008_g 0.0442167f $X=0.402 $Y=1.96 $X2=0 $Y2=0
cc_167 N_SCE_M1015_g N_GATE_M1014_g 0.020509f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_168 N_SCE_c_168_n N_GATE_M1014_g 0.0168557f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_169 N_SCE_c_169_n N_GATE_M1014_g 0.00149764f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_170 N_SCE_c_166_n N_GATE_c_199_n 0.0442167f $X=0.402 $Y=1.778 $X2=0 $Y2=0
cc_171 N_SCE_c_169_n N_GATE_c_199_n 0.00108715f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_172 N_SCE_c_166_n N_GATE_c_200_n 0.00240586f $X=0.402 $Y=1.778 $X2=0 $Y2=0
cc_173 N_SCE_c_169_n N_GATE_c_200_n 0.0194621f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_174 N_SCE_M1022_g N_VPWR_c_837_n 0.023455f $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_175 N_SCE_c_172_n N_VPWR_c_837_n 0.0047928f $X=0.402 $Y=1.96 $X2=0 $Y2=0
cc_176 N_SCE_c_169_n N_VPWR_c_837_n 0.0246159f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_177 N_SCE_M1022_g N_VPWR_c_846_n 0.00460063f $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_178 N_SCE_M1022_g N_VPWR_c_835_n 0.00908061f $X=0.495 $Y=2.54 $X2=0 $Y2=0
cc_179 N_SCE_M1015_g N_A_114_112#_c_927_n 0.00819024f $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_180 N_SCE_c_168_n N_A_114_112#_c_927_n 0.00147346f $X=0.385 $Y=1.455 $X2=0
+ $Y2=0
cc_181 N_SCE_c_169_n N_A_114_112#_c_927_n 0.00895228f $X=0.385 $Y=1.455 $X2=0
+ $Y2=0
cc_182 N_SCE_M1015_g N_A_114_112#_c_942_n 0.00257503f $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_183 N_SCE_M1015_g N_A_114_112#_c_929_n 0.00333944f $X=0.495 $Y=0.835 $X2=0
+ $Y2=0
cc_184 N_SCE_M1022_g N_A_114_112#_c_937_n 0.00179754f $X=0.495 $Y=2.54 $X2=0
+ $Y2=0
cc_185 N_SCE_M1015_g N_VGND_c_1063_n 0.00819878f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_186 N_SCE_c_168_n N_VGND_c_1063_n 0.00386581f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_187 N_SCE_c_169_n N_VGND_c_1063_n 0.0216167f $X=0.385 $Y=1.455 $X2=0 $Y2=0
cc_188 N_SCE_M1015_g N_VGND_c_1073_n 0.00432822f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_189 N_SCE_M1015_g N_VGND_c_1078_n 0.00487769f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_190 N_GATE_M1014_g N_A_318_74#_c_242_n 5.25064e-19 $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_191 N_GATE_M1014_g N_A_288_48#_c_319_n 0.024928f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_192 N_GATE_M1008_g N_VPWR_c_837_n 0.00322322f $X=0.885 $Y=2.54 $X2=0 $Y2=0
cc_193 N_GATE_c_200_n N_VPWR_c_837_n 8.49317e-19 $X=0.96 $Y=1.795 $X2=0 $Y2=0
cc_194 N_GATE_M1008_g N_VPWR_c_838_n 0.00343721f $X=0.885 $Y=2.54 $X2=0 $Y2=0
cc_195 N_GATE_M1008_g N_VPWR_c_846_n 0.005209f $X=0.885 $Y=2.54 $X2=0 $Y2=0
cc_196 N_GATE_M1008_g N_VPWR_c_835_n 0.00988003f $X=0.885 $Y=2.54 $X2=0 $Y2=0
cc_197 N_GATE_c_200_n N_A_114_112#_M1008_d 0.00238772f $X=0.96 $Y=1.795 $X2=0
+ $Y2=0
cc_198 N_GATE_M1014_g N_A_114_112#_c_927_n 0.0100761f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_199 N_GATE_c_199_n N_A_114_112#_c_927_n 4.05655e-19 $X=0.96 $Y=1.795 $X2=0
+ $Y2=0
cc_200 N_GATE_c_200_n N_A_114_112#_c_927_n 0.00615564f $X=0.96 $Y=1.795 $X2=0
+ $Y2=0
cc_201 N_GATE_M1014_g N_A_114_112#_c_942_n 0.00513644f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_202 N_GATE_M1014_g N_A_114_112#_c_928_n 0.00867681f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_203 N_GATE_M1014_g N_A_114_112#_c_929_n 0.00231761f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_204 N_GATE_M1014_g N_A_114_112#_c_930_n 0.00909975f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_205 N_GATE_c_199_n N_A_114_112#_c_930_n 8.19427e-19 $X=0.96 $Y=1.795 $X2=0
+ $Y2=0
cc_206 N_GATE_c_200_n N_A_114_112#_c_930_n 0.025014f $X=0.96 $Y=1.795 $X2=0
+ $Y2=0
cc_207 N_GATE_c_200_n N_A_114_112#_c_933_n 0.00194498f $X=0.96 $Y=1.795 $X2=0
+ $Y2=0
cc_208 N_GATE_M1008_g N_A_114_112#_c_931_n 0.00350508f $X=0.885 $Y=2.54 $X2=0
+ $Y2=0
cc_209 N_GATE_M1014_g N_A_114_112#_c_931_n 0.00596863f $X=0.925 $Y=0.835 $X2=0
+ $Y2=0
cc_210 N_GATE_c_199_n N_A_114_112#_c_931_n 0.00153099f $X=0.96 $Y=1.795 $X2=0
+ $Y2=0
cc_211 N_GATE_c_200_n N_A_114_112#_c_931_n 0.0426645f $X=0.96 $Y=1.795 $X2=0
+ $Y2=0
cc_212 N_GATE_M1008_g N_A_114_112#_c_937_n 0.0132669f $X=0.885 $Y=2.54 $X2=0
+ $Y2=0
cc_213 N_GATE_c_199_n N_A_114_112#_c_937_n 6.37845e-19 $X=0.96 $Y=1.795 $X2=0
+ $Y2=0
cc_214 N_GATE_c_200_n N_A_114_112#_c_937_n 0.0239778f $X=0.96 $Y=1.795 $X2=0
+ $Y2=0
cc_215 N_GATE_M1014_g N_VGND_c_1073_n 0.0034063f $X=0.925 $Y=0.835 $X2=0 $Y2=0
cc_216 N_GATE_M1014_g N_VGND_c_1078_n 0.00487769f $X=0.925 $Y=0.835 $X2=0 $Y2=0
cc_217 N_A_318_74#_c_240_n N_A_288_48#_c_319_n 0.00317258f $X=1.895 $Y=1.545
+ $X2=0 $Y2=0
cc_218 N_A_318_74#_c_242_n N_A_288_48#_c_319_n 0.00411406f $X=1.895 $Y=0.965
+ $X2=0 $Y2=0
cc_219 N_A_318_74#_c_240_n N_A_288_48#_c_320_n 0.00469377f $X=1.895 $Y=1.545
+ $X2=0 $Y2=0
cc_220 N_A_318_74#_c_242_n N_A_288_48#_c_320_n 0.00535941f $X=1.895 $Y=0.965
+ $X2=0 $Y2=0
cc_221 N_A_318_74#_c_243_n N_A_288_48#_c_320_n 2.27576e-19 $X=2.34 $Y=1.847
+ $X2=0 $Y2=0
cc_222 N_A_318_74#_c_240_n N_A_288_48#_M1012_g 0.012674f $X=1.895 $Y=1.545 $X2=0
+ $Y2=0
cc_223 N_A_318_74#_c_243_n N_A_288_48#_M1012_g 0.0308895f $X=2.34 $Y=1.847 $X2=0
+ $Y2=0
cc_224 N_A_318_74#_c_244_n N_A_288_48#_M1012_g 5.65608e-19 $X=2.855 $Y=1.55
+ $X2=0 $Y2=0
cc_225 N_A_318_74#_c_245_n N_A_288_48#_M1012_g 0.00401978f $X=2.94 $Y=1.455
+ $X2=0 $Y2=0
cc_226 N_A_318_74#_M1005_g N_A_288_48#_c_339_n 0.0123772f $X=2.94 $Y=2.315 $X2=0
+ $Y2=0
cc_227 N_A_318_74#_c_241_n N_A_288_48#_c_323_n 0.00115318f $X=2.69 $Y=1.63 $X2=0
+ $Y2=0
cc_228 N_A_318_74#_c_244_n N_A_288_48#_c_323_n 0.00135102f $X=2.855 $Y=1.55
+ $X2=0 $Y2=0
cc_229 N_A_318_74#_c_245_n N_A_288_48#_c_323_n 0.0116215f $X=2.94 $Y=1.455 $X2=0
+ $Y2=0
cc_230 N_A_318_74#_c_240_n N_A_288_48#_c_324_n 0.00644266f $X=1.895 $Y=1.545
+ $X2=0 $Y2=0
cc_231 N_A_318_74#_c_242_n N_A_288_48#_c_324_n 6.5359e-19 $X=1.895 $Y=0.965
+ $X2=0 $Y2=0
cc_232 N_A_318_74#_c_243_n N_A_288_48#_c_324_n 0.00740977f $X=2.34 $Y=1.847
+ $X2=0 $Y2=0
cc_233 N_A_318_74#_c_245_n N_A_288_48#_c_324_n 0.00214647f $X=2.94 $Y=1.455
+ $X2=0 $Y2=0
cc_234 N_A_318_74#_M1018_g N_A_288_48#_c_325_n 0.0202664f $X=3.35 $Y=0.615 $X2=0
+ $Y2=0
cc_235 N_A_318_74#_M1005_g N_A_288_48#_M1013_g 0.0172848f $X=2.94 $Y=2.315 $X2=0
+ $Y2=0
cc_236 N_A_318_74#_c_242_n N_A_288_48#_c_326_n 0.00502799f $X=1.895 $Y=0.965
+ $X2=0 $Y2=0
cc_237 N_A_318_74#_M1018_g N_A_288_48#_c_327_n 0.0119709f $X=3.35 $Y=0.615 $X2=0
+ $Y2=0
cc_238 N_A_318_74#_M1018_g N_A_288_48#_c_329_n 0.00550364f $X=3.35 $Y=0.615
+ $X2=0 $Y2=0
cc_239 N_A_318_74#_M1018_g N_A_288_48#_c_331_n 0.00115488f $X=3.35 $Y=0.615
+ $X2=0 $Y2=0
cc_240 N_A_318_74#_M1018_g N_A_288_48#_c_335_n 3.86166e-19 $X=3.35 $Y=0.615
+ $X2=0 $Y2=0
cc_241 N_A_318_74#_c_240_n N_A_288_48#_c_335_n 0.023335f $X=1.895 $Y=1.545 $X2=0
+ $Y2=0
cc_242 N_A_318_74#_c_241_n N_A_288_48#_c_335_n 0.0104963f $X=2.69 $Y=1.63 $X2=0
+ $Y2=0
cc_243 N_A_318_74#_c_242_n N_A_288_48#_c_335_n 0.00160791f $X=1.895 $Y=0.965
+ $X2=0 $Y2=0
cc_244 N_A_318_74#_c_243_n N_A_288_48#_c_335_n 0.0247748f $X=2.34 $Y=1.847 $X2=0
+ $Y2=0
cc_245 N_A_318_74#_c_244_n N_A_288_48#_c_335_n 0.00190778f $X=2.855 $Y=1.55
+ $X2=0 $Y2=0
cc_246 N_A_318_74#_c_245_n N_A_288_48#_c_335_n 9.77176e-19 $X=2.94 $Y=1.455
+ $X2=0 $Y2=0
cc_247 N_A_318_74#_M1018_g N_A_706_317#_M1019_g 0.0547363f $X=3.35 $Y=0.615
+ $X2=0 $Y2=0
cc_248 N_A_318_74#_c_245_n N_A_706_317#_M1019_g 0.00691964f $X=2.94 $Y=1.455
+ $X2=0 $Y2=0
cc_249 N_A_318_74#_M1005_g N_A_706_317#_c_484_n 0.00327975f $X=2.94 $Y=2.315
+ $X2=0 $Y2=0
cc_250 N_A_318_74#_c_245_n N_A_706_317#_c_484_n 0.00698703f $X=2.94 $Y=1.455
+ $X2=0 $Y2=0
cc_251 N_A_318_74#_M1018_g N_A_580_74#_c_619_n 0.00840926f $X=3.35 $Y=0.615
+ $X2=0 $Y2=0
cc_252 N_A_318_74#_c_244_n N_A_580_74#_c_619_n 0.00316115f $X=2.855 $Y=1.55
+ $X2=0 $Y2=0
cc_253 N_A_318_74#_c_245_n N_A_580_74#_c_619_n 0.00541836f $X=2.94 $Y=1.455
+ $X2=0 $Y2=0
cc_254 N_A_318_74#_M1018_g N_A_580_74#_c_608_n 0.00883344f $X=3.35 $Y=0.615
+ $X2=0 $Y2=0
cc_255 N_A_318_74#_c_245_n N_A_580_74#_c_608_n 0.00508821f $X=2.94 $Y=1.455
+ $X2=0 $Y2=0
cc_256 N_A_318_74#_c_245_n N_A_580_74#_c_609_n 0.00543726f $X=2.94 $Y=1.455
+ $X2=0 $Y2=0
cc_257 N_A_318_74#_M1005_g N_A_580_74#_c_615_n 0.00809131f $X=2.94 $Y=2.315
+ $X2=0 $Y2=0
cc_258 N_A_318_74#_c_244_n N_A_580_74#_c_615_n 5.57966e-19 $X=2.855 $Y=1.55
+ $X2=0 $Y2=0
cc_259 N_A_318_74#_c_245_n N_A_580_74#_c_615_n 0.00388244f $X=2.94 $Y=1.455
+ $X2=0 $Y2=0
cc_260 N_A_318_74#_M1005_g N_A_580_74#_c_610_n 0.00998648f $X=2.94 $Y=2.315
+ $X2=0 $Y2=0
cc_261 N_A_318_74#_c_244_n N_A_580_74#_c_610_n 0.0213899f $X=2.855 $Y=1.55 $X2=0
+ $Y2=0
cc_262 N_A_318_74#_c_245_n N_A_580_74#_c_610_n 0.0110999f $X=2.94 $Y=1.455 $X2=0
+ $Y2=0
cc_263 N_A_318_74#_c_244_n N_A_580_74#_c_631_n 0.00239474f $X=2.855 $Y=1.55
+ $X2=0 $Y2=0
cc_264 N_A_318_74#_c_245_n N_A_580_74#_c_631_n 0.0116105f $X=2.94 $Y=1.455 $X2=0
+ $Y2=0
cc_265 N_A_318_74#_M1005_g N_VPWR_c_835_n 0.00112709f $X=2.94 $Y=2.315 $X2=0
+ $Y2=0
cc_266 N_A_318_74#_c_242_n N_A_114_112#_c_927_n 0.00245013f $X=1.895 $Y=0.965
+ $X2=0 $Y2=0
cc_267 N_A_318_74#_c_242_n N_A_114_112#_c_942_n 0.00161039f $X=1.895 $Y=0.965
+ $X2=0 $Y2=0
cc_268 N_A_318_74#_M1006_d N_A_114_112#_c_928_n 0.00669515f $X=1.59 $Y=0.37
+ $X2=0 $Y2=0
cc_269 N_A_318_74#_c_242_n N_A_114_112#_c_928_n 0.0261275f $X=1.895 $Y=0.965
+ $X2=0 $Y2=0
cc_270 N_A_318_74#_c_240_n N_A_114_112#_c_930_n 0.0131979f $X=1.895 $Y=1.545
+ $X2=0 $Y2=0
cc_271 N_A_318_74#_c_242_n N_A_114_112#_c_930_n 0.00393441f $X=1.895 $Y=0.965
+ $X2=0 $Y2=0
cc_272 N_A_318_74#_c_240_n N_A_114_112#_c_931_n 0.0116322f $X=1.895 $Y=1.545
+ $X2=0 $Y2=0
cc_273 N_A_318_74#_c_243_n N_A_114_112#_c_931_n 0.0358396f $X=2.34 $Y=1.847
+ $X2=0 $Y2=0
cc_274 N_A_318_74#_M1012_d N_A_114_112#_c_935_n 0.00534086f $X=2.04 $Y=1.84
+ $X2=0 $Y2=0
cc_275 N_A_318_74#_M1005_g N_A_114_112#_c_935_n 0.00232122f $X=2.94 $Y=2.315
+ $X2=0 $Y2=0
cc_276 N_A_318_74#_c_241_n N_A_114_112#_c_935_n 0.00650951f $X=2.69 $Y=1.63
+ $X2=0 $Y2=0
cc_277 N_A_318_74#_c_243_n N_A_114_112#_c_935_n 0.0330524f $X=2.34 $Y=1.847
+ $X2=0 $Y2=0
cc_278 N_A_318_74#_M1005_g N_A_114_112#_c_936_n 0.001764f $X=2.94 $Y=2.315 $X2=0
+ $Y2=0
cc_279 N_A_318_74#_c_241_n N_A_114_112#_c_936_n 0.01174f $X=2.69 $Y=1.63 $X2=0
+ $Y2=0
cc_280 N_A_318_74#_c_243_n N_A_114_112#_c_936_n 0.0193404f $X=2.34 $Y=1.847
+ $X2=0 $Y2=0
cc_281 N_A_318_74#_c_244_n N_A_114_112#_c_936_n 0.00915244f $X=2.855 $Y=1.55
+ $X2=0 $Y2=0
cc_282 N_A_318_74#_c_245_n N_A_114_112#_c_936_n 8.54792e-19 $X=2.94 $Y=1.455
+ $X2=0 $Y2=0
cc_283 N_A_318_74#_M1018_g N_VGND_c_1069_n 9.15902e-19 $X=3.35 $Y=0.615 $X2=0
+ $Y2=0
cc_284 N_A_288_48#_c_332_n N_A_706_317#_M1004_d 0.00253411f $X=4.995 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_285 N_A_288_48#_c_327_n N_A_706_317#_M1019_g 0.00371294f $X=3.53 $Y=0.34
+ $X2=0 $Y2=0
cc_286 N_A_288_48#_c_329_n N_A_706_317#_M1019_g 0.00954024f $X=3.615 $Y=0.905
+ $X2=0 $Y2=0
cc_287 N_A_288_48#_c_330_n N_A_706_317#_M1019_g 0.0112741f $X=4.21 $Y=0.99 $X2=0
+ $Y2=0
cc_288 N_A_288_48#_c_331_n N_A_706_317#_M1019_g 0.00209968f $X=3.7 $Y=0.99 $X2=0
+ $Y2=0
cc_289 N_A_288_48#_c_380_p N_A_706_317#_M1019_g 0.00167035f $X=4.295 $Y=0.905
+ $X2=0 $Y2=0
cc_290 N_A_288_48#_M1013_g N_A_706_317#_M1007_g 0.0412085f $X=3.465 $Y=2.465
+ $X2=0 $Y2=0
cc_291 N_A_288_48#_c_342_n N_A_706_317#_c_489_n 0.0104522f $X=5.145 $Y=1.885
+ $X2=0 $Y2=0
cc_292 N_A_288_48#_c_332_n N_A_706_317#_c_477_n 0.0206246f $X=4.995 $Y=0.34
+ $X2=0 $Y2=0
cc_293 N_A_288_48#_c_334_n N_A_706_317#_c_477_n 0.0307524f $X=5.195 $Y=0.515
+ $X2=0 $Y2=0
cc_294 N_A_288_48#_c_337_n N_A_706_317#_c_478_n 0.0307524f $X=5.152 $Y=1.72
+ $X2=0 $Y2=0
cc_295 N_A_288_48#_M1010_s N_A_706_317#_c_492_n 0.0112283f $X=5.01 $Y=1.74 $X2=0
+ $Y2=0
cc_296 N_A_288_48#_c_342_n N_A_706_317#_c_492_n 0.0202912f $X=5.145 $Y=1.885
+ $X2=0 $Y2=0
cc_297 N_A_288_48#_c_342_n N_A_706_317#_c_479_n 0.00932987f $X=5.145 $Y=1.885
+ $X2=0 $Y2=0
cc_298 N_A_288_48#_c_337_n N_A_706_317#_c_479_n 9.85805e-19 $X=5.152 $Y=1.72
+ $X2=0 $Y2=0
cc_299 N_A_288_48#_c_337_n N_A_706_317#_c_480_n 0.00218999f $X=5.152 $Y=1.72
+ $X2=0 $Y2=0
cc_300 N_A_288_48#_M1013_g N_A_706_317#_c_482_n 5.57125e-19 $X=3.465 $Y=2.465
+ $X2=0 $Y2=0
cc_301 N_A_288_48#_c_342_n N_A_706_317#_c_495_n 0.0149883f $X=5.145 $Y=1.885
+ $X2=0 $Y2=0
cc_302 N_A_288_48#_c_336_n N_A_706_317#_c_483_n 0.0307524f $X=5.177 $Y=1.01
+ $X2=0 $Y2=0
cc_303 N_A_288_48#_M1013_g N_A_706_317#_c_484_n 0.00167735f $X=3.465 $Y=2.465
+ $X2=0 $Y2=0
cc_304 N_A_288_48#_c_327_n N_A_580_74#_M1023_d 0.00281472f $X=3.53 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_305 N_A_288_48#_c_342_n N_A_580_74#_M1000_g 4.42753e-19 $X=5.145 $Y=1.885
+ $X2=0 $Y2=0
cc_306 N_A_288_48#_c_337_n N_A_580_74#_M1000_g 8.28864e-19 $X=5.152 $Y=1.72
+ $X2=0 $Y2=0
cc_307 N_A_288_48#_c_325_n N_A_580_74#_c_619_n 0.00294277f $X=2.825 $Y=0.995
+ $X2=0 $Y2=0
cc_308 N_A_288_48#_c_327_n N_A_580_74#_c_619_n 0.0254752f $X=3.53 $Y=0.34 $X2=0
+ $Y2=0
cc_309 N_A_288_48#_c_329_n N_A_580_74#_c_619_n 0.0191208f $X=3.615 $Y=0.905
+ $X2=0 $Y2=0
cc_310 N_A_288_48#_c_325_n N_A_580_74#_c_608_n 0.0024498f $X=2.825 $Y=0.995
+ $X2=0 $Y2=0
cc_311 N_A_288_48#_c_326_n N_A_580_74#_c_608_n 0.0051404f $X=2.63 $Y=1.03 $X2=0
+ $Y2=0
cc_312 N_A_288_48#_c_329_n N_A_580_74#_c_608_n 0.00421956f $X=3.615 $Y=0.905
+ $X2=0 $Y2=0
cc_313 N_A_288_48#_c_331_n N_A_580_74#_c_608_n 0.0137149f $X=3.7 $Y=0.99 $X2=0
+ $Y2=0
cc_314 N_A_288_48#_c_335_n N_A_580_74#_c_608_n 0.00638342f $X=2.315 $Y=1.195
+ $X2=0 $Y2=0
cc_315 N_A_288_48#_c_330_n N_A_580_74#_c_609_n 0.0332831f $X=4.21 $Y=0.99 $X2=0
+ $Y2=0
cc_316 N_A_288_48#_c_331_n N_A_580_74#_c_609_n 0.0140682f $X=3.7 $Y=0.99 $X2=0
+ $Y2=0
cc_317 N_A_288_48#_c_339_n N_A_580_74#_c_615_n 0.00462717f $X=3.375 $Y=3.15
+ $X2=0 $Y2=0
cc_318 N_A_288_48#_M1013_g N_A_580_74#_c_610_n 0.00465976f $X=3.465 $Y=2.465
+ $X2=0 $Y2=0
cc_319 N_A_288_48#_c_330_n N_A_580_74#_c_611_n 0.0162324f $X=4.21 $Y=0.99 $X2=0
+ $Y2=0
cc_320 N_A_288_48#_c_330_n N_A_580_74#_c_612_n 0.00123174f $X=4.21 $Y=0.99 $X2=0
+ $Y2=0
cc_321 N_A_288_48#_c_329_n N_A_580_74#_c_613_n 2.03258e-19 $X=3.615 $Y=0.905
+ $X2=0 $Y2=0
cc_322 N_A_288_48#_c_330_n N_A_580_74#_c_613_n 0.00554025f $X=4.21 $Y=0.99 $X2=0
+ $Y2=0
cc_323 N_A_288_48#_c_380_p N_A_580_74#_c_613_n 0.0128024f $X=4.295 $Y=0.905
+ $X2=0 $Y2=0
cc_324 N_A_288_48#_c_332_n N_A_580_74#_c_613_n 0.011853f $X=4.995 $Y=0.34 $X2=0
+ $Y2=0
cc_325 N_A_288_48#_c_333_n N_A_580_74#_c_613_n 0.00273646f $X=4.38 $Y=0.34 $X2=0
+ $Y2=0
cc_326 N_A_288_48#_c_334_n N_A_580_74#_c_613_n 0.00468553f $X=5.195 $Y=0.515
+ $X2=0 $Y2=0
cc_327 N_A_288_48#_c_342_n N_CLK_M1010_g 0.00828728f $X=5.145 $Y=1.885 $X2=0
+ $Y2=0
cc_328 N_A_288_48#_c_332_n N_CLK_c_693_n 0.00462641f $X=4.995 $Y=0.34 $X2=0
+ $Y2=0
cc_329 N_A_288_48#_c_334_n N_CLK_c_693_n 0.00451642f $X=5.195 $Y=0.515 $X2=0
+ $Y2=0
cc_330 N_A_288_48#_c_336_n N_CLK_c_693_n 0.00219347f $X=5.177 $Y=1.01 $X2=0
+ $Y2=0
cc_331 N_A_288_48#_c_337_n N_CLK_c_693_n 0.00401029f $X=5.152 $Y=1.72 $X2=0
+ $Y2=0
cc_332 N_A_288_48#_c_342_n N_CLK_M1021_g 9.75393e-19 $X=5.145 $Y=1.885 $X2=0
+ $Y2=0
cc_333 N_A_288_48#_c_336_n CLK 0.00186086f $X=5.177 $Y=1.01 $X2=0 $Y2=0
cc_334 N_A_288_48#_c_337_n CLK 0.0277686f $X=5.152 $Y=1.72 $X2=0 $Y2=0
cc_335 N_A_288_48#_c_337_n N_CLK_c_697_n 0.0124174f $X=5.152 $Y=1.72 $X2=0 $Y2=0
cc_336 N_A_288_48#_M1012_g N_VPWR_c_838_n 0.0240893f $X=1.95 $Y=2.26 $X2=0 $Y2=0
cc_337 N_A_288_48#_M1013_g N_VPWR_c_839_n 0.011579f $X=3.465 $Y=2.465 $X2=0
+ $Y2=0
cc_338 N_A_288_48#_c_340_n N_VPWR_c_847_n 0.0551463f $X=2.04 $Y=3.15 $X2=0 $Y2=0
cc_339 N_A_288_48#_c_339_n N_VPWR_c_835_n 0.0535024f $X=3.375 $Y=3.15 $X2=0
+ $Y2=0
cc_340 N_A_288_48#_c_340_n N_VPWR_c_835_n 0.00797315f $X=2.04 $Y=3.15 $X2=0
+ $Y2=0
cc_341 N_A_288_48#_c_326_n N_A_114_112#_M1023_s 0.0122448f $X=2.63 $Y=1.03 $X2=0
+ $Y2=0
cc_342 N_A_288_48#_c_328_n N_A_114_112#_M1023_s 6.86248e-19 $X=2.715 $Y=0.34
+ $X2=0 $Y2=0
cc_343 N_A_288_48#_c_319_n N_A_114_112#_c_927_n 0.00112866f $X=1.515 $Y=1.21
+ $X2=0 $Y2=0
cc_344 N_A_288_48#_c_319_n N_A_114_112#_c_942_n 0.00100301f $X=1.515 $Y=1.21
+ $X2=0 $Y2=0
cc_345 N_A_288_48#_c_319_n N_A_114_112#_c_928_n 0.0150312f $X=1.515 $Y=1.21
+ $X2=0 $Y2=0
cc_346 N_A_288_48#_c_324_n N_A_114_112#_c_928_n 0.00226467f $X=2.48 $Y=1.07
+ $X2=0 $Y2=0
cc_347 N_A_288_48#_c_320_n N_A_114_112#_c_930_n 0.00461745f $X=1.86 $Y=1.285
+ $X2=0 $Y2=0
cc_348 N_A_288_48#_c_321_n N_A_114_112#_c_930_n 0.011085f $X=1.59 $Y=1.285 $X2=0
+ $Y2=0
cc_349 N_A_288_48#_M1012_g N_A_114_112#_c_930_n 2.01632e-19 $X=1.95 $Y=2.26
+ $X2=0 $Y2=0
cc_350 N_A_288_48#_M1012_g N_A_114_112#_c_931_n 0.0103431f $X=1.95 $Y=2.26 $X2=0
+ $Y2=0
cc_351 N_A_288_48#_M1012_g N_A_114_112#_c_935_n 0.0245763f $X=1.95 $Y=2.26 $X2=0
+ $Y2=0
cc_352 N_A_288_48#_c_339_n N_A_114_112#_c_935_n 0.0144075f $X=3.375 $Y=3.15
+ $X2=0 $Y2=0
cc_353 N_A_288_48#_M1012_g N_A_114_112#_c_936_n 0.00398344f $X=1.95 $Y=2.26
+ $X2=0 $Y2=0
cc_354 N_A_288_48#_M1012_g N_A_114_112#_c_937_n 0.00463211f $X=1.95 $Y=2.26
+ $X2=0 $Y2=0
cc_355 N_A_288_48#_c_319_n N_A_114_112#_c_932_n 0.00504475f $X=1.515 $Y=1.21
+ $X2=0 $Y2=0
cc_356 N_A_288_48#_c_324_n N_A_114_112#_c_932_n 0.00493278f $X=2.48 $Y=1.07
+ $X2=0 $Y2=0
cc_357 N_A_288_48#_c_325_n N_A_114_112#_c_932_n 8.15455e-19 $X=2.825 $Y=0.995
+ $X2=0 $Y2=0
cc_358 N_A_288_48#_c_326_n N_A_114_112#_c_932_n 0.0212796f $X=2.63 $Y=1.03 $X2=0
+ $Y2=0
cc_359 N_A_288_48#_c_328_n N_A_114_112#_c_932_n 0.00632876f $X=2.715 $Y=0.34
+ $X2=0 $Y2=0
cc_360 N_A_288_48#_c_335_n N_A_114_112#_c_932_n 0.0108433f $X=2.315 $Y=1.195
+ $X2=0 $Y2=0
cc_361 N_A_288_48#_c_330_n N_VGND_M1019_d 0.00676444f $X=4.21 $Y=0.99 $X2=0
+ $Y2=0
cc_362 N_A_288_48#_c_380_p N_VGND_M1019_d 0.00511615f $X=4.295 $Y=0.905 $X2=0
+ $Y2=0
cc_363 N_A_288_48#_c_327_n N_VGND_c_1064_n 0.0128817f $X=3.53 $Y=0.34 $X2=0
+ $Y2=0
cc_364 N_A_288_48#_c_330_n N_VGND_c_1064_n 0.013847f $X=4.21 $Y=0.99 $X2=0 $Y2=0
cc_365 N_A_288_48#_c_380_p N_VGND_c_1064_n 0.0224799f $X=4.295 $Y=0.905 $X2=0
+ $Y2=0
cc_366 N_A_288_48#_c_333_n N_VGND_c_1064_n 0.0142952f $X=4.38 $Y=0.34 $X2=0
+ $Y2=0
cc_367 N_A_288_48#_c_332_n N_VGND_c_1065_n 0.011924f $X=4.995 $Y=0.34 $X2=0
+ $Y2=0
cc_368 N_A_288_48#_c_319_n N_VGND_c_1069_n 0.00315544f $X=1.515 $Y=1.21 $X2=0
+ $Y2=0
cc_369 N_A_288_48#_c_325_n N_VGND_c_1069_n 0.00278271f $X=2.825 $Y=0.995 $X2=0
+ $Y2=0
cc_370 N_A_288_48#_c_327_n N_VGND_c_1069_n 0.0641927f $X=3.53 $Y=0.34 $X2=0
+ $Y2=0
cc_371 N_A_288_48#_c_328_n N_VGND_c_1069_n 0.0121867f $X=2.715 $Y=0.34 $X2=0
+ $Y2=0
cc_372 N_A_288_48#_c_332_n N_VGND_c_1071_n 0.0656368f $X=4.995 $Y=0.34 $X2=0
+ $Y2=0
cc_373 N_A_288_48#_c_333_n N_VGND_c_1071_n 0.0121867f $X=4.38 $Y=0.34 $X2=0
+ $Y2=0
cc_374 N_A_288_48#_c_319_n N_VGND_c_1076_n 0.00542971f $X=1.515 $Y=1.21 $X2=0
+ $Y2=0
cc_375 N_A_288_48#_c_319_n N_VGND_c_1078_n 0.00400711f $X=1.515 $Y=1.21 $X2=0
+ $Y2=0
cc_376 N_A_288_48#_c_325_n N_VGND_c_1078_n 0.00363426f $X=2.825 $Y=0.995 $X2=0
+ $Y2=0
cc_377 N_A_288_48#_c_327_n N_VGND_c_1078_n 0.0365608f $X=3.53 $Y=0.34 $X2=0
+ $Y2=0
cc_378 N_A_288_48#_c_328_n N_VGND_c_1078_n 0.00660921f $X=2.715 $Y=0.34 $X2=0
+ $Y2=0
cc_379 N_A_288_48#_c_332_n N_VGND_c_1078_n 0.0371906f $X=4.995 $Y=0.34 $X2=0
+ $Y2=0
cc_380 N_A_288_48#_c_333_n N_VGND_c_1078_n 0.00660921f $X=4.38 $Y=0.34 $X2=0
+ $Y2=0
cc_381 N_A_288_48#_c_327_n A_685_81# 0.00179331f $X=3.53 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_382 N_A_288_48#_c_329_n A_685_81# 0.00376627f $X=3.615 $Y=0.905 $X2=-0.19
+ $Y2=-0.245
cc_383 N_A_706_317#_c_488_n N_A_580_74#_M1000_g 0.0133018f $X=4.44 $Y=1.84 $X2=0
+ $Y2=0
cc_384 N_A_706_317#_c_489_n N_A_580_74#_M1000_g 0.00548407f $X=4.632 $Y=2.22
+ $X2=0 $Y2=0
cc_385 N_A_706_317#_c_490_n N_A_580_74#_M1000_g 0.00766689f $X=4.605 $Y=2.755
+ $X2=0 $Y2=0
cc_386 N_A_706_317#_c_478_n N_A_580_74#_M1000_g 0.00410983f $X=4.74 $Y=1.755
+ $X2=0 $Y2=0
cc_387 N_A_706_317#_c_482_n N_A_580_74#_M1000_g 9.71511e-19 $X=3.695 $Y=1.75
+ $X2=0 $Y2=0
cc_388 N_A_706_317#_c_495_n N_A_580_74#_M1000_g 0.00140227f $X=4.632 $Y=1.84
+ $X2=0 $Y2=0
cc_389 N_A_706_317#_c_496_n N_A_580_74#_M1000_g 0.00205065f $X=4.632 $Y=2.305
+ $X2=0 $Y2=0
cc_390 N_A_706_317#_c_484_n N_A_580_74#_M1000_g 0.0292862f $X=3.855 $Y=1.75
+ $X2=0 $Y2=0
cc_391 N_A_706_317#_M1019_g N_A_580_74#_c_619_n 2.25119e-19 $X=3.74 $Y=0.615
+ $X2=0 $Y2=0
cc_392 N_A_706_317#_M1019_g N_A_580_74#_c_608_n 0.00116521f $X=3.74 $Y=0.615
+ $X2=0 $Y2=0
cc_393 N_A_706_317#_M1019_g N_A_580_74#_c_609_n 0.0107958f $X=3.74 $Y=0.615
+ $X2=0 $Y2=0
cc_394 N_A_706_317#_c_488_n N_A_580_74#_c_609_n 0.0134189f $X=4.44 $Y=1.84 $X2=0
+ $Y2=0
cc_395 N_A_706_317#_c_482_n N_A_580_74#_c_609_n 0.0242682f $X=3.695 $Y=1.75
+ $X2=0 $Y2=0
cc_396 N_A_706_317#_c_484_n N_A_580_74#_c_609_n 0.00369392f $X=3.855 $Y=1.75
+ $X2=0 $Y2=0
cc_397 N_A_706_317#_M1019_g N_A_580_74#_c_610_n 0.00310402f $X=3.74 $Y=0.615
+ $X2=0 $Y2=0
cc_398 N_A_706_317#_M1007_g N_A_580_74#_c_610_n 0.00620393f $X=3.855 $Y=2.465
+ $X2=0 $Y2=0
cc_399 N_A_706_317#_c_482_n N_A_580_74#_c_610_n 0.0255945f $X=3.695 $Y=1.75
+ $X2=0 $Y2=0
cc_400 N_A_706_317#_c_484_n N_A_580_74#_c_610_n 0.00258641f $X=3.855 $Y=1.75
+ $X2=0 $Y2=0
cc_401 N_A_706_317#_M1019_g N_A_580_74#_c_611_n 0.00113382f $X=3.74 $Y=0.615
+ $X2=0 $Y2=0
cc_402 N_A_706_317#_c_488_n N_A_580_74#_c_611_n 0.0209034f $X=4.44 $Y=1.84 $X2=0
+ $Y2=0
cc_403 N_A_706_317#_c_478_n N_A_580_74#_c_611_n 0.0255154f $X=4.74 $Y=1.755
+ $X2=0 $Y2=0
cc_404 N_A_706_317#_c_495_n N_A_580_74#_c_611_n 0.00360126f $X=4.632 $Y=1.84
+ $X2=0 $Y2=0
cc_405 N_A_706_317#_M1019_g N_A_580_74#_c_612_n 0.012245f $X=3.74 $Y=0.615 $X2=0
+ $Y2=0
cc_406 N_A_706_317#_c_488_n N_A_580_74#_c_612_n 9.4463e-19 $X=4.44 $Y=1.84 $X2=0
+ $Y2=0
cc_407 N_A_706_317#_c_495_n N_A_580_74#_c_612_n 6.41724e-19 $X=4.632 $Y=1.84
+ $X2=0 $Y2=0
cc_408 N_A_706_317#_M1019_g N_A_580_74#_c_613_n 0.0154325f $X=3.74 $Y=0.615
+ $X2=0 $Y2=0
cc_409 N_A_706_317#_c_478_n N_A_580_74#_c_613_n 0.0118613f $X=4.74 $Y=1.755
+ $X2=0 $Y2=0
cc_410 N_A_706_317#_c_489_n N_CLK_M1010_g 0.0044461f $X=4.632 $Y=2.22 $X2=0
+ $Y2=0
cc_411 N_A_706_317#_c_490_n N_CLK_M1010_g 0.0091196f $X=4.605 $Y=2.755 $X2=0
+ $Y2=0
cc_412 N_A_706_317#_c_478_n N_CLK_M1010_g 0.001416f $X=4.74 $Y=1.755 $X2=0 $Y2=0
cc_413 N_A_706_317#_c_492_n N_CLK_M1010_g 0.0216723f $X=5.835 $Y=2.305 $X2=0
+ $Y2=0
cc_414 N_A_706_317#_c_479_n N_CLK_M1010_g 0.00267871f $X=5.92 $Y=2.22 $X2=0
+ $Y2=0
cc_415 N_A_706_317#_c_480_n N_CLK_M1010_g 3.09558e-19 $X=6.005 $Y=1.465 $X2=0
+ $Y2=0
cc_416 N_A_706_317#_c_477_n N_CLK_c_693_n 5.87969e-19 $X=4.635 $Y=0.835 $X2=0
+ $Y2=0
cc_417 N_A_706_317#_M1020_g N_CLK_M1021_g 0.0173598f $X=6.565 $Y=2.37 $X2=0
+ $Y2=0
cc_418 N_A_706_317#_c_492_n N_CLK_M1021_g 0.0153829f $X=5.835 $Y=2.305 $X2=0
+ $Y2=0
cc_419 N_A_706_317#_c_479_n N_CLK_M1021_g 0.0206291f $X=5.92 $Y=2.22 $X2=0 $Y2=0
cc_420 N_A_706_317#_c_480_n N_CLK_M1021_g 0.0030238f $X=6.005 $Y=1.465 $X2=0
+ $Y2=0
cc_421 N_A_706_317#_M1011_g N_CLK_c_695_n 0.042261f $X=6.275 $Y=0.74 $X2=0 $Y2=0
cc_422 N_A_706_317#_M1011_g CLK 2.78077e-19 $X=6.275 $Y=0.74 $X2=0 $Y2=0
cc_423 N_A_706_317#_c_492_n CLK 0.00722814f $X=5.835 $Y=2.305 $X2=0 $Y2=0
cc_424 N_A_706_317#_c_480_n CLK 0.0199911f $X=6.005 $Y=1.465 $X2=0 $Y2=0
cc_425 N_A_706_317#_c_492_n N_CLK_c_697_n 0.00180527f $X=5.835 $Y=2.305 $X2=0
+ $Y2=0
cc_426 N_A_706_317#_c_480_n N_CLK_c_697_n 0.0168212f $X=6.005 $Y=1.465 $X2=0
+ $Y2=0
cc_427 N_A_706_317#_c_485_n N_CLK_c_697_n 0.042261f $X=6.565 $Y=1.465 $X2=0
+ $Y2=0
cc_428 N_A_706_317#_M1020_g N_A_1198_374#_M1001_g 0.0224304f $X=6.565 $Y=2.37
+ $X2=0 $Y2=0
cc_429 N_A_706_317#_M1020_g N_A_1198_374#_c_758_n 0.0133662f $X=6.565 $Y=2.37
+ $X2=0 $Y2=0
cc_430 N_A_706_317#_M1011_g N_A_1198_374#_c_749_n 0.0115865f $X=6.275 $Y=0.74
+ $X2=0 $Y2=0
cc_431 N_A_706_317#_M1020_g N_A_1198_374#_c_759_n 0.0148982f $X=6.565 $Y=2.37
+ $X2=0 $Y2=0
cc_432 N_A_706_317#_c_481_n N_A_1198_374#_c_759_n 0.00175142f $X=6.365 $Y=1.465
+ $X2=0 $Y2=0
cc_433 N_A_706_317#_M1020_g N_A_1198_374#_c_760_n 0.00189286f $X=6.565 $Y=2.37
+ $X2=0 $Y2=0
cc_434 N_A_706_317#_c_479_n N_A_1198_374#_c_760_n 0.0103611f $X=5.92 $Y=2.22
+ $X2=0 $Y2=0
cc_435 N_A_706_317#_c_481_n N_A_1198_374#_c_760_n 0.0277979f $X=6.365 $Y=1.465
+ $X2=0 $Y2=0
cc_436 N_A_706_317#_c_485_n N_A_1198_374#_c_760_n 0.00699793f $X=6.565 $Y=1.465
+ $X2=0 $Y2=0
cc_437 N_A_706_317#_M1011_g N_A_1198_374#_c_751_n 0.0038748f $X=6.275 $Y=0.74
+ $X2=0 $Y2=0
cc_438 N_A_706_317#_c_481_n N_A_1198_374#_c_751_n 0.0171756f $X=6.365 $Y=1.465
+ $X2=0 $Y2=0
cc_439 N_A_706_317#_c_485_n N_A_1198_374#_c_751_n 0.0086752f $X=6.565 $Y=1.465
+ $X2=0 $Y2=0
cc_440 N_A_706_317#_M1020_g N_A_1198_374#_c_752_n 0.00307306f $X=6.565 $Y=2.37
+ $X2=0 $Y2=0
cc_441 N_A_706_317#_c_481_n N_A_1198_374#_c_753_n 0.0164832f $X=6.365 $Y=1.465
+ $X2=0 $Y2=0
cc_442 N_A_706_317#_c_485_n N_A_1198_374#_c_753_n 0.00307306f $X=6.565 $Y=1.465
+ $X2=0 $Y2=0
cc_443 N_A_706_317#_M1011_g N_A_1198_374#_c_754_n 0.00399952f $X=6.275 $Y=0.74
+ $X2=0 $Y2=0
cc_444 N_A_706_317#_c_481_n N_A_1198_374#_c_755_n 3.30771e-19 $X=6.365 $Y=1.465
+ $X2=0 $Y2=0
cc_445 N_A_706_317#_c_485_n N_A_1198_374#_c_755_n 0.0180242f $X=6.565 $Y=1.465
+ $X2=0 $Y2=0
cc_446 N_A_706_317#_c_488_n N_VPWR_M1007_d 0.00226423f $X=4.44 $Y=1.84 $X2=0
+ $Y2=0
cc_447 N_A_706_317#_c_492_n N_VPWR_M1010_d 0.00755771f $X=5.835 $Y=2.305 $X2=0
+ $Y2=0
cc_448 N_A_706_317#_M1007_g N_VPWR_c_839_n 0.00787223f $X=3.855 $Y=2.465 $X2=0
+ $Y2=0
cc_449 N_A_706_317#_c_488_n N_VPWR_c_839_n 0.0197787f $X=4.44 $Y=1.84 $X2=0
+ $Y2=0
cc_450 N_A_706_317#_c_490_n N_VPWR_c_839_n 0.0185201f $X=4.605 $Y=2.755 $X2=0
+ $Y2=0
cc_451 N_A_706_317#_M1020_g N_VPWR_c_840_n 5.85824e-19 $X=6.565 $Y=2.37 $X2=0
+ $Y2=0
cc_452 N_A_706_317#_c_492_n N_VPWR_c_840_n 0.0210288f $X=5.835 $Y=2.305 $X2=0
+ $Y2=0
cc_453 N_A_706_317#_M1020_g N_VPWR_c_841_n 0.00776968f $X=6.565 $Y=2.37 $X2=0
+ $Y2=0
cc_454 N_A_706_317#_M1020_g N_VPWR_c_844_n 0.00589836f $X=6.565 $Y=2.37 $X2=0
+ $Y2=0
cc_455 N_A_706_317#_M1007_g N_VPWR_c_847_n 0.00479829f $X=3.855 $Y=2.465 $X2=0
+ $Y2=0
cc_456 N_A_706_317#_c_490_n N_VPWR_c_848_n 0.0136788f $X=4.605 $Y=2.755 $X2=0
+ $Y2=0
cc_457 N_A_706_317#_M1007_g N_VPWR_c_835_n 0.00553463f $X=3.855 $Y=2.465 $X2=0
+ $Y2=0
cc_458 N_A_706_317#_M1020_g N_VPWR_c_835_n 0.00620995f $X=6.565 $Y=2.37 $X2=0
+ $Y2=0
cc_459 N_A_706_317#_c_490_n N_VPWR_c_835_n 0.0135953f $X=4.605 $Y=2.755 $X2=0
+ $Y2=0
cc_460 N_A_706_317#_M1020_g GCLK 0.0010233f $X=6.565 $Y=2.37 $X2=0 $Y2=0
cc_461 N_A_706_317#_M1019_g N_VGND_c_1064_n 0.0012897f $X=3.74 $Y=0.615 $X2=0
+ $Y2=0
cc_462 N_A_706_317#_M1011_g N_VGND_c_1065_n 0.00234521f $X=6.275 $Y=0.74 $X2=0
+ $Y2=0
cc_463 N_A_706_317#_c_480_n N_VGND_c_1065_n 0.00115537f $X=6.005 $Y=1.465 $X2=0
+ $Y2=0
cc_464 N_A_706_317#_M1011_g N_VGND_c_1066_n 0.00356081f $X=6.275 $Y=0.74 $X2=0
+ $Y2=0
cc_465 N_A_706_317#_M1019_g N_VGND_c_1069_n 0.00444804f $X=3.74 $Y=0.615 $X2=0
+ $Y2=0
cc_466 N_A_706_317#_M1011_g N_VGND_c_1074_n 0.00434272f $X=6.275 $Y=0.74 $X2=0
+ $Y2=0
cc_467 N_A_706_317#_M1019_g N_VGND_c_1078_n 0.00409911f $X=3.74 $Y=0.615 $X2=0
+ $Y2=0
cc_468 N_A_706_317#_M1011_g N_VGND_c_1078_n 0.00825669f $X=6.275 $Y=0.74 $X2=0
+ $Y2=0
cc_469 N_A_580_74#_M1000_g N_VPWR_c_839_n 0.00561192f $X=4.38 $Y=2.34 $X2=0
+ $Y2=0
cc_470 N_A_580_74#_c_610_n N_VPWR_c_839_n 0.00549938f $X=3.18 $Y=2.235 $X2=0
+ $Y2=0
cc_471 N_A_580_74#_c_615_n N_VPWR_c_847_n 0.00630871f $X=3.165 $Y=2.465 $X2=0
+ $Y2=0
cc_472 N_A_580_74#_M1000_g N_VPWR_c_848_n 0.00612719f $X=4.38 $Y=2.34 $X2=0
+ $Y2=0
cc_473 N_A_580_74#_M1000_g N_VPWR_c_835_n 0.00632145f $X=4.38 $Y=2.34 $X2=0
+ $Y2=0
cc_474 N_A_580_74#_c_615_n N_VPWR_c_835_n 0.00932018f $X=3.165 $Y=2.465 $X2=0
+ $Y2=0
cc_475 N_A_580_74#_c_610_n N_A_114_112#_c_936_n 0.00708697f $X=3.18 $Y=2.235
+ $X2=0 $Y2=0
cc_476 N_A_580_74#_c_613_n N_VGND_c_1064_n 0.00126464f $X=4.325 $Y=1.255 $X2=0
+ $Y2=0
cc_477 N_A_580_74#_c_613_n N_VGND_c_1071_n 9.34772e-19 $X=4.325 $Y=1.255 $X2=0
+ $Y2=0
cc_478 N_CLK_M1021_g N_A_1198_374#_c_758_n 0.00926161f $X=5.9 $Y=2.37 $X2=0
+ $Y2=0
cc_479 N_CLK_c_695_n N_A_1198_374#_c_749_n 0.0016642f $X=5.915 $Y=1.22 $X2=0
+ $Y2=0
cc_480 N_CLK_M1021_g N_A_1198_374#_c_760_n 7.54259e-19 $X=5.9 $Y=2.37 $X2=0
+ $Y2=0
cc_481 N_CLK_c_695_n N_A_1198_374#_c_751_n 7.31697e-19 $X=5.915 $Y=1.22 $X2=0
+ $Y2=0
cc_482 N_CLK_M1010_g N_VPWR_c_840_n 0.00377698f $X=5.37 $Y=2.16 $X2=0 $Y2=0
cc_483 N_CLK_M1021_g N_VPWR_c_840_n 0.0111311f $X=5.9 $Y=2.37 $X2=0 $Y2=0
cc_484 N_CLK_M1021_g N_VPWR_c_844_n 0.00512593f $X=5.9 $Y=2.37 $X2=0 $Y2=0
cc_485 N_CLK_M1010_g N_VPWR_c_848_n 0.00426167f $X=5.37 $Y=2.16 $X2=0 $Y2=0
cc_486 N_CLK_M1010_g N_VPWR_c_835_n 0.00523464f $X=5.37 $Y=2.16 $X2=0 $Y2=0
cc_487 N_CLK_M1021_g N_VPWR_c_835_n 0.00520946f $X=5.9 $Y=2.37 $X2=0 $Y2=0
cc_488 N_CLK_c_693_n N_VGND_c_1065_n 0.00475792f $X=5.41 $Y=1.22 $X2=0 $Y2=0
cc_489 N_CLK_c_695_n N_VGND_c_1065_n 0.0147865f $X=5.915 $Y=1.22 $X2=0 $Y2=0
cc_490 CLK N_VGND_c_1065_n 0.0111858f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_491 N_CLK_c_697_n N_VGND_c_1065_n 0.00440608f $X=5.915 $Y=1.385 $X2=0 $Y2=0
cc_492 N_CLK_c_693_n N_VGND_c_1071_n 0.00430908f $X=5.41 $Y=1.22 $X2=0 $Y2=0
cc_493 N_CLK_c_695_n N_VGND_c_1074_n 0.00398535f $X=5.915 $Y=1.22 $X2=0 $Y2=0
cc_494 N_CLK_c_693_n N_VGND_c_1078_n 0.00821159f $X=5.41 $Y=1.22 $X2=0 $Y2=0
cc_495 N_CLK_c_695_n N_VGND_c_1078_n 0.00786935f $X=5.915 $Y=1.22 $X2=0 $Y2=0
cc_496 N_A_1198_374#_c_759_n N_VPWR_M1020_d 0.00434052f $X=6.87 $Y=1.885 $X2=0
+ $Y2=0
cc_497 N_A_1198_374#_c_758_n N_VPWR_c_840_n 0.0152573f $X=6.34 $Y=2.015 $X2=0
+ $Y2=0
cc_498 N_A_1198_374#_M1001_g N_VPWR_c_841_n 0.00554989f $X=7.15 $Y=2.4 $X2=0
+ $Y2=0
cc_499 N_A_1198_374#_c_758_n N_VPWR_c_841_n 0.0249197f $X=6.34 $Y=2.015 $X2=0
+ $Y2=0
cc_500 N_A_1198_374#_c_759_n N_VPWR_c_841_n 0.0248097f $X=6.87 $Y=1.885 $X2=0
+ $Y2=0
cc_501 N_A_1198_374#_c_755_n N_VPWR_c_841_n 4.97899e-19 $X=7.6 $Y=1.465 $X2=0
+ $Y2=0
cc_502 N_A_1198_374#_M1003_g N_VPWR_c_843_n 0.0064767f $X=7.6 $Y=2.4 $X2=0 $Y2=0
cc_503 N_A_1198_374#_c_755_n N_VPWR_c_843_n 3.5215e-19 $X=7.6 $Y=1.465 $X2=0
+ $Y2=0
cc_504 N_A_1198_374#_c_758_n N_VPWR_c_844_n 0.0106486f $X=6.34 $Y=2.015 $X2=0
+ $Y2=0
cc_505 N_A_1198_374#_M1001_g N_VPWR_c_849_n 0.005209f $X=7.15 $Y=2.4 $X2=0 $Y2=0
cc_506 N_A_1198_374#_M1003_g N_VPWR_c_849_n 0.00492575f $X=7.6 $Y=2.4 $X2=0
+ $Y2=0
cc_507 N_A_1198_374#_M1001_g N_VPWR_c_835_n 0.00986727f $X=7.15 $Y=2.4 $X2=0
+ $Y2=0
cc_508 N_A_1198_374#_M1003_g N_VPWR_c_835_n 0.00894467f $X=7.6 $Y=2.4 $X2=0
+ $Y2=0
cc_509 N_A_1198_374#_c_758_n N_VPWR_c_835_n 0.0114079f $X=6.34 $Y=2.015 $X2=0
+ $Y2=0
cc_510 N_A_1198_374#_M1009_g N_GCLK_c_1025_n 0.00969649f $X=7.245 $Y=0.74 $X2=0
+ $Y2=0
cc_511 N_A_1198_374#_M1017_g N_GCLK_c_1025_n 0.00788704f $X=7.675 $Y=0.74 $X2=0
+ $Y2=0
cc_512 N_A_1198_374#_c_749_n N_GCLK_c_1025_n 0.00490352f $X=6.49 $Y=0.515 $X2=0
+ $Y2=0
cc_513 N_A_1198_374#_c_750_n N_GCLK_c_1025_n 0.0103299f $X=6.87 $Y=1.045 $X2=0
+ $Y2=0
cc_514 N_A_1198_374#_M1009_g N_GCLK_c_1026_n 0.00359373f $X=7.245 $Y=0.74 $X2=0
+ $Y2=0
cc_515 N_A_1198_374#_M1017_g N_GCLK_c_1026_n 0.00327512f $X=7.675 $Y=0.74 $X2=0
+ $Y2=0
cc_516 N_A_1198_374#_M1001_g GCLK 0.00352266f $X=7.15 $Y=2.4 $X2=0 $Y2=0
cc_517 N_A_1198_374#_M1003_g GCLK 0.00263013f $X=7.6 $Y=2.4 $X2=0 $Y2=0
cc_518 N_A_1198_374#_c_759_n GCLK 0.0066044f $X=6.87 $Y=1.885 $X2=0 $Y2=0
cc_519 N_A_1198_374#_c_753_n GCLK 9.53215e-19 $X=7.06 $Y=1.465 $X2=0 $Y2=0
cc_520 N_A_1198_374#_c_755_n GCLK 0.00307792f $X=7.6 $Y=1.465 $X2=0 $Y2=0
cc_521 N_A_1198_374#_M1001_g GCLK 0.0136822f $X=7.15 $Y=2.4 $X2=0 $Y2=0
cc_522 N_A_1198_374#_M1003_g GCLK 0.0146989f $X=7.6 $Y=2.4 $X2=0 $Y2=0
cc_523 N_A_1198_374#_M1001_g N_GCLK_c_1027_n 0.00148164f $X=7.15 $Y=2.4 $X2=0
+ $Y2=0
cc_524 N_A_1198_374#_M1009_g N_GCLK_c_1027_n 0.00154761f $X=7.245 $Y=0.74 $X2=0
+ $Y2=0
cc_525 N_A_1198_374#_M1003_g N_GCLK_c_1027_n 0.00929518f $X=7.6 $Y=2.4 $X2=0
+ $Y2=0
cc_526 N_A_1198_374#_M1017_g N_GCLK_c_1027_n 0.00413752f $X=7.675 $Y=0.74 $X2=0
+ $Y2=0
cc_527 N_A_1198_374#_c_759_n N_GCLK_c_1027_n 9.86568e-19 $X=6.87 $Y=1.885 $X2=0
+ $Y2=0
cc_528 N_A_1198_374#_c_752_n N_GCLK_c_1027_n 0.00762005f $X=6.955 $Y=1.8 $X2=0
+ $Y2=0
cc_529 N_A_1198_374#_c_753_n N_GCLK_c_1027_n 0.0237053f $X=7.06 $Y=1.465 $X2=0
+ $Y2=0
cc_530 N_A_1198_374#_c_754_n N_GCLK_c_1027_n 0.00759747f $X=7.047 $Y=1.3 $X2=0
+ $Y2=0
cc_531 N_A_1198_374#_c_755_n N_GCLK_c_1027_n 0.0255254f $X=7.6 $Y=1.465 $X2=0
+ $Y2=0
cc_532 N_A_1198_374#_c_750_n N_VGND_M1009_s 0.00432991f $X=6.87 $Y=1.045 $X2=0
+ $Y2=0
cc_533 N_A_1198_374#_c_749_n N_VGND_c_1065_n 0.0202037f $X=6.49 $Y=0.515 $X2=0
+ $Y2=0
cc_534 N_A_1198_374#_c_751_n N_VGND_c_1065_n 0.001765f $X=6.655 $Y=1.045 $X2=0
+ $Y2=0
cc_535 N_A_1198_374#_M1009_g N_VGND_c_1066_n 0.00545557f $X=7.245 $Y=0.74 $X2=0
+ $Y2=0
cc_536 N_A_1198_374#_c_749_n N_VGND_c_1066_n 0.0309452f $X=6.49 $Y=0.515 $X2=0
+ $Y2=0
cc_537 N_A_1198_374#_c_750_n N_VGND_c_1066_n 0.0154159f $X=6.87 $Y=1.045 $X2=0
+ $Y2=0
cc_538 N_A_1198_374#_c_753_n N_VGND_c_1066_n 0.00258618f $X=7.06 $Y=1.465 $X2=0
+ $Y2=0
cc_539 N_A_1198_374#_c_755_n N_VGND_c_1066_n 0.00104545f $X=7.6 $Y=1.465 $X2=0
+ $Y2=0
cc_540 N_A_1198_374#_M1017_g N_VGND_c_1068_n 0.00647412f $X=7.675 $Y=0.74 $X2=0
+ $Y2=0
cc_541 N_A_1198_374#_c_749_n N_VGND_c_1074_n 0.0145639f $X=6.49 $Y=0.515 $X2=0
+ $Y2=0
cc_542 N_A_1198_374#_M1009_g N_VGND_c_1075_n 0.00434272f $X=7.245 $Y=0.74 $X2=0
+ $Y2=0
cc_543 N_A_1198_374#_M1017_g N_VGND_c_1075_n 0.00434272f $X=7.675 $Y=0.74 $X2=0
+ $Y2=0
cc_544 N_A_1198_374#_M1009_g N_VGND_c_1078_n 0.00825283f $X=7.245 $Y=0.74 $X2=0
+ $Y2=0
cc_545 N_A_1198_374#_M1017_g N_VGND_c_1078_n 0.00823907f $X=7.675 $Y=0.74 $X2=0
+ $Y2=0
cc_546 N_A_1198_374#_c_749_n N_VGND_c_1078_n 0.0119984f $X=6.49 $Y=0.515 $X2=0
+ $Y2=0
cc_547 N_VPWR_c_835_n N_A_114_112#_c_933_n 0.00670752f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_548 N_VPWR_M1012_s N_A_114_112#_c_931_n 0.00795928f $X=1.515 $Y=1.84 $X2=0
+ $Y2=0
cc_549 N_VPWR_M1012_s N_A_114_112#_c_935_n 0.0082426f $X=1.515 $Y=1.84 $X2=0
+ $Y2=0
cc_550 N_VPWR_c_838_n N_A_114_112#_c_935_n 0.0129362f $X=1.65 $Y=2.825 $X2=0
+ $Y2=0
cc_551 N_VPWR_c_847_n N_A_114_112#_c_935_n 0.00575553f $X=3.99 $Y=3.33 $X2=0
+ $Y2=0
cc_552 N_VPWR_c_835_n N_A_114_112#_c_935_n 0.0296734f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_553 N_VPWR_c_837_n N_A_114_112#_c_937_n 0.0204878f $X=0.27 $Y=2.295 $X2=0
+ $Y2=0
cc_554 N_VPWR_c_838_n N_A_114_112#_c_937_n 0.0229788f $X=1.65 $Y=2.825 $X2=0
+ $Y2=0
cc_555 N_VPWR_c_846_n N_A_114_112#_c_937_n 0.0145175f $X=1.485 $Y=3.33 $X2=0
+ $Y2=0
cc_556 N_VPWR_c_835_n N_A_114_112#_c_937_n 0.0119619f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_557 N_VPWR_M1012_s N_A_114_112#_c_938_n 0.00252977f $X=1.515 $Y=1.84 $X2=0
+ $Y2=0
cc_558 N_VPWR_c_838_n N_A_114_112#_c_938_n 0.0136075f $X=1.65 $Y=2.825 $X2=0
+ $Y2=0
cc_559 N_VPWR_c_835_n N_A_114_112#_c_938_n 0.00116919f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_560 N_VPWR_c_843_n GCLK 0.0444514f $X=7.825 $Y=1.985 $X2=0 $Y2=0
cc_561 N_VPWR_c_841_n GCLK 0.0326636f $X=6.875 $Y=2.305 $X2=0 $Y2=0
cc_562 N_VPWR_c_849_n GCLK 0.0155031f $X=7.74 $Y=3.33 $X2=0 $Y2=0
cc_563 N_VPWR_c_835_n GCLK 0.0126371f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_564 N_A_114_112#_c_928_n N_VGND_M1014_d 0.00932283f $X=2.125 $Y=0.625 $X2=0
+ $Y2=0
cc_565 N_A_114_112#_c_927_n N_VGND_c_1063_n 0.00658627f $X=0.717 $Y=0.948 $X2=0
+ $Y2=0
cc_566 N_A_114_112#_c_929_n N_VGND_c_1063_n 0.00756924f $X=0.89 $Y=0.625 $X2=0
+ $Y2=0
cc_567 N_A_114_112#_c_928_n N_VGND_c_1069_n 0.0151441f $X=2.125 $Y=0.625 $X2=0
+ $Y2=0
cc_568 N_A_114_112#_c_932_n N_VGND_c_1069_n 0.0105752f $X=2.29 $Y=0.53 $X2=0
+ $Y2=0
cc_569 N_A_114_112#_c_928_n N_VGND_c_1073_n 0.00350553f $X=2.125 $Y=0.625 $X2=0
+ $Y2=0
cc_570 N_A_114_112#_c_929_n N_VGND_c_1073_n 0.00842441f $X=0.89 $Y=0.625 $X2=0
+ $Y2=0
cc_571 N_A_114_112#_c_928_n N_VGND_c_1076_n 0.0242087f $X=2.125 $Y=0.625 $X2=0
+ $Y2=0
cc_572 N_A_114_112#_c_928_n N_VGND_c_1078_n 0.0288276f $X=2.125 $Y=0.625 $X2=0
+ $Y2=0
cc_573 N_A_114_112#_c_929_n N_VGND_c_1078_n 0.0111078f $X=0.89 $Y=0.625 $X2=0
+ $Y2=0
cc_574 N_A_114_112#_c_932_n N_VGND_c_1078_n 0.00897192f $X=2.29 $Y=0.53 $X2=0
+ $Y2=0
cc_575 N_GCLK_c_1025_n N_VGND_c_1066_n 0.0164982f $X=7.46 $Y=0.515 $X2=0 $Y2=0
cc_576 N_GCLK_c_1025_n N_VGND_c_1068_n 0.0293763f $X=7.46 $Y=0.515 $X2=0 $Y2=0
cc_577 N_GCLK_c_1025_n N_VGND_c_1075_n 0.0144922f $X=7.46 $Y=0.515 $X2=0 $Y2=0
cc_578 N_GCLK_c_1025_n N_VGND_c_1078_n 0.0118826f $X=7.46 $Y=0.515 $X2=0 $Y2=0

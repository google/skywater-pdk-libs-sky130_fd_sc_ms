# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__a2bb2o_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.264000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 1.350000 2.850000 1.780000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.264000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.360000 1.350000 3.685000 1.780000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 1.260000 7.075000 1.780000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.492000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405000 1.260000 6.115000 1.780000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.086400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.960000 2.045000 1.130000 ;
        RECT 0.125000 1.130000 0.835000 1.780000 ;
        RECT 0.665000 1.780000 0.835000 1.800000 ;
        RECT 0.665000 1.800000 2.240000 1.970000 ;
        RECT 0.935000 0.350000 1.185000 0.960000 ;
        RECT 1.010000 1.970000 1.340000 2.980000 ;
        RECT 1.795000 0.350000 2.045000 0.960000 ;
        RECT 1.910000 1.970000 2.240000 2.980000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.505000  0.085000 0.755000 0.790000 ;
      RECT 0.560000  2.140000 0.810000 3.245000 ;
      RECT 1.035000  1.300000 2.385000 1.630000 ;
      RECT 1.365000  0.085000 1.615000 0.790000 ;
      RECT 1.540000  2.140000 1.710000 3.245000 ;
      RECT 2.215000  1.010000 2.815000 1.180000 ;
      RECT 2.215000  1.180000 2.385000 1.300000 ;
      RECT 2.225000  0.085000 2.475000 0.840000 ;
      RECT 2.410000  1.950000 2.780000 3.245000 ;
      RECT 2.645000  0.255000 3.530000 0.425000 ;
      RECT 2.645000  0.425000 2.815000 1.010000 ;
      RECT 2.985000  0.595000 3.190000 1.130000 ;
      RECT 3.020000  1.130000 3.190000 1.950000 ;
      RECT 3.020000  1.950000 4.150000 2.120000 ;
      RECT 3.290000  2.120000 3.620000 2.980000 ;
      RECT 3.360000  0.425000 3.530000 1.010000 ;
      RECT 3.360000  1.010000 4.815000 1.180000 ;
      RECT 3.700000  0.085000 4.385000 0.840000 ;
      RECT 3.855000  1.470000 4.150000 1.950000 ;
      RECT 4.060000  2.290000 4.390000 2.905000 ;
      RECT 4.060000  2.905000 5.210000 3.075000 ;
      RECT 4.565000  0.350000 5.765000 0.600000 ;
      RECT 4.565000  0.600000 4.815000 1.010000 ;
      RECT 4.565000  1.180000 4.760000 2.735000 ;
      RECT 4.960000  1.950000 7.090000 2.120000 ;
      RECT 4.960000  2.120000 5.210000 2.905000 ;
      RECT 5.005000  0.770000 6.115000 0.920000 ;
      RECT 5.005000  0.920000 7.095000 1.090000 ;
      RECT 5.410000  2.290000 5.660000 3.245000 ;
      RECT 5.860000  2.120000 6.190000 2.980000 ;
      RECT 5.945000  0.350000 6.115000 0.770000 ;
      RECT 6.295000  0.350000 6.665000 0.750000 ;
      RECT 6.390000  2.290000 6.560000 3.245000 ;
      RECT 6.495000  0.085000 6.665000 0.350000 ;
      RECT 6.760000  2.120000 7.090000 2.980000 ;
      RECT 6.845000  0.350000 7.095000 0.920000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_ms__a2bb2o_4

* File: sky130_fd_sc_ms__a2111o_2.pex.spice
* Created: Wed Sep  2 11:49:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A2111O_2%A_91_244# 1 2 3 4 15 17 19 22 24 26 27 28
+ 29 31 32 33 35 39 41 45 47 51 56 59 60
c116 60 0 1.10806e-19 $X=2.885 $Y=1.095
c117 27 0 1.60145e-19 $X=1.275 $Y=1.55
r118 64 65 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=0.99 $Y=1.385
+ $X2=0.995 $Y2=1.385
r119 63 64 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.56 $Y=1.385
+ $X2=0.99 $Y2=1.385
r120 61 63 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.545 $Y=1.385
+ $X2=0.56 $Y2=1.385
r121 56 65 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=1.195 $Y=1.385
+ $X2=0.995 $Y2=1.385
r122 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.195
+ $Y=1.385 $X2=1.195 $Y2=1.385
r123 53 55 13.2509 $w=2.67e-07 $l=2.9e-07 $layer=LI1_cond $X=1.195 $Y=1.095
+ $X2=1.195 $Y2=1.385
r124 49 51 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.355 $Y=1.01
+ $X2=4.355 $Y2=0.515
r125 48 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.01 $Y=1.095
+ $X2=2.885 $Y2=1.095
r126 47 49 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.19 $Y=1.095
+ $X2=4.355 $Y2=1.01
r127 47 48 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=4.19 $Y=1.095
+ $X2=3.01 $Y2=1.095
r128 43 60 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.885 $Y=1.01
+ $X2=2.885 $Y2=1.095
r129 43 45 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=2.885 $Y=1.01
+ $X2=2.885 $Y2=0.515
r130 42 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.03 $Y=1.095
+ $X2=1.905 $Y2=1.095
r131 41 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.76 $Y=1.095
+ $X2=2.885 $Y2=1.095
r132 41 42 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.76 $Y=1.095
+ $X2=2.03 $Y2=1.095
r133 37 59 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.905 $Y=1.01
+ $X2=1.905 $Y2=1.095
r134 37 39 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.905 $Y=1.01
+ $X2=1.905 $Y2=0.515
r135 33 58 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.92 $Y=2.12 $X2=1.92
+ $Y2=2.035
r136 33 35 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.92 $Y=2.12
+ $X2=1.92 $Y2=2.815
r137 31 58 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.755 $Y=2.035
+ $X2=1.92 $Y2=2.035
r138 31 32 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.755 $Y=2.035
+ $X2=1.36 $Y2=2.035
r139 30 53 3.37873 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.36 $Y=1.095
+ $X2=1.195 $Y2=1.095
r140 29 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.78 $Y=1.095
+ $X2=1.905 $Y2=1.095
r141 29 30 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.78 $Y=1.095
+ $X2=1.36 $Y2=1.095
r142 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.275 $Y=1.95
+ $X2=1.36 $Y2=2.035
r143 27 55 9.14344 $w=2.67e-07 $l=2.0106e-07 $layer=LI1_cond $X=1.275 $Y=1.55
+ $X2=1.195 $Y2=1.385
r144 27 28 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.275 $Y=1.55
+ $X2=1.275 $Y2=1.95
r145 24 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=1.22
+ $X2=0.99 $Y2=1.385
r146 24 26 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.99 $Y=1.22
+ $X2=0.99 $Y2=0.74
r147 20 65 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.55
+ $X2=0.995 $Y2=1.385
r148 20 22 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.995 $Y=1.55
+ $X2=0.995 $Y2=2.4
r149 17 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.56 $Y=1.22
+ $X2=0.56 $Y2=1.385
r150 17 19 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.56 $Y=1.22
+ $X2=0.56 $Y2=0.74
r151 13 61 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.55
+ $X2=0.545 $Y2=1.385
r152 13 15 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.545 $Y=1.55
+ $X2=0.545 $Y2=2.4
r153 4 58 400 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=1.795
+ $Y=1.84 $X2=1.92 $Y2=2.115
r154 4 35 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=1.795
+ $Y=1.84 $X2=1.92 $Y2=2.815
r155 3 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.215
+ $Y=0.37 $X2=4.355 $Y2=0.515
r156 2 45 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.705
+ $Y=0.37 $X2=2.845 $Y2=0.515
r157 1 39 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.82
+ $Y=0.37 $X2=1.945 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A2111O_2%D1 3 7 9 10 14
c37 14 0 1.60145e-19 $X=2.07 $Y=1.515
r38 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.07 $Y=1.515
+ $X2=2.07 $Y2=1.68
r39 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.07 $Y=1.515
+ $X2=2.07 $Y2=1.35
r40 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.07
+ $Y=1.515 $X2=2.07 $Y2=1.515
r41 10 15 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=2.16 $Y=1.565 $X2=2.07
+ $Y2=1.565
r42 9 15 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=2.07 $Y2=1.565
r43 7 16 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.16 $Y=0.74 $X2=2.16
+ $Y2=1.35
r44 3 17 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.145 $Y=2.4
+ $X2=2.145 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__A2111O_2%C1 3 7 9 10 11 12 18 19
c40 18 0 1.10806e-19 $X=2.61 $Y=1.515
c41 3 0 2.48122e-19 $X=2.535 $Y=2.4
r42 18 21 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.61 $Y=1.515
+ $X2=2.61 $Y2=1.68
r43 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.61 $Y=1.515
+ $X2=2.61 $Y2=1.35
r44 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.515 $X2=2.61 $Y2=1.515
r45 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.61 $Y=2.405
+ $X2=2.61 $Y2=2.775
r46 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.61 $Y=2.035
+ $X2=2.61 $Y2=2.405
r47 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=2.035
r48 9 19 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=1.515
r49 7 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.63 $Y=0.74 $X2=2.63
+ $Y2=1.35
r50 3 21 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.535 $Y=2.4
+ $X2=2.535 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__A2111O_2%B1 3 7 9 12 13
c38 13 0 1.02106e-19 $X=3.15 $Y=1.515
r39 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=1.515
+ $X2=3.15 $Y2=1.68
r40 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=1.515
+ $X2=3.15 $Y2=1.35
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.15
+ $Y=1.515 $X2=3.15 $Y2=1.515
r42 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.15 $Y=1.665
+ $X2=3.15 $Y2=1.515
r43 7 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.075 $Y=2.4
+ $X2=3.075 $Y2=1.68
r44 3 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.06 $Y=0.74 $X2=3.06
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__A2111O_2%A2 3 7 9 10 14
c36 14 0 1.56668e-19 $X=3.69 $Y=1.515
r37 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.69 $Y=1.515
+ $X2=3.69 $Y2=1.68
r38 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.69 $Y=1.515
+ $X2=3.69 $Y2=1.35
r39 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.69
+ $Y=1.515 $X2=3.69 $Y2=1.515
r40 10 15 10.4524 $w=4.28e-07 $l=3.9e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=3.69 $Y2=1.565
r41 9 15 2.41209 $w=4.28e-07 $l=9e-08 $layer=LI1_cond $X=3.6 $Y=1.565 $X2=3.69
+ $Y2=1.565
r42 7 16 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.78 $Y=0.74 $X2=3.78
+ $Y2=1.35
r43 3 17 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.615 $Y=2.4
+ $X2=3.615 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__A2111O_2%A1 3 7 10 11 14 15
c30 15 0 1.56668e-19 $X=4.53 $Y=1.515
r31 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.53
+ $Y=1.515 $X2=4.53 $Y2=1.515
r32 11 15 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.53 $Y=1.665
+ $X2=4.53 $Y2=1.515
r33 9 14 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=4.245 $Y=1.515
+ $X2=4.53 $Y2=1.515
r34 9 10 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.245 $Y=1.515
+ $X2=4.155 $Y2=1.515
r35 5 10 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=4.155 $Y=1.68
+ $X2=4.155 $Y2=1.515
r36 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.155 $Y=1.68
+ $X2=4.155 $Y2=2.4
r37 1 10 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=4.14 $Y=1.35
+ $X2=4.155 $Y2=1.515
r38 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.14 $Y=1.35 $X2=4.14
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A2111O_2%VPWR 1 2 3 10 12 18 22 25 26 27 29 42 43 49
r53 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r54 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r55 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r56 40 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r57 39 40 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r58 37 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r59 36 39 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r60 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r61 34 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=3.33
+ $X2=1.22 $Y2=3.33
r62 34 36 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 33 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r64 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r65 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r66 30 46 3.96192 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=3.33
+ $X2=0.202 $Y2=3.33
r67 30 32 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.405 $Y=3.33
+ $X2=0.72 $Y2=3.33
r68 29 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.22 $Y2=3.33
r69 29 32 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.72 $Y2=3.33
r70 27 40 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=3.6
+ $Y2=3.33
r71 27 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=1.68 $Y2=3.33
r72 25 39 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.675 $Y=3.33
+ $X2=3.6 $Y2=3.33
r73 25 26 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.675 $Y=3.33
+ $X2=3.86 $Y2=3.33
r74 24 42 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=4.56 $Y2=3.33
r75 24 26 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=3.86 $Y2=3.33
r76 20 26 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.86 $Y=3.245
+ $X2=3.86 $Y2=3.33
r77 20 22 24.6062 $w=3.68e-07 $l=7.9e-07 $layer=LI1_cond $X=3.86 $Y=3.245
+ $X2=3.86 $Y2=2.455
r78 16 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=3.245
+ $X2=1.22 $Y2=3.33
r79 16 18 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.22 $Y=3.245
+ $X2=1.22 $Y2=2.455
r80 12 15 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r81 10 46 3.18124 $w=2.5e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.202 $Y2=3.33
r82 10 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r83 3 22 300 $w=1.7e-07 $l=6.8815e-07 $layer=licon1_PDIFF $count=2 $X=3.705
+ $Y=1.84 $X2=3.86 $Y2=2.455
r84 2 18 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=1.84 $X2=1.22 $Y2=2.455
r85 1 15 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.84 $X2=0.32 $Y2=2.815
r86 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.84 $X2=0.32 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__A2111O_2%X 1 2 9 11 12 13 14 34
c19 11 0 1.2388e-19 $X=0.635 $Y=1.58
r20 20 34 0.542326 $w=2.53e-07 $l=1.2e-08 $layer=LI1_cond $X=0.732 $Y=1.677
+ $X2=0.732 $Y2=1.665
r21 13 14 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.732 $Y=2.405
+ $X2=0.732 $Y2=2.775
r22 12 13 18.9814 $w=2.53e-07 $l=4.2e-07 $layer=LI1_cond $X=0.732 $Y=1.985
+ $X2=0.732 $Y2=2.405
r23 11 34 1.67217 $w=2.53e-07 $l=3.7e-08 $layer=LI1_cond $X=0.732 $Y=1.628
+ $X2=0.732 $Y2=1.665
r24 11 32 4.80861 $w=2.53e-07 $l=7.8e-08 $layer=LI1_cond $X=0.732 $Y=1.628
+ $X2=0.732 $Y2=1.55
r25 11 12 12.2927 $w=2.53e-07 $l=2.72e-07 $layer=LI1_cond $X=0.732 $Y=1.713
+ $X2=0.732 $Y2=1.985
r26 11 20 1.62698 $w=2.53e-07 $l=3.6e-08 $layer=LI1_cond $X=0.732 $Y=1.713
+ $X2=0.732 $Y2=1.677
r27 9 32 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=0.775 $Y=0.515
+ $X2=0.775 $Y2=1.55
r28 2 14 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.635
+ $Y=1.84 $X2=0.77 $Y2=2.815
r29 2 12 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.635
+ $Y=1.84 $X2=0.77 $Y2=1.985
r30 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.635
+ $Y=0.37 $X2=0.775 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A2111O_2%A_633_368# 1 2 7 9 11 13 15
c28 7 0 1.46017e-19 $X=3.32 $Y=2.12
r29 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.38 $Y=2.12 $X2=4.38
+ $Y2=2.035
r30 13 15 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.38 $Y=2.12
+ $X2=4.38 $Y2=2.815
r31 12 18 5.55669 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.505 $Y=2.035
+ $X2=3.32 $Y2=2.035
r32 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.215 $Y=2.035
+ $X2=4.38 $Y2=2.035
r33 11 12 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.215 $Y=2.035
+ $X2=3.505 $Y2=2.035
r34 7 18 2.55307 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.32 $Y=2.12 $X2=3.32
+ $Y2=2.035
r35 7 9 21.6472 $w=3.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.32 $Y=2.12 $X2=3.32
+ $Y2=2.815
r36 2 20 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=4.245
+ $Y=1.84 $X2=4.38 $Y2=2.115
r37 2 15 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.245
+ $Y=1.84 $X2=4.38 $Y2=2.815
r38 1 18 400 $w=1.7e-07 $l=3.43875e-07 $layer=licon1_PDIFF $count=1 $X=3.165
+ $Y=1.84 $X2=3.32 $Y2=2.115
r39 1 9 400 $w=1.7e-07 $l=1.04964e-06 $layer=licon1_PDIFF $count=1 $X=3.165
+ $Y=1.84 $X2=3.32 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__A2111O_2%VGND 1 2 3 4 13 15 19 23 27 30 31 32 34 43
+ 49 50 56 59
r61 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r62 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r63 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r64 50 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r65 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r66 47 59 11.9488 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=3.73 $Y=0 $X2=3.455
+ $Y2=0
r67 47 49 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.73 $Y=0 $X2=4.56
+ $Y2=0
r68 46 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r69 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r70 43 59 11.9488 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=3.18 $Y=0 $X2=3.455
+ $Y2=0
r71 43 45 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.18 $Y=0 $X2=3.12
+ $Y2=0
r72 42 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r73 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r74 39 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.37 $Y=0 $X2=1.205
+ $Y2=0
r75 39 41 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.37 $Y=0 $X2=2.16
+ $Y2=0
r76 38 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r77 38 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r78 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r79 35 53 4.60552 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.51 $Y=0 $X2=0.255
+ $Y2=0
r80 35 37 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.51 $Y=0 $X2=0.72
+ $Y2=0
r81 34 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.04 $Y=0 $X2=1.205
+ $Y2=0
r82 34 37 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.04 $Y=0 $X2=0.72
+ $Y2=0
r83 32 46 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r84 32 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r85 30 41 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.16
+ $Y2=0
r86 30 31 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.21 $Y=0 $X2=2.395
+ $Y2=0
r87 29 45 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.58 $Y=0 $X2=3.12
+ $Y2=0
r88 29 31 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.58 $Y=0 $X2=2.395
+ $Y2=0
r89 25 59 2.31338 $w=5.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.455 $Y=0.085
+ $X2=3.455 $Y2=0
r90 25 27 12.8307 $w=5.48e-07 $l=5.9e-07 $layer=LI1_cond $X=3.455 $Y=0.085
+ $X2=3.455 $Y2=0.675
r91 21 31 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.395 $Y=0.085
+ $X2=2.395 $Y2=0
r92 21 23 18.3768 $w=3.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.395 $Y=0.085
+ $X2=2.395 $Y2=0.675
r93 17 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0.085
+ $X2=1.205 $Y2=0
r94 17 19 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.205 $Y=0.085
+ $X2=1.205 $Y2=0.675
r95 13 53 3.16065 $w=3.3e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.345 $Y=0.085
+ $X2=0.255 $Y2=0
r96 13 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.345 $Y=0.085
+ $X2=0.345 $Y2=0.515
r97 4 27 182 $w=1.7e-07 $l=4.36635e-07 $layer=licon1_NDIFF $count=1 $X=3.135
+ $Y=0.37 $X2=3.445 $Y2=0.675
r98 3 23 182 $w=1.7e-07 $l=3.76597e-07 $layer=licon1_NDIFF $count=1 $X=2.235
+ $Y=0.37 $X2=2.395 $Y2=0.675
r99 2 19 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.37 $X2=1.205 $Y2=0.675
r100 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.22
+ $Y=0.37 $X2=0.345 $Y2=0.515
.ends


* File: sky130_fd_sc_ms__nor3_2.pxi.spice
* Created: Wed Sep  2 12:16:04 2020
* 
x_PM_SKY130_FD_SC_MS__NOR3_2%C N_C_c_59_n N_C_M1000_g N_C_c_56_n N_C_M1006_g
+ N_C_c_60_n N_C_M1002_g C N_C_c_58_n PM_SKY130_FD_SC_MS__NOR3_2%C
x_PM_SKY130_FD_SC_MS__NOR3_2%B N_B_M1001_g N_B_M1008_g N_B_c_95_n N_B_M1004_g
+ N_B_c_96_n N_B_c_97_n N_B_c_98_n B N_B_c_100_n PM_SKY130_FD_SC_MS__NOR3_2%B
x_PM_SKY130_FD_SC_MS__NOR3_2%A N_A_M1003_g N_A_c_158_n N_A_M1007_g N_A_c_159_n
+ N_A_M1005_g N_A_c_161_n N_A_c_162_n N_A_c_163_n N_A_c_164_n A N_A_c_166_n
+ PM_SKY130_FD_SC_MS__NOR3_2%A
x_PM_SKY130_FD_SC_MS__NOR3_2%A_27_368# N_A_27_368#_M1000_d N_A_27_368#_M1002_d
+ N_A_27_368#_M1004_s N_A_27_368#_c_215_n N_A_27_368#_c_216_n
+ N_A_27_368#_c_217_n N_A_27_368#_c_218_n N_A_27_368#_c_219_n
+ N_A_27_368#_c_220_n PM_SKY130_FD_SC_MS__NOR3_2%A_27_368#
x_PM_SKY130_FD_SC_MS__NOR3_2%Y N_Y_M1006_s N_Y_M1008_d N_Y_M1000_s N_Y_c_262_n
+ N_Y_c_269_n N_Y_c_272_n N_Y_c_258_n Y Y Y Y N_Y_c_264_n Y
+ PM_SKY130_FD_SC_MS__NOR3_2%Y
x_PM_SKY130_FD_SC_MS__NOR3_2%A_309_368# N_A_309_368#_M1001_d
+ N_A_309_368#_M1005_d N_A_309_368#_c_304_n N_A_309_368#_c_302_n
+ N_A_309_368#_c_309_n N_A_309_368#_c_306_n N_A_309_368#_c_303_n
+ PM_SKY130_FD_SC_MS__NOR3_2%A_309_368#
x_PM_SKY130_FD_SC_MS__NOR3_2%VPWR N_VPWR_M1003_s N_VPWR_c_328_n VPWR
+ N_VPWR_c_329_n N_VPWR_c_330_n N_VPWR_c_327_n N_VPWR_c_332_n
+ PM_SKY130_FD_SC_MS__NOR3_2%VPWR
x_PM_SKY130_FD_SC_MS__NOR3_2%VGND N_VGND_M1006_d N_VGND_M1007_d N_VGND_c_364_n
+ N_VGND_c_365_n VGND N_VGND_c_366_n N_VGND_c_367_n N_VGND_c_368_n
+ N_VGND_c_369_n N_VGND_c_370_n PM_SKY130_FD_SC_MS__NOR3_2%VGND
cc_1 VNB N_C_c_56_n 0.0238316f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_2 VNB C 0.0064001f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_C_c_58_n 0.0618864f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=1.385
cc_4 VNB N_B_M1001_g 0.00632357f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_5 VNB N_B_c_95_n 0.0638178f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_6 VNB N_B_c_96_n 0.0196703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_B_c_97_n 0.00315176f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=1.49
cc_8 VNB N_B_c_98_n 0.0307722f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=1.385
cc_9 VNB B 0.00742405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B_c_100_n 0.0218521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_M1003_g 0.0159305f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_12 VNB N_A_c_158_n 0.0171724f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_13 VNB N_A_c_159_n 0.00880223f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.4
cc_14 VNB N_A_M1005_g 0.0176973f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_15 VNB N_A_c_161_n 0.0171751f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=1.385
cc_16 VNB N_A_c_162_n 0.00955942f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=1.385
cc_17 VNB N_A_c_163_n 0.0169275f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.295
cc_18 VNB N_A_c_164_n 0.029959f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.385
cc_19 VNB A 0.0323167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_c_166_n 0.0558262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_258_n 0.00280505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB Y 0.0212531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB Y 0.00704942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB Y 0.033575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_327_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.385
cc_26 VNB N_VGND_c_364_n 0.0185359f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.76
cc_27 VNB N_VGND_c_365_n 0.0188688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_366_n 0.0252139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_367_n 0.206462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_368_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_369_n 0.0280581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_370_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VPB N_C_c_59_n 0.0193495f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.76
cc_34 VPB N_C_c_60_n 0.0164225f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.76
cc_35 VPB N_C_c_58_n 0.0157671f $X=-0.19 $Y=1.66 $X2=0.81 $Y2=1.385
cc_36 VPB N_B_M1001_g 0.0223633f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_37 VPB N_B_c_95_n 0.0335044f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_38 VPB N_A_M1003_g 0.0218496f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_39 VPB N_A_M1005_g 0.0214006f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_40 VPB N_A_27_368#_c_215_n 0.0322259f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.22
cc_41 VPB N_A_27_368#_c_216_n 0.00512891f $X=-0.19 $Y=1.66 $X2=0.81 $Y2=1.385
cc_42 VPB N_A_27_368#_c_217_n 0.00965139f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=1.49
cc_43 VPB N_A_27_368#_c_218_n 0.0151346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A_27_368#_c_219_n 0.00751347f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A_27_368#_c_220_n 0.0432118f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_Y_c_262_n 0.00202686f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_47 VPB Y 0.00293411f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_Y_c_264_n 0.00767133f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_309_368#_c_302_n 0.00281193f $X=-0.19 $Y=1.66 $X2=1.005 $Y2=2.4
cc_50 VPB N_A_309_368#_c_303_n 0.00233516f $X=-0.19 $Y=1.66 $X2=0.81 $Y2=1.385
cc_51 VPB N_VPWR_c_328_n 0.00396467f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_52 VPB N_VPWR_c_329_n 0.0518789f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_53 VPB N_VPWR_c_330_n 0.0298982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_327_n 0.0613443f $X=-0.19 $Y=1.66 $X2=0.79 $Y2=1.385
cc_55 VPB N_VPWR_c_332_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 N_C_c_58_n N_B_M1001_g 0.0230263f $X=0.81 $Y=1.385 $X2=0 $Y2=0
cc_57 C N_B_c_97_n 0.0146852f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_58 N_C_c_58_n N_B_c_97_n 0.00140882f $X=0.81 $Y=1.385 $X2=0 $Y2=0
cc_59 C N_B_c_98_n 9.60045e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_60 N_C_c_58_n N_B_c_98_n 0.0216281f $X=0.81 $Y=1.385 $X2=0 $Y2=0
cc_61 C N_B_c_100_n 0.00107469f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_62 N_C_c_59_n N_A_27_368#_c_215_n 0.0112976f $X=0.505 $Y=1.76 $X2=0 $Y2=0
cc_63 N_C_c_60_n N_A_27_368#_c_215_n 5.42618e-19 $X=1.005 $Y=1.76 $X2=0 $Y2=0
cc_64 N_C_c_59_n N_A_27_368#_c_216_n 0.0119307f $X=0.505 $Y=1.76 $X2=0 $Y2=0
cc_65 N_C_c_60_n N_A_27_368#_c_216_n 0.0139536f $X=1.005 $Y=1.76 $X2=0 $Y2=0
cc_66 N_C_c_59_n N_A_27_368#_c_217_n 0.00291744f $X=0.505 $Y=1.76 $X2=0 $Y2=0
cc_67 N_C_c_58_n N_A_27_368#_c_219_n 0.00110907f $X=0.81 $Y=1.385 $X2=0 $Y2=0
cc_68 N_C_c_59_n N_Y_c_262_n 0.0128115f $X=0.505 $Y=1.76 $X2=0 $Y2=0
cc_69 N_C_c_60_n N_Y_c_262_n 0.00257327f $X=1.005 $Y=1.76 $X2=0 $Y2=0
cc_70 C N_Y_c_262_n 0.0274789f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_71 N_C_c_58_n N_Y_c_262_n 0.0151636f $X=0.81 $Y=1.385 $X2=0 $Y2=0
cc_72 N_C_c_56_n N_Y_c_269_n 0.0112f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_73 C N_Y_c_269_n 0.028324f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_74 N_C_c_58_n N_Y_c_269_n 0.00755208f $X=0.81 $Y=1.385 $X2=0 $Y2=0
cc_75 N_C_c_60_n N_Y_c_272_n 0.0104219f $X=1.005 $Y=1.76 $X2=0 $Y2=0
cc_76 N_C_c_56_n Y 0.0124397f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_77 N_C_c_56_n Y 8.87593e-19 $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_78 N_C_c_56_n Y 0.01042f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_79 C Y 0.0225409f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_80 N_C_c_58_n Y 0.0056331f $X=0.81 $Y=1.385 $X2=0 $Y2=0
cc_81 N_C_c_59_n N_VPWR_c_329_n 0.00333896f $X=0.505 $Y=1.76 $X2=0 $Y2=0
cc_82 N_C_c_60_n N_VPWR_c_329_n 0.00333926f $X=1.005 $Y=1.76 $X2=0 $Y2=0
cc_83 N_C_c_59_n N_VPWR_c_327_n 0.00426915f $X=0.505 $Y=1.76 $X2=0 $Y2=0
cc_84 N_C_c_60_n N_VPWR_c_327_n 0.00423286f $X=1.005 $Y=1.76 $X2=0 $Y2=0
cc_85 N_C_c_56_n N_VGND_c_367_n 0.00453471f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_86 N_C_c_56_n N_VGND_c_368_n 0.00434272f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_87 N_C_c_56_n N_VGND_c_369_n 0.0110054f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_88 N_B_M1001_g N_A_M1003_g 0.0231675f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_89 N_B_c_96_n N_A_M1003_g 0.0129333f $X=2.925 $Y=1.465 $X2=0 $Y2=0
cc_90 N_B_c_100_n N_A_c_158_n 0.0179489f $X=1.47 $Y=1.22 $X2=0 $Y2=0
cc_91 N_B_c_96_n N_A_c_159_n 0.00380862f $X=2.925 $Y=1.465 $X2=0 $Y2=0
cc_92 N_B_c_95_n N_A_M1005_g 0.0318297f $X=2.855 $Y=1.725 $X2=0 $Y2=0
cc_93 N_B_c_96_n N_A_M1005_g 0.0129019f $X=2.925 $Y=1.465 $X2=0 $Y2=0
cc_94 B N_A_M1005_g 3.6606e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_95 B N_A_c_161_n 0.00159669f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_96 N_B_c_97_n N_A_c_162_n 0.0011932f $X=1.47 $Y=1.385 $X2=0 $Y2=0
cc_97 N_B_c_98_n N_A_c_162_n 0.0221136f $X=1.47 $Y=1.385 $X2=0 $Y2=0
cc_98 N_B_c_100_n N_A_c_162_n 0.00228878f $X=1.47 $Y=1.22 $X2=0 $Y2=0
cc_99 N_B_c_95_n N_A_c_163_n 0.00713314f $X=2.855 $Y=1.725 $X2=0 $Y2=0
cc_100 N_B_c_96_n N_A_c_163_n 0.00855379f $X=2.925 $Y=1.465 $X2=0 $Y2=0
cc_101 B N_A_c_163_n 8.70735e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_102 N_B_c_95_n N_A_c_164_n 0.00551673f $X=2.855 $Y=1.725 $X2=0 $Y2=0
cc_103 N_B_c_96_n N_A_c_164_n 0.00317985f $X=2.925 $Y=1.465 $X2=0 $Y2=0
cc_104 B N_A_c_164_n 3.63484e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_105 N_B_c_95_n A 0.00183654f $X=2.855 $Y=1.725 $X2=0 $Y2=0
cc_106 N_B_c_96_n A 0.0114949f $X=2.925 $Y=1.465 $X2=0 $Y2=0
cc_107 B A 0.0242925f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_108 N_B_M1001_g N_A_27_368#_c_216_n 0.00297009f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_109 N_B_M1001_g N_A_27_368#_c_218_n 0.0154114f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_110 N_B_c_95_n N_A_27_368#_c_218_n 0.0220621f $X=2.855 $Y=1.725 $X2=0 $Y2=0
cc_111 N_B_c_96_n N_A_27_368#_c_218_n 0.093824f $X=2.925 $Y=1.465 $X2=0 $Y2=0
cc_112 N_B_c_97_n N_A_27_368#_c_218_n 0.0233821f $X=1.47 $Y=1.385 $X2=0 $Y2=0
cc_113 N_B_c_98_n N_A_27_368#_c_218_n 9.72046e-19 $X=1.47 $Y=1.385 $X2=0 $Y2=0
cc_114 B N_A_27_368#_c_218_n 0.0262111f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_115 N_B_c_97_n N_A_27_368#_c_219_n 7.62703e-19 $X=1.47 $Y=1.385 $X2=0 $Y2=0
cc_116 N_B_c_95_n N_A_27_368#_c_220_n 0.00151667f $X=2.855 $Y=1.725 $X2=0 $Y2=0
cc_117 N_B_c_96_n N_Y_c_269_n 0.0144587f $X=2.925 $Y=1.465 $X2=0 $Y2=0
cc_118 N_B_c_97_n N_Y_c_269_n 0.0176193f $X=1.47 $Y=1.385 $X2=0 $Y2=0
cc_119 N_B_c_98_n N_Y_c_269_n 8.56939e-19 $X=1.47 $Y=1.385 $X2=0 $Y2=0
cc_120 N_B_c_100_n N_Y_c_269_n 0.0142961f $X=1.47 $Y=1.22 $X2=0 $Y2=0
cc_121 N_B_c_100_n N_Y_c_258_n 0.00261686f $X=1.47 $Y=1.22 $X2=0 $Y2=0
cc_122 N_B_M1001_g N_A_309_368#_c_304_n 0.00244698f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_123 N_B_M1001_g N_A_309_368#_c_302_n 0.0095906f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_124 N_B_c_95_n N_A_309_368#_c_306_n 0.00242423f $X=2.855 $Y=1.725 $X2=0 $Y2=0
cc_125 N_B_c_95_n N_A_309_368#_c_303_n 0.00977276f $X=2.855 $Y=1.725 $X2=0 $Y2=0
cc_126 N_B_M1001_g N_VPWR_c_328_n 6.19643e-19 $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_127 N_B_c_95_n N_VPWR_c_328_n 6.62524e-19 $X=2.855 $Y=1.725 $X2=0 $Y2=0
cc_128 N_B_M1001_g N_VPWR_c_329_n 0.00520636f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_129 N_B_c_95_n N_VPWR_c_330_n 0.00520636f $X=2.855 $Y=1.725 $X2=0 $Y2=0
cc_130 N_B_M1001_g N_VPWR_c_327_n 0.00983669f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_131 N_B_c_95_n N_VPWR_c_327_n 0.00987022f $X=2.855 $Y=1.725 $X2=0 $Y2=0
cc_132 N_B_c_100_n N_VGND_c_364_n 0.00383152f $X=1.47 $Y=1.22 $X2=0 $Y2=0
cc_133 N_B_c_96_n N_VGND_c_365_n 0.0204916f $X=2.925 $Y=1.465 $X2=0 $Y2=0
cc_134 N_B_c_100_n N_VGND_c_367_n 0.00383029f $X=1.47 $Y=1.22 $X2=0 $Y2=0
cc_135 N_B_c_100_n N_VGND_c_369_n 0.00924883f $X=1.47 $Y=1.22 $X2=0 $Y2=0
cc_136 N_A_M1003_g N_A_27_368#_c_218_n 0.0119241f $X=1.935 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A_M1005_g N_A_27_368#_c_218_n 0.0117481f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_138 N_A_c_158_n N_Y_c_269_n 0.00265815f $X=2.03 $Y=1.185 $X2=0 $Y2=0
cc_139 N_A_c_162_n N_Y_c_269_n 0.00307701f $X=1.975 $Y=1.26 $X2=0 $Y2=0
cc_140 N_A_c_158_n N_Y_c_258_n 0.0055158f $X=2.03 $Y=1.185 $X2=0 $Y2=0
cc_141 N_A_M1003_g N_A_309_368#_c_302_n 2.57325e-19 $X=1.935 $Y=2.4 $X2=0 $Y2=0
cc_142 N_A_M1003_g N_A_309_368#_c_309_n 0.0149911f $X=1.935 $Y=2.4 $X2=0 $Y2=0
cc_143 N_A_M1005_g N_A_309_368#_c_309_n 0.0143795f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A_M1005_g N_A_309_368#_c_303_n 2.34582e-19 $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_145 N_A_M1003_g N_VPWR_c_328_n 0.00951846f $X=1.935 $Y=2.4 $X2=0 $Y2=0
cc_146 N_A_M1005_g N_VPWR_c_328_n 0.0111228f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_147 N_A_M1003_g N_VPWR_c_329_n 0.00521592f $X=1.935 $Y=2.4 $X2=0 $Y2=0
cc_148 N_A_M1005_g N_VPWR_c_330_n 0.00460063f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_149 N_A_M1003_g N_VPWR_c_327_n 0.0102937f $X=1.935 $Y=2.4 $X2=0 $Y2=0
cc_150 N_A_M1005_g N_VPWR_c_327_n 0.00908665f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_151 N_A_c_158_n N_VGND_c_364_n 0.00434272f $X=2.03 $Y=1.185 $X2=0 $Y2=0
cc_152 N_A_c_158_n N_VGND_c_365_n 0.0080629f $X=2.03 $Y=1.185 $X2=0 $Y2=0
cc_153 N_A_c_159_n N_VGND_c_365_n 0.00795019f $X=2.315 $Y=1.26 $X2=0 $Y2=0
cc_154 A N_VGND_c_365_n 0.0553698f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_155 N_A_c_166_n N_VGND_c_365_n 0.0117383f $X=2.815 $Y=0.475 $X2=0 $Y2=0
cc_156 A N_VGND_c_366_n 0.0298314f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_157 N_A_c_166_n N_VGND_c_366_n 0.0120882f $X=2.815 $Y=0.475 $X2=0 $Y2=0
cc_158 N_A_c_158_n N_VGND_c_367_n 0.00825771f $X=2.03 $Y=1.185 $X2=0 $Y2=0
cc_159 A N_VGND_c_367_n 0.0218461f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_160 N_A_c_166_n N_VGND_c_367_n 0.0154157f $X=2.815 $Y=0.475 $X2=0 $Y2=0
cc_161 N_A_c_158_n N_VGND_c_369_n 4.24281e-19 $X=2.03 $Y=1.185 $X2=0 $Y2=0
cc_162 N_A_27_368#_c_216_n N_Y_M1000_s 0.00218982f $X=1.145 $Y=2.99 $X2=0 $Y2=0
cc_163 N_A_27_368#_c_215_n N_Y_c_262_n 0.0023016f $X=0.28 $Y=2.145 $X2=0 $Y2=0
cc_164 N_A_27_368#_c_219_n N_Y_c_262_n 0.0112335f $X=1.315 $Y=1.805 $X2=0 $Y2=0
cc_165 N_A_27_368#_c_216_n N_Y_c_272_n 0.0177084f $X=1.145 $Y=2.99 $X2=0 $Y2=0
cc_166 N_A_27_368#_M1000_d N_Y_c_264_n 0.00271132f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_167 N_A_27_368#_c_215_n N_Y_c_264_n 0.0216158f $X=0.28 $Y=2.145 $X2=0 $Y2=0
cc_168 N_A_27_368#_c_218_n N_A_309_368#_M1001_d 0.00197722f $X=2.965 $Y=1.805
+ $X2=-0.19 $Y2=1.66
cc_169 N_A_27_368#_c_218_n N_A_309_368#_M1005_d 0.00165831f $X=2.965 $Y=1.805
+ $X2=0 $Y2=0
cc_170 N_A_27_368#_c_218_n N_A_309_368#_c_304_n 0.0173758f $X=2.965 $Y=1.805
+ $X2=0 $Y2=0
cc_171 N_A_27_368#_c_216_n N_A_309_368#_c_302_n 0.00401662f $X=1.145 $Y=2.99
+ $X2=0 $Y2=0
cc_172 N_A_27_368#_c_218_n N_A_309_368#_c_309_n 0.0371166f $X=2.965 $Y=1.805
+ $X2=0 $Y2=0
cc_173 N_A_27_368#_c_218_n N_A_309_368#_c_306_n 0.0149351f $X=2.965 $Y=1.805
+ $X2=0 $Y2=0
cc_174 N_A_27_368#_c_220_n N_A_309_368#_c_303_n 0.0281768f $X=3.08 $Y=1.985
+ $X2=0 $Y2=0
cc_175 N_A_27_368#_c_218_n N_VPWR_M1003_s 0.00187547f $X=2.965 $Y=1.805
+ $X2=-0.19 $Y2=1.66
cc_176 N_A_27_368#_c_216_n N_VPWR_c_329_n 0.0562636f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_177 N_A_27_368#_c_217_n N_VPWR_c_329_n 0.023515f $X=0.445 $Y=2.99 $X2=0 $Y2=0
cc_178 N_A_27_368#_c_220_n N_VPWR_c_330_n 0.0124046f $X=3.08 $Y=1.985 $X2=0
+ $Y2=0
cc_179 N_A_27_368#_c_216_n N_VPWR_c_327_n 0.0314185f $X=1.145 $Y=2.99 $X2=0
+ $Y2=0
cc_180 N_A_27_368#_c_217_n N_VPWR_c_327_n 0.0126871f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_181 N_A_27_368#_c_220_n N_VPWR_c_327_n 0.0102675f $X=3.08 $Y=1.985 $X2=0
+ $Y2=0
cc_182 N_Y_c_269_n N_VGND_M1006_d 0.0266486f $X=1.65 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_183 N_Y_c_258_n N_VGND_c_364_n 0.0145947f $X=1.815 $Y=0.515 $X2=0 $Y2=0
cc_184 N_Y_c_258_n N_VGND_c_365_n 0.0191389f $X=1.815 $Y=0.515 $X2=0 $Y2=0
cc_185 N_Y_c_269_n N_VGND_c_367_n 0.0128359f $X=1.65 $Y=0.925 $X2=0 $Y2=0
cc_186 N_Y_c_258_n N_VGND_c_367_n 0.0120104f $X=1.815 $Y=0.515 $X2=0 $Y2=0
cc_187 Y N_VGND_c_367_n 0.011995f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_188 Y N_VGND_c_368_n 0.0145556f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_189 N_Y_c_269_n N_VGND_c_369_n 0.0573941f $X=1.65 $Y=0.925 $X2=0 $Y2=0
cc_190 N_Y_c_258_n N_VGND_c_369_n 0.0133889f $X=1.815 $Y=0.515 $X2=0 $Y2=0
cc_191 Y N_VGND_c_369_n 0.0121582f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_192 N_A_309_368#_c_309_n N_VPWR_M1003_s 0.00374639f $X=2.515 $Y=2.145
+ $X2=-0.19 $Y2=1.66
cc_193 N_A_309_368#_c_302_n N_VPWR_c_328_n 0.0466429f $X=1.68 $Y=2.825 $X2=0
+ $Y2=0
cc_194 N_A_309_368#_c_309_n N_VPWR_c_328_n 0.0171295f $X=2.515 $Y=2.145 $X2=0
+ $Y2=0
cc_195 N_A_309_368#_c_303_n N_VPWR_c_328_n 0.0233151f $X=2.63 $Y=2.485 $X2=0
+ $Y2=0
cc_196 N_A_309_368#_c_302_n N_VPWR_c_329_n 0.0151586f $X=1.68 $Y=2.825 $X2=0
+ $Y2=0
cc_197 N_A_309_368#_c_303_n N_VPWR_c_330_n 0.0128344f $X=2.63 $Y=2.485 $X2=0
+ $Y2=0
cc_198 N_A_309_368#_c_302_n N_VPWR_c_327_n 0.0120472f $X=1.68 $Y=2.825 $X2=0
+ $Y2=0
cc_199 N_A_309_368#_c_303_n N_VPWR_c_327_n 0.0101895f $X=2.63 $Y=2.485 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__nor2b_4.pxi.spice
* Created: Wed Sep  2 12:15:51 2020
* 
x_PM_SKY130_FD_SC_MS__NOR2B_4%A N_A_M1004_g N_A_M1005_g N_A_M1007_g N_A_c_80_n
+ N_A_M1003_g N_A_M1012_g N_A_c_82_n N_A_M1008_g N_A_c_83_n N_A_c_84_n
+ N_A_c_85_n N_A_c_86_n A A N_A_c_87_n PM_SKY130_FD_SC_MS__NOR2B_4%A
x_PM_SKY130_FD_SC_MS__NOR2B_4%A_353_323# N_A_353_323#_M1001_d
+ N_A_353_323#_M1000_d N_A_353_323#_c_185_n N_A_353_323#_M1009_g
+ N_A_353_323#_c_180_n N_A_353_323#_M1006_g N_A_353_323#_c_186_n
+ N_A_353_323#_M1010_g N_A_353_323#_c_181_n N_A_353_323#_M1014_g
+ N_A_353_323#_c_187_n N_A_353_323#_M1011_g N_A_353_323#_c_188_n
+ N_A_353_323#_M1013_g N_A_353_323#_c_189_n N_A_353_323#_c_190_n
+ N_A_353_323#_c_191_n N_A_353_323#_c_182_n N_A_353_323#_c_183_n
+ N_A_353_323#_c_184_n PM_SKY130_FD_SC_MS__NOR2B_4%A_353_323#
x_PM_SKY130_FD_SC_MS__NOR2B_4%B_N N_B_N_c_285_n N_B_N_M1000_g N_B_N_M1001_g
+ N_B_N_c_286_n N_B_N_M1002_g B_N B_N N_B_N_c_284_n
+ PM_SKY130_FD_SC_MS__NOR2B_4%B_N
x_PM_SKY130_FD_SC_MS__NOR2B_4%VPWR N_VPWR_M1004_s N_VPWR_M1005_s N_VPWR_M1012_s
+ N_VPWR_M1002_s N_VPWR_c_317_n N_VPWR_c_318_n N_VPWR_c_319_n N_VPWR_c_320_n
+ N_VPWR_c_321_n N_VPWR_c_322_n N_VPWR_c_323_n N_VPWR_c_324_n VPWR
+ N_VPWR_c_325_n N_VPWR_c_326_n N_VPWR_c_327_n N_VPWR_c_316_n
+ PM_SKY130_FD_SC_MS__NOR2B_4%VPWR
x_PM_SKY130_FD_SC_MS__NOR2B_4%A_119_368# N_A_119_368#_M1004_d
+ N_A_119_368#_M1007_d N_A_119_368#_M1010_s N_A_119_368#_M1013_s
+ N_A_119_368#_c_386_n N_A_119_368#_c_381_n N_A_119_368#_c_391_n
+ N_A_119_368#_c_393_n N_A_119_368#_c_394_n N_A_119_368#_c_382_n
+ N_A_119_368#_c_383_n N_A_119_368#_c_402_n N_A_119_368#_c_384_n
+ N_A_119_368#_c_398_n N_A_119_368#_c_385_n
+ PM_SKY130_FD_SC_MS__NOR2B_4%A_119_368#
x_PM_SKY130_FD_SC_MS__NOR2B_4%Y N_Y_M1006_d N_Y_M1003_d N_Y_M1009_d N_Y_M1011_d
+ N_Y_c_438_n N_Y_c_439_n N_Y_c_440_n N_Y_c_481_n N_Y_c_482_n N_Y_c_460_n
+ N_Y_c_487_n N_Y_c_490_n N_Y_c_441_n N_Y_c_442_n N_Y_c_443_n N_Y_c_492_n
+ N_Y_c_468_n Y Y Y PM_SKY130_FD_SC_MS__NOR2B_4%Y
x_PM_SKY130_FD_SC_MS__NOR2B_4%VGND N_VGND_M1006_s N_VGND_M1014_s N_VGND_M1008_s
+ N_VGND_c_523_n N_VGND_c_524_n VGND N_VGND_c_525_n N_VGND_c_526_n
+ N_VGND_c_527_n N_VGND_c_528_n N_VGND_c_529_n N_VGND_c_530_n N_VGND_c_531_n
+ N_VGND_c_532_n PM_SKY130_FD_SC_MS__NOR2B_4%VGND
cc_1 VNB N_A_M1004_g 0.0188384f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A_M1005_g 0.0162349f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_3 VNB N_A_M1007_g 0.0176514f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_4 VNB N_A_c_80_n 0.0193643f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=1.22
cc_5 VNB N_A_M1012_g 0.00737533f $X=-0.19 $Y=-0.245 $X2=3.705 $Y2=2.4
cc_6 VNB N_A_c_82_n 0.016198f $X=-0.19 $Y=-0.245 $X2=3.94 $Y2=1.22
cc_7 VNB N_A_c_83_n 0.0136474f $X=-0.19 $Y=-0.245 $X2=3.645 $Y2=1.095
cc_8 VNB N_A_c_84_n 0.0161986f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.095
cc_9 VNB N_A_c_85_n 0.00205904f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=1.385
cc_10 VNB N_A_c_86_n 0.0447165f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=1.385
cc_11 VNB N_A_c_87_n 0.0863864f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=1.175
cc_12 VNB N_A_353_323#_c_180_n 0.0180618f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_13 VNB N_A_353_323#_c_181_n 0.0197816f $X=-0.19 $Y=-0.245 $X2=3.705 $Y2=1.55
cc_14 VNB N_A_353_323#_c_182_n 0.00529851f $X=-0.19 $Y=-0.245 $X2=1.295
+ $Y2=1.175
cc_15 VNB N_A_353_323#_c_183_n 0.107436f $X=-0.19 $Y=-0.245 $X2=3.705 $Y2=1.385
cc_16 VNB N_A_353_323#_c_184_n 0.0346171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B_N_M1001_g 0.0395613f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_18 VNB B_N 0.0261981f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_19 VNB N_B_N_c_284_n 0.0405493f $X=-0.19 $Y=-0.245 $X2=3.705 $Y2=2.4
cc_20 VNB N_VPWR_c_316_n 0.223389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_438_n 0.0115493f $X=-0.19 $Y=-0.245 $X2=3.51 $Y2=0.74
cc_22 VNB N_Y_c_439_n 0.00816012f $X=-0.19 $Y=-0.245 $X2=3.705 $Y2=2.4
cc_23 VNB N_Y_c_440_n 6.68229e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_441_n 8.97027e-19 $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_25 VNB N_Y_c_442_n 0.00230198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_443_n 0.032652f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.175
cc_27 VNB Y 0.0283086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB Y 0.0173879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_523_n 0.0166025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_524_n 0.00489167f $X=-0.19 $Y=-0.245 $X2=3.705 $Y2=2.4
cc_31 VNB N_VGND_c_525_n 0.0455645f $X=-0.19 $Y=-0.245 $X2=3.94 $Y2=0.74
cc_32 VNB N_VGND_c_526_n 0.0170209f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_33 VNB N_VGND_c_527_n 0.0292937f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=1.175
cc_34 VNB N_VGND_c_528_n 0.303426f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=1.175
cc_35 VNB N_VGND_c_529_n 0.00631651f $X=-0.19 $Y=-0.245 $X2=3.705 $Y2=1.385
cc_36 VNB N_VGND_c_530_n 0.0186046f $X=-0.19 $Y=-0.245 $X2=1.295 $Y2=1.21
cc_37 VNB N_VGND_c_531_n 0.0247843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_532_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_A_M1004_g 0.0279777f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_40 VPB N_A_M1005_g 0.0216908f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_41 VPB N_A_M1007_g 0.0214722f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_42 VPB N_A_M1012_g 0.0237814f $X=-0.19 $Y=1.66 $X2=3.705 $Y2=2.4
cc_43 VPB N_A_353_323#_c_185_n 0.0157733f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_44 VPB N_A_353_323#_c_186_n 0.0159149f $X=-0.19 $Y=1.66 $X2=3.51 $Y2=1.22
cc_45 VPB N_A_353_323#_c_187_n 0.0159175f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A_353_323#_c_188_n 0.0157059f $X=-0.19 $Y=1.66 $X2=3.94 $Y2=0.74
cc_47 VPB N_A_353_323#_c_189_n 7.4105e-19 $X=-0.19 $Y=1.66 $X2=3.81 $Y2=1.18
cc_48 VPB N_A_353_323#_c_190_n 0.017297f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.21
cc_49 VPB N_A_353_323#_c_191_n 0.00612873f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.175
cc_50 VPB N_A_353_323#_c_183_n 0.027815f $X=-0.19 $Y=1.66 $X2=3.705 $Y2=1.385
cc_51 VPB N_B_N_c_285_n 0.0166837f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.34
cc_52 VPB N_B_N_c_286_n 0.0179902f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB B_N 0.00796315f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_54 VPB N_B_N_c_284_n 0.0536259f $X=-0.19 $Y=1.66 $X2=3.705 $Y2=2.4
cc_55 VPB N_VPWR_c_317_n 0.0106521f $X=-0.19 $Y=1.66 $X2=3.51 $Y2=1.22
cc_56 VPB N_VPWR_c_318_n 0.0535771f $X=-0.19 $Y=1.66 $X2=3.51 $Y2=0.74
cc_57 VPB N_VPWR_c_319_n 0.00768031f $X=-0.19 $Y=1.66 $X2=3.94 $Y2=0.74
cc_58 VPB N_VPWR_c_320_n 0.0132011f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=1.18
cc_59 VPB N_VPWR_c_321_n 0.0117686f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_322_n 0.0541822f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.21
cc_61 VPB N_VPWR_c_323_n 0.0597948f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.175
cc_62 VPB N_VPWR_c_324_n 0.00631788f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.175
cc_63 VPB N_VPWR_c_325_n 0.0206041f $X=-0.19 $Y=1.66 $X2=1.295 $Y2=1.175
cc_64 VPB N_VPWR_c_326_n 0.0212408f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.21
cc_65 VPB N_VPWR_c_327_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_316_n 0.0780916f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_A_119_368#_c_381_n 0.00231613f $X=-0.19 $Y=1.66 $X2=3.51 $Y2=0.74
cc_68 VPB N_A_119_368#_c_382_n 0.00227131f $X=-0.19 $Y=1.66 $X2=3.645 $Y2=1.095
cc_69 VPB N_A_119_368#_c_383_n 0.00160153f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.095
cc_70 VPB N_A_119_368#_c_384_n 0.00424161f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_A_119_368#_c_385_n 0.00196526f $X=-0.19 $Y=1.66 $X2=3.705 $Y2=1.385
cc_72 VPB N_Y_c_439_n 0.00767295f $X=-0.19 $Y=1.66 $X2=3.705 $Y2=2.4
cc_73 VPB N_Y_c_440_n 7.1566e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_Y_c_441_n 0.00182538f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.21
cc_75 VPB N_Y_c_442_n 0.00101457f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB Y 0.00244476f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 N_A_c_83_n N_A_353_323#_c_180_n 0.0125877f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_78 N_A_c_84_n N_A_353_323#_c_180_n 0.00632392f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_79 N_A_c_87_n N_A_353_323#_c_180_n 0.00840639f $X=1.295 $Y=1.175 $X2=0 $Y2=0
cc_80 N_A_c_83_n N_A_353_323#_c_181_n 0.0125331f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_81 N_A_c_83_n N_A_353_323#_c_189_n 0.0749937f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_82 N_A_c_84_n N_A_353_323#_c_189_n 0.00262271f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_83 N_A_c_85_n N_A_353_323#_c_189_n 0.00688023f $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_84 N_A_c_86_n N_A_353_323#_c_189_n 0.00184555f $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_85 N_A_M1012_g N_A_353_323#_c_190_n 0.017669f $X=3.705 $Y=2.4 $X2=0 $Y2=0
cc_86 N_A_c_83_n N_A_353_323#_c_190_n 0.0132262f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_87 N_A_c_85_n N_A_353_323#_c_190_n 0.0251788f $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_88 N_A_c_86_n N_A_353_323#_c_190_n 0.0073225f $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_89 N_A_M1012_g N_A_353_323#_c_191_n 5.22703e-19 $X=3.705 $Y=2.4 $X2=0 $Y2=0
cc_90 N_A_M1012_g N_A_353_323#_c_182_n 7.73468e-19 $X=3.705 $Y=2.4 $X2=0 $Y2=0
cc_91 N_A_c_82_n N_A_353_323#_c_182_n 0.00177623f $X=3.94 $Y=1.22 $X2=0 $Y2=0
cc_92 N_A_c_83_n N_A_353_323#_c_182_n 0.00603876f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_93 N_A_c_85_n N_A_353_323#_c_182_n 0.0123049f $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_94 N_A_M1007_g N_A_353_323#_c_183_n 0.0279017f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_95 N_A_M1012_g N_A_353_323#_c_183_n 0.0190407f $X=3.705 $Y=2.4 $X2=0 $Y2=0
cc_96 N_A_c_83_n N_A_353_323#_c_183_n 0.0276696f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_97 N_A_c_84_n N_A_353_323#_c_183_n 2.03013e-19 $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_98 N_A_c_85_n N_A_353_323#_c_183_n 0.00151745f $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_99 N_A_c_86_n N_A_353_323#_c_183_n 0.019063f $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_100 N_A_c_82_n N_A_353_323#_c_184_n 9.69162e-19 $X=3.94 $Y=1.22 $X2=0 $Y2=0
cc_101 N_A_c_82_n N_B_N_M1001_g 0.0194276f $X=3.94 $Y=1.22 $X2=0 $Y2=0
cc_102 N_A_c_83_n N_B_N_M1001_g 5.68631e-19 $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_103 N_A_c_85_n N_B_N_M1001_g 0.001297f $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_104 N_A_M1012_g N_B_N_c_284_n 0.0231272f $X=3.705 $Y=2.4 $X2=0 $Y2=0
cc_105 N_A_c_86_n N_B_N_c_284_n 0.0194276f $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_106 N_A_M1004_g N_VPWR_c_318_n 0.00542061f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_107 N_A_M1005_g N_VPWR_c_319_n 0.0027763f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_108 N_A_M1007_g N_VPWR_c_319_n 0.00120619f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_109 N_A_M1012_g N_VPWR_c_320_n 0.00305677f $X=3.705 $Y=2.4 $X2=0 $Y2=0
cc_110 N_A_M1007_g N_VPWR_c_323_n 0.00517089f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_111 N_A_M1012_g N_VPWR_c_323_n 0.00517089f $X=3.705 $Y=2.4 $X2=0 $Y2=0
cc_112 N_A_M1004_g N_VPWR_c_325_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_113 N_A_M1005_g N_VPWR_c_325_n 0.005209f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_114 N_A_M1004_g N_VPWR_c_316_n 0.00986008f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_115 N_A_M1005_g N_VPWR_c_316_n 0.00982266f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_116 N_A_M1007_g N_VPWR_c_316_n 0.00977588f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_117 N_A_M1012_g N_VPWR_c_316_n 0.00982505f $X=3.705 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A_M1004_g N_A_119_368#_c_386_n 0.0025567f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A_M1005_g N_A_119_368#_c_386_n 8.84614e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A_M1004_g N_A_119_368#_c_381_n 0.0116401f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_121 N_A_M1005_g N_A_119_368#_c_381_n 0.0122944f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_122 N_A_M1007_g N_A_119_368#_c_381_n 6.60002e-19 $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_123 N_A_M1005_g N_A_119_368#_c_391_n 0.0128923f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_124 N_A_M1007_g N_A_119_368#_c_391_n 0.012931f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_125 N_A_M1007_g N_A_119_368#_c_393_n 8.84614e-19 $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_126 N_A_M1005_g N_A_119_368#_c_394_n 6.38352e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_127 N_A_M1007_g N_A_119_368#_c_394_n 0.0108845f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_128 N_A_M1007_g N_A_119_368#_c_383_n 0.00347836f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_129 N_A_M1012_g N_A_119_368#_c_384_n 0.00362176f $X=3.705 $Y=2.4 $X2=0 $Y2=0
cc_130 N_A_M1012_g N_A_119_368#_c_398_n 0.0100211f $X=3.705 $Y=2.4 $X2=0 $Y2=0
cc_131 N_A_c_83_n N_Y_M1006_d 0.00176891f $X=3.645 $Y=1.095 $X2=-0.19 $Y2=-0.245
cc_132 N_A_c_83_n N_Y_M1003_d 0.00178017f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_133 N_A_M1005_g N_Y_c_439_n 0.0121287f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_134 N_A_M1007_g N_Y_c_439_n 0.0117857f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_135 N_A_c_83_n N_Y_c_439_n 0.0037097f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_136 N_A_c_84_n N_Y_c_439_n 0.0724897f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_137 N_A_c_87_n N_Y_c_439_n 0.00294898f $X=1.295 $Y=1.175 $X2=0 $Y2=0
cc_138 N_A_M1007_g N_Y_c_440_n 7.92833e-19 $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A_c_83_n N_Y_c_440_n 0.0100147f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_140 N_A_c_80_n N_Y_c_460_n 0.0110659f $X=3.51 $Y=1.22 $X2=0 $Y2=0
cc_141 N_A_M1004_g N_Y_c_441_n 0.0133495f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_142 N_A_M1004_g N_Y_c_442_n 0.0101629f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_143 N_A_M1005_g N_Y_c_442_n 0.00180432f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A_c_87_n N_Y_c_442_n 5.58672e-19 $X=1.295 $Y=1.175 $X2=0 $Y2=0
cc_145 N_A_c_83_n N_Y_c_443_n 0.105987f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_146 N_A_c_84_n N_Y_c_443_n 0.0773139f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_147 N_A_c_87_n N_Y_c_443_n 0.0169737f $X=1.295 $Y=1.175 $X2=0 $Y2=0
cc_148 N_A_c_80_n N_Y_c_468_n 0.00837425f $X=3.51 $Y=1.22 $X2=0 $Y2=0
cc_149 N_A_c_83_n N_Y_c_468_n 0.0155098f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_150 N_A_c_86_n N_Y_c_468_n 4.50695e-19 $X=3.81 $Y=1.385 $X2=0 $Y2=0
cc_151 N_A_c_84_n Y 0.0114186f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_152 N_A_c_87_n Y 0.00943558f $X=1.295 $Y=1.175 $X2=0 $Y2=0
cc_153 N_A_c_84_n Y 0.00181037f $X=1.795 $Y=1.095 $X2=0 $Y2=0
cc_154 N_A_c_87_n Y 0.0083228f $X=1.295 $Y=1.175 $X2=0 $Y2=0
cc_155 N_A_c_83_n N_VGND_M1006_s 8.73801e-19 $X=3.645 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_156 N_A_c_84_n N_VGND_M1006_s 0.00289875f $X=1.795 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_157 N_A_c_83_n N_VGND_M1014_s 0.0116574f $X=3.645 $Y=1.095 $X2=0 $Y2=0
cc_158 N_A_c_80_n N_VGND_c_524_n 7.7967e-19 $X=3.51 $Y=1.22 $X2=0 $Y2=0
cc_159 N_A_c_82_n N_VGND_c_524_n 0.0122954f $X=3.94 $Y=1.22 $X2=0 $Y2=0
cc_160 N_A_c_80_n N_VGND_c_526_n 0.00327917f $X=3.51 $Y=1.22 $X2=0 $Y2=0
cc_161 N_A_c_82_n N_VGND_c_526_n 0.00383152f $X=3.94 $Y=1.22 $X2=0 $Y2=0
cc_162 N_A_c_80_n N_VGND_c_528_n 0.00418901f $X=3.51 $Y=1.22 $X2=0 $Y2=0
cc_163 N_A_c_82_n N_VGND_c_528_n 0.0075754f $X=3.94 $Y=1.22 $X2=0 $Y2=0
cc_164 N_A_c_80_n N_VGND_c_531_n 0.00641807f $X=3.51 $Y=1.22 $X2=0 $Y2=0
cc_165 N_A_353_323#_c_191_n N_B_N_c_285_n 0.0155689f $X=4.515 $Y=2.16 $X2=-0.19
+ $Y2=-0.245
cc_166 N_A_353_323#_c_182_n N_B_N_M1001_g 0.0158316f $X=4.495 $Y=1.72 $X2=0
+ $Y2=0
cc_167 N_A_353_323#_c_184_n N_B_N_M1001_g 0.00981473f $X=5 $Y=0.505 $X2=0 $Y2=0
cc_168 N_A_353_323#_c_191_n N_B_N_c_286_n 0.0165147f $X=4.515 $Y=2.16 $X2=0
+ $Y2=0
cc_169 N_A_353_323#_c_191_n B_N 0.0085076f $X=4.515 $Y=2.16 $X2=0 $Y2=0
cc_170 N_A_353_323#_c_182_n B_N 0.0416881f $X=4.495 $Y=1.72 $X2=0 $Y2=0
cc_171 N_A_353_323#_c_184_n B_N 0.0366877f $X=5 $Y=0.505 $X2=0 $Y2=0
cc_172 N_A_353_323#_c_190_n N_B_N_c_284_n 0.0150009f $X=4.35 $Y=1.805 $X2=0
+ $Y2=0
cc_173 N_A_353_323#_c_191_n N_B_N_c_284_n 0.0178372f $X=4.515 $Y=2.16 $X2=0
+ $Y2=0
cc_174 N_A_353_323#_c_182_n N_B_N_c_284_n 0.0133442f $X=4.495 $Y=1.72 $X2=0
+ $Y2=0
cc_175 N_A_353_323#_c_184_n N_B_N_c_284_n 0.00745702f $X=5 $Y=0.505 $X2=0 $Y2=0
cc_176 N_A_353_323#_c_190_n N_VPWR_M1012_s 0.00302409f $X=4.35 $Y=1.805 $X2=0
+ $Y2=0
cc_177 N_A_353_323#_c_190_n N_VPWR_c_320_n 0.0237371f $X=4.35 $Y=1.805 $X2=0
+ $Y2=0
cc_178 N_A_353_323#_c_191_n N_VPWR_c_320_n 0.0237568f $X=4.515 $Y=2.16 $X2=0
+ $Y2=0
cc_179 N_A_353_323#_c_191_n N_VPWR_c_322_n 0.0303402f $X=4.515 $Y=2.16 $X2=0
+ $Y2=0
cc_180 N_A_353_323#_c_185_n N_VPWR_c_323_n 0.00333926f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_181 N_A_353_323#_c_186_n N_VPWR_c_323_n 0.00333896f $X=2.305 $Y=1.765 $X2=0
+ $Y2=0
cc_182 N_A_353_323#_c_187_n N_VPWR_c_323_n 0.00333896f $X=2.755 $Y=1.765 $X2=0
+ $Y2=0
cc_183 N_A_353_323#_c_188_n N_VPWR_c_323_n 0.00333926f $X=3.205 $Y=1.765 $X2=0
+ $Y2=0
cc_184 N_A_353_323#_c_191_n N_VPWR_c_326_n 0.0101104f $X=4.515 $Y=2.16 $X2=0
+ $Y2=0
cc_185 N_A_353_323#_c_185_n N_VPWR_c_316_n 0.00422798f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_186 N_A_353_323#_c_186_n N_VPWR_c_316_n 0.00422685f $X=2.305 $Y=1.765 $X2=0
+ $Y2=0
cc_187 N_A_353_323#_c_187_n N_VPWR_c_316_n 0.00422685f $X=2.755 $Y=1.765 $X2=0
+ $Y2=0
cc_188 N_A_353_323#_c_188_n N_VPWR_c_316_n 0.00423254f $X=3.205 $Y=1.765 $X2=0
+ $Y2=0
cc_189 N_A_353_323#_c_191_n N_VPWR_c_316_n 0.0112627f $X=4.515 $Y=2.16 $X2=0
+ $Y2=0
cc_190 N_A_353_323#_c_190_n N_A_119_368#_M1013_s 0.00218982f $X=4.35 $Y=1.805
+ $X2=0 $Y2=0
cc_191 N_A_353_323#_c_185_n N_A_119_368#_c_382_n 0.0130344f $X=1.855 $Y=1.765
+ $X2=0 $Y2=0
cc_192 N_A_353_323#_c_186_n N_A_119_368#_c_382_n 0.00936332f $X=2.305 $Y=1.765
+ $X2=0 $Y2=0
cc_193 N_A_353_323#_c_185_n N_A_119_368#_c_402_n 4.47651e-19 $X=1.855 $Y=1.765
+ $X2=0 $Y2=0
cc_194 N_A_353_323#_c_186_n N_A_119_368#_c_402_n 0.00781935f $X=2.305 $Y=1.765
+ $X2=0 $Y2=0
cc_195 N_A_353_323#_c_187_n N_A_119_368#_c_402_n 0.00774767f $X=2.755 $Y=1.765
+ $X2=0 $Y2=0
cc_196 N_A_353_323#_c_188_n N_A_119_368#_c_402_n 4.41999e-19 $X=3.205 $Y=1.765
+ $X2=0 $Y2=0
cc_197 N_A_353_323#_c_187_n N_A_119_368#_c_384_n 0.00936332f $X=2.755 $Y=1.765
+ $X2=0 $Y2=0
cc_198 N_A_353_323#_c_188_n N_A_119_368#_c_384_n 0.0141392f $X=3.205 $Y=1.765
+ $X2=0 $Y2=0
cc_199 N_A_353_323#_c_190_n N_A_119_368#_c_398_n 0.0189268f $X=4.35 $Y=1.805
+ $X2=0 $Y2=0
cc_200 N_A_353_323#_c_186_n N_A_119_368#_c_385_n 0.00193733f $X=2.305 $Y=1.765
+ $X2=0 $Y2=0
cc_201 N_A_353_323#_c_187_n N_A_119_368#_c_385_n 0.00193733f $X=2.755 $Y=1.765
+ $X2=0 $Y2=0
cc_202 N_A_353_323#_c_189_n N_Y_M1011_d 5.96688e-19 $X=3.055 $Y=1.515 $X2=0
+ $Y2=0
cc_203 N_A_353_323#_c_183_n N_Y_c_439_n 0.0100577f $X=3.06 $Y=1.515 $X2=0 $Y2=0
cc_204 N_A_353_323#_c_185_n N_Y_c_440_n 0.00798552f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_205 N_A_353_323#_c_186_n N_Y_c_440_n 0.00175036f $X=2.305 $Y=1.765 $X2=0
+ $Y2=0
cc_206 N_A_353_323#_c_189_n N_Y_c_440_n 0.00838044f $X=3.055 $Y=1.515 $X2=0
+ $Y2=0
cc_207 N_A_353_323#_c_183_n N_Y_c_440_n 0.0160804f $X=3.06 $Y=1.515 $X2=0 $Y2=0
cc_208 N_A_353_323#_c_185_n N_Y_c_481_n 0.00877682f $X=1.855 $Y=1.765 $X2=0
+ $Y2=0
cc_209 N_A_353_323#_c_186_n N_Y_c_482_n 0.0137546f $X=2.305 $Y=1.765 $X2=0 $Y2=0
cc_210 N_A_353_323#_c_187_n N_Y_c_482_n 0.0132973f $X=2.755 $Y=1.765 $X2=0 $Y2=0
cc_211 N_A_353_323#_c_189_n N_Y_c_482_n 0.0224947f $X=3.055 $Y=1.515 $X2=0 $Y2=0
cc_212 N_A_353_323#_c_183_n N_Y_c_482_n 0.00214309f $X=3.06 $Y=1.515 $X2=0 $Y2=0
cc_213 N_A_353_323#_c_181_n N_Y_c_460_n 0.0105158f $X=2.44 $Y=1.225 $X2=0 $Y2=0
cc_214 N_A_353_323#_c_188_n N_Y_c_487_n 0.00232812f $X=3.205 $Y=1.765 $X2=0
+ $Y2=0
cc_215 N_A_353_323#_c_189_n N_Y_c_487_n 0.00938901f $X=3.055 $Y=1.515 $X2=0
+ $Y2=0
cc_216 N_A_353_323#_c_183_n N_Y_c_487_n 0.00222422f $X=3.06 $Y=1.515 $X2=0 $Y2=0
cc_217 N_A_353_323#_c_188_n N_Y_c_490_n 0.00638746f $X=3.205 $Y=1.765 $X2=0
+ $Y2=0
cc_218 N_A_353_323#_c_180_n N_Y_c_443_n 0.0105158f $X=2.01 $Y=1.225 $X2=0 $Y2=0
cc_219 N_A_353_323#_c_180_n N_Y_c_492_n 0.00718488f $X=2.01 $Y=1.225 $X2=0 $Y2=0
cc_220 N_A_353_323#_c_181_n N_Y_c_492_n 0.00718488f $X=2.44 $Y=1.225 $X2=0 $Y2=0
cc_221 N_A_353_323#_c_180_n N_VGND_c_523_n 0.00789696f $X=2.01 $Y=1.225 $X2=0
+ $Y2=0
cc_222 N_A_353_323#_c_184_n N_VGND_c_524_n 0.0217307f $X=5 $Y=0.505 $X2=0 $Y2=0
cc_223 N_A_353_323#_c_184_n N_VGND_c_527_n 0.0340697f $X=5 $Y=0.505 $X2=0 $Y2=0
cc_224 N_A_353_323#_c_180_n N_VGND_c_528_n 0.00420785f $X=2.01 $Y=1.225 $X2=0
+ $Y2=0
cc_225 N_A_353_323#_c_181_n N_VGND_c_528_n 0.00420763f $X=2.44 $Y=1.225 $X2=0
+ $Y2=0
cc_226 N_A_353_323#_c_184_n N_VGND_c_528_n 0.027759f $X=5 $Y=0.505 $X2=0 $Y2=0
cc_227 N_A_353_323#_c_180_n N_VGND_c_530_n 0.00327334f $X=2.01 $Y=1.225 $X2=0
+ $Y2=0
cc_228 N_A_353_323#_c_181_n N_VGND_c_530_n 0.00327334f $X=2.44 $Y=1.225 $X2=0
+ $Y2=0
cc_229 N_A_353_323#_c_181_n N_VGND_c_531_n 0.00845421f $X=2.44 $Y=1.225 $X2=0
+ $Y2=0
cc_230 N_B_N_c_285_n N_VPWR_c_320_n 0.00816104f $X=4.29 $Y=1.94 $X2=0 $Y2=0
cc_231 N_B_N_c_286_n N_VPWR_c_322_n 0.00873548f $X=4.74 $Y=1.94 $X2=0 $Y2=0
cc_232 B_N N_VPWR_c_322_n 0.0223353f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_233 N_B_N_c_284_n N_VPWR_c_322_n 0.00508612f $X=4.74 $Y=1.717 $X2=0 $Y2=0
cc_234 N_B_N_c_285_n N_VPWR_c_326_n 0.00578748f $X=4.29 $Y=1.94 $X2=0 $Y2=0
cc_235 N_B_N_c_286_n N_VPWR_c_326_n 0.00578748f $X=4.74 $Y=1.94 $X2=0 $Y2=0
cc_236 N_B_N_c_285_n N_VPWR_c_316_n 0.00615499f $X=4.29 $Y=1.94 $X2=0 $Y2=0
cc_237 N_B_N_c_286_n N_VPWR_c_316_n 0.00615499f $X=4.74 $Y=1.94 $X2=0 $Y2=0
cc_238 N_B_N_M1001_g N_VGND_c_524_n 0.00333403f $X=4.37 $Y=0.74 $X2=0 $Y2=0
cc_239 N_B_N_M1001_g N_VGND_c_527_n 0.00421682f $X=4.37 $Y=0.74 $X2=0 $Y2=0
cc_240 N_B_N_M1001_g N_VGND_c_528_n 0.00784929f $X=4.37 $Y=0.74 $X2=0 $Y2=0
cc_241 N_VPWR_c_318_n N_A_119_368#_c_381_n 0.0299644f $X=0.28 $Y=2.015 $X2=0
+ $Y2=0
cc_242 N_VPWR_c_319_n N_A_119_368#_c_381_n 0.0243582f $X=1.18 $Y=2.425 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_325_n N_A_119_368#_c_381_n 0.0144623f $X=1.095 $Y=3.33 $X2=0
+ $Y2=0
cc_244 N_VPWR_c_316_n N_A_119_368#_c_381_n 0.0118344f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_245 N_VPWR_M1005_s N_A_119_368#_c_391_n 0.00323401f $X=1.045 $Y=1.84 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_319_n N_A_119_368#_c_391_n 0.0126919f $X=1.18 $Y=2.425 $X2=0
+ $Y2=0
cc_247 N_VPWR_c_323_n N_A_119_368#_c_382_n 0.0408559f $X=3.815 $Y=3.33 $X2=0
+ $Y2=0
cc_248 N_VPWR_c_316_n N_A_119_368#_c_382_n 0.0229294f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_249 N_VPWR_c_319_n N_A_119_368#_c_383_n 0.0101219f $X=1.18 $Y=2.425 $X2=0
+ $Y2=0
cc_250 N_VPWR_c_323_n N_A_119_368#_c_383_n 0.0178163f $X=3.815 $Y=3.33 $X2=0
+ $Y2=0
cc_251 N_VPWR_c_316_n N_A_119_368#_c_383_n 0.00958215f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_252 N_VPWR_c_320_n N_A_119_368#_c_384_n 0.0119238f $X=3.98 $Y=2.145 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_323_n N_A_119_368#_c_384_n 0.0624483f $X=3.815 $Y=3.33 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_316_n N_A_119_368#_c_384_n 0.0344904f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_323_n N_A_119_368#_c_385_n 0.0234328f $X=3.815 $Y=3.33 $X2=0
+ $Y2=0
cc_256 N_VPWR_c_316_n N_A_119_368#_c_385_n 0.0125526f $X=5.04 $Y=3.33 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_318_n N_Y_c_441_n 4.37108e-19 $X=0.28 $Y=2.015 $X2=0 $Y2=0
cc_258 N_VPWR_c_318_n Y 0.0184311f $X=0.28 $Y=2.015 $X2=0 $Y2=0
cc_259 N_A_119_368#_c_382_n N_Y_M1009_d 0.00165831f $X=2.365 $Y=2.99 $X2=0 $Y2=0
cc_260 N_A_119_368#_c_384_n N_Y_M1011_d 0.00163705f $X=3.315 $Y=2.99 $X2=0 $Y2=0
cc_261 N_A_119_368#_c_391_n N_Y_c_439_n 0.0360974f $X=1.465 $Y=2.005 $X2=0 $Y2=0
cc_262 N_A_119_368#_c_393_n N_Y_c_439_n 0.0175624f $X=1.59 $Y=2.09 $X2=0 $Y2=0
cc_263 N_A_119_368#_c_382_n N_Y_c_481_n 0.0160403f $X=2.365 $Y=2.99 $X2=0 $Y2=0
cc_264 N_A_119_368#_M1010_s N_Y_c_482_n 0.00379761f $X=2.395 $Y=1.84 $X2=0 $Y2=0
cc_265 N_A_119_368#_c_382_n N_Y_c_482_n 0.00319714f $X=2.365 $Y=2.99 $X2=0 $Y2=0
cc_266 N_A_119_368#_c_402_n N_Y_c_482_n 0.0170155f $X=2.53 $Y=2.485 $X2=0 $Y2=0
cc_267 N_A_119_368#_c_384_n N_Y_c_482_n 0.00318644f $X=3.315 $Y=2.99 $X2=0 $Y2=0
cc_268 N_A_119_368#_c_384_n N_Y_c_490_n 0.0137427f $X=3.315 $Y=2.99 $X2=0 $Y2=0
cc_269 N_A_119_368#_c_386_n N_Y_c_442_n 0.0219373f $X=0.73 $Y=2.09 $X2=0 $Y2=0
cc_270 N_Y_c_443_n N_VGND_M1006_s 0.00811085f $X=2.06 $Y=0.685 $X2=-0.19
+ $Y2=-0.245
cc_271 N_Y_c_460_n N_VGND_M1014_s 0.0210657f $X=3.56 $Y=0.755 $X2=0 $Y2=0
cc_272 N_Y_c_443_n N_VGND_c_523_n 0.0252515f $X=2.06 $Y=0.685 $X2=0 $Y2=0
cc_273 N_Y_c_438_n N_VGND_c_525_n 0.00433932f $X=0.355 $Y=0.755 $X2=0 $Y2=0
cc_274 N_Y_c_443_n N_VGND_c_525_n 0.0202416f $X=2.06 $Y=0.685 $X2=0 $Y2=0
cc_275 N_Y_c_460_n N_VGND_c_526_n 0.0023667f $X=3.56 $Y=0.755 $X2=0 $Y2=0
cc_276 N_Y_c_468_n N_VGND_c_526_n 0.00544924f $X=3.725 $Y=0.675 $X2=0 $Y2=0
cc_277 N_Y_c_438_n N_VGND_c_528_n 0.00680159f $X=0.355 $Y=0.755 $X2=0 $Y2=0
cc_278 N_Y_c_460_n N_VGND_c_528_n 0.0121701f $X=3.56 $Y=0.755 $X2=0 $Y2=0
cc_279 N_Y_c_443_n N_VGND_c_528_n 0.0390596f $X=2.06 $Y=0.685 $X2=0 $Y2=0
cc_280 N_Y_c_492_n N_VGND_c_528_n 0.0101808f $X=2.39 $Y=0.685 $X2=0 $Y2=0
cc_281 N_Y_c_468_n N_VGND_c_528_n 0.00786294f $X=3.725 $Y=0.675 $X2=0 $Y2=0
cc_282 N_Y_c_460_n N_VGND_c_530_n 0.00236055f $X=3.56 $Y=0.755 $X2=0 $Y2=0
cc_283 N_Y_c_443_n N_VGND_c_530_n 0.00236055f $X=2.06 $Y=0.685 $X2=0 $Y2=0
cc_284 N_Y_c_492_n N_VGND_c_530_n 0.00642607f $X=2.39 $Y=0.685 $X2=0 $Y2=0
cc_285 N_Y_c_460_n N_VGND_c_531_n 0.061776f $X=3.56 $Y=0.755 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__ha_1.spice
* Created: Fri Aug 28 17:37:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__ha_1.pex.spice"
.subckt sky130_fd_sc_ms__ha_1  VNB VPB B A SUM VPWR COUT VGND
* 
* VGND	VGND
* COUT	COUT
* VPWR	VPWR
* SUM	SUM
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A_83_260#_M1011_g N_SUM_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.19515 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_A_305_130#_M1007_d N_A_239_294#_M1007_g N_A_83_260#_M1007_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.1726 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1009 N_VGND_M1009_d N_B_M1009_g N_A_305_130#_M1007_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.125537 AS=0.0896 PD=1.065 PS=0.92 NRD=1.872 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1013 N_A_305_130#_M1013_d N_A_M1013_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.125537 PD=1.85 PS=1.065 NRD=0 NRS=16.872 M=1 R=4.26667
+ SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 A_695_119# N_B_M1001_g N_A_239_294#_M1001_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1824 PD=0.85 PS=1.85 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1010 N_VGND_M1010_d N_A_M1010_g A_695_119# VNB NLOWVT L=0.15 W=0.64
+ AD=0.115478 AS=0.0672 PD=1.01101 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667
+ SA=75000.6 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1004 N_COUT_M1004_d N_A_239_294#_M1004_g N_VGND_M1010_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.133522 PD=2.05 PS=1.16899 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_A_83_260#_M1005_g N_SUM_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.390286 AS=0.3136 PD=2.04 PS=2.8 NRD=32.5247 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90002.8 A=0.2016 P=2.6 MULT=1
MM1006 N_A_83_260#_M1006_d N_A_239_294#_M1006_g N_VPWR_M1005_d VPB PSHORT L=0.18
+ W=0.84 AD=0.142891 AS=0.292714 PD=1.20978 PS=1.53 NRD=0 NRS=48.068 M=1
+ R=4.66667 SA=90001 SB=90002.7 A=0.1512 P=2.04 MULT=1
MM1003 A_389_392# N_B_M1003_g N_A_83_260#_M1006_d VPB PSHORT L=0.18 W=1 AD=0.195
+ AS=0.170109 PD=1.39 PS=1.44022 NRD=27.5603 NRS=9.8303 M=1 R=5.55556 SA=90001.3
+ SB=90002.3 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g A_389_392# VPB PSHORT L=0.18 W=1 AD=0.316196
+ AS=0.195 PD=1.78804 PS=1.39 NRD=0 NRS=27.5603 M=1 R=5.55556 SA=90001.9
+ SB=90001.7 A=0.18 P=2.36 MULT=1
MM1012 N_A_239_294#_M1012_d N_B_M1012_g N_VPWR_M1002_d VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.265604 PD=1.11 PS=1.50196 NRD=0 NRS=0 M=1 R=4.66667 SA=90002.7
+ SB=90001.2 A=0.1512 P=2.04 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_239_294#_M1012_d VPB PSHORT L=0.18 W=0.84
+ AD=0.1632 AS=0.1134 PD=1.27714 PS=1.11 NRD=10.5395 NRS=0 M=1 R=4.66667
+ SA=90003.1 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1008 N_COUT_M1008_d N_A_239_294#_M1008_g N_VPWR_M1000_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.2176 PD=2.8 PS=1.70286 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90002.8 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.471 P=14.32
c_88 VPB 0 2.55746e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__ha_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__nand3b_2.spice
* Created: Fri Aug 28 17:44:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nand3b_2.pex.spice"
.subckt sky130_fd_sc_ms__nand3b_2  VNB VPB A_N C B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* C	C
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_N_M1002_g N_A_27_94#_M1002_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.108058 AS=0.1728 PD=0.987826 PS=1.82 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1001 N_A_206_74#_M1001_d N_C_M1001_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.124942 PD=1.02 PS=1.14217 NRD=0 NRS=7.296 M=1 R=4.93333
+ SA=75000.6 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1008 N_A_206_74#_M1001_d N_C_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.19445 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_Y_M1006_d N_A_27_94#_M1006_g N_A_403_54#_M1006_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.24845 PD=1.02 PS=2.6 NRD=0 NRS=45.516 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1007 N_Y_M1006_d N_A_27_94#_M1007_g N_A_403_54#_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1816 PD=1.02 PS=1.38 NRD=0 NRS=30.876 M=1 R=4.93333
+ SA=75000.6 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1010 N_A_206_74#_M1010_d N_B_M1010_g N_A_403_54#_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1816 PD=1.02 PS=1.38 NRD=0 NRS=30.876 M=1 R=4.93333
+ SA=75001.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1011 N_A_206_74#_M1010_d N_B_M1011_g N_A_403_54#_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1998 PD=1.02 PS=2.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_A_N_M1000_g N_A_27_94#_M1000_s VPB PSHORT L=0.18 W=1
+ AD=0.167453 AS=0.28 PD=1.36321 PS=2.56 NRD=4.9053 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90003.3 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1000_d N_C_M1003_g N_Y_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.187547 AS=0.1764 PD=1.52679 PS=1.435 NRD=3.5066 NRS=2.6201 M=1 R=6.22222
+ SA=90000.6 SB=90002.8 A=0.2016 P=2.6 MULT=1
MM1013 N_VPWR_M1013_d N_C_M1013_g N_Y_M1003_s VPB PSHORT L=0.18 W=1.12 AD=0.1792
+ AS=0.1764 PD=1.44 PS=1.435 NRD=7.8997 NRS=3.5066 M=1 R=6.22222 SA=90001.1
+ SB=90002.3 A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1004_d N_A_27_94#_M1004_g N_VPWR_M1013_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.6
+ SB=90001.8 A=0.2016 P=2.6 MULT=1
MM1005 N_Y_M1004_d N_A_27_94#_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2688 PD=1.39 PS=1.6 NRD=0 NRS=14.0658 M=1 R=6.22222 SA=90002.1
+ SB=90001.4 A=0.2016 P=2.6 MULT=1
MM1009 N_Y_M1009_d N_B_M1009_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12 AD=0.1848
+ AS=0.2688 PD=1.45 PS=1.6 NRD=0 NRS=21.0987 M=1 R=6.22222 SA=90002.7 SB=90000.7
+ A=0.2016 P=2.6 MULT=1
MM1012 N_Y_M1009_d N_B_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12 AD=0.1848
+ AS=0.3136 PD=1.45 PS=2.8 NRD=9.6727 NRS=0 M=1 R=6.22222 SA=90003.3 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__nand3b_2.pxi.spice"
*
.ends
*
*

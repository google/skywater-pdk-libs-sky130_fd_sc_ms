* File: sky130_fd_sc_ms__a2bb2oi_2.pex.spice
* Created: Fri Aug 28 17:04:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A2BB2OI_2%A1_N 1 3 5 10 12 14 18
r27 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=0.45 $X2=0.27 $Y2=0.45
r28 14 17 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.27 $Y=0.36 $X2=0.27
+ $Y2=0.45
r29 12 18 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=0.27 $Y=0.555
+ $X2=0.27 $Y2=0.45
r30 10 11 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.985 $Y=0.83
+ $X2=0.985 $Y2=1.225
r31 7 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.985 $Y=0.435
+ $X2=0.985 $Y2=0.83
r32 3 11 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.97 $Y=1.315 $X2=0.97
+ $Y2=1.225
r33 3 5 445.073 $w=1.8e-07 $l=1.145e-06 $layer=POLY_cond $X=0.97 $Y=1.315
+ $X2=0.97 $Y2=2.46
r34 2 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.435 $Y=0.36
+ $X2=0.27 $Y2=0.36
r35 1 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.91 $Y=0.36
+ $X2=0.985 $Y2=0.435
r36 1 2 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=0.91 $Y=0.36
+ $X2=0.435 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_2%A2_N 3 7 9 12 13
c35 13 0 1.88217e-19 $X=1.435 $Y=1.615
c36 7 0 1.77687e-19 $X=1.46 $Y=0.83
r37 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.435 $Y=1.615
+ $X2=1.435 $Y2=1.78
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.435 $Y=1.615
+ $X2=1.435 $Y2=1.45
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.435
+ $Y=1.615 $X2=1.435 $Y2=1.615
r40 9 13 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=1.435 $Y2=1.615
r41 7 14 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=1.46 $Y=0.83 $X2=1.46
+ $Y2=1.45
r42 3 15 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=1.36 $Y=2.46 $X2=1.36
+ $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_2%A_212_102# 1 2 9 13 17 19 20 23 27 29 30
+ 33 35 38 39
c91 39 0 1.56524e-19 $X=1.665 $Y=1.95
c92 27 0 1.77687e-19 $X=1.22 $Y=0.655
c93 20 0 1.88217e-19 $X=2.56 $Y=1.575
c94 17 0 1.0233e-19 $X=2.47 $Y=2.4
r95 43 46 54.2649 $w=3.02e-07 $l=3.4e-07 $layer=POLY_cond $X=2.04 $Y=1.485
+ $X2=2.38 $Y2=1.485
r96 43 44 14.3642 $w=3.02e-07 $l=9e-08 $layer=POLY_cond $X=2.04 $Y=1.485
+ $X2=1.95 $Y2=1.485
r97 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.04
+ $Y=1.485 $X2=2.04 $Y2=1.485
r98 38 39 9.45624 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.665 $Y=2.115
+ $X2=1.665 $Y2=1.95
r99 35 42 8.98608 $w=3.5e-07 $l=2.26892e-07 $layer=LI1_cond $X=1.825 $Y=1.65
+ $X2=1.972 $Y2=1.485
r100 35 39 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.825 $Y=1.65
+ $X2=1.825 $Y2=1.95
r101 31 38 1.95278 $w=4.88e-07 $l=8e-08 $layer=LI1_cond $X=1.665 $Y=2.195
+ $X2=1.665 $Y2=2.115
r102 31 33 15.1341 $w=4.88e-07 $l=6.2e-07 $layer=LI1_cond $X=1.665 $Y=2.195
+ $X2=1.665 $Y2=2.815
r103 29 42 10.1086 $w=3.5e-07 $l=3.89076e-07 $layer=LI1_cond $X=1.74 $Y=1.195
+ $X2=1.972 $Y2=1.485
r104 29 30 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.74 $Y=1.195
+ $X2=1.33 $Y2=1.195
r105 25 30 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=1.182 $Y=1.11
+ $X2=1.33 $Y2=1.195
r106 25 27 17.775 $w=2.93e-07 $l=4.55e-07 $layer=LI1_cond $X=1.182 $Y=1.11
+ $X2=1.182 $Y2=0.655
r107 21 23 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=2.92 $Y=1.65
+ $X2=2.92 $Y2=2.4
r108 19 21 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.83 $Y=1.575
+ $X2=2.92 $Y2=1.65
r109 19 20 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.83 $Y=1.575
+ $X2=2.56 $Y2=1.575
r110 15 20 26.5744 $w=3.02e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.47 $Y=1.65
+ $X2=2.56 $Y2=1.575
r111 15 46 14.3642 $w=3.02e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.47 $Y=1.65
+ $X2=2.38 $Y2=1.485
r112 15 17 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=2.47 $Y=1.65
+ $X2=2.47 $Y2=2.4
r113 11 46 19.1248 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.38 $Y=1.32
+ $X2=2.38 $Y2=1.485
r114 11 13 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.38 $Y=1.32
+ $X2=2.38 $Y2=0.78
r115 7 44 19.1248 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.95 $Y=1.32
+ $X2=1.95 $Y2=1.485
r116 7 9 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.95 $Y=1.32 $X2=1.95
+ $Y2=0.78
r117 2 38 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=1.45
+ $Y=1.96 $X2=1.585 $Y2=2.115
r118 2 33 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.45
+ $Y=1.96 $X2=1.585 $Y2=2.815
r119 1 27 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=1.06
+ $Y=0.51 $X2=1.22 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_2%B2 3 7 11 15 17 23 24
c52 23 0 1.29225e-19 $X=3.57 $Y=1.485
c53 15 0 2.40437e-20 $X=3.845 $Y=0.74
c54 11 0 1.47716e-19 $X=3.82 $Y=2.4
r55 24 25 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=3.82 $Y=1.485
+ $X2=3.845 $Y2=1.485
r56 22 24 36.8502 $w=3.27e-07 $l=2.5e-07 $layer=POLY_cond $X=3.57 $Y=1.485
+ $X2=3.82 $Y2=1.485
r57 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.57
+ $Y=1.485 $X2=3.57 $Y2=1.485
r58 20 22 22.8471 $w=3.27e-07 $l=1.55e-07 $layer=POLY_cond $X=3.415 $Y=1.485
+ $X2=3.57 $Y2=1.485
r59 19 20 6.63303 $w=3.27e-07 $l=4.5e-08 $layer=POLY_cond $X=3.37 $Y=1.485
+ $X2=3.415 $Y2=1.485
r60 17 23 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.57 $Y=1.665
+ $X2=3.57 $Y2=1.485
r61 13 25 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.845 $Y=1.32
+ $X2=3.845 $Y2=1.485
r62 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.845 $Y=1.32
+ $X2=3.845 $Y2=0.74
r63 9 24 16.7191 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.82 $Y=1.65
+ $X2=3.82 $Y2=1.485
r64 9 11 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=3.82 $Y=1.65 $X2=3.82
+ $Y2=2.4
r65 5 20 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.415 $Y=1.32
+ $X2=3.415 $Y2=1.485
r66 5 7 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.415 $Y=1.32
+ $X2=3.415 $Y2=0.74
r67 1 19 16.7191 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.37 $Y=1.65
+ $X2=3.37 $Y2=1.485
r68 1 3 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=3.37 $Y=1.65 $X2=3.37
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_2%B1 3 7 11 15 17 18 28
c41 7 0 3.50294e-19 $X=4.275 $Y=0.74
c42 3 0 1.47716e-19 $X=4.27 $Y=2.4
r43 27 28 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.705 $Y=1.515
+ $X2=4.72 $Y2=1.515
r44 25 27 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=4.345 $Y=1.515
+ $X2=4.705 $Y2=1.515
r45 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.345
+ $Y=1.515 $X2=4.345 $Y2=1.515
r46 23 25 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=4.275 $Y=1.515
+ $X2=4.345 $Y2=1.515
r47 21 23 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=4.27 $Y=1.515
+ $X2=4.275 $Y2=1.515
r48 18 26 5.76222 $w=4.28e-07 $l=2.15e-07 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.345 $Y2=1.565
r49 17 26 7.10226 $w=4.28e-07 $l=2.65e-07 $layer=LI1_cond $X=4.08 $Y=1.565
+ $X2=4.345 $Y2=1.565
r50 13 28 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.72 $Y=1.68
+ $X2=4.72 $Y2=1.515
r51 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.72 $Y=1.68
+ $X2=4.72 $Y2=2.4
r52 9 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.705 $Y=1.35
+ $X2=4.705 $Y2=1.515
r53 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.705 $Y=1.35
+ $X2=4.705 $Y2=0.74
r54 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.275 $Y=1.35
+ $X2=4.275 $Y2=1.515
r55 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.275 $Y=1.35
+ $X2=4.275 $Y2=0.74
r56 1 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.27 $Y=1.68
+ $X2=4.27 $Y2=1.515
r57 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.27 $Y=1.68 $X2=4.27
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_2%VPWR 1 2 3 12 18 22 24 26 31 39 46 47 50
+ 53 56
r56 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r57 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r58 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 47 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r60 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r61 44 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.66 $Y=3.33
+ $X2=4.495 $Y2=3.33
r62 44 46 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.66 $Y=3.33
+ $X2=5.04 $Y2=3.33
r63 43 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r64 43 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r65 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r66 40 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=3.33
+ $X2=3.595 $Y2=3.33
r67 40 42 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.76 $Y=3.33 $X2=4.08
+ $Y2=3.33
r68 39 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=3.33
+ $X2=4.495 $Y2=3.33
r69 39 42 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.33 $Y=3.33
+ $X2=4.08 $Y2=3.33
r70 38 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r71 37 38 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r72 35 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r73 34 37 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r74 34 35 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r75 32 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.91 $Y=3.33
+ $X2=0.745 $Y2=3.33
r76 32 34 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.91 $Y=3.33 $X2=1.2
+ $Y2=3.33
r77 31 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.43 $Y=3.33
+ $X2=3.595 $Y2=3.33
r78 31 37 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.43 $Y=3.33
+ $X2=3.12 $Y2=3.33
r79 29 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r80 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r81 26 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.58 $Y=3.33
+ $X2=0.745 $Y2=3.33
r82 26 28 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.58 $Y=3.33
+ $X2=0.24 $Y2=3.33
r83 24 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r84 24 35 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.2 $Y2=3.33
r85 20 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.495 $Y=3.245
+ $X2=4.495 $Y2=3.33
r86 20 22 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=4.495 $Y=3.245
+ $X2=4.495 $Y2=2.455
r87 16 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=3.245
+ $X2=3.595 $Y2=3.33
r88 16 18 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=3.595 $Y=3.245
+ $X2=3.595 $Y2=2.455
r89 12 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.745 $Y=2.105
+ $X2=0.745 $Y2=2.815
r90 10 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=3.245
+ $X2=0.745 $Y2=3.33
r91 10 15 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.745 $Y=3.245
+ $X2=0.745 $Y2=2.815
r92 3 22 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=4.36
+ $Y=1.84 $X2=4.495 $Y2=2.455
r93 2 18 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=3.46
+ $Y=1.84 $X2=3.595 $Y2=2.455
r94 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.96 $X2=0.745 $Y2=2.815
r95 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.96 $X2=0.745 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_2%A_424_368# 1 2 3 4 15 19 20 21 24 25 29 31
+ 33 35 40
c56 29 0 2.95431e-19 $X=4.045 $Y=2.815
c57 21 0 1.0233e-19 $X=3.105 $Y=2.12
r58 33 42 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=4.985 $Y=2.12
+ $X2=4.985 $Y2=1.97
r59 33 35 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=4.985 $Y=2.12
+ $X2=4.985 $Y2=2.4
r60 32 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=2.035
+ $X2=4.045 $Y2=2.035
r61 31 42 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=4.86 $Y=2.035
+ $X2=4.985 $Y2=1.97
r62 31 32 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.86 $Y=2.035
+ $X2=4.13 $Y2=2.035
r63 27 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.045 $Y=2.12
+ $X2=4.045 $Y2=2.035
r64 27 29 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.045 $Y=2.12
+ $X2=4.045 $Y2=2.815
r65 26 38 3.99177 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=3.23 $Y=2.035
+ $X2=3.105 $Y2=1.97
r66 25 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.96 $Y=2.035
+ $X2=4.045 $Y2=2.035
r67 25 26 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.96 $Y=2.035
+ $X2=3.23 $Y2=2.035
r68 22 24 23.2793 $w=2.48e-07 $l=5.05e-07 $layer=LI1_cond $X=3.105 $Y=2.905
+ $X2=3.105 $Y2=2.4
r69 21 38 3.1514 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=3.105 $Y=2.12
+ $X2=3.105 $Y2=1.97
r70 21 24 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=3.105 $Y=2.12
+ $X2=3.105 $Y2=2.4
r71 19 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.98 $Y=2.99
+ $X2=3.105 $Y2=2.905
r72 19 20 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.98 $Y=2.99
+ $X2=2.33 $Y2=2.99
r73 15 18 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=2.205 $Y=1.985
+ $X2=2.205 $Y2=2.815
r74 13 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.205 $Y=2.905
+ $X2=2.33 $Y2=2.99
r75 13 18 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=2.205 $Y=2.905
+ $X2=2.205 $Y2=2.815
r76 4 42 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.81
+ $Y=1.84 $X2=4.945 $Y2=1.985
r77 4 35 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=4.81
+ $Y=1.84 $X2=4.945 $Y2=2.4
r78 3 40 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=3.91
+ $Y=1.84 $X2=4.045 $Y2=2.115
r79 3 29 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.91
+ $Y=1.84 $X2=4.045 $Y2=2.815
r80 2 38 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.01
+ $Y=1.84 $X2=3.145 $Y2=1.985
r81 2 24 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=3.01
+ $Y=1.84 $X2=3.145 $Y2=2.4
r82 1 18 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=2.12
+ $Y=1.84 $X2=2.245 $Y2=2.815
r83 1 15 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.12
+ $Y=1.84 $X2=2.245 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_2%Y 1 2 3 12 14 15 18 20 22 25 29 30 37
c57 25 0 5.94286e-20 $X=3.63 $Y=0.95
c58 22 0 2.40437e-20 $X=3.465 $Y=1.065
r59 30 37 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=1.195
+ $X2=3.235 $Y2=1.195
r60 25 27 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.63 $Y=0.95
+ $X2=3.63 $Y2=1.065
r61 22 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.465 $Y=1.065
+ $X2=3.63 $Y2=1.065
r62 22 37 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.465 $Y=1.065
+ $X2=3.235 $Y2=1.065
r63 21 29 4.50329 $w=3e-07 $l=1.28e-07 $layer=LI1_cond $X=2.78 $Y=1.195
+ $X2=2.652 $Y2=1.195
r64 20 30 2.6801 $w=4.28e-07 $l=1e-07 $layer=LI1_cond $X=3.02 $Y=1.195 $X2=3.12
+ $Y2=1.195
r65 20 21 6.43224 $w=4.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.02 $Y=1.195
+ $X2=2.78 $Y2=1.195
r66 16 29 1.93381 $w=2.55e-07 $l=2.15e-07 $layer=LI1_cond $X=2.652 $Y=1.41
+ $X2=2.652 $Y2=1.195
r67 16 18 25.9865 $w=2.53e-07 $l=5.75e-07 $layer=LI1_cond $X=2.652 $Y=1.41
+ $X2=2.652 $Y2=1.985
r68 14 29 4.50329 $w=3e-07 $l=1.82784e-07 $layer=LI1_cond $X=2.525 $Y=1.065
+ $X2=2.652 $Y2=1.195
r69 14 15 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.525 $Y=1.065
+ $X2=2.25 $Y2=1.065
r70 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.165 $Y=0.98
+ $X2=2.25 $Y2=1.065
r71 10 12 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.165 $Y=0.98
+ $X2=2.165 $Y2=0.555
r72 3 18 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.56
+ $Y=1.84 $X2=2.695 $Y2=1.985
r73 2 25 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=3.49
+ $Y=0.37 $X2=3.63 $Y2=0.95
r74 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.025
+ $Y=0.41 $X2=2.165 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_2%VGND 1 2 3 4 15 19 23 27 30 31 32 34 39 44
+ 57 58 61 64 67
r77 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r78 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r79 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r80 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r81 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r82 52 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r83 51 54 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r84 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r85 49 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.76 $Y=0 $X2=2.595
+ $Y2=0
r86 49 51 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.76 $Y=0 $X2=3.12
+ $Y2=0
r87 48 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r88 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r89 45 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.9 $Y=0 $X2=1.735
+ $Y2=0
r90 45 47 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.9 $Y=0 $X2=2.16
+ $Y2=0
r91 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.43 $Y=0 $X2=2.595
+ $Y2=0
r92 44 47 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.43 $Y=0 $X2=2.16
+ $Y2=0
r93 43 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r94 43 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r95 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r96 40 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.73
+ $Y2=0
r97 40 42 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r98 39 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.57 $Y=0 $X2=1.735
+ $Y2=0
r99 39 42 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.57 $Y=0 $X2=1.2
+ $Y2=0
r100 37 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r101 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r102 34 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.73
+ $Y2=0
r103 34 36 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.605 $Y=0
+ $X2=0.24 $Y2=0
r104 32 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r105 32 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r106 32 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r107 30 54 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.325 $Y=0 $X2=4.08
+ $Y2=0
r108 30 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.325 $Y=0 $X2=4.45
+ $Y2=0
r109 29 57 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=4.575 $Y=0
+ $X2=5.04 $Y2=0
r110 29 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.575 $Y=0 $X2=4.45
+ $Y2=0
r111 25 31 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.45 $Y=0.085
+ $X2=4.45 $Y2=0
r112 25 27 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=4.45 $Y=0.085
+ $X2=4.45 $Y2=0.595
r113 21 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=0.085
+ $X2=2.595 $Y2=0
r114 21 23 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=2.595 $Y=0.085
+ $X2=2.595 $Y2=0.645
r115 17 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.735 $Y=0.085
+ $X2=1.735 $Y2=0
r116 17 19 23.0489 $w=3.28e-07 $l=6.6e-07 $layer=LI1_cond $X=1.735 $Y=0.085
+ $X2=1.735 $Y2=0.745
r117 13 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r118 13 15 26.7367 $w=2.48e-07 $l=5.8e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.665
r119 4 27 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=4.35
+ $Y=0.37 $X2=4.49 $Y2=0.595
r120 3 23 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=2.455
+ $Y=0.41 $X2=2.595 $Y2=0.645
r121 2 19 182 $w=1.7e-07 $l=3.19726e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.51 $X2=1.735 $Y2=0.745
r122 1 15 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.645
+ $Y=0.51 $X2=0.77 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_MS__A2BB2OI_2%A_615_74# 1 2 3 10 14 18 19 22
c34 14 0 1.6164e-19 $X=4.06 $Y=0.6
r35 20 22 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=4.92 $Y=1.01
+ $X2=4.92 $Y2=0.515
r36 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.755 $Y=1.095
+ $X2=4.92 $Y2=1.01
r37 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.755 $Y=1.095
+ $X2=4.145 $Y2=1.095
r38 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.06 $Y=1.01
+ $X2=4.145 $Y2=1.095
r39 15 17 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.06 $Y=1.01
+ $X2=4.06 $Y2=0.965
r40 14 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.06 $Y=0.6 $X2=4.06
+ $Y2=0.475
r41 14 17 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.06 $Y=0.6
+ $X2=4.06 $Y2=0.965
r42 10 25 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.975 $Y=0.475
+ $X2=4.06 $Y2=0.475
r43 10 12 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=3.975 $Y=0.475
+ $X2=3.2 $Y2=0.475
r44 3 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.78
+ $Y=0.37 $X2=4.92 $Y2=0.515
r45 2 25 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.92
+ $Y=0.37 $X2=4.06 $Y2=0.515
r46 2 17 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=3.92
+ $Y=0.37 $X2=4.06 $Y2=0.965
r47 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.075
+ $Y=0.37 $X2=3.2 $Y2=0.515
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and3_2 A B C VGND VNB VPB VPWR X
M1000 X a_41_384# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.368e+11p pd=2.12e+06u as=6.9565e+11p ps=5.12e+06u
M1001 X a_41_384# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.2592e+12p ps=8.72e+06u
M1002 VPWR a_41_384# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND C a_247_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1004 a_247_136# B a_133_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.688e+11p ps=2.12e+06u
M1005 a_133_136# A a_41_384# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1006 VPWR A a_41_384# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=4.62e+11p ps=4.46e+06u
M1007 a_41_384# B VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR C a_41_384# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_41_384# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

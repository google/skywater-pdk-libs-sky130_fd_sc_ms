* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o2bb2ai_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_857_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_857_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 Y a_117_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 Y a_117_368# a_857_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VPWR A1_N a_117_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 VGND A1_N a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_857_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VPWR A2_N a_117_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 Y a_117_368# a_857_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 VPWR A2_N a_117_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X10 VGND A1_N a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 a_117_368# A2_N a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 a_1215_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X13 VPWR a_117_368# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X14 a_1215_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 a_27_74# A2_N a_117_368# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 Y a_117_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X17 a_1215_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X18 a_1215_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X19 a_117_368# A1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X20 VPWR B1 a_1215_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X21 a_857_74# a_117_368# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 a_117_368# A1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X23 a_117_368# A2_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X24 a_27_74# A2_N a_117_368# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 VGND B2 a_857_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 VGND B2 a_857_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 a_117_368# A2_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X28 Y B2 a_1215_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X29 a_117_368# A2_N a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X30 a_857_74# a_117_368# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X31 Y B2 a_1215_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X32 a_27_74# A1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X33 VGND B1 a_857_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X34 VGND B1 a_857_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X35 VPWR A1_N a_117_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X36 VPWR a_117_368# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X37 VPWR B1 a_1215_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X38 a_27_74# A1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X39 a_857_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

* File: sky130_fd_sc_ms__a2111o_2.pxi.spice
* Created: Fri Aug 28 16:55:31 2020
* 
x_PM_SKY130_FD_SC_MS__A2111O_2%A_91_244# N_A_91_244#_M1013_s N_A_91_244#_M1003_d
+ N_A_91_244#_M1011_d N_A_91_244#_M1001_s N_A_91_244#_M1004_g N_A_91_244#_c_87_n
+ N_A_91_244#_M1008_g N_A_91_244#_M1005_g N_A_91_244#_c_89_n N_A_91_244#_M1009_g
+ N_A_91_244#_c_90_n N_A_91_244#_c_91_n N_A_91_244#_c_92_n N_A_91_244#_c_104_n
+ N_A_91_244#_c_105_n N_A_91_244#_c_106_n N_A_91_244#_c_107_n N_A_91_244#_c_93_n
+ N_A_91_244#_c_94_n N_A_91_244#_c_95_n N_A_91_244#_c_96_n N_A_91_244#_c_97_n
+ N_A_91_244#_c_98_n N_A_91_244#_c_99_n N_A_91_244#_c_100_n
+ PM_SKY130_FD_SC_MS__A2111O_2%A_91_244#
x_PM_SKY130_FD_SC_MS__A2111O_2%D1 N_D1_M1001_g N_D1_M1013_g D1 D1 N_D1_c_204_n
+ PM_SKY130_FD_SC_MS__A2111O_2%D1
x_PM_SKY130_FD_SC_MS__A2111O_2%C1 N_C1_M1006_g N_C1_M1003_g C1 C1 C1 C1
+ N_C1_c_240_n N_C1_c_241_n PM_SKY130_FD_SC_MS__A2111O_2%C1
x_PM_SKY130_FD_SC_MS__A2111O_2%B1 N_B1_M1012_g N_B1_M1000_g B1 N_B1_c_280_n
+ N_B1_c_281_n PM_SKY130_FD_SC_MS__A2111O_2%B1
x_PM_SKY130_FD_SC_MS__A2111O_2%A2 N_A2_M1002_g N_A2_M1010_g A2 A2 N_A2_c_319_n
+ PM_SKY130_FD_SC_MS__A2111O_2%A2
x_PM_SKY130_FD_SC_MS__A2111O_2%A1 N_A1_M1011_g N_A1_M1007_g N_A1_c_354_n A1
+ N_A1_c_355_n N_A1_c_356_n PM_SKY130_FD_SC_MS__A2111O_2%A1
x_PM_SKY130_FD_SC_MS__A2111O_2%VPWR N_VPWR_M1004_s N_VPWR_M1005_s N_VPWR_M1002_d
+ N_VPWR_c_384_n N_VPWR_c_385_n N_VPWR_c_386_n N_VPWR_c_387_n N_VPWR_c_388_n
+ N_VPWR_c_389_n VPWR N_VPWR_c_390_n N_VPWR_c_391_n N_VPWR_c_383_n
+ N_VPWR_c_393_n PM_SKY130_FD_SC_MS__A2111O_2%VPWR
x_PM_SKY130_FD_SC_MS__A2111O_2%X N_X_M1008_s N_X_M1004_d N_X_c_436_n X X X X X
+ PM_SKY130_FD_SC_MS__A2111O_2%X
x_PM_SKY130_FD_SC_MS__A2111O_2%A_633_368# N_A_633_368#_M1000_d
+ N_A_633_368#_M1007_d N_A_633_368#_c_459_n N_A_633_368#_c_456_n
+ N_A_633_368#_c_467_n N_A_633_368#_c_457_n N_A_633_368#_c_458_n
+ PM_SKY130_FD_SC_MS__A2111O_2%A_633_368#
x_PM_SKY130_FD_SC_MS__A2111O_2%VGND N_VGND_M1008_d N_VGND_M1009_d N_VGND_M1013_d
+ N_VGND_M1012_d N_VGND_c_484_n N_VGND_c_485_n N_VGND_c_486_n N_VGND_c_487_n
+ N_VGND_c_488_n N_VGND_c_489_n N_VGND_c_490_n VGND N_VGND_c_491_n
+ N_VGND_c_492_n N_VGND_c_493_n N_VGND_c_494_n N_VGND_c_495_n N_VGND_c_496_n
+ PM_SKY130_FD_SC_MS__A2111O_2%VGND
cc_1 VNB N_A_91_244#_M1004_g 0.00871317f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_2 VNB N_A_91_244#_c_87_n 0.021272f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.22
cc_3 VNB N_A_91_244#_M1005_g 0.00630758f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.4
cc_4 VNB N_A_91_244#_c_89_n 0.0189136f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=1.22
cc_5 VNB N_A_91_244#_c_90_n 0.0144821f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=1.55
cc_6 VNB N_A_91_244#_c_91_n 0.00164528f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=1.95
cc_7 VNB N_A_91_244#_c_92_n 0.0247935f $X=-0.19 $Y=-0.245 $X2=1.78 $Y2=1.095
cc_8 VNB N_A_91_244#_c_93_n 0.0159334f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=0.515
cc_9 VNB N_A_91_244#_c_94_n 0.00754392f $X=-0.19 $Y=-0.245 $X2=2.76 $Y2=1.095
cc_10 VNB N_A_91_244#_c_95_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=0.515
cc_11 VNB N_A_91_244#_c_96_n 0.0208031f $X=-0.19 $Y=-0.245 $X2=4.19 $Y2=1.095
cc_12 VNB N_A_91_244#_c_97_n 0.0281813f $X=-0.19 $Y=-0.245 $X2=4.355 $Y2=0.515
cc_13 VNB N_A_91_244#_c_98_n 0.0802753f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=1.385
cc_14 VNB N_A_91_244#_c_99_n 0.00237125f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.095
cc_15 VNB N_A_91_244#_c_100_n 0.0086793f $X=-0.19 $Y=-0.245 $X2=2.885 $Y2=1.095
cc_16 VNB N_D1_M1013_g 0.0327351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB D1 0.00943624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_D1_c_204_n 0.0257661f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_19 VNB N_C1_M1003_g 0.0238646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_C1_c_240_n 0.0262087f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_21 VNB N_C1_c_241_n 0.00167125f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_22 VNB N_B1_M1012_g 0.0272326f $X=-0.19 $Y=-0.245 $X2=4.215 $Y2=0.37
cc_23 VNB N_B1_c_280_n 0.0262412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B1_c_281_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.55
cc_25 VNB N_A2_M1010_g 0.0254699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB A2 0.00423229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A2_c_319_n 0.021856f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_28 VNB N_A1_M1011_g 0.0321165f $X=-0.19 $Y=-0.245 $X2=4.215 $Y2=0.37
cc_29 VNB N_A1_c_354_n 0.00984469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A1_c_355_n 0.0439496f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_31 VNB N_A1_c_356_n 0.00813406f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_32 VNB N_VPWR_c_383_n 0.203486f $X=-0.19 $Y=-0.245 $X2=2.885 $Y2=1.01
cc_33 VNB N_X_c_436_n 0.00350677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB X 8.01576e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_484_n 0.0141006f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.55
cc_36 VNB N_VGND_c_485_n 0.0502297f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.4
cc_37 VNB N_VGND_c_486_n 0.016021f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.74
cc_38 VNB N_VGND_c_487_n 0.00333244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_488_n 0.00790127f $X=-0.19 $Y=-0.245 $X2=1.275 $Y2=1.55
cc_40 VNB N_VGND_c_489_n 0.0245715f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=1.095
cc_41 VNB N_VGND_c_490_n 0.00677473f $X=-0.19 $Y=-0.245 $X2=1.755 $Y2=2.035
cc_42 VNB N_VGND_c_491_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=2.815
cc_43 VNB N_VGND_c_492_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=2.885 $Y2=1.01
cc_44 VNB N_VGND_c_493_n 0.0334725f $X=-0.19 $Y=-0.245 $X2=4.355 $Y2=1.01
cc_45 VNB N_VGND_c_494_n 0.302009f $X=-0.19 $Y=-0.245 $X2=4.355 $Y2=0.515
cc_46 VNB N_VGND_c_495_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=1.385
cc_47 VNB N_VGND_c_496_n 0.0103896f $X=-0.19 $Y=-0.245 $X2=1.905 $Y2=1.095
cc_48 VPB N_A_91_244#_M1004_g 0.0274058f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_49 VPB N_A_91_244#_M1005_g 0.0247066f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=2.4
cc_50 VPB N_A_91_244#_c_91_n 0.00560051f $X=-0.19 $Y=1.66 $X2=1.275 $Y2=1.95
cc_51 VPB N_A_91_244#_c_104_n 0.0241081f $X=-0.19 $Y=1.66 $X2=1.755 $Y2=2.035
cc_52 VPB N_A_91_244#_c_105_n 2.25523e-19 $X=-0.19 $Y=1.66 $X2=1.36 $Y2=2.035
cc_53 VPB N_A_91_244#_c_106_n 6.27129e-19 $X=-0.19 $Y=1.66 $X2=1.92 $Y2=2.12
cc_54 VPB N_A_91_244#_c_107_n 0.0137435f $X=-0.19 $Y=1.66 $X2=1.92 $Y2=2.815
cc_55 VPB N_D1_M1001_g 0.024618f $X=-0.19 $Y=1.66 $X2=4.215 $Y2=0.37
cc_56 VPB D1 0.00846085f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_D1_c_204_n 0.00576404f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_58 VPB N_C1_M1006_g 0.0217532f $X=-0.19 $Y=1.66 $X2=4.215 $Y2=0.37
cc_59 VPB N_C1_c_240_n 0.00561973f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_60 VPB N_C1_c_241_n 0.00130499f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_61 VPB N_B1_M1000_g 0.0236127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_B1_c_280_n 0.00562372f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_B1_c_281_n 0.00199771f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.55
cc_64 VPB N_A2_M1002_g 0.0223054f $X=-0.19 $Y=1.66 $X2=4.215 $Y2=0.37
cc_65 VPB A2 0.00451479f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A2_c_319_n 0.00538829f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_67 VPB N_A1_M1007_g 0.0281996f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_A1_c_354_n 5.8517e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_A1_c_355_n 0.0145157f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_70 VPB N_A1_c_356_n 0.0117191f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_71 VPB N_VPWR_c_384_n 0.011928f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_385_n 0.0646893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_386_n 0.0148803f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.74
cc_74 VPB N_VPWR_c_387_n 0.0067963f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=2.4
cc_75 VPB N_VPWR_c_388_n 0.0650536f $X=-0.19 $Y=1.66 $X2=0.99 $Y2=0.74
cc_76 VPB N_VPWR_c_389_n 0.00689679f $X=-0.19 $Y=1.66 $X2=0.99 $Y2=0.74
cc_77 VPB N_VPWR_c_390_n 0.0184862f $X=-0.19 $Y=1.66 $X2=1.78 $Y2=1.095
cc_78 VPB N_VPWR_c_391_n 0.0236066f $X=-0.19 $Y=1.66 $X2=2.03 $Y2=1.095
cc_79 VPB N_VPWR_c_383_n 0.100755f $X=-0.19 $Y=1.66 $X2=2.885 $Y2=1.01
cc_80 VPB N_VPWR_c_393_n 0.0061274f $X=-0.19 $Y=1.66 $X2=4.355 $Y2=1.01
cc_81 VPB X 0.00342209f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_633_368#_c_456_n 0.00312968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_A_633_368#_c_457_n 0.00743317f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=1.55
cc_84 VPB N_A_633_368#_c_458_n 0.0358769f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.4
cc_85 N_A_91_244#_c_91_n N_D1_M1001_g 0.00343373f $X=1.275 $Y=1.95 $X2=0 $Y2=0
cc_86 N_A_91_244#_c_106_n N_D1_M1001_g 0.00300739f $X=1.92 $Y=2.12 $X2=0 $Y2=0
cc_87 N_A_91_244#_c_107_n N_D1_M1001_g 0.0139742f $X=1.92 $Y=2.815 $X2=0 $Y2=0
cc_88 N_A_91_244#_c_93_n N_D1_M1013_g 0.00159319f $X=1.945 $Y=0.515 $X2=0 $Y2=0
cc_89 N_A_91_244#_c_94_n N_D1_M1013_g 0.0140963f $X=2.76 $Y=1.095 $X2=0 $Y2=0
cc_90 N_A_91_244#_c_90_n D1 0.0146967f $X=1.275 $Y=1.55 $X2=0 $Y2=0
cc_91 N_A_91_244#_c_91_n D1 0.0169761f $X=1.275 $Y=1.95 $X2=0 $Y2=0
cc_92 N_A_91_244#_c_92_n D1 0.0173741f $X=1.78 $Y=1.095 $X2=0 $Y2=0
cc_93 N_A_91_244#_c_104_n D1 0.0153495f $X=1.755 $Y=2.035 $X2=0 $Y2=0
cc_94 N_A_91_244#_c_106_n D1 0.0264311f $X=1.92 $Y=2.12 $X2=0 $Y2=0
cc_95 N_A_91_244#_c_94_n D1 0.0183652f $X=2.76 $Y=1.095 $X2=0 $Y2=0
cc_96 N_A_91_244#_c_98_n D1 9.56934e-19 $X=1.195 $Y=1.385 $X2=0 $Y2=0
cc_97 N_A_91_244#_c_99_n D1 0.0220075f $X=1.905 $Y=1.095 $X2=0 $Y2=0
cc_98 N_A_91_244#_c_91_n N_D1_c_204_n 4.43363e-19 $X=1.275 $Y=1.95 $X2=0 $Y2=0
cc_99 N_A_91_244#_c_106_n N_D1_c_204_n 7.81657e-19 $X=1.92 $Y=2.12 $X2=0 $Y2=0
cc_100 N_A_91_244#_c_94_n N_D1_c_204_n 0.00134913f $X=2.76 $Y=1.095 $X2=0 $Y2=0
cc_101 N_A_91_244#_c_98_n N_D1_c_204_n 0.0033277f $X=1.195 $Y=1.385 $X2=0 $Y2=0
cc_102 N_A_91_244#_c_99_n N_D1_c_204_n 0.00291196f $X=1.905 $Y=1.095 $X2=0 $Y2=0
cc_103 N_A_91_244#_c_106_n N_C1_M1006_g 4.24617e-19 $X=1.92 $Y=2.12 $X2=0 $Y2=0
cc_104 N_A_91_244#_c_107_n N_C1_M1006_g 0.00236546f $X=1.92 $Y=2.815 $X2=0 $Y2=0
cc_105 N_A_91_244#_c_94_n N_C1_M1003_g 0.0132453f $X=2.76 $Y=1.095 $X2=0 $Y2=0
cc_106 N_A_91_244#_c_95_n N_C1_M1003_g 3.97481e-19 $X=2.845 $Y=0.515 $X2=0 $Y2=0
cc_107 N_A_91_244#_c_94_n N_C1_c_240_n 0.00114367f $X=2.76 $Y=1.095 $X2=0 $Y2=0
cc_108 N_A_91_244#_c_106_n N_C1_c_241_n 0.00741114f $X=1.92 $Y=2.12 $X2=0 $Y2=0
cc_109 N_A_91_244#_c_107_n N_C1_c_241_n 0.0316148f $X=1.92 $Y=2.815 $X2=0 $Y2=0
cc_110 N_A_91_244#_c_94_n N_C1_c_241_n 0.0244947f $X=2.76 $Y=1.095 $X2=0 $Y2=0
cc_111 N_A_91_244#_c_100_n N_C1_c_241_n 0.00124816f $X=2.885 $Y=1.095 $X2=0
+ $Y2=0
cc_112 N_A_91_244#_c_95_n N_B1_M1012_g 0.00979642f $X=2.845 $Y=0.515 $X2=0 $Y2=0
cc_113 N_A_91_244#_c_96_n N_B1_M1012_g 0.0123033f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_114 N_A_91_244#_c_100_n N_B1_M1012_g 0.00154264f $X=2.885 $Y=1.095 $X2=0
+ $Y2=0
cc_115 N_A_91_244#_c_96_n N_B1_c_280_n 0.00125903f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_116 N_A_91_244#_c_96_n N_B1_c_281_n 0.0229301f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_117 N_A_91_244#_c_100_n N_B1_c_281_n 0.00196319f $X=2.885 $Y=1.095 $X2=0
+ $Y2=0
cc_118 N_A_91_244#_c_95_n N_A2_M1010_g 9.95982e-19 $X=2.845 $Y=0.515 $X2=0 $Y2=0
cc_119 N_A_91_244#_c_96_n N_A2_M1010_g 0.0149964f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_120 N_A_91_244#_c_97_n N_A2_M1010_g 0.00218322f $X=4.355 $Y=0.515 $X2=0 $Y2=0
cc_121 N_A_91_244#_c_96_n A2 0.0544915f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_122 N_A_91_244#_c_96_n N_A2_c_319_n 0.00474488f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_123 N_A_91_244#_c_96_n N_A1_M1011_g 0.0135439f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_124 N_A_91_244#_c_97_n N_A1_M1011_g 0.0125612f $X=4.355 $Y=0.515 $X2=0 $Y2=0
cc_125 N_A_91_244#_c_96_n N_A1_c_354_n 0.00680871f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_126 N_A_91_244#_c_96_n N_A1_c_355_n 0.00121887f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_127 N_A_91_244#_c_96_n N_A1_c_356_n 0.0132907f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_128 N_A_91_244#_c_91_n N_VPWR_M1005_s 0.00210234f $X=1.275 $Y=1.95 $X2=0
+ $Y2=0
cc_129 N_A_91_244#_c_105_n N_VPWR_M1005_s 0.00503276f $X=1.36 $Y=2.035 $X2=0
+ $Y2=0
cc_130 N_A_91_244#_M1004_g N_VPWR_c_385_n 0.00517389f $X=0.545 $Y=2.4 $X2=0
+ $Y2=0
cc_131 N_A_91_244#_M1004_g N_VPWR_c_386_n 5.65601e-19 $X=0.545 $Y=2.4 $X2=0
+ $Y2=0
cc_132 N_A_91_244#_M1005_g N_VPWR_c_386_n 0.0149818f $X=0.995 $Y=2.4 $X2=0 $Y2=0
cc_133 N_A_91_244#_c_104_n N_VPWR_c_386_n 0.00198924f $X=1.755 $Y=2.035 $X2=0
+ $Y2=0
cc_134 N_A_91_244#_c_105_n N_VPWR_c_386_n 0.0152886f $X=1.36 $Y=2.035 $X2=0
+ $Y2=0
cc_135 N_A_91_244#_c_107_n N_VPWR_c_386_n 0.033566f $X=1.92 $Y=2.815 $X2=0 $Y2=0
cc_136 N_A_91_244#_c_107_n N_VPWR_c_388_n 0.014549f $X=1.92 $Y=2.815 $X2=0 $Y2=0
cc_137 N_A_91_244#_M1004_g N_VPWR_c_390_n 0.005209f $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_138 N_A_91_244#_M1005_g N_VPWR_c_390_n 0.00460063f $X=0.995 $Y=2.4 $X2=0
+ $Y2=0
cc_139 N_A_91_244#_M1004_g N_VPWR_c_383_n 0.00986139f $X=0.545 $Y=2.4 $X2=0
+ $Y2=0
cc_140 N_A_91_244#_M1005_g N_VPWR_c_383_n 0.00908554f $X=0.995 $Y=2.4 $X2=0
+ $Y2=0
cc_141 N_A_91_244#_c_107_n N_VPWR_c_383_n 0.0119743f $X=1.92 $Y=2.815 $X2=0
+ $Y2=0
cc_142 N_A_91_244#_c_87_n N_X_c_436_n 0.00267578f $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_143 N_A_91_244#_c_89_n N_X_c_436_n 0.00139568f $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_144 N_A_91_244#_c_90_n N_X_c_436_n 0.0319992f $X=1.275 $Y=1.55 $X2=0 $Y2=0
cc_145 N_A_91_244#_c_98_n N_X_c_436_n 0.0251153f $X=1.195 $Y=1.385 $X2=0 $Y2=0
cc_146 N_A_91_244#_M1004_g X 0.029482f $X=0.545 $Y=2.4 $X2=0 $Y2=0
cc_147 N_A_91_244#_M1005_g X 0.00324126f $X=0.995 $Y=2.4 $X2=0 $Y2=0
cc_148 N_A_91_244#_c_91_n X 0.016544f $X=1.275 $Y=1.95 $X2=0 $Y2=0
cc_149 N_A_91_244#_c_98_n X 0.00657588f $X=1.195 $Y=1.385 $X2=0 $Y2=0
cc_150 N_A_91_244#_c_90_n N_VGND_M1009_d 0.00288214f $X=1.275 $Y=1.55 $X2=0
+ $Y2=0
cc_151 N_A_91_244#_c_94_n N_VGND_M1013_d 0.00218982f $X=2.76 $Y=1.095 $X2=0
+ $Y2=0
cc_152 N_A_91_244#_c_96_n N_VGND_M1012_d 0.0059981f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_153 N_A_91_244#_c_87_n N_VGND_c_485_n 0.0159149f $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_154 N_A_91_244#_c_89_n N_VGND_c_485_n 5.58177e-19 $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_155 N_A_91_244#_c_98_n N_VGND_c_485_n 0.00158354f $X=1.195 $Y=1.385 $X2=0
+ $Y2=0
cc_156 N_A_91_244#_c_87_n N_VGND_c_486_n 4.71636e-19 $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_157 N_A_91_244#_c_89_n N_VGND_c_486_n 0.0128397f $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_158 N_A_91_244#_c_90_n N_VGND_c_486_n 0.020572f $X=1.275 $Y=1.55 $X2=0 $Y2=0
cc_159 N_A_91_244#_c_92_n N_VGND_c_486_n 7.22336e-19 $X=1.78 $Y=1.095 $X2=0
+ $Y2=0
cc_160 N_A_91_244#_c_93_n N_VGND_c_486_n 0.0217548f $X=1.945 $Y=0.515 $X2=0
+ $Y2=0
cc_161 N_A_91_244#_c_98_n N_VGND_c_486_n 0.00147764f $X=1.195 $Y=1.385 $X2=0
+ $Y2=0
cc_162 N_A_91_244#_c_93_n N_VGND_c_487_n 0.0186004f $X=1.945 $Y=0.515 $X2=0
+ $Y2=0
cc_163 N_A_91_244#_c_94_n N_VGND_c_487_n 0.020332f $X=2.76 $Y=1.095 $X2=0 $Y2=0
cc_164 N_A_91_244#_c_95_n N_VGND_c_487_n 0.0186004f $X=2.845 $Y=0.515 $X2=0
+ $Y2=0
cc_165 N_A_91_244#_c_95_n N_VGND_c_488_n 0.018474f $X=2.845 $Y=0.515 $X2=0 $Y2=0
cc_166 N_A_91_244#_c_96_n N_VGND_c_488_n 0.0389277f $X=4.19 $Y=1.095 $X2=0 $Y2=0
cc_167 N_A_91_244#_c_97_n N_VGND_c_488_n 0.01706f $X=4.355 $Y=0.515 $X2=0 $Y2=0
cc_168 N_A_91_244#_c_93_n N_VGND_c_489_n 0.011066f $X=1.945 $Y=0.515 $X2=0 $Y2=0
cc_169 N_A_91_244#_c_87_n N_VGND_c_491_n 0.00383152f $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_170 N_A_91_244#_c_89_n N_VGND_c_491_n 0.00383152f $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_171 N_A_91_244#_c_95_n N_VGND_c_492_n 0.0109942f $X=2.845 $Y=0.515 $X2=0
+ $Y2=0
cc_172 N_A_91_244#_c_97_n N_VGND_c_493_n 0.0145639f $X=4.355 $Y=0.515 $X2=0
+ $Y2=0
cc_173 N_A_91_244#_c_87_n N_VGND_c_494_n 0.0075754f $X=0.56 $Y=1.22 $X2=0 $Y2=0
cc_174 N_A_91_244#_c_89_n N_VGND_c_494_n 0.0075754f $X=0.99 $Y=1.22 $X2=0 $Y2=0
cc_175 N_A_91_244#_c_93_n N_VGND_c_494_n 0.00915947f $X=1.945 $Y=0.515 $X2=0
+ $Y2=0
cc_176 N_A_91_244#_c_95_n N_VGND_c_494_n 0.00904371f $X=2.845 $Y=0.515 $X2=0
+ $Y2=0
cc_177 N_A_91_244#_c_97_n N_VGND_c_494_n 0.0119984f $X=4.355 $Y=0.515 $X2=0
+ $Y2=0
cc_178 N_A_91_244#_c_96_n A_771_74# 0.00366293f $X=4.19 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_179 N_D1_M1001_g N_C1_M1006_g 0.0519644f $X=2.145 $Y=2.4 $X2=0 $Y2=0
cc_180 N_D1_M1013_g N_C1_M1003_g 0.0281796f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_181 D1 N_C1_c_240_n 0.00257845f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_182 N_D1_c_204_n N_C1_c_240_n 0.0519644f $X=2.07 $Y=1.515 $X2=0 $Y2=0
cc_183 N_D1_M1001_g N_C1_c_241_n 0.00445369f $X=2.145 $Y=2.4 $X2=0 $Y2=0
cc_184 D1 N_C1_c_241_n 0.0361869f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_185 N_D1_c_204_n N_C1_c_241_n 4.92305e-19 $X=2.07 $Y=1.515 $X2=0 $Y2=0
cc_186 N_D1_M1001_g N_VPWR_c_386_n 0.00395159f $X=2.145 $Y=2.4 $X2=0 $Y2=0
cc_187 N_D1_M1001_g N_VPWR_c_388_n 0.005209f $X=2.145 $Y=2.4 $X2=0 $Y2=0
cc_188 N_D1_M1001_g N_VPWR_c_383_n 0.00988003f $X=2.145 $Y=2.4 $X2=0 $Y2=0
cc_189 N_D1_M1013_g N_VGND_c_487_n 0.0140324f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_190 N_D1_M1013_g N_VGND_c_489_n 0.00383152f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_191 N_D1_M1013_g N_VGND_c_494_n 0.00762539f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_192 N_C1_M1003_g N_B1_M1012_g 0.0195038f $X=2.63 $Y=0.74 $X2=0 $Y2=0
cc_193 N_C1_M1006_g N_B1_M1000_g 0.0432729f $X=2.535 $Y=2.4 $X2=0 $Y2=0
cc_194 N_C1_c_241_n N_B1_M1000_g 0.0127978f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_195 N_C1_c_240_n N_B1_c_280_n 0.0201104f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_196 N_C1_c_241_n N_B1_c_280_n 0.00114936f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_197 N_C1_c_240_n N_B1_c_281_n 0.00114936f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_198 N_C1_c_241_n N_B1_c_281_n 0.0276388f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_199 N_C1_M1006_g N_VPWR_c_388_n 0.00365007f $X=2.535 $Y=2.4 $X2=0 $Y2=0
cc_200 N_C1_c_241_n N_VPWR_c_388_n 0.00925382f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_201 N_C1_M1006_g N_VPWR_c_383_n 0.00443968f $X=2.535 $Y=2.4 $X2=0 $Y2=0
cc_202 N_C1_c_241_n N_VPWR_c_383_n 0.0105443f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_203 N_C1_c_241_n A_525_368# 0.0138299f $X=2.61 $Y=1.515 $X2=-0.19 $Y2=-0.245
cc_204 N_C1_c_241_n N_A_633_368#_c_459_n 0.00784414f $X=2.61 $Y=1.515 $X2=0
+ $Y2=0
cc_205 N_C1_M1006_g N_A_633_368#_c_456_n 0.00107927f $X=2.535 $Y=2.4 $X2=0 $Y2=0
cc_206 N_C1_c_241_n N_A_633_368#_c_456_n 0.0338545f $X=2.61 $Y=1.515 $X2=0 $Y2=0
cc_207 N_C1_M1003_g N_VGND_c_487_n 0.0110514f $X=2.63 $Y=0.74 $X2=0 $Y2=0
cc_208 N_C1_M1003_g N_VGND_c_492_n 0.00383152f $X=2.63 $Y=0.74 $X2=0 $Y2=0
cc_209 N_C1_M1003_g N_VGND_c_494_n 0.00757637f $X=2.63 $Y=0.74 $X2=0 $Y2=0
cc_210 N_B1_M1000_g N_A2_M1002_g 0.0273612f $X=3.075 $Y=2.4 $X2=0 $Y2=0
cc_211 N_B1_c_281_n N_A2_M1002_g 3.34283e-19 $X=3.15 $Y=1.515 $X2=0 $Y2=0
cc_212 N_B1_M1012_g N_A2_M1010_g 0.0187776f $X=3.06 $Y=0.74 $X2=0 $Y2=0
cc_213 N_B1_M1000_g A2 2.9613e-19 $X=3.075 $Y=2.4 $X2=0 $Y2=0
cc_214 N_B1_c_280_n A2 0.00201442f $X=3.15 $Y=1.515 $X2=0 $Y2=0
cc_215 N_B1_c_281_n A2 0.0366314f $X=3.15 $Y=1.515 $X2=0 $Y2=0
cc_216 N_B1_c_280_n N_A2_c_319_n 0.0206382f $X=3.15 $Y=1.515 $X2=0 $Y2=0
cc_217 N_B1_c_281_n N_A2_c_319_n 3.7859e-19 $X=3.15 $Y=1.515 $X2=0 $Y2=0
cc_218 N_B1_M1000_g N_VPWR_c_387_n 6.73475e-19 $X=3.075 $Y=2.4 $X2=0 $Y2=0
cc_219 N_B1_M1000_g N_VPWR_c_388_n 0.005209f $X=3.075 $Y=2.4 $X2=0 $Y2=0
cc_220 N_B1_M1000_g N_VPWR_c_383_n 0.00985168f $X=3.075 $Y=2.4 $X2=0 $Y2=0
cc_221 N_B1_M1000_g N_A_633_368#_c_459_n 0.0030919f $X=3.075 $Y=2.4 $X2=0 $Y2=0
cc_222 N_B1_c_280_n N_A_633_368#_c_459_n 7.74224e-19 $X=3.15 $Y=1.515 $X2=0
+ $Y2=0
cc_223 N_B1_c_281_n N_A_633_368#_c_459_n 0.0130747f $X=3.15 $Y=1.515 $X2=0 $Y2=0
cc_224 N_B1_M1000_g N_A_633_368#_c_456_n 0.0144438f $X=3.075 $Y=2.4 $X2=0 $Y2=0
cc_225 N_B1_M1012_g N_VGND_c_487_n 5.17244e-19 $X=3.06 $Y=0.74 $X2=0 $Y2=0
cc_226 N_B1_M1012_g N_VGND_c_488_n 0.00589272f $X=3.06 $Y=0.74 $X2=0 $Y2=0
cc_227 N_B1_M1012_g N_VGND_c_492_n 0.00434272f $X=3.06 $Y=0.74 $X2=0 $Y2=0
cc_228 N_B1_M1012_g N_VGND_c_494_n 0.0082236f $X=3.06 $Y=0.74 $X2=0 $Y2=0
cc_229 N_A2_M1010_g N_A1_M1011_g 0.0442642f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_230 N_A2_M1002_g N_A1_M1007_g 0.0327166f $X=3.615 $Y=2.4 $X2=0 $Y2=0
cc_231 A2 N_A1_M1007_g 0.00506992f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_232 A2 N_A1_c_354_n 0.0136716f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_233 N_A2_c_319_n N_A1_c_354_n 0.0442642f $X=3.69 $Y=1.515 $X2=0 $Y2=0
cc_234 A2 N_A1_c_356_n 0.0346458f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_235 N_A2_M1002_g N_VPWR_c_387_n 0.0127556f $X=3.615 $Y=2.4 $X2=0 $Y2=0
cc_236 N_A2_M1002_g N_VPWR_c_388_n 0.00460063f $X=3.615 $Y=2.4 $X2=0 $Y2=0
cc_237 N_A2_M1002_g N_VPWR_c_383_n 0.00909457f $X=3.615 $Y=2.4 $X2=0 $Y2=0
cc_238 N_A2_M1002_g N_A_633_368#_c_456_n 0.00510762f $X=3.615 $Y=2.4 $X2=0 $Y2=0
cc_239 N_A2_M1002_g N_A_633_368#_c_467_n 0.0171755f $X=3.615 $Y=2.4 $X2=0 $Y2=0
cc_240 A2 N_A_633_368#_c_467_n 0.0480196f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_241 N_A2_c_319_n N_A_633_368#_c_467_n 7.04415e-19 $X=3.69 $Y=1.515 $X2=0
+ $Y2=0
cc_242 N_A2_M1002_g N_A_633_368#_c_458_n 8.67149e-19 $X=3.615 $Y=2.4 $X2=0 $Y2=0
cc_243 N_A2_M1010_g N_VGND_c_488_n 0.0215908f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A2_M1010_g N_VGND_c_493_n 0.00383152f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_245 N_A2_M1010_g N_VGND_c_494_n 0.0075694f $X=3.78 $Y=0.74 $X2=0 $Y2=0
cc_246 N_A1_M1007_g N_VPWR_c_387_n 0.00741529f $X=4.155 $Y=2.4 $X2=0 $Y2=0
cc_247 N_A1_M1007_g N_VPWR_c_391_n 0.005209f $X=4.155 $Y=2.4 $X2=0 $Y2=0
cc_248 N_A1_M1007_g N_VPWR_c_383_n 0.00986635f $X=4.155 $Y=2.4 $X2=0 $Y2=0
cc_249 N_A1_M1007_g N_A_633_368#_c_467_n 0.013962f $X=4.155 $Y=2.4 $X2=0 $Y2=0
cc_250 N_A1_M1007_g N_A_633_368#_c_457_n 0.00190089f $X=4.155 $Y=2.4 $X2=0 $Y2=0
cc_251 N_A1_c_355_n N_A_633_368#_c_457_n 0.00467488f $X=4.53 $Y=1.515 $X2=0
+ $Y2=0
cc_252 N_A1_c_356_n N_A_633_368#_c_457_n 0.0159673f $X=4.53 $Y=1.515 $X2=0 $Y2=0
cc_253 N_A1_M1007_g N_A_633_368#_c_458_n 0.0119414f $X=4.155 $Y=2.4 $X2=0 $Y2=0
cc_254 N_A1_M1011_g N_VGND_c_488_n 0.00189477f $X=4.14 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A1_M1011_g N_VGND_c_493_n 0.00434272f $X=4.14 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A1_M1011_g N_VGND_c_494_n 0.00824773f $X=4.14 $Y=0.74 $X2=0 $Y2=0
cc_257 N_VPWR_c_385_n X 0.0380882f $X=0.32 $Y=1.985 $X2=0 $Y2=0
cc_258 N_VPWR_c_386_n X 0.0238869f $X=1.22 $Y=2.455 $X2=0 $Y2=0
cc_259 N_VPWR_c_390_n X 0.0112024f $X=1.055 $Y=3.33 $X2=0 $Y2=0
cc_260 N_VPWR_c_383_n X 0.00920426f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_261 N_VPWR_c_387_n N_A_633_368#_c_456_n 0.0271521f $X=3.86 $Y=2.455 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_388_n N_A_633_368#_c_456_n 0.0163338f $X=3.675 $Y=3.33 $X2=0
+ $Y2=0
cc_263 N_VPWR_c_383_n N_A_633_368#_c_456_n 0.0134516f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_264 N_VPWR_M1002_d N_A_633_368#_c_467_n 0.00505363f $X=3.705 $Y=1.84 $X2=0
+ $Y2=0
cc_265 N_VPWR_c_387_n N_A_633_368#_c_467_n 0.0221812f $X=3.86 $Y=2.455 $X2=0
+ $Y2=0
cc_266 N_VPWR_c_387_n N_A_633_368#_c_458_n 0.0266947f $X=3.86 $Y=2.455 $X2=0
+ $Y2=0
cc_267 N_VPWR_c_391_n N_A_633_368#_c_458_n 0.014549f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_268 N_VPWR_c_383_n N_A_633_368#_c_458_n 0.0119743f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_269 N_X_c_436_n N_VGND_c_485_n 0.0293294f $X=0.775 $Y=0.515 $X2=0 $Y2=0
cc_270 N_X_c_436_n N_VGND_c_486_n 0.0182488f $X=0.775 $Y=0.515 $X2=0 $Y2=0
cc_271 N_X_c_436_n N_VGND_c_491_n 0.00749631f $X=0.775 $Y=0.515 $X2=0 $Y2=0
cc_272 N_X_c_436_n N_VGND_c_494_n 0.0062048f $X=0.775 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__o2111ai_4.pex.spice
* Created: Fri Aug 28 17:52:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O2111AI_4%D1 1 3 4 6 9 11 13 14 16 18 20 21 22 23
c60 18 0 2.41904e-19 $X=1.855 $Y=1.185
c61 16 0 7.64129e-20 $X=1.81 $Y=2.4
r62 35 36 16.6033 $w=4.79e-07 $l=1.65e-07 $layer=POLY_cond $X=1.26 $Y=1.432
+ $X2=1.425 $Y2=1.432
r63 33 35 7.54697 $w=4.79e-07 $l=7.5e-08 $layer=POLY_cond $X=1.185 $Y=1.432
+ $X2=1.26 $Y2=1.432
r64 33 34 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.185
+ $Y=1.515 $X2=1.185 $Y2=1.515
r65 31 33 19.119 $w=4.79e-07 $l=1.9e-07 $layer=POLY_cond $X=0.995 $Y=1.432
+ $X2=1.185 $Y2=1.432
r66 29 31 49.3069 $w=4.79e-07 $l=4.9e-07 $layer=POLY_cond $X=0.505 $Y=1.432
+ $X2=0.995 $Y2=1.432
r67 29 30 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.505
+ $Y=1.515 $X2=0.505 $Y2=1.515
r68 27 29 1.00626 $w=4.79e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.432
+ $X2=0.505 $Y2=1.432
r69 23 34 0.402015 $w=4.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.185 $Y2=1.565
r70 22 34 12.4625 $w=4.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.185 $Y2=1.565
r71 22 30 5.76222 $w=4.28e-07 $l=2.15e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.505 $Y2=1.565
r72 21 30 7.10226 $w=4.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.505 $Y2=1.565
r73 18 38 30.3274 $w=1.5e-07 $l=2.47e-07 $layer=POLY_cond $X=1.855 $Y=1.185
+ $X2=1.855 $Y2=1.432
r74 18 20 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.855 $Y=1.185
+ $X2=1.855 $Y2=0.74
r75 14 38 4.52818 $w=4.79e-07 $l=4.5e-08 $layer=POLY_cond $X=1.81 $Y=1.432
+ $X2=1.855 $Y2=1.432
r76 14 36 38.7411 $w=4.79e-07 $l=3.85e-07 $layer=POLY_cond $X=1.81 $Y=1.432
+ $X2=1.425 $Y2=1.432
r77 14 16 289.589 $w=1.8e-07 $l=7.45e-07 $layer=POLY_cond $X=1.81 $Y=1.655
+ $X2=1.81 $Y2=2.4
r78 11 36 30.3274 $w=1.5e-07 $l=2.47e-07 $layer=POLY_cond $X=1.425 $Y=1.185
+ $X2=1.425 $Y2=1.432
r79 11 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.425 $Y=1.185
+ $X2=1.425 $Y2=0.74
r80 7 35 25.811 $w=1.8e-07 $l=2.48e-07 $layer=POLY_cond $X=1.26 $Y=1.68 $X2=1.26
+ $Y2=1.432
r81 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.26 $Y=1.68 $X2=1.26
+ $Y2=2.4
r82 4 31 30.3274 $w=1.5e-07 $l=2.47e-07 $layer=POLY_cond $X=0.995 $Y=1.185
+ $X2=0.995 $Y2=1.432
r83 4 6 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.995 $Y=1.185
+ $X2=0.995 $Y2=0.74
r84 1 27 30.3274 $w=1.5e-07 $l=2.47e-07 $layer=POLY_cond $X=0.495 $Y=1.185
+ $X2=0.495 $Y2=1.432
r85 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.495 $Y=1.185
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_4%C1 1 3 4 6 7 9 10 12 13 15 16 17 18 20 29
+ 39
c74 16 0 6.98451e-20 $X=3.5 $Y=1.26
c75 4 0 2.84156e-19 $X=2.285 $Y=1.185
r76 36 37 1.37714 $w=5.25e-07 $l=1.5e-08 $layer=POLY_cond $X=3.13 $Y=1.455
+ $X2=3.145 $Y2=1.455
r77 31 32 2.29524 $w=5.25e-07 $l=2.5e-08 $layer=POLY_cond $X=2.26 $Y=1.455
+ $X2=2.285 $Y2=1.455
r78 29 39 4.04332 $w=4.78e-07 $l=1.15e-07 $layer=LI1_cond $X=4.08 $Y=1.54
+ $X2=3.965 $Y2=1.54
r79 28 36 6.88571 $w=5.25e-07 $l=7.5e-08 $layer=POLY_cond $X=3.055 $Y=1.455
+ $X2=3.13 $Y2=1.455
r80 28 34 31.2152 $w=5.25e-07 $l=3.4e-07 $layer=POLY_cond $X=3.055 $Y=1.455
+ $X2=2.715 $Y2=1.455
r81 27 39 31.7795 $w=3.28e-07 $l=9.1e-07 $layer=LI1_cond $X=3.055 $Y=1.465
+ $X2=3.965 $Y2=1.465
r82 27 28 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.055
+ $Y=1.465 $X2=3.055 $Y2=1.465
r83 24 34 31.2152 $w=5.25e-07 $l=3.4e-07 $layer=POLY_cond $X=2.375 $Y=1.455
+ $X2=2.715 $Y2=1.455
r84 24 32 8.26286 $w=5.25e-07 $l=9e-08 $layer=POLY_cond $X=2.375 $Y=1.455
+ $X2=2.285 $Y2=1.455
r85 23 27 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.375 $Y=1.465
+ $X2=3.055 $Y2=1.465
r86 23 24 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.375
+ $Y=1.465 $X2=2.375 $Y2=1.465
r87 18 20 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.575 $Y=1.185
+ $X2=3.575 $Y2=0.74
r88 17 37 34.3153 $w=5.25e-07 $l=2.29456e-07 $layer=POLY_cond $X=3.22 $Y=1.26
+ $X2=3.145 $Y2=1.455
r89 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.5 $Y=1.26
+ $X2=3.575 $Y2=1.185
r90 16 17 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.5 $Y=1.26 $X2=3.22
+ $Y2=1.26
r91 13 37 32.6451 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.145 $Y=1.185
+ $X2=3.145 $Y2=1.455
r92 13 15 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.145 $Y=1.185
+ $X2=3.145 $Y2=0.74
r93 10 36 28.0673 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=3.13 $Y=1.725
+ $X2=3.13 $Y2=1.455
r94 10 12 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.13 $Y=1.725
+ $X2=3.13 $Y2=2.4
r95 7 34 32.6451 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.715 $Y=1.185
+ $X2=2.715 $Y2=1.455
r96 7 9 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.715 $Y=1.185
+ $X2=2.715 $Y2=0.74
r97 4 32 32.6451 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.285 $Y=1.185
+ $X2=2.285 $Y2=1.455
r98 4 6 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.285 $Y=1.185
+ $X2=2.285 $Y2=0.74
r99 1 31 28.0673 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=2.26 $Y=1.725
+ $X2=2.26 $Y2=1.455
r100 1 3 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=2.26 $Y=1.725
+ $X2=2.26 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_4%B1 1 3 4 5 6 8 13 17 21 23 25 27 28 29 30
+ 31 37
c86 37 0 1.99442e-19 $X=4.49 $Y=1.537
c87 17 0 3.32178e-19 $X=4.995 $Y=0.74
c88 1 0 2.35345e-20 $X=3.58 $Y=1.725
r89 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.675
+ $Y=1.515 $X2=5.675 $Y2=1.515
r90 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.655
+ $Y=1.515 $X2=4.655 $Y2=1.515
r91 31 45 8.71033 $w=4.28e-07 $l=3.25e-07 $layer=LI1_cond $X=6 $Y=1.565
+ $X2=5.675 $Y2=1.565
r92 30 45 4.15415 $w=4.28e-07 $l=1.55e-07 $layer=LI1_cond $X=5.52 $Y=1.565
+ $X2=5.675 $Y2=1.565
r93 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=5.52 $Y2=1.565
r94 29 40 10.3184 $w=4.28e-07 $l=3.85e-07 $layer=LI1_cond $X=5.04 $Y=1.565
+ $X2=4.655 $Y2=1.565
r95 28 40 2.54609 $w=4.28e-07 $l=9.5e-08 $layer=LI1_cond $X=4.56 $Y=1.565
+ $X2=4.655 $Y2=1.565
r96 23 44 26.6954 $w=3.75e-07 $l=1.8e-07 $layer=POLY_cond $X=5.855 $Y=1.537
+ $X2=5.675 $Y2=1.537
r97 23 25 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.855 $Y=1.35
+ $X2=5.855 $Y2=0.74
r98 19 44 37.0769 $w=3.75e-07 $l=2.5e-07 $layer=POLY_cond $X=5.425 $Y=1.537
+ $X2=5.675 $Y2=1.537
r99 19 21 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.425 $Y=1.35
+ $X2=5.425 $Y2=0.74
r100 15 19 63.7723 $w=3.75e-07 $l=4.3e-07 $layer=POLY_cond $X=4.995 $Y=1.537
+ $X2=5.425 $Y2=1.537
r101 15 39 50.4246 $w=3.75e-07 $l=3.4e-07 $layer=POLY_cond $X=4.995 $Y=1.537
+ $X2=4.655 $Y2=1.537
r102 15 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.995 $Y=1.35
+ $X2=4.995 $Y2=0.74
r103 11 39 13.3477 $w=3.75e-07 $l=9e-08 $layer=POLY_cond $X=4.565 $Y=1.537
+ $X2=4.655 $Y2=1.537
r104 11 37 31.8081 $w=3.75e-07 $l=7.5e-08 $layer=POLY_cond $X=4.565 $Y=1.537
+ $X2=4.49 $Y2=1.537
r105 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.565 $Y=1.35
+ $X2=4.565 $Y2=0.74
r106 10 27 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.22 $Y=1.65 $X2=4.13
+ $Y2=1.65
r107 10 37 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.22 $Y=1.65
+ $X2=4.49 $Y2=1.65
r108 6 27 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.13 $Y=1.725
+ $X2=4.13 $Y2=1.65
r109 6 8 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=4.13 $Y=1.725
+ $X2=4.13 $Y2=2.4
r110 4 27 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.04 $Y=1.65 $X2=4.13
+ $Y2=1.65
r111 4 5 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.04 $Y=1.65 $X2=3.67
+ $Y2=1.65
r112 1 5 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.58 $Y=1.725
+ $X2=3.67 $Y2=1.65
r113 1 3 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.58 $Y=1.725
+ $X2=3.58 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_4%A1 3 7 11 15 19 23 27 31 33 34 35 50 51
c87 15 0 1.61888e-19 $X=6.855 $Y=0.74
c88 7 0 8.45991e-20 $X=6.355 $Y=0.74
r89 51 52 12.3943 $w=3.5e-07 $l=9e-08 $layer=POLY_cond $X=7.625 $Y=1.5 $X2=7.715
+ $Y2=1.5
r90 49 51 21.3457 $w=3.5e-07 $l=1.55e-07 $layer=POLY_cond $X=7.47 $Y=1.5
+ $X2=7.625 $Y2=1.5
r91 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.47
+ $Y=1.515 $X2=7.47 $Y2=1.515
r92 47 49 25.4771 $w=3.5e-07 $l=1.85e-07 $layer=POLY_cond $X=7.285 $Y=1.5
+ $X2=7.47 $Y2=1.5
r93 46 47 15.1486 $w=3.5e-07 $l=1.1e-07 $layer=POLY_cond $X=7.175 $Y=1.5
+ $X2=7.285 $Y2=1.5
r94 45 46 44.0686 $w=3.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.855 $Y=1.5
+ $X2=7.175 $Y2=1.5
r95 44 45 17.9029 $w=3.5e-07 $l=1.3e-07 $layer=POLY_cond $X=6.725 $Y=1.5
+ $X2=6.855 $Y2=1.5
r96 42 44 37.8714 $w=3.5e-07 $l=2.75e-07 $layer=POLY_cond $X=6.45 $Y=1.5
+ $X2=6.725 $Y2=1.5
r97 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.45
+ $Y=1.515 $X2=6.45 $Y2=1.515
r98 40 42 13.0829 $w=3.5e-07 $l=9.5e-08 $layer=POLY_cond $X=6.355 $Y=1.5
+ $X2=6.45 $Y2=1.5
r99 39 40 13.0829 $w=3.5e-07 $l=9.5e-08 $layer=POLY_cond $X=6.26 $Y=1.5
+ $X2=6.355 $Y2=1.5
r100 35 50 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.47 $Y2=1.565
r101 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.44 $Y2=1.565
r102 33 34 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.96 $Y2=1.565
r103 33 43 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.45 $Y2=1.565
r104 29 52 22.6286 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.715 $Y=1.32
+ $X2=7.715 $Y2=1.5
r105 29 31 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.715 $Y=1.32
+ $X2=7.715 $Y2=0.74
r106 25 51 18.307 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=7.625 $Y=1.68
+ $X2=7.625 $Y2=1.5
r107 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.625 $Y=1.68
+ $X2=7.625 $Y2=2.4
r108 21 47 22.6286 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.285 $Y=1.32
+ $X2=7.285 $Y2=1.5
r109 21 23 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.285 $Y=1.32
+ $X2=7.285 $Y2=0.74
r110 17 46 18.307 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=7.175 $Y=1.68
+ $X2=7.175 $Y2=1.5
r111 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.175 $Y=1.68
+ $X2=7.175 $Y2=2.4
r112 13 45 22.6286 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.855 $Y=1.32
+ $X2=6.855 $Y2=1.5
r113 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.855 $Y=1.32
+ $X2=6.855 $Y2=0.74
r114 9 44 18.307 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=6.725 $Y=1.68
+ $X2=6.725 $Y2=1.5
r115 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.725 $Y=1.68
+ $X2=6.725 $Y2=2.4
r116 5 40 22.6286 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.355 $Y=1.32
+ $X2=6.355 $Y2=1.5
r117 5 7 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.355 $Y=1.32
+ $X2=6.355 $Y2=0.74
r118 1 39 18.307 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=6.26 $Y=1.68 $X2=6.26
+ $Y2=1.5
r119 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.26 $Y=1.68 $X2=6.26
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_4%A2 3 5 7 10 12 14 15 17 18 20 21 23 24 26
+ 27 28 29 30 46 47
c86 10 0 6.66039e-20 $X=8.575 $Y=2.4
r87 47 48 0.985685 $w=4.89e-07 $l=1e-08 $layer=POLY_cond $X=9.575 $Y=1.495
+ $X2=9.585 $Y2=1.495
r88 45 47 16.7566 $w=4.89e-07 $l=1.7e-07 $layer=POLY_cond $X=9.405 $Y=1.495
+ $X2=9.575 $Y2=1.495
r89 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.405
+ $Y=1.515 $X2=9.405 $Y2=1.515
r90 43 45 24.6421 $w=4.89e-07 $l=2.5e-07 $layer=POLY_cond $X=9.155 $Y=1.495
+ $X2=9.405 $Y2=1.495
r91 42 43 7.88548 $w=4.89e-07 $l=8e-08 $layer=POLY_cond $X=9.075 $Y=1.495
+ $X2=9.155 $Y2=1.495
r92 41 42 42.3845 $w=4.89e-07 $l=4.3e-07 $layer=POLY_cond $X=8.645 $Y=1.495
+ $X2=9.075 $Y2=1.495
r93 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.385
+ $Y=1.515 $X2=8.385 $Y2=1.515
r94 36 38 23.6564 $w=4.89e-07 $l=2.4e-07 $layer=POLY_cond $X=8.145 $Y=1.495
+ $X2=8.385 $Y2=1.495
r95 30 46 1.20605 $w=4.28e-07 $l=4.5e-08 $layer=LI1_cond $X=9.36 $Y=1.565
+ $X2=9.405 $Y2=1.565
r96 29 30 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.565
+ $X2=9.36 $Y2=1.565
r97 28 29 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.4 $Y=1.565
+ $X2=8.88 $Y2=1.565
r98 28 39 0.402015 $w=4.28e-07 $l=1.5e-08 $layer=LI1_cond $X=8.4 $Y=1.565
+ $X2=8.385 $Y2=1.565
r99 27 39 12.4625 $w=4.28e-07 $l=4.65e-07 $layer=LI1_cond $X=7.92 $Y=1.565
+ $X2=8.385 $Y2=1.565
r100 24 48 30.8469 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.585 $Y=1.225
+ $X2=9.585 $Y2=1.495
r101 24 26 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=9.585 $Y=1.225
+ $X2=9.585 $Y2=0.74
r102 21 47 26.3167 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=9.575 $Y=1.765
+ $X2=9.575 $Y2=1.495
r103 21 23 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=9.575 $Y=1.765
+ $X2=9.575 $Y2=2.4
r104 18 43 30.8469 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.155 $Y=1.225
+ $X2=9.155 $Y2=1.495
r105 18 20 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=9.155 $Y=1.225
+ $X2=9.155 $Y2=0.74
r106 15 42 26.3167 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=9.075 $Y=1.765
+ $X2=9.075 $Y2=1.495
r107 15 17 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=9.075 $Y=1.765
+ $X2=9.075 $Y2=2.4
r108 12 41 30.8469 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=8.645 $Y=1.225
+ $X2=8.645 $Y2=1.495
r109 12 14 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=8.645 $Y=1.225
+ $X2=8.645 $Y2=0.74
r110 8 41 6.8998 $w=4.89e-07 $l=7e-08 $layer=POLY_cond $X=8.575 $Y=1.495
+ $X2=8.645 $Y2=1.495
r111 8 38 18.728 $w=4.89e-07 $l=1.9e-07 $layer=POLY_cond $X=8.575 $Y=1.495
+ $X2=8.385 $Y2=1.495
r112 8 10 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.575 $Y=1.68
+ $X2=8.575 $Y2=2.4
r113 5 36 30.8469 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=8.145 $Y=1.225
+ $X2=8.145 $Y2=1.495
r114 5 7 155.847 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=8.145 $Y=1.225
+ $X2=8.145 $Y2=0.74
r115 1 36 5.42127 $w=4.89e-07 $l=5.5e-08 $layer=POLY_cond $X=8.09 $Y=1.495
+ $X2=8.145 $Y2=1.495
r116 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.09 $Y=1.68 $X2=8.09
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_4%Y 1 2 3 4 5 6 7 8 25 29 31 32 35 37 38 41
+ 43 47 49 53 65 68 74 76 78 79
c131 43 0 6.98451e-20 $X=4.19 $Y=2.035
c132 37 0 2.35345e-20 $X=3.19 $Y=1.885
c133 31 0 9.95308e-20 $X=1.685 $Y=1.13
r134 71 72 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=3.355 $Y=1.985
+ $X2=3.355 $Y2=2.035
r135 68 71 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=3.355 $Y=1.885
+ $X2=3.355 $Y2=1.985
r136 64 65 13.0168 $w=1.028e-06 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=2.465
+ $X2=1.2 $Y2=2.465
r137 61 64 4.50097 $w=1.028e-06 $l=3.8e-07 $layer=LI1_cond $X=0.655 $Y=2.465
+ $X2=1.035 $Y2=2.465
r138 58 61 4.44175 $w=1.028e-06 $l=3.75e-07 $layer=LI1_cond $X=0.28 $Y=2.465
+ $X2=0.655 $Y2=2.465
r139 54 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.515 $Y=2.035
+ $X2=8.35 $Y2=2.035
r140 53 78 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.185 $Y=2.035
+ $X2=9.35 $Y2=2.035
r141 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.185 $Y=2.035
+ $X2=8.515 $Y2=2.035
r142 50 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.52 $Y=2.035
+ $X2=4.355 $Y2=2.035
r143 49 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.185 $Y=2.035
+ $X2=8.35 $Y2=2.035
r144 49 50 239.107 $w=1.68e-07 $l=3.665e-06 $layer=LI1_cond $X=8.185 $Y=2.035
+ $X2=4.52 $Y2=2.035
r145 45 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.355 $Y=2.12
+ $X2=4.355 $Y2=2.035
r146 45 47 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.355 $Y=2.12
+ $X2=4.355 $Y2=2.815
r147 44 72 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.52 $Y=2.035
+ $X2=3.355 $Y2=2.035
r148 43 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.19 $Y=2.035
+ $X2=4.355 $Y2=2.035
r149 43 44 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.19 $Y=2.035
+ $X2=3.52 $Y2=2.035
r150 39 72 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=2.12
+ $X2=3.355 $Y2=2.035
r151 39 41 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.355 $Y=2.12
+ $X2=3.355 $Y2=2.815
r152 38 85 8.97309 $w=3.43e-07 $l=1.88348e-07 $layer=LI1_cond $X=2.2 $Y=1.885
+ $X2=2.035 $Y2=1.835
r153 37 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.19 $Y=1.885
+ $X2=3.355 $Y2=1.885
r154 37 38 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=3.19 $Y=1.885
+ $X2=2.2 $Y2=1.885
r155 33 85 0.950996 $w=3.3e-07 $l=2.85e-07 $layer=LI1_cond $X=2.035 $Y=2.12
+ $X2=2.035 $Y2=1.835
r156 33 35 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.035 $Y=2.12
+ $X2=2.035 $Y2=2.815
r157 32 85 12.449 $w=3.43e-07 $l=4.71434e-07 $layer=LI1_cond $X=1.685 $Y=1.55
+ $X2=2.035 $Y2=1.835
r158 32 79 0.177843 $w=3.43e-07 $l=1.17473e-07 $layer=LI1_cond $X=1.685 $Y=1.55
+ $X2=1.68 $Y2=1.665
r159 31 67 4.30634 $w=2.4e-07 $l=1.8e-07 $layer=LI1_cond $X=1.685 $Y=1.13
+ $X2=1.685 $Y2=0.95
r160 31 32 20.1678 $w=2.38e-07 $l=4.2e-07 $layer=LI1_cond $X=1.685 $Y=1.13
+ $X2=1.685 $Y2=1.55
r161 29 79 9.8623 $w=3.43e-07 $l=4.55192e-07 $layer=LI1_cond $X=1.87 $Y=2.035
+ $X2=1.68 $Y2=1.665
r162 29 65 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.87 $Y=2.035
+ $X2=1.2 $Y2=2.035
r163 25 67 2.87089 $w=3.6e-07 $l=1.2e-07 $layer=LI1_cond $X=1.565 $Y=0.95
+ $X2=1.685 $Y2=0.95
r164 25 27 25.1297 $w=3.58e-07 $l=7.85e-07 $layer=LI1_cond $X=1.565 $Y=0.95
+ $X2=0.78 $Y2=0.95
r165 8 78 300 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=2 $X=9.165
+ $Y=1.84 $X2=9.35 $Y2=2.115
r166 7 76 300 $w=1.7e-07 $l=3.49821e-07 $layer=licon1_PDIFF $count=2 $X=8.18
+ $Y=1.84 $X2=8.35 $Y2=2.115
r167 6 74 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=4.22
+ $Y=1.84 $X2=4.355 $Y2=2.115
r168 6 47 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.22
+ $Y=1.84 $X2=4.355 $Y2=2.815
r169 5 71 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.22
+ $Y=1.84 $X2=3.355 $Y2=1.985
r170 5 41 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.22
+ $Y=1.84 $X2=3.355 $Y2=2.815
r171 4 85 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.9
+ $Y=1.84 $X2=2.035 $Y2=1.985
r172 4 35 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.9
+ $Y=1.84 $X2=2.035 $Y2=2.815
r173 3 64 266.667 $w=1.7e-07 $l=1.1463e-06 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=1.035 $Y2=2.4
r174 3 61 266.667 $w=1.7e-07 $l=1.20732e-06 $layer=licon1_PDIFF $count=2
+ $X=0.135 $Y=1.84 $X2=0.655 $Y2=2.815
r175 3 61 266.667 $w=1.7e-07 $l=6.09754e-07 $layer=licon1_PDIFF $count=2
+ $X=0.135 $Y=1.84 $X2=0.655 $Y2=2.035
r176 3 58 266.667 $w=1.7e-07 $l=6.28331e-07 $layer=licon1_PDIFF $count=2
+ $X=0.135 $Y=1.84 $X2=0.28 $Y2=2.4
r177 2 67 182 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.64 $Y2=0.91
r178 1 27 182 $w=1.7e-07 $l=6.76905e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_4%VPWR 1 2 3 4 5 18 22 26 30 34 37 38 40 41
+ 42 51 59 66 73 74 77 80 83
r98 83 84 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r99 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r100 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r101 74 84 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=7.44 $Y2=3.33
r102 73 74 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r103 71 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.485 $Y=3.33
+ $X2=7.4 $Y2=3.33
r104 71 73 153.642 $w=1.68e-07 $l=2.355e-06 $layer=LI1_cond $X=7.485 $Y=3.33
+ $X2=9.84 $Y2=3.33
r105 70 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r106 70 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r107 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r108 67 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.585 $Y=3.33
+ $X2=6.46 $Y2=3.33
r109 67 69 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.585 $Y=3.33
+ $X2=6.96 $Y2=3.33
r110 66 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.315 $Y=3.33
+ $X2=7.4 $Y2=3.33
r111 66 69 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.315 $Y=3.33
+ $X2=6.96 $Y2=3.33
r112 65 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r113 64 65 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r114 61 64 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=3.33 $X2=6
+ $Y2=3.33
r115 61 62 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r116 59 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.335 $Y=3.33
+ $X2=6.46 $Y2=3.33
r117 59 64 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.335 $Y=3.33
+ $X2=6 $Y2=3.33
r118 58 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r119 58 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r120 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r121 55 77 13.1282 $w=1.7e-07 $l=3.25e-07 $layer=LI1_cond $X=3.02 $Y=3.33
+ $X2=2.695 $Y2=3.33
r122 55 57 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.02 $Y=3.33
+ $X2=3.6 $Y2=3.33
r123 54 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r124 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r125 51 77 13.1282 $w=1.7e-07 $l=3.25e-07 $layer=LI1_cond $X=2.37 $Y=3.33
+ $X2=2.695 $Y2=3.33
r126 51 53 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.37 $Y=3.33
+ $X2=2.16 $Y2=3.33
r127 50 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r128 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r129 46 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r130 45 49 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r131 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r132 42 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r133 42 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.08 $Y2=3.33
r134 40 57 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.69 $Y=3.33 $X2=3.6
+ $Y2=3.33
r135 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.69 $Y=3.33
+ $X2=3.855 $Y2=3.33
r136 39 61 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=4.02 $Y=3.33 $X2=4.08
+ $Y2=3.33
r137 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.02 $Y=3.33
+ $X2=3.855 $Y2=3.33
r138 37 49 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.37 $Y=3.33
+ $X2=1.2 $Y2=3.33
r139 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.37 $Y=3.33
+ $X2=1.535 $Y2=3.33
r140 36 53 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=1.7 $Y=3.33
+ $X2=2.16 $Y2=3.33
r141 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.7 $Y=3.33
+ $X2=1.535 $Y2=3.33
r142 32 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.4 $Y=3.245 $X2=7.4
+ $Y2=3.33
r143 32 34 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=7.4 $Y=3.245
+ $X2=7.4 $Y2=2.805
r144 28 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.46 $Y=3.245
+ $X2=6.46 $Y2=3.33
r145 28 30 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=6.46 $Y=3.245
+ $X2=6.46 $Y2=2.805
r146 24 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.855 $Y=3.245
+ $X2=3.855 $Y2=3.33
r147 24 26 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=3.855 $Y=3.245
+ $X2=3.855 $Y2=2.455
r148 20 77 2.7021 $w=6.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=3.245
+ $X2=2.695 $Y2=3.33
r149 20 22 17.2971 $w=6.48e-07 $l=9.4e-07 $layer=LI1_cond $X=2.695 $Y=3.245
+ $X2=2.695 $Y2=2.305
r150 16 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=3.245
+ $X2=1.535 $Y2=3.33
r151 16 18 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.535 $Y=3.245
+ $X2=1.535 $Y2=2.455
r152 5 34 600 $w=1.7e-07 $l=1.03029e-06 $layer=licon1_PDIFF $count=1 $X=7.265
+ $Y=1.84 $X2=7.4 $Y2=2.805
r153 4 30 600 $w=1.7e-07 $l=1.03729e-06 $layer=licon1_PDIFF $count=1 $X=6.35
+ $Y=1.84 $X2=6.5 $Y2=2.805
r154 3 26 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=3.67
+ $Y=1.84 $X2=3.855 $Y2=2.455
r155 2 22 150 $w=1.7e-07 $l=7.52396e-07 $layer=licon1_PDIFF $count=4 $X=2.35
+ $Y=1.84 $X2=2.905 $Y2=2.305
r156 1 18 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=1.35
+ $Y=1.84 $X2=1.535 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_4%A_954_368# 1 2 3 4 5 16 22 26 28 29 30 31
+ 34 36 40 46 48 51
c69 28 0 6.66039e-20 $X=7.85 $Y=2.46
r70 45 46 10.2208 $w=6.88e-07 $l=1.35e-07 $layer=LI1_cond $X=6.03 $Y=2.635
+ $X2=6.165 $Y2=2.635
r71 40 43 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=9.84 $Y=1.985
+ $X2=9.84 $Y2=2.815
r72 38 43 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=9.84 $Y=2.905 $X2=9.84
+ $Y2=2.815
r73 37 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.015 $Y=2.99
+ $X2=8.85 $Y2=2.99
r74 36 38 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.715 $Y=2.99
+ $X2=9.84 $Y2=2.905
r75 36 37 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=9.715 $Y=2.99
+ $X2=9.015 $Y2=2.99
r76 32 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.85 $Y=2.905
+ $X2=8.85 $Y2=2.99
r77 32 34 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=8.85 $Y=2.905
+ $X2=8.85 $Y2=2.455
r78 30 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.685 $Y=2.99
+ $X2=8.85 $Y2=2.99
r79 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.685 $Y=2.99
+ $X2=8.015 $Y2=2.99
r80 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.85 $Y=2.905
+ $X2=8.015 $Y2=2.99
r81 28 50 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.85 $Y=2.46 $X2=7.85
+ $Y2=2.375
r82 28 29 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=7.85 $Y=2.46
+ $X2=7.85 $Y2=2.905
r83 27 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.115 $Y=2.375
+ $X2=6.95 $Y2=2.375
r84 26 50 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.685 $Y=2.375
+ $X2=7.85 $Y2=2.375
r85 26 27 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=7.685 $Y=2.375
+ $X2=7.115 $Y2=2.375
r86 22 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.785 $Y=2.375
+ $X2=6.95 $Y2=2.375
r87 22 46 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=6.785 $Y=2.375
+ $X2=6.165 $Y2=2.375
r88 18 21 12.5675 $w=6.88e-07 $l=7.25e-07 $layer=LI1_cond $X=4.945 $Y=2.635
+ $X2=5.67 $Y2=2.635
r89 16 45 3.64024 $w=6.88e-07 $l=2.1e-07 $layer=LI1_cond $X=5.82 $Y=2.635
+ $X2=6.03 $Y2=2.635
r90 16 21 2.60017 $w=6.88e-07 $l=1.5e-07 $layer=LI1_cond $X=5.82 $Y=2.635
+ $X2=5.67 $Y2=2.635
r91 5 43 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.665
+ $Y=1.84 $X2=9.8 $Y2=2.815
r92 5 40 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.665
+ $Y=1.84 $X2=9.8 $Y2=1.985
r93 4 34 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=8.665
+ $Y=1.84 $X2=8.85 $Y2=2.455
r94 3 50 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=7.715
+ $Y=1.84 $X2=7.85 $Y2=2.455
r95 2 48 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=6.815
+ $Y=1.84 $X2=6.95 $Y2=2.455
r96 1 45 300 $w=1.7e-07 $l=1.50389e-06 $layer=licon1_PDIFF $count=2 $X=4.77
+ $Y=1.84 $X2=6.03 $Y2=2.375
r97 1 21 200 $w=1.7e-07 $l=1.13644e-06 $layer=licon1_PDIFF $count=3 $X=4.77
+ $Y=1.84 $X2=5.67 $Y2=2.375
r98 1 18 200 $w=1.7e-07 $l=6.1632e-07 $layer=licon1_PDIFF $count=3 $X=4.77
+ $Y=1.84 $X2=4.945 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_4%A_27_74# 1 2 3 4 5 18 22 23 28 31
c47 23 0 1.61246e-19 $X=2.07 $Y=0.815
c48 22 0 1.84625e-19 $X=2.07 $Y=0.6
r49 26 28 31.4635 $w=3.13e-07 $l=8.6e-07 $layer=LI1_cond $X=2.93 $Y=0.972
+ $X2=3.79 $Y2=0.972
r50 24 35 2.68365 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=0.972
+ $X2=2.07 $Y2=0.972
r51 24 26 28.3538 $w=3.13e-07 $l=7.75e-07 $layer=LI1_cond $X=2.155 $Y=0.972
+ $X2=2.93 $Y2=0.972
r52 23 35 4.95685 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=2.07 $Y=0.815
+ $X2=2.07 $Y2=0.972
r53 22 33 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.07 $Y=0.6 $X2=2.07
+ $Y2=0.475
r54 22 23 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.07 $Y=0.6
+ $X2=2.07 $Y2=0.815
r55 19 31 3.97509 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=0.475
+ $X2=0.28 $Y2=0.475
r56 19 21 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=0.445 $Y=0.475
+ $X2=1.21 $Y2=0.475
r57 18 33 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=0.475
+ $X2=2.07 $Y2=0.475
r58 18 21 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=1.985 $Y=0.475
+ $X2=1.21 $Y2=0.475
r59 5 28 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=3.65
+ $Y=0.37 $X2=3.79 $Y2=0.95
r60 4 26 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=2.79
+ $Y=0.37 $X2=2.93 $Y2=0.95
r61 3 35 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.37 $X2=2.07 $Y2=0.965
r62 3 33 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.37 $X2=2.07 $Y2=0.515
r63 2 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.21 $Y2=0.515
r64 1 31 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_4%A_472_74# 1 2 3 4 22 23
c28 23 0 8.0658e-20 $X=5.475 $Y=0.515
c29 22 0 2.50688e-19 $X=5.64 $Y=0.515
r30 22 23 5.91831 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.64 $Y=0.515
+ $X2=5.475 $Y2=0.515
r31 20 23 27.1508 $w=2.93e-07 $l=6.95e-07 $layer=LI1_cond $X=4.78 $Y=0.497
+ $X2=5.475 $Y2=0.497
r32 18 20 55.4735 $w=2.93e-07 $l=1.42e-06 $layer=LI1_cond $X=3.36 $Y=0.497
+ $X2=4.78 $Y2=0.497
r33 15 18 33.5966 $w=2.93e-07 $l=8.6e-07 $layer=LI1_cond $X=2.5 $Y=0.497
+ $X2=3.36 $Y2=0.497
r34 4 22 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.5
+ $Y=0.37 $X2=5.64 $Y2=0.515
r35 3 20 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.64
+ $Y=0.37 $X2=4.78 $Y2=0.515
r36 2 18 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.22
+ $Y=0.37 $X2=3.36 $Y2=0.515
r37 1 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.36
+ $Y=0.37 $X2=2.5 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_4%A_841_74# 1 2 3 4 5 6 7 24 27 30 32 36 38
+ 42 44 48 50 54 59 60 62 63 64 65
c108 59 0 3.65531e-19 $X=4.515 $Y=0.972
c109 30 0 1.61888e-19 $X=6.14 $Y=0.515
r110 59 60 21.8141 $w=2.78e-07 $l=5.3e-07 $layer=LI1_cond $X=4.515 $Y=0.99
+ $X2=5.045 $Y2=0.99
r111 57 59 6.20639 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=4.35 $Y=0.972
+ $X2=4.515 $Y2=0.972
r112 52 54 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=9.84 $Y=1.01
+ $X2=9.84 $Y2=0.515
r113 51 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.025 $Y=1.095
+ $X2=8.9 $Y2=1.095
r114 50 52 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.715 $Y=1.095
+ $X2=9.84 $Y2=1.01
r115 50 51 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.715 $Y=1.095
+ $X2=9.025 $Y2=1.095
r116 46 65 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.9 $Y=1.01
+ $X2=8.9 $Y2=1.095
r117 46 48 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=8.9 $Y=1.01
+ $X2=8.9 $Y2=0.515
r118 45 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.095 $Y=1.095
+ $X2=7.97 $Y2=1.095
r119 44 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.775 $Y=1.095
+ $X2=8.9 $Y2=1.095
r120 44 45 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.775 $Y=1.095
+ $X2=8.095 $Y2=1.095
r121 40 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.97 $Y=1.01
+ $X2=7.97 $Y2=1.095
r122 40 42 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=7.97 $Y=1.01
+ $X2=7.97 $Y2=0.515
r123 39 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.155 $Y=1.095
+ $X2=7.07 $Y2=1.095
r124 38 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.845 $Y=1.095
+ $X2=7.97 $Y2=1.095
r125 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.845 $Y=1.095
+ $X2=7.155 $Y2=1.095
r126 34 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.07 $Y=1.01
+ $X2=7.07 $Y2=1.095
r127 34 36 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=7.07 $Y=1.01
+ $X2=7.07 $Y2=0.515
r128 33 62 6.46576 $w=2.5e-07 $l=2.0106e-07 $layer=LI1_cond $X=6.305 $Y=1.095
+ $X2=6.14 $Y2=1.015
r129 32 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.985 $Y=1.095
+ $X2=7.07 $Y2=1.095
r130 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.985 $Y=1.095
+ $X2=6.305 $Y2=1.095
r131 28 62 0.364692 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=6.14 $Y=0.85
+ $X2=6.14 $Y2=1.015
r132 28 30 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.14 $Y=0.85
+ $X2=6.14 $Y2=0.515
r133 27 60 6.05995 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.21 $Y=1.015
+ $X2=5.045 $Y2=1.015
r134 24 62 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=5.975 $Y=1.015
+ $X2=6.14 $Y2=1.015
r135 24 27 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=5.975 $Y=1.015
+ $X2=5.21 $Y2=1.015
r136 7 54 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.66
+ $Y=0.37 $X2=9.8 $Y2=0.515
r137 6 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.72
+ $Y=0.37 $X2=8.86 $Y2=0.515
r138 5 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.79
+ $Y=0.37 $X2=7.93 $Y2=0.515
r139 4 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.93
+ $Y=0.37 $X2=7.07 $Y2=0.515
r140 3 62 182 $w=1.7e-07 $l=6.9208e-07 $layer=licon1_NDIFF $count=1 $X=5.93
+ $Y=0.37 $X2=6.14 $Y2=0.965
r141 3 30 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.93
+ $Y=0.37 $X2=6.14 $Y2=0.515
r142 2 27 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=5.07
+ $Y=0.37 $X2=5.21 $Y2=0.95
r143 1 57 182 $w=1.7e-07 $l=6.4846e-07 $layer=licon1_NDIFF $count=1 $X=4.205
+ $Y=0.37 $X2=4.35 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_MS__O2111AI_4%VGND 1 2 3 4 15 19 23 27 29 31 36 41 46 53
+ 54 57 60 63 66
r103 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r104 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r105 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r106 57 58 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r107 54 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r108 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r109 51 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.535 $Y=0 $X2=9.37
+ $Y2=0
r110 51 53 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.535 $Y=0
+ $X2=9.84 $Y2=0
r111 50 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r112 50 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r113 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r114 47 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.595 $Y=0 $X2=8.43
+ $Y2=0
r115 47 49 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.595 $Y=0
+ $X2=8.88 $Y2=0
r116 46 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.205 $Y=0 $X2=9.37
+ $Y2=0
r117 46 49 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.205 $Y=0
+ $X2=8.88 $Y2=0
r118 45 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r119 45 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r120 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r121 42 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.665 $Y=0 $X2=7.5
+ $Y2=0
r122 42 44 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.665 $Y=0
+ $X2=7.92 $Y2=0
r123 41 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.265 $Y=0 $X2=8.43
+ $Y2=0
r124 41 44 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.265 $Y=0 $X2=7.92
+ $Y2=0
r125 40 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r126 40 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r127 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r128 37 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.805 $Y=0 $X2=6.64
+ $Y2=0
r129 37 39 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=6.805 $Y=0
+ $X2=6.96 $Y2=0
r130 36 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.335 $Y=0 $X2=7.5
+ $Y2=0
r131 36 39 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.335 $Y=0
+ $X2=6.96 $Y2=0
r132 33 34 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r133 31 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.475 $Y=0 $X2=6.64
+ $Y2=0
r134 31 33 406.775 $w=1.68e-07 $l=6.235e-06 $layer=LI1_cond $X=6.475 $Y=0
+ $X2=0.24 $Y2=0
r135 29 58 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.48 $Y2=0
r136 29 34 1.33793 $w=4.9e-07 $l=4.8e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=0.24
+ $Y2=0
r137 25 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.37 $Y=0.085
+ $X2=9.37 $Y2=0
r138 25 27 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=9.37 $Y=0.085
+ $X2=9.37 $Y2=0.655
r139 21 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.43 $Y=0.085
+ $X2=8.43 $Y2=0
r140 21 23 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=8.43 $Y=0.085
+ $X2=8.43 $Y2=0.655
r141 17 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.5 $Y=0.085 $X2=7.5
+ $Y2=0
r142 17 19 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=7.5 $Y=0.085
+ $X2=7.5 $Y2=0.655
r143 13 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.64 $Y=0.085
+ $X2=6.64 $Y2=0
r144 13 15 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=6.64 $Y=0.085
+ $X2=6.64 $Y2=0.655
r145 4 27 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=9.23
+ $Y=0.37 $X2=9.37 $Y2=0.655
r146 3 23 182 $w=1.7e-07 $l=3.756e-07 $layer=licon1_NDIFF $count=1 $X=8.22
+ $Y=0.37 $X2=8.43 $Y2=0.655
r147 2 19 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=7.36
+ $Y=0.37 $X2=7.5 $Y2=0.655
r148 1 15 182 $w=1.7e-07 $l=3.756e-07 $layer=licon1_NDIFF $count=1 $X=6.43
+ $Y=0.37 $X2=6.64 $Y2=0.655
.ends


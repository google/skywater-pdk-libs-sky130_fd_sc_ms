* File: sky130_fd_sc_ms__maj3_2.spice
* Created: Fri Aug 28 17:38:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__maj3_2.pex.spice"
.subckt sky130_fd_sc_ms__maj3_2  VNB VPB B C A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* C	C
* B	B
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A_87_264#_M1011_g N_X_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75004 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1014_d N_A_87_264#_M1014_g N_X_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.33115 AS=0.1036 PD=1.635 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1008 A_413_74# N_A_M1008_g N_VGND_M1014_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.33115 PD=0.98 PS=1.635 NRD=10.536 NRS=10.536 M=1 R=4.93333 SA=75001.7
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1009 N_A_87_264#_M1009_d N_B_M1009_g A_413_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.0888 PD=1.02 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75002.1
+ SB=75002.1 A=0.111 P=1.78 MULT=1
MM1002 A_577_74# N_B_M1002_g N_A_87_264#_M1009_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1221 AS=0.1036 PD=1.07 PS=1.02 NRD=17.832 NRS=0 M=1 R=4.93333 SA=75002.5
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_C_M1003_g A_577_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1665
+ AS=0.1221 PD=1.19 PS=1.07 NRD=13.776 NRS=17.832 M=1 R=4.93333 SA=75003
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1012 A_793_74# N_A_M1012_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.1665 PD=0.98 PS=1.19 NRD=10.536 NRS=13.776 M=1 R=4.93333 SA=75003.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1013 N_A_87_264#_M1013_d N_C_M1013_g A_793_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.0888 PD=2.05 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75004
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_VPWR_M1004_d N_A_87_264#_M1004_g N_X_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003.4 A=0.2016 P=2.6 MULT=1
MM1005 N_VPWR_M1005_d N_A_87_264#_M1005_g N_X_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.409223 AS=0.1512 PD=1.96 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90002.9 A=0.2016 P=2.6 MULT=1
MM1000 A_396_368# N_A_M1000_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=1 AD=0.171687
+ AS=0.365377 PD=1.43 PS=1.75 NRD=22.9702 NRS=0 M=1 R=5.55556 SA=90001.6
+ SB=90002.3 A=0.18 P=2.36 MULT=1
MM1007 N_A_87_264#_M1007_d N_B_M1007_g A_396_368# VPB PSHORT L=0.18 W=1 AD=0.135
+ AS=0.171687 PD=1.27 PS=1.43 NRD=0 NRS=22.9702 M=1 R=5.55556 SA=90001.9
+ SB=90002 A=0.18 P=2.36 MULT=1
MM1010 A_587_347# N_B_M1010_g N_A_87_264#_M1007_d VPB PSHORT L=0.18 W=1 AD=0.14
+ AS=0.135 PD=1.28 PS=1.27 NRD=16.7253 NRS=0 M=1 R=5.55556 SA=90002.3 SB=90001.5
+ A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_C_M1001_g A_587_347# VPB PSHORT L=0.18 W=1 AD=0.2034
+ AS=0.14 PD=1.495 PS=1.28 NRD=23.1278 NRS=16.7253 M=1 R=5.55556 SA=90002.8
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1006 A_793_368# N_A_M1006_g N_VPWR_M1001_d VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.2034 PD=1.24 PS=1.495 NRD=12.7853 NRS=0 M=1 R=5.55556 SA=90003.2
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1015 N_A_87_264#_M1015_d N_C_M1015_g A_793_368# VPB PSHORT L=0.18 W=1 AD=0.28
+ AS=0.12 PD=2.56 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556 SA=90003.6 SB=90000.2
+ A=0.18 P=2.36 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.83955 P=14.29
*
.include "sky130_fd_sc_ms__maj3_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__dlrtn_4.pxi.spice
* Created: Wed Sep  2 12:05:36 2020
* 
x_PM_SKY130_FD_SC_MS__DLRTN_4%D N_D_M1024_g N_D_M1013_g D N_D_c_174_n
+ PM_SKY130_FD_SC_MS__DLRTN_4%D
x_PM_SKY130_FD_SC_MS__DLRTN_4%GATE_N N_GATE_N_M1007_g N_GATE_N_M1003_g GATE_N
+ N_GATE_N_c_206_n PM_SKY130_FD_SC_MS__DLRTN_4%GATE_N
x_PM_SKY130_FD_SC_MS__DLRTN_4%A_232_98# N_A_232_98#_M1003_d N_A_232_98#_M1007_d
+ N_A_232_98#_M1008_g N_A_232_98#_M1020_g N_A_232_98#_M1017_g
+ N_A_232_98#_M1000_g N_A_232_98#_c_244_n N_A_232_98#_c_245_n
+ N_A_232_98#_c_254_n N_A_232_98#_c_246_n N_A_232_98#_c_255_n
+ N_A_232_98#_c_256_n N_A_232_98#_c_257_n N_A_232_98#_c_258_n
+ N_A_232_98#_c_259_n N_A_232_98#_c_260_n N_A_232_98#_c_261_n
+ N_A_232_98#_c_247_n N_A_232_98#_c_248_n PM_SKY130_FD_SC_MS__DLRTN_4%A_232_98#
x_PM_SKY130_FD_SC_MS__DLRTN_4%A_27_136# N_A_27_136#_M1024_s N_A_27_136#_M1013_s
+ N_A_27_136#_c_361_n N_A_27_136#_M1005_g N_A_27_136#_c_362_n
+ N_A_27_136#_c_363_n N_A_27_136#_M1018_g N_A_27_136#_c_364_n
+ N_A_27_136#_c_365_n N_A_27_136#_c_366_n N_A_27_136#_c_367_n
+ N_A_27_136#_c_368_n N_A_27_136#_c_373_n N_A_27_136#_c_369_n
+ PM_SKY130_FD_SC_MS__DLRTN_4%A_27_136#
x_PM_SKY130_FD_SC_MS__DLRTN_4%A_348_392# N_A_348_392#_M1020_s
+ N_A_348_392#_M1008_s N_A_348_392#_M1028_g N_A_348_392#_M1006_g
+ N_A_348_392#_c_443_n N_A_348_392#_c_451_n N_A_348_392#_c_452_n
+ N_A_348_392#_c_444_n N_A_348_392#_c_445_n N_A_348_392#_c_446_n
+ N_A_348_392#_c_447_n N_A_348_392#_c_448_n N_A_348_392#_c_454_n
+ PM_SKY130_FD_SC_MS__DLRTN_4%A_348_392#
x_PM_SKY130_FD_SC_MS__DLRTN_4%A_888_406# N_A_888_406#_M1009_s
+ N_A_888_406#_M1012_d N_A_888_406#_M1014_d N_A_888_406#_M1010_g
+ N_A_888_406#_M1015_g N_A_888_406#_c_556_n N_A_888_406#_M1019_g
+ N_A_888_406#_c_538_n N_A_888_406#_c_539_n N_A_888_406#_M1001_g
+ N_A_888_406#_M1023_g N_A_888_406#_M1004_g N_A_888_406#_M1025_g
+ N_A_888_406#_M1011_g N_A_888_406#_M1027_g N_A_888_406#_M1022_g
+ N_A_888_406#_c_561_n N_A_888_406#_c_562_n N_A_888_406#_c_583_p
+ N_A_888_406#_c_547_n N_A_888_406#_c_548_n N_A_888_406#_c_564_n
+ N_A_888_406#_c_549_n N_A_888_406#_c_594_p N_A_888_406#_c_565_n
+ N_A_888_406#_c_550_n N_A_888_406#_c_551_n N_A_888_406#_c_552_n
+ N_A_888_406#_c_568_n N_A_888_406#_c_553_n
+ PM_SKY130_FD_SC_MS__DLRTN_4%A_888_406#
x_PM_SKY130_FD_SC_MS__DLRTN_4%A_642_392# N_A_642_392#_M1017_d
+ N_A_642_392#_M1028_d N_A_642_392#_M1012_g N_A_642_392#_c_722_n
+ N_A_642_392#_M1009_g N_A_642_392#_M1016_g N_A_642_392#_c_723_n
+ N_A_642_392#_M1026_g N_A_642_392#_c_731_n N_A_642_392#_c_732_n
+ N_A_642_392#_c_733_n N_A_642_392#_c_734_n N_A_642_392#_c_765_n
+ N_A_642_392#_c_724_n N_A_642_392#_c_725_n N_A_642_392#_c_726_n
+ N_A_642_392#_c_727_n N_A_642_392#_c_728_n
+ PM_SKY130_FD_SC_MS__DLRTN_4%A_642_392#
x_PM_SKY130_FD_SC_MS__DLRTN_4%RESET_B N_RESET_B_M1014_g N_RESET_B_c_839_n
+ N_RESET_B_M1002_g N_RESET_B_c_840_n N_RESET_B_M1021_g N_RESET_B_M1029_g
+ RESET_B RESET_B RESET_B N_RESET_B_c_843_n PM_SKY130_FD_SC_MS__DLRTN_4%RESET_B
x_PM_SKY130_FD_SC_MS__DLRTN_4%VPWR N_VPWR_M1013_d N_VPWR_M1008_d N_VPWR_M1010_d
+ N_VPWR_M1016_s N_VPWR_M1029_s N_VPWR_M1023_d N_VPWR_M1027_d N_VPWR_c_895_n
+ N_VPWR_c_896_n N_VPWR_c_897_n N_VPWR_c_898_n N_VPWR_c_899_n N_VPWR_c_900_n
+ N_VPWR_c_901_n N_VPWR_c_902_n N_VPWR_c_903_n N_VPWR_c_904_n N_VPWR_c_905_n
+ N_VPWR_c_906_n N_VPWR_c_907_n VPWR N_VPWR_c_908_n N_VPWR_c_909_n
+ N_VPWR_c_910_n N_VPWR_c_911_n N_VPWR_c_912_n N_VPWR_c_894_n
+ PM_SKY130_FD_SC_MS__DLRTN_4%VPWR
x_PM_SKY130_FD_SC_MS__DLRTN_4%Q N_Q_M1001_s N_Q_M1011_s N_Q_M1019_s N_Q_M1025_s
+ N_Q_c_1016_n N_Q_c_1011_n N_Q_c_1023_n N_Q_c_1005_n N_Q_c_1006_n N_Q_c_1012_n
+ N_Q_c_1007_n N_Q_c_1013_n N_Q_c_1014_n Q Q Q N_Q_c_1010_n
+ PM_SKY130_FD_SC_MS__DLRTN_4%Q
x_PM_SKY130_FD_SC_MS__DLRTN_4%VGND N_VGND_M1024_d N_VGND_M1020_d N_VGND_M1015_d
+ N_VGND_M1002_s N_VGND_M1001_d N_VGND_M1004_d N_VGND_M1022_d N_VGND_c_1079_n
+ N_VGND_c_1080_n N_VGND_c_1081_n N_VGND_c_1082_n N_VGND_c_1083_n
+ N_VGND_c_1084_n N_VGND_c_1085_n N_VGND_c_1086_n N_VGND_c_1087_n
+ N_VGND_c_1088_n VGND N_VGND_c_1089_n N_VGND_c_1090_n N_VGND_c_1091_n
+ N_VGND_c_1092_n N_VGND_c_1093_n N_VGND_c_1094_n N_VGND_c_1095_n
+ N_VGND_c_1096_n N_VGND_c_1097_n N_VGND_c_1098_n N_VGND_c_1099_n
+ PM_SKY130_FD_SC_MS__DLRTN_4%VGND
x_PM_SKY130_FD_SC_MS__DLRTN_4%A_1035_74# N_A_1035_74#_M1009_d
+ N_A_1035_74#_M1026_d N_A_1035_74#_M1021_d N_A_1035_74#_c_1198_n
+ N_A_1035_74#_c_1199_n N_A_1035_74#_c_1200_n N_A_1035_74#_c_1207_n
+ N_A_1035_74#_c_1218_n N_A_1035_74#_c_1221_n N_A_1035_74#_c_1201_n
+ N_A_1035_74#_c_1202_n PM_SKY130_FD_SC_MS__DLRTN_4%A_1035_74#
cc_1 VNB N_D_M1024_g 0.0308051f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.955
cc_2 VNB D 0.0020826f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_3 VNB N_D_c_174_n 0.0209411f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_4 VNB N_GATE_N_M1003_g 0.0293544f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.39
cc_5 VNB N_GATE_N_c_206_n 0.0194391f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_6 VNB N_A_232_98#_M1020_g 0.0274357f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_7 VNB N_A_232_98#_M1017_g 0.0488807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_232_98#_c_244_n 0.0283723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_232_98#_c_245_n 0.0133008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_232_98#_c_246_n 0.0101216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_232_98#_c_247_n 0.00493468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_232_98#_c_248_n 0.00341963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_136#_c_361_n 0.0436194f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.39
cc_14 VNB N_A_27_136#_c_362_n 0.0319058f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.615
cc_15 VNB N_A_27_136#_c_363_n 0.016625f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_16 VNB N_A_27_136#_c_364_n 0.00939626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_136#_c_365_n 0.00892374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_136#_c_366_n 0.0118837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_136#_c_367_n 0.00172991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_136#_c_368_n 0.013789f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_136#_c_369_n 0.0194302f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_348_392#_M1006_g 0.0321721f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_23 VNB N_A_348_392#_c_443_n 0.00310365f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_24 VNB N_A_348_392#_c_444_n 0.0176286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_348_392#_c_445_n 0.00312853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_348_392#_c_446_n 0.0216723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_348_392#_c_447_n 0.0311398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_348_392#_c_448_n 0.00437346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_888_406#_M1015_g 0.064354f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_30 VNB N_A_888_406#_M1019_g 0.00144121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_888_406#_c_538_n 0.0098246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_888_406#_c_539_n 0.0111631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_888_406#_M1001_g 0.0237608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_888_406#_M1023_g 0.00148032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_888_406#_M1004_g 0.0203648f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_888_406#_M1025_g 0.0017134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_888_406#_M1011_g 0.0203434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_888_406#_M1027_g 0.00182109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_888_406#_M1022_g 0.0232586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_888_406#_c_547_n 0.00197983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_888_406#_c_548_n 0.00514849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_888_406#_c_549_n 0.0016809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_888_406#_c_550_n 0.00244605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_888_406#_c_551_n 0.00378547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_888_406#_c_552_n 0.00283662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_888_406#_c_553_n 0.0828531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_642_392#_c_722_n 0.0192663f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.615
cc_48 VNB N_A_642_392#_c_723_n 0.0163945f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.615
cc_49 VNB N_A_642_392#_c_724_n 0.0130544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_642_392#_c_725_n 0.00257326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_642_392#_c_726_n 0.0163589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_642_392#_c_727_n 0.00339515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_642_392#_c_728_n 0.101808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_RESET_B_M1014_g 0.00370409f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.955
cc_55 VNB N_RESET_B_c_839_n 0.016867f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.78
cc_56 VNB N_RESET_B_c_840_n 0.0211591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_RESET_B_M1029_g 0.00392107f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_58 VNB RESET_B 0.0270615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_RESET_B_c_843_n 0.0651696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VPWR_c_894_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_Q_c_1005_n 0.00180794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_Q_c_1006_n 0.00165555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_Q_c_1007_n 0.0017948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB Q 0.0171365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB Q 0.0270077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_Q_c_1010_n 0.00306278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1079_n 0.0205322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1080_n 0.00928694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1081_n 0.00340259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1082_n 0.0187851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1083_n 0.0106146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1084_n 0.00250542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1085_n 0.012003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1086_n 0.0195864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1087_n 0.0442338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1088_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1089_n 0.0197505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1090_n 0.0374084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1091_n 0.0150459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1092_n 0.0150459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1093_n 0.00631593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1094_n 0.0373356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1095_n 0.0305963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1096_n 0.00601668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1097_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1098_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1099_n 0.523604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1035_74#_c_1198_n 0.0057158f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_89 VNB N_A_1035_74#_c_1199_n 0.00450979f $X=-0.19 $Y=-0.245 $X2=0.587
+ $Y2=1.45
cc_90 VNB N_A_1035_74#_c_1200_n 0.00418613f $X=-0.19 $Y=-0.245 $X2=0.587
+ $Y2=1.78
cc_91 VNB N_A_1035_74#_c_1201_n 0.00179342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1035_74#_c_1202_n 0.0060844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VPB N_D_M1013_g 0.0298454f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.39
cc_94 VPB D 0.00118268f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_95 VPB N_D_c_174_n 0.0127318f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_96 VPB N_GATE_N_M1007_g 0.0288566f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.955
cc_97 VPB N_GATE_N_c_206_n 0.0126865f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_98 VPB N_A_232_98#_M1008_g 0.0299536f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_99 VPB N_A_232_98#_M1017_g 0.0256345f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_232_98#_M1000_g 0.0250425f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_232_98#_c_244_n 0.0188163f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_232_98#_c_245_n 0.00334934f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_232_98#_c_254_n 0.0124407f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_232_98#_c_255_n 0.00647598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_232_98#_c_256_n 0.00569032f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_232_98#_c_257_n 0.00733803f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_232_98#_c_258_n 0.00560999f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_232_98#_c_259_n 0.0441499f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_232_98#_c_260_n 0.0107399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_232_98#_c_261_n 0.00380672f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_232_98#_c_247_n 0.00748064f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_27_136#_c_361_n 0.00497416f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=2.39
cc_113 VPB N_A_27_136#_M1005_g 0.0303887f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_114 VPB N_A_27_136#_c_367_n 0.00161498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_27_136#_c_373_n 0.0469784f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_27_136#_c_369_n 0.0138202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_348_392#_M1028_g 0.0232753f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_118 VPB N_A_348_392#_c_443_n 0.00309752f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_119 VPB N_A_348_392#_c_451_n 0.0132079f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_348_392#_c_452_n 8.9109e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_348_392#_c_444_n 0.0121213f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_348_392#_c_454_n 0.0021356f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_888_406#_M1010_g 0.0273942f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_124 VPB N_A_888_406#_M1015_g 0.00498254f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_125 VPB N_A_888_406#_c_556_n 0.00661911f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_126 VPB N_A_888_406#_M1019_g 0.0231542f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_888_406#_M1023_g 0.0225055f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_888_406#_M1025_g 0.0236122f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_888_406#_M1027_g 0.0260681f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_888_406#_c_561_n 0.0122435f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_888_406#_c_562_n 0.0300752f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_888_406#_c_548_n 0.00473446f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_888_406#_c_564_n 0.00625609f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_888_406#_c_565_n 0.00239598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_888_406#_c_551_n 0.00791229f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_888_406#_c_552_n 0.00112048f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_888_406#_c_568_n 0.019113f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_642_392#_M1012_g 0.0318905f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_139 VPB N_A_642_392#_M1016_g 0.028201f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_140 VPB N_A_642_392#_c_731_n 0.00185598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_642_392#_c_732_n 0.00332253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_642_392#_c_733_n 0.0295182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_642_392#_c_734_n 0.00146234f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_642_392#_c_727_n 3.15148e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_642_392#_c_728_n 0.0336549f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_RESET_B_M1014_g 0.0363653f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.955
cc_147 VPB N_RESET_B_M1029_g 0.0375452f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_148 VPB N_VPWR_c_895_n 0.0305181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_896_n 0.0187933f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_897_n 0.0102803f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_898_n 0.0110347f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_899_n 0.00510895f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_900_n 0.0155055f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_901_n 0.0407013f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_902_n 0.0184575f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_903_n 0.0346264f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_904_n 0.0205172f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_905_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_906_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_907_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_908_n 0.0183788f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_909_n 0.0267333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_910_n 0.0554149f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_911_n 0.0252234f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_912_n 0.00628274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_894_n 0.125449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_Q_c_1011_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.587 $Y2=1.78
cc_168 VPB N_Q_c_1012_n 0.00326394f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_Q_c_1013_n 0.0141772f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_Q_c_1014_n 0.00292772f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB Q 0.00746653f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 N_D_M1013_g N_GATE_N_M1007_g 0.0141966f $X=0.535 $Y=2.39 $X2=0 $Y2=0
cc_173 N_D_M1024_g N_GATE_N_M1003_g 0.0253063f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_174 D GATE_N 0.0264214f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_175 N_D_c_174_n GATE_N 3.64022e-19 $X=0.59 $Y=1.615 $X2=0 $Y2=0
cc_176 D N_GATE_N_c_206_n 0.00190882f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_177 N_D_c_174_n N_GATE_N_c_206_n 0.0206217f $X=0.59 $Y=1.615 $X2=0 $Y2=0
cc_178 N_D_M1024_g N_A_232_98#_c_246_n 0.00111637f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_179 N_D_M1024_g N_A_27_136#_c_364_n 0.00496207f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_180 N_D_M1024_g N_A_27_136#_c_365_n 0.0102665f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_181 D N_A_27_136#_c_365_n 0.00871068f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_182 N_D_c_174_n N_A_27_136#_c_365_n 0.00288484f $X=0.59 $Y=1.615 $X2=0 $Y2=0
cc_183 N_D_M1024_g N_A_27_136#_c_366_n 0.00286883f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_184 N_D_M1024_g N_A_27_136#_c_368_n 0.00636483f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_185 D N_A_27_136#_c_368_n 0.00131568f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_186 N_D_M1013_g N_A_27_136#_c_373_n 0.0149549f $X=0.535 $Y=2.39 $X2=0 $Y2=0
cc_187 D N_A_27_136#_c_373_n 0.00400158f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_188 N_D_c_174_n N_A_27_136#_c_373_n 7.86724e-19 $X=0.59 $Y=1.615 $X2=0 $Y2=0
cc_189 N_D_M1024_g N_A_27_136#_c_369_n 0.0126381f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_190 N_D_M1013_g N_A_27_136#_c_369_n 0.00408775f $X=0.535 $Y=2.39 $X2=0 $Y2=0
cc_191 D N_A_27_136#_c_369_n 0.0250413f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_192 N_D_M1013_g N_VPWR_c_895_n 0.00460946f $X=0.535 $Y=2.39 $X2=0 $Y2=0
cc_193 D N_VPWR_c_895_n 0.0136154f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_194 N_D_c_174_n N_VPWR_c_895_n 0.00253923f $X=0.59 $Y=1.615 $X2=0 $Y2=0
cc_195 N_D_M1013_g N_VPWR_c_909_n 0.00546844f $X=0.535 $Y=2.39 $X2=0 $Y2=0
cc_196 N_D_M1013_g N_VPWR_c_894_n 0.00599321f $X=0.535 $Y=2.39 $X2=0 $Y2=0
cc_197 N_D_M1024_g N_VGND_c_1089_n 0.00301898f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_198 N_D_M1024_g N_VGND_c_1099_n 0.00454494f $X=0.495 $Y=0.955 $X2=0 $Y2=0
cc_199 N_GATE_N_M1003_g N_A_232_98#_c_244_n 8.31894e-19 $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_200 GATE_N N_A_232_98#_c_244_n 3.22315e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_201 N_GATE_N_c_206_n N_A_232_98#_c_244_n 0.0158557f $X=1.13 $Y=1.615 $X2=0
+ $Y2=0
cc_202 N_GATE_N_M1003_g N_A_232_98#_c_246_n 0.00648185f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_203 GATE_N N_A_232_98#_c_246_n 0.0105236f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_204 N_GATE_N_c_206_n N_A_232_98#_c_246_n 0.00313382f $X=1.13 $Y=1.615 $X2=0
+ $Y2=0
cc_205 N_GATE_N_M1007_g N_A_232_98#_c_255_n 0.00815489f $X=1.085 $Y=2.39 $X2=0
+ $Y2=0
cc_206 N_GATE_N_M1007_g N_A_232_98#_c_257_n 0.00344538f $X=1.085 $Y=2.39 $X2=0
+ $Y2=0
cc_207 N_GATE_N_M1007_g N_A_232_98#_c_260_n 0.00358739f $X=1.085 $Y=2.39 $X2=0
+ $Y2=0
cc_208 GATE_N N_A_232_98#_c_260_n 0.0120132f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_209 N_GATE_N_c_206_n N_A_232_98#_c_260_n 0.00290121f $X=1.13 $Y=1.615 $X2=0
+ $Y2=0
cc_210 N_GATE_N_M1007_g N_A_232_98#_c_261_n 0.00522341f $X=1.085 $Y=2.39 $X2=0
+ $Y2=0
cc_211 GATE_N N_A_232_98#_c_247_n 0.0262364f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_212 N_GATE_N_c_206_n N_A_232_98#_c_247_n 0.00256913f $X=1.13 $Y=1.615 $X2=0
+ $Y2=0
cc_213 N_GATE_N_M1003_g N_A_232_98#_c_248_n 0.00568622f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_214 N_GATE_N_M1003_g N_A_27_136#_c_364_n 0.00189038f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_215 N_GATE_N_M1003_g N_A_27_136#_c_365_n 0.0160857f $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_216 GATE_N N_A_27_136#_c_365_n 0.00350057f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_217 N_GATE_N_M1003_g N_A_348_392#_c_448_n 3.18666e-19 $X=1.085 $Y=0.86 $X2=0
+ $Y2=0
cc_218 N_GATE_N_M1007_g N_A_348_392#_c_454_n 8.4935e-19 $X=1.085 $Y=2.39 $X2=0
+ $Y2=0
cc_219 N_GATE_N_M1007_g N_VPWR_c_895_n 0.0046091f $X=1.085 $Y=2.39 $X2=0 $Y2=0
cc_220 N_GATE_N_c_206_n N_VPWR_c_895_n 3.99972e-19 $X=1.13 $Y=1.615 $X2=0 $Y2=0
cc_221 N_GATE_N_M1007_g N_VPWR_c_903_n 0.00546038f $X=1.085 $Y=2.39 $X2=0 $Y2=0
cc_222 N_GATE_N_M1007_g N_VPWR_c_894_n 0.00599321f $X=1.085 $Y=2.39 $X2=0 $Y2=0
cc_223 N_GATE_N_M1003_g N_VGND_c_1079_n 0.00546687f $X=1.085 $Y=0.86 $X2=0 $Y2=0
cc_224 N_GATE_N_M1003_g N_VGND_c_1094_n 0.0038134f $X=1.085 $Y=0.86 $X2=0 $Y2=0
cc_225 N_GATE_N_M1003_g N_VGND_c_1099_n 0.00508379f $X=1.085 $Y=0.86 $X2=0 $Y2=0
cc_226 N_A_232_98#_M1020_g N_A_27_136#_c_361_n 0.0186166f $X=2.18 $Y=0.86 $X2=0
+ $Y2=0
cc_227 N_A_232_98#_c_245_n N_A_27_136#_c_361_n 0.0042319f $X=2.02 $Y=1.42 $X2=0
+ $Y2=0
cc_228 N_A_232_98#_c_245_n N_A_27_136#_M1005_g 0.0332771f $X=2.02 $Y=1.42 $X2=0
+ $Y2=0
cc_229 N_A_232_98#_c_256_n N_A_27_136#_M1005_g 0.0150059f $X=3.87 $Y=2.685 $X2=0
+ $Y2=0
cc_230 N_A_232_98#_M1017_g N_A_27_136#_c_363_n 0.0548797f $X=3.645 $Y=0.69 $X2=0
+ $Y2=0
cc_231 N_A_232_98#_M1003_d N_A_27_136#_c_365_n 0.0113826f $X=1.16 $Y=0.49 $X2=0
+ $Y2=0
cc_232 N_A_232_98#_M1020_g N_A_27_136#_c_365_n 0.016975f $X=2.18 $Y=0.86 $X2=0
+ $Y2=0
cc_233 N_A_232_98#_c_244_n N_A_27_136#_c_365_n 0.00121652f $X=2.02 $Y=1.585
+ $X2=0 $Y2=0
cc_234 N_A_232_98#_c_246_n N_A_27_136#_c_365_n 0.0339256f $X=1.46 $Y=1.125 $X2=0
+ $Y2=0
cc_235 N_A_232_98#_c_247_n N_A_27_136#_c_365_n 0.00498546f $X=1.7 $Y=1.585 $X2=0
+ $Y2=0
cc_236 N_A_232_98#_M1020_g N_A_27_136#_c_367_n 0.0104291f $X=2.18 $Y=0.86 $X2=0
+ $Y2=0
cc_237 N_A_232_98#_c_256_n N_A_348_392#_M1008_s 0.00849365f $X=3.87 $Y=2.685
+ $X2=0 $Y2=0
cc_238 N_A_232_98#_M1017_g N_A_348_392#_M1028_g 0.0390614f $X=3.645 $Y=0.69
+ $X2=0 $Y2=0
cc_239 N_A_232_98#_c_256_n N_A_348_392#_M1028_g 0.0142695f $X=3.87 $Y=2.685
+ $X2=0 $Y2=0
cc_240 N_A_232_98#_M1017_g N_A_348_392#_M1006_g 0.0217567f $X=3.645 $Y=0.69
+ $X2=0 $Y2=0
cc_241 N_A_232_98#_M1008_g N_A_348_392#_c_443_n 0.00608517f $X=2.11 $Y=2.38
+ $X2=0 $Y2=0
cc_242 N_A_232_98#_M1020_g N_A_348_392#_c_443_n 0.0059554f $X=2.18 $Y=0.86 $X2=0
+ $Y2=0
cc_243 N_A_232_98#_c_245_n N_A_348_392#_c_443_n 0.0129609f $X=2.02 $Y=1.42 $X2=0
+ $Y2=0
cc_244 N_A_232_98#_c_261_n N_A_348_392#_c_443_n 0.00633443f $X=1.387 $Y=1.95
+ $X2=0 $Y2=0
cc_245 N_A_232_98#_c_247_n N_A_348_392#_c_443_n 0.0239603f $X=1.7 $Y=1.585 $X2=0
+ $Y2=0
cc_246 N_A_232_98#_c_248_n N_A_348_392#_c_443_n 0.00698482f $X=1.662 $Y=1.42
+ $X2=0 $Y2=0
cc_247 N_A_232_98#_M1017_g N_A_348_392#_c_451_n 6.53392e-19 $X=3.645 $Y=0.69
+ $X2=0 $Y2=0
cc_248 N_A_232_98#_c_245_n N_A_348_392#_c_451_n 0.00171935f $X=2.02 $Y=1.42
+ $X2=0 $Y2=0
cc_249 N_A_232_98#_c_256_n N_A_348_392#_c_451_n 0.023167f $X=3.87 $Y=2.685 $X2=0
+ $Y2=0
cc_250 N_A_232_98#_M1017_g N_A_348_392#_c_452_n 0.00172099f $X=3.645 $Y=0.69
+ $X2=0 $Y2=0
cc_251 N_A_232_98#_M1017_g N_A_348_392#_c_444_n 0.021052f $X=3.645 $Y=0.69 $X2=0
+ $Y2=0
cc_252 N_A_232_98#_M1017_g N_A_348_392#_c_446_n 0.0227514f $X=3.645 $Y=0.69
+ $X2=0 $Y2=0
cc_253 N_A_232_98#_M1017_g N_A_348_392#_c_447_n 0.021337f $X=3.645 $Y=0.69 $X2=0
+ $Y2=0
cc_254 N_A_232_98#_c_259_n N_A_348_392#_c_447_n 0.00489746f $X=4.035 $Y=2.195
+ $X2=0 $Y2=0
cc_255 N_A_232_98#_M1020_g N_A_348_392#_c_448_n 0.00658026f $X=2.18 $Y=0.86
+ $X2=0 $Y2=0
cc_256 N_A_232_98#_c_244_n N_A_348_392#_c_448_n 0.00532403f $X=2.02 $Y=1.585
+ $X2=0 $Y2=0
cc_257 N_A_232_98#_c_245_n N_A_348_392#_c_448_n 3.30391e-19 $X=2.02 $Y=1.42
+ $X2=0 $Y2=0
cc_258 N_A_232_98#_c_246_n N_A_348_392#_c_448_n 0.0218242f $X=1.46 $Y=1.125
+ $X2=0 $Y2=0
cc_259 N_A_232_98#_c_247_n N_A_348_392#_c_448_n 0.0049796f $X=1.7 $Y=1.585 $X2=0
+ $Y2=0
cc_260 N_A_232_98#_M1008_g N_A_348_392#_c_454_n 0.0191654f $X=2.11 $Y=2.38 $X2=0
+ $Y2=0
cc_261 N_A_232_98#_c_244_n N_A_348_392#_c_454_n 0.00505569f $X=2.02 $Y=1.585
+ $X2=0 $Y2=0
cc_262 N_A_232_98#_c_256_n N_A_348_392#_c_454_n 0.0262142f $X=3.87 $Y=2.685
+ $X2=0 $Y2=0
cc_263 N_A_232_98#_c_261_n N_A_348_392#_c_454_n 0.0439828f $X=1.387 $Y=1.95
+ $X2=0 $Y2=0
cc_264 N_A_232_98#_c_247_n N_A_348_392#_c_454_n 0.00527154f $X=1.7 $Y=1.585
+ $X2=0 $Y2=0
cc_265 N_A_232_98#_M1000_g N_A_888_406#_M1010_g 0.0106116f $X=3.66 $Y=2.73 $X2=0
+ $Y2=0
cc_266 N_A_232_98#_c_256_n N_A_888_406#_M1010_g 0.00258283f $X=3.87 $Y=2.685
+ $X2=0 $Y2=0
cc_267 N_A_232_98#_c_258_n N_A_888_406#_M1010_g 0.00603301f $X=4.035 $Y=2.195
+ $X2=0 $Y2=0
cc_268 N_A_232_98#_c_258_n N_A_888_406#_c_561_n 0.0198487f $X=4.035 $Y=2.195
+ $X2=0 $Y2=0
cc_269 N_A_232_98#_c_259_n N_A_888_406#_c_561_n 0.00136396f $X=4.035 $Y=2.195
+ $X2=0 $Y2=0
cc_270 N_A_232_98#_c_258_n N_A_888_406#_c_562_n 4.19484e-19 $X=4.035 $Y=2.195
+ $X2=0 $Y2=0
cc_271 N_A_232_98#_c_259_n N_A_888_406#_c_562_n 0.0185169f $X=4.035 $Y=2.195
+ $X2=0 $Y2=0
cc_272 N_A_232_98#_c_256_n N_A_642_392#_M1028_d 0.00652375f $X=3.87 $Y=2.685
+ $X2=0 $Y2=0
cc_273 N_A_232_98#_M1000_g N_A_642_392#_c_731_n 0.00414328f $X=3.66 $Y=2.73
+ $X2=0 $Y2=0
cc_274 N_A_232_98#_c_254_n N_A_642_392#_c_731_n 0.00409691f $X=3.66 $Y=2.195
+ $X2=0 $Y2=0
cc_275 N_A_232_98#_c_256_n N_A_642_392#_c_731_n 0.0322626f $X=3.87 $Y=2.685
+ $X2=0 $Y2=0
cc_276 N_A_232_98#_c_258_n N_A_642_392#_c_731_n 0.0135326f $X=4.035 $Y=2.195
+ $X2=0 $Y2=0
cc_277 N_A_232_98#_M1017_g N_A_642_392#_c_732_n 0.00920521f $X=3.645 $Y=0.69
+ $X2=0 $Y2=0
cc_278 N_A_232_98#_c_254_n N_A_642_392#_c_732_n 0.00727416f $X=3.66 $Y=2.195
+ $X2=0 $Y2=0
cc_279 N_A_232_98#_c_258_n N_A_642_392#_c_732_n 0.016391f $X=4.035 $Y=2.195
+ $X2=0 $Y2=0
cc_280 N_A_232_98#_M1017_g N_A_642_392#_c_733_n 0.00544814f $X=3.645 $Y=0.69
+ $X2=0 $Y2=0
cc_281 N_A_232_98#_c_254_n N_A_642_392#_c_733_n 0.00577048f $X=3.66 $Y=2.195
+ $X2=0 $Y2=0
cc_282 N_A_232_98#_c_258_n N_A_642_392#_c_733_n 0.0262124f $X=4.035 $Y=2.195
+ $X2=0 $Y2=0
cc_283 N_A_232_98#_c_259_n N_A_642_392#_c_733_n 0.0014355f $X=4.035 $Y=2.195
+ $X2=0 $Y2=0
cc_284 N_A_232_98#_M1017_g N_A_642_392#_c_734_n 0.00468408f $X=3.645 $Y=0.69
+ $X2=0 $Y2=0
cc_285 N_A_232_98#_M1017_g N_A_642_392#_c_725_n 0.00113438f $X=3.645 $Y=0.69
+ $X2=0 $Y2=0
cc_286 N_A_232_98#_c_256_n N_VPWR_M1008_d 0.00997142f $X=3.87 $Y=2.685 $X2=0
+ $Y2=0
cc_287 N_A_232_98#_c_257_n N_VPWR_c_895_n 0.0103557f $X=1.63 $Y=2.685 $X2=0
+ $Y2=0
cc_288 N_A_232_98#_c_260_n N_VPWR_c_895_n 0.0265799f $X=1.31 $Y=2.115 $X2=0
+ $Y2=0
cc_289 N_A_232_98#_c_256_n N_VPWR_c_902_n 0.0242954f $X=3.87 $Y=2.685 $X2=0
+ $Y2=0
cc_290 N_A_232_98#_M1008_g N_VPWR_c_903_n 0.00425923f $X=2.11 $Y=2.38 $X2=0
+ $Y2=0
cc_291 N_A_232_98#_c_256_n N_VPWR_c_903_n 0.0118623f $X=3.87 $Y=2.685 $X2=0
+ $Y2=0
cc_292 N_A_232_98#_c_257_n N_VPWR_c_903_n 0.0133379f $X=1.63 $Y=2.685 $X2=0
+ $Y2=0
cc_293 N_A_232_98#_M1000_g N_VPWR_c_910_n 0.00508505f $X=3.66 $Y=2.73 $X2=0
+ $Y2=0
cc_294 N_A_232_98#_c_256_n N_VPWR_c_910_n 0.0305694f $X=3.87 $Y=2.685 $X2=0
+ $Y2=0
cc_295 N_A_232_98#_c_256_n N_VPWR_c_911_n 0.0063817f $X=3.87 $Y=2.685 $X2=0
+ $Y2=0
cc_296 N_A_232_98#_M1008_g N_VPWR_c_894_n 0.00595788f $X=2.11 $Y=2.38 $X2=0
+ $Y2=0
cc_297 N_A_232_98#_M1000_g N_VPWR_c_894_n 0.00647345f $X=3.66 $Y=2.73 $X2=0
+ $Y2=0
cc_298 N_A_232_98#_c_256_n N_VPWR_c_894_n 0.0680058f $X=3.87 $Y=2.685 $X2=0
+ $Y2=0
cc_299 N_A_232_98#_c_257_n N_VPWR_c_894_n 0.0161941f $X=1.63 $Y=2.685 $X2=0
+ $Y2=0
cc_300 N_A_232_98#_c_256_n A_564_392# 0.00327529f $X=3.87 $Y=2.685 $X2=-0.19
+ $Y2=-0.245
cc_301 N_A_232_98#_c_256_n A_750_504# 0.0119402f $X=3.87 $Y=2.685 $X2=-0.19
+ $Y2=-0.245
cc_302 N_A_232_98#_c_258_n A_750_504# 0.00288822f $X=4.035 $Y=2.195 $X2=-0.19
+ $Y2=-0.245
cc_303 N_A_232_98#_M1017_g N_VGND_c_1087_n 0.00461464f $X=3.645 $Y=0.69 $X2=0
+ $Y2=0
cc_304 N_A_232_98#_M1020_g N_VGND_c_1094_n 0.0038134f $X=2.18 $Y=0.86 $X2=0
+ $Y2=0
cc_305 N_A_232_98#_M1020_g N_VGND_c_1095_n 0.0060117f $X=2.18 $Y=0.86 $X2=0
+ $Y2=0
cc_306 N_A_232_98#_M1020_g N_VGND_c_1099_n 0.00508379f $X=2.18 $Y=0.86 $X2=0
+ $Y2=0
cc_307 N_A_232_98#_M1017_g N_VGND_c_1099_n 0.00909529f $X=3.645 $Y=0.69 $X2=0
+ $Y2=0
cc_308 N_A_27_136#_c_365_n N_A_348_392#_M1020_s 0.00727646f $X=2.49 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_309 N_A_27_136#_M1005_g N_A_348_392#_M1028_g 0.0532408f $X=2.73 $Y=2.46 $X2=0
+ $Y2=0
cc_310 N_A_27_136#_c_361_n N_A_348_392#_c_443_n 0.00147873f $X=2.73 $Y=1.67
+ $X2=0 $Y2=0
cc_311 N_A_27_136#_M1005_g N_A_348_392#_c_443_n 0.00407445f $X=2.73 $Y=2.46
+ $X2=0 $Y2=0
cc_312 N_A_27_136#_c_367_n N_A_348_392#_c_443_n 0.0205894f $X=2.655 $Y=1.505
+ $X2=0 $Y2=0
cc_313 N_A_27_136#_c_361_n N_A_348_392#_c_451_n 9.68515e-19 $X=2.73 $Y=1.67
+ $X2=0 $Y2=0
cc_314 N_A_27_136#_M1005_g N_A_348_392#_c_451_n 0.0146091f $X=2.73 $Y=2.46 $X2=0
+ $Y2=0
cc_315 N_A_27_136#_c_362_n N_A_348_392#_c_451_n 0.00421244f $X=3.18 $Y=1.16
+ $X2=0 $Y2=0
cc_316 N_A_27_136#_c_367_n N_A_348_392#_c_451_n 0.0189066f $X=2.655 $Y=1.505
+ $X2=0 $Y2=0
cc_317 N_A_27_136#_c_361_n N_A_348_392#_c_452_n 0.0022027f $X=2.73 $Y=1.67 $X2=0
+ $Y2=0
cc_318 N_A_27_136#_c_367_n N_A_348_392#_c_452_n 0.00947434f $X=2.655 $Y=1.505
+ $X2=0 $Y2=0
cc_319 N_A_27_136#_c_361_n N_A_348_392#_c_444_n 0.0532408f $X=2.73 $Y=1.67 $X2=0
+ $Y2=0
cc_320 N_A_27_136#_c_362_n N_A_348_392#_c_444_n 0.0194807f $X=3.18 $Y=1.16 $X2=0
+ $Y2=0
cc_321 N_A_27_136#_c_367_n N_A_348_392#_c_444_n 6.17168e-19 $X=2.655 $Y=1.505
+ $X2=0 $Y2=0
cc_322 N_A_27_136#_c_361_n N_A_348_392#_c_445_n 0.00471724f $X=2.73 $Y=1.67
+ $X2=0 $Y2=0
cc_323 N_A_27_136#_c_362_n N_A_348_392#_c_445_n 0.0195998f $X=3.18 $Y=1.16 $X2=0
+ $Y2=0
cc_324 N_A_27_136#_c_367_n N_A_348_392#_c_445_n 0.0231983f $X=2.655 $Y=1.505
+ $X2=0 $Y2=0
cc_325 N_A_27_136#_c_365_n N_A_348_392#_c_448_n 0.0255532f $X=2.49 $Y=0.745
+ $X2=0 $Y2=0
cc_326 N_A_27_136#_c_367_n N_A_348_392#_c_448_n 0.0132245f $X=2.655 $Y=1.505
+ $X2=0 $Y2=0
cc_327 N_A_27_136#_M1005_g N_A_642_392#_c_731_n 8.09912e-19 $X=2.73 $Y=2.46
+ $X2=0 $Y2=0
cc_328 N_A_27_136#_c_373_n N_VPWR_c_895_n 0.0354172f $X=0.31 $Y=2.115 $X2=0
+ $Y2=0
cc_329 N_A_27_136#_M1005_g N_VPWR_c_902_n 0.00590973f $X=2.73 $Y=2.46 $X2=0
+ $Y2=0
cc_330 N_A_27_136#_c_373_n N_VPWR_c_909_n 0.0106578f $X=0.31 $Y=2.115 $X2=0
+ $Y2=0
cc_331 N_A_27_136#_M1005_g N_VPWR_c_910_n 0.00381426f $X=2.73 $Y=2.46 $X2=0
+ $Y2=0
cc_332 N_A_27_136#_M1005_g N_VPWR_c_894_n 0.00477601f $X=2.73 $Y=2.46 $X2=0
+ $Y2=0
cc_333 N_A_27_136#_c_373_n N_VPWR_c_894_n 0.01295f $X=0.31 $Y=2.115 $X2=0 $Y2=0
cc_334 N_A_27_136#_c_365_n N_VGND_M1024_d 0.0128101f $X=2.49 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_335 N_A_27_136#_c_365_n N_VGND_M1020_d 0.0184416f $X=2.49 $Y=0.745 $X2=0
+ $Y2=0
cc_336 N_A_27_136#_c_367_n N_VGND_M1020_d 0.00868742f $X=2.655 $Y=1.505 $X2=0
+ $Y2=0
cc_337 N_A_27_136#_c_365_n N_VGND_c_1079_n 0.0252207f $X=2.49 $Y=0.745 $X2=0
+ $Y2=0
cc_338 N_A_27_136#_c_363_n N_VGND_c_1087_n 0.00461464f $X=3.255 $Y=1.085 $X2=0
+ $Y2=0
cc_339 N_A_27_136#_c_365_n N_VGND_c_1089_n 0.00286374f $X=2.49 $Y=0.745 $X2=0
+ $Y2=0
cc_340 N_A_27_136#_c_366_n N_VGND_c_1089_n 0.00683196f $X=0.445 $Y=0.745 $X2=0
+ $Y2=0
cc_341 N_A_27_136#_c_365_n N_VGND_c_1094_n 0.0206111f $X=2.49 $Y=0.745 $X2=0
+ $Y2=0
cc_342 N_A_27_136#_c_361_n N_VGND_c_1095_n 0.00827409f $X=2.73 $Y=1.67 $X2=0
+ $Y2=0
cc_343 N_A_27_136#_c_363_n N_VGND_c_1095_n 0.00826245f $X=3.255 $Y=1.085 $X2=0
+ $Y2=0
cc_344 N_A_27_136#_c_365_n N_VGND_c_1095_n 0.0415433f $X=2.49 $Y=0.745 $X2=0
+ $Y2=0
cc_345 N_A_27_136#_c_363_n N_VGND_c_1099_n 0.00913019f $X=3.255 $Y=1.085 $X2=0
+ $Y2=0
cc_346 N_A_27_136#_c_365_n N_VGND_c_1099_n 0.0464148f $X=2.49 $Y=0.745 $X2=0
+ $Y2=0
cc_347 N_A_27_136#_c_366_n N_VGND_c_1099_n 0.0106568f $X=0.445 $Y=0.745 $X2=0
+ $Y2=0
cc_348 N_A_348_392#_M1006_g N_A_888_406#_M1015_g 0.0429601f $X=4.12 $Y=0.58
+ $X2=0 $Y2=0
cc_349 N_A_348_392#_c_446_n N_A_888_406#_M1015_g 0.00125688f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_350 N_A_348_392#_c_447_n N_A_888_406#_M1015_g 0.0196496f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_351 N_A_348_392#_c_451_n N_A_642_392#_M1028_d 0.00218043f $X=3.03 $Y=2.005
+ $X2=0 $Y2=0
cc_352 N_A_348_392#_M1028_g N_A_642_392#_c_731_n 0.0040106f $X=3.12 $Y=2.46
+ $X2=0 $Y2=0
cc_353 N_A_348_392#_c_451_n N_A_642_392#_c_731_n 0.00981755f $X=3.03 $Y=2.005
+ $X2=0 $Y2=0
cc_354 N_A_348_392#_c_444_n N_A_642_392#_c_731_n 4.60641e-19 $X=3.195 $Y=1.61
+ $X2=0 $Y2=0
cc_355 N_A_348_392#_M1028_g N_A_642_392#_c_732_n 0.00323747f $X=3.12 $Y=2.46
+ $X2=0 $Y2=0
cc_356 N_A_348_392#_c_451_n N_A_642_392#_c_732_n 0.0141265f $X=3.03 $Y=2.005
+ $X2=0 $Y2=0
cc_357 N_A_348_392#_c_452_n N_A_642_392#_c_732_n 0.00467676f $X=3.195 $Y=1.61
+ $X2=0 $Y2=0
cc_358 N_A_348_392#_c_446_n N_A_642_392#_c_733_n 0.0428459f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_359 N_A_348_392#_c_447_n N_A_642_392#_c_733_n 0.00393734f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_360 N_A_348_392#_M1028_g N_A_642_392#_c_734_n 2.54769e-19 $X=3.12 $Y=2.46
+ $X2=0 $Y2=0
cc_361 N_A_348_392#_c_452_n N_A_642_392#_c_734_n 0.0146859f $X=3.195 $Y=1.61
+ $X2=0 $Y2=0
cc_362 N_A_348_392#_c_444_n N_A_642_392#_c_734_n 5.21268e-19 $X=3.195 $Y=1.61
+ $X2=0 $Y2=0
cc_363 N_A_348_392#_c_446_n N_A_642_392#_c_734_n 0.0139157f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_364 N_A_348_392#_M1006_g N_A_642_392#_c_765_n 0.00924174f $X=4.12 $Y=0.58
+ $X2=0 $Y2=0
cc_365 N_A_348_392#_M1006_g N_A_642_392#_c_724_n 0.00848162f $X=4.12 $Y=0.58
+ $X2=0 $Y2=0
cc_366 N_A_348_392#_c_446_n N_A_642_392#_c_724_n 0.0137779f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_367 N_A_348_392#_c_447_n N_A_642_392#_c_724_n 0.00145734f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_368 N_A_348_392#_M1006_g N_A_642_392#_c_725_n 0.00270114f $X=4.12 $Y=0.58
+ $X2=0 $Y2=0
cc_369 N_A_348_392#_c_446_n N_A_642_392#_c_725_n 0.0282919f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_370 N_A_348_392#_c_447_n N_A_642_392#_c_725_n 0.00266725f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_371 N_A_348_392#_c_446_n N_A_642_392#_c_726_n 0.00454193f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_372 N_A_348_392#_c_446_n N_A_642_392#_c_727_n 0.00679878f $X=4.095 $Y=1.355
+ $X2=0 $Y2=0
cc_373 N_A_348_392#_c_451_n N_VPWR_M1008_d 0.00652215f $X=3.03 $Y=2.005 $X2=0
+ $Y2=0
cc_374 N_A_348_392#_M1028_g N_VPWR_c_910_n 0.00381426f $X=3.12 $Y=2.46 $X2=0
+ $Y2=0
cc_375 N_A_348_392#_M1028_g N_VPWR_c_894_n 0.00478587f $X=3.12 $Y=2.46 $X2=0
+ $Y2=0
cc_376 N_A_348_392#_c_451_n A_564_392# 0.00175242f $X=3.03 $Y=2.005 $X2=-0.19
+ $Y2=-0.245
cc_377 N_A_348_392#_M1006_g N_VGND_c_1080_n 0.00161704f $X=4.12 $Y=0.58 $X2=0
+ $Y2=0
cc_378 N_A_348_392#_M1006_g N_VGND_c_1087_n 0.00435336f $X=4.12 $Y=0.58 $X2=0
+ $Y2=0
cc_379 N_A_348_392#_M1006_g N_VGND_c_1099_n 0.00449679f $X=4.12 $Y=0.58 $X2=0
+ $Y2=0
cc_380 N_A_888_406#_M1010_g N_A_642_392#_M1012_g 0.00628999f $X=4.53 $Y=2.73
+ $X2=0 $Y2=0
cc_381 N_A_888_406#_c_556_n N_A_642_392#_M1012_g 0.00448553f $X=4.56 $Y=1.825
+ $X2=0 $Y2=0
cc_382 N_A_888_406#_c_561_n N_A_642_392#_M1012_g 0.0250304f $X=5.49 $Y=2.195
+ $X2=0 $Y2=0
cc_383 N_A_888_406#_c_562_n N_A_642_392#_M1012_g 0.00501306f $X=4.605 $Y=2.195
+ $X2=0 $Y2=0
cc_384 N_A_888_406#_c_583_p N_A_642_392#_M1012_g 0.0112228f $X=5.655 $Y=2.03
+ $X2=0 $Y2=0
cc_385 N_A_888_406#_c_565_n N_A_642_392#_M1012_g 0.0198646f $X=5.655 $Y=2.245
+ $X2=0 $Y2=0
cc_386 N_A_888_406#_c_547_n N_A_642_392#_c_722_n 0.00270654f $X=5.75 $Y=0.81
+ $X2=0 $Y2=0
cc_387 N_A_888_406#_c_583_p N_A_642_392#_M1016_g 0.00775472f $X=5.655 $Y=2.03
+ $X2=0 $Y2=0
cc_388 N_A_888_406#_c_565_n N_A_642_392#_M1016_g 0.01416f $X=5.655 $Y=2.245
+ $X2=0 $Y2=0
cc_389 N_A_888_406#_c_547_n N_A_642_392#_c_723_n 0.00270654f $X=5.75 $Y=0.81
+ $X2=0 $Y2=0
cc_390 N_A_888_406#_M1015_g N_A_642_392#_c_733_n 0.00639399f $X=4.545 $Y=0.58
+ $X2=0 $Y2=0
cc_391 N_A_888_406#_c_556_n N_A_642_392#_c_733_n 0.00540326f $X=4.56 $Y=1.825
+ $X2=0 $Y2=0
cc_392 N_A_888_406#_c_561_n N_A_642_392#_c_733_n 0.0634347f $X=5.49 $Y=2.195
+ $X2=0 $Y2=0
cc_393 N_A_888_406#_c_562_n N_A_642_392#_c_733_n 0.00348128f $X=4.605 $Y=2.195
+ $X2=0 $Y2=0
cc_394 N_A_888_406#_c_583_p N_A_642_392#_c_733_n 0.00415403f $X=5.655 $Y=2.03
+ $X2=0 $Y2=0
cc_395 N_A_888_406#_c_594_p N_A_642_392#_c_733_n 0.00582853f $X=5.662 $Y=1.705
+ $X2=0 $Y2=0
cc_396 N_A_888_406#_c_568_n N_A_642_392#_c_733_n 0.00447383f $X=4.605 $Y=2.03
+ $X2=0 $Y2=0
cc_397 N_A_888_406#_M1015_g N_A_642_392#_c_765_n 0.00164878f $X=4.545 $Y=0.58
+ $X2=0 $Y2=0
cc_398 N_A_888_406#_M1015_g N_A_642_392#_c_724_n 0.0153705f $X=4.545 $Y=0.58
+ $X2=0 $Y2=0
cc_399 N_A_888_406#_M1015_g N_A_642_392#_c_726_n 0.00636966f $X=4.545 $Y=0.58
+ $X2=0 $Y2=0
cc_400 N_A_888_406#_c_547_n N_A_642_392#_c_726_n 0.00674443f $X=5.75 $Y=0.81
+ $X2=0 $Y2=0
cc_401 N_A_888_406#_M1015_g N_A_642_392#_c_727_n 0.00603966f $X=4.545 $Y=0.58
+ $X2=0 $Y2=0
cc_402 N_A_888_406#_c_547_n N_A_642_392#_c_727_n 0.00989338f $X=5.75 $Y=0.81
+ $X2=0 $Y2=0
cc_403 N_A_888_406#_c_594_p N_A_642_392#_c_727_n 0.00388535f $X=5.662 $Y=1.705
+ $X2=0 $Y2=0
cc_404 N_A_888_406#_M1015_g N_A_642_392#_c_728_n 0.0267316f $X=4.545 $Y=0.58
+ $X2=0 $Y2=0
cc_405 N_A_888_406#_c_556_n N_A_642_392#_c_728_n 0.00302799f $X=4.56 $Y=1.825
+ $X2=0 $Y2=0
cc_406 N_A_888_406#_c_561_n N_A_642_392#_c_728_n 0.00690333f $X=5.49 $Y=2.195
+ $X2=0 $Y2=0
cc_407 N_A_888_406#_c_547_n N_A_642_392#_c_728_n 0.0295448f $X=5.75 $Y=0.81
+ $X2=0 $Y2=0
cc_408 N_A_888_406#_c_548_n N_A_642_392#_c_728_n 0.018384f $X=6.49 $Y=1.705
+ $X2=0 $Y2=0
cc_409 N_A_888_406#_c_594_p N_A_642_392#_c_728_n 0.0208109f $X=5.662 $Y=1.705
+ $X2=0 $Y2=0
cc_410 N_A_888_406#_c_583_p N_RESET_B_M1014_g 7.37301e-19 $X=5.655 $Y=2.03 $X2=0
+ $Y2=0
cc_411 N_A_888_406#_c_548_n N_RESET_B_M1014_g 0.017283f $X=6.49 $Y=1.705 $X2=0
+ $Y2=0
cc_412 N_A_888_406#_c_564_n N_RESET_B_M1014_g 0.00604301f $X=6.655 $Y=2.245
+ $X2=0 $Y2=0
cc_413 N_A_888_406#_c_565_n N_RESET_B_M1014_g 4.48115e-19 $X=5.655 $Y=2.245
+ $X2=0 $Y2=0
cc_414 N_A_888_406#_M1019_g N_RESET_B_M1029_g 0.0161669f $X=7.485 $Y=2.4 $X2=0
+ $Y2=0
cc_415 N_A_888_406#_c_564_n N_RESET_B_M1029_g 0.0216315f $X=6.655 $Y=2.245 $X2=0
+ $Y2=0
cc_416 N_A_888_406#_c_550_n N_RESET_B_M1029_g 0.00268108f $X=6.655 $Y=1.705
+ $X2=0 $Y2=0
cc_417 N_A_888_406#_c_551_n N_RESET_B_M1029_g 0.0150612f $X=7.725 $Y=1.545 $X2=0
+ $Y2=0
cc_418 N_A_888_406#_c_539_n RESET_B 0.00505214f $X=7.575 $Y=1.555 $X2=0 $Y2=0
cc_419 N_A_888_406#_M1001_g RESET_B 0.0071116f $X=7.815 $Y=0.74 $X2=0 $Y2=0
cc_420 N_A_888_406#_c_547_n RESET_B 0.0106111f $X=5.75 $Y=0.81 $X2=0 $Y2=0
cc_421 N_A_888_406#_c_548_n RESET_B 0.0121777f $X=6.49 $Y=1.705 $X2=0 $Y2=0
cc_422 N_A_888_406#_c_550_n RESET_B 0.0277859f $X=6.655 $Y=1.705 $X2=0 $Y2=0
cc_423 N_A_888_406#_c_551_n RESET_B 0.056296f $X=7.725 $Y=1.545 $X2=0 $Y2=0
cc_424 N_A_888_406#_c_552_n RESET_B 0.0138646f $X=7.895 $Y=1.545 $X2=0 $Y2=0
cc_425 N_A_888_406#_c_553_n RESET_B 0.00110961f $X=8.985 $Y=1.465 $X2=0 $Y2=0
cc_426 N_A_888_406#_c_539_n N_RESET_B_c_843_n 0.0161669f $X=7.575 $Y=1.555 $X2=0
+ $Y2=0
cc_427 N_A_888_406#_c_547_n N_RESET_B_c_843_n 0.00126612f $X=5.75 $Y=0.81 $X2=0
+ $Y2=0
cc_428 N_A_888_406#_c_550_n N_RESET_B_c_843_n 0.00490094f $X=6.655 $Y=1.705
+ $X2=0 $Y2=0
cc_429 N_A_888_406#_c_561_n N_VPWR_M1010_d 0.00359259f $X=5.49 $Y=2.195 $X2=0
+ $Y2=0
cc_430 N_A_888_406#_c_565_n N_VPWR_c_896_n 0.0133787f $X=5.655 $Y=2.245 $X2=0
+ $Y2=0
cc_431 N_A_888_406#_c_548_n N_VPWR_c_897_n 0.0188408f $X=6.49 $Y=1.705 $X2=0
+ $Y2=0
cc_432 N_A_888_406#_c_564_n N_VPWR_c_897_n 0.0346006f $X=6.655 $Y=2.245 $X2=0
+ $Y2=0
cc_433 N_A_888_406#_c_565_n N_VPWR_c_897_n 0.0358549f $X=5.655 $Y=2.245 $X2=0
+ $Y2=0
cc_434 N_A_888_406#_M1019_g N_VPWR_c_898_n 0.00341102f $X=7.485 $Y=2.4 $X2=0
+ $Y2=0
cc_435 N_A_888_406#_c_564_n N_VPWR_c_898_n 0.0276905f $X=6.655 $Y=2.245 $X2=0
+ $Y2=0
cc_436 N_A_888_406#_c_551_n N_VPWR_c_898_n 0.0175657f $X=7.725 $Y=1.545 $X2=0
+ $Y2=0
cc_437 N_A_888_406#_M1023_g N_VPWR_c_899_n 0.00194999f $X=7.935 $Y=2.4 $X2=0
+ $Y2=0
cc_438 N_A_888_406#_M1025_g N_VPWR_c_899_n 0.012491f $X=8.435 $Y=2.4 $X2=0 $Y2=0
cc_439 N_A_888_406#_M1027_g N_VPWR_c_899_n 4.84307e-19 $X=8.985 $Y=2.4 $X2=0
+ $Y2=0
cc_440 N_A_888_406#_M1025_g N_VPWR_c_901_n 5.18084e-19 $X=8.435 $Y=2.4 $X2=0
+ $Y2=0
cc_441 N_A_888_406#_M1027_g N_VPWR_c_901_n 0.0178683f $X=8.985 $Y=2.4 $X2=0
+ $Y2=0
cc_442 N_A_888_406#_c_564_n N_VPWR_c_904_n 0.0135207f $X=6.655 $Y=2.245 $X2=0
+ $Y2=0
cc_443 N_A_888_406#_M1019_g N_VPWR_c_906_n 0.005209f $X=7.485 $Y=2.4 $X2=0 $Y2=0
cc_444 N_A_888_406#_M1023_g N_VPWR_c_906_n 0.005209f $X=7.935 $Y=2.4 $X2=0 $Y2=0
cc_445 N_A_888_406#_M1025_g N_VPWR_c_908_n 0.00460063f $X=8.435 $Y=2.4 $X2=0
+ $Y2=0
cc_446 N_A_888_406#_M1027_g N_VPWR_c_908_n 0.00460063f $X=8.985 $Y=2.4 $X2=0
+ $Y2=0
cc_447 N_A_888_406#_M1010_g N_VPWR_c_910_n 0.00562069f $X=4.53 $Y=2.73 $X2=0
+ $Y2=0
cc_448 N_A_888_406#_M1010_g N_VPWR_c_911_n 0.0206426f $X=4.53 $Y=2.73 $X2=0
+ $Y2=0
cc_449 N_A_888_406#_c_561_n N_VPWR_c_911_n 0.0399366f $X=5.49 $Y=2.195 $X2=0
+ $Y2=0
cc_450 N_A_888_406#_c_562_n N_VPWR_c_911_n 0.00316881f $X=4.605 $Y=2.195 $X2=0
+ $Y2=0
cc_451 N_A_888_406#_c_565_n N_VPWR_c_911_n 0.0132892f $X=5.655 $Y=2.245 $X2=0
+ $Y2=0
cc_452 N_A_888_406#_M1010_g N_VPWR_c_894_n 0.00539454f $X=4.53 $Y=2.73 $X2=0
+ $Y2=0
cc_453 N_A_888_406#_M1019_g N_VPWR_c_894_n 0.00986727f $X=7.485 $Y=2.4 $X2=0
+ $Y2=0
cc_454 N_A_888_406#_M1023_g N_VPWR_c_894_n 0.00982082f $X=7.935 $Y=2.4 $X2=0
+ $Y2=0
cc_455 N_A_888_406#_M1025_g N_VPWR_c_894_n 0.00909486f $X=8.435 $Y=2.4 $X2=0
+ $Y2=0
cc_456 N_A_888_406#_M1027_g N_VPWR_c_894_n 0.00909486f $X=8.985 $Y=2.4 $X2=0
+ $Y2=0
cc_457 N_A_888_406#_c_564_n N_VPWR_c_894_n 0.0119594f $X=6.655 $Y=2.245 $X2=0
+ $Y2=0
cc_458 N_A_888_406#_c_565_n N_VPWR_c_894_n 0.0119176f $X=5.655 $Y=2.245 $X2=0
+ $Y2=0
cc_459 N_A_888_406#_M1019_g N_Q_c_1016_n 0.00373184f $X=7.485 $Y=2.4 $X2=0 $Y2=0
cc_460 N_A_888_406#_c_538_n N_Q_c_1016_n 4.99328e-19 $X=7.74 $Y=1.555 $X2=0
+ $Y2=0
cc_461 N_A_888_406#_M1023_g N_Q_c_1016_n 8.84614e-19 $X=7.935 $Y=2.4 $X2=0 $Y2=0
cc_462 N_A_888_406#_c_551_n N_Q_c_1016_n 0.022627f $X=7.725 $Y=1.545 $X2=0 $Y2=0
cc_463 N_A_888_406#_M1019_g N_Q_c_1011_n 0.0101797f $X=7.485 $Y=2.4 $X2=0 $Y2=0
cc_464 N_A_888_406#_M1023_g N_Q_c_1011_n 0.0117052f $X=7.935 $Y=2.4 $X2=0 $Y2=0
cc_465 N_A_888_406#_M1025_g N_Q_c_1011_n 6.25418e-19 $X=8.435 $Y=2.4 $X2=0 $Y2=0
cc_466 N_A_888_406#_M1023_g N_Q_c_1023_n 0.0139523f $X=7.935 $Y=2.4 $X2=0 $Y2=0
cc_467 N_A_888_406#_M1025_g N_Q_c_1023_n 0.0156182f $X=8.435 $Y=2.4 $X2=0 $Y2=0
cc_468 N_A_888_406#_c_549_n N_Q_c_1023_n 0.0250657f $X=8.91 $Y=1.465 $X2=0 $Y2=0
cc_469 N_A_888_406#_c_552_n N_Q_c_1023_n 0.00144113f $X=7.895 $Y=1.545 $X2=0
+ $Y2=0
cc_470 N_A_888_406#_c_553_n N_Q_c_1023_n 0.00326676f $X=8.985 $Y=1.465 $X2=0
+ $Y2=0
cc_471 N_A_888_406#_M1001_g N_Q_c_1005_n 2.84024e-19 $X=7.815 $Y=0.74 $X2=0
+ $Y2=0
cc_472 N_A_888_406#_M1004_g N_Q_c_1005_n 2.84024e-19 $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_473 N_A_888_406#_M1001_g N_Q_c_1006_n 4.35498e-19 $X=7.815 $Y=0.74 $X2=0
+ $Y2=0
cc_474 N_A_888_406#_c_549_n N_Q_c_1006_n 0.0160251f $X=8.91 $Y=1.465 $X2=0 $Y2=0
cc_475 N_A_888_406#_c_553_n N_Q_c_1006_n 0.00272398f $X=8.985 $Y=1.465 $X2=0
+ $Y2=0
cc_476 N_A_888_406#_M1025_g N_Q_c_1012_n 4.86047e-19 $X=8.435 $Y=2.4 $X2=0 $Y2=0
cc_477 N_A_888_406#_M1027_g N_Q_c_1012_n 4.86047e-19 $X=8.985 $Y=2.4 $X2=0 $Y2=0
cc_478 N_A_888_406#_M1011_g N_Q_c_1007_n 2.84024e-19 $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_479 N_A_888_406#_M1022_g N_Q_c_1007_n 2.84024e-19 $X=9.105 $Y=0.74 $X2=0
+ $Y2=0
cc_480 N_A_888_406#_M1027_g N_Q_c_1013_n 0.0161477f $X=8.985 $Y=2.4 $X2=0 $Y2=0
cc_481 N_A_888_406#_c_549_n N_Q_c_1013_n 0.0143577f $X=8.91 $Y=1.465 $X2=0 $Y2=0
cc_482 N_A_888_406#_c_553_n N_Q_c_1013_n 0.00263964f $X=8.985 $Y=1.465 $X2=0
+ $Y2=0
cc_483 N_A_888_406#_M1025_g N_Q_c_1014_n 0.00116804f $X=8.435 $Y=2.4 $X2=0 $Y2=0
cc_484 N_A_888_406#_c_549_n N_Q_c_1014_n 0.0276641f $X=8.91 $Y=1.465 $X2=0 $Y2=0
cc_485 N_A_888_406#_c_553_n N_Q_c_1014_n 0.00517557f $X=8.985 $Y=1.465 $X2=0
+ $Y2=0
cc_486 N_A_888_406#_M1022_g Q 0.0178501f $X=9.105 $Y=0.74 $X2=0 $Y2=0
cc_487 N_A_888_406#_c_553_n Q 0.00267222f $X=8.985 $Y=1.465 $X2=0 $Y2=0
cc_488 N_A_888_406#_M1022_g Q 0.0112629f $X=9.105 $Y=0.74 $X2=0 $Y2=0
cc_489 N_A_888_406#_c_549_n Q 0.0267934f $X=8.91 $Y=1.465 $X2=0 $Y2=0
cc_490 N_A_888_406#_c_553_n Q 0.00743463f $X=8.985 $Y=1.465 $X2=0 $Y2=0
cc_491 N_A_888_406#_M1004_g N_Q_c_1010_n 0.0124418f $X=8.245 $Y=0.74 $X2=0 $Y2=0
cc_492 N_A_888_406#_M1011_g N_Q_c_1010_n 0.0124434f $X=8.675 $Y=0.74 $X2=0 $Y2=0
cc_493 N_A_888_406#_c_549_n N_Q_c_1010_n 0.071138f $X=8.91 $Y=1.465 $X2=0 $Y2=0
cc_494 N_A_888_406#_c_553_n N_Q_c_1010_n 0.00263605f $X=8.985 $Y=1.465 $X2=0
+ $Y2=0
cc_495 N_A_888_406#_M1015_g N_VGND_c_1080_n 0.011225f $X=4.545 $Y=0.58 $X2=0
+ $Y2=0
cc_496 N_A_888_406#_c_539_n N_VGND_c_1083_n 0.00338089f $X=7.575 $Y=1.555 $X2=0
+ $Y2=0
cc_497 N_A_888_406#_M1001_g N_VGND_c_1083_n 0.0116379f $X=7.815 $Y=0.74 $X2=0
+ $Y2=0
cc_498 N_A_888_406#_M1004_g N_VGND_c_1083_n 5.21765e-19 $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_499 N_A_888_406#_c_551_n N_VGND_c_1083_n 0.003848f $X=7.725 $Y=1.545 $X2=0
+ $Y2=0
cc_500 N_A_888_406#_c_552_n N_VGND_c_1083_n 0.00148206f $X=7.895 $Y=1.545 $X2=0
+ $Y2=0
cc_501 N_A_888_406#_M1001_g N_VGND_c_1084_n 4.765e-19 $X=7.815 $Y=0.74 $X2=0
+ $Y2=0
cc_502 N_A_888_406#_M1004_g N_VGND_c_1084_n 0.00952924f $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_503 N_A_888_406#_M1011_g N_VGND_c_1084_n 0.00952924f $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_504 N_A_888_406#_M1022_g N_VGND_c_1084_n 4.765e-19 $X=9.105 $Y=0.74 $X2=0
+ $Y2=0
cc_505 N_A_888_406#_M1011_g N_VGND_c_1086_n 4.31235e-19 $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_506 N_A_888_406#_M1022_g N_VGND_c_1086_n 0.00824245f $X=9.105 $Y=0.74 $X2=0
+ $Y2=0
cc_507 N_A_888_406#_M1015_g N_VGND_c_1087_n 0.00383152f $X=4.545 $Y=0.58 $X2=0
+ $Y2=0
cc_508 N_A_888_406#_M1001_g N_VGND_c_1091_n 0.00383152f $X=7.815 $Y=0.74 $X2=0
+ $Y2=0
cc_509 N_A_888_406#_M1004_g N_VGND_c_1091_n 0.00383152f $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_510 N_A_888_406#_M1011_g N_VGND_c_1092_n 0.00383152f $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_511 N_A_888_406#_M1022_g N_VGND_c_1092_n 0.00383152f $X=9.105 $Y=0.74 $X2=0
+ $Y2=0
cc_512 N_A_888_406#_M1015_g N_VGND_c_1099_n 0.00386109f $X=4.545 $Y=0.58 $X2=0
+ $Y2=0
cc_513 N_A_888_406#_M1001_g N_VGND_c_1099_n 0.0075754f $X=7.815 $Y=0.74 $X2=0
+ $Y2=0
cc_514 N_A_888_406#_M1004_g N_VGND_c_1099_n 0.0075754f $X=8.245 $Y=0.74 $X2=0
+ $Y2=0
cc_515 N_A_888_406#_M1011_g N_VGND_c_1099_n 0.0075754f $X=8.675 $Y=0.74 $X2=0
+ $Y2=0
cc_516 N_A_888_406#_M1022_g N_VGND_c_1099_n 0.00375577f $X=9.105 $Y=0.74 $X2=0
+ $Y2=0
cc_517 N_A_888_406#_M1015_g N_A_1035_74#_c_1198_n 0.00431882f $X=4.545 $Y=0.58
+ $X2=0 $Y2=0
cc_518 N_A_888_406#_M1009_s N_A_1035_74#_c_1199_n 0.00169477f $X=5.61 $Y=0.37
+ $X2=0 $Y2=0
cc_519 N_A_888_406#_c_547_n N_A_1035_74#_c_1199_n 0.0126348f $X=5.75 $Y=0.81
+ $X2=0 $Y2=0
cc_520 N_A_888_406#_M1015_g N_A_1035_74#_c_1200_n 6.04331e-19 $X=4.545 $Y=0.58
+ $X2=0 $Y2=0
cc_521 N_A_888_406#_c_548_n N_A_1035_74#_c_1207_n 0.00658578f $X=6.49 $Y=1.705
+ $X2=0 $Y2=0
cc_522 N_A_888_406#_M1001_g N_A_1035_74#_c_1202_n 7.13159e-19 $X=7.815 $Y=0.74
+ $X2=0 $Y2=0
cc_523 N_A_642_392#_M1016_g N_RESET_B_M1014_g 0.0179708f $X=5.88 $Y=2.52 $X2=0
+ $Y2=0
cc_524 N_A_642_392#_c_723_n N_RESET_B_c_839_n 0.00870882f $X=5.965 $Y=1.12 $X2=0
+ $Y2=0
cc_525 N_A_642_392#_c_728_n RESET_B 0.00162569f $X=5.88 $Y=1.455 $X2=0 $Y2=0
cc_526 N_A_642_392#_c_728_n N_RESET_B_c_843_n 0.0330602f $X=5.88 $Y=1.455 $X2=0
+ $Y2=0
cc_527 N_A_642_392#_M1012_g N_VPWR_c_896_n 0.00644749f $X=5.43 $Y=2.52 $X2=0
+ $Y2=0
cc_528 N_A_642_392#_M1016_g N_VPWR_c_896_n 0.00644749f $X=5.88 $Y=2.52 $X2=0
+ $Y2=0
cc_529 N_A_642_392#_M1016_g N_VPWR_c_897_n 0.00298275f $X=5.88 $Y=2.52 $X2=0
+ $Y2=0
cc_530 N_A_642_392#_M1012_g N_VPWR_c_911_n 0.00283737f $X=5.43 $Y=2.52 $X2=0
+ $Y2=0
cc_531 N_A_642_392#_M1012_g N_VPWR_c_894_n 0.00647345f $X=5.43 $Y=2.52 $X2=0
+ $Y2=0
cc_532 N_A_642_392#_M1016_g N_VPWR_c_894_n 0.00647345f $X=5.88 $Y=2.52 $X2=0
+ $Y2=0
cc_533 N_A_642_392#_c_722_n N_VGND_c_1080_n 0.00131584f $X=5.535 $Y=1.12 $X2=0
+ $Y2=0
cc_534 N_A_642_392#_c_765_n N_VGND_c_1080_n 0.00834935f $X=3.905 $Y=0.565 $X2=0
+ $Y2=0
cc_535 N_A_642_392#_c_724_n N_VGND_c_1080_n 0.0149311f $X=4.815 $Y=0.935 $X2=0
+ $Y2=0
cc_536 N_A_642_392#_c_726_n N_VGND_c_1080_n 0.00981709f $X=5.017 $Y=1.322 $X2=0
+ $Y2=0
cc_537 N_A_642_392#_c_723_n N_VGND_c_1081_n 2.42234e-19 $X=5.965 $Y=1.12 $X2=0
+ $Y2=0
cc_538 N_A_642_392#_c_765_n N_VGND_c_1087_n 0.0101443f $X=3.905 $Y=0.565 $X2=0
+ $Y2=0
cc_539 N_A_642_392#_c_722_n N_VGND_c_1090_n 0.00278247f $X=5.535 $Y=1.12 $X2=0
+ $Y2=0
cc_540 N_A_642_392#_c_723_n N_VGND_c_1090_n 0.00278247f $X=5.965 $Y=1.12 $X2=0
+ $Y2=0
cc_541 N_A_642_392#_c_722_n N_VGND_c_1099_n 0.00358425f $X=5.535 $Y=1.12 $X2=0
+ $Y2=0
cc_542 N_A_642_392#_c_723_n N_VGND_c_1099_n 0.00353524f $X=5.965 $Y=1.12 $X2=0
+ $Y2=0
cc_543 N_A_642_392#_c_765_n N_VGND_c_1099_n 0.0115712f $X=3.905 $Y=0.565 $X2=0
+ $Y2=0
cc_544 N_A_642_392#_c_724_n N_VGND_c_1099_n 0.0168958f $X=4.815 $Y=0.935 $X2=0
+ $Y2=0
cc_545 N_A_642_392#_c_726_n N_VGND_c_1099_n 0.00277523f $X=5.017 $Y=1.322 $X2=0
+ $Y2=0
cc_546 N_A_642_392#_c_722_n N_A_1035_74#_c_1198_n 0.00781452f $X=5.535 $Y=1.12
+ $X2=0 $Y2=0
cc_547 N_A_642_392#_c_723_n N_A_1035_74#_c_1198_n 6.05606e-19 $X=5.965 $Y=1.12
+ $X2=0 $Y2=0
cc_548 N_A_642_392#_c_726_n N_A_1035_74#_c_1198_n 0.0144827f $X=5.017 $Y=1.322
+ $X2=0 $Y2=0
cc_549 N_A_642_392#_c_728_n N_A_1035_74#_c_1198_n 0.0106502f $X=5.88 $Y=1.455
+ $X2=0 $Y2=0
cc_550 N_A_642_392#_c_722_n N_A_1035_74#_c_1199_n 0.0100245f $X=5.535 $Y=1.12
+ $X2=0 $Y2=0
cc_551 N_A_642_392#_c_723_n N_A_1035_74#_c_1199_n 0.0116238f $X=5.965 $Y=1.12
+ $X2=0 $Y2=0
cc_552 N_A_642_392#_c_728_n N_A_1035_74#_c_1199_n 2.49111e-19 $X=5.88 $Y=1.455
+ $X2=0 $Y2=0
cc_553 N_A_642_392#_c_722_n N_A_1035_74#_c_1200_n 0.00281658f $X=5.535 $Y=1.12
+ $X2=0 $Y2=0
cc_554 N_A_642_392#_c_723_n N_A_1035_74#_c_1207_n 0.00243926f $X=5.965 $Y=1.12
+ $X2=0 $Y2=0
cc_555 N_A_642_392#_c_722_n N_A_1035_74#_c_1218_n 5.52887e-19 $X=5.535 $Y=1.12
+ $X2=0 $Y2=0
cc_556 N_A_642_392#_c_723_n N_A_1035_74#_c_1218_n 0.00474692f $X=5.965 $Y=1.12
+ $X2=0 $Y2=0
cc_557 N_RESET_B_M1014_g N_VPWR_c_897_n 0.0168315f $X=6.38 $Y=2.52 $X2=0 $Y2=0
cc_558 N_RESET_B_M1029_g N_VPWR_c_897_n 7.97061e-19 $X=6.9 $Y=2.52 $X2=0 $Y2=0
cc_559 N_RESET_B_M1029_g N_VPWR_c_898_n 0.00863803f $X=6.9 $Y=2.52 $X2=0 $Y2=0
cc_560 N_RESET_B_M1014_g N_VPWR_c_904_n 0.00562069f $X=6.38 $Y=2.52 $X2=0 $Y2=0
cc_561 N_RESET_B_M1029_g N_VPWR_c_904_n 0.00666374f $X=6.9 $Y=2.52 $X2=0 $Y2=0
cc_562 N_RESET_B_M1014_g N_VPWR_c_894_n 0.0054305f $X=6.38 $Y=2.52 $X2=0 $Y2=0
cc_563 N_RESET_B_M1029_g N_VPWR_c_894_n 0.00647345f $X=6.9 $Y=2.52 $X2=0 $Y2=0
cc_564 N_RESET_B_M1029_g N_Q_c_1016_n 5.4687e-19 $X=6.9 $Y=2.52 $X2=0 $Y2=0
cc_565 RESET_B N_Q_c_1006_n 4.79428e-19 $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_566 N_RESET_B_c_839_n N_VGND_c_1081_n 0.00623004f $X=6.395 $Y=1.12 $X2=0
+ $Y2=0
cc_567 N_RESET_B_c_840_n N_VGND_c_1081_n 0.00749966f $X=6.825 $Y=1.12 $X2=0
+ $Y2=0
cc_568 N_RESET_B_c_840_n N_VGND_c_1082_n 0.00383152f $X=6.825 $Y=1.12 $X2=0
+ $Y2=0
cc_569 N_RESET_B_c_840_n N_VGND_c_1083_n 0.00252276f $X=6.825 $Y=1.12 $X2=0
+ $Y2=0
cc_570 RESET_B N_VGND_c_1083_n 0.0103498f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_571 N_RESET_B_c_839_n N_VGND_c_1090_n 0.00383152f $X=6.395 $Y=1.12 $X2=0
+ $Y2=0
cc_572 N_RESET_B_c_839_n N_VGND_c_1099_n 0.00369368f $X=6.395 $Y=1.12 $X2=0
+ $Y2=0
cc_573 N_RESET_B_c_840_n N_VGND_c_1099_n 0.00374269f $X=6.825 $Y=1.12 $X2=0
+ $Y2=0
cc_574 N_RESET_B_c_839_n N_A_1035_74#_c_1199_n 9.48753e-19 $X=6.395 $Y=1.12
+ $X2=0 $Y2=0
cc_575 N_RESET_B_c_839_n N_A_1035_74#_c_1221_n 0.00969758f $X=6.395 $Y=1.12
+ $X2=0 $Y2=0
cc_576 N_RESET_B_c_840_n N_A_1035_74#_c_1221_n 0.00969758f $X=6.825 $Y=1.12
+ $X2=0 $Y2=0
cc_577 RESET_B N_A_1035_74#_c_1221_n 0.0397203f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_578 N_RESET_B_c_843_n N_A_1035_74#_c_1221_n 0.0024149f $X=6.825 $Y=1.285
+ $X2=0 $Y2=0
cc_579 RESET_B N_A_1035_74#_c_1201_n 0.0216332f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_580 N_RESET_B_c_843_n N_A_1035_74#_c_1201_n 0.00118495f $X=6.825 $Y=1.285
+ $X2=0 $Y2=0
cc_581 N_RESET_B_c_840_n N_A_1035_74#_c_1202_n 3.34329e-19 $X=6.825 $Y=1.12
+ $X2=0 $Y2=0
cc_582 N_VPWR_c_898_n N_Q_c_1011_n 0.032647f $X=7.21 $Y=2.245 $X2=0 $Y2=0
cc_583 N_VPWR_c_899_n N_Q_c_1011_n 0.0263057f $X=8.21 $Y=2.465 $X2=0 $Y2=0
cc_584 N_VPWR_c_906_n N_Q_c_1011_n 0.0144623f $X=8.045 $Y=3.33 $X2=0 $Y2=0
cc_585 N_VPWR_c_894_n N_Q_c_1011_n 0.0118344f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_586 N_VPWR_M1023_d N_Q_c_1023_n 0.00479311f $X=8.025 $Y=1.84 $X2=0 $Y2=0
cc_587 N_VPWR_c_899_n N_Q_c_1023_n 0.0189268f $X=8.21 $Y=2.465 $X2=0 $Y2=0
cc_588 N_VPWR_c_899_n N_Q_c_1012_n 0.0263057f $X=8.21 $Y=2.465 $X2=0 $Y2=0
cc_589 N_VPWR_c_901_n N_Q_c_1012_n 0.0323093f $X=9.21 $Y=2.305 $X2=0 $Y2=0
cc_590 N_VPWR_c_908_n N_Q_c_1012_n 0.0146357f $X=9.045 $Y=3.33 $X2=0 $Y2=0
cc_591 N_VPWR_c_894_n N_Q_c_1012_n 0.0121141f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_592 N_VPWR_M1027_d N_Q_c_1013_n 0.00312742f $X=9.075 $Y=1.84 $X2=0 $Y2=0
cc_593 N_VPWR_c_901_n N_Q_c_1013_n 0.023022f $X=9.21 $Y=2.305 $X2=0 $Y2=0
cc_594 N_Q_c_1010_n N_VGND_M1004_d 0.00176461f $X=8.795 $Y=0.965 $X2=0 $Y2=0
cc_595 Q N_VGND_M1022_d 0.0042279f $X=9.275 $Y=0.84 $X2=0 $Y2=0
cc_596 N_Q_c_1005_n N_VGND_c_1083_n 0.0224826f $X=8.03 $Y=0.525 $X2=0 $Y2=0
cc_597 N_Q_c_1005_n N_VGND_c_1084_n 0.016479f $X=8.03 $Y=0.525 $X2=0 $Y2=0
cc_598 N_Q_c_1007_n N_VGND_c_1084_n 0.016479f $X=8.89 $Y=0.525 $X2=0 $Y2=0
cc_599 N_Q_c_1010_n N_VGND_c_1084_n 0.0170777f $X=8.795 $Y=0.965 $X2=0 $Y2=0
cc_600 N_Q_c_1007_n N_VGND_c_1086_n 0.0104754f $X=8.89 $Y=0.525 $X2=0 $Y2=0
cc_601 Q N_VGND_c_1086_n 0.0216656f $X=9.275 $Y=0.84 $X2=0 $Y2=0
cc_602 N_Q_c_1005_n N_VGND_c_1091_n 0.00806491f $X=8.03 $Y=0.525 $X2=0 $Y2=0
cc_603 N_Q_c_1007_n N_VGND_c_1092_n 0.00781705f $X=8.89 $Y=0.525 $X2=0 $Y2=0
cc_604 N_Q_c_1005_n N_VGND_c_1099_n 0.00690154f $X=8.03 $Y=0.525 $X2=0 $Y2=0
cc_605 N_Q_c_1007_n N_VGND_c_1099_n 0.00680101f $X=8.89 $Y=0.525 $X2=0 $Y2=0
cc_606 Q N_VGND_c_1099_n 0.00669281f $X=9.275 $Y=0.84 $X2=0 $Y2=0
cc_607 N_VGND_c_1080_n N_A_1035_74#_c_1198_n 0.017158f $X=4.76 $Y=0.515 $X2=0
+ $Y2=0
cc_608 N_VGND_c_1081_n N_A_1035_74#_c_1199_n 0.0112234f $X=6.61 $Y=0.515 $X2=0
+ $Y2=0
cc_609 N_VGND_c_1090_n N_A_1035_74#_c_1199_n 0.0512248f $X=6.445 $Y=0 $X2=0
+ $Y2=0
cc_610 N_VGND_c_1099_n N_A_1035_74#_c_1199_n 0.0283929f $X=9.36 $Y=0 $X2=0 $Y2=0
cc_611 N_VGND_c_1080_n N_A_1035_74#_c_1200_n 0.0121616f $X=4.76 $Y=0.515 $X2=0
+ $Y2=0
cc_612 N_VGND_c_1090_n N_A_1035_74#_c_1200_n 0.0236075f $X=6.445 $Y=0 $X2=0
+ $Y2=0
cc_613 N_VGND_c_1099_n N_A_1035_74#_c_1200_n 0.0127226f $X=9.36 $Y=0 $X2=0 $Y2=0
cc_614 N_VGND_M1002_s N_A_1035_74#_c_1221_n 0.0032758f $X=6.47 $Y=0.37 $X2=0
+ $Y2=0
cc_615 N_VGND_c_1081_n N_A_1035_74#_c_1221_n 0.0166614f $X=6.61 $Y=0.515 $X2=0
+ $Y2=0
cc_616 N_VGND_c_1099_n N_A_1035_74#_c_1221_n 0.0122318f $X=9.36 $Y=0 $X2=0 $Y2=0
cc_617 N_VGND_c_1083_n N_A_1035_74#_c_1201_n 0.012877f $X=7.6 $Y=0.525 $X2=0
+ $Y2=0
cc_618 N_VGND_c_1081_n N_A_1035_74#_c_1202_n 0.00975481f $X=6.61 $Y=0.515 $X2=0
+ $Y2=0
cc_619 N_VGND_c_1082_n N_A_1035_74#_c_1202_n 0.0111768f $X=7.435 $Y=0 $X2=0
+ $Y2=0
cc_620 N_VGND_c_1083_n N_A_1035_74#_c_1202_n 0.0274502f $X=7.6 $Y=0.525 $X2=0
+ $Y2=0
cc_621 N_VGND_c_1099_n N_A_1035_74#_c_1202_n 0.00945682f $X=9.36 $Y=0 $X2=0
+ $Y2=0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfbbn_2 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR
+ Q Q_N
X0 VPWR a_1007_366# a_1989_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X1 a_1989_424# a_871_368# a_1997_82# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X2 VPWR a_2216_410# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 a_1007_366# a_1157_464# a_1595_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X4 a_1157_464# a_871_368# a_197_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X5 Q a_3272_94# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_688_98# CLK_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 a_1997_82# a_688_98# a_2174_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X8 a_1643_257# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X9 a_1473_73# a_1157_464# a_1007_366# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X10 a_1997_82# a_871_368# a_2247_82# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X11 a_209_464# D a_197_119# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X12 a_1473_73# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X13 a_2174_508# a_2216_410# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X14 a_3272_94# a_2216_410# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X15 a_27_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X16 VGND SCE a_341_410# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X17 VGND a_688_98# a_871_368# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 VGND SET_B a_2452_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 VPWR a_3272_94# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X20 a_1007_366# a_1643_257# a_1473_73# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X21 VGND SCD a_119_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X22 a_363_119# a_341_410# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X23 VGND a_1007_366# a_1185_125# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X24 a_1185_125# a_688_98# a_1157_464# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X25 VGND a_1007_366# a_1902_125# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X26 a_1157_464# a_688_98# a_197_119# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X27 VPWR a_1643_257# a_2559_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X28 Q_N a_2216_410# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X29 VPWR a_688_98# a_871_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X30 Q_N a_2216_410# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X31 a_1073_464# a_871_368# a_1157_464# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X32 a_1902_125# a_688_98# a_1997_82# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X33 a_2452_74# a_1643_257# a_2216_410# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X34 a_2559_392# a_1997_82# a_2216_410# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X35 a_1595_424# a_1643_257# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X36 a_688_98# CLK_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X37 a_2216_410# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X38 a_3272_94# a_2216_410# VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X39 VGND a_2216_410# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X40 a_197_119# a_341_410# a_27_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X41 VPWR SCE a_341_410# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X42 VGND a_3272_94# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X43 a_2247_82# a_2216_410# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X44 a_1643_257# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X45 a_2216_410# a_1997_82# a_2452_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X46 a_197_119# D a_363_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X47 Q a_3272_94# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X48 VPWR SCE a_209_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X49 VPWR a_1007_366# a_1073_464# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X50 VPWR SET_B a_1007_366# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X51 a_119_119# SCE a_197_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
.ends

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfrbp_2 CLK D RESET_B VGND VNB VPB VPWR Q Q_N
M1000 Q a_2366_352# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=3.6099e+12p ps=2.652e+07u
M1001 Q a_2366_352# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=2.19475e+12p ps=1.777e+07u
M1002 a_1800_291# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1003 VPWR a_2366_352# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR RESET_B a_70_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=3.864e+11p ps=3.52e+06u
M1005 a_1758_389# a_818_418# a_1586_149# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=3.55e+11p ps=3e+06u
M1006 a_298_294# a_728_331# a_70_74# VNB nlowvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=2.632e+11p ps=3.03e+06u
M1007 a_728_331# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1008 VGND a_1800_291# a_1499_149# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.8e+06u
M1009 a_728_331# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1010 VGND a_1586_149# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.072e+11p ps=2.04e+06u
M1011 VPWR RESET_B a_298_294# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=2.247e+11p ps=2.75e+06u
M1012 a_156_74# D a_70_74# VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1013 a_686_485# a_334_119# VPWR VPB pshort w=420000u l=180000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1014 VPWR a_1800_291# a_1758_389# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_614_81# a_334_119# a_536_81# VNB nlowvt w=420000u l=150000u
+  ad=3.465e+11p pd=3.33e+06u as=1.008e+11p ps=1.32e+06u
M1016 VGND a_2366_352# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1586_149# a_728_331# a_1499_149# VNB nlowvt w=420000u l=150000u
+  ad=2.165e+11p pd=2.13e+06u as=0p ps=0u
M1018 a_1800_291# a_1586_149# a_1974_74# VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1019 VPWR a_1586_149# a_1800_291# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_2366_352# a_1586_149# VPWR VPB pshort w=1e+06u l=180000u
+  ad=3.75e+11p pd=2.75e+06u as=0p ps=0u
M1021 a_1974_74# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_2366_352# a_1586_149# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1023 a_334_119# a_298_294# VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.45e+11p pd=5.09e+06u as=0p ps=0u
M1024 a_298_294# a_728_331# a_686_485# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_334_119# a_818_418# a_1586_149# VNB nlowvt w=740000u l=150000u
+  ad=5.2345e+11p pd=4.67e+06u as=0p ps=0u
M1026 a_70_74# a_818_418# a_298_294# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1586_149# a_728_331# a_334_119# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_536_81# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND a_728_331# a_818_418# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.998e+11p ps=2.02e+06u
M1030 Q_N a_1586_149# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1031 a_334_119# a_298_294# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_614_81# a_818_418# a_298_294# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Q_N a_1586_149# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR a_728_331# a_818_418# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1035 VPWR a_1586_149# Q_N VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_70_74# D VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND RESET_B a_156_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

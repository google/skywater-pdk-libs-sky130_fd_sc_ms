* File: sky130_fd_sc_ms__nor4_4.spice
* Created: Fri Aug 28 17:49:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nor4_4.pex.spice"
.subckt sky130_fd_sc_ms__nor4_4  VNB VPB D C B A Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_D_M1001_g N_Y_M1001_s VNB NLOWVT L=0.15 W=0.74 AD=0.2442
+ AS=0.4329 PD=2.14 PS=1.91 NRD=7.296 NRS=0 M=1 R=4.93333 SA=75000.3 SB=75007.6
+ A=0.111 P=1.78 MULT=1
MM1022 N_VGND_M1022_d N_D_M1022_g N_Y_M1001_s VNB NLOWVT L=0.15 W=0.74 AD=0.1295
+ AS=0.4329 PD=1.09 PS=1.91 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6 SB=75006.3
+ A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1022_d N_C_M1014_g N_Y_M1014_s VNB NLOWVT L=0.15 W=0.74 AD=0.1295
+ AS=0.444 PD=1.09 PS=1.94 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.1 SB=75005.8
+ A=0.111 P=1.78 MULT=1
MM1023 N_VGND_M1023_d N_C_M1023_g N_Y_M1014_s VNB NLOWVT L=0.15 W=0.74 AD=0.1295
+ AS=0.444 PD=1.09 PS=1.94 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.4 SB=75004.5
+ A=0.111 P=1.78 MULT=1
MM1009 N_Y_M1009_d N_B_M1009_g N_VGND_M1023_d VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003.9 SB=75004
+ A=0.111 P=1.78 MULT=1
MM1020 N_Y_M1009_d N_B_M1020_g N_VGND_M1020_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.8621 PD=1.02 PS=3.07 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.4 SB=75003.5
+ A=0.111 P=1.78 MULT=1
MM1016 N_Y_M1016_d N_A_M1016_g N_VGND_M1020_s VNB NLOWVT L=0.15 W=0.74 AD=0.2627
+ AS=0.8621 PD=1.45 PS=3.07 NRD=48.648 NRS=0 M=1 R=4.93333 SA=75006.8 SB=75001.1
+ A=0.111 P=1.78 MULT=1
MM1021 N_Y_M1016_d N_A_M1021_g N_VGND_M1021_s VNB NLOWVT L=0.15 W=0.74 AD=0.2627
+ AS=0.2109 PD=1.45 PS=2.05 NRD=48.648 NRS=0 M=1 R=4.93333 SA=75007.7 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_D_M1002_g N_A_27_368#_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.2
+ SB=90003.4 A=0.2016 P=2.6 MULT=1
MM1003 N_Y_M1002_d N_D_M1003_g N_A_27_368#_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.7
+ SB=90002.9 A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1004_d N_D_M1004_g N_A_27_368#_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90002.5 A=0.2016 P=2.6 MULT=1
MM1006 N_Y_M1004_d N_D_M1006_g N_A_27_368#_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.6
+ SB=90002 A=0.2016 P=2.6 MULT=1
MM1007 N_A_499_368#_M1007_d N_C_M1007_g N_A_27_368#_M1006_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90002.1 SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1012 N_A_499_368#_M1007_d N_C_M1012_g N_A_27_368#_M1012_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90002.5 SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1015 N_A_499_368#_M1015_d N_C_M1015_g N_A_27_368#_M1012_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1017 N_A_499_368#_M1015_d N_C_M1017_g N_A_27_368#_M1017_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.4
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1000 N_A_499_368#_M1000_d N_B_M1000_g N_A_879_368#_M1000_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003.6 A=0.2016 P=2.6 MULT=1
MM1005 N_A_499_368#_M1000_d N_B_M1005_g N_A_879_368#_M1005_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1624 PD=1.39 PS=1.41 NRD=0 NRS=0.8668 M=1 R=6.22222
+ SA=90000.6 SB=90003.1 A=0.2016 P=2.6 MULT=1
MM1010 N_A_499_368#_M1010_d N_B_M1010_g N_A_879_368#_M1005_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1624 PD=1.39 PS=1.41 NRD=0 NRS=0.8668 M=1 R=6.22222
+ SA=90001.1 SB=90002.6 A=0.2016 P=2.6 MULT=1
MM1013 N_A_499_368#_M1010_d N_B_M1013_g N_A_879_368#_M1013_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.6 SB=90002.2 A=0.2016 P=2.6 MULT=1
MM1008 N_A_879_368#_M1013_s N_A_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002
+ SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1011 N_A_879_368#_M1011_d N_A_M1011_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.6
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1018 N_A_879_368#_M1011_d N_A_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1019 N_A_879_368#_M1019_d N_A_M1019_g N_VPWR_M1018_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.2072 PD=2.8 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX24_noxref VNB VPB NWDIODE A=16.7772 P=21.76
*
.include "sky130_fd_sc_ms__nor4_4.pxi.spice"
*
.ends
*
*

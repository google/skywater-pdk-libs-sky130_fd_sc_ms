* NGSPICE file created from sky130_fd_sc_ms__and4_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__and4_1 A B C D VGND VNB VPB VPWR X
M1000 VPWR B a_96_74# VPB pshort w=840000u l=180000u
+  ad=1.1326e+12p pd=8.13e+06u as=5.376e+11p ps=4.64e+06u
M1001 VPWR D a_96_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1002 a_96_74# C VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND D a_335_74# VNB nlowvt w=640000u l=150000u
+  ad=2.554e+11p pd=2.2e+06u as=2.688e+11p ps=2.12e+06u
M1004 a_96_74# A VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_96_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1006 X a_96_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1007 a_257_74# B a_179_74# VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.536e+11p ps=1.76e+06u
M1008 a_335_74# C a_257_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_179_74# A a_96_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
.ends


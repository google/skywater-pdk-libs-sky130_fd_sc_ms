* File: sky130_fd_sc_ms__a31oi_1.spice
* Created: Wed Sep  2 11:55:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a31oi_1.pex.spice"
.subckt sky130_fd_sc_ms__a31oi_1  VNB VPB A3 A2 A1 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1006 A_145_74# N_A3_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.3182 PD=0.98 PS=2.34 NRD=10.536 NRS=23.508 M=1 R=4.93333 SA=75000.4
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1004 A_223_74# N_A2_M1004_g A_145_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.0888 PD=1.16 PS=0.98 NRD=25.128 NRS=10.536 M=1 R=4.93333 SA=75000.7
+ SB=75001.4 A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1003_d N_A1_M1003_g A_223_74# VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.1554 PD=1.16 PS=1.16 NRD=11.34 NRS=25.128 M=1 R=4.93333 SA=75001.3
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_B1_M1005_g N_Y_M1003_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.9
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_A_139_368#_M1007_d N_A3_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.4144 PD=1.39 PS=2.98 NRD=0 NRS=14.9326 M=1 R=6.22222 SA=90000.3
+ SB=90001.8 A=0.2016 P=2.6 MULT=1
MM1000 N_VPWR_M1000_d N_A2_M1000_g N_A_139_368#_M1007_d VPB PSHORT L=0.18 W=1.12
+ AD=0.2576 AS=0.1512 PD=1.58 PS=1.39 NRD=14.9326 NRS=0 M=1 R=6.22222 SA=90000.7
+ SB=90001.3 A=0.2016 P=2.6 MULT=1
MM1001 N_A_139_368#_M1001_d N_A1_M1001_g N_VPWR_M1000_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.2576 PD=1.44 PS=1.58 NRD=0 NRS=16.7056 M=1 R=6.22222 SA=90001.4
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1002 N_Y_M1002_d N_B1_M1002_g N_A_139_368#_M1001_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1792 PD=2.8 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.9
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0636 P=10.24
*
.include "sky130_fd_sc_ms__a31oi_1.pxi.spice"
*
.ends
*
*

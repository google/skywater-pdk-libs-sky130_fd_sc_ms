* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfbbn_1 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR
+ Q Q_N
X0 a_2091_508# a_2133_410# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X1 a_197_119# a_353_93# a_27_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X2 a_1162_497# a_867_82# a_197_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 a_977_243# a_1579_258# a_1434_78# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X4 a_2133_410# a_1954_119# a_2392_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_1579_258# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X6 a_1151_119# a_662_82# a_1162_497# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X7 VPWR a_662_82# a_867_82# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 VPWR a_977_243# a_1084_497# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X9 VPWR a_1579_258# a_2512_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X10 VPWR a_3078_384# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X11 VGND a_3078_384# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X12 a_1434_78# a_1162_497# a_977_243# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X13 a_977_243# a_1162_497# a_1531_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X14 VPWR SCE a_353_93# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X15 a_3078_384# a_2133_410# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X16 a_2133_410# SET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X17 a_1579_258# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X18 a_27_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X19 VGND a_2133_410# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 a_1084_497# a_867_82# a_1162_497# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X21 a_1531_424# a_1579_258# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X22 a_1906_424# a_867_82# a_1954_119# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X23 a_305_119# a_353_93# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X24 a_662_82# CLK_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 a_215_464# D a_197_119# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X26 VGND SCD a_119_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X27 VGND SCE a_353_93# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X28 a_2164_119# a_2133_410# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X29 a_1876_119# a_662_82# a_1954_119# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X30 a_662_82# CLK_N VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X31 VGND a_977_243# a_1151_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X32 VGND a_662_82# a_867_82# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X33 a_1954_119# a_867_82# a_2164_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X34 a_3078_384# a_2133_410# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X35 VPWR a_977_243# a_1906_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X36 a_2392_74# a_1579_258# a_2133_410# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X37 a_1954_119# a_662_82# a_2091_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X38 a_2512_392# a_1954_119# a_2133_410# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X39 VGND SET_B a_2392_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X40 VPWR SCE a_215_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X41 a_1434_78# SET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X42 a_197_119# D a_305_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X43 VPWR SET_B a_977_243# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X44 VPWR a_2133_410# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X45 a_1162_497# a_662_82# a_197_119# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X46 VGND a_977_243# a_1876_119# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X47 a_119_119# SCE a_197_119# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
.ends

* File: sky130_fd_sc_ms__fahcon_1.spice
* Created: Fri Aug 28 17:36:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__fahcon_1.pex.spice"
.subckt sky130_fd_sc_ms__fahcon_1  VNB VPB A B CI VPWR COUT_N SUM VGND
* 
* VGND	VGND
* SUM	SUM
* COUT_N	COUT_N
* VPWR	VPWR
* CI	CI
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1014 N_VGND_M1014_d N_A_M1014_g N_A_27_100#_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.263987 AS=0.2109 PD=1.5658 PS=2.05 NRD=2.424 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.6 A=0.111 P=1.78 MULT=1
MM1002 N_A_244_368#_M1002_d N_A_27_100#_M1002_g N_VGND_M1014_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.228313 PD=0.92 PS=1.3542 NRD=0 NRS=80.616 M=1 R=4.26667
+ SA=75001.1 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1003 N_A_374_120#_M1003_d N_A_336_263#_M1003_g N_A_244_368#_M1002_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.150225 AS=0.0896 PD=1.145 PS=0.92 NRD=14.988 NRS=0 M=1
+ R=4.26667 SA=75001.5 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1013 N_A_27_100#_M1013_d N_B_M1013_g N_A_374_120#_M1003_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.0928 AS=0.150225 PD=0.93 PS=1.145 NRD=1.872 NRS=14.988 M=1
+ R=4.26667 SA=75001.9 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1030 N_A_372_365#_M1030_d N_A_336_263#_M1030_g N_A_27_100#_M1013_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1456 AS=0.0928 PD=1.095 PS=0.93 NRD=13.116 NRS=0 M=1
+ R=4.26667 SA=75002.4 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1015 N_A_244_368#_M1015_d N_B_M1015_g N_A_372_365#_M1030_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.1456 PD=1.85 PS=1.095 NRD=0 NRS=19.68 M=1 R=4.26667
+ SA=75003 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1024 N_VGND_M1024_d N_B_M1024_g N_A_336_263#_M1024_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.124942 AS=0.4662 PD=1.14217 PS=2.74 NRD=7.296 NRS=2.016 M=1 R=4.93333
+ SA=75000.6 SB=75005.2 A=0.111 P=1.78 MULT=1
MM1031 N_A_1026_389#_M1031_d N_B_M1031_g N_VGND_M1024_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.2496 AS=0.108058 PD=1.42 PS=0.987826 NRD=0 NRS=0 M=1 R=4.26667 SA=75001
+ SB=75005.5 A=0.096 P=1.58 MULT=1
MM1016 N_COUT_N_M1016_d N_A_372_365#_M1016_g N_A_1026_389#_M1031_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1792 AS=0.2496 PD=1.2 PS=1.42 NRD=10.308 NRS=2.808 M=1
+ R=4.26667 SA=75002 SB=75004.6 A=0.096 P=1.58 MULT=1
MM1018 N_A_1264_421#_M1018_d N_A_374_120#_M1018_g N_COUT_N_M1016_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.176 AS=0.1792 PD=1.19 PS=1.2 NRD=50.616 NRS=42.18 M=1
+ R=4.26667 SA=75002.7 SB=75003.9 A=0.096 P=1.58 MULT=1
MM1025 N_VGND_M1025_d N_CI_M1025_g N_A_1264_421#_M1018_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.118446 AS=0.176 PD=1.02029 PS=1.19 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75003.4 SB=75003.2 A=0.096 P=1.58 MULT=1
MM1004 N_A_1609_368#_M1004_d N_CI_M1004_g N_VGND_M1025_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.13883 AS=0.136954 PD=1.17971 PS=1.17971 NRD=0 NRS=1.62 M=1
+ R=4.93333 SA=75003.4 SB=75002.7 A=0.111 P=1.78 MULT=1
MM1026 N_A_1744_94#_M1026_d N_A_372_365#_M1026_g N_A_1609_368#_M1004_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.2112 AS=0.12007 PD=1.3 PS=1.02029 NRD=14.988
+ NRS=15.468 M=1 R=4.26667 SA=75003.8 SB=75002.6 A=0.096 P=1.58 MULT=1
MM1022 N_A_1719_368#_M1022_d N_A_374_120#_M1022_g N_A_1744_94#_M1026_d VNB
+ NLOWVT L=0.15 W=0.64 AD=0.1632 AS=0.2112 PD=1.15 PS=1.3 NRD=43.116 NRS=56.244
+ M=1 R=4.26667 SA=75004.6 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1017 N_VGND_M1017_d N_A_1609_368#_M1017_g N_A_1719_368#_M1022_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.277472 AS=0.1632 PD=1.56754 PS=1.15 NRD=70.968 NRS=0 M=1
+ R=4.26667 SA=75005.3 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1009 N_SUM_M1009_d N_A_1744_94#_M1009_g N_VGND_M1017_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.320828 PD=2.05 PS=1.81246 NRD=0 NRS=61.38 M=1 R=4.93333
+ SA=75005.4 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1020 N_VPWR_M1020_d N_A_M1020_g N_A_27_100#_M1020_s VPB PSHORT L=0.18 W=1.12
+ AD=0.234883 AS=0.3136 PD=1.61132 PS=2.8 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1021 N_A_244_368#_M1021_d N_A_27_100#_M1021_g N_VPWR_M1020_d VPB PSHORT L=0.18
+ W=1 AD=0.234918 AS=0.209717 PD=1.60326 PS=1.43868 NRD=0 NRS=16.0752 M=1
+ R=5.55556 SA=90000.8 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1000 N_A_372_365#_M1000_d N_A_336_263#_M1000_g N_A_244_368#_M1021_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.1638 AS=0.197332 PD=1.23 PS=1.34674 NRD=26.9693 NRS=43.7734
+ M=1 R=4.66667 SA=90001.4 SB=90001.8 A=0.1512 P=2.04 MULT=1
MM1008 N_A_27_100#_M1008_d N_B_M1008_g N_A_372_365#_M1000_d VPB PSHORT L=0.18
+ W=0.84 AD=0.1134 AS=0.1638 PD=1.11 PS=1.23 NRD=0 NRS=0 M=1 R=4.66667 SA=90002
+ SB=90001.2 A=0.1512 P=2.04 MULT=1
MM1011 N_A_374_120#_M1011_d N_A_336_263#_M1011_g N_A_27_100#_M1008_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.1988 AS=0.1134 PD=1.4 PS=1.11 NRD=18.7544 NRS=0 M=1
+ R=4.66667 SA=90002.4 SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1019 N_A_244_368#_M1019_d N_B_M1019_g N_A_374_120#_M1011_d VPB PSHORT L=0.18
+ W=0.84 AD=0.231 AS=0.1988 PD=2.23 PS=1.4 NRD=0 NRS=18.7544 M=1 R=4.66667
+ SA=90003 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1027 N_VPWR_M1027_d N_B_M1027_g N_A_336_263#_M1027_s VPB PSHORT L=0.18 W=1.12
+ AD=0.245449 AS=0.3136 PD=1.63245 PS=2.8 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90002.9 A=0.2016 P=2.6 MULT=1
MM1001 N_A_1026_389#_M1001_d N_B_M1001_g N_VPWR_M1027_d VPB PSHORT L=0.18 W=1
+ AD=0.186413 AS=0.219151 PD=1.47283 PS=1.45755 NRD=0 NRS=20.0152 M=1 R=5.55556
+ SA=90000.8 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1012 N_COUT_N_M1012_d N_A_374_120#_M1012_g N_A_1026_389#_M1001_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.1995 AS=0.156587 PD=1.315 PS=1.23717 NRD=35.1645
+ NRS=19.1484 M=1 R=4.66667 SA=90001.3 SB=90002.6 A=0.1512 P=2.04 MULT=1
MM1023 N_A_1264_421#_M1023_d N_A_372_365#_M1023_g N_COUT_N_M1012_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.417078 AS=0.1995 PD=1.86261 PS=1.315 NRD=0 NRS=10.5395 M=1
+ R=4.66667 SA=90002 SB=90001.9 A=0.1512 P=2.04 MULT=1
MM1005 N_VPWR_M1005_d N_CI_M1005_g N_A_1264_421#_M1023_d VPB PSHORT L=0.18 W=1
+ AD=0.167453 AS=0.496522 PD=1.36321 PS=2.21739 NRD=9.8303 NRS=0 M=1 R=5.55556
+ SA=90002.7 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1006 N_A_1609_368#_M1006_d N_CI_M1006_g N_VPWR_M1005_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.187547 PD=2.8 PS=1.52679 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90002.9 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1007 N_A_1744_94#_M1007_d N_A_372_365#_M1007_g N_A_1719_368#_M1007_s VPB
+ PSHORT L=0.18 W=0.84 AD=0.1134 AS=0.3907 PD=1.11 PS=2.99 NRD=0 NRS=96.1754 M=1
+ R=4.66667 SA=90000.3 SB=90000.6 A=0.1512 P=2.04 MULT=1
MM1010 N_A_1609_368#_M1010_d N_A_374_120#_M1010_g N_A_1744_94#_M1007_d VPB
+ PSHORT L=0.18 W=0.84 AD=0.2352 AS=0.1134 PD=2.24 PS=1.11 NRD=0 NRS=0 M=1
+ R=4.66667 SA=90000.7 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1028 N_VPWR_M1028_d N_A_1609_368#_M1028_g N_A_1719_368#_M1028_s VPB PSHORT
+ L=0.18 W=1 AD=0.167453 AS=0.28 PD=1.36321 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1029 N_SUM_M1029_d N_A_1744_94#_M1029_g N_VPWR_M1028_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.187547 PD=2.8 PS=1.52679 NRD=0 NRS=8.7862 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX32_noxref VNB VPB NWDIODE A=22.1908 P=27.55
c_221 VPB 0 2.78883e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__fahcon_1.pxi.spice"
*
.ends
*
*

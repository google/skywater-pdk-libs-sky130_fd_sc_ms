* File: sky130_fd_sc_ms__o21bai_1.pxi.spice
* Created: Fri Aug 28 17:56:05 2020
* 
x_PM_SKY130_FD_SC_MS__O21BAI_1%B1_N N_B1_N_M1001_g N_B1_N_c_61_n N_B1_N_M1005_g
+ B1_N N_B1_N_c_62_n PM_SKY130_FD_SC_MS__O21BAI_1%B1_N
x_PM_SKY130_FD_SC_MS__O21BAI_1%A_27_74# N_A_27_74#_M1001_s N_A_27_74#_M1005_s
+ N_A_27_74#_c_91_n N_A_27_74#_M1006_g N_A_27_74#_M1003_g N_A_27_74#_c_94_n
+ N_A_27_74#_c_95_n N_A_27_74#_c_102_n N_A_27_74#_c_96_n N_A_27_74#_c_97_n
+ N_A_27_74#_c_103_n N_A_27_74#_c_104_n N_A_27_74#_c_98_n N_A_27_74#_c_99_n
+ N_A_27_74#_c_100_n PM_SKY130_FD_SC_MS__O21BAI_1%A_27_74#
x_PM_SKY130_FD_SC_MS__O21BAI_1%A2 N_A2_M1007_g N_A2_M1004_g A2 A2 A2 A2
+ N_A2_c_168_n A2 PM_SKY130_FD_SC_MS__O21BAI_1%A2
x_PM_SKY130_FD_SC_MS__O21BAI_1%A1 N_A1_M1000_g N_A1_M1002_g A1 N_A1_c_210_n
+ N_A1_c_211_n PM_SKY130_FD_SC_MS__O21BAI_1%A1
x_PM_SKY130_FD_SC_MS__O21BAI_1%VPWR N_VPWR_M1005_d N_VPWR_M1000_d N_VPWR_c_236_n
+ N_VPWR_c_237_n N_VPWR_c_238_n VPWR N_VPWR_c_239_n N_VPWR_c_240_n
+ N_VPWR_c_241_n N_VPWR_c_235_n PM_SKY130_FD_SC_MS__O21BAI_1%VPWR
x_PM_SKY130_FD_SC_MS__O21BAI_1%Y N_Y_M1003_s N_Y_M1006_d N_Y_c_268_n N_Y_c_269_n
+ Y Y Y Y N_Y_c_270_n PM_SKY130_FD_SC_MS__O21BAI_1%Y
x_PM_SKY130_FD_SC_MS__O21BAI_1%VGND N_VGND_M1001_d N_VGND_M1004_d N_VGND_c_311_n
+ N_VGND_c_312_n VGND N_VGND_c_313_n N_VGND_c_314_n N_VGND_c_315_n
+ N_VGND_c_316_n N_VGND_c_317_n N_VGND_c_318_n PM_SKY130_FD_SC_MS__O21BAI_1%VGND
x_PM_SKY130_FD_SC_MS__O21BAI_1%A_308_74# N_A_308_74#_M1003_d N_A_308_74#_M1002_d
+ N_A_308_74#_c_349_n N_A_308_74#_c_350_n N_A_308_74#_c_351_n
+ N_A_308_74#_c_352_n PM_SKY130_FD_SC_MS__O21BAI_1%A_308_74#
cc_1 VNB N_B1_N_M1001_g 0.0548074f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.645
cc_2 VNB N_B1_N_c_61_n 0.0206119f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.02
cc_3 VNB N_B1_N_c_62_n 0.0105252f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.615
cc_4 VNB N_A_27_74#_c_91_n 0.0183564f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.54
cc_5 VNB N_A_27_74#_M1006_g 0.0102546f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.615
cc_6 VNB N_A_27_74#_M1003_g 0.0258899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_74#_c_94_n 0.00624997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_74#_c_95_n 0.0328912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_74#_c_96_n 0.00635589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_74#_c_97_n 0.0100794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_74#_c_98_n 0.0194928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_c_99_n 4.49976e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_74#_c_100_n 0.0361426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_M1007_g 0.00166758f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.645
cc_15 VNB N_A2_M1004_g 0.0218673f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.54
cc_16 VNB A2 0.00676042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A2_c_168_n 0.0281251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB A2 9.9768e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_M1000_g 0.00195314f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.645
cc_20 VNB N_A1_M1002_g 0.0294024f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.54
cc_21 VNB N_A1_c_210_n 0.0581712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A1_c_211_n 0.00431187f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.615
cc_23 VNB N_VPWR_c_235_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_268_n 0.00782665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_269_n 0.00507195f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_26 VNB N_Y_c_270_n 0.00363505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_311_n 0.014848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_312_n 0.00396562f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.615
cc_29 VNB N_VGND_c_313_n 0.0172318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_314_n 0.0312347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_315_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_316_n 0.196523f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_317_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_318_n 0.00622543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_308_74#_c_349_n 0.00178852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_308_74#_c_350_n 0.0121113f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.615
cc_37 VNB N_A_308_74#_c_351_n 0.0048099f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.615
cc_38 VNB N_A_308_74#_c_352_n 0.0247745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_B1_N_c_61_n 0.0629316f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.02
cc_40 VPB N_B1_N_c_62_n 0.0070275f $X=-0.19 $Y=1.66 $X2=0.4 $Y2=1.615
cc_41 VPB N_A_27_74#_M1006_g 0.0255498f $X=-0.19 $Y=1.66 $X2=0.4 $Y2=1.615
cc_42 VPB N_A_27_74#_c_102_n 0.0352562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_A_27_74#_c_103_n 0.0062701f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_A_27_74#_c_104_n 0.00956337f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_A_27_74#_c_99_n 0.00567328f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_A2_M1007_g 0.0236842f $X=-0.19 $Y=1.66 $X2=0.49 $Y2=0.645
cc_47 VPB A2 0.00308878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A1_M1000_g 0.0273412f $X=-0.19 $Y=1.66 $X2=0.49 $Y2=0.645
cc_49 VPB N_A1_c_211_n 0.00896873f $X=-0.19 $Y=1.66 $X2=0.4 $Y2=1.615
cc_50 VPB N_VPWR_c_236_n 0.0134879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_237_n 0.0103902f $X=-0.19 $Y=1.66 $X2=0.4 $Y2=1.615
cc_52 VPB N_VPWR_c_238_n 0.0498087f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.615
cc_53 VPB N_VPWR_c_239_n 0.0197879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_240_n 0.0342718f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_241_n 0.0128614f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_235_n 0.0599833f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB Y 0.0091875f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB Y 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_Y_c_270_n 0.00204394f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 N_B1_N_M1001_g N_A_27_74#_c_95_n 0.0108396f $X=0.49 $Y=0.645 $X2=0 $Y2=0
cc_61 N_B1_N_c_61_n N_A_27_74#_c_102_n 0.0194634f $X=0.525 $Y=2.02 $X2=0 $Y2=0
cc_62 N_B1_N_M1001_g N_A_27_74#_c_96_n 0.0172243f $X=0.49 $Y=0.645 $X2=0 $Y2=0
cc_63 N_B1_N_c_61_n N_A_27_74#_c_96_n 0.00218706f $X=0.525 $Y=2.02 $X2=0 $Y2=0
cc_64 N_B1_N_c_62_n N_A_27_74#_c_96_n 0.0148079f $X=0.4 $Y=1.615 $X2=0 $Y2=0
cc_65 N_B1_N_c_61_n N_A_27_74#_c_97_n 0.00291196f $X=0.525 $Y=2.02 $X2=0 $Y2=0
cc_66 N_B1_N_c_62_n N_A_27_74#_c_97_n 0.0202724f $X=0.4 $Y=1.615 $X2=0 $Y2=0
cc_67 N_B1_N_c_61_n N_A_27_74#_c_103_n 0.0146029f $X=0.525 $Y=2.02 $X2=0 $Y2=0
cc_68 N_B1_N_c_62_n N_A_27_74#_c_103_n 0.00710736f $X=0.4 $Y=1.615 $X2=0 $Y2=0
cc_69 N_B1_N_c_61_n N_A_27_74#_c_104_n 0.00938905f $X=0.525 $Y=2.02 $X2=0 $Y2=0
cc_70 N_B1_N_c_62_n N_A_27_74#_c_104_n 0.0280174f $X=0.4 $Y=1.615 $X2=0 $Y2=0
cc_71 N_B1_N_M1001_g N_A_27_74#_c_98_n 0.00425012f $X=0.49 $Y=0.645 $X2=0 $Y2=0
cc_72 N_B1_N_c_61_n N_A_27_74#_c_98_n 6.31941e-19 $X=0.525 $Y=2.02 $X2=0 $Y2=0
cc_73 N_B1_N_c_62_n N_A_27_74#_c_98_n 0.014171f $X=0.4 $Y=1.615 $X2=0 $Y2=0
cc_74 N_B1_N_c_61_n N_A_27_74#_c_99_n 0.00705846f $X=0.525 $Y=2.02 $X2=0 $Y2=0
cc_75 N_B1_N_c_62_n N_A_27_74#_c_99_n 0.0109803f $X=0.4 $Y=1.615 $X2=0 $Y2=0
cc_76 N_B1_N_M1001_g N_A_27_74#_c_100_n 0.0173988f $X=0.49 $Y=0.645 $X2=0 $Y2=0
cc_77 N_B1_N_c_62_n N_A_27_74#_c_100_n 2.01862e-19 $X=0.4 $Y=1.615 $X2=0 $Y2=0
cc_78 N_B1_N_c_61_n N_VPWR_c_236_n 0.00580638f $X=0.525 $Y=2.02 $X2=0 $Y2=0
cc_79 N_B1_N_c_61_n N_VPWR_c_239_n 0.005209f $X=0.525 $Y=2.02 $X2=0 $Y2=0
cc_80 N_B1_N_c_61_n N_VPWR_c_235_n 0.00990536f $X=0.525 $Y=2.02 $X2=0 $Y2=0
cc_81 N_B1_N_M1001_g N_Y_c_268_n 0.0014725f $X=0.49 $Y=0.645 $X2=0 $Y2=0
cc_82 N_B1_N_M1001_g N_Y_c_269_n 0.00454738f $X=0.49 $Y=0.645 $X2=0 $Y2=0
cc_83 N_B1_N_M1001_g N_VGND_c_311_n 0.018223f $X=0.49 $Y=0.645 $X2=0 $Y2=0
cc_84 N_B1_N_M1001_g N_VGND_c_313_n 0.00383152f $X=0.49 $Y=0.645 $X2=0 $Y2=0
cc_85 N_B1_N_M1001_g N_VGND_c_316_n 0.0076118f $X=0.49 $Y=0.645 $X2=0 $Y2=0
cc_86 N_A_27_74#_M1006_g N_A2_M1007_g 0.0180396f $X=1.45 $Y=2.4 $X2=0 $Y2=0
cc_87 N_A_27_74#_M1003_g N_A2_M1004_g 0.0135343f $X=1.465 $Y=0.74 $X2=0 $Y2=0
cc_88 N_A_27_74#_c_94_n A2 0.00121312f $X=1.45 $Y=1.375 $X2=0 $Y2=0
cc_89 N_A_27_74#_c_94_n N_A2_c_168_n 0.0208451f $X=1.45 $Y=1.375 $X2=0 $Y2=0
cc_90 N_A_27_74#_c_103_n N_VPWR_M1005_d 0.00188126f $X=0.745 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_91 N_A_27_74#_M1006_g N_VPWR_c_236_n 0.0189584f $X=1.45 $Y=2.4 $X2=0 $Y2=0
cc_92 N_A_27_74#_c_102_n N_VPWR_c_236_n 0.0267701f $X=0.3 $Y=2.265 $X2=0 $Y2=0
cc_93 N_A_27_74#_c_103_n N_VPWR_c_236_n 0.0226871f $X=0.745 $Y=2.035 $X2=0 $Y2=0
cc_94 N_A_27_74#_c_98_n N_VPWR_c_236_n 0.00622181f $X=0.83 $Y=1.63 $X2=0 $Y2=0
cc_95 N_A_27_74#_c_100_n N_VPWR_c_236_n 0.00166955f $X=0.97 $Y=1.375 $X2=0 $Y2=0
cc_96 N_A_27_74#_c_102_n N_VPWR_c_239_n 0.014549f $X=0.3 $Y=2.265 $X2=0 $Y2=0
cc_97 N_A_27_74#_M1006_g N_VPWR_c_240_n 0.00481245f $X=1.45 $Y=2.4 $X2=0 $Y2=0
cc_98 N_A_27_74#_M1006_g N_VPWR_c_235_n 0.00859218f $X=1.45 $Y=2.4 $X2=0 $Y2=0
cc_99 N_A_27_74#_c_102_n N_VPWR_c_235_n 0.0119743f $X=0.3 $Y=2.265 $X2=0 $Y2=0
cc_100 N_A_27_74#_M1003_g N_Y_c_268_n 0.0107219f $X=1.465 $Y=0.74 $X2=0 $Y2=0
cc_101 N_A_27_74#_c_91_n N_Y_c_269_n 0.00697146f $X=1.36 $Y=1.375 $X2=0 $Y2=0
cc_102 N_A_27_74#_M1003_g N_Y_c_269_n 0.00313748f $X=1.465 $Y=0.74 $X2=0 $Y2=0
cc_103 N_A_27_74#_c_98_n N_Y_c_269_n 0.00594309f $X=0.83 $Y=1.63 $X2=0 $Y2=0
cc_104 N_A_27_74#_c_100_n N_Y_c_269_n 3.87822e-19 $X=0.97 $Y=1.375 $X2=0 $Y2=0
cc_105 N_A_27_74#_M1006_g Y 0.0149474f $X=1.45 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A_27_74#_M1006_g Y 0.0223073f $X=1.45 $Y=2.4 $X2=0 $Y2=0
cc_107 N_A_27_74#_c_103_n Y 0.00448678f $X=0.745 $Y=2.035 $X2=0 $Y2=0
cc_108 N_A_27_74#_c_91_n N_Y_c_270_n 0.00528353f $X=1.36 $Y=1.375 $X2=0 $Y2=0
cc_109 N_A_27_74#_M1006_g N_Y_c_270_n 0.0116052f $X=1.45 $Y=2.4 $X2=0 $Y2=0
cc_110 N_A_27_74#_M1003_g N_Y_c_270_n 0.00642503f $X=1.465 $Y=0.74 $X2=0 $Y2=0
cc_111 N_A_27_74#_c_94_n N_Y_c_270_n 0.00362889f $X=1.45 $Y=1.375 $X2=0 $Y2=0
cc_112 N_A_27_74#_c_98_n N_Y_c_270_n 0.0326327f $X=0.83 $Y=1.63 $X2=0 $Y2=0
cc_113 N_A_27_74#_c_99_n N_Y_c_270_n 0.0112316f $X=0.83 $Y=1.95 $X2=0 $Y2=0
cc_114 N_A_27_74#_c_100_n N_Y_c_270_n 5.3485e-19 $X=0.97 $Y=1.375 $X2=0 $Y2=0
cc_115 N_A_27_74#_M1003_g N_VGND_c_311_n 0.00394308f $X=1.465 $Y=0.74 $X2=0
+ $Y2=0
cc_116 N_A_27_74#_c_95_n N_VGND_c_311_n 0.0226023f $X=0.275 $Y=0.645 $X2=0 $Y2=0
cc_117 N_A_27_74#_c_96_n N_VGND_c_311_n 0.0169933f $X=0.745 $Y=1.195 $X2=0 $Y2=0
cc_118 N_A_27_74#_c_98_n N_VGND_c_311_n 0.0116183f $X=0.83 $Y=1.63 $X2=0 $Y2=0
cc_119 N_A_27_74#_c_100_n N_VGND_c_311_n 3.25717e-19 $X=0.97 $Y=1.375 $X2=0
+ $Y2=0
cc_120 N_A_27_74#_M1003_g N_VGND_c_312_n 6.23092e-19 $X=1.465 $Y=0.74 $X2=0
+ $Y2=0
cc_121 N_A_27_74#_c_95_n N_VGND_c_313_n 0.011066f $X=0.275 $Y=0.645 $X2=0 $Y2=0
cc_122 N_A_27_74#_M1003_g N_VGND_c_314_n 0.00366292f $X=1.465 $Y=0.74 $X2=0
+ $Y2=0
cc_123 N_A_27_74#_M1003_g N_VGND_c_316_n 0.00606692f $X=1.465 $Y=0.74 $X2=0
+ $Y2=0
cc_124 N_A_27_74#_c_95_n N_VGND_c_316_n 0.00915947f $X=0.275 $Y=0.645 $X2=0
+ $Y2=0
cc_125 N_A_27_74#_M1003_g N_A_308_74#_c_349_n 0.00187536f $X=1.465 $Y=0.74 $X2=0
+ $Y2=0
cc_126 N_A_27_74#_M1003_g N_A_308_74#_c_351_n 6.78975e-19 $X=1.465 $Y=0.74 $X2=0
+ $Y2=0
cc_127 N_A2_M1007_g N_A1_M1000_g 0.0493347f $X=1.9 $Y=2.4 $X2=0 $Y2=0
cc_128 A2 N_A1_M1000_g 0.00816475f $X=2.16 $Y=1.665 $X2=0 $Y2=0
cc_129 N_A2_M1004_g N_A1_M1002_g 0.031308f $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_130 A2 N_A1_c_210_n 0.00280484f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_131 N_A2_c_168_n N_A1_c_210_n 0.0209448f $X=1.915 $Y=1.465 $X2=0 $Y2=0
cc_132 A2 N_A1_c_211_n 0.0270733f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_133 N_A2_c_168_n N_A1_c_211_n 2.28131e-19 $X=1.915 $Y=1.465 $X2=0 $Y2=0
cc_134 A2 N_A1_c_211_n 0.0114994f $X=2.16 $Y=1.665 $X2=0 $Y2=0
cc_135 N_A2_M1007_g N_VPWR_c_240_n 0.005209f $X=1.9 $Y=2.4 $X2=0 $Y2=0
cc_136 A2 N_VPWR_c_240_n 0.00659295f $X=2.16 $Y=1.665 $X2=0 $Y2=0
cc_137 N_A2_M1007_g N_VPWR_c_235_n 0.00983863f $X=1.9 $Y=2.4 $X2=0 $Y2=0
cc_138 A2 N_VPWR_c_235_n 0.0079425f $X=2.16 $Y=1.665 $X2=0 $Y2=0
cc_139 N_A2_M1004_g N_Y_c_269_n 9.65872e-19 $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A2_M1007_g Y 0.00271154f $X=1.9 $Y=2.4 $X2=0 $Y2=0
cc_141 A2 Y 0.00677064f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_142 N_A2_c_168_n Y 0.00138377f $X=1.915 $Y=1.465 $X2=0 $Y2=0
cc_143 A2 Y 0.0360598f $X=2.16 $Y=1.665 $X2=0 $Y2=0
cc_144 N_A2_M1007_g Y 0.0136842f $X=1.9 $Y=2.4 $X2=0 $Y2=0
cc_145 N_A2_M1007_g N_Y_c_270_n 6.60313e-19 $X=1.9 $Y=2.4 $X2=0 $Y2=0
cc_146 A2 N_Y_c_270_n 0.0165956f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_147 N_A2_c_168_n N_Y_c_270_n 3.78425e-19 $X=1.915 $Y=1.465 $X2=0 $Y2=0
cc_148 A2 N_Y_c_270_n 0.00555067f $X=2.16 $Y=1.665 $X2=0 $Y2=0
cc_149 A2 A_398_368# 0.0133933f $X=2.16 $Y=1.665 $X2=-0.19 $Y2=-0.245
cc_150 N_A2_M1004_g N_VGND_c_312_n 0.00803907f $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A2_M1004_g N_VGND_c_314_n 0.00383152f $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A2_M1004_g N_VGND_c_316_n 0.00758084f $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A2_M1004_g N_A_308_74#_c_349_n 4.4413e-19 $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A2_M1004_g N_A_308_74#_c_350_n 0.0125718f $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_155 A2 N_A_308_74#_c_350_n 0.0347779f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_156 N_A2_c_168_n N_A_308_74#_c_350_n 0.00279286f $X=1.915 $Y=1.465 $X2=0
+ $Y2=0
cc_157 A2 N_A_308_74#_c_351_n 0.00548166f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_158 N_A2_c_168_n N_A_308_74#_c_351_n 0.00153394f $X=1.915 $Y=1.465 $X2=0
+ $Y2=0
cc_159 N_A1_M1000_g N_VPWR_c_238_n 0.00536186f $X=2.38 $Y=2.4 $X2=0 $Y2=0
cc_160 N_A1_c_210_n N_VPWR_c_238_n 0.00135527f $X=2.61 $Y=1.465 $X2=0 $Y2=0
cc_161 N_A1_c_211_n N_VPWR_c_238_n 0.0219775f $X=2.61 $Y=1.465 $X2=0 $Y2=0
cc_162 N_A1_M1000_g N_VPWR_c_240_n 0.00553757f $X=2.38 $Y=2.4 $X2=0 $Y2=0
cc_163 N_A1_M1000_g N_VPWR_c_235_n 0.0109277f $X=2.38 $Y=2.4 $X2=0 $Y2=0
cc_164 N_A1_M1000_g Y 7.41969e-19 $X=2.38 $Y=2.4 $X2=0 $Y2=0
cc_165 N_A1_M1002_g N_VGND_c_312_n 0.0107652f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A1_M1002_g N_VGND_c_315_n 0.00383152f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A1_M1002_g N_VGND_c_316_n 0.00761198f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A1_M1002_g N_A_308_74#_c_350_n 0.0169051f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A1_c_210_n N_A_308_74#_c_350_n 0.00319341f $X=2.61 $Y=1.465 $X2=0 $Y2=0
cc_170 N_A1_c_211_n N_A_308_74#_c_350_n 0.0270164f $X=2.61 $Y=1.465 $X2=0 $Y2=0
cc_171 N_A1_M1002_g N_A_308_74#_c_352_n 0.00159319f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_172 N_VPWR_c_236_n Y 0.0271727f $X=1.14 $Y=2.455 $X2=0 $Y2=0
cc_173 N_VPWR_c_240_n Y 0.0159194f $X=2.52 $Y=3.33 $X2=0 $Y2=0
cc_174 N_VPWR_c_235_n Y 0.0129582f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_175 N_Y_c_268_n N_VGND_c_311_n 0.0421766f $X=1.25 $Y=0.515 $X2=0 $Y2=0
cc_176 N_Y_c_268_n N_VGND_c_314_n 0.0170618f $X=1.25 $Y=0.515 $X2=0 $Y2=0
cc_177 N_Y_c_268_n N_VGND_c_316_n 0.013925f $X=1.25 $Y=0.515 $X2=0 $Y2=0
cc_178 N_Y_c_268_n N_A_308_74#_c_349_n 0.0455845f $X=1.25 $Y=0.515 $X2=0 $Y2=0
cc_179 N_Y_c_269_n N_A_308_74#_c_351_n 0.0142394f $X=1.28 $Y=1.13 $X2=0 $Y2=0
cc_180 N_VGND_c_312_n N_A_308_74#_c_349_n 0.0125684f $X=2.165 $Y=0.515 $X2=0
+ $Y2=0
cc_181 N_VGND_c_314_n N_A_308_74#_c_349_n 0.00749631f $X=1.995 $Y=0 $X2=0 $Y2=0
cc_182 N_VGND_c_316_n N_A_308_74#_c_349_n 0.0062048f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_183 N_VGND_M1004_d N_A_308_74#_c_350_n 0.00234908f $X=2.02 $Y=0.37 $X2=0
+ $Y2=0
cc_184 N_VGND_c_312_n N_A_308_74#_c_350_n 0.0122946f $X=2.165 $Y=0.515 $X2=0
+ $Y2=0
cc_185 N_VGND_c_312_n N_A_308_74#_c_352_n 0.0126098f $X=2.165 $Y=0.515 $X2=0
+ $Y2=0
cc_186 N_VGND_c_315_n N_A_308_74#_c_352_n 0.011066f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_187 N_VGND_c_316_n N_A_308_74#_c_352_n 0.00915947f $X=2.64 $Y=0 $X2=0 $Y2=0

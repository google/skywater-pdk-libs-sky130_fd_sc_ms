* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dlygate4sd2_1 A VGND VNB VPB VPWR X
M1000 X a_405_138# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.968e+11p pd=2.77e+06u as=9.174e+11p ps=6.14e+06u
M1001 VPWR A a_28_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1002 a_288_74# a_28_74# VGND VNB nlowvt w=420000u l=180000u
+  ad=1.113e+11p pd=1.37e+06u as=5.258e+11p ps=4.42e+06u
M1003 VGND A a_28_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1004 VGND a_288_74# a_405_138# VNB nlowvt w=420000u l=180000u
+  ad=0p pd=0u as=2.436e+11p ps=2e+06u
M1005 X a_405_138# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1006 VPWR a_288_74# a_405_138# VPB pshort w=1e+06u l=250000u
+  ad=0p pd=0u as=5.1e+11p ps=3.02e+06u
M1007 a_288_74# a_28_74# VPWR VPB pshort w=1e+06u l=250000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
.ends

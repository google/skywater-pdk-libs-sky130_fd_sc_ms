* File: sky130_fd_sc_ms__o31a_2.pxi.spice
* Created: Wed Sep  2 12:25:35 2020
* 
x_PM_SKY130_FD_SC_MS__O31A_2%A_55_264# N_A_55_264#_M1003_d N_A_55_264#_M1000_d
+ N_A_55_264#_M1004_g N_A_55_264#_M1005_g N_A_55_264#_c_72_n N_A_55_264#_M1006_g
+ N_A_55_264#_M1011_g N_A_55_264#_c_75_n N_A_55_264#_c_76_n N_A_55_264#_c_91_p
+ N_A_55_264#_c_123_p N_A_55_264#_c_77_n N_A_55_264#_c_78_n N_A_55_264#_c_79_n
+ N_A_55_264#_c_85_n N_A_55_264#_c_80_n N_A_55_264#_c_87_n N_A_55_264#_c_81_n
+ PM_SKY130_FD_SC_MS__O31A_2%A_55_264#
x_PM_SKY130_FD_SC_MS__O31A_2%A1 N_A1_M1010_g N_A1_M1007_g A1 A1 N_A1_c_178_n
+ N_A1_c_179_n PM_SKY130_FD_SC_MS__O31A_2%A1
x_PM_SKY130_FD_SC_MS__O31A_2%A2 N_A2_M1002_g N_A2_M1009_g A2 A2 N_A2_c_219_n
+ PM_SKY130_FD_SC_MS__O31A_2%A2
x_PM_SKY130_FD_SC_MS__O31A_2%A3 N_A3_M1008_g N_A3_M1000_g A3 N_A3_c_255_n
+ N_A3_c_256_n PM_SKY130_FD_SC_MS__O31A_2%A3
x_PM_SKY130_FD_SC_MS__O31A_2%B1 N_B1_c_295_n N_B1_M1001_g N_B1_M1003_g
+ N_B1_c_292_n B1 N_B1_c_293_n N_B1_c_294_n PM_SKY130_FD_SC_MS__O31A_2%B1
x_PM_SKY130_FD_SC_MS__O31A_2%VPWR N_VPWR_M1004_s N_VPWR_M1011_s N_VPWR_M1001_d
+ N_VPWR_c_324_n N_VPWR_c_325_n N_VPWR_c_326_n N_VPWR_c_327_n N_VPWR_c_328_n
+ VPWR N_VPWR_c_329_n N_VPWR_c_330_n N_VPWR_c_331_n N_VPWR_c_323_n
+ PM_SKY130_FD_SC_MS__O31A_2%VPWR
x_PM_SKY130_FD_SC_MS__O31A_2%X N_X_M1005_s N_X_M1004_d N_X_c_366_n N_X_c_367_n
+ N_X_c_368_n X N_X_c_370_n PM_SKY130_FD_SC_MS__O31A_2%X
x_PM_SKY130_FD_SC_MS__O31A_2%VGND N_VGND_M1005_d N_VGND_M1006_d N_VGND_M1002_d
+ N_VGND_c_405_n N_VGND_c_406_n N_VGND_c_407_n N_VGND_c_408_n N_VGND_c_409_n
+ VGND N_VGND_c_410_n N_VGND_c_411_n N_VGND_c_412_n N_VGND_c_413_n
+ N_VGND_c_414_n PM_SKY130_FD_SC_MS__O31A_2%VGND
x_PM_SKY130_FD_SC_MS__O31A_2%A_328_74# N_A_328_74#_M1010_d N_A_328_74#_M1008_d
+ N_A_328_74#_c_453_n N_A_328_74#_c_454_n N_A_328_74#_c_463_n
+ N_A_328_74#_c_456_n PM_SKY130_FD_SC_MS__O31A_2%A_328_74#
cc_1 VNB N_A_55_264#_M1004_g 5.36566e-19 $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A_55_264#_M1005_g 0.028293f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_3 VNB N_A_55_264#_c_72_n 0.0148764f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.395
cc_4 VNB N_A_55_264#_M1006_g 0.0234109f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_5 VNB N_A_55_264#_M1011_g 0.00998306f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=2.4
cc_6 VNB N_A_55_264#_c_75_n 0.00779835f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=1.395
cc_7 VNB N_A_55_264#_c_76_n 5.59499e-19 $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=2.32
cc_8 VNB N_A_55_264#_c_77_n 0.0100559f $X=-0.19 $Y=-0.245 $X2=3.56 $Y2=0.96
cc_9 VNB N_A_55_264#_c_78_n 0.0264193f $X=-0.19 $Y=-0.245 $X2=3.56 $Y2=0.515
cc_10 VNB N_A_55_264#_c_79_n 0.0130668f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=1.485
cc_11 VNB N_A_55_264#_c_80_n 0.00441108f $X=-0.19 $Y=-0.245 $X2=2.995 $Y2=1.94
cc_12 VNB N_A_55_264#_c_81_n 0.0372417f $X=-0.19 $Y=-0.245 $X2=0.457 $Y2=1.395
cc_13 VNB N_A1_M1010_g 0.0273181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A1_c_178_n 0.026037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A1_c_179_n 0.00624344f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.395
cc_16 VNB N_A2_M1002_g 0.0336545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB A2 0.00275083f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_18 VNB N_A2_c_219_n 0.01856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A3_M1000_g 0.00649324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB A3 0.0105601f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_21 VNB N_A3_c_255_n 0.0324935f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.32
cc_22 VNB N_A3_c_256_n 0.0202699f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_23 VNB N_B1_M1003_g 0.0309473f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_24 VNB N_B1_c_292_n 0.00159338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_B1_c_293_n 0.0716888f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.32
cc_26 VNB N_B1_c_294_n 0.00435854f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_27 VNB N_VPWR_c_323_n 0.163682f $X=-0.19 $Y=-0.245 $X2=2.995 $Y2=2.405
cc_28 VNB N_X_c_366_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_29 VNB N_X_c_367_n 0.00291266f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_30 VNB N_X_c_368_n 0.00418437f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_31 VNB N_VGND_c_405_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_406_n 0.0477751f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_33 VNB N_VGND_c_407_n 0.021169f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.395
cc_34 VNB N_VGND_c_408_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=0.74
cc_35 VNB N_VGND_c_409_n 0.00673484f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=2.4
cc_36 VNB N_VGND_c_410_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.65
cc_37 VNB N_VGND_c_411_n 0.0384742f $X=-0.19 $Y=-0.245 $X2=3.56 $Y2=0.515
cc_38 VNB N_VGND_c_412_n 0.228611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_413_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_414_n 0.0073872f $X=-0.19 $Y=-0.245 $X2=2.995 $Y2=1.94
cc_41 VNB N_A_328_74#_c_453_n 0.00760749f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.65
cc_42 VNB N_A_328_74#_c_454_n 0.00280429f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_43 VPB N_A_55_264#_M1004_g 0.0252005f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_44 VPB N_A_55_264#_M1011_g 0.0239348f $X=-0.19 $Y=1.66 $X2=1.01 $Y2=2.4
cc_45 VPB N_A_55_264#_c_76_n 0.00756788f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=2.32
cc_46 VPB N_A_55_264#_c_85_n 0.00833193f $X=-0.19 $Y=1.66 $X2=2.93 $Y2=2.105
cc_47 VPB N_A_55_264#_c_80_n 0.00302977f $X=-0.19 $Y=1.66 $X2=2.995 $Y2=1.94
cc_48 VPB N_A_55_264#_c_87_n 0.0031255f $X=-0.19 $Y=1.66 $X2=2.93 $Y2=2.46
cc_49 VPB N_A1_M1007_g 0.0270884f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.65
cc_50 VPB N_A1_c_178_n 0.00560598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A1_c_179_n 0.00455356f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.395
cc_52 VPB N_A2_M1009_g 0.022375f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.65
cc_53 VPB A2 0.00171577f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_54 VPB N_A2_c_219_n 0.014176f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A3_M1000_g 0.0329816f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_B1_c_295_n 0.0288995f $X=-0.19 $Y=1.66 $X2=3.35 $Y2=0.37
cc_57 VPB N_B1_c_292_n 0.00731593f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_B1_c_294_n 0.00824274f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_59 VPB N_VPWR_c_324_n 0.0119967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_325_n 0.0214998f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_61 VPB N_VPWR_c_326_n 0.00447196f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.395
cc_62 VPB N_VPWR_c_327_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=0.74
cc_63 VPB N_VPWR_c_328_n 0.054016f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_329_n 0.0195091f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.65
cc_65 VPB N_VPWR_c_330_n 0.0534801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_331_n 0.009684f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_323_n 0.0651418f $X=-0.19 $Y=1.66 $X2=2.995 $Y2=2.405
cc_68 VPB N_X_c_367_n 0.00168814f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_69 VPB N_X_c_370_n 0.00237832f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 N_A_55_264#_M1006_g N_A1_M1010_g 0.0226424f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_71 N_A_55_264#_c_75_n N_A1_M1010_g 0.00111862f $X=1.01 $Y=1.395 $X2=0 $Y2=0
cc_72 N_A_55_264#_M1011_g N_A1_M1007_g 0.0339027f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_73 N_A_55_264#_c_91_p N_A1_M1007_g 0.0137395f $X=2.765 $Y=2.405 $X2=0 $Y2=0
cc_74 N_A_55_264#_c_75_n N_A1_c_178_n 0.0126756f $X=1.01 $Y=1.395 $X2=0 $Y2=0
cc_75 N_A_55_264#_c_91_p N_A1_c_178_n 3.5342e-19 $X=2.765 $Y=2.405 $X2=0 $Y2=0
cc_76 N_A_55_264#_M1011_g N_A1_c_179_n 0.00428383f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_77 N_A_55_264#_c_75_n N_A1_c_179_n 0.00139906f $X=1.01 $Y=1.395 $X2=0 $Y2=0
cc_78 N_A_55_264#_c_91_p N_A1_c_179_n 0.0211965f $X=2.765 $Y=2.405 $X2=0 $Y2=0
cc_79 N_A_55_264#_c_91_p N_A2_M1009_g 0.0136742f $X=2.765 $Y=2.405 $X2=0 $Y2=0
cc_80 N_A_55_264#_c_91_p A2 0.0211204f $X=2.765 $Y=2.405 $X2=0 $Y2=0
cc_81 N_A_55_264#_c_85_n A2 0.00455394f $X=2.93 $Y=2.105 $X2=0 $Y2=0
cc_82 N_A_55_264#_c_91_p N_A2_c_219_n 4.33455e-19 $X=2.765 $Y=2.405 $X2=0 $Y2=0
cc_83 N_A_55_264#_c_91_p N_A3_M1000_g 0.0174176f $X=2.765 $Y=2.405 $X2=0 $Y2=0
cc_84 N_A_55_264#_c_85_n N_A3_M1000_g 2.77713e-19 $X=2.93 $Y=2.105 $X2=0 $Y2=0
cc_85 N_A_55_264#_c_80_n N_A3_M1000_g 0.00708267f $X=2.995 $Y=1.94 $X2=0 $Y2=0
cc_86 N_A_55_264#_c_87_n N_A3_M1000_g 5.9741e-19 $X=2.93 $Y=2.46 $X2=0 $Y2=0
cc_87 N_A_55_264#_c_85_n A3 0.00541843f $X=2.93 $Y=2.105 $X2=0 $Y2=0
cc_88 N_A_55_264#_c_80_n A3 0.0281608f $X=2.995 $Y=1.94 $X2=0 $Y2=0
cc_89 N_A_55_264#_c_85_n N_A3_c_255_n 8.3549e-19 $X=2.93 $Y=2.105 $X2=0 $Y2=0
cc_90 N_A_55_264#_c_80_n N_A3_c_255_n 0.00194886f $X=2.995 $Y=1.94 $X2=0 $Y2=0
cc_91 N_A_55_264#_c_77_n N_A3_c_256_n 0.00396327f $X=3.56 $Y=0.96 $X2=0 $Y2=0
cc_92 N_A_55_264#_c_80_n N_A3_c_256_n 0.00100883f $X=2.995 $Y=1.94 $X2=0 $Y2=0
cc_93 N_A_55_264#_c_85_n N_B1_c_295_n 0.0107372f $X=2.93 $Y=2.105 $X2=-0.19
+ $Y2=-0.245
cc_94 N_A_55_264#_c_80_n N_B1_c_295_n 0.00887889f $X=2.995 $Y=1.94 $X2=-0.19
+ $Y2=-0.245
cc_95 N_A_55_264#_c_87_n N_B1_c_295_n 0.0105298f $X=2.93 $Y=2.46 $X2=-0.19
+ $Y2=-0.245
cc_96 N_A_55_264#_c_77_n N_B1_M1003_g 0.0191744f $X=3.56 $Y=0.96 $X2=0 $Y2=0
cc_97 N_A_55_264#_c_78_n N_B1_M1003_g 0.0122539f $X=3.56 $Y=0.515 $X2=0 $Y2=0
cc_98 N_A_55_264#_c_80_n N_B1_M1003_g 0.00855406f $X=2.995 $Y=1.94 $X2=0 $Y2=0
cc_99 N_A_55_264#_c_80_n N_B1_c_292_n 0.00394106f $X=2.995 $Y=1.94 $X2=0 $Y2=0
cc_100 N_A_55_264#_c_77_n N_B1_c_293_n 0.0043993f $X=3.56 $Y=0.96 $X2=0 $Y2=0
cc_101 N_A_55_264#_c_80_n N_B1_c_293_n 0.0105781f $X=2.995 $Y=1.94 $X2=0 $Y2=0
cc_102 N_A_55_264#_c_77_n N_B1_c_294_n 0.0254991f $X=3.56 $Y=0.96 $X2=0 $Y2=0
cc_103 N_A_55_264#_c_80_n N_B1_c_294_n 0.0348575f $X=2.995 $Y=1.94 $X2=0 $Y2=0
cc_104 N_A_55_264#_c_76_n N_VPWR_M1004_s 0.0205644f $X=0.31 $Y=2.32 $X2=-0.19
+ $Y2=-0.245
cc_105 N_A_55_264#_c_123_p N_VPWR_M1004_s 0.00920379f $X=0.395 $Y=2.405
+ $X2=-0.19 $Y2=-0.245
cc_106 N_A_55_264#_c_91_p N_VPWR_M1011_s 0.0154423f $X=2.765 $Y=2.405 $X2=0
+ $Y2=0
cc_107 N_A_55_264#_M1004_g N_VPWR_c_325_n 0.0123108f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_108 N_A_55_264#_M1011_g N_VPWR_c_325_n 0.00130701f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_109 N_A_55_264#_c_91_p N_VPWR_c_325_n 0.0021187f $X=2.765 $Y=2.405 $X2=0
+ $Y2=0
cc_110 N_A_55_264#_c_123_p N_VPWR_c_325_n 0.0116597f $X=0.395 $Y=2.405 $X2=0
+ $Y2=0
cc_111 N_A_55_264#_M1004_g N_VPWR_c_326_n 0.00130368f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_112 N_A_55_264#_M1011_g N_VPWR_c_326_n 0.0170227f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_113 N_A_55_264#_c_91_p N_VPWR_c_326_n 0.0322528f $X=2.765 $Y=2.405 $X2=0
+ $Y2=0
cc_114 N_A_55_264#_c_85_n N_VPWR_c_328_n 0.0819739f $X=2.93 $Y=2.105 $X2=0 $Y2=0
cc_115 N_A_55_264#_M1004_g N_VPWR_c_329_n 0.00460063f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_116 N_A_55_264#_M1011_g N_VPWR_c_329_n 0.00460063f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_117 N_A_55_264#_c_87_n N_VPWR_c_330_n 0.0200508f $X=2.93 $Y=2.46 $X2=0 $Y2=0
cc_118 N_A_55_264#_M1004_g N_VPWR_c_323_n 0.00461394f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_119 N_A_55_264#_M1011_g N_VPWR_c_323_n 0.00461394f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A_55_264#_c_91_p N_VPWR_c_323_n 0.058057f $X=2.765 $Y=2.405 $X2=0 $Y2=0
cc_121 N_A_55_264#_c_123_p N_VPWR_c_323_n 6.15054e-19 $X=0.395 $Y=2.405 $X2=0
+ $Y2=0
cc_122 N_A_55_264#_c_87_n N_VPWR_c_323_n 0.0162933f $X=2.93 $Y=2.46 $X2=0 $Y2=0
cc_123 N_A_55_264#_c_91_p N_X_M1004_d 0.00649057f $X=2.765 $Y=2.405 $X2=0 $Y2=0
cc_124 N_A_55_264#_M1005_g N_X_c_366_n 0.00772833f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A_55_264#_M1006_g N_X_c_366_n 0.00752022f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A_55_264#_M1004_g N_X_c_367_n 0.00140903f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_127 N_A_55_264#_M1005_g N_X_c_367_n 0.00408016f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A_55_264#_c_72_n N_X_c_367_n 0.00833621f $X=0.92 $Y=1.395 $X2=0 $Y2=0
cc_129 N_A_55_264#_M1006_g N_X_c_367_n 0.00495702f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A_55_264#_M1011_g N_X_c_367_n 0.00893795f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_131 N_A_55_264#_c_75_n N_X_c_367_n 0.00266977f $X=1.01 $Y=1.395 $X2=0 $Y2=0
cc_132 N_A_55_264#_c_76_n N_X_c_367_n 0.00731129f $X=0.31 $Y=2.32 $X2=0 $Y2=0
cc_133 N_A_55_264#_c_79_n N_X_c_367_n 0.0244835f $X=0.44 $Y=1.485 $X2=0 $Y2=0
cc_134 N_A_55_264#_c_81_n N_X_c_367_n 0.001226f $X=0.457 $Y=1.395 $X2=0 $Y2=0
cc_135 N_A_55_264#_M1005_g N_X_c_368_n 0.00316168f $X=0.565 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A_55_264#_c_72_n N_X_c_368_n 0.00181038f $X=0.92 $Y=1.395 $X2=0 $Y2=0
cc_137 N_A_55_264#_M1006_g N_X_c_368_n 0.00193058f $X=0.995 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A_55_264#_M1004_g N_X_c_370_n 0.00494228f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A_55_264#_c_72_n N_X_c_370_n 0.00512017f $X=0.92 $Y=1.395 $X2=0 $Y2=0
cc_140 N_A_55_264#_M1011_g N_X_c_370_n 0.00697918f $X=1.01 $Y=2.4 $X2=0 $Y2=0
cc_141 N_A_55_264#_c_76_n N_X_c_370_n 0.013351f $X=0.31 $Y=2.32 $X2=0 $Y2=0
cc_142 N_A_55_264#_c_91_p N_X_c_370_n 0.0203347f $X=2.765 $Y=2.405 $X2=0 $Y2=0
cc_143 N_A_55_264#_c_79_n N_X_c_370_n 0.00304274f $X=0.44 $Y=1.485 $X2=0 $Y2=0
cc_144 N_A_55_264#_c_81_n N_X_c_370_n 0.00182001f $X=0.457 $Y=1.395 $X2=0 $Y2=0
cc_145 N_A_55_264#_c_91_p A_349_392# 0.00734082f $X=2.765 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_146 N_A_55_264#_c_91_p A_433_392# 0.0137232f $X=2.765 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_147 N_A_55_264#_M1005_g N_VGND_c_406_n 0.0184907f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_148 N_A_55_264#_c_79_n N_VGND_c_406_n 0.0171976f $X=0.44 $Y=1.485 $X2=0 $Y2=0
cc_149 N_A_55_264#_c_81_n N_VGND_c_406_n 0.00400955f $X=0.457 $Y=1.395 $X2=0
+ $Y2=0
cc_150 N_A_55_264#_M1006_g N_VGND_c_407_n 0.00666821f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_151 N_A_55_264#_M1005_g N_VGND_c_410_n 0.00434272f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_152 N_A_55_264#_M1006_g N_VGND_c_410_n 0.00434272f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_153 N_A_55_264#_c_78_n N_VGND_c_411_n 0.0145203f $X=3.56 $Y=0.515 $X2=0 $Y2=0
cc_154 N_A_55_264#_M1005_g N_VGND_c_412_n 0.00823934f $X=0.565 $Y=0.74 $X2=0
+ $Y2=0
cc_155 N_A_55_264#_M1006_g N_VGND_c_412_n 0.00821312f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_156 N_A_55_264#_c_78_n N_VGND_c_412_n 0.0120696f $X=3.56 $Y=0.515 $X2=0 $Y2=0
cc_157 N_A_55_264#_c_77_n N_A_328_74#_M1008_d 0.00329864f $X=3.56 $Y=0.96 $X2=0
+ $Y2=0
cc_158 N_A_55_264#_c_77_n N_A_328_74#_c_456_n 0.00855261f $X=3.56 $Y=0.96 $X2=0
+ $Y2=0
cc_159 N_A1_M1010_g N_A2_M1002_g 0.0252626f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A1_c_178_n N_A2_M1002_g 0.0472489f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_161 N_A1_c_179_n N_A2_M1002_g 0.00627802f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_162 N_A1_c_178_n A2 7.90645e-19 $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_163 N_A1_c_179_n A2 0.0425296f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_164 N_A1_M1007_g N_A2_c_219_n 0.0472489f $X=1.655 $Y=2.46 $X2=0 $Y2=0
cc_165 N_A1_c_179_n N_VPWR_M1011_s 0.00365787f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_166 N_A1_M1007_g N_VPWR_c_326_n 0.0167351f $X=1.655 $Y=2.46 $X2=0 $Y2=0
cc_167 N_A1_M1007_g N_VPWR_c_330_n 0.00460063f $X=1.655 $Y=2.46 $X2=0 $Y2=0
cc_168 N_A1_M1007_g N_VPWR_c_323_n 0.00460677f $X=1.655 $Y=2.46 $X2=0 $Y2=0
cc_169 N_A1_M1010_g N_X_c_366_n 0.00115542f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A1_c_178_n N_X_c_367_n 0.00104954f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_171 N_A1_c_179_n N_X_c_367_n 0.015435f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_172 N_A1_M1007_g N_X_c_370_n 2.80273e-19 $X=1.655 $Y=2.46 $X2=0 $Y2=0
cc_173 N_A1_c_179_n N_X_c_370_n 0.0122114f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_174 N_A1_M1010_g N_VGND_c_407_n 0.00666787f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A1_c_178_n N_VGND_c_407_n 2.14662e-19 $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_176 N_A1_c_179_n N_VGND_c_407_n 0.00205464f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_177 N_A1_M1010_g N_VGND_c_408_n 0.00434272f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A1_M1010_g N_VGND_c_409_n 4.1081e-19 $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A1_M1010_g N_VGND_c_412_n 0.00821983f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_180 N_A1_M1010_g N_A_328_74#_c_453_n 0.00437183f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_181 N_A1_c_178_n N_A_328_74#_c_453_n 7.965e-19 $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_182 N_A1_c_179_n N_A_328_74#_c_453_n 0.0132489f $X=1.58 $Y=1.515 $X2=0 $Y2=0
cc_183 N_A1_M1010_g N_A_328_74#_c_454_n 0.00549371f $X=1.565 $Y=0.74 $X2=0 $Y2=0
cc_184 N_A2_M1009_g N_A3_M1000_g 0.0407802f $X=2.075 $Y=2.46 $X2=0 $Y2=0
cc_185 A2 N_A3_M1000_g 0.0068079f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_186 N_A2_M1002_g A3 0.00565381f $X=2.06 $Y=0.74 $X2=0 $Y2=0
cc_187 A2 A3 0.00544377f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_188 N_A2_c_219_n A3 4.91538e-19 $X=2.15 $Y=1.635 $X2=0 $Y2=0
cc_189 N_A2_c_219_n N_A3_c_255_n 0.018352f $X=2.15 $Y=1.635 $X2=0 $Y2=0
cc_190 N_A2_M1002_g N_A3_c_256_n 0.0270404f $X=2.06 $Y=0.74 $X2=0 $Y2=0
cc_191 N_A2_M1009_g N_VPWR_c_326_n 0.00206847f $X=2.075 $Y=2.46 $X2=0 $Y2=0
cc_192 N_A2_M1009_g N_VPWR_c_330_n 0.00553757f $X=2.075 $Y=2.46 $X2=0 $Y2=0
cc_193 N_A2_M1009_g N_VPWR_c_323_n 0.00557035f $X=2.075 $Y=2.46 $X2=0 $Y2=0
cc_194 A2 A_433_392# 0.00353488f $X=2.075 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_195 N_A2_M1002_g N_VGND_c_408_n 0.00398535f $X=2.06 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A2_M1002_g N_VGND_c_409_n 0.00710985f $X=2.06 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A2_M1002_g N_VGND_c_412_n 0.00384527f $X=2.06 $Y=0.74 $X2=0 $Y2=0
cc_198 N_A2_M1002_g N_A_328_74#_c_453_n 0.00143395f $X=2.06 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A2_M1002_g N_A_328_74#_c_454_n 0.00224861f $X=2.06 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A2_M1002_g N_A_328_74#_c_463_n 0.0142189f $X=2.06 $Y=0.74 $X2=0 $Y2=0
cc_201 A2 N_A_328_74#_c_463_n 0.00933039f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_202 N_A2_c_219_n N_A_328_74#_c_463_n 7.71987e-19 $X=2.15 $Y=1.635 $X2=0 $Y2=0
cc_203 N_A2_M1002_g N_A_328_74#_c_456_n 5.02222e-19 $X=2.06 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A3_M1000_g N_B1_c_295_n 0.00979394f $X=2.645 $Y=2.46 $X2=-0.19
+ $Y2=-0.245
cc_205 N_A3_c_255_n N_B1_M1003_g 0.002904f $X=2.72 $Y=1.385 $X2=0 $Y2=0
cc_206 N_A3_c_256_n N_B1_M1003_g 0.0197735f $X=2.72 $Y=1.22 $X2=0 $Y2=0
cc_207 N_A3_M1000_g N_B1_c_293_n 0.00641549f $X=2.645 $Y=2.46 $X2=0 $Y2=0
cc_208 A3 N_B1_c_293_n 2.74107e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_209 N_A3_c_255_n N_B1_c_293_n 0.0132146f $X=2.72 $Y=1.385 $X2=0 $Y2=0
cc_210 N_A3_M1000_g N_VPWR_c_330_n 0.00553757f $X=2.645 $Y=2.46 $X2=0 $Y2=0
cc_211 N_A3_M1000_g N_VPWR_c_323_n 0.00558121f $X=2.645 $Y=2.46 $X2=0 $Y2=0
cc_212 N_A3_c_256_n N_VGND_c_409_n 0.0052684f $X=2.72 $Y=1.22 $X2=0 $Y2=0
cc_213 N_A3_c_256_n N_VGND_c_411_n 0.0043552f $X=2.72 $Y=1.22 $X2=0 $Y2=0
cc_214 N_A3_c_256_n N_VGND_c_412_n 0.00436921f $X=2.72 $Y=1.22 $X2=0 $Y2=0
cc_215 A3 N_A_328_74#_c_463_n 0.0078091f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_216 N_A3_c_256_n N_A_328_74#_c_463_n 0.00931502f $X=2.72 $Y=1.22 $X2=0 $Y2=0
cc_217 A3 N_A_328_74#_c_456_n 0.010823f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_218 N_A3_c_255_n N_A_328_74#_c_456_n 9.87449e-19 $X=2.72 $Y=1.385 $X2=0 $Y2=0
cc_219 N_A3_c_256_n N_A_328_74#_c_456_n 0.01381f $X=2.72 $Y=1.22 $X2=0 $Y2=0
cc_220 N_B1_c_295_n N_VPWR_c_328_n 0.0264142f $X=3.185 $Y=1.88 $X2=0 $Y2=0
cc_221 N_B1_c_293_n N_VPWR_c_328_n 0.00181048f $X=3.56 $Y=1.465 $X2=0 $Y2=0
cc_222 N_B1_c_294_n N_VPWR_c_328_n 0.0299469f $X=3.56 $Y=1.465 $X2=0 $Y2=0
cc_223 N_B1_c_295_n N_VPWR_c_330_n 0.00407599f $X=3.185 $Y=1.88 $X2=0 $Y2=0
cc_224 N_B1_c_295_n N_VPWR_c_323_n 0.00621559f $X=3.185 $Y=1.88 $X2=0 $Y2=0
cc_225 N_B1_M1003_g N_VGND_c_411_n 0.0043552f $X=3.275 $Y=0.74 $X2=0 $Y2=0
cc_226 N_B1_M1003_g N_VGND_c_412_n 0.00825941f $X=3.275 $Y=0.74 $X2=0 $Y2=0
cc_227 N_B1_M1003_g N_A_328_74#_c_456_n 0.0115428f $X=3.275 $Y=0.74 $X2=0 $Y2=0
cc_228 N_X_c_366_n N_VGND_c_406_n 0.0308109f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_229 N_X_c_366_n N_VGND_c_407_n 0.0308109f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_230 N_X_c_366_n N_VGND_c_410_n 0.0144922f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_231 N_X_c_366_n N_VGND_c_412_n 0.0118826f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_232 N_VGND_c_407_n N_A_328_74#_c_453_n 0.0151247f $X=1.28 $Y=0.515 $X2=0
+ $Y2=0
cc_233 N_VGND_c_407_n N_A_328_74#_c_454_n 0.0165124f $X=1.28 $Y=0.515 $X2=0
+ $Y2=0
cc_234 N_VGND_c_408_n N_A_328_74#_c_454_n 0.0145639f $X=2.115 $Y=0 $X2=0 $Y2=0
cc_235 N_VGND_c_409_n N_A_328_74#_c_454_n 0.0104328f $X=2.31 $Y=0.515 $X2=0
+ $Y2=0
cc_236 N_VGND_c_412_n N_A_328_74#_c_454_n 0.0119984f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_237 N_VGND_M1002_d N_A_328_74#_c_463_n 0.0126964f $X=2.135 $Y=0.37 $X2=0
+ $Y2=0
cc_238 N_VGND_c_409_n N_A_328_74#_c_463_n 0.0255658f $X=2.31 $Y=0.515 $X2=0
+ $Y2=0
cc_239 N_VGND_c_412_n N_A_328_74#_c_463_n 0.0120739f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_240 N_VGND_c_411_n N_A_328_74#_c_456_n 0.0140542f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_241 N_VGND_c_412_n N_A_328_74#_c_456_n 0.0180651f $X=3.6 $Y=0 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__a21boi_2.pxi.spice
* Created: Fri Aug 28 16:58:47 2020
* 
x_PM_SKY130_FD_SC_MS__A21BOI_2%B1_N N_B1_N_M1010_g N_B1_N_M1003_g N_B1_N_c_84_n
+ N_B1_N_c_85_n B1_N PM_SKY130_FD_SC_MS__A21BOI_2%B1_N
x_PM_SKY130_FD_SC_MS__A21BOI_2%A_62_94# N_A_62_94#_M1003_s N_A_62_94#_M1010_d
+ N_A_62_94#_M1006_g N_A_62_94#_c_124_n N_A_62_94#_M1001_g N_A_62_94#_M1011_g
+ N_A_62_94#_c_118_n N_A_62_94#_c_119_n N_A_62_94#_c_127_n N_A_62_94#_M1002_g
+ N_A_62_94#_c_120_n N_A_62_94#_c_121_n N_A_62_94#_c_122_n N_A_62_94#_c_128_n
+ N_A_62_94#_c_129_n N_A_62_94#_c_123_n N_A_62_94#_c_130_n
+ PM_SKY130_FD_SC_MS__A21BOI_2%A_62_94#
x_PM_SKY130_FD_SC_MS__A21BOI_2%A1 N_A1_M1004_g N_A1_M1000_g N_A1_M1005_g
+ N_A1_M1012_g A1 N_A1_c_200_n N_A1_c_201_n PM_SKY130_FD_SC_MS__A21BOI_2%A1
x_PM_SKY130_FD_SC_MS__A21BOI_2%A2 N_A2_M1008_g N_A2_c_255_n N_A2_M1007_g
+ N_A2_c_256_n N_A2_M1013_g N_A2_M1009_g A2 N_A2_c_259_n
+ PM_SKY130_FD_SC_MS__A21BOI_2%A2
x_PM_SKY130_FD_SC_MS__A21BOI_2%VPWR N_VPWR_M1010_s N_VPWR_M1004_d N_VPWR_M1008_d
+ N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_302_n VPWR
+ N_VPWR_c_303_n N_VPWR_c_304_n N_VPWR_c_305_n N_VPWR_c_298_n N_VPWR_c_307_n
+ N_VPWR_c_308_n PM_SKY130_FD_SC_MS__A21BOI_2%VPWR
x_PM_SKY130_FD_SC_MS__A21BOI_2%A_241_368# N_A_241_368#_M1001_s
+ N_A_241_368#_M1002_s N_A_241_368#_M1005_s N_A_241_368#_M1009_s
+ N_A_241_368#_c_351_n N_A_241_368#_c_352_n N_A_241_368#_c_353_n
+ N_A_241_368#_c_354_n N_A_241_368#_c_370_n N_A_241_368#_c_355_n
+ N_A_241_368#_c_356_n N_A_241_368#_c_357_n N_A_241_368#_c_358_n
+ PM_SKY130_FD_SC_MS__A21BOI_2%A_241_368#
x_PM_SKY130_FD_SC_MS__A21BOI_2%Y N_Y_M1006_d N_Y_M1000_s N_Y_M1001_d N_Y_c_410_n
+ N_Y_c_411_n N_Y_c_412_n N_Y_c_413_n N_Y_c_414_n Y N_Y_c_415_n N_Y_c_416_n
+ PM_SKY130_FD_SC_MS__A21BOI_2%Y
x_PM_SKY130_FD_SC_MS__A21BOI_2%VGND N_VGND_M1003_d N_VGND_M1011_s N_VGND_M1007_d
+ N_VGND_c_466_n N_VGND_c_467_n N_VGND_c_468_n N_VGND_c_469_n N_VGND_c_470_n
+ N_VGND_c_471_n VGND N_VGND_c_472_n N_VGND_c_473_n N_VGND_c_474_n
+ N_VGND_c_475_n N_VGND_c_476_n PM_SKY130_FD_SC_MS__A21BOI_2%VGND
x_PM_SKY130_FD_SC_MS__A21BOI_2%A_436_74# N_A_436_74#_M1000_d N_A_436_74#_M1012_d
+ N_A_436_74#_M1013_s N_A_436_74#_c_525_n N_A_436_74#_c_526_n
+ N_A_436_74#_c_538_n N_A_436_74#_c_532_n N_A_436_74#_c_527_n
+ N_A_436_74#_c_528_n PM_SKY130_FD_SC_MS__A21BOI_2%A_436_74#
cc_1 VNB N_B1_N_M1003_g 0.0389049f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.79
cc_2 VNB N_B1_N_c_84_n 0.0255356f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.615
cc_3 VNB N_B1_N_c_85_n 0.0118108f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.615
cc_4 VNB B1_N 0.0085963f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_5 VNB N_A_62_94#_M1006_g 0.0238777f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.615
cc_6 VNB N_A_62_94#_M1011_g 0.0256721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_62_94#_c_118_n 0.0155409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_62_94#_c_119_n 0.0485631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_62_94#_c_120_n 0.0274788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_62_94#_c_121_n 0.00519287f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_62_94#_c_122_n 0.00946887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_62_94#_c_123_n 0.0170134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_M1004_g 4.57023e-19 $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.46
cc_14 VNB N_A1_M1000_g 0.0246159f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=0.79
cc_15 VNB N_A1_M1005_g 4.92602e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_16 VNB N_A1_M1012_g 0.0222596f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.615
cc_17 VNB N_A1_c_200_n 0.00102877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_c_201_n 0.0474278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A2_M1008_g 0.00608326f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.46
cc_20 VNB N_A2_c_255_n 0.0168884f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.45
cc_21 VNB N_A2_c_256_n 0.0224993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A2_M1009_g 0.00926004f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.615
cc_23 VNB A2 0.00752679f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.615
cc_24 VNB N_A2_c_259_n 0.0526892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_298_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_410_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_411_n 0.00252401f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.615
cc_28 VNB N_Y_c_412_n 0.00316101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_413_n 0.00314005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_414_n 0.00402553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_415_n 0.00185509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_416_n 0.0220781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_466_n 0.00948899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_467_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_468_n 0.0117687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_469_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_470_n 0.0247362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_471_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_472_n 0.0382181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_473_n 0.0178682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_474_n 0.267893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_475_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_476_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_436_74#_c_525_n 0.00820512f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.615
cc_45 VNB N_A_436_74#_c_526_n 0.00160668f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.615
cc_46 VNB N_A_436_74#_c_527_n 0.0159805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_436_74#_c_528_n 0.0207145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VPB N_B1_N_M1010_g 0.0312046f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=2.46
cc_49 VPB N_B1_N_c_84_n 0.0189871f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.615
cc_50 VPB N_B1_N_c_85_n 0.00718035f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.615
cc_51 VPB B1_N 0.00521552f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_52 VPB N_A_62_94#_c_124_n 0.0185501f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_53 VPB N_A_62_94#_c_118_n 0.00961598f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_62_94#_c_119_n 0.00541458f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_62_94#_c_127_n 0.0157683f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_62_94#_c_128_n 0.00317516f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_62_94#_c_129_n 0.0104044f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_62_94#_c_130_n 0.00596926f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A1_M1004_g 0.0218312f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=2.46
cc_60 VPB N_A1_M1005_g 0.0222953f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_61 VPB N_A1_c_200_n 0.00347442f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A2_M1008_g 0.0213936f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=2.46
cc_63 VPB N_A2_M1009_g 0.0282484f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.615
cc_64 VPB N_VPWR_c_299_n 0.013204f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.615
cc_65 VPB N_VPWR_c_300_n 0.0517177f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_301_n 0.00329129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_302_n 0.00329222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_303_n 0.0519887f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_304_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_305_n 0.0177091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_298_n 0.0777528f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_307_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_308_n 0.00638264f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_241_368#_c_351_n 0.0113975f $X=-0.19 $Y=1.66 $X2=0.31 $Y2=1.615
cc_75 VPB N_A_241_368#_c_352_n 0.00474121f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_241_368#_c_353_n 0.00440836f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_241_368#_c_354_n 0.00318834f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_241_368#_c_355_n 0.00179594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_241_368#_c_356_n 0.0175857f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_A_241_368#_c_357_n 0.0431963f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_A_241_368#_c_358_n 0.00491856f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 N_B1_N_M1003_g N_A_62_94#_M1006_g 0.0146457f $X=0.65 $Y=0.79 $X2=0 $Y2=0
cc_83 N_B1_N_c_85_n N_A_62_94#_c_119_n 0.0146457f $X=0.61 $Y=1.615 $X2=0 $Y2=0
cc_84 N_B1_N_M1003_g N_A_62_94#_c_120_n 4.61877e-19 $X=0.65 $Y=0.79 $X2=0 $Y2=0
cc_85 N_B1_N_M1003_g N_A_62_94#_c_121_n 0.0194717f $X=0.65 $Y=0.79 $X2=0 $Y2=0
cc_86 N_B1_N_c_85_n N_A_62_94#_c_121_n 0.0022655f $X=0.61 $Y=1.615 $X2=0 $Y2=0
cc_87 N_B1_N_c_84_n N_A_62_94#_c_122_n 0.00685382f $X=0.495 $Y=1.615 $X2=0 $Y2=0
cc_88 B1_N N_A_62_94#_c_122_n 0.0172883f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_89 N_B1_N_M1010_g N_A_62_94#_c_128_n 0.00358321f $X=0.585 $Y=2.46 $X2=0 $Y2=0
cc_90 N_B1_N_c_85_n N_A_62_94#_c_128_n 0.0017226f $X=0.61 $Y=1.615 $X2=0 $Y2=0
cc_91 N_B1_N_M1010_g N_A_62_94#_c_129_n 0.0116145f $X=0.585 $Y=2.46 $X2=0 $Y2=0
cc_92 N_B1_N_M1003_g N_A_62_94#_c_123_n 0.00745999f $X=0.65 $Y=0.79 $X2=0 $Y2=0
cc_93 B1_N N_A_62_94#_c_123_n 0.0101785f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_94 N_B1_N_M1010_g N_A_62_94#_c_130_n 0.00580403f $X=0.585 $Y=2.46 $X2=0 $Y2=0
cc_95 N_B1_N_c_85_n N_A_62_94#_c_130_n 0.0039252f $X=0.61 $Y=1.615 $X2=0 $Y2=0
cc_96 B1_N N_A_62_94#_c_130_n 0.00592225f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_97 N_B1_N_M1010_g N_VPWR_c_300_n 0.00525184f $X=0.585 $Y=2.46 $X2=0 $Y2=0
cc_98 N_B1_N_c_84_n N_VPWR_c_300_n 0.00577732f $X=0.495 $Y=1.615 $X2=0 $Y2=0
cc_99 B1_N N_VPWR_c_300_n 0.0209147f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_100 N_B1_N_M1010_g N_VPWR_c_303_n 0.005209f $X=0.585 $Y=2.46 $X2=0 $Y2=0
cc_101 N_B1_N_M1010_g N_VPWR_c_298_n 0.00991388f $X=0.585 $Y=2.46 $X2=0 $Y2=0
cc_102 N_B1_N_M1010_g N_A_241_368#_c_351_n 0.00146587f $X=0.585 $Y=2.46 $X2=0
+ $Y2=0
cc_103 N_B1_N_M1010_g N_A_241_368#_c_353_n 0.00302726f $X=0.585 $Y=2.46 $X2=0
+ $Y2=0
cc_104 N_B1_N_M1003_g N_VGND_c_466_n 0.00577735f $X=0.65 $Y=0.79 $X2=0 $Y2=0
cc_105 N_B1_N_M1003_g N_VGND_c_470_n 0.00507111f $X=0.65 $Y=0.79 $X2=0 $Y2=0
cc_106 N_B1_N_M1003_g N_VGND_c_474_n 0.00514438f $X=0.65 $Y=0.79 $X2=0 $Y2=0
cc_107 N_A_62_94#_c_127_n N_A1_M1004_g 0.00912097f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_108 N_A_62_94#_c_118_n N_A1_c_200_n 6.16883e-19 $X=1.915 $Y=1.69 $X2=0 $Y2=0
cc_109 N_A_62_94#_c_118_n N_A1_c_201_n 0.00912097f $X=1.915 $Y=1.69 $X2=0 $Y2=0
cc_110 N_A_62_94#_c_119_n N_A1_c_201_n 0.00305683f $X=1.645 $Y=1.69 $X2=0 $Y2=0
cc_111 N_A_62_94#_c_128_n N_VPWR_c_300_n 0.034897f $X=0.81 $Y=2.105 $X2=0 $Y2=0
cc_112 N_A_62_94#_c_124_n N_VPWR_c_303_n 0.00333926f $X=1.555 $Y=1.765 $X2=0
+ $Y2=0
cc_113 N_A_62_94#_c_127_n N_VPWR_c_303_n 0.00333926f $X=2.005 $Y=1.765 $X2=0
+ $Y2=0
cc_114 N_A_62_94#_c_129_n N_VPWR_c_303_n 0.014549f $X=0.81 $Y=2.815 $X2=0 $Y2=0
cc_115 N_A_62_94#_c_124_n N_VPWR_c_298_n 0.0042782f $X=1.555 $Y=1.765 $X2=0
+ $Y2=0
cc_116 N_A_62_94#_c_127_n N_VPWR_c_298_n 0.00422798f $X=2.005 $Y=1.765 $X2=0
+ $Y2=0
cc_117 N_A_62_94#_c_129_n N_VPWR_c_298_n 0.0119743f $X=0.81 $Y=2.815 $X2=0 $Y2=0
cc_118 N_A_62_94#_c_124_n N_A_241_368#_c_351_n 0.00147311f $X=1.555 $Y=1.765
+ $X2=0 $Y2=0
cc_119 N_A_62_94#_c_119_n N_A_241_368#_c_351_n 0.00240798f $X=1.645 $Y=1.69
+ $X2=0 $Y2=0
cc_120 N_A_62_94#_c_123_n N_A_241_368#_c_351_n 0.0194066f $X=0.89 $Y=1.65 $X2=0
+ $Y2=0
cc_121 N_A_62_94#_c_130_n N_A_241_368#_c_351_n 0.0812754f $X=0.81 $Y=1.94 $X2=0
+ $Y2=0
cc_122 N_A_62_94#_c_124_n N_A_241_368#_c_352_n 0.01495f $X=1.555 $Y=1.765 $X2=0
+ $Y2=0
cc_123 N_A_62_94#_c_127_n N_A_241_368#_c_352_n 0.0137017f $X=2.005 $Y=1.765
+ $X2=0 $Y2=0
cc_124 N_A_62_94#_c_129_n N_A_241_368#_c_353_n 0.00613234f $X=0.81 $Y=2.815
+ $X2=0 $Y2=0
cc_125 N_A_62_94#_M1006_g N_Y_c_410_n 3.92313e-19 $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A_62_94#_M1011_g N_Y_c_410_n 3.92313e-19 $X=1.57 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A_62_94#_M1006_g N_Y_c_411_n 4.14962e-19 $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_128 N_A_62_94#_c_119_n N_Y_c_411_n 0.00101398f $X=1.645 $Y=1.69 $X2=0 $Y2=0
cc_129 N_A_62_94#_c_123_n N_Y_c_411_n 0.0131103f $X=0.89 $Y=1.65 $X2=0 $Y2=0
cc_130 N_A_62_94#_c_124_n N_Y_c_412_n 0.013941f $X=1.555 $Y=1.765 $X2=0 $Y2=0
cc_131 N_A_62_94#_c_118_n N_Y_c_412_n 0.014258f $X=1.915 $Y=1.69 $X2=0 $Y2=0
cc_132 N_A_62_94#_c_119_n N_Y_c_412_n 0.0107456f $X=1.645 $Y=1.69 $X2=0 $Y2=0
cc_133 N_A_62_94#_c_127_n N_Y_c_412_n 0.0124932f $X=2.005 $Y=1.765 $X2=0 $Y2=0
cc_134 N_A_62_94#_c_123_n N_Y_c_412_n 0.0153964f $X=0.89 $Y=1.65 $X2=0 $Y2=0
cc_135 N_A_62_94#_c_130_n N_Y_c_412_n 0.00462333f $X=0.81 $Y=1.94 $X2=0 $Y2=0
cc_136 N_A_62_94#_M1011_g N_Y_c_415_n 0.0126976f $X=1.57 $Y=0.74 $X2=0 $Y2=0
cc_137 N_A_62_94#_M1006_g N_Y_c_416_n 5.22898e-19 $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A_62_94#_M1011_g N_Y_c_416_n 0.0124603f $X=1.57 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A_62_94#_c_118_n N_Y_c_416_n 0.00792266f $X=1.915 $Y=1.69 $X2=0 $Y2=0
cc_140 N_A_62_94#_c_119_n N_Y_c_416_n 0.00363407f $X=1.645 $Y=1.69 $X2=0 $Y2=0
cc_141 N_A_62_94#_c_123_n N_Y_c_416_n 0.0113438f $X=0.89 $Y=1.65 $X2=0 $Y2=0
cc_142 N_A_62_94#_c_123_n N_VGND_M1003_d 0.00188126f $X=0.89 $Y=1.65 $X2=-0.19
+ $Y2=-0.245
cc_143 N_A_62_94#_M1006_g N_VGND_c_466_n 0.0113786f $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A_62_94#_M1011_g N_VGND_c_466_n 5.01478e-19 $X=1.57 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A_62_94#_c_120_n N_VGND_c_466_n 0.00121634f $X=0.435 $Y=0.615 $X2=0
+ $Y2=0
cc_146 N_A_62_94#_c_121_n N_VGND_c_466_n 0.00265802f $X=0.805 $Y=1.195 $X2=0
+ $Y2=0
cc_147 N_A_62_94#_c_123_n N_VGND_c_466_n 0.0192874f $X=0.89 $Y=1.65 $X2=0 $Y2=0
cc_148 N_A_62_94#_M1006_g N_VGND_c_467_n 0.00383152f $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A_62_94#_M1011_g N_VGND_c_467_n 0.00383152f $X=1.57 $Y=0.74 $X2=0 $Y2=0
cc_150 N_A_62_94#_M1006_g N_VGND_c_468_n 4.62684e-19 $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_151 N_A_62_94#_M1011_g N_VGND_c_468_n 0.0117356f $X=1.57 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A_62_94#_c_120_n N_VGND_c_470_n 0.00787252f $X=0.435 $Y=0.615 $X2=0
+ $Y2=0
cc_153 N_A_62_94#_M1006_g N_VGND_c_474_n 0.0075754f $X=1.14 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A_62_94#_M1011_g N_VGND_c_474_n 0.0075754f $X=1.57 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A_62_94#_c_120_n N_VGND_c_474_n 0.0085887f $X=0.435 $Y=0.615 $X2=0
+ $Y2=0
cc_156 N_A_62_94#_M1011_g N_A_436_74#_c_525_n 6.92543e-19 $X=1.57 $Y=0.74 $X2=0
+ $Y2=0
cc_157 N_A1_M1005_g N_A2_M1008_g 0.012693f $X=2.905 $Y=2.4 $X2=0 $Y2=0
cc_158 N_A1_c_200_n N_A2_M1008_g 4.48724e-19 $X=2.65 $Y=1.485 $X2=0 $Y2=0
cc_159 N_A1_M1012_g N_A2_c_255_n 0.0123753f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A1_M1012_g A2 0.00134497f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A1_c_200_n A2 0.00804954f $X=2.65 $Y=1.485 $X2=0 $Y2=0
cc_162 N_A1_c_201_n A2 3.7708e-19 $X=2.905 $Y=1.485 $X2=0 $Y2=0
cc_163 N_A1_M1012_g N_A2_c_259_n 0.0135068f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A1_c_200_n N_A2_c_259_n 2.20158e-19 $X=2.65 $Y=1.485 $X2=0 $Y2=0
cc_165 N_A1_c_201_n N_A2_c_259_n 0.012693f $X=2.905 $Y=1.485 $X2=0 $Y2=0
cc_166 N_A1_M1004_g N_VPWR_c_301_n 0.0126906f $X=2.455 $Y=2.4 $X2=0 $Y2=0
cc_167 N_A1_M1005_g N_VPWR_c_301_n 0.0133668f $X=2.905 $Y=2.4 $X2=0 $Y2=0
cc_168 N_A1_M1005_g N_VPWR_c_302_n 5.94799e-19 $X=2.905 $Y=2.4 $X2=0 $Y2=0
cc_169 N_A1_M1004_g N_VPWR_c_303_n 0.00460063f $X=2.455 $Y=2.4 $X2=0 $Y2=0
cc_170 N_A1_M1005_g N_VPWR_c_304_n 0.00460063f $X=2.905 $Y=2.4 $X2=0 $Y2=0
cc_171 N_A1_M1004_g N_VPWR_c_298_n 0.00908665f $X=2.455 $Y=2.4 $X2=0 $Y2=0
cc_172 N_A1_M1005_g N_VPWR_c_298_n 0.00908665f $X=2.905 $Y=2.4 $X2=0 $Y2=0
cc_173 N_A1_M1004_g N_A_241_368#_c_352_n 0.00101073f $X=2.455 $Y=2.4 $X2=0 $Y2=0
cc_174 N_A1_M1004_g N_A_241_368#_c_354_n 4.77247e-19 $X=2.455 $Y=2.4 $X2=0 $Y2=0
cc_175 N_A1_M1004_g N_A_241_368#_c_370_n 0.0177554f $X=2.455 $Y=2.4 $X2=0 $Y2=0
cc_176 N_A1_M1005_g N_A_241_368#_c_370_n 0.0196844f $X=2.905 $Y=2.4 $X2=0 $Y2=0
cc_177 N_A1_c_200_n N_A_241_368#_c_370_n 0.0218744f $X=2.65 $Y=1.485 $X2=0 $Y2=0
cc_178 N_A1_c_201_n N_A_241_368#_c_370_n 4.54857e-19 $X=2.905 $Y=1.485 $X2=0
+ $Y2=0
cc_179 N_A1_M1005_g N_A_241_368#_c_355_n 3.62369e-19 $X=2.905 $Y=2.4 $X2=0 $Y2=0
cc_180 N_A1_M1005_g N_A_241_368#_c_358_n 0.00190277f $X=2.905 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A1_c_200_n N_A_241_368#_c_358_n 0.00384603f $X=2.65 $Y=1.485 $X2=0
+ $Y2=0
cc_182 N_A1_c_200_n N_Y_c_412_n 0.011574f $X=2.65 $Y=1.485 $X2=0 $Y2=0
cc_183 N_A1_c_201_n N_Y_c_412_n 0.00299935f $X=2.905 $Y=1.485 $X2=0 $Y2=0
cc_184 N_A1_M1000_g N_Y_c_413_n 0.0126181f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_185 N_A1_c_200_n N_Y_c_413_n 0.00619439f $X=2.65 $Y=1.485 $X2=0 $Y2=0
cc_186 N_A1_c_201_n N_Y_c_413_n 0.0033205f $X=2.905 $Y=1.485 $X2=0 $Y2=0
cc_187 N_A1_M1000_g N_Y_c_414_n 0.0103649f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_188 N_A1_M1012_g N_Y_c_414_n 0.00672659f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A1_c_200_n N_Y_c_414_n 0.0200194f $X=2.65 $Y=1.485 $X2=0 $Y2=0
cc_190 N_A1_c_201_n N_Y_c_414_n 7.44695e-19 $X=2.905 $Y=1.485 $X2=0 $Y2=0
cc_191 N_A1_M1000_g N_Y_c_416_n 0.00689063f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A1_c_200_n N_Y_c_416_n 0.00638885f $X=2.65 $Y=1.485 $X2=0 $Y2=0
cc_193 N_A1_c_201_n N_Y_c_416_n 0.00143746f $X=2.905 $Y=1.485 $X2=0 $Y2=0
cc_194 N_A1_M1000_g N_VGND_c_468_n 0.00714008f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A1_M1012_g N_VGND_c_469_n 6.35276e-19 $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A1_M1000_g N_VGND_c_472_n 0.00291649f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A1_M1012_g N_VGND_c_472_n 0.00291649f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_198 N_A1_M1000_g N_VGND_c_474_n 0.0036412f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A1_M1012_g N_VGND_c_474_n 0.00359219f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A1_M1000_g N_A_436_74#_c_525_n 0.01124f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_201 N_A1_M1012_g N_A_436_74#_c_525_n 0.0142063f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_202 N_A2_M1008_g N_VPWR_c_301_n 5.41206e-19 $X=3.355 $Y=2.4 $X2=0 $Y2=0
cc_203 N_A2_M1008_g N_VPWR_c_302_n 0.0156093f $X=3.355 $Y=2.4 $X2=0 $Y2=0
cc_204 N_A2_M1009_g N_VPWR_c_302_n 0.0188964f $X=3.825 $Y=2.4 $X2=0 $Y2=0
cc_205 N_A2_M1008_g N_VPWR_c_304_n 0.00460063f $X=3.355 $Y=2.4 $X2=0 $Y2=0
cc_206 N_A2_M1009_g N_VPWR_c_305_n 0.00460063f $X=3.825 $Y=2.4 $X2=0 $Y2=0
cc_207 N_A2_M1008_g N_VPWR_c_298_n 0.00908665f $X=3.355 $Y=2.4 $X2=0 $Y2=0
cc_208 N_A2_M1009_g N_VPWR_c_298_n 0.00912261f $X=3.825 $Y=2.4 $X2=0 $Y2=0
cc_209 N_A2_M1008_g N_A_241_368#_c_355_n 3.62369e-19 $X=3.355 $Y=2.4 $X2=0 $Y2=0
cc_210 N_A2_M1008_g N_A_241_368#_c_356_n 0.0149087f $X=3.355 $Y=2.4 $X2=0 $Y2=0
cc_211 N_A2_M1009_g N_A_241_368#_c_356_n 0.0221599f $X=3.825 $Y=2.4 $X2=0 $Y2=0
cc_212 A2 N_A_241_368#_c_356_n 0.0334689f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_213 N_A2_c_259_n N_A_241_368#_c_356_n 7.74501e-19 $X=3.825 $Y=1.385 $X2=0
+ $Y2=0
cc_214 N_A2_M1009_g N_A_241_368#_c_357_n 0.00147311f $X=3.825 $Y=2.4 $X2=0 $Y2=0
cc_215 N_A2_M1008_g N_A_241_368#_c_358_n 2.3892e-19 $X=3.355 $Y=2.4 $X2=0 $Y2=0
cc_216 N_A2_c_255_n N_Y_c_414_n 4.34981e-19 $X=3.38 $Y=1.22 $X2=0 $Y2=0
cc_217 N_A2_c_255_n N_VGND_c_469_n 0.00768902f $X=3.38 $Y=1.22 $X2=0 $Y2=0
cc_218 N_A2_c_256_n N_VGND_c_469_n 0.010528f $X=3.81 $Y=1.22 $X2=0 $Y2=0
cc_219 N_A2_c_255_n N_VGND_c_472_n 0.00383152f $X=3.38 $Y=1.22 $X2=0 $Y2=0
cc_220 N_A2_c_256_n N_VGND_c_473_n 0.00383152f $X=3.81 $Y=1.22 $X2=0 $Y2=0
cc_221 N_A2_c_255_n N_VGND_c_474_n 0.00384065f $X=3.38 $Y=1.22 $X2=0 $Y2=0
cc_222 N_A2_c_256_n N_VGND_c_474_n 0.00387675f $X=3.81 $Y=1.22 $X2=0 $Y2=0
cc_223 N_A2_c_255_n N_A_436_74#_c_532_n 0.00985057f $X=3.38 $Y=1.22 $X2=0 $Y2=0
cc_224 N_A2_c_256_n N_A_436_74#_c_532_n 0.0141214f $X=3.81 $Y=1.22 $X2=0 $Y2=0
cc_225 A2 N_A_436_74#_c_532_n 0.0271317f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_226 N_A2_c_259_n N_A_436_74#_c_532_n 6.30401e-19 $X=3.825 $Y=1.385 $X2=0
+ $Y2=0
cc_227 N_A2_c_256_n N_A_436_74#_c_527_n 7.92899e-19 $X=3.81 $Y=1.22 $X2=0 $Y2=0
cc_228 N_A2_c_256_n N_A_436_74#_c_528_n 0.00159319f $X=3.81 $Y=1.22 $X2=0 $Y2=0
cc_229 N_VPWR_c_301_n N_A_241_368#_c_352_n 0.0103602f $X=2.68 $Y=2.375 $X2=0
+ $Y2=0
cc_230 N_VPWR_c_303_n N_A_241_368#_c_352_n 0.0583239f $X=2.515 $Y=3.33 $X2=0
+ $Y2=0
cc_231 N_VPWR_c_298_n N_A_241_368#_c_352_n 0.0324477f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_232 N_VPWR_c_303_n N_A_241_368#_c_353_n 0.0179217f $X=2.515 $Y=3.33 $X2=0
+ $Y2=0
cc_233 N_VPWR_c_298_n N_A_241_368#_c_353_n 0.00971942f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_234 N_VPWR_M1004_d N_A_241_368#_c_370_n 0.0031498f $X=2.545 $Y=1.84 $X2=0
+ $Y2=0
cc_235 N_VPWR_c_301_n N_A_241_368#_c_370_n 0.0170259f $X=2.68 $Y=2.375 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_301_n N_A_241_368#_c_355_n 0.0233699f $X=2.68 $Y=2.375 $X2=0
+ $Y2=0
cc_237 N_VPWR_c_302_n N_A_241_368#_c_355_n 0.0312215f $X=3.59 $Y=2.145 $X2=0
+ $Y2=0
cc_238 N_VPWR_c_304_n N_A_241_368#_c_355_n 0.00749631f $X=3.415 $Y=3.33 $X2=0
+ $Y2=0
cc_239 N_VPWR_c_298_n N_A_241_368#_c_355_n 0.0062048f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_240 N_VPWR_M1008_d N_A_241_368#_c_356_n 0.00187091f $X=3.445 $Y=1.84 $X2=0
+ $Y2=0
cc_241 N_VPWR_c_302_n N_A_241_368#_c_356_n 0.018653f $X=3.59 $Y=2.145 $X2=0
+ $Y2=0
cc_242 N_VPWR_c_302_n N_A_241_368#_c_357_n 0.03126f $X=3.59 $Y=2.145 $X2=0 $Y2=0
cc_243 N_VPWR_c_305_n N_A_241_368#_c_357_n 0.011066f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_244 N_VPWR_c_298_n N_A_241_368#_c_357_n 0.00915947f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_245 N_A_241_368#_c_352_n N_Y_M1001_d 0.00165831f $X=2.115 $Y=2.99 $X2=0 $Y2=0
cc_246 N_A_241_368#_c_351_n N_Y_c_411_n 6.70242e-19 $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_247 N_A_241_368#_c_351_n N_Y_c_412_n 0.030821f $X=1.33 $Y=1.985 $X2=0 $Y2=0
cc_248 N_A_241_368#_c_352_n N_Y_c_412_n 0.0159318f $X=2.115 $Y=2.99 $X2=0 $Y2=0
cc_249 N_A_241_368#_c_354_n N_Y_c_412_n 0.0120471f $X=2.215 $Y=2.12 $X2=0 $Y2=0
cc_250 N_A_241_368#_c_354_n N_Y_c_413_n 0.00127772f $X=2.215 $Y=2.12 $X2=0 $Y2=0
cc_251 N_A_241_368#_c_354_n N_Y_c_416_n 0.00783425f $X=2.215 $Y=2.12 $X2=0 $Y2=0
cc_252 N_A_241_368#_c_356_n N_A_436_74#_c_538_n 0.00103389f $X=3.965 $Y=1.805
+ $X2=0 $Y2=0
cc_253 N_A_241_368#_c_358_n N_A_436_74#_c_538_n 0.00450741f $X=3.13 $Y=1.805
+ $X2=0 $Y2=0
cc_254 N_A_241_368#_c_356_n N_A_436_74#_c_527_n 0.00969915f $X=3.965 $Y=1.805
+ $X2=0 $Y2=0
cc_255 N_Y_c_416_n N_VGND_M1011_s 0.00288199f $X=2.275 $Y=1.195 $X2=0 $Y2=0
cc_256 N_Y_c_410_n N_VGND_c_466_n 0.0218329f $X=1.355 $Y=0.515 $X2=0 $Y2=0
cc_257 N_Y_c_410_n N_VGND_c_467_n 0.00749631f $X=1.355 $Y=0.515 $X2=0 $Y2=0
cc_258 N_Y_c_410_n N_VGND_c_468_n 0.0171736f $X=1.355 $Y=0.515 $X2=0 $Y2=0
cc_259 N_Y_c_414_n N_VGND_c_468_n 0.0011882f $X=2.735 $Y=0.91 $X2=0 $Y2=0
cc_260 N_Y_c_416_n N_VGND_c_468_n 0.023479f $X=2.275 $Y=1.195 $X2=0 $Y2=0
cc_261 N_Y_c_410_n N_VGND_c_474_n 0.0062048f $X=1.355 $Y=0.515 $X2=0 $Y2=0
cc_262 N_Y_c_413_n N_A_436_74#_M1000_d 0.00174919f $X=2.57 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_263 N_Y_c_416_n N_A_436_74#_M1000_d 0.00213669f $X=2.275 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_264 N_Y_M1000_s N_A_436_74#_c_525_n 0.00178571f $X=2.595 $Y=0.37 $X2=0 $Y2=0
cc_265 N_Y_c_414_n N_A_436_74#_c_525_n 0.0162079f $X=2.735 $Y=0.91 $X2=0 $Y2=0
cc_266 N_Y_c_416_n N_A_436_74#_c_525_n 0.0153378f $X=2.275 $Y=1.195 $X2=0 $Y2=0
cc_267 N_VGND_c_468_n N_A_436_74#_c_525_n 0.0202776f $X=1.785 $Y=0.645 $X2=0
+ $Y2=0
cc_268 N_VGND_c_472_n N_A_436_74#_c_525_n 0.038121f $X=3.43 $Y=0 $X2=0 $Y2=0
cc_269 N_VGND_c_474_n N_A_436_74#_c_525_n 0.0321651f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_270 N_VGND_c_469_n N_A_436_74#_c_526_n 0.00985092f $X=3.595 $Y=0.55 $X2=0
+ $Y2=0
cc_271 N_VGND_c_472_n N_A_436_74#_c_526_n 0.00760167f $X=3.43 $Y=0 $X2=0 $Y2=0
cc_272 N_VGND_c_474_n N_A_436_74#_c_526_n 0.00628491f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_273 N_VGND_M1007_d N_A_436_74#_c_532_n 0.00328934f $X=3.455 $Y=0.37 $X2=0
+ $Y2=0
cc_274 N_VGND_c_469_n N_A_436_74#_c_532_n 0.0167019f $X=3.595 $Y=0.55 $X2=0
+ $Y2=0
cc_275 N_VGND_c_474_n N_A_436_74#_c_532_n 0.0116543f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_276 N_VGND_c_469_n N_A_436_74#_c_528_n 0.0121972f $X=3.595 $Y=0.55 $X2=0
+ $Y2=0
cc_277 N_VGND_c_473_n N_A_436_74#_c_528_n 0.011066f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_278 N_VGND_c_474_n N_A_436_74#_c_528_n 0.00915947f $X=4.08 $Y=0 $X2=0 $Y2=0

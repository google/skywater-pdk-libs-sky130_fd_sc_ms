* File: sky130_fd_sc_ms__o2bb2ai_4.pxi.spice
* Created: Wed Sep  2 12:24:42 2020
* 
x_PM_SKY130_FD_SC_MS__O2BB2AI_4%A1_N N_A1_N_M1026_g N_A1_N_M1012_g
+ N_A1_N_M1032_g N_A1_N_M1027_g N_A1_N_M1033_g N_A1_N_M1030_g N_A1_N_M1034_g
+ N_A1_N_M1036_g A1_N A1_N A1_N A1_N N_A1_N_c_175_n N_A1_N_c_176_n
+ PM_SKY130_FD_SC_MS__O2BB2AI_4%A1_N
x_PM_SKY130_FD_SC_MS__O2BB2AI_4%A2_N N_A2_N_M1008_g N_A2_N_M1000_g
+ N_A2_N_M1017_g N_A2_N_M1003_g N_A2_N_M1022_g N_A2_N_M1005_g N_A2_N_c_258_n
+ N_A2_N_M1010_g N_A2_N_M1039_g N_A2_N_c_261_n A2_N A2_N N_A2_N_c_262_n
+ PM_SKY130_FD_SC_MS__O2BB2AI_4%A2_N
x_PM_SKY130_FD_SC_MS__O2BB2AI_4%A_117_368# N_A_117_368#_M1008_s
+ N_A_117_368#_M1022_s N_A_117_368#_M1026_d N_A_117_368#_M1030_d
+ N_A_117_368#_M1000_d N_A_117_368#_M1005_d N_A_117_368#_M1014_g
+ N_A_117_368#_M1019_g N_A_117_368#_M1009_g N_A_117_368#_M1021_g
+ N_A_117_368#_M1018_g N_A_117_368#_M1028_g N_A_117_368#_M1023_g
+ N_A_117_368#_c_359_n N_A_117_368#_c_360_n N_A_117_368#_M1029_g
+ N_A_117_368#_c_375_n N_A_117_368#_c_370_n N_A_117_368#_c_382_n
+ N_A_117_368#_c_371_n N_A_117_368#_c_389_n N_A_117_368#_c_402_n
+ N_A_117_368#_c_372_n N_A_117_368#_c_362_n N_A_117_368#_c_363_n
+ N_A_117_368#_c_416_n N_A_117_368#_c_373_n N_A_117_368#_c_423_n
+ N_A_117_368#_c_364_n N_A_117_368#_c_374_n N_A_117_368#_c_365_n
+ N_A_117_368#_c_392_n N_A_117_368#_c_437_n N_A_117_368#_c_441_n
+ PM_SKY130_FD_SC_MS__O2BB2AI_4%A_117_368#
x_PM_SKY130_FD_SC_MS__O2BB2AI_4%B2 N_B2_M1002_g N_B2_M1001_g N_B2_M1024_g
+ N_B2_M1004_g N_B2_M1025_g N_B2_M1031_g N_B2_M1037_g N_B2_M1038_g B2 B2 B2 B2
+ N_B2_c_563_n N_B2_c_564_n PM_SKY130_FD_SC_MS__O2BB2AI_4%B2
x_PM_SKY130_FD_SC_MS__O2BB2AI_4%B1 N_B1_M1007_g N_B1_M1006_g N_B1_M1013_g
+ N_B1_M1011_g N_B1_M1016_g N_B1_M1015_g N_B1_M1020_g N_B1_M1035_g B1 B1 B1 B1
+ N_B1_c_654_n PM_SKY130_FD_SC_MS__O2BB2AI_4%B1
x_PM_SKY130_FD_SC_MS__O2BB2AI_4%VPWR N_VPWR_M1026_s N_VPWR_M1027_s
+ N_VPWR_M1036_s N_VPWR_M1003_s N_VPWR_M1010_s N_VPWR_M1019_s N_VPWR_M1028_s
+ N_VPWR_M1007_d N_VPWR_M1015_d N_VPWR_c_731_n N_VPWR_c_732_n N_VPWR_c_733_n
+ N_VPWR_c_734_n N_VPWR_c_735_n N_VPWR_c_736_n N_VPWR_c_737_n N_VPWR_c_738_n
+ N_VPWR_c_739_n N_VPWR_c_740_n N_VPWR_c_741_n N_VPWR_c_742_n N_VPWR_c_743_n
+ N_VPWR_c_744_n N_VPWR_c_745_n N_VPWR_c_746_n N_VPWR_c_747_n N_VPWR_c_748_n
+ N_VPWR_c_749_n N_VPWR_c_750_n N_VPWR_c_751_n VPWR N_VPWR_c_752_n
+ N_VPWR_c_753_n N_VPWR_c_754_n N_VPWR_c_730_n N_VPWR_c_756_n N_VPWR_c_757_n
+ N_VPWR_c_758_n PM_SKY130_FD_SC_MS__O2BB2AI_4%VPWR
x_PM_SKY130_FD_SC_MS__O2BB2AI_4%Y N_Y_M1009_s N_Y_M1023_s N_Y_M1014_d
+ N_Y_M1021_d N_Y_M1001_d N_Y_M1031_d N_Y_c_884_n N_Y_c_885_n N_Y_c_886_n
+ N_Y_c_903_n N_Y_c_880_n N_Y_c_881_n N_Y_c_887_n N_Y_c_916_n N_Y_c_882_n
+ N_Y_c_889_n N_Y_c_890_n N_Y_c_940_n N_Y_c_883_n N_Y_c_944_n N_Y_c_949_n Y
+ PM_SKY130_FD_SC_MS__O2BB2AI_4%Y
x_PM_SKY130_FD_SC_MS__O2BB2AI_4%A_1215_368# N_A_1215_368#_M1001_s
+ N_A_1215_368#_M1004_s N_A_1215_368#_M1037_s N_A_1215_368#_M1011_s
+ N_A_1215_368#_M1020_s N_A_1215_368#_c_988_n N_A_1215_368#_c_989_n
+ N_A_1215_368#_c_990_n N_A_1215_368#_c_1051_n N_A_1215_368#_c_991_n
+ N_A_1215_368#_c_1003_n N_A_1215_368#_c_992_n N_A_1215_368#_c_1011_n
+ N_A_1215_368#_c_993_n N_A_1215_368#_c_994_n N_A_1215_368#_c_995_n
+ N_A_1215_368#_c_1020_n PM_SKY130_FD_SC_MS__O2BB2AI_4%A_1215_368#
x_PM_SKY130_FD_SC_MS__O2BB2AI_4%A_27_74# N_A_27_74#_M1012_d N_A_27_74#_M1032_d
+ N_A_27_74#_M1034_d N_A_27_74#_M1017_d N_A_27_74#_M1039_d N_A_27_74#_c_1054_n
+ N_A_27_74#_c_1055_n N_A_27_74#_c_1056_n N_A_27_74#_c_1057_n
+ N_A_27_74#_c_1058_n N_A_27_74#_c_1059_n N_A_27_74#_c_1060_n
+ N_A_27_74#_c_1093_n N_A_27_74#_c_1061_n N_A_27_74#_c_1062_n
+ N_A_27_74#_c_1063_n N_A_27_74#_c_1064_n PM_SKY130_FD_SC_MS__O2BB2AI_4%A_27_74#
x_PM_SKY130_FD_SC_MS__O2BB2AI_4%VGND N_VGND_M1012_s N_VGND_M1033_s
+ N_VGND_M1002_d N_VGND_M1025_d N_VGND_M1006_s N_VGND_M1016_s N_VGND_c_1122_n
+ N_VGND_c_1123_n N_VGND_c_1124_n N_VGND_c_1125_n N_VGND_c_1126_n
+ N_VGND_c_1127_n N_VGND_c_1128_n VGND N_VGND_c_1129_n N_VGND_c_1130_n
+ N_VGND_c_1131_n N_VGND_c_1132_n N_VGND_c_1133_n N_VGND_c_1134_n
+ N_VGND_c_1135_n N_VGND_c_1136_n N_VGND_c_1137_n N_VGND_c_1138_n
+ N_VGND_c_1139_n N_VGND_c_1140_n N_VGND_c_1141_n
+ PM_SKY130_FD_SC_MS__O2BB2AI_4%VGND
x_PM_SKY130_FD_SC_MS__O2BB2AI_4%A_857_74# N_A_857_74#_M1009_d
+ N_A_857_74#_M1018_d N_A_857_74#_M1029_d N_A_857_74#_M1024_s
+ N_A_857_74#_M1038_s N_A_857_74#_M1013_d N_A_857_74#_M1035_d
+ N_A_857_74#_c_1251_n N_A_857_74#_c_1252_n N_A_857_74#_c_1253_n
+ N_A_857_74#_c_1318_n N_A_857_74#_c_1254_n N_A_857_74#_c_1255_n
+ N_A_857_74#_c_1256_n N_A_857_74#_c_1257_n N_A_857_74#_c_1258_n
+ N_A_857_74#_c_1259_n N_A_857_74#_c_1260_n N_A_857_74#_c_1261_n
+ N_A_857_74#_c_1262_n N_A_857_74#_c_1263_n N_A_857_74#_c_1264_n
+ N_A_857_74#_c_1265_n N_A_857_74#_c_1266_n N_A_857_74#_c_1267_n
+ PM_SKY130_FD_SC_MS__O2BB2AI_4%A_857_74#
cc_1 VNB N_A1_N_M1012_g 0.0318708f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A1_N_M1032_g 0.0226407f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_3 VNB N_A1_N_M1033_g 0.0226407f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.74
cc_4 VNB N_A1_N_M1034_g 0.0229726f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.74
cc_5 VNB N_A1_N_c_175_n 0.0160224f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.515
cc_6 VNB N_A1_N_c_176_n 0.0812712f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.515
cc_7 VNB N_A2_N_M1008_g 0.0213573f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_8 VNB N_A2_N_M1017_g 0.0218695f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_9 VNB N_A2_N_M1022_g 0.0224304f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.74
cc_10 VNB N_A2_N_c_258_n 0.0106061f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.35
cc_11 VNB N_A2_N_M1010_g 0.00459789f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.68
cc_12 VNB N_A2_N_M1039_g 0.0282424f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_13 VNB N_A2_N_c_261_n 0.00935952f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_14 VNB N_A2_N_c_262_n 0.0574705f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.515
cc_15 VNB N_A_117_368#_M1014_g 0.00159413f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=1.68
cc_16 VNB N_A_117_368#_M1019_g 0.00154301f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.35
cc_17 VNB N_A_117_368#_M1009_g 0.027434f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=1.68
cc_18 VNB N_A_117_368#_M1021_g 0.00154166f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_19 VNB N_A_117_368#_M1018_g 0.0200535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_117_368#_M1028_g 0.00167336f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=1.515
cc_21 VNB N_A_117_368#_M1023_g 0.0193643f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_22 VNB N_A_117_368#_c_359_n 0.0243374f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.515
cc_23 VNB N_A_117_368#_c_360_n 0.0979322f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=1.515
cc_24 VNB N_A_117_368#_M1029_g 0.020471f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.515
cc_25 VNB N_A_117_368#_c_362_n 0.00349695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_117_368#_c_363_n 0.00229069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_117_368#_c_364_n 0.00589432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_117_368#_c_365_n 0.0113354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B2_M1002_g 0.0239651f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_30 VNB N_B2_M1024_g 0.0240453f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_31 VNB N_B2_M1025_g 0.0234895f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.74
cc_32 VNB N_B2_M1038_g 0.0245189f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_33 VNB N_B2_c_563_n 0.00585801f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.515
cc_34 VNB N_B2_c_564_n 0.0759749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_B1_M1006_g 0.0230003f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_36 VNB N_B1_M1013_g 0.0224928f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_37 VNB N_B1_M1016_g 0.0240453f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.74
cc_38 VNB N_B1_M1035_g 0.0328675f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_39 VNB B1 0.0153948f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_40 VNB N_B1_c_654_n 0.0831493f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.515
cc_41 VNB N_VPWR_c_730_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_Y_c_880_n 0.00258452f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_43 VNB N_Y_c_881_n 0.00229484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_Y_c_882_n 0.00349117f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=1.515
cc_45 VNB N_Y_c_883_n 0.00416741f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.515
cc_46 VNB N_A_27_74#_c_1054_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.74
cc_47 VNB N_A_27_74#_c_1055_n 0.00307486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_27_74#_c_1056_n 0.00955057f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=1.68
cc_49 VNB N_A_27_74#_c_1057_n 0.00188248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_27_74#_c_1058_n 0.0101688f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.74
cc_51 VNB N_A_27_74#_c_1059_n 0.0026914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_27_74#_c_1060_n 0.00211517f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_53 VNB N_A_27_74#_c_1061_n 0.00647211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_27_74#_c_1062_n 0.00865153f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=1.515
cc_55 VNB N_A_27_74#_c_1063_n 0.00133271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_27_74#_c_1064_n 0.00244965f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_57 VNB N_VGND_c_1122_n 0.00324953f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=1.68
cc_58 VNB N_VGND_c_1123_n 0.00324953f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.35
cc_59 VNB N_VGND_c_1124_n 0.108794f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.74
cc_60 VNB N_VGND_c_1125_n 0.00558127f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.4
cc_61 VNB N_VGND_c_1126_n 0.00494723f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_62 VNB N_VGND_c_1127_n 0.00269659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1128_n 0.00558127f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=1.515
cc_64 VNB N_VGND_c_1129_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.515
cc_65 VNB N_VGND_c_1130_n 0.0154137f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.515
cc_66 VNB N_VGND_c_1131_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1132_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_68 VNB N_VGND_c_1133_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1134_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1135_n 0.534813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1136_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1137_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1138_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1139_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1140_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1141_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_857_74#_c_1251_n 0.00792168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_857_74#_c_1252_n 0.0027626f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.74
cc_79 VNB N_A_857_74#_c_1253_n 0.00377359f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.74
cc_80 VNB N_A_857_74#_c_1254_n 0.00487777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_857_74#_c_1255_n 0.00317099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_857_74#_c_1256_n 0.00219196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_857_74#_c_1257_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.41 $Y2=1.515
cc_84 VNB N_A_857_74#_c_1258_n 0.00518435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_857_74#_c_1259_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=1.365
+ $Y2=1.515
cc_86 VNB N_A_857_74#_c_1260_n 0.00448959f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.515
cc_87 VNB N_A_857_74#_c_1261_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=1.845
+ $Y2=1.515
cc_88 VNB N_A_857_74#_c_1262_n 0.0125337f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_89 VNB N_A_857_74#_c_1263_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_90 VNB N_A_857_74#_c_1264_n 0.00121798f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_91 VNB N_A_857_74#_c_1265_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_857_74#_c_1266_n 0.0090169f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.565
cc_93 VNB N_A_857_74#_c_1267_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VPB N_A1_N_M1026_g 0.0246451f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_95 VPB N_A1_N_M1027_g 0.020498f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_96 VPB N_A1_N_M1030_g 0.020498f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_97 VPB N_A1_N_M1036_g 0.0208438f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_98 VPB N_A1_N_c_175_n 0.017403f $X=-0.19 $Y=1.66 $X2=1.77 $Y2=1.515
cc_99 VPB N_A1_N_c_176_n 0.0166563f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.515
cc_100 VPB N_A2_N_M1000_g 0.0214106f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_101 VPB N_A2_N_M1003_g 0.0204968f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_102 VPB N_A2_N_M1005_g 0.0208684f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_103 VPB N_A2_N_M1010_g 0.0222147f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.68
cc_104 VPB A2_N 0.00503583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A2_N_c_262_n 0.00976784f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.515
cc_106 VPB N_A_117_368#_M1014_g 0.0227918f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.68
cc_107 VPB N_A_117_368#_M1019_g 0.0220607f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.35
cc_108 VPB N_A_117_368#_M1021_g 0.0220515f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_109 VPB N_A_117_368#_M1028_g 0.0247319f $X=-0.19 $Y=1.66 $X2=0.41 $Y2=1.515
cc_110 VPB N_A_117_368#_c_370_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_117_368#_c_371_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_117_368#_c_372_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_117_368#_c_373_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_117_368#_c_374_n 0.00128541f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_B2_M1001_g 0.0240703f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_116 VPB N_B2_M1004_g 0.0196385f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_117 VPB N_B2_M1031_g 0.0196385f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_118 VPB N_B2_M1037_g 0.0207362f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=0.74
cc_119 VPB N_B2_c_563_n 0.0139997f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.515
cc_120 VPB N_B2_c_564_n 0.0136118f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_B1_M1007_g 0.0207956f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_122 VPB N_B1_M1011_g 0.0204971f $X=-0.19 $Y=1.66 $X2=0.945 $Y2=2.4
cc_123 VPB N_B1_M1015_g 0.0204971f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=2.4
cc_124 VPB N_B1_M1020_g 0.0275823f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=0.74
cc_125 VPB B1 0.0150114f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_126 VPB N_B1_c_654_n 0.0169943f $X=-0.19 $Y=1.66 $X2=1.77 $Y2=1.515
cc_127 VPB N_VPWR_c_731_n 0.0103331f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_732_n 0.0506396f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=2.4
cc_129 VPB N_VPWR_c_733_n 0.00797179f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_130 VPB N_VPWR_c_734_n 0.00797179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_735_n 0.00797179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_736_n 0.00996599f $X=-0.19 $Y=1.66 $X2=1.365 $Y2=1.515
cc_133 VPB N_VPWR_c_737_n 0.00732691f $X=-0.19 $Y=1.66 $X2=1.845 $Y2=1.515
cc_134 VPB N_VPWR_c_738_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_135 VPB N_VPWR_c_739_n 0.0116901f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_136 VPB N_VPWR_c_740_n 0.00570462f $X=-0.19 $Y=1.66 $X2=1.68 $Y2=1.565
cc_137 VPB N_VPWR_c_741_n 0.00837583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_742_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_743_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_744_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_745_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_746_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_747_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_748_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_749_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_750_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_751_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_752_n 0.0581001f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_753_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_754_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_730_n 0.109455f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_756_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_757_n 0.00487714f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_758_n 0.00391723f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_Y_c_884_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.68
cc_156 VPB N_Y_c_885_n 0.00219429f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.35
cc_157 VPB N_Y_c_886_n 0.00224287f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=0.74
cc_158 VPB N_Y_c_887_n 0.00202354f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_159 VPB N_Y_c_882_n 0.00243906f $X=-0.19 $Y=1.66 $X2=0.41 $Y2=1.515
cc_160 VPB N_Y_c_889_n 0.0120271f $X=-0.19 $Y=1.66 $X2=0.41 $Y2=1.515
cc_161 VPB N_Y_c_890_n 0.00300835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_A_1215_368#_c_988_n 0.00587698f $X=-0.19 $Y=1.66 $X2=1.365 $Y2=0.74
cc_163 VPB N_A_1215_368#_c_989_n 0.00240659f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_1215_368#_c_990_n 0.00384043f $X=-0.19 $Y=1.66 $X2=1.395 $Y2=1.68
cc_165 VPB N_A_1215_368#_c_991_n 0.00478582f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=0.74
cc_166 VPB N_A_1215_368#_c_992_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_167 VPB N_A_1215_368#_c_993_n 0.00802076f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_1215_368#_c_994_n 0.0355666f $X=-0.19 $Y=1.66 $X2=0.41 $Y2=1.515
cc_169 VPB N_A_1215_368#_c_995_n 0.00145593f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 N_A1_N_M1034_g N_A2_N_M1008_g 0.0189918f $X=1.795 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A1_N_M1036_g N_A2_N_M1000_g 0.0327168f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_172 N_A1_N_c_175_n N_A2_N_M1000_g 3.39254e-19 $X=1.77 $Y=1.515 $X2=0 $Y2=0
cc_173 N_A1_N_c_175_n A2_N 0.0234915f $X=1.77 $Y=1.515 $X2=0 $Y2=0
cc_174 N_A1_N_c_176_n A2_N 4.87369e-19 $X=1.845 $Y=1.515 $X2=0 $Y2=0
cc_175 N_A1_N_c_175_n N_A2_N_c_262_n 0.00140344f $X=1.77 $Y=1.515 $X2=0 $Y2=0
cc_176 N_A1_N_c_176_n N_A2_N_c_262_n 0.0214891f $X=1.845 $Y=1.515 $X2=0 $Y2=0
cc_177 N_A1_N_M1026_g N_A_117_368#_c_375_n 0.0025567f $X=0.495 $Y=2.4 $X2=0
+ $Y2=0
cc_178 N_A1_N_M1027_g N_A_117_368#_c_375_n 8.84614e-19 $X=0.945 $Y=2.4 $X2=0
+ $Y2=0
cc_179 N_A1_N_c_175_n N_A_117_368#_c_375_n 0.0235495f $X=1.77 $Y=1.515 $X2=0
+ $Y2=0
cc_180 N_A1_N_c_176_n N_A_117_368#_c_375_n 5.54423e-19 $X=1.845 $Y=1.515 $X2=0
+ $Y2=0
cc_181 N_A1_N_M1026_g N_A_117_368#_c_370_n 0.0114394f $X=0.495 $Y=2.4 $X2=0
+ $Y2=0
cc_182 N_A1_N_M1027_g N_A_117_368#_c_370_n 0.0121132f $X=0.945 $Y=2.4 $X2=0
+ $Y2=0
cc_183 N_A1_N_M1030_g N_A_117_368#_c_370_n 6.50516e-19 $X=1.395 $Y=2.4 $X2=0
+ $Y2=0
cc_184 N_A1_N_M1027_g N_A_117_368#_c_382_n 0.012931f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_185 N_A1_N_M1030_g N_A_117_368#_c_382_n 0.012931f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_186 N_A1_N_c_175_n N_A_117_368#_c_382_n 0.0391869f $X=1.77 $Y=1.515 $X2=0
+ $Y2=0
cc_187 N_A1_N_c_176_n N_A_117_368#_c_382_n 4.89709e-19 $X=1.845 $Y=1.515 $X2=0
+ $Y2=0
cc_188 N_A1_N_M1027_g N_A_117_368#_c_371_n 6.50516e-19 $X=0.945 $Y=2.4 $X2=0
+ $Y2=0
cc_189 N_A1_N_M1030_g N_A_117_368#_c_371_n 0.0121132f $X=1.395 $Y=2.4 $X2=0
+ $Y2=0
cc_190 N_A1_N_M1036_g N_A_117_368#_c_371_n 0.0121132f $X=1.845 $Y=2.4 $X2=0
+ $Y2=0
cc_191 N_A1_N_M1036_g N_A_117_368#_c_389_n 0.0128923f $X=1.845 $Y=2.4 $X2=0
+ $Y2=0
cc_192 N_A1_N_c_175_n N_A_117_368#_c_389_n 0.0109106f $X=1.77 $Y=1.515 $X2=0
+ $Y2=0
cc_193 N_A1_N_M1036_g N_A_117_368#_c_372_n 6.50516e-19 $X=1.845 $Y=2.4 $X2=0
+ $Y2=0
cc_194 N_A1_N_M1030_g N_A_117_368#_c_392_n 8.84614e-19 $X=1.395 $Y=2.4 $X2=0
+ $Y2=0
cc_195 N_A1_N_M1036_g N_A_117_368#_c_392_n 8.84614e-19 $X=1.845 $Y=2.4 $X2=0
+ $Y2=0
cc_196 N_A1_N_c_175_n N_A_117_368#_c_392_n 0.0235495f $X=1.77 $Y=1.515 $X2=0
+ $Y2=0
cc_197 N_A1_N_c_176_n N_A_117_368#_c_392_n 5.52302e-19 $X=1.845 $Y=1.515 $X2=0
+ $Y2=0
cc_198 N_A1_N_M1026_g N_VPWR_c_732_n 0.00501904f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_199 N_A1_N_c_175_n N_VPWR_c_732_n 0.0199914f $X=1.77 $Y=1.515 $X2=0 $Y2=0
cc_200 N_A1_N_c_176_n N_VPWR_c_732_n 6.56847e-19 $X=1.845 $Y=1.515 $X2=0 $Y2=0
cc_201 N_A1_N_M1027_g N_VPWR_c_733_n 0.0027763f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_202 N_A1_N_M1030_g N_VPWR_c_733_n 0.0027763f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_203 N_A1_N_M1036_g N_VPWR_c_734_n 0.0027763f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_204 N_A1_N_M1026_g N_VPWR_c_742_n 0.005209f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_205 N_A1_N_M1027_g N_VPWR_c_742_n 0.005209f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_206 N_A1_N_M1030_g N_VPWR_c_744_n 0.005209f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_207 N_A1_N_M1036_g N_VPWR_c_744_n 0.005209f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_208 N_A1_N_M1026_g N_VPWR_c_730_n 0.00985972f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_209 N_A1_N_M1027_g N_VPWR_c_730_n 0.00982266f $X=0.945 $Y=2.4 $X2=0 $Y2=0
cc_210 N_A1_N_M1030_g N_VPWR_c_730_n 0.00982266f $X=1.395 $Y=2.4 $X2=0 $Y2=0
cc_211 N_A1_N_M1036_g N_VPWR_c_730_n 0.00982376f $X=1.845 $Y=2.4 $X2=0 $Y2=0
cc_212 N_A1_N_M1012_g N_A_27_74#_c_1054_n 0.00159319f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_213 N_A1_N_M1012_g N_A_27_74#_c_1055_n 0.0136535f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_214 N_A1_N_M1032_g N_A_27_74#_c_1055_n 0.0131164f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_215 N_A1_N_c_175_n N_A_27_74#_c_1055_n 0.0517333f $X=1.77 $Y=1.515 $X2=0
+ $Y2=0
cc_216 N_A1_N_c_176_n N_A_27_74#_c_1055_n 0.00359119f $X=1.845 $Y=1.515 $X2=0
+ $Y2=0
cc_217 N_A1_N_c_175_n N_A_27_74#_c_1056_n 0.0211272f $X=1.77 $Y=1.515 $X2=0
+ $Y2=0
cc_218 N_A1_N_c_176_n N_A_27_74#_c_1056_n 0.00279548f $X=1.845 $Y=1.515 $X2=0
+ $Y2=0
cc_219 N_A1_N_M1032_g N_A_27_74#_c_1057_n 4.03599e-19 $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_220 N_A1_N_M1033_g N_A_27_74#_c_1057_n 4.03599e-19 $X=1.365 $Y=0.74 $X2=0
+ $Y2=0
cc_221 N_A1_N_M1033_g N_A_27_74#_c_1058_n 0.0130699f $X=1.365 $Y=0.74 $X2=0
+ $Y2=0
cc_222 N_A1_N_M1034_g N_A_27_74#_c_1058_n 0.0128967f $X=1.795 $Y=0.74 $X2=0
+ $Y2=0
cc_223 N_A1_N_c_175_n N_A_27_74#_c_1058_n 0.0525922f $X=1.77 $Y=1.515 $X2=0
+ $Y2=0
cc_224 N_A1_N_c_176_n N_A_27_74#_c_1058_n 0.00413938f $X=1.845 $Y=1.515 $X2=0
+ $Y2=0
cc_225 N_A1_N_M1034_g N_A_27_74#_c_1060_n 9.48753e-19 $X=1.795 $Y=0.74 $X2=0
+ $Y2=0
cc_226 N_A1_N_c_175_n N_A_27_74#_c_1063_n 0.0154618f $X=1.77 $Y=1.515 $X2=0
+ $Y2=0
cc_227 N_A1_N_c_176_n N_A_27_74#_c_1063_n 0.00270057f $X=1.845 $Y=1.515 $X2=0
+ $Y2=0
cc_228 N_A1_N_M1012_g N_VGND_c_1122_n 0.0133724f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_229 N_A1_N_M1032_g N_VGND_c_1122_n 0.0103611f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_230 N_A1_N_M1033_g N_VGND_c_1122_n 4.7018e-19 $X=1.365 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A1_N_M1032_g N_VGND_c_1123_n 4.7018e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A1_N_M1033_g N_VGND_c_1123_n 0.0103611f $X=1.365 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A1_N_M1034_g N_VGND_c_1123_n 0.00968343f $X=1.795 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A1_N_M1034_g N_VGND_c_1124_n 0.00383152f $X=1.795 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A1_N_M1012_g N_VGND_c_1129_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A1_N_M1032_g N_VGND_c_1130_n 0.00383152f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A1_N_M1033_g N_VGND_c_1130_n 0.00383152f $X=1.365 $Y=0.74 $X2=0 $Y2=0
cc_238 N_A1_N_M1012_g N_VGND_c_1135_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_239 N_A1_N_M1032_g N_VGND_c_1135_n 0.0075764f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A1_N_M1033_g N_VGND_c_1135_n 0.0075764f $X=1.365 $Y=0.74 $X2=0 $Y2=0
cc_241 N_A1_N_M1034_g N_VGND_c_1135_n 0.00757637f $X=1.795 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A2_N_M1010_g N_A_117_368#_M1014_g 0.0119658f $X=3.645 $Y=2.4 $X2=0
+ $Y2=0
cc_243 N_A2_N_M1039_g N_A_117_368#_c_360_n 0.00590113f $X=3.655 $Y=0.74 $X2=0
+ $Y2=0
cc_244 N_A2_N_c_261_n N_A_117_368#_c_360_n 0.012318f $X=3.555 $Y=1.32 $X2=0
+ $Y2=0
cc_245 N_A2_N_M1000_g N_A_117_368#_c_371_n 6.50516e-19 $X=2.295 $Y=2.4 $X2=0
+ $Y2=0
cc_246 N_A2_N_M1000_g N_A_117_368#_c_389_n 0.0135031f $X=2.295 $Y=2.4 $X2=0
+ $Y2=0
cc_247 A2_N N_A_117_368#_c_389_n 0.00945133f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_248 N_A2_N_M1008_g N_A_117_368#_c_402_n 0.00498003f $X=2.225 $Y=0.74 $X2=0
+ $Y2=0
cc_249 N_A2_N_M1017_g N_A_117_368#_c_402_n 0.00661392f $X=2.655 $Y=0.74 $X2=0
+ $Y2=0
cc_250 N_A2_N_M1022_g N_A_117_368#_c_402_n 5.87434e-19 $X=3.18 $Y=0.74 $X2=0
+ $Y2=0
cc_251 N_A2_N_M1000_g N_A_117_368#_c_372_n 0.0121132f $X=2.295 $Y=2.4 $X2=0
+ $Y2=0
cc_252 N_A2_N_M1003_g N_A_117_368#_c_372_n 0.0121132f $X=2.745 $Y=2.4 $X2=0
+ $Y2=0
cc_253 N_A2_N_M1005_g N_A_117_368#_c_372_n 6.50516e-19 $X=3.195 $Y=2.4 $X2=0
+ $Y2=0
cc_254 N_A2_N_M1017_g N_A_117_368#_c_362_n 0.00952207f $X=2.655 $Y=0.74 $X2=0
+ $Y2=0
cc_255 N_A2_N_M1022_g N_A_117_368#_c_362_n 0.0132432f $X=3.18 $Y=0.74 $X2=0
+ $Y2=0
cc_256 A2_N N_A_117_368#_c_362_n 0.0473393f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_257 N_A2_N_c_262_n N_A_117_368#_c_362_n 0.00499391f $X=3.285 $Y=1.5 $X2=0
+ $Y2=0
cc_258 N_A2_N_M1008_g N_A_117_368#_c_363_n 0.00407645f $X=2.225 $Y=0.74 $X2=0
+ $Y2=0
cc_259 N_A2_N_M1017_g N_A_117_368#_c_363_n 0.00271614f $X=2.655 $Y=0.74 $X2=0
+ $Y2=0
cc_260 A2_N N_A_117_368#_c_363_n 0.027784f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_261 N_A2_N_c_262_n N_A_117_368#_c_363_n 0.00275304f $X=3.285 $Y=1.5 $X2=0
+ $Y2=0
cc_262 N_A2_N_M1003_g N_A_117_368#_c_416_n 0.012931f $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_263 N_A2_N_M1005_g N_A_117_368#_c_416_n 0.0135113f $X=3.195 $Y=2.4 $X2=0
+ $Y2=0
cc_264 A2_N N_A_117_368#_c_416_n 0.0377615f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_265 N_A2_N_c_262_n N_A_117_368#_c_416_n 4.90053e-19 $X=3.285 $Y=1.5 $X2=0
+ $Y2=0
cc_266 N_A2_N_M1003_g N_A_117_368#_c_373_n 6.50516e-19 $X=2.745 $Y=2.4 $X2=0
+ $Y2=0
cc_267 N_A2_N_M1005_g N_A_117_368#_c_373_n 0.0121132f $X=3.195 $Y=2.4 $X2=0
+ $Y2=0
cc_268 N_A2_N_M1010_g N_A_117_368#_c_373_n 0.0108828f $X=3.645 $Y=2.4 $X2=0
+ $Y2=0
cc_269 N_A2_N_M1039_g N_A_117_368#_c_423_n 0.00567006f $X=3.655 $Y=0.74 $X2=0
+ $Y2=0
cc_270 N_A2_N_M1022_g N_A_117_368#_c_364_n 0.00319592f $X=3.18 $Y=0.74 $X2=0
+ $Y2=0
cc_271 N_A2_N_c_258_n N_A_117_368#_c_364_n 0.0114992f $X=3.555 $Y=1.395 $X2=0
+ $Y2=0
cc_272 N_A2_N_M1010_g N_A_117_368#_c_364_n 0.0018418f $X=3.645 $Y=2.4 $X2=0
+ $Y2=0
cc_273 N_A2_N_M1039_g N_A_117_368#_c_364_n 0.0115523f $X=3.655 $Y=0.74 $X2=0
+ $Y2=0
cc_274 N_A2_N_c_261_n N_A_117_368#_c_364_n 0.00175427f $X=3.555 $Y=1.32 $X2=0
+ $Y2=0
cc_275 A2_N N_A_117_368#_c_364_n 0.0232738f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_276 N_A2_N_c_262_n N_A_117_368#_c_364_n 0.00135651f $X=3.285 $Y=1.5 $X2=0
+ $Y2=0
cc_277 N_A2_N_M1010_g N_A_117_368#_c_374_n 0.00639039f $X=3.645 $Y=2.4 $X2=0
+ $Y2=0
cc_278 A2_N N_A_117_368#_c_374_n 0.0113234f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_279 N_A2_N_c_262_n N_A_117_368#_c_374_n 0.0042775f $X=3.285 $Y=1.5 $X2=0
+ $Y2=0
cc_280 N_A2_N_M1010_g N_A_117_368#_c_365_n 0.00775752f $X=3.645 $Y=2.4 $X2=0
+ $Y2=0
cc_281 N_A2_N_M1039_g N_A_117_368#_c_365_n 0.00637964f $X=3.655 $Y=0.74 $X2=0
+ $Y2=0
cc_282 N_A2_N_c_261_n N_A_117_368#_c_365_n 0.006096f $X=3.555 $Y=1.32 $X2=0
+ $Y2=0
cc_283 N_A2_N_M1000_g N_A_117_368#_c_437_n 8.84614e-19 $X=2.295 $Y=2.4 $X2=0
+ $Y2=0
cc_284 N_A2_N_M1003_g N_A_117_368#_c_437_n 8.84614e-19 $X=2.745 $Y=2.4 $X2=0
+ $Y2=0
cc_285 A2_N N_A_117_368#_c_437_n 0.0235495f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_286 N_A2_N_c_262_n N_A_117_368#_c_437_n 5.49354e-19 $X=3.285 $Y=1.5 $X2=0
+ $Y2=0
cc_287 N_A2_N_M1005_g N_A_117_368#_c_441_n 0.00196977f $X=3.195 $Y=2.4 $X2=0
+ $Y2=0
cc_288 N_A2_N_c_258_n N_A_117_368#_c_441_n 0.00118718f $X=3.555 $Y=1.395 $X2=0
+ $Y2=0
cc_289 N_A2_N_M1010_g N_A_117_368#_c_441_n 0.0020266f $X=3.645 $Y=2.4 $X2=0
+ $Y2=0
cc_290 N_A2_N_M1000_g N_VPWR_c_734_n 0.0027763f $X=2.295 $Y=2.4 $X2=0 $Y2=0
cc_291 N_A2_N_M1003_g N_VPWR_c_735_n 0.0027763f $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_292 N_A2_N_M1005_g N_VPWR_c_735_n 0.0027763f $X=3.195 $Y=2.4 $X2=0 $Y2=0
cc_293 N_A2_N_M1010_g N_VPWR_c_736_n 0.00313866f $X=3.645 $Y=2.4 $X2=0 $Y2=0
cc_294 N_A2_N_M1000_g N_VPWR_c_746_n 0.005209f $X=2.295 $Y=2.4 $X2=0 $Y2=0
cc_295 N_A2_N_M1003_g N_VPWR_c_746_n 0.005209f $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_296 N_A2_N_M1005_g N_VPWR_c_748_n 0.005209f $X=3.195 $Y=2.4 $X2=0 $Y2=0
cc_297 N_A2_N_M1010_g N_VPWR_c_748_n 0.005209f $X=3.645 $Y=2.4 $X2=0 $Y2=0
cc_298 N_A2_N_M1000_g N_VPWR_c_730_n 0.00982376f $X=2.295 $Y=2.4 $X2=0 $Y2=0
cc_299 N_A2_N_M1003_g N_VPWR_c_730_n 0.00982266f $X=2.745 $Y=2.4 $X2=0 $Y2=0
cc_300 N_A2_N_M1005_g N_VPWR_c_730_n 0.00982266f $X=3.195 $Y=2.4 $X2=0 $Y2=0
cc_301 N_A2_N_M1010_g N_VPWR_c_730_n 0.00982376f $X=3.645 $Y=2.4 $X2=0 $Y2=0
cc_302 N_A2_N_M1008_g N_A_27_74#_c_1058_n 5.7448e-19 $X=2.225 $Y=0.74 $X2=0
+ $Y2=0
cc_303 N_A2_N_M1008_g N_A_27_74#_c_1059_n 0.0120041f $X=2.225 $Y=0.74 $X2=0
+ $Y2=0
cc_304 N_A2_N_M1017_g N_A_27_74#_c_1059_n 0.0112986f $X=2.655 $Y=0.74 $X2=0
+ $Y2=0
cc_305 N_A2_N_M1022_g N_A_27_74#_c_1061_n 0.00938114f $X=3.18 $Y=0.74 $X2=0
+ $Y2=0
cc_306 N_A2_N_M1039_g N_A_27_74#_c_1061_n 0.0135229f $X=3.655 $Y=0.74 $X2=0
+ $Y2=0
cc_307 N_A2_N_M1039_g N_A_27_74#_c_1062_n 0.00159289f $X=3.655 $Y=0.74 $X2=0
+ $Y2=0
cc_308 N_A2_N_M1022_g N_A_27_74#_c_1064_n 0.00217786f $X=3.18 $Y=0.74 $X2=0
+ $Y2=0
cc_309 N_A2_N_M1008_g N_VGND_c_1124_n 0.00278271f $X=2.225 $Y=0.74 $X2=0 $Y2=0
cc_310 N_A2_N_M1017_g N_VGND_c_1124_n 0.00278271f $X=2.655 $Y=0.74 $X2=0 $Y2=0
cc_311 N_A2_N_M1022_g N_VGND_c_1124_n 0.00278271f $X=3.18 $Y=0.74 $X2=0 $Y2=0
cc_312 N_A2_N_M1039_g N_VGND_c_1124_n 0.00278271f $X=3.655 $Y=0.74 $X2=0 $Y2=0
cc_313 N_A2_N_M1008_g N_VGND_c_1135_n 0.00353526f $X=2.225 $Y=0.74 $X2=0 $Y2=0
cc_314 N_A2_N_M1017_g N_VGND_c_1135_n 0.00354301f $X=2.655 $Y=0.74 $X2=0 $Y2=0
cc_315 N_A2_N_M1022_g N_VGND_c_1135_n 0.00354734f $X=3.18 $Y=0.74 $X2=0 $Y2=0
cc_316 N_A2_N_M1039_g N_VGND_c_1135_n 0.0035886f $X=3.655 $Y=0.74 $X2=0 $Y2=0
cc_317 N_A2_N_M1039_g N_A_857_74#_c_1253_n 5.96586e-19 $X=3.655 $Y=0.74 $X2=0
+ $Y2=0
cc_318 N_A_117_368#_M1029_g N_B2_M1002_g 0.0115453f $X=5.935 $Y=0.74 $X2=0 $Y2=0
cc_319 N_A_117_368#_c_359_n N_B2_c_563_n 0.0125083f $X=5.86 $Y=1.375 $X2=0 $Y2=0
cc_320 N_A_117_368#_c_360_n N_B2_c_563_n 5.44913e-19 $X=5.58 $Y=1.375 $X2=0
+ $Y2=0
cc_321 N_A_117_368#_c_359_n N_B2_c_564_n 0.0115453f $X=5.86 $Y=1.375 $X2=0 $Y2=0
cc_322 N_A_117_368#_c_360_n N_B2_c_564_n 0.00141988f $X=5.58 $Y=1.375 $X2=0
+ $Y2=0
cc_323 N_A_117_368#_c_382_n N_VPWR_M1027_s 0.00314376f $X=1.455 $Y=2.035 $X2=0
+ $Y2=0
cc_324 N_A_117_368#_c_389_n N_VPWR_M1036_s 0.00761058f $X=2.355 $Y=2.035 $X2=0
+ $Y2=0
cc_325 N_A_117_368#_c_416_n N_VPWR_M1003_s 0.00314376f $X=3.255 $Y=2.035 $X2=0
+ $Y2=0
cc_326 N_A_117_368#_c_370_n N_VPWR_c_732_n 0.0289761f $X=0.72 $Y=2.815 $X2=0
+ $Y2=0
cc_327 N_A_117_368#_c_370_n N_VPWR_c_733_n 0.0233699f $X=0.72 $Y=2.815 $X2=0
+ $Y2=0
cc_328 N_A_117_368#_c_382_n N_VPWR_c_733_n 0.0126919f $X=1.455 $Y=2.035 $X2=0
+ $Y2=0
cc_329 N_A_117_368#_c_371_n N_VPWR_c_733_n 0.0233699f $X=1.62 $Y=2.815 $X2=0
+ $Y2=0
cc_330 N_A_117_368#_c_371_n N_VPWR_c_734_n 0.0233699f $X=1.62 $Y=2.815 $X2=0
+ $Y2=0
cc_331 N_A_117_368#_c_389_n N_VPWR_c_734_n 0.0126919f $X=2.355 $Y=2.035 $X2=0
+ $Y2=0
cc_332 N_A_117_368#_c_372_n N_VPWR_c_734_n 0.0233699f $X=2.52 $Y=2.815 $X2=0
+ $Y2=0
cc_333 N_A_117_368#_c_372_n N_VPWR_c_735_n 0.0233699f $X=2.52 $Y=2.815 $X2=0
+ $Y2=0
cc_334 N_A_117_368#_c_416_n N_VPWR_c_735_n 0.0126919f $X=3.255 $Y=2.035 $X2=0
+ $Y2=0
cc_335 N_A_117_368#_c_373_n N_VPWR_c_735_n 0.0233699f $X=3.42 $Y=2.815 $X2=0
+ $Y2=0
cc_336 N_A_117_368#_M1014_g N_VPWR_c_736_n 0.00313838f $X=4.095 $Y=2.4 $X2=0
+ $Y2=0
cc_337 N_A_117_368#_c_373_n N_VPWR_c_736_n 0.0289376f $X=3.42 $Y=2.815 $X2=0
+ $Y2=0
cc_338 N_A_117_368#_c_374_n N_VPWR_c_736_n 0.00447613f $X=3.5 $Y=1.95 $X2=0
+ $Y2=0
cc_339 N_A_117_368#_c_365_n N_VPWR_c_736_n 0.0137368f $X=5.26 $Y=1.465 $X2=0
+ $Y2=0
cc_340 N_A_117_368#_M1019_g N_VPWR_c_737_n 0.00329146f $X=4.545 $Y=2.4 $X2=0
+ $Y2=0
cc_341 N_A_117_368#_M1021_g N_VPWR_c_737_n 0.00208338f $X=4.995 $Y=2.4 $X2=0
+ $Y2=0
cc_342 N_A_117_368#_M1021_g N_VPWR_c_738_n 0.005209f $X=4.995 $Y=2.4 $X2=0 $Y2=0
cc_343 N_A_117_368#_M1028_g N_VPWR_c_738_n 0.00460063f $X=5.445 $Y=2.4 $X2=0
+ $Y2=0
cc_344 N_A_117_368#_M1021_g N_VPWR_c_739_n 5.61186e-19 $X=4.995 $Y=2.4 $X2=0
+ $Y2=0
cc_345 N_A_117_368#_M1028_g N_VPWR_c_739_n 0.0140603f $X=5.445 $Y=2.4 $X2=0
+ $Y2=0
cc_346 N_A_117_368#_c_370_n N_VPWR_c_742_n 0.0144623f $X=0.72 $Y=2.815 $X2=0
+ $Y2=0
cc_347 N_A_117_368#_c_371_n N_VPWR_c_744_n 0.0144623f $X=1.62 $Y=2.815 $X2=0
+ $Y2=0
cc_348 N_A_117_368#_c_372_n N_VPWR_c_746_n 0.0144623f $X=2.52 $Y=2.815 $X2=0
+ $Y2=0
cc_349 N_A_117_368#_c_373_n N_VPWR_c_748_n 0.0144623f $X=3.42 $Y=2.815 $X2=0
+ $Y2=0
cc_350 N_A_117_368#_M1014_g N_VPWR_c_750_n 0.005209f $X=4.095 $Y=2.4 $X2=0 $Y2=0
cc_351 N_A_117_368#_M1019_g N_VPWR_c_750_n 0.005209f $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_352 N_A_117_368#_M1014_g N_VPWR_c_730_n 0.00982376f $X=4.095 $Y=2.4 $X2=0
+ $Y2=0
cc_353 N_A_117_368#_M1019_g N_VPWR_c_730_n 0.00982266f $X=4.545 $Y=2.4 $X2=0
+ $Y2=0
cc_354 N_A_117_368#_M1021_g N_VPWR_c_730_n 0.00982266f $X=4.995 $Y=2.4 $X2=0
+ $Y2=0
cc_355 N_A_117_368#_M1028_g N_VPWR_c_730_n 0.00908554f $X=5.445 $Y=2.4 $X2=0
+ $Y2=0
cc_356 N_A_117_368#_c_370_n N_VPWR_c_730_n 0.0118344f $X=0.72 $Y=2.815 $X2=0
+ $Y2=0
cc_357 N_A_117_368#_c_371_n N_VPWR_c_730_n 0.0118344f $X=1.62 $Y=2.815 $X2=0
+ $Y2=0
cc_358 N_A_117_368#_c_372_n N_VPWR_c_730_n 0.0118344f $X=2.52 $Y=2.815 $X2=0
+ $Y2=0
cc_359 N_A_117_368#_c_373_n N_VPWR_c_730_n 0.0118344f $X=3.42 $Y=2.815 $X2=0
+ $Y2=0
cc_360 N_A_117_368#_M1014_g N_Y_c_884_n 0.0130723f $X=4.095 $Y=2.4 $X2=0 $Y2=0
cc_361 N_A_117_368#_M1019_g N_Y_c_884_n 0.0143001f $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_362 N_A_117_368#_M1021_g N_Y_c_884_n 6.9775e-19 $X=4.995 $Y=2.4 $X2=0 $Y2=0
cc_363 N_A_117_368#_M1019_g N_Y_c_885_n 0.012931f $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_364 N_A_117_368#_M1021_g N_Y_c_885_n 0.012931f $X=4.995 $Y=2.4 $X2=0 $Y2=0
cc_365 N_A_117_368#_c_360_n N_Y_c_885_n 0.00235274f $X=5.58 $Y=1.375 $X2=0 $Y2=0
cc_366 N_A_117_368#_c_365_n N_Y_c_885_n 0.0416512f $X=5.26 $Y=1.465 $X2=0 $Y2=0
cc_367 N_A_117_368#_M1014_g N_Y_c_886_n 0.0030623f $X=4.095 $Y=2.4 $X2=0 $Y2=0
cc_368 N_A_117_368#_M1019_g N_Y_c_886_n 0.00135419f $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_369 N_A_117_368#_c_360_n N_Y_c_886_n 0.00209661f $X=5.58 $Y=1.375 $X2=0 $Y2=0
cc_370 N_A_117_368#_c_374_n N_Y_c_886_n 5.60546e-19 $X=3.5 $Y=1.95 $X2=0 $Y2=0
cc_371 N_A_117_368#_c_365_n N_Y_c_886_n 0.0275631f $X=5.26 $Y=1.465 $X2=0 $Y2=0
cc_372 N_A_117_368#_M1009_g N_Y_c_903_n 0.00515339f $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_373 N_A_117_368#_M1018_g N_Y_c_903_n 0.00611761f $X=5.075 $Y=0.74 $X2=0 $Y2=0
cc_374 N_A_117_368#_M1023_g N_Y_c_903_n 5.55764e-19 $X=5.505 $Y=0.74 $X2=0 $Y2=0
cc_375 N_A_117_368#_M1018_g N_Y_c_880_n 0.00885064f $X=5.075 $Y=0.74 $X2=0 $Y2=0
cc_376 N_A_117_368#_M1023_g N_Y_c_880_n 0.00995138f $X=5.505 $Y=0.74 $X2=0 $Y2=0
cc_377 N_A_117_368#_c_360_n N_Y_c_880_n 0.00253755f $X=5.58 $Y=1.375 $X2=0 $Y2=0
cc_378 N_A_117_368#_c_365_n N_Y_c_880_n 0.0258049f $X=5.26 $Y=1.465 $X2=0 $Y2=0
cc_379 N_A_117_368#_M1009_g N_Y_c_881_n 0.00310933f $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_380 N_A_117_368#_M1018_g N_Y_c_881_n 0.00163137f $X=5.075 $Y=0.74 $X2=0 $Y2=0
cc_381 N_A_117_368#_c_360_n N_Y_c_881_n 0.0026843f $X=5.58 $Y=1.375 $X2=0 $Y2=0
cc_382 N_A_117_368#_c_365_n N_Y_c_881_n 0.0270731f $X=5.26 $Y=1.465 $X2=0 $Y2=0
cc_383 N_A_117_368#_M1021_g N_Y_c_887_n 0.0107378f $X=4.995 $Y=2.4 $X2=0 $Y2=0
cc_384 N_A_117_368#_M1028_g N_Y_c_887_n 3.68116e-19 $X=5.445 $Y=2.4 $X2=0 $Y2=0
cc_385 N_A_117_368#_M1018_g N_Y_c_916_n 5.64138e-19 $X=5.075 $Y=0.74 $X2=0 $Y2=0
cc_386 N_A_117_368#_M1023_g N_Y_c_916_n 0.00646632f $X=5.505 $Y=0.74 $X2=0 $Y2=0
cc_387 N_A_117_368#_M1029_g N_Y_c_916_n 0.00494352f $X=5.935 $Y=0.74 $X2=0 $Y2=0
cc_388 N_A_117_368#_M1018_g N_Y_c_882_n 8.44792e-19 $X=5.075 $Y=0.74 $X2=0 $Y2=0
cc_389 N_A_117_368#_M1023_g N_Y_c_882_n 0.00419028f $X=5.505 $Y=0.74 $X2=0 $Y2=0
cc_390 N_A_117_368#_c_359_n N_Y_c_882_n 0.00830694f $X=5.86 $Y=1.375 $X2=0 $Y2=0
cc_391 N_A_117_368#_c_360_n N_Y_c_882_n 0.0158931f $X=5.58 $Y=1.375 $X2=0 $Y2=0
cc_392 N_A_117_368#_M1029_g N_Y_c_882_n 0.00294584f $X=5.935 $Y=0.74 $X2=0 $Y2=0
cc_393 N_A_117_368#_c_365_n N_Y_c_882_n 0.0250936f $X=5.26 $Y=1.465 $X2=0 $Y2=0
cc_394 N_A_117_368#_c_359_n N_Y_c_889_n 0.00510836f $X=5.86 $Y=1.375 $X2=0 $Y2=0
cc_395 N_A_117_368#_M1019_g N_Y_c_890_n 4.34352e-19 $X=4.545 $Y=2.4 $X2=0 $Y2=0
cc_396 N_A_117_368#_M1021_g N_Y_c_890_n 0.00472982f $X=4.995 $Y=2.4 $X2=0 $Y2=0
cc_397 N_A_117_368#_M1028_g N_Y_c_890_n 0.026106f $X=5.445 $Y=2.4 $X2=0 $Y2=0
cc_398 N_A_117_368#_c_360_n N_Y_c_890_n 0.00266697f $X=5.58 $Y=1.375 $X2=0 $Y2=0
cc_399 N_A_117_368#_c_365_n N_Y_c_890_n 0.0264621f $X=5.26 $Y=1.465 $X2=0 $Y2=0
cc_400 N_A_117_368#_M1023_g N_Y_c_883_n 0.00144713f $X=5.505 $Y=0.74 $X2=0 $Y2=0
cc_401 N_A_117_368#_c_359_n N_Y_c_883_n 0.00217378f $X=5.86 $Y=1.375 $X2=0 $Y2=0
cc_402 N_A_117_368#_M1029_g N_Y_c_883_n 0.00375789f $X=5.935 $Y=0.74 $X2=0 $Y2=0
cc_403 N_A_117_368#_M1028_g N_A_1215_368#_c_988_n 9.69578e-19 $X=5.445 $Y=2.4
+ $X2=0 $Y2=0
cc_404 N_A_117_368#_M1028_g N_A_1215_368#_c_990_n 5.99495e-19 $X=5.445 $Y=2.4
+ $X2=0 $Y2=0
cc_405 N_A_117_368#_c_362_n N_A_27_74#_M1017_d 0.00285668f $X=3.275 $Y=1.095
+ $X2=0 $Y2=0
cc_406 N_A_117_368#_c_363_n N_A_27_74#_c_1058_n 0.00997012f $X=2.605 $Y=1.095
+ $X2=0 $Y2=0
cc_407 N_A_117_368#_M1008_s N_A_27_74#_c_1059_n 0.00176461f $X=2.3 $Y=0.37 $X2=0
+ $Y2=0
cc_408 N_A_117_368#_c_402_n N_A_27_74#_c_1059_n 0.0158692f $X=2.44 $Y=0.82 $X2=0
+ $Y2=0
cc_409 N_A_117_368#_c_362_n N_A_27_74#_c_1059_n 0.00304353f $X=3.275 $Y=1.095
+ $X2=0 $Y2=0
cc_410 N_A_117_368#_c_362_n N_A_27_74#_c_1093_n 0.020976f $X=3.275 $Y=1.095
+ $X2=0 $Y2=0
cc_411 N_A_117_368#_M1022_s N_A_27_74#_c_1061_n 0.00224297f $X=3.255 $Y=0.37
+ $X2=0 $Y2=0
cc_412 N_A_117_368#_M1009_g N_A_27_74#_c_1061_n 5.96586e-19 $X=4.645 $Y=0.74
+ $X2=0 $Y2=0
cc_413 N_A_117_368#_c_362_n N_A_27_74#_c_1061_n 0.00364245f $X=3.275 $Y=1.095
+ $X2=0 $Y2=0
cc_414 N_A_117_368#_c_423_n N_A_27_74#_c_1061_n 0.0176798f $X=3.44 $Y=0.86 $X2=0
+ $Y2=0
cc_415 N_A_117_368#_c_364_n N_A_27_74#_c_1062_n 0.00555794f $X=3.5 $Y=1.63 $X2=0
+ $Y2=0
cc_416 N_A_117_368#_c_365_n N_A_27_74#_c_1062_n 0.0219383f $X=5.26 $Y=1.465
+ $X2=0 $Y2=0
cc_417 N_A_117_368#_M1009_g N_VGND_c_1124_n 0.00278271f $X=4.645 $Y=0.74 $X2=0
+ $Y2=0
cc_418 N_A_117_368#_M1018_g N_VGND_c_1124_n 0.00278271f $X=5.075 $Y=0.74 $X2=0
+ $Y2=0
cc_419 N_A_117_368#_M1023_g N_VGND_c_1124_n 0.00278271f $X=5.505 $Y=0.74 $X2=0
+ $Y2=0
cc_420 N_A_117_368#_M1029_g N_VGND_c_1124_n 0.00278271f $X=5.935 $Y=0.74 $X2=0
+ $Y2=0
cc_421 N_A_117_368#_M1009_g N_VGND_c_1135_n 0.00358427f $X=4.645 $Y=0.74 $X2=0
+ $Y2=0
cc_422 N_A_117_368#_M1018_g N_VGND_c_1135_n 0.00353428f $X=5.075 $Y=0.74 $X2=0
+ $Y2=0
cc_423 N_A_117_368#_M1023_g N_VGND_c_1135_n 0.00353428f $X=5.505 $Y=0.74 $X2=0
+ $Y2=0
cc_424 N_A_117_368#_M1029_g N_VGND_c_1135_n 0.00353526f $X=5.935 $Y=0.74 $X2=0
+ $Y2=0
cc_425 N_A_117_368#_M1009_g N_A_857_74#_c_1251_n 0.00159289f $X=4.645 $Y=0.74
+ $X2=0 $Y2=0
cc_426 N_A_117_368#_c_360_n N_A_857_74#_c_1251_n 0.0064005f $X=5.58 $Y=1.375
+ $X2=0 $Y2=0
cc_427 N_A_117_368#_c_365_n N_A_857_74#_c_1251_n 0.0209147f $X=5.26 $Y=1.465
+ $X2=0 $Y2=0
cc_428 N_A_117_368#_M1009_g N_A_857_74#_c_1252_n 0.0132617f $X=4.645 $Y=0.74
+ $X2=0 $Y2=0
cc_429 N_A_117_368#_M1018_g N_A_857_74#_c_1252_n 0.0100569f $X=5.075 $Y=0.74
+ $X2=0 $Y2=0
cc_430 N_A_117_368#_M1023_g N_A_857_74#_c_1254_n 0.00988997f $X=5.505 $Y=0.74
+ $X2=0 $Y2=0
cc_431 N_A_117_368#_M1029_g N_A_857_74#_c_1254_n 0.0120041f $X=5.935 $Y=0.74
+ $X2=0 $Y2=0
cc_432 N_A_117_368#_M1029_g N_A_857_74#_c_1256_n 7.38995e-19 $X=5.935 $Y=0.74
+ $X2=0 $Y2=0
cc_433 N_B2_M1037_g N_B1_M1007_g 0.012736f $X=7.785 $Y=2.4 $X2=0 $Y2=0
cc_434 N_B2_M1038_g N_B1_M1006_g 0.0195038f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_435 N_B2_c_563_n B1 0.0150955f $X=7.475 $Y=1.515 $X2=0 $Y2=0
cc_436 N_B2_c_564_n B1 0.00199057f $X=7.795 $Y=1.515 $X2=0 $Y2=0
cc_437 N_B2_c_563_n N_B1_c_654_n 6.26242e-19 $X=7.475 $Y=1.515 $X2=0 $Y2=0
cc_438 N_B2_c_564_n N_B1_c_654_n 0.0213985f $X=7.795 $Y=1.515 $X2=0 $Y2=0
cc_439 N_B2_M1001_g N_VPWR_c_739_n 8.9486e-19 $X=6.435 $Y=2.4 $X2=0 $Y2=0
cc_440 N_B2_M1001_g N_VPWR_c_752_n 0.00333926f $X=6.435 $Y=2.4 $X2=0 $Y2=0
cc_441 N_B2_M1004_g N_VPWR_c_752_n 0.00333926f $X=6.885 $Y=2.4 $X2=0 $Y2=0
cc_442 N_B2_M1031_g N_VPWR_c_752_n 0.00333926f $X=7.335 $Y=2.4 $X2=0 $Y2=0
cc_443 N_B2_M1037_g N_VPWR_c_752_n 0.00333926f $X=7.785 $Y=2.4 $X2=0 $Y2=0
cc_444 N_B2_M1001_g N_VPWR_c_730_n 0.0042782f $X=6.435 $Y=2.4 $X2=0 $Y2=0
cc_445 N_B2_M1004_g N_VPWR_c_730_n 0.00422687f $X=6.885 $Y=2.4 $X2=0 $Y2=0
cc_446 N_B2_M1031_g N_VPWR_c_730_n 0.00422687f $X=7.335 $Y=2.4 $X2=0 $Y2=0
cc_447 N_B2_M1037_g N_VPWR_c_730_n 0.00422798f $X=7.785 $Y=2.4 $X2=0 $Y2=0
cc_448 N_B2_M1001_g N_Y_c_882_n 7.22654e-19 $X=6.435 $Y=2.4 $X2=0 $Y2=0
cc_449 N_B2_c_563_n N_Y_c_882_n 0.035327f $X=7.475 $Y=1.515 $X2=0 $Y2=0
cc_450 N_B2_c_564_n N_Y_c_882_n 5.42229e-19 $X=7.795 $Y=1.515 $X2=0 $Y2=0
cc_451 N_B2_M1001_g N_Y_c_889_n 0.0150541f $X=6.435 $Y=2.4 $X2=0 $Y2=0
cc_452 N_B2_c_563_n N_Y_c_889_n 0.0457335f $X=7.475 $Y=1.515 $X2=0 $Y2=0
cc_453 N_B2_M1001_g N_Y_c_890_n 0.00389737f $X=6.435 $Y=2.4 $X2=0 $Y2=0
cc_454 N_B2_M1004_g N_Y_c_940_n 0.012931f $X=6.885 $Y=2.4 $X2=0 $Y2=0
cc_455 N_B2_M1031_g N_Y_c_940_n 0.012931f $X=7.335 $Y=2.4 $X2=0 $Y2=0
cc_456 N_B2_c_563_n N_Y_c_940_n 0.0391869f $X=7.475 $Y=1.515 $X2=0 $Y2=0
cc_457 N_B2_c_564_n N_Y_c_940_n 4.89004e-19 $X=7.795 $Y=1.515 $X2=0 $Y2=0
cc_458 N_B2_M1001_g N_Y_c_944_n 0.0159493f $X=6.435 $Y=2.4 $X2=0 $Y2=0
cc_459 N_B2_M1004_g N_Y_c_944_n 0.01146f $X=6.885 $Y=2.4 $X2=0 $Y2=0
cc_460 N_B2_M1031_g N_Y_c_944_n 5.63205e-19 $X=7.335 $Y=2.4 $X2=0 $Y2=0
cc_461 N_B2_c_563_n N_Y_c_944_n 0.0235495f $X=7.475 $Y=1.515 $X2=0 $Y2=0
cc_462 N_B2_c_564_n N_Y_c_944_n 5.54423e-19 $X=7.795 $Y=1.515 $X2=0 $Y2=0
cc_463 N_B2_M1004_g N_Y_c_949_n 5.63205e-19 $X=6.885 $Y=2.4 $X2=0 $Y2=0
cc_464 N_B2_M1031_g N_Y_c_949_n 0.01146f $X=7.335 $Y=2.4 $X2=0 $Y2=0
cc_465 N_B2_M1037_g N_Y_c_949_n 0.0127383f $X=7.785 $Y=2.4 $X2=0 $Y2=0
cc_466 N_B2_c_563_n N_Y_c_949_n 0.0187567f $X=7.475 $Y=1.515 $X2=0 $Y2=0
cc_467 N_B2_c_564_n N_Y_c_949_n 5.54777e-19 $X=7.795 $Y=1.515 $X2=0 $Y2=0
cc_468 N_B2_M1001_g N_A_1215_368#_c_989_n 0.0149887f $X=6.435 $Y=2.4 $X2=0 $Y2=0
cc_469 N_B2_M1004_g N_A_1215_368#_c_989_n 0.0140221f $X=6.885 $Y=2.4 $X2=0 $Y2=0
cc_470 N_B2_M1031_g N_A_1215_368#_c_991_n 0.0139834f $X=7.335 $Y=2.4 $X2=0 $Y2=0
cc_471 N_B2_M1037_g N_A_1215_368#_c_991_n 0.0137347f $X=7.785 $Y=2.4 $X2=0 $Y2=0
cc_472 N_B2_M1002_g N_VGND_c_1124_n 0.00383152f $X=6.365 $Y=0.74 $X2=0 $Y2=0
cc_473 N_B2_M1002_g N_VGND_c_1125_n 0.00964869f $X=6.365 $Y=0.74 $X2=0 $Y2=0
cc_474 N_B2_M1024_g N_VGND_c_1125_n 0.00418685f $X=6.865 $Y=0.74 $X2=0 $Y2=0
cc_475 N_B2_M1024_g N_VGND_c_1126_n 5.14838e-19 $X=6.865 $Y=0.74 $X2=0 $Y2=0
cc_476 N_B2_M1025_g N_VGND_c_1126_n 0.010415f $X=7.295 $Y=0.74 $X2=0 $Y2=0
cc_477 N_B2_M1038_g N_VGND_c_1126_n 0.00418685f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_478 N_B2_M1038_g N_VGND_c_1127_n 5.14838e-19 $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_479 N_B2_M1024_g N_VGND_c_1131_n 0.00434272f $X=6.865 $Y=0.74 $X2=0 $Y2=0
cc_480 N_B2_M1025_g N_VGND_c_1131_n 0.00383152f $X=7.295 $Y=0.74 $X2=0 $Y2=0
cc_481 N_B2_M1038_g N_VGND_c_1132_n 0.00434272f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_482 N_B2_M1002_g N_VGND_c_1135_n 0.00757637f $X=6.365 $Y=0.74 $X2=0 $Y2=0
cc_483 N_B2_M1024_g N_VGND_c_1135_n 0.00820718f $X=6.865 $Y=0.74 $X2=0 $Y2=0
cc_484 N_B2_M1025_g N_VGND_c_1135_n 0.0075754f $X=7.295 $Y=0.74 $X2=0 $Y2=0
cc_485 N_B2_M1038_g N_VGND_c_1135_n 0.00820816f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_486 N_B2_M1002_g N_A_857_74#_c_1254_n 9.48753e-19 $X=6.365 $Y=0.74 $X2=0
+ $Y2=0
cc_487 N_B2_M1002_g N_A_857_74#_c_1255_n 0.0132997f $X=6.365 $Y=0.74 $X2=0 $Y2=0
cc_488 N_B2_M1024_g N_A_857_74#_c_1255_n 0.0115433f $X=6.865 $Y=0.74 $X2=0 $Y2=0
cc_489 N_B2_c_563_n N_A_857_74#_c_1255_n 0.051298f $X=7.475 $Y=1.515 $X2=0 $Y2=0
cc_490 N_B2_c_564_n N_A_857_74#_c_1255_n 0.00414639f $X=7.795 $Y=1.515 $X2=0
+ $Y2=0
cc_491 N_B2_c_563_n N_A_857_74#_c_1256_n 0.0153286f $X=7.475 $Y=1.515 $X2=0
+ $Y2=0
cc_492 N_B2_M1002_g N_A_857_74#_c_1257_n 9.78807e-19 $X=6.365 $Y=0.74 $X2=0
+ $Y2=0
cc_493 N_B2_M1024_g N_A_857_74#_c_1257_n 0.00922099f $X=6.865 $Y=0.74 $X2=0
+ $Y2=0
cc_494 N_B2_M1025_g N_A_857_74#_c_1257_n 3.97481e-19 $X=7.295 $Y=0.74 $X2=0
+ $Y2=0
cc_495 N_B2_M1025_g N_A_857_74#_c_1258_n 0.0134949f $X=7.295 $Y=0.74 $X2=0 $Y2=0
cc_496 N_B2_M1038_g N_A_857_74#_c_1258_n 0.0153304f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_497 N_B2_c_563_n N_A_857_74#_c_1258_n 0.0358392f $X=7.475 $Y=1.515 $X2=0
+ $Y2=0
cc_498 N_B2_c_564_n N_A_857_74#_c_1258_n 0.00412669f $X=7.795 $Y=1.515 $X2=0
+ $Y2=0
cc_499 N_B2_M1025_g N_A_857_74#_c_1259_n 9.78807e-19 $X=7.295 $Y=0.74 $X2=0
+ $Y2=0
cc_500 N_B2_M1038_g N_A_857_74#_c_1259_n 0.00922099f $X=7.795 $Y=0.74 $X2=0
+ $Y2=0
cc_501 N_B2_M1024_g N_A_857_74#_c_1265_n 0.00157732f $X=6.865 $Y=0.74 $X2=0
+ $Y2=0
cc_502 N_B2_c_563_n N_A_857_74#_c_1265_n 0.0213626f $X=7.475 $Y=1.515 $X2=0
+ $Y2=0
cc_503 N_B2_c_564_n N_A_857_74#_c_1265_n 0.00246761f $X=7.795 $Y=1.515 $X2=0
+ $Y2=0
cc_504 N_B2_M1038_g N_A_857_74#_c_1266_n 0.00249368f $X=7.795 $Y=0.74 $X2=0
+ $Y2=0
cc_505 N_B2_c_564_n N_A_857_74#_c_1266_n 2.41927e-19 $X=7.795 $Y=1.515 $X2=0
+ $Y2=0
cc_506 N_B1_M1007_g N_VPWR_c_740_n 0.0115016f $X=8.235 $Y=2.4 $X2=0 $Y2=0
cc_507 N_B1_M1011_g N_VPWR_c_740_n 0.0030671f $X=8.685 $Y=2.4 $X2=0 $Y2=0
cc_508 N_B1_M1015_g N_VPWR_c_741_n 0.0029264f $X=9.135 $Y=2.4 $X2=0 $Y2=0
cc_509 N_B1_M1020_g N_VPWR_c_741_n 0.00294462f $X=9.585 $Y=2.4 $X2=0 $Y2=0
cc_510 N_B1_M1007_g N_VPWR_c_752_n 0.00460063f $X=8.235 $Y=2.4 $X2=0 $Y2=0
cc_511 N_B1_M1011_g N_VPWR_c_753_n 0.005209f $X=8.685 $Y=2.4 $X2=0 $Y2=0
cc_512 N_B1_M1015_g N_VPWR_c_753_n 0.005209f $X=9.135 $Y=2.4 $X2=0 $Y2=0
cc_513 N_B1_M1020_g N_VPWR_c_754_n 0.005209f $X=9.585 $Y=2.4 $X2=0 $Y2=0
cc_514 N_B1_M1007_g N_VPWR_c_730_n 0.00908665f $X=8.235 $Y=2.4 $X2=0 $Y2=0
cc_515 N_B1_M1011_g N_VPWR_c_730_n 0.0098193f $X=8.685 $Y=2.4 $X2=0 $Y2=0
cc_516 N_B1_M1015_g N_VPWR_c_730_n 0.0098193f $X=9.135 $Y=2.4 $X2=0 $Y2=0
cc_517 N_B1_M1020_g N_VPWR_c_730_n 0.00985524f $X=9.585 $Y=2.4 $X2=0 $Y2=0
cc_518 N_B1_M1007_g N_A_1215_368#_c_991_n 0.00100669f $X=8.235 $Y=2.4 $X2=0
+ $Y2=0
cc_519 N_B1_M1007_g N_A_1215_368#_c_1003_n 0.0140245f $X=8.235 $Y=2.4 $X2=0
+ $Y2=0
cc_520 N_B1_M1011_g N_A_1215_368#_c_1003_n 0.0128923f $X=8.685 $Y=2.4 $X2=0
+ $Y2=0
cc_521 B1 N_A_1215_368#_c_1003_n 0.0410448f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_522 N_B1_c_654_n N_A_1215_368#_c_1003_n 4.89709e-19 $X=9.585 $Y=1.515 $X2=0
+ $Y2=0
cc_523 N_B1_M1007_g N_A_1215_368#_c_992_n 6.56158e-19 $X=8.235 $Y=2.4 $X2=0
+ $Y2=0
cc_524 N_B1_M1011_g N_A_1215_368#_c_992_n 0.011979f $X=8.685 $Y=2.4 $X2=0 $Y2=0
cc_525 N_B1_M1015_g N_A_1215_368#_c_992_n 0.0118161f $X=9.135 $Y=2.4 $X2=0 $Y2=0
cc_526 N_B1_M1020_g N_A_1215_368#_c_992_n 6.35255e-19 $X=9.585 $Y=2.4 $X2=0
+ $Y2=0
cc_527 N_B1_M1015_g N_A_1215_368#_c_1011_n 0.012931f $X=9.135 $Y=2.4 $X2=0 $Y2=0
cc_528 N_B1_M1020_g N_A_1215_368#_c_1011_n 0.012931f $X=9.585 $Y=2.4 $X2=0 $Y2=0
cc_529 B1 N_A_1215_368#_c_1011_n 0.0391869f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_530 N_B1_c_654_n N_A_1215_368#_c_1011_n 4.90767e-19 $X=9.585 $Y=1.515 $X2=0
+ $Y2=0
cc_531 N_B1_M1020_g N_A_1215_368#_c_993_n 8.84614e-19 $X=9.585 $Y=2.4 $X2=0
+ $Y2=0
cc_532 B1 N_A_1215_368#_c_993_n 0.02461f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_533 N_B1_c_654_n N_A_1215_368#_c_993_n 8.7412e-19 $X=9.585 $Y=1.515 $X2=0
+ $Y2=0
cc_534 N_B1_M1015_g N_A_1215_368#_c_994_n 6.30136e-19 $X=9.135 $Y=2.4 $X2=0
+ $Y2=0
cc_535 N_B1_M1020_g N_A_1215_368#_c_994_n 0.0119841f $X=9.585 $Y=2.4 $X2=0 $Y2=0
cc_536 N_B1_M1011_g N_A_1215_368#_c_1020_n 8.84614e-19 $X=8.685 $Y=2.4 $X2=0
+ $Y2=0
cc_537 N_B1_M1015_g N_A_1215_368#_c_1020_n 8.84614e-19 $X=9.135 $Y=2.4 $X2=0
+ $Y2=0
cc_538 B1 N_A_1215_368#_c_1020_n 0.0235495f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_539 N_B1_c_654_n N_A_1215_368#_c_1020_n 5.52302e-19 $X=9.585 $Y=1.515 $X2=0
+ $Y2=0
cc_540 N_B1_M1006_g N_VGND_c_1127_n 0.0104021f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_541 N_B1_M1013_g N_VGND_c_1127_n 0.0104021f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_542 N_B1_M1016_g N_VGND_c_1127_n 5.14838e-19 $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_543 N_B1_M1016_g N_VGND_c_1128_n 0.00418685f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_544 N_B1_M1035_g N_VGND_c_1128_n 0.0133319f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_545 N_B1_M1006_g N_VGND_c_1132_n 0.00383152f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_546 N_B1_M1013_g N_VGND_c_1133_n 0.00383152f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_547 N_B1_M1016_g N_VGND_c_1133_n 0.00434272f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_548 N_B1_M1035_g N_VGND_c_1134_n 0.00383152f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_549 N_B1_M1006_g N_VGND_c_1135_n 0.00757637f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_550 N_B1_M1013_g N_VGND_c_1135_n 0.0075754f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_551 N_B1_M1016_g N_VGND_c_1135_n 0.00820718f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_552 N_B1_M1035_g N_VGND_c_1135_n 0.00761198f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_553 N_B1_M1006_g N_A_857_74#_c_1259_n 3.97481e-19 $X=8.225 $Y=0.74 $X2=0
+ $Y2=0
cc_554 N_B1_M1006_g N_A_857_74#_c_1260_n 0.0130828f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_555 N_B1_M1013_g N_A_857_74#_c_1260_n 0.0131017f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_556 B1 N_A_857_74#_c_1260_n 0.0475521f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_557 N_B1_c_654_n N_A_857_74#_c_1260_n 0.00251192f $X=9.585 $Y=1.515 $X2=0
+ $Y2=0
cc_558 N_B1_M1013_g N_A_857_74#_c_1261_n 3.97481e-19 $X=8.655 $Y=0.74 $X2=0
+ $Y2=0
cc_559 N_B1_M1016_g N_A_857_74#_c_1261_n 0.00922099f $X=9.085 $Y=0.74 $X2=0
+ $Y2=0
cc_560 N_B1_M1035_g N_A_857_74#_c_1261_n 9.78807e-19 $X=9.585 $Y=0.74 $X2=0
+ $Y2=0
cc_561 N_B1_M1016_g N_A_857_74#_c_1262_n 0.0115433f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_562 N_B1_M1035_g N_A_857_74#_c_1262_n 0.0140566f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_563 B1 N_A_857_74#_c_1262_n 0.0721685f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_564 N_B1_c_654_n N_A_857_74#_c_1262_n 0.00832868f $X=9.585 $Y=1.515 $X2=0
+ $Y2=0
cc_565 N_B1_M1035_g N_A_857_74#_c_1263_n 0.00159319f $X=9.585 $Y=0.74 $X2=0
+ $Y2=0
cc_566 N_B1_M1016_g N_A_857_74#_c_1267_n 0.00157732f $X=9.085 $Y=0.74 $X2=0
+ $Y2=0
cc_567 B1 N_A_857_74#_c_1267_n 0.0213626f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_568 N_B1_c_654_n N_A_857_74#_c_1267_n 0.00250705f $X=9.585 $Y=1.515 $X2=0
+ $Y2=0
cc_569 N_VPWR_c_736_n N_Y_c_884_n 0.0338794f $X=3.87 $Y=1.985 $X2=0 $Y2=0
cc_570 N_VPWR_c_737_n N_Y_c_884_n 0.0283117f $X=4.77 $Y=2.305 $X2=0 $Y2=0
cc_571 N_VPWR_c_750_n N_Y_c_884_n 0.0144623f $X=4.685 $Y=3.33 $X2=0 $Y2=0
cc_572 N_VPWR_c_730_n N_Y_c_884_n 0.0118344f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_573 N_VPWR_M1019_s N_Y_c_885_n 0.00165831f $X=4.635 $Y=1.84 $X2=0 $Y2=0
cc_574 N_VPWR_c_737_n N_Y_c_885_n 0.0126919f $X=4.77 $Y=2.305 $X2=0 $Y2=0
cc_575 N_VPWR_c_736_n N_Y_c_886_n 0.00618362f $X=3.87 $Y=1.985 $X2=0 $Y2=0
cc_576 N_VPWR_c_737_n N_Y_c_887_n 0.0268116f $X=4.77 $Y=2.305 $X2=0 $Y2=0
cc_577 N_VPWR_c_738_n N_Y_c_887_n 0.0109793f $X=5.505 $Y=3.33 $X2=0 $Y2=0
cc_578 N_VPWR_c_739_n N_Y_c_887_n 0.0224199f $X=5.67 $Y=2.405 $X2=0 $Y2=0
cc_579 N_VPWR_c_730_n N_Y_c_887_n 0.00901959f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_580 N_VPWR_M1028_s N_Y_c_889_n 0.00321299f $X=5.535 $Y=1.84 $X2=0 $Y2=0
cc_581 N_VPWR_c_739_n N_Y_c_889_n 0.00863845f $X=5.67 $Y=2.405 $X2=0 $Y2=0
cc_582 N_VPWR_M1028_s N_Y_c_890_n 0.00498517f $X=5.535 $Y=1.84 $X2=0 $Y2=0
cc_583 N_VPWR_c_739_n N_Y_c_890_n 0.0125571f $X=5.67 $Y=2.405 $X2=0 $Y2=0
cc_584 N_VPWR_c_739_n N_A_1215_368#_c_988_n 0.0412869f $X=5.67 $Y=2.405 $X2=0
+ $Y2=0
cc_585 N_VPWR_c_752_n N_A_1215_368#_c_989_n 0.0439866f $X=8.295 $Y=3.33 $X2=0
+ $Y2=0
cc_586 N_VPWR_c_730_n N_A_1215_368#_c_989_n 0.0246722f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_587 N_VPWR_c_739_n N_A_1215_368#_c_990_n 0.0129574f $X=5.67 $Y=2.405 $X2=0
+ $Y2=0
cc_588 N_VPWR_c_752_n N_A_1215_368#_c_990_n 0.018997f $X=8.295 $Y=3.33 $X2=0
+ $Y2=0
cc_589 N_VPWR_c_730_n N_A_1215_368#_c_990_n 0.0103026f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_590 N_VPWR_c_740_n N_A_1215_368#_c_991_n 0.0107937f $X=8.46 $Y=2.455 $X2=0
+ $Y2=0
cc_591 N_VPWR_c_752_n N_A_1215_368#_c_991_n 0.0583239f $X=8.295 $Y=3.33 $X2=0
+ $Y2=0
cc_592 N_VPWR_c_730_n N_A_1215_368#_c_991_n 0.0324477f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_593 N_VPWR_M1007_d N_A_1215_368#_c_1003_n 0.00314376f $X=8.325 $Y=1.84 $X2=0
+ $Y2=0
cc_594 N_VPWR_c_740_n N_A_1215_368#_c_1003_n 0.0148589f $X=8.46 $Y=2.455 $X2=0
+ $Y2=0
cc_595 N_VPWR_c_740_n N_A_1215_368#_c_992_n 0.0249143f $X=8.46 $Y=2.455 $X2=0
+ $Y2=0
cc_596 N_VPWR_c_741_n N_A_1215_368#_c_992_n 0.0248868f $X=9.36 $Y=2.455 $X2=0
+ $Y2=0
cc_597 N_VPWR_c_753_n N_A_1215_368#_c_992_n 0.0144623f $X=9.26 $Y=3.33 $X2=0
+ $Y2=0
cc_598 N_VPWR_c_730_n N_A_1215_368#_c_992_n 0.0118344f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_599 N_VPWR_M1015_d N_A_1215_368#_c_1011_n 0.00314376f $X=9.225 $Y=1.84 $X2=0
+ $Y2=0
cc_600 N_VPWR_c_741_n N_A_1215_368#_c_1011_n 0.0126919f $X=9.36 $Y=2.455 $X2=0
+ $Y2=0
cc_601 N_VPWR_c_741_n N_A_1215_368#_c_994_n 0.0254369f $X=9.36 $Y=2.455 $X2=0
+ $Y2=0
cc_602 N_VPWR_c_754_n N_A_1215_368#_c_994_n 0.014549f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_603 N_VPWR_c_730_n N_A_1215_368#_c_994_n 0.0119743f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_604 N_VPWR_c_752_n N_A_1215_368#_c_995_n 0.0143373f $X=8.295 $Y=3.33 $X2=0
+ $Y2=0
cc_605 N_VPWR_c_730_n N_A_1215_368#_c_995_n 0.00777554f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_606 N_Y_c_889_n N_A_1215_368#_M1001_s 0.00537088f $X=6.495 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_607 N_Y_c_940_n N_A_1215_368#_M1004_s 0.00314376f $X=7.395 $Y=2.035 $X2=0
+ $Y2=0
cc_608 N_Y_c_889_n N_A_1215_368#_c_988_n 0.0197787f $X=6.495 $Y=2.035 $X2=0
+ $Y2=0
cc_609 N_Y_M1001_d N_A_1215_368#_c_989_n 0.00165831f $X=6.525 $Y=1.84 $X2=0
+ $Y2=0
cc_610 N_Y_c_944_n N_A_1215_368#_c_989_n 0.0159318f $X=6.66 $Y=2.055 $X2=0 $Y2=0
cc_611 N_Y_c_940_n N_A_1215_368#_c_1051_n 0.0126919f $X=7.395 $Y=2.035 $X2=0
+ $Y2=0
cc_612 N_Y_M1031_d N_A_1215_368#_c_991_n 0.00165831f $X=7.425 $Y=1.84 $X2=0
+ $Y2=0
cc_613 N_Y_c_949_n N_A_1215_368#_c_991_n 0.0159318f $X=7.56 $Y=2.055 $X2=0 $Y2=0
cc_614 N_Y_c_880_n N_A_857_74#_M1018_d 0.00176461f $X=5.545 $Y=1.045 $X2=0 $Y2=0
cc_615 N_Y_c_881_n N_A_857_74#_c_1251_n 0.00756924f $X=5.025 $Y=1.045 $X2=0
+ $Y2=0
cc_616 N_Y_M1009_s N_A_857_74#_c_1252_n 0.00176461f $X=4.72 $Y=0.37 $X2=0 $Y2=0
cc_617 N_Y_c_903_n N_A_857_74#_c_1252_n 0.0157609f $X=4.86 $Y=0.86 $X2=0 $Y2=0
cc_618 N_Y_c_880_n N_A_857_74#_c_1252_n 0.0032855f $X=5.545 $Y=1.045 $X2=0 $Y2=0
cc_619 N_Y_c_880_n N_A_857_74#_c_1318_n 0.0132452f $X=5.545 $Y=1.045 $X2=0 $Y2=0
cc_620 N_Y_M1023_s N_A_857_74#_c_1254_n 0.00176461f $X=5.58 $Y=0.37 $X2=0 $Y2=0
cc_621 N_Y_c_880_n N_A_857_74#_c_1254_n 0.00302054f $X=5.545 $Y=1.045 $X2=0
+ $Y2=0
cc_622 N_Y_c_916_n N_A_857_74#_c_1254_n 0.0166135f $X=5.72 $Y=0.86 $X2=0 $Y2=0
cc_623 N_Y_c_882_n N_A_857_74#_c_1256_n 0.00252526f $X=5.63 $Y=1.8 $X2=0 $Y2=0
cc_624 N_Y_c_883_n N_A_857_74#_c_1256_n 0.00570271f $X=5.715 $Y=1.045 $X2=0
+ $Y2=0
cc_625 N_A_27_74#_c_1055_n N_VGND_M1012_s 0.00176461f $X=1.055 $Y=1.095
+ $X2=-0.19 $Y2=-0.245
cc_626 N_A_27_74#_c_1058_n N_VGND_M1033_s 0.00176461f $X=1.925 $Y=1.095 $X2=0
+ $Y2=0
cc_627 N_A_27_74#_c_1054_n N_VGND_c_1122_n 0.0182902f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_628 N_A_27_74#_c_1055_n N_VGND_c_1122_n 0.0171619f $X=1.055 $Y=1.095 $X2=0
+ $Y2=0
cc_629 N_A_27_74#_c_1057_n N_VGND_c_1122_n 0.0182548f $X=1.145 $Y=0.515 $X2=0
+ $Y2=0
cc_630 N_A_27_74#_c_1057_n N_VGND_c_1123_n 0.0182548f $X=1.145 $Y=0.515 $X2=0
+ $Y2=0
cc_631 N_A_27_74#_c_1058_n N_VGND_c_1123_n 0.0171619f $X=1.925 $Y=1.095 $X2=0
+ $Y2=0
cc_632 N_A_27_74#_c_1060_n N_VGND_c_1123_n 0.0112234f $X=2.095 $Y=0.34 $X2=0
+ $Y2=0
cc_633 N_A_27_74#_c_1059_n N_VGND_c_1124_n 0.0428729f $X=2.775 $Y=0.34 $X2=0
+ $Y2=0
cc_634 N_A_27_74#_c_1060_n N_VGND_c_1124_n 0.0121867f $X=2.095 $Y=0.34 $X2=0
+ $Y2=0
cc_635 N_A_27_74#_c_1061_n N_VGND_c_1124_n 0.0607975f $X=3.785 $Y=0.34 $X2=0
+ $Y2=0
cc_636 N_A_27_74#_c_1064_n N_VGND_c_1124_n 0.023391f $X=2.94 $Y=0.34 $X2=0 $Y2=0
cc_637 N_A_27_74#_c_1054_n N_VGND_c_1129_n 0.011066f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_638 N_A_27_74#_c_1057_n N_VGND_c_1130_n 0.00794252f $X=1.145 $Y=0.515 $X2=0
+ $Y2=0
cc_639 N_A_27_74#_c_1054_n N_VGND_c_1135_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_640 N_A_27_74#_c_1057_n N_VGND_c_1135_n 0.00657413f $X=1.145 $Y=0.515 $X2=0
+ $Y2=0
cc_641 N_A_27_74#_c_1059_n N_VGND_c_1135_n 0.0241933f $X=2.775 $Y=0.34 $X2=0
+ $Y2=0
cc_642 N_A_27_74#_c_1060_n N_VGND_c_1135_n 0.00660921f $X=2.095 $Y=0.34 $X2=0
+ $Y2=0
cc_643 N_A_27_74#_c_1061_n N_VGND_c_1135_n 0.0339133f $X=3.785 $Y=0.34 $X2=0
+ $Y2=0
cc_644 N_A_27_74#_c_1064_n N_VGND_c_1135_n 0.0127797f $X=2.94 $Y=0.34 $X2=0
+ $Y2=0
cc_645 N_A_27_74#_c_1062_n N_A_857_74#_c_1251_n 0.0455088f $X=3.87 $Y=0.515
+ $X2=0 $Y2=0
cc_646 N_A_27_74#_c_1061_n N_A_857_74#_c_1253_n 0.0128665f $X=3.785 $Y=0.34
+ $X2=0 $Y2=0
cc_647 N_VGND_c_1124_n N_A_857_74#_c_1252_n 0.043517f $X=6.415 $Y=0 $X2=0 $Y2=0
cc_648 N_VGND_c_1135_n N_A_857_74#_c_1252_n 0.0245693f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_649 N_VGND_c_1124_n N_A_857_74#_c_1253_n 0.0179217f $X=6.415 $Y=0 $X2=0 $Y2=0
cc_650 N_VGND_c_1135_n N_A_857_74#_c_1253_n 0.00971942f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_651 N_VGND_c_1124_n N_A_857_74#_c_1254_n 0.0557038f $X=6.415 $Y=0 $X2=0 $Y2=0
cc_652 N_VGND_c_1125_n N_A_857_74#_c_1254_n 0.0112234f $X=6.58 $Y=0.65 $X2=0
+ $Y2=0
cc_653 N_VGND_c_1135_n N_A_857_74#_c_1254_n 0.0311785f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_654 N_VGND_M1002_d N_A_857_74#_c_1255_n 0.00256964f $X=6.44 $Y=0.37 $X2=0
+ $Y2=0
cc_655 N_VGND_c_1125_n N_A_857_74#_c_1255_n 0.0201026f $X=6.58 $Y=0.65 $X2=0
+ $Y2=0
cc_656 N_VGND_c_1125_n N_A_857_74#_c_1257_n 0.018051f $X=6.58 $Y=0.65 $X2=0
+ $Y2=0
cc_657 N_VGND_c_1126_n N_A_857_74#_c_1257_n 0.0179318f $X=7.51 $Y=0.65 $X2=0
+ $Y2=0
cc_658 N_VGND_c_1131_n N_A_857_74#_c_1257_n 0.0109942f $X=7.345 $Y=0 $X2=0 $Y2=0
cc_659 N_VGND_c_1135_n N_A_857_74#_c_1257_n 0.00904371f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_660 N_VGND_M1025_d N_A_857_74#_c_1258_n 0.00256964f $X=7.37 $Y=0.37 $X2=0
+ $Y2=0
cc_661 N_VGND_c_1126_n N_A_857_74#_c_1258_n 0.0201026f $X=7.51 $Y=0.65 $X2=0
+ $Y2=0
cc_662 N_VGND_c_1126_n N_A_857_74#_c_1259_n 0.018051f $X=7.51 $Y=0.65 $X2=0
+ $Y2=0
cc_663 N_VGND_c_1127_n N_A_857_74#_c_1259_n 0.0179318f $X=8.44 $Y=0.65 $X2=0
+ $Y2=0
cc_664 N_VGND_c_1132_n N_A_857_74#_c_1259_n 0.0109942f $X=8.275 $Y=0 $X2=0 $Y2=0
cc_665 N_VGND_c_1135_n N_A_857_74#_c_1259_n 0.00904371f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_666 N_VGND_M1006_s N_A_857_74#_c_1260_n 0.00180746f $X=8.3 $Y=0.37 $X2=0
+ $Y2=0
cc_667 N_VGND_c_1127_n N_A_857_74#_c_1260_n 0.0163515f $X=8.44 $Y=0.65 $X2=0
+ $Y2=0
cc_668 N_VGND_c_1127_n N_A_857_74#_c_1261_n 0.0179318f $X=8.44 $Y=0.65 $X2=0
+ $Y2=0
cc_669 N_VGND_c_1128_n N_A_857_74#_c_1261_n 0.018051f $X=9.37 $Y=0.65 $X2=0
+ $Y2=0
cc_670 N_VGND_c_1133_n N_A_857_74#_c_1261_n 0.0109942f $X=9.205 $Y=0 $X2=0 $Y2=0
cc_671 N_VGND_c_1135_n N_A_857_74#_c_1261_n 0.00904371f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_672 N_VGND_M1016_s N_A_857_74#_c_1262_n 0.00256964f $X=9.16 $Y=0.37 $X2=0
+ $Y2=0
cc_673 N_VGND_c_1128_n N_A_857_74#_c_1262_n 0.0201026f $X=9.37 $Y=0.65 $X2=0
+ $Y2=0
cc_674 N_VGND_c_1128_n N_A_857_74#_c_1263_n 0.0179318f $X=9.37 $Y=0.65 $X2=0
+ $Y2=0
cc_675 N_VGND_c_1134_n N_A_857_74#_c_1263_n 0.011066f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_676 N_VGND_c_1135_n N_A_857_74#_c_1263_n 0.00915947f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_677 N_VGND_c_1124_n N_A_857_74#_c_1264_n 0.0119713f $X=6.415 $Y=0 $X2=0 $Y2=0
cc_678 N_VGND_c_1135_n N_A_857_74#_c_1264_n 0.00656877f $X=9.84 $Y=0 $X2=0 $Y2=0

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__nor4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__nor4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.310000 1.350000 7.075000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.860000 1.350000 6.115000 1.635000 ;
        RECT 5.405000 1.635000 6.115000 1.780000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.470000 1.315000 1.800000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495000 1.470000 1.825000 1.800000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  1.164500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.890000 0.350000 3.220000 0.670000 ;
        RECT 2.890000 0.670000 4.285000 0.840000 ;
        RECT 2.975000 1.850000 4.285000 2.020000 ;
        RECT 2.975000 2.020000 3.225000 2.735000 ;
        RECT 3.955000 0.350000 4.285000 0.670000 ;
        RECT 3.955000 0.840000 4.285000 1.010000 ;
        RECT 3.955000 1.010000 6.575000 1.180000 ;
        RECT 4.115000 1.180000 4.285000 1.550000 ;
        RECT 4.115000 1.550000 4.675000 1.780000 ;
        RECT 4.115000 1.780000 4.285000 1.850000 ;
        RECT 4.965000 0.350000 5.215000 1.010000 ;
        RECT 6.325000 0.350000 6.575000 1.010000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.115000  1.130000 0.815000 1.300000 ;
      RECT 0.115000  1.300000 0.285000 1.970000 ;
      RECT 0.115000  1.970000 0.445000 2.980000 ;
      RECT 0.485000  0.360000 0.815000 0.710000 ;
      RECT 0.485000  0.710000 2.665000 0.880000 ;
      RECT 0.485000  0.880000 0.815000 1.130000 ;
      RECT 0.615000  1.970000 1.715000 3.245000 ;
      RECT 0.990000  0.085000 1.515000 0.540000 ;
      RECT 1.620000  1.050000 2.325000 1.300000 ;
      RECT 1.885000  1.970000 2.325000 2.140000 ;
      RECT 1.885000  2.140000 2.215000 2.980000 ;
      RECT 2.155000  1.300000 2.325000 1.350000 ;
      RECT 2.155000  1.350000 3.165000 1.680000 ;
      RECT 2.155000  1.680000 2.325000 1.970000 ;
      RECT 2.195000  0.085000 2.710000 0.540000 ;
      RECT 2.495000  0.880000 2.665000 1.010000 ;
      RECT 2.495000  1.010000 3.785000 1.180000 ;
      RECT 2.495000  1.850000 2.775000 2.905000 ;
      RECT 2.495000  2.905000 3.725000 3.075000 ;
      RECT 3.395000  2.190000 4.675000 2.360000 ;
      RECT 3.395000  2.360000 3.725000 2.905000 ;
      RECT 3.400000  0.085000 3.775000 0.500000 ;
      RECT 3.615000  1.180000 3.785000 1.350000 ;
      RECT 3.615000  1.350000 3.945000 1.680000 ;
      RECT 3.895000  2.530000 4.175000 2.905000 ;
      RECT 3.895000  2.905000 5.685000 3.075000 ;
      RECT 4.345000  2.360000 4.675000 2.735000 ;
      RECT 4.455000  0.085000 4.785000 0.840000 ;
      RECT 4.905000  1.820000 5.155000 1.950000 ;
      RECT 4.905000  1.950000 7.085000 2.120000 ;
      RECT 4.905000  2.120000 5.155000 2.735000 ;
      RECT 5.355000  2.290000 5.685000 2.905000 ;
      RECT 5.385000  0.085000 6.155000 0.840000 ;
      RECT 5.855000  2.120000 6.185000 2.980000 ;
      RECT 6.385000  2.290000 6.555000 3.245000 ;
      RECT 6.755000  0.085000 7.085000 1.130000 ;
      RECT 6.755000  2.120000 7.085000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_ms__nor4bb_2
END LIBRARY

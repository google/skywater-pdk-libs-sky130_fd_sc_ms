* File: sky130_fd_sc_ms__or3b_4.pex.spice
* Created: Fri Aug 28 18:08:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__OR3B_4%C_N 1 3 8 10 12 19 20
c34 3 0 1.18961e-19 $X=0.5 $Y=2.46
r35 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.61
+ $Y=0.405 $X2=0.61 $Y2=0.405
r36 17 19 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=0.515 $Y=0.405
+ $X2=0.61 $Y2=0.405
r37 15 20 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=0.27 $Y=0.447
+ $X2=0.61 $Y2=0.447
r38 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=0.405 $X2=0.27 $Y2=0.405
r39 12 17 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.44 $Y=0.405
+ $X2=0.515 $Y2=0.405
r40 12 14 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=0.44 $Y=0.405
+ $X2=0.27 $Y2=0.405
r41 10 15 0.898008 $w=3.83e-07 $l=3e-08 $layer=LI1_cond $X=0.24 $Y=0.447
+ $X2=0.27 $Y2=0.447
r42 8 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.515 $Y=1 $X2=0.515
+ $Y2=1.395
r43 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=0.57
+ $X2=0.515 $Y2=0.405
r44 5 8 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.515 $Y=0.57
+ $X2=0.515 $Y2=1
r45 1 9 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.5 $Y=1.485 $X2=0.5
+ $Y2=1.395
r46 1 3 378.992 $w=1.8e-07 $l=9.75e-07 $layer=POLY_cond $X=0.5 $Y=1.485 $X2=0.5
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__OR3B_4%A 3 7 10 14 15 17 18 19 25 27
c93 10 0 7.15249e-20 $X=3.405 $Y=2.46
r94 25 28 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.45 $Y=1.385
+ $X2=3.45 $Y2=1.55
r95 25 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.45 $Y=1.385
+ $X2=3.45 $Y2=1.22
r96 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.45
+ $Y=1.385 $X2=3.45 $Y2=1.385
r97 19 26 12.9453 $w=3.11e-07 $l=3.3e-07 $layer=LI1_cond $X=3.12 $Y=1.35
+ $X2=3.45 $Y2=1.35
r98 17 19 7.00102 $w=3.11e-07 $l=1.62635e-07 $layer=LI1_cond $X=3.005 $Y=1.235
+ $X2=3.12 $Y2=1.35
r99 17 18 122.326 $w=1.68e-07 $l=1.875e-06 $layer=LI1_cond $X=3.005 $Y=1.235
+ $X2=1.13 $Y2=1.235
r100 15 23 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.595
+ $X2=0.965 $Y2=1.76
r101 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.595 $X2=0.965 $Y2=1.595
r102 12 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.965 $Y=1.32
+ $X2=1.13 $Y2=1.235
r103 12 14 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.965 $Y=1.32
+ $X2=0.965 $Y2=1.595
r104 10 28 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=3.405 $Y=2.46
+ $X2=3.405 $Y2=1.55
r105 7 27 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.39 $Y=0.74 $X2=3.39
+ $Y2=1.22
r106 3 23 272.097 $w=1.8e-07 $l=7e-07 $layer=POLY_cond $X=1.01 $Y=2.46 $X2=1.01
+ $Y2=1.76
.ends

.subckt PM_SKY130_FD_SC_MS__OR3B_4%B 3 7 11 13 14 15 21 26 27 32 43
c67 11 0 1.44963e-19 $X=2.96 $Y=0.74
c68 7 0 1.95106e-19 $X=2.895 $Y=2.46
c69 3 0 1.78721e-19 $X=1.46 $Y=2.46
r70 32 43 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=1.68 $Y=1.675
+ $X2=1.67 $Y2=1.675
r71 26 29 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.91 $Y=1.635
+ $X2=2.91 $Y2=1.8
r72 26 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.91 $Y=1.635
+ $X2=2.91 $Y2=1.47
r73 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.91
+ $Y=1.635 $X2=2.91 $Y2=1.635
r74 21 24 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.505 $Y=1.635
+ $X2=1.505 $Y2=1.8
r75 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.505
+ $Y=1.635 $X2=1.505 $Y2=1.635
r76 15 27 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=2.64 $Y=1.675
+ $X2=2.91 $Y2=1.675
r77 14 15 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.675
+ $X2=2.64 $Y2=1.675
r78 13 43 1.87799 $w=3.08e-07 $l=3.8e-08 $layer=LI1_cond $X=1.632 $Y=1.645
+ $X2=1.67 $Y2=1.645
r79 13 22 4.7213 $w=3.08e-07 $l=1.27e-07 $layer=LI1_cond $X=1.632 $Y=1.645
+ $X2=1.505 $Y2=1.645
r80 13 14 20.4213 $w=2.48e-07 $l=4.43e-07 $layer=LI1_cond $X=1.717 $Y=1.675
+ $X2=2.16 $Y2=1.675
r81 13 32 1.70562 $w=2.48e-07 $l=3.7e-08 $layer=LI1_cond $X=1.717 $Y=1.675
+ $X2=1.68 $Y2=1.675
r82 11 28 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.96 $Y=0.74
+ $X2=2.96 $Y2=1.47
r83 7 29 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.895 $Y=2.46
+ $X2=2.895 $Y2=1.8
r84 3 24 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.46 $Y=2.46 $X2=1.46
+ $Y2=1.8
.ends

.subckt PM_SKY130_FD_SC_MS__OR3B_4%A_27_392# 1 2 8 11 13 17 19 21 22 23 27 30 34
+ 35 38 39 41
r88 39 44 88.9594 $w=4.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.805 $Y=0.475
+ $X2=1.805 $Y2=0.98
r89 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.745
+ $Y=0.475 $X2=1.745 $Y2=0.475
r90 36 38 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.745 $Y=0.81
+ $X2=1.745 $Y2=0.475
r91 34 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.58 $Y=0.895
+ $X2=1.745 $Y2=0.81
r92 34 35 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=1.58 $Y=0.895
+ $X2=0.465 $Y2=0.895
r93 30 32 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=0.235 $Y=2.105
+ $X2=0.235 $Y2=2.815
r94 30 41 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=0.235 $Y=2.105
+ $X2=0.235 $Y2=1.34
r95 25 41 6.76842 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=0.287 $Y=1.163
+ $X2=0.287 $Y2=1.34
r96 25 27 2.85676 $w=3.53e-07 $l=8.8e-08 $layer=LI1_cond $X=0.287 $Y=1.163
+ $X2=0.287 $Y2=1.075
r97 24 35 7.97992 $w=1.7e-07 $l=2.16365e-07 $layer=LI1_cond $X=0.287 $Y=0.98
+ $X2=0.465 $Y2=0.895
r98 24 27 3.084 $w=3.53e-07 $l=9.5e-08 $layer=LI1_cond $X=0.287 $Y=0.98
+ $X2=0.287 $Y2=1.075
r99 19 23 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=2.46 $Y=1.185
+ $X2=2.445 $Y2=1.26
r100 19 21 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.46 $Y=1.185
+ $X2=2.46 $Y2=0.74
r101 15 23 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=2.445 $Y=1.335
+ $X2=2.445 $Y2=1.26
r102 15 17 437.298 $w=1.8e-07 $l=1.125e-06 $layer=POLY_cond $X=2.445 $Y=1.335
+ $X2=2.445 $Y2=2.46
r103 14 22 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.06 $Y=1.26 $X2=1.97
+ $Y2=1.26
r104 13 23 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.355 $Y=1.26
+ $X2=2.445 $Y2=1.26
r105 13 14 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=2.355 $Y=1.26
+ $X2=2.06 $Y2=1.26
r106 9 22 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=1.97 $Y=1.335
+ $X2=1.97 $Y2=1.26
r107 9 11 437.298 $w=1.8e-07 $l=1.125e-06 $layer=POLY_cond $X=1.97 $Y=1.335
+ $X2=1.97 $Y2=2.46
r108 8 22 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=1.955 $Y=1.185
+ $X2=1.97 $Y2=1.26
r109 8 44 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=1.955 $Y=1.185
+ $X2=1.955 $Y2=0.98
r110 2 32 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.275 $Y2=2.815
r111 2 30 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.275 $Y2=2.105
r112 1 27 182 $w=1.7e-07 $l=4.61844e-07 $layer=licon1_NDIFF $count=1 $X=0.155
+ $Y=0.68 $X2=0.3 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_MS__OR3B_4%A_412_392# 1 2 3 12 16 20 24 28 32 36 40 44
+ 46 48 49 52 54 57 59 65 71 73 74 84
c159 52 0 1.44963e-19 $X=3.175 $Y=0.515
c160 16 0 1.10433e-19 $X=3.915 $Y=2.4
r161 81 82 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.815 $Y=1.465
+ $X2=4.835 $Y2=1.465
r162 80 81 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=4.365 $Y=1.465
+ $X2=4.815 $Y2=1.465
r163 79 80 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=4.355 $Y=1.465
+ $X2=4.365 $Y2=1.465
r164 75 77 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.9 $Y=1.465
+ $X2=3.915 $Y2=1.465
r165 69 71 10.0544 $w=2.18e-07 $l=1.8e-07 $layer=LI1_cond $X=2.205 $Y=2.08
+ $X2=2.385 $Y2=2.08
r166 66 84 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=5.01 $Y=1.465
+ $X2=5.265 $Y2=1.465
r167 66 82 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=5.01 $Y=1.465
+ $X2=4.835 $Y2=1.465
r168 65 66 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.01
+ $Y=1.465 $X2=5.01 $Y2=1.465
r169 63 79 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=3.99 $Y=1.465
+ $X2=4.355 $Y2=1.465
r170 63 77 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.99 $Y=1.465
+ $X2=3.915 $Y2=1.465
r171 62 65 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=3.99 $Y=1.465
+ $X2=5.01 $Y2=1.465
r172 62 63 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.99
+ $Y=1.465 $X2=3.99 $Y2=1.465
r173 60 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.885 $Y=1.465
+ $X2=3.8 $Y2=1.465
r174 60 62 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.885 $Y=1.465
+ $X2=3.99 $Y2=1.465
r175 58 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.8 $Y=1.63 $X2=3.8
+ $Y2=1.465
r176 58 59 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.8 $Y=1.63 $X2=3.8
+ $Y2=1.97
r177 57 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.8 $Y=1.3 $X2=3.8
+ $Y2=1.465
r178 56 57 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.8 $Y=0.98 $X2=3.8
+ $Y2=1.3
r179 55 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.34 $Y=0.895
+ $X2=3.215 $Y2=0.895
r180 54 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.715 $Y=0.895
+ $X2=3.8 $Y2=0.98
r181 54 55 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.715 $Y=0.895
+ $X2=3.34 $Y2=0.895
r182 50 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=0.81
+ $X2=3.215 $Y2=0.895
r183 50 52 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.215 $Y=0.81
+ $X2=3.215 $Y2=0.515
r184 48 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.09 $Y=0.895
+ $X2=3.215 $Y2=0.895
r185 48 49 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.09 $Y=0.895
+ $X2=2.41 $Y2=0.895
r186 46 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.715 $Y=2.055
+ $X2=3.8 $Y2=1.97
r187 46 71 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=3.715 $Y=2.055
+ $X2=2.385 $Y2=2.055
r188 42 49 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.245 $Y=0.81
+ $X2=2.41 $Y2=0.895
r189 42 44 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.245 $Y=0.81
+ $X2=2.245 $Y2=0.515
r190 38 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.265 $Y=1.3
+ $X2=5.265 $Y2=1.465
r191 38 40 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.265 $Y=1.3
+ $X2=5.265 $Y2=0.74
r192 34 84 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.265 $Y=1.63
+ $X2=5.265 $Y2=1.465
r193 34 36 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=5.265 $Y=1.63
+ $X2=5.265 $Y2=2.4
r194 30 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.835 $Y=1.3
+ $X2=4.835 $Y2=1.465
r195 30 32 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.835 $Y=1.3
+ $X2=4.835 $Y2=0.74
r196 26 81 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.815 $Y=1.63
+ $X2=4.815 $Y2=1.465
r197 26 28 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.815 $Y=1.63
+ $X2=4.815 $Y2=2.4
r198 22 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.355 $Y=1.3
+ $X2=4.355 $Y2=1.465
r199 22 24 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=4.355 $Y=1.3
+ $X2=4.355 $Y2=0.74
r200 18 80 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.365 $Y=1.63
+ $X2=4.365 $Y2=1.465
r201 18 20 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=4.365 $Y=1.63
+ $X2=4.365 $Y2=2.4
r202 14 77 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.915 $Y=1.63
+ $X2=3.915 $Y2=1.465
r203 14 16 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=3.915 $Y=1.63
+ $X2=3.915 $Y2=2.4
r204 10 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.9 $Y=1.3 $X2=3.9
+ $Y2=1.465
r205 10 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.9 $Y=1.3 $X2=3.9
+ $Y2=0.74
r206 3 69 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.06
+ $Y=1.96 $X2=2.205 $Y2=2.105
r207 2 73 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=3.035
+ $Y=0.37 $X2=3.175 $Y2=0.895
r208 2 52 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.035
+ $Y=0.37 $X2=3.175 $Y2=0.515
r209 1 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.105
+ $Y=0.37 $X2=2.245 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR3B_4%VPWR 1 2 3 4 15 21 25 27 29 31 33 38 46 51 57
+ 60 63 67
r74 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r75 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r76 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r77 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r78 55 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r79 55 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r80 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r81 52 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.675 $Y=3.33
+ $X2=4.55 $Y2=3.33
r82 52 54 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.675 $Y=3.33
+ $X2=5.04 $Y2=3.33
r83 51 66 4.02656 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=5.405 $Y=3.33
+ $X2=5.582 $Y2=3.33
r84 51 54 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.405 $Y=3.33
+ $X2=5.04 $Y2=3.33
r85 50 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r86 50 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r87 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r88 47 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.835 $Y=3.33
+ $X2=3.67 $Y2=3.33
r89 47 49 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.835 $Y=3.33
+ $X2=4.08 $Y2=3.33
r90 46 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.55 $Y2=3.33
r91 46 49 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.425 $Y=3.33
+ $X2=4.08 $Y2=3.33
r92 45 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r93 44 45 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r94 42 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r95 41 44 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r96 41 42 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r97 39 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=3.33
+ $X2=0.725 $Y2=3.33
r98 39 41 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.89 $Y=3.33 $X2=1.2
+ $Y2=3.33
r99 38 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.505 $Y=3.33
+ $X2=3.67 $Y2=3.33
r100 38 44 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.505 $Y=3.33
+ $X2=3.12 $Y2=3.33
r101 36 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r102 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r103 33 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.725 $Y2=3.33
r104 33 35 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.24 $Y2=3.33
r105 31 45 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r106 31 42 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=1.2 $Y2=3.33
r107 27 66 3.1166 $w=2.5e-07 $l=1.07912e-07 $layer=LI1_cond $X=5.53 $Y=3.245
+ $X2=5.582 $Y2=3.33
r108 27 29 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=5.53 $Y=3.245
+ $X2=5.53 $Y2=2.305
r109 23 63 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.55 $Y=3.245
+ $X2=4.55 $Y2=3.33
r110 23 25 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=4.55 $Y=3.245
+ $X2=4.55 $Y2=2.305
r111 19 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=3.245
+ $X2=3.67 $Y2=3.33
r112 19 21 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=3.67 $Y=3.245
+ $X2=3.67 $Y2=2.475
r113 15 18 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.725 $Y=2.105
+ $X2=0.725 $Y2=2.815
r114 13 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=3.33
r115 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=2.815
r116 4 29 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=5.355
+ $Y=1.84 $X2=5.49 $Y2=2.305
r117 3 25 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=4.455
+ $Y=1.84 $X2=4.59 $Y2=2.305
r118 2 21 300 $w=1.7e-07 $l=5.96112e-07 $layer=licon1_PDIFF $count=2 $X=3.495
+ $Y=1.96 $X2=3.67 $Y2=2.475
r119 1 18 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.96 $X2=0.725 $Y2=2.815
r120 1 15 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.96 $X2=0.725 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_MS__OR3B_4%A_220_392# 1 2 9 13 15 19 21
c38 21 0 3.0554e-19 $X=3.17 $Y=2.475
c39 13 0 1.18961e-19 $X=1.235 $Y=2.815
r40 16 19 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.4 $Y=2.445
+ $X2=1.235 $Y2=2.445
r41 15 21 4.91858 $w=1.7e-07 $l=1.77059e-07 $layer=LI1_cond $X=3.005 $Y=2.445
+ $X2=3.17 $Y2=2.42
r42 15 16 104.711 $w=1.68e-07 $l=1.605e-06 $layer=LI1_cond $X=3.005 $Y=2.445
+ $X2=1.4 $Y2=2.445
r43 11 19 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=2.53
+ $X2=1.235 $Y2=2.445
r44 11 13 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.235 $Y=2.53
+ $X2=1.235 $Y2=2.815
r45 7 19 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=2.36
+ $X2=1.235 $Y2=2.445
r46 7 9 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=1.235 $Y=2.36
+ $X2=1.235 $Y2=2.135
r47 2 21 300 $w=1.7e-07 $l=6.00417e-07 $layer=licon1_PDIFF $count=2 $X=2.985
+ $Y=1.96 $X2=3.17 $Y2=2.475
r48 1 13 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.1
+ $Y=1.96 $X2=1.235 $Y2=2.815
r49 1 9 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.1
+ $Y=1.96 $X2=1.235 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_MS__OR3B_4%A_310_392# 1 2 11
c13 11 0 2.50246e-19 $X=2.67 $Y=2.8
r14 8 11 38.0718 $w=2.78e-07 $l=9.25e-07 $layer=LI1_cond $X=1.745 $Y=2.84
+ $X2=2.67 $Y2=2.84
r15 2 11 600 $w=1.7e-07 $l=9.04986e-07 $layer=licon1_PDIFF $count=1 $X=2.535
+ $Y=1.96 $X2=2.67 $Y2=2.8
r16 1 8 600 $w=1.7e-07 $l=9.32416e-07 $layer=licon1_PDIFF $count=1 $X=1.55
+ $Y=1.96 $X2=1.745 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_MS__OR3B_4%X 1 2 3 4 15 19 23 24 25 26 29 35 37 39 41 42
+ 45 46
r80 45 46 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=5.52 $Y=1.295
+ $X2=5.52 $Y2=1.665
r81 44 46 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=5.52 $Y=1.8
+ $X2=5.52 $Y2=1.665
r82 43 45 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.52 $Y=1.13
+ $X2=5.52 $Y2=1.295
r83 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.205 $Y=1.885
+ $X2=5.04 $Y2=1.885
r84 39 44 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=5.405 $Y=1.885
+ $X2=5.52 $Y2=1.8
r85 39 40 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=5.405 $Y=1.885
+ $X2=5.205 $Y2=1.885
r86 38 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.135 $Y=1.045
+ $X2=5.01 $Y2=1.045
r87 37 43 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=5.405 $Y=1.045
+ $X2=5.52 $Y2=1.13
r88 37 38 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.405 $Y=1.045
+ $X2=5.135 $Y2=1.045
r89 33 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.01 $Y=0.96
+ $X2=5.01 $Y2=1.045
r90 33 35 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=5.01 $Y=0.96
+ $X2=5.01 $Y2=0.515
r91 29 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=5.04 $Y=1.985
+ $X2=5.04 $Y2=2.815
r92 27 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.04 $Y=1.97 $X2=5.04
+ $Y2=1.885
r93 27 29 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.04 $Y=1.97
+ $X2=5.04 $Y2=1.985
r94 25 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.875 $Y=1.885
+ $X2=5.04 $Y2=1.885
r95 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.875 $Y=1.885
+ $X2=4.225 $Y2=1.885
r96 23 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.885 $Y=1.045
+ $X2=5.01 $Y2=1.045
r97 23 24 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=4.885 $Y=1.045
+ $X2=4.225 $Y2=1.045
r98 19 21 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.14 $Y=1.985
+ $X2=4.14 $Y2=2.815
r99 17 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.14 $Y=1.97
+ $X2=4.225 $Y2=1.885
r100 17 19 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=4.14 $Y=1.97
+ $X2=4.14 $Y2=1.985
r101 13 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.14 $Y=0.96
+ $X2=4.225 $Y2=1.045
r102 13 15 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=4.14 $Y=0.96
+ $X2=4.14 $Y2=0.515
r103 4 31 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.905
+ $Y=1.84 $X2=5.04 $Y2=2.815
r104 4 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.905
+ $Y=1.84 $X2=5.04 $Y2=1.985
r105 3 21 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.84 $X2=4.14 $Y2=2.815
r106 3 19 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.84 $X2=4.14 $Y2=1.985
r107 2 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.91
+ $Y=0.37 $X2=5.05 $Y2=0.515
r108 1 15 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=3.975
+ $Y=0.37 $X2=4.14 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR3B_4%VGND 1 2 3 4 5 18 22 26 30 32 34 36 38 43 48
+ 53 58 64 67 70 73 77
r87 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r88 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r89 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r90 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r91 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r92 62 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r93 62 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r94 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r95 59 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.655 $Y=0 $X2=4.53
+ $Y2=0
r96 59 61 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.655 $Y=0 $X2=5.04
+ $Y2=0
r97 58 76 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.537
+ $Y2=0
r98 58 61 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.04
+ $Y2=0
r99 57 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r100 57 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r101 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r102 54 70 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.85 $Y=0 $X2=3.68
+ $Y2=0
r103 54 56 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.85 $Y=0 $X2=4.08
+ $Y2=0
r104 53 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.405 $Y=0 $X2=4.53
+ $Y2=0
r105 53 56 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.405 $Y=0
+ $X2=4.08 $Y2=0
r106 52 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r107 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r108 49 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.91 $Y=0 $X2=2.745
+ $Y2=0
r109 49 51 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.91 $Y=0 $X2=3.12
+ $Y2=0
r110 48 70 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.51 $Y=0 $X2=3.68
+ $Y2=0
r111 48 51 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.51 $Y=0 $X2=3.12
+ $Y2=0
r112 47 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r113 47 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r114 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r115 44 64 10.8012 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.177
+ $Y2=0
r116 44 46 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.41 $Y=0 $X2=1.68
+ $Y2=0
r117 43 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.58 $Y=0 $X2=2.745
+ $Y2=0
r118 43 46 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=2.58 $Y=0 $X2=1.68
+ $Y2=0
r119 41 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r120 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r121 38 64 10.8012 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=0.945 $Y=0
+ $X2=1.177 $Y2=0
r122 38 40 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.945 $Y=0
+ $X2=0.72 $Y2=0
r123 36 52 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=3.12 $Y2=0
r124 36 68 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=2.64 $Y2=0
r125 32 76 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.537 $Y2=0
r126 32 34 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0.625
r127 28 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.53 $Y=0.085
+ $X2=4.53 $Y2=0
r128 28 30 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=4.53 $Y=0.085
+ $X2=4.53 $Y2=0.595
r129 24 70 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.68 $Y=0.085
+ $X2=3.68 $Y2=0
r130 24 26 14.575 $w=3.38e-07 $l=4.3e-07 $layer=LI1_cond $X=3.68 $Y=0.085
+ $X2=3.68 $Y2=0.515
r131 20 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.745 $Y=0.085
+ $X2=2.745 $Y2=0
r132 20 22 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.745 $Y=0.085
+ $X2=2.745 $Y2=0.535
r133 16 64 1.88438 $w=4.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.177 $Y=0.085
+ $X2=1.177 $Y2=0
r134 16 18 10.0316 $w=4.63e-07 $l=3.9e-07 $layer=LI1_cond $X=1.177 $Y=0.085
+ $X2=1.177 $Y2=0.475
r135 5 34 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=5.34
+ $Y=0.37 $X2=5.48 $Y2=0.625
r136 4 30 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.37 $X2=4.57 $Y2=0.595
r137 3 26 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=3.465
+ $Y=0.37 $X2=3.68 $Y2=0.515
r138 2 22 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=2.535
+ $Y=0.37 $X2=2.745 $Y2=0.535
r139 1 18 182 $w=1.7e-07 $l=6.79816e-07 $layer=licon1_NDIFF $count=1 $X=0.59
+ $Y=0.68 $X2=1.175 $Y2=0.475
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__dfrtn_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__dfrtn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.960000 0.370000 2.150000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.517000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.590000 0.440000 10.955000 1.150000 ;
        RECT 10.605000 1.820000 10.955000 2.980000 ;
        RECT 10.785000 1.150000 10.955000 1.820000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.415800 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.880000 1.350000 1.285000 1.780000 ;
        RECT 4.820000 1.470000 5.155000 1.800000 ;
        RECT 8.285000 1.465000 8.710000 1.795000 ;
      LAYER mcon ;
        RECT 1.115000 1.580000 1.285000 1.750000 ;
        RECT 4.955000 1.580000 5.125000 1.750000 ;
        RECT 8.315000 1.580000 8.485000 1.750000 ;
      LAYER met1 ;
        RECT 1.055000 1.550000 1.345000 1.595000 ;
        RECT 1.055000 1.595000 8.545000 1.735000 ;
        RECT 1.055000 1.735000 1.345000 1.780000 ;
        RECT 4.895000 1.550000 5.185000 1.595000 ;
        RECT 4.895000 1.735000 5.185000 1.780000 ;
        RECT 8.255000 1.550000 8.545000 1.595000 ;
        RECT 8.255000 1.735000 8.545000 1.780000 ;
    END
  END RESET_B
  PIN CLK_N
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.455000 1.180000 1.765000 1.550000 ;
        RECT 1.515000 1.550000 1.765000 1.575000 ;
    END
  END CLK_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 11.040000 0.085000 ;
        RECT  1.045000  0.085000  1.245000 0.810000 ;
        RECT  2.035000  0.085000  2.365000 0.640000 ;
        RECT  5.025000  0.085000  5.355000 0.620000 ;
        RECT  8.115000  0.085000  8.555000 0.905000 ;
        RECT 10.160000  0.085000 10.410000 1.130000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 11.040000 3.415000 ;
        RECT  0.110000 2.520000  0.440000 3.245000 ;
        RECT  1.060000 2.550000  1.390000 3.245000 ;
        RECT  2.045000 2.550000  2.375000 3.245000 ;
        RECT  4.490000 2.360000  4.820000 3.245000 ;
        RECT  5.490000 2.360000  5.820000 3.245000 ;
        RECT  8.140000 2.520000  8.470000 3.245000 ;
        RECT  9.210000 2.520000  9.460000 3.245000 ;
        RECT 10.150000 2.100000 10.400000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.145000 0.350000  0.710000 0.790000 ;
      RECT 0.540000 0.790000  0.710000 2.180000 ;
      RECT 0.540000 2.180000  3.440000 2.350000 ;
      RECT 0.640000 2.350000  3.440000 2.380000 ;
      RECT 0.640000 2.380000  0.890000 2.980000 ;
      RECT 1.515000 1.820000  2.395000 2.010000 ;
      RECT 1.530000 0.395000  1.865000 0.810000 ;
      RECT 1.530000 0.810000  2.475000 1.010000 ;
      RECT 2.145000 1.010000  2.475000 1.220000 ;
      RECT 2.145000 1.220000  2.505000 1.575000 ;
      RECT 2.145000 1.575000  2.395000 1.820000 ;
      RECT 2.565000 1.745000  2.940000 2.010000 ;
      RECT 2.645000 0.255000  4.465000 0.465000 ;
      RECT 2.645000 0.465000  2.940000 1.090000 ;
      RECT 2.675000 1.090000  2.940000 1.745000 ;
      RECT 3.115000 0.635000  3.365000 1.840000 ;
      RECT 3.115000 1.840000  3.440000 2.180000 ;
      RECT 3.170000 2.380000  3.440000 2.705000 ;
      RECT 3.535000 0.465000  3.705000 1.670000 ;
      RECT 3.620000 2.275000  4.055000 2.705000 ;
      RECT 3.875000 0.635000  4.125000 1.075000 ;
      RECT 3.875000 1.075000  4.055000 2.020000 ;
      RECT 3.875000 2.020000  5.695000 2.190000 ;
      RECT 3.875000 2.190000  4.055000 2.275000 ;
      RECT 4.280000 1.470000  4.610000 1.800000 ;
      RECT 4.295000 0.465000  4.465000 0.790000 ;
      RECT 4.295000 0.790000  5.695000 0.960000 ;
      RECT 4.440000 1.130000  6.195000 1.300000 ;
      RECT 4.440000 1.300000  4.610000 1.470000 ;
      RECT 4.990000 2.190000  5.300000 2.705000 ;
      RECT 5.365000 1.470000  5.695000 2.020000 ;
      RECT 5.525000 0.255000  6.535000 0.425000 ;
      RECT 5.525000 0.425000  5.695000 0.790000 ;
      RECT 5.865000 0.595000  6.195000 1.130000 ;
      RECT 5.865000 1.300000  6.035000 1.970000 ;
      RECT 5.865000 1.970000  6.700000 2.140000 ;
      RECT 5.990000 2.140000  6.700000 2.980000 ;
      RECT 6.205000 1.470000  6.510000 1.630000 ;
      RECT 6.205000 1.630000  7.560000 1.800000 ;
      RECT 6.365000 0.425000  6.535000 1.125000 ;
      RECT 6.365000 1.125000  7.420000 1.295000 ;
      RECT 6.705000 0.625000  7.900000 0.955000 ;
      RECT 6.750000 1.295000  7.420000 1.455000 ;
      RECT 6.870000 2.535000  7.900000 2.705000 ;
      RECT 6.870000 2.705000  7.600000 2.865000 ;
      RECT 7.310000 1.800000  7.560000 2.365000 ;
      RECT 7.730000 0.955000  7.900000 1.125000 ;
      RECT 7.730000 1.125000  9.220000 1.295000 ;
      RECT 7.730000 1.295000  7.900000 2.535000 ;
      RECT 8.070000 1.965000  9.560000 2.135000 ;
      RECT 8.070000 2.135000  9.050000 2.335000 ;
      RECT 8.680000 2.335000  9.010000 2.980000 ;
      RECT 8.920000 1.295000  9.220000 1.795000 ;
      RECT 9.045000 0.575000  9.560000 0.955000 ;
      RECT 9.390000 0.955000  9.560000 1.965000 ;
      RECT 9.650000 2.305000  9.980000 2.980000 ;
      RECT 9.730000 0.530000  9.980000 1.320000 ;
      RECT 9.730000 1.320000 10.615000 1.650000 ;
      RECT 9.730000 1.650000  9.980000 2.305000 ;
  END
END sky130_fd_sc_ms__dfrtn_1

* File: sky130_fd_sc_ms__dlxtn_2.pxi.spice
* Created: Fri Aug 28 17:29:42 2020
* 
x_PM_SKY130_FD_SC_MS__DLXTN_2%D N_D_M1016_g N_D_M1001_g D N_D_c_135_n
+ N_D_c_136_n PM_SKY130_FD_SC_MS__DLXTN_2%D
x_PM_SKY130_FD_SC_MS__DLXTN_2%GATE_N N_GATE_N_M1004_g N_GATE_N_M1017_g GATE_N
+ N_GATE_N_c_164_n PM_SKY130_FD_SC_MS__DLXTN_2%GATE_N
x_PM_SKY130_FD_SC_MS__DLXTN_2%A_232_82# N_A_232_82#_M1004_d N_A_232_82#_M1017_d
+ N_A_232_82#_c_206_n N_A_232_82#_M1018_g N_A_232_82#_c_208_n
+ N_A_232_82#_M1008_g N_A_232_82#_c_209_n N_A_232_82#_M1002_g
+ N_A_232_82#_c_210_n N_A_232_82#_M1015_g N_A_232_82#_c_211_n
+ N_A_232_82#_c_212_n N_A_232_82#_c_213_n N_A_232_82#_c_214_n
+ N_A_232_82#_c_215_n N_A_232_82#_c_216_n N_A_232_82#_c_224_n
+ N_A_232_82#_c_254_p N_A_232_82#_c_225_n N_A_232_82#_c_226_n
+ N_A_232_82#_c_227_n N_A_232_82#_c_228_n N_A_232_82#_c_229_n
+ N_A_232_82#_c_217_n N_A_232_82#_c_218_n N_A_232_82#_c_219_n
+ N_A_232_82#_c_220_n N_A_232_82#_c_221_n PM_SKY130_FD_SC_MS__DLXTN_2%A_232_82#
x_PM_SKY130_FD_SC_MS__DLXTN_2%A_27_120# N_A_27_120#_M1016_s N_A_27_120#_M1001_s
+ N_A_27_120#_c_364_n N_A_27_120#_M1009_g N_A_27_120#_c_366_n
+ N_A_27_120#_c_367_n N_A_27_120#_M1003_g N_A_27_120#_c_375_n
+ N_A_27_120#_c_368_n N_A_27_120#_c_395_n N_A_27_120#_c_383_n
+ N_A_27_120#_c_369_n N_A_27_120#_c_370_n N_A_27_120#_c_371_n
+ N_A_27_120#_c_372_n N_A_27_120#_c_377_n N_A_27_120#_c_373_n
+ PM_SKY130_FD_SC_MS__DLXTN_2%A_27_120#
x_PM_SKY130_FD_SC_MS__DLXTN_2%A_369_392# N_A_369_392#_M1008_s
+ N_A_369_392#_M1018_s N_A_369_392#_M1012_g N_A_369_392#_M1013_g
+ N_A_369_392#_c_478_n N_A_369_392#_c_488_n N_A_369_392#_c_489_n
+ N_A_369_392#_c_479_n N_A_369_392#_c_480_n N_A_369_392#_c_481_n
+ N_A_369_392#_c_482_n N_A_369_392#_c_483_n N_A_369_392#_c_484_n
+ N_A_369_392#_c_485_n PM_SKY130_FD_SC_MS__DLXTN_2%A_369_392#
x_PM_SKY130_FD_SC_MS__DLXTN_2%A_842_405# N_A_842_405#_M1011_d
+ N_A_842_405#_M1014_d N_A_842_405#_M1007_g N_A_842_405#_M1006_g
+ N_A_842_405#_M1005_g N_A_842_405#_M1000_g N_A_842_405#_M1010_g
+ N_A_842_405#_M1019_g N_A_842_405#_c_588_n N_A_842_405#_c_589_n
+ N_A_842_405#_c_598_n N_A_842_405#_c_599_n N_A_842_405#_c_600_n
+ N_A_842_405#_c_590_n N_A_842_405#_c_591_n N_A_842_405#_c_601_n
+ N_A_842_405#_c_641_p N_A_842_405#_c_592_n N_A_842_405#_c_593_n
+ N_A_842_405#_c_602_n PM_SKY130_FD_SC_MS__DLXTN_2%A_842_405#
x_PM_SKY130_FD_SC_MS__DLXTN_2%A_672_392# N_A_672_392#_M1002_d
+ N_A_672_392#_M1012_d N_A_672_392#_M1014_g N_A_672_392#_M1011_g
+ N_A_672_392#_c_686_n N_A_672_392#_c_687_n N_A_672_392#_c_699_n
+ N_A_672_392#_c_688_n N_A_672_392#_c_689_n
+ PM_SKY130_FD_SC_MS__DLXTN_2%A_672_392#
x_PM_SKY130_FD_SC_MS__DLXTN_2%VPWR N_VPWR_M1001_d N_VPWR_M1018_d N_VPWR_M1007_d
+ N_VPWR_M1005_d N_VPWR_M1019_d N_VPWR_c_759_n N_VPWR_c_760_n N_VPWR_c_761_n
+ N_VPWR_c_762_n N_VPWR_c_763_n N_VPWR_c_764_n N_VPWR_c_765_n N_VPWR_c_766_n
+ N_VPWR_c_767_n VPWR N_VPWR_c_768_n N_VPWR_c_769_n N_VPWR_c_770_n
+ N_VPWR_c_771_n N_VPWR_c_772_n N_VPWR_c_758_n PM_SKY130_FD_SC_MS__DLXTN_2%VPWR
x_PM_SKY130_FD_SC_MS__DLXTN_2%Q N_Q_M1000_d N_Q_M1005_s N_Q_c_841_n N_Q_c_842_n
+ Q Q Q N_Q_c_843_n Q PM_SKY130_FD_SC_MS__DLXTN_2%Q
x_PM_SKY130_FD_SC_MS__DLXTN_2%VGND N_VGND_M1016_d N_VGND_M1008_d N_VGND_M1006_d
+ N_VGND_M1000_s N_VGND_M1010_s N_VGND_c_864_n N_VGND_c_865_n N_VGND_c_866_n
+ N_VGND_c_867_n N_VGND_c_868_n VGND N_VGND_c_869_n N_VGND_c_870_n
+ N_VGND_c_871_n N_VGND_c_872_n N_VGND_c_873_n N_VGND_c_874_n N_VGND_c_875_n
+ N_VGND_c_876_n N_VGND_c_877_n N_VGND_c_878_n PM_SKY130_FD_SC_MS__DLXTN_2%VGND
cc_1 VNB N_D_M1016_g 0.0283486f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.875
cc_2 VNB N_D_M1001_g 0.0015305f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.54
cc_3 VNB N_D_c_135_n 0.00404056f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_4 VNB N_D_c_136_n 0.0694963f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.465
cc_5 VNB N_GATE_N_M1004_g 0.0303764f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.875
cc_6 VNB GATE_N 0.00262174f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_GATE_N_c_164_n 0.0199144f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_8 VNB N_A_232_82#_c_206_n 0.011531f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.54
cc_9 VNB N_A_232_82#_M1018_g 0.0168108f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_10 VNB N_A_232_82#_c_208_n 0.0183869f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_11 VNB N_A_232_82#_c_209_n 0.0142471f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.465
cc_12 VNB N_A_232_82#_c_210_n 0.0167029f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.665
cc_13 VNB N_A_232_82#_c_211_n 0.00785913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_232_82#_c_212_n 0.0137619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_232_82#_c_213_n 0.0286494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_232_82#_c_214_n 0.00787851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_232_82#_c_215_n 0.00927555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_232_82#_c_216_n 0.00410622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_232_82#_c_217_n 0.039075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_232_82#_c_218_n 5.48748e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_232_82#_c_219_n 0.020808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_232_82#_c_220_n 0.00429395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_232_82#_c_221_n 0.0275096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_120#_c_364_n 0.0484273f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.54
cc_25 VNB N_A_27_120#_M1009_g 0.00179016f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_26 VNB N_A_27_120#_c_366_n 0.0194095f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_27 VNB N_A_27_120#_c_367_n 0.0158242f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_28 VNB N_A_27_120#_c_368_n 0.00560545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_120#_c_369_n 0.0218103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_120#_c_370_n 0.00147483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_120#_c_371_n 0.00304925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_120#_c_372_n 0.0278554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_120#_c_373_n 0.00714823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_369_392#_c_478_n 0.00241858f $X=-0.19 $Y=-0.245 $X2=0.655
+ $Y2=1.465
cc_35 VNB N_A_369_392#_c_479_n 0.00222566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_369_392#_c_480_n 0.00974233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_369_392#_c_481_n 0.0388791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_369_392#_c_482_n 0.00315129f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_369_392#_c_483_n 0.0205788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_369_392#_c_484_n 0.0080822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_369_392#_c_485_n 0.0145211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_842_405#_M1006_g 0.0414386f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_43 VNB N_A_842_405#_M1005_g 0.00221276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_842_405#_M1000_g 0.02472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_842_405#_M1010_g 0.0271225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_842_405#_M1019_g 0.00290854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_842_405#_c_588_n 0.0597619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_842_405#_c_589_n 0.0504497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_842_405#_c_590_n 0.00795778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_842_405#_c_591_n 0.0034055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_842_405#_c_592_n 0.0084286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_842_405#_c_593_n 0.00202256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_672_392#_M1014_g 5.7532e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_54 VNB N_A_672_392#_M1011_g 0.024451f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_55 VNB N_A_672_392#_c_686_n 0.0399447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_672_392#_c_687_n 0.00298842f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_57 VNB N_A_672_392#_c_688_n 0.00379072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_672_392#_c_689_n 0.0286454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VPWR_c_758_n 0.302998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_Q_c_841_n 0.00267235f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_61 VNB N_Q_c_842_n 0.00227864f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_62 VNB N_Q_c_843_n 0.00373325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_864_n 0.0103486f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_64 VNB N_VGND_c_865_n 0.0103936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_866_n 0.00786656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_867_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_868_n 0.0542709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_869_n 0.0195351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_870_n 0.0439744f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_871_n 0.0430783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_872_n 0.0200091f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_873_n 0.0172943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_874_n 0.0196327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_875_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_876_n 0.00619583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_877_n 0.0054847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_878_n 0.422042f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VPB N_D_M1001_g 0.0486432f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.54
cc_79 VPB N_D_c_135_n 0.0123656f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_80 VPB N_GATE_N_M1017_g 0.0390372f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=2.54
cc_81 VPB GATE_N 0.00260948f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_82 VPB N_GATE_N_c_164_n 0.0127652f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_83 VPB N_A_232_82#_M1018_g 0.0334551f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_84 VPB N_A_232_82#_M1015_g 0.0521586f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_232_82#_c_224_n 0.00641506f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_A_232_82#_c_225_n 0.00818583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_232_82#_c_226_n 7.63471e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_232_82#_c_227_n 0.0127742f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_232_82#_c_228_n 0.0232178f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_232_82#_c_229_n 0.00682609f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_232_82#_c_218_n 0.00380583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_232_82#_c_219_n 0.0162329f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_232_82#_c_220_n 0.00223583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_232_82#_c_221_n 0.0252921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_A_27_120#_M1009_g 0.0295937f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_96 VPB N_A_27_120#_c_375_n 0.0358457f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_97 VPB N_A_27_120#_c_368_n 0.00273869f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_27_120#_c_377_n 0.0136666f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_369_392#_M1012_g 0.0207809f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_100 VPB N_A_369_392#_c_478_n 0.00104552f $X=-0.19 $Y=1.66 $X2=0.655 $Y2=1.465
cc_101 VPB N_A_369_392#_c_488_n 0.00879291f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_102 VPB N_A_369_392#_c_489_n 0.0101735f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_369_392#_c_482_n 0.00102696f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_369_392#_c_483_n 0.0141739f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_842_405#_M1007_g 0.0235219f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_106 VPB N_A_842_405#_M1006_g 0.0233314f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_107 VPB N_A_842_405#_M1005_g 0.0255102f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_842_405#_M1019_g 0.0287837f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_842_405#_c_598_n 0.00410771f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_842_405#_c_599_n 0.0124508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_842_405#_c_600_n 0.00829389f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_842_405#_c_601_n 0.00351153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_842_405#_c_602_n 0.0564811f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_672_392#_M1014_g 0.0264986f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_115 VPB N_A_672_392#_c_688_n 0.00187511f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_759_n 0.00969617f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_117 VPB N_VPWR_c_760_n 0.0140952f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_761_n 0.011478f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_762_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_763_n 0.0646317f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_764_n 0.0239248f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_765_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_766_n 0.0218405f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_767_n 0.00410958f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_768_n 0.0345071f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_769_n 0.0221566f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_770_n 0.00660399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_771_n 0.0393527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_772_n 0.0263687f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_758_n 0.104095f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_Q_c_843_n 0.00321419f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 N_D_M1016_g N_GATE_N_M1004_g 0.0184595f $X=0.495 $Y=0.875 $X2=0 $Y2=0
cc_133 N_D_c_136_n N_GATE_N_M1004_g 0.00663446f $X=0.655 $Y=1.465 $X2=0 $Y2=0
cc_134 N_D_M1001_g N_GATE_N_M1017_g 0.0161448f $X=0.655 $Y=2.54 $X2=0 $Y2=0
cc_135 N_D_c_136_n GATE_N 3.81053e-19 $X=0.655 $Y=1.465 $X2=0 $Y2=0
cc_136 N_D_c_136_n N_GATE_N_c_164_n 0.0174277f $X=0.655 $Y=1.465 $X2=0 $Y2=0
cc_137 N_D_M1001_g N_A_232_82#_c_228_n 4.79724e-19 $X=0.655 $Y=2.54 $X2=0 $Y2=0
cc_138 N_D_M1001_g N_A_27_120#_c_375_n 0.0154244f $X=0.655 $Y=2.54 $X2=0 $Y2=0
cc_139 N_D_M1016_g N_A_27_120#_c_368_n 0.00397398f $X=0.495 $Y=0.875 $X2=0 $Y2=0
cc_140 N_D_M1001_g N_A_27_120#_c_368_n 0.0129118f $X=0.655 $Y=2.54 $X2=0 $Y2=0
cc_141 N_D_c_135_n N_A_27_120#_c_368_n 0.0348574f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_142 N_D_c_136_n N_A_27_120#_c_368_n 0.0116014f $X=0.655 $Y=1.465 $X2=0 $Y2=0
cc_143 N_D_M1016_g N_A_27_120#_c_383_n 4.90322e-19 $X=0.495 $Y=0.875 $X2=0 $Y2=0
cc_144 N_D_M1016_g N_A_27_120#_c_372_n 0.0266287f $X=0.495 $Y=0.875 $X2=0 $Y2=0
cc_145 N_D_c_135_n N_A_27_120#_c_372_n 0.024806f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_146 N_D_c_136_n N_A_27_120#_c_372_n 0.0026784f $X=0.655 $Y=1.465 $X2=0 $Y2=0
cc_147 N_D_M1001_g N_A_27_120#_c_377_n 0.0170813f $X=0.655 $Y=2.54 $X2=0 $Y2=0
cc_148 N_D_c_135_n N_A_27_120#_c_377_n 0.0155123f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_149 N_D_c_136_n N_A_27_120#_c_377_n 0.00484569f $X=0.655 $Y=1.465 $X2=0 $Y2=0
cc_150 N_D_M1001_g N_VPWR_c_759_n 0.00361707f $X=0.655 $Y=2.54 $X2=0 $Y2=0
cc_151 N_D_M1001_g N_VPWR_c_764_n 0.005209f $X=0.655 $Y=2.54 $X2=0 $Y2=0
cc_152 N_D_M1001_g N_VPWR_c_758_n 0.00986738f $X=0.655 $Y=2.54 $X2=0 $Y2=0
cc_153 N_D_M1016_g N_VGND_c_869_n 0.00327294f $X=0.495 $Y=0.875 $X2=0 $Y2=0
cc_154 N_D_M1016_g N_VGND_c_878_n 0.00476395f $X=0.495 $Y=0.875 $X2=0 $Y2=0
cc_155 N_GATE_N_M1004_g N_A_232_82#_c_214_n 0.00461345f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_156 GATE_N N_A_232_82#_c_214_n 0.00948482f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_157 N_GATE_N_c_164_n N_A_232_82#_c_214_n 0.00100798f $X=1.15 $Y=1.615 $X2=0
+ $Y2=0
cc_158 N_GATE_N_M1004_g N_A_232_82#_c_215_n 0.00303911f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_159 N_GATE_N_M1004_g N_A_232_82#_c_216_n 0.00593761f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_160 GATE_N N_A_232_82#_c_216_n 0.0263887f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_161 N_GATE_N_c_164_n N_A_232_82#_c_216_n 0.00218737f $X=1.15 $Y=1.615 $X2=0
+ $Y2=0
cc_162 N_GATE_N_M1017_g N_A_232_82#_c_224_n 4.52945e-19 $X=1.205 $Y=2.54 $X2=0
+ $Y2=0
cc_163 N_GATE_N_M1017_g N_A_232_82#_c_228_n 0.0168272f $X=1.205 $Y=2.54 $X2=0
+ $Y2=0
cc_164 GATE_N N_A_232_82#_c_228_n 0.00240021f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_165 N_GATE_N_M1017_g N_A_232_82#_c_229_n 0.0109124f $X=1.205 $Y=2.54 $X2=0
+ $Y2=0
cc_166 N_GATE_N_M1004_g N_A_232_82#_c_217_n 0.014014f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_167 GATE_N N_A_232_82#_c_219_n 3.56619e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_168 N_GATE_N_c_164_n N_A_232_82#_c_219_n 0.0168587f $X=1.15 $Y=1.615 $X2=0
+ $Y2=0
cc_169 N_GATE_N_M1017_g N_A_27_120#_c_375_n 4.57948e-19 $X=1.205 $Y=2.54 $X2=0
+ $Y2=0
cc_170 N_GATE_N_M1004_g N_A_27_120#_c_368_n 0.0059942f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_171 N_GATE_N_M1017_g N_A_27_120#_c_368_n 0.00308057f $X=1.205 $Y=2.54 $X2=0
+ $Y2=0
cc_172 GATE_N N_A_27_120#_c_368_n 0.0228108f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_173 N_GATE_N_c_164_n N_A_27_120#_c_368_n 0.00187493f $X=1.15 $Y=1.615 $X2=0
+ $Y2=0
cc_174 N_GATE_N_M1004_g N_A_27_120#_c_395_n 0.0164833f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_175 N_GATE_N_M1004_g N_A_27_120#_c_383_n 0.00644004f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_176 N_GATE_N_M1004_g N_A_27_120#_c_370_n 0.00578481f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_177 N_GATE_N_M1004_g N_A_27_120#_c_372_n 0.00668497f $X=1.085 $Y=0.78 $X2=0
+ $Y2=0
cc_178 N_GATE_N_M1017_g N_A_27_120#_c_377_n 0.00353156f $X=1.205 $Y=2.54 $X2=0
+ $Y2=0
cc_179 N_GATE_N_M1017_g N_A_369_392#_c_489_n 2.77935e-19 $X=1.205 $Y=2.54 $X2=0
+ $Y2=0
cc_180 N_GATE_N_M1017_g N_VPWR_c_759_n 0.00361707f $X=1.205 $Y=2.54 $X2=0 $Y2=0
cc_181 GATE_N N_VPWR_c_759_n 0.00308887f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_182 N_GATE_N_c_164_n N_VPWR_c_759_n 5.55981e-19 $X=1.15 $Y=1.615 $X2=0 $Y2=0
cc_183 N_GATE_N_M1017_g N_VPWR_c_768_n 0.005209f $X=1.205 $Y=2.54 $X2=0 $Y2=0
cc_184 N_GATE_N_M1017_g N_VPWR_c_758_n 0.00987709f $X=1.205 $Y=2.54 $X2=0 $Y2=0
cc_185 N_GATE_N_M1004_g N_VGND_c_870_n 0.00382493f $X=1.085 $Y=0.78 $X2=0 $Y2=0
cc_186 N_GATE_N_M1004_g N_VGND_c_874_n 0.0029536f $X=1.085 $Y=0.78 $X2=0 $Y2=0
cc_187 N_GATE_N_M1004_g N_VGND_c_878_n 0.00479772f $X=1.085 $Y=0.78 $X2=0 $Y2=0
cc_188 N_A_232_82#_M1018_g N_A_27_120#_c_364_n 0.00952668f $X=2.215 $Y=2.38
+ $X2=0 $Y2=0
cc_189 N_A_232_82#_c_208_n N_A_27_120#_c_364_n 0.00378548f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_190 N_A_232_82#_c_212_n N_A_27_120#_c_364_n 0.00491582f $X=2.355 $Y=1.26
+ $X2=0 $Y2=0
cc_191 N_A_232_82#_M1018_g N_A_27_120#_M1009_g 0.0339985f $X=2.215 $Y=2.38 $X2=0
+ $Y2=0
cc_192 N_A_232_82#_c_224_n N_A_27_120#_M1009_g 0.013675f $X=2.875 $Y=2.525 $X2=0
+ $Y2=0
cc_193 N_A_232_82#_c_254_p N_A_27_120#_M1009_g 0.00717936f $X=2.96 $Y=2.905
+ $X2=0 $Y2=0
cc_194 N_A_232_82#_c_226_n N_A_27_120#_M1009_g 0.00447908f $X=3.045 $Y=2.99
+ $X2=0 $Y2=0
cc_195 N_A_232_82#_c_213_n N_A_27_120#_c_366_n 0.0229627f $X=3.825 $Y=1.185
+ $X2=0 $Y2=0
cc_196 N_A_232_82#_c_208_n N_A_27_120#_c_367_n 0.00442582f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_197 N_A_232_82#_c_209_n N_A_27_120#_c_367_n 0.0229627f $X=3.605 $Y=1.11 $X2=0
+ $Y2=0
cc_198 N_A_232_82#_c_228_n N_A_27_120#_c_375_n 0.00410401f $X=1.43 $Y=2.265
+ $X2=0 $Y2=0
cc_199 N_A_232_82#_c_214_n N_A_27_120#_c_368_n 0.00182037f $X=1.485 $Y=1.045
+ $X2=0 $Y2=0
cc_200 N_A_232_82#_M1004_d N_A_27_120#_c_395_n 0.00866525f $X=1.16 $Y=0.41 $X2=0
+ $Y2=0
cc_201 N_A_232_82#_c_214_n N_A_27_120#_c_395_n 0.00975585f $X=1.485 $Y=1.045
+ $X2=0 $Y2=0
cc_202 N_A_232_82#_M1004_d N_A_27_120#_c_383_n 0.0058378f $X=1.16 $Y=0.41 $X2=0
+ $Y2=0
cc_203 N_A_232_82#_M1004_d N_A_27_120#_c_369_n 0.00239893f $X=1.16 $Y=0.41 $X2=0
+ $Y2=0
cc_204 N_A_232_82#_c_208_n N_A_27_120#_c_369_n 0.0157054f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_205 N_A_232_82#_c_214_n N_A_27_120#_c_369_n 0.00585336f $X=1.485 $Y=1.045
+ $X2=0 $Y2=0
cc_206 N_A_232_82#_c_215_n N_A_27_120#_c_369_n 0.0169889f $X=1.685 $Y=1.17 $X2=0
+ $Y2=0
cc_207 N_A_232_82#_c_217_n N_A_27_120#_c_369_n 0.00199179f $X=1.72 $Y=0.925
+ $X2=0 $Y2=0
cc_208 N_A_232_82#_c_208_n N_A_27_120#_c_371_n 0.00800558f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_209 N_A_232_82#_c_214_n N_A_27_120#_c_372_n 0.0106332f $X=1.485 $Y=1.045
+ $X2=0 $Y2=0
cc_210 N_A_232_82#_c_228_n N_A_27_120#_c_377_n 7.41183e-19 $X=1.43 $Y=2.265
+ $X2=0 $Y2=0
cc_211 N_A_232_82#_M1018_g N_A_27_120#_c_373_n 0.00202018f $X=2.215 $Y=2.38
+ $X2=0 $Y2=0
cc_212 N_A_232_82#_c_212_n N_A_27_120#_c_373_n 2.84937e-19 $X=2.355 $Y=1.26
+ $X2=0 $Y2=0
cc_213 N_A_232_82#_c_224_n N_A_369_392#_M1018_s 0.00752555f $X=2.875 $Y=2.525
+ $X2=0 $Y2=0
cc_214 N_A_232_82#_M1015_g N_A_369_392#_M1012_g 0.0221739f $X=3.88 $Y=2.725
+ $X2=0 $Y2=0
cc_215 N_A_232_82#_c_224_n N_A_369_392#_M1012_g 0.00144159f $X=2.875 $Y=2.525
+ $X2=0 $Y2=0
cc_216 N_A_232_82#_c_254_p N_A_369_392#_M1012_g 0.00446725f $X=2.96 $Y=2.905
+ $X2=0 $Y2=0
cc_217 N_A_232_82#_c_225_n N_A_369_392#_M1012_g 0.0152619f $X=4.02 $Y=2.99 $X2=0
+ $Y2=0
cc_218 N_A_232_82#_c_221_n N_A_369_392#_M1012_g 4.19954e-19 $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_219 N_A_232_82#_c_206_n N_A_369_392#_c_478_n 0.00462651f $X=2.125 $Y=1.26
+ $X2=0 $Y2=0
cc_220 N_A_232_82#_M1018_g N_A_369_392#_c_478_n 0.0139947f $X=2.215 $Y=2.38
+ $X2=0 $Y2=0
cc_221 N_A_232_82#_c_208_n N_A_369_392#_c_478_n 0.0094035f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_222 N_A_232_82#_c_212_n N_A_369_392#_c_478_n 0.00522206f $X=2.355 $Y=1.26
+ $X2=0 $Y2=0
cc_223 N_A_232_82#_c_215_n N_A_369_392#_c_478_n 0.0326777f $X=1.685 $Y=1.17
+ $X2=0 $Y2=0
cc_224 N_A_232_82#_c_216_n N_A_369_392#_c_478_n 0.046382f $X=1.685 $Y=1.57 $X2=0
+ $Y2=0
cc_225 N_A_232_82#_c_229_n N_A_369_392#_c_478_n 0.00124535f $X=1.46 $Y=2.1 $X2=0
+ $Y2=0
cc_226 N_A_232_82#_c_217_n N_A_369_392#_c_478_n 0.00162222f $X=1.72 $Y=0.925
+ $X2=0 $Y2=0
cc_227 N_A_232_82#_c_219_n N_A_369_392#_c_478_n 0.00255297f $X=1.72 $Y=1.605
+ $X2=0 $Y2=0
cc_228 N_A_232_82#_c_212_n N_A_369_392#_c_488_n 0.00379117f $X=2.355 $Y=1.26
+ $X2=0 $Y2=0
cc_229 N_A_232_82#_c_224_n N_A_369_392#_c_488_n 0.0190563f $X=2.875 $Y=2.525
+ $X2=0 $Y2=0
cc_230 N_A_232_82#_c_206_n N_A_369_392#_c_489_n 0.00141981f $X=2.125 $Y=1.26
+ $X2=0 $Y2=0
cc_231 N_A_232_82#_M1018_g N_A_369_392#_c_489_n 0.0199656f $X=2.215 $Y=2.38
+ $X2=0 $Y2=0
cc_232 N_A_232_82#_c_224_n N_A_369_392#_c_489_n 0.0289802f $X=2.875 $Y=2.525
+ $X2=0 $Y2=0
cc_233 N_A_232_82#_c_229_n N_A_369_392#_c_489_n 0.0341526f $X=1.46 $Y=2.1 $X2=0
+ $Y2=0
cc_234 N_A_232_82#_c_218_n N_A_369_392#_c_489_n 0.00497552f $X=1.72 $Y=1.605
+ $X2=0 $Y2=0
cc_235 N_A_232_82#_c_219_n N_A_369_392#_c_489_n 4.32246e-19 $X=1.72 $Y=1.605
+ $X2=0 $Y2=0
cc_236 N_A_232_82#_c_209_n N_A_369_392#_c_480_n 0.0198684f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_237 N_A_232_82#_c_213_n N_A_369_392#_c_480_n 0.0014907f $X=3.825 $Y=1.185
+ $X2=0 $Y2=0
cc_238 N_A_232_82#_c_209_n N_A_369_392#_c_481_n 0.0101699f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_239 N_A_232_82#_c_210_n N_A_369_392#_c_482_n 3.61841e-19 $X=3.825 $Y=1.485
+ $X2=0 $Y2=0
cc_240 N_A_232_82#_M1015_g N_A_369_392#_c_482_n 4.66392e-19 $X=3.88 $Y=2.725
+ $X2=0 $Y2=0
cc_241 N_A_232_82#_c_210_n N_A_369_392#_c_483_n 0.0174101f $X=3.825 $Y=1.485
+ $X2=0 $Y2=0
cc_242 N_A_232_82#_c_209_n N_A_369_392#_c_484_n 0.00336691f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_243 N_A_232_82#_c_210_n N_A_369_392#_c_484_n 0.00121983f $X=3.825 $Y=1.485
+ $X2=0 $Y2=0
cc_244 N_A_232_82#_c_209_n N_A_369_392#_c_485_n 0.0109494f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_245 N_A_232_82#_c_213_n N_A_369_392#_c_485_n 0.00477162f $X=3.825 $Y=1.185
+ $X2=0 $Y2=0
cc_246 N_A_232_82#_c_221_n N_A_369_392#_c_485_n 0.00690996f $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_247 N_A_232_82#_c_225_n N_A_842_405#_M1007_g 0.00119414f $X=4.02 $Y=2.99
+ $X2=0 $Y2=0
cc_248 N_A_232_82#_M1015_g N_A_842_405#_M1006_g 0.00224512f $X=3.88 $Y=2.725
+ $X2=0 $Y2=0
cc_249 N_A_232_82#_c_213_n N_A_842_405#_M1006_g 0.00421996f $X=3.825 $Y=1.185
+ $X2=0 $Y2=0
cc_250 N_A_232_82#_c_227_n N_A_842_405#_M1006_g 0.00366868f $X=4.105 $Y=2.905
+ $X2=0 $Y2=0
cc_251 N_A_232_82#_c_220_n N_A_842_405#_M1006_g 0.00176725f $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_252 N_A_232_82#_c_221_n N_A_842_405#_M1006_g 0.0170611f $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_253 N_A_232_82#_c_227_n N_A_842_405#_c_598_n 0.0262086f $X=4.105 $Y=2.905
+ $X2=0 $Y2=0
cc_254 N_A_232_82#_M1015_g N_A_842_405#_c_602_n 0.0484491f $X=3.88 $Y=2.725
+ $X2=0 $Y2=0
cc_255 N_A_232_82#_c_227_n N_A_842_405#_c_602_n 0.00828434f $X=4.105 $Y=2.905
+ $X2=0 $Y2=0
cc_256 N_A_232_82#_c_220_n N_A_842_405#_c_602_n 0.00107151f $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_257 N_A_232_82#_c_221_n N_A_842_405#_c_602_n 0.00935259f $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_258 N_A_232_82#_c_225_n N_A_672_392#_M1012_d 0.00356836f $X=4.02 $Y=2.99
+ $X2=0 $Y2=0
cc_259 N_A_232_82#_c_220_n N_A_672_392#_c_686_n 0.0114859f $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_260 N_A_232_82#_c_221_n N_A_672_392#_c_686_n 2.9672e-19 $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_261 N_A_232_82#_c_209_n N_A_672_392#_c_687_n 0.00856348f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_262 N_A_232_82#_c_213_n N_A_672_392#_c_687_n 0.00190905f $X=3.825 $Y=1.185
+ $X2=0 $Y2=0
cc_263 N_A_232_82#_c_220_n N_A_672_392#_c_687_n 0.0149091f $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_264 N_A_232_82#_c_221_n N_A_672_392#_c_687_n 0.00507885f $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_265 N_A_232_82#_M1015_g N_A_672_392#_c_699_n 0.0183269f $X=3.88 $Y=2.725
+ $X2=0 $Y2=0
cc_266 N_A_232_82#_c_224_n N_A_672_392#_c_699_n 0.00974321f $X=2.875 $Y=2.525
+ $X2=0 $Y2=0
cc_267 N_A_232_82#_c_254_p N_A_672_392#_c_699_n 0.00640505f $X=2.96 $Y=2.905
+ $X2=0 $Y2=0
cc_268 N_A_232_82#_c_225_n N_A_672_392#_c_699_n 0.0300593f $X=4.02 $Y=2.99 $X2=0
+ $Y2=0
cc_269 N_A_232_82#_c_227_n N_A_672_392#_c_699_n 0.0423538f $X=4.105 $Y=2.905
+ $X2=0 $Y2=0
cc_270 N_A_232_82#_c_209_n N_A_672_392#_c_688_n 6.33047e-19 $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_271 N_A_232_82#_c_210_n N_A_672_392#_c_688_n 0.0120805f $X=3.825 $Y=1.485
+ $X2=0 $Y2=0
cc_272 N_A_232_82#_M1015_g N_A_672_392#_c_688_n 0.0074333f $X=3.88 $Y=2.725
+ $X2=0 $Y2=0
cc_273 N_A_232_82#_c_213_n N_A_672_392#_c_688_n 0.00989251f $X=3.825 $Y=1.185
+ $X2=0 $Y2=0
cc_274 N_A_232_82#_c_220_n N_A_672_392#_c_688_n 0.0423538f $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_275 N_A_232_82#_c_221_n N_A_672_392#_c_688_n 0.0100291f $X=4.185 $Y=1.65
+ $X2=0 $Y2=0
cc_276 N_A_232_82#_c_224_n N_VPWR_M1018_d 0.0103748f $X=2.875 $Y=2.525 $X2=0
+ $Y2=0
cc_277 N_A_232_82#_c_228_n N_VPWR_c_759_n 0.0273513f $X=1.43 $Y=2.265 $X2=0
+ $Y2=0
cc_278 N_A_232_82#_M1018_g N_VPWR_c_760_n 0.00397791f $X=2.215 $Y=2.38 $X2=0
+ $Y2=0
cc_279 N_A_232_82#_c_224_n N_VPWR_c_760_n 0.0266399f $X=2.875 $Y=2.525 $X2=0
+ $Y2=0
cc_280 N_A_232_82#_c_226_n N_VPWR_c_760_n 0.0119562f $X=3.045 $Y=2.99 $X2=0
+ $Y2=0
cc_281 N_A_232_82#_M1018_g N_VPWR_c_768_n 0.00440215f $X=2.215 $Y=2.38 $X2=0
+ $Y2=0
cc_282 N_A_232_82#_c_224_n N_VPWR_c_768_n 0.00946875f $X=2.875 $Y=2.525 $X2=0
+ $Y2=0
cc_283 N_A_232_82#_c_228_n N_VPWR_c_768_n 0.0172262f $X=1.43 $Y=2.265 $X2=0
+ $Y2=0
cc_284 N_A_232_82#_M1015_g N_VPWR_c_771_n 0.00113339f $X=3.88 $Y=2.725 $X2=0
+ $Y2=0
cc_285 N_A_232_82#_c_224_n N_VPWR_c_771_n 0.00197169f $X=2.875 $Y=2.525 $X2=0
+ $Y2=0
cc_286 N_A_232_82#_c_225_n N_VPWR_c_771_n 0.0743861f $X=4.02 $Y=2.99 $X2=0 $Y2=0
cc_287 N_A_232_82#_c_226_n N_VPWR_c_771_n 0.0118974f $X=3.045 $Y=2.99 $X2=0
+ $Y2=0
cc_288 N_A_232_82#_c_225_n N_VPWR_c_772_n 0.0138114f $X=4.02 $Y=2.99 $X2=0 $Y2=0
cc_289 N_A_232_82#_M1018_g N_VPWR_c_758_n 0.00595788f $X=2.215 $Y=2.38 $X2=0
+ $Y2=0
cc_290 N_A_232_82#_c_224_n N_VPWR_c_758_n 0.0240232f $X=2.875 $Y=2.525 $X2=0
+ $Y2=0
cc_291 N_A_232_82#_c_225_n N_VPWR_c_758_n 0.0424364f $X=4.02 $Y=2.99 $X2=0 $Y2=0
cc_292 N_A_232_82#_c_226_n N_VPWR_c_758_n 0.00629995f $X=3.045 $Y=2.99 $X2=0
+ $Y2=0
cc_293 N_A_232_82#_c_228_n N_VPWR_c_758_n 0.0141903f $X=1.43 $Y=2.265 $X2=0
+ $Y2=0
cc_294 N_A_232_82#_c_224_n A_588_392# 0.00268432f $X=2.875 $Y=2.525 $X2=-0.19
+ $Y2=-0.245
cc_295 N_A_232_82#_c_254_p A_588_392# 0.00318252f $X=2.96 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_296 N_A_232_82#_c_225_n A_588_392# 0.00293798f $X=4.02 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_297 N_A_232_82#_c_227_n A_794_503# 0.00147774f $X=4.105 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_298 N_A_232_82#_c_208_n N_VGND_c_864_n 0.00196494f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_299 N_A_232_82#_c_209_n N_VGND_c_864_n 3.70241e-19 $X=3.605 $Y=1.11 $X2=0
+ $Y2=0
cc_300 N_A_232_82#_c_208_n N_VGND_c_870_n 0.00278271f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_301 N_A_232_82#_c_209_n N_VGND_c_871_n 9.44495e-19 $X=3.605 $Y=1.11 $X2=0
+ $Y2=0
cc_302 N_A_232_82#_c_208_n N_VGND_c_878_n 0.00363426f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_303 N_A_27_120#_c_369_n N_A_369_392#_M1008_s 0.00441657f $X=2.475 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_304 N_A_27_120#_c_364_n N_A_369_392#_c_478_n 3.44763e-19 $X=2.85 $Y=1.63
+ $X2=0 $Y2=0
cc_305 N_A_27_120#_M1009_g N_A_369_392#_c_478_n 9.58777e-19 $X=2.85 $Y=2.46
+ $X2=0 $Y2=0
cc_306 N_A_27_120#_c_369_n N_A_369_392#_c_478_n 0.0144209f $X=2.475 $Y=0.34
+ $X2=0 $Y2=0
cc_307 N_A_27_120#_c_371_n N_A_369_392#_c_478_n 0.0324263f $X=2.56 $Y=1.3 $X2=0
+ $Y2=0
cc_308 N_A_27_120#_c_373_n N_A_369_392#_c_478_n 0.0263966f $X=2.805 $Y=1.465
+ $X2=0 $Y2=0
cc_309 N_A_27_120#_c_364_n N_A_369_392#_c_488_n 0.00349359f $X=2.85 $Y=1.63
+ $X2=0 $Y2=0
cc_310 N_A_27_120#_M1009_g N_A_369_392#_c_488_n 0.0141343f $X=2.85 $Y=2.46 $X2=0
+ $Y2=0
cc_311 N_A_27_120#_c_366_n N_A_369_392#_c_488_n 0.0050599f $X=3.14 $Y=1.185
+ $X2=0 $Y2=0
cc_312 N_A_27_120#_c_373_n N_A_369_392#_c_488_n 0.0372099f $X=2.805 $Y=1.465
+ $X2=0 $Y2=0
cc_313 N_A_27_120#_M1009_g N_A_369_392#_c_489_n 0.00147976f $X=2.85 $Y=2.46
+ $X2=0 $Y2=0
cc_314 N_A_27_120#_c_367_n N_A_369_392#_c_479_n 0.00178439f $X=3.215 $Y=1.11
+ $X2=0 $Y2=0
cc_315 N_A_27_120#_c_364_n N_A_369_392#_c_482_n 2.00831e-19 $X=2.85 $Y=1.63
+ $X2=0 $Y2=0
cc_316 N_A_27_120#_M1009_g N_A_369_392#_c_482_n 0.0012292f $X=2.85 $Y=2.46 $X2=0
+ $Y2=0
cc_317 N_A_27_120#_c_366_n N_A_369_392#_c_482_n 8.35401e-19 $X=3.14 $Y=1.185
+ $X2=0 $Y2=0
cc_318 N_A_27_120#_c_373_n N_A_369_392#_c_482_n 0.0104417f $X=2.805 $Y=1.465
+ $X2=0 $Y2=0
cc_319 N_A_27_120#_c_364_n N_A_369_392#_c_483_n 0.0100759f $X=2.85 $Y=1.63 $X2=0
+ $Y2=0
cc_320 N_A_27_120#_M1009_g N_A_369_392#_c_483_n 0.0790361f $X=2.85 $Y=2.46 $X2=0
+ $Y2=0
cc_321 N_A_27_120#_c_366_n N_A_369_392#_c_483_n 0.00738423f $X=3.14 $Y=1.185
+ $X2=0 $Y2=0
cc_322 N_A_27_120#_c_373_n N_A_369_392#_c_483_n 5.53572e-19 $X=2.805 $Y=1.465
+ $X2=0 $Y2=0
cc_323 N_A_27_120#_c_364_n N_A_369_392#_c_484_n 0.00193199f $X=2.85 $Y=1.63
+ $X2=0 $Y2=0
cc_324 N_A_27_120#_c_367_n N_A_369_392#_c_484_n 0.0047803f $X=3.215 $Y=1.11
+ $X2=0 $Y2=0
cc_325 N_A_27_120#_c_371_n N_A_369_392#_c_484_n 0.00674121f $X=2.56 $Y=1.3 $X2=0
+ $Y2=0
cc_326 N_A_27_120#_c_373_n N_A_369_392#_c_484_n 0.00771809f $X=2.805 $Y=1.465
+ $X2=0 $Y2=0
cc_327 N_A_27_120#_M1009_g N_A_672_392#_c_699_n 0.00169208f $X=2.85 $Y=2.46
+ $X2=0 $Y2=0
cc_328 N_A_27_120#_c_375_n N_VPWR_c_759_n 0.0266809f $X=0.43 $Y=2.265 $X2=0
+ $Y2=0
cc_329 N_A_27_120#_M1009_g N_VPWR_c_760_n 0.00486648f $X=2.85 $Y=2.46 $X2=0
+ $Y2=0
cc_330 N_A_27_120#_c_375_n N_VPWR_c_764_n 0.014549f $X=0.43 $Y=2.265 $X2=0 $Y2=0
cc_331 N_A_27_120#_M1009_g N_VPWR_c_771_n 0.0037741f $X=2.85 $Y=2.46 $X2=0 $Y2=0
cc_332 N_A_27_120#_M1009_g N_VPWR_c_758_n 0.00488877f $X=2.85 $Y=2.46 $X2=0
+ $Y2=0
cc_333 N_A_27_120#_c_375_n N_VPWR_c_758_n 0.0119743f $X=0.43 $Y=2.265 $X2=0
+ $Y2=0
cc_334 N_A_27_120#_c_368_n N_VGND_M1016_d 7.20017e-19 $X=0.71 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_335 N_A_27_120#_c_395_n N_VGND_M1016_d 0.00789213f $X=1.145 $Y=0.665
+ $X2=-0.19 $Y2=-0.245
cc_336 N_A_27_120#_c_372_n N_VGND_M1016_d 0.00822019f $X=0.795 $Y=0.855
+ $X2=-0.19 $Y2=-0.245
cc_337 N_A_27_120#_c_369_n N_VGND_M1008_d 6.47853e-19 $X=2.475 $Y=0.34 $X2=0
+ $Y2=0
cc_338 N_A_27_120#_c_371_n N_VGND_M1008_d 0.0113692f $X=2.56 $Y=1.3 $X2=0 $Y2=0
cc_339 N_A_27_120#_c_364_n N_VGND_c_864_n 0.0127456f $X=2.85 $Y=1.63 $X2=0 $Y2=0
cc_340 N_A_27_120#_c_367_n N_VGND_c_864_n 0.00940057f $X=3.215 $Y=1.11 $X2=0
+ $Y2=0
cc_341 N_A_27_120#_c_369_n N_VGND_c_864_n 0.0148948f $X=2.475 $Y=0.34 $X2=0
+ $Y2=0
cc_342 N_A_27_120#_c_371_n N_VGND_c_864_n 0.0481399f $X=2.56 $Y=1.3 $X2=0 $Y2=0
cc_343 N_A_27_120#_c_373_n N_VGND_c_864_n 0.00988174f $X=2.805 $Y=1.465 $X2=0
+ $Y2=0
cc_344 N_A_27_120#_c_372_n N_VGND_c_869_n 0.0110697f $X=0.795 $Y=0.855 $X2=0
+ $Y2=0
cc_345 N_A_27_120#_c_395_n N_VGND_c_870_n 0.00313112f $X=1.145 $Y=0.665 $X2=0
+ $Y2=0
cc_346 N_A_27_120#_c_369_n N_VGND_c_870_n 0.086417f $X=2.475 $Y=0.34 $X2=0 $Y2=0
cc_347 N_A_27_120#_c_370_n N_VGND_c_870_n 0.0118998f $X=1.315 $Y=0.34 $X2=0
+ $Y2=0
cc_348 N_A_27_120#_c_367_n N_VGND_c_871_n 0.00539704f $X=3.215 $Y=1.11 $X2=0
+ $Y2=0
cc_349 N_A_27_120#_c_370_n N_VGND_c_874_n 0.0120702f $X=1.315 $Y=0.34 $X2=0
+ $Y2=0
cc_350 N_A_27_120#_c_372_n N_VGND_c_874_n 0.0255806f $X=0.795 $Y=0.855 $X2=0
+ $Y2=0
cc_351 N_A_27_120#_c_367_n N_VGND_c_878_n 0.0052351f $X=3.215 $Y=1.11 $X2=0
+ $Y2=0
cc_352 N_A_27_120#_c_395_n N_VGND_c_878_n 0.00556468f $X=1.145 $Y=0.665 $X2=0
+ $Y2=0
cc_353 N_A_27_120#_c_369_n N_VGND_c_878_n 0.049532f $X=2.475 $Y=0.34 $X2=0 $Y2=0
cc_354 N_A_27_120#_c_370_n N_VGND_c_878_n 0.00655543f $X=1.315 $Y=0.34 $X2=0
+ $Y2=0
cc_355 N_A_27_120#_c_372_n N_VGND_c_878_n 0.0175471f $X=0.795 $Y=0.855 $X2=0
+ $Y2=0
cc_356 N_A_369_392#_c_481_n N_A_842_405#_M1006_g 0.0358316f $X=4.21 $Y=0.42
+ $X2=0 $Y2=0
cc_357 N_A_369_392#_c_480_n N_A_672_392#_M1002_d 0.00217732f $X=4.21 $Y=0.42
+ $X2=-0.19 $Y2=-0.245
cc_358 N_A_369_392#_c_482_n N_A_672_392#_M1012_d 0.00110467f $X=3.345 $Y=1.635
+ $X2=0 $Y2=0
cc_359 N_A_369_392#_c_480_n N_A_672_392#_c_686_n 0.00333692f $X=4.21 $Y=0.42
+ $X2=0 $Y2=0
cc_360 N_A_369_392#_c_485_n N_A_672_392#_c_686_n 0.00622744f $X=4.21 $Y=0.585
+ $X2=0 $Y2=0
cc_361 N_A_369_392#_c_480_n N_A_672_392#_c_687_n 0.032399f $X=4.21 $Y=0.42 $X2=0
+ $Y2=0
cc_362 N_A_369_392#_c_481_n N_A_672_392#_c_687_n 0.00386148f $X=4.21 $Y=0.42
+ $X2=0 $Y2=0
cc_363 N_A_369_392#_c_484_n N_A_672_392#_c_687_n 0.011037f $X=3.345 $Y=1.47
+ $X2=0 $Y2=0
cc_364 N_A_369_392#_c_485_n N_A_672_392#_c_687_n 0.0132252f $X=4.21 $Y=0.585
+ $X2=0 $Y2=0
cc_365 N_A_369_392#_M1012_g N_A_672_392#_c_699_n 0.0112636f $X=3.27 $Y=2.46
+ $X2=0 $Y2=0
cc_366 N_A_369_392#_c_482_n N_A_672_392#_c_699_n 0.010554f $X=3.345 $Y=1.635
+ $X2=0 $Y2=0
cc_367 N_A_369_392#_c_483_n N_A_672_392#_c_699_n 6.56002e-19 $X=3.345 $Y=1.635
+ $X2=0 $Y2=0
cc_368 N_A_369_392#_M1012_g N_A_672_392#_c_688_n 0.00314789f $X=3.27 $Y=2.46
+ $X2=0 $Y2=0
cc_369 N_A_369_392#_c_482_n N_A_672_392#_c_688_n 0.0382495f $X=3.345 $Y=1.635
+ $X2=0 $Y2=0
cc_370 N_A_369_392#_c_483_n N_A_672_392#_c_688_n 0.00187211f $X=3.345 $Y=1.635
+ $X2=0 $Y2=0
cc_371 N_A_369_392#_c_484_n N_A_672_392#_c_688_n 0.0277249f $X=3.345 $Y=1.47
+ $X2=0 $Y2=0
cc_372 N_A_369_392#_c_485_n N_A_672_392#_c_688_n 2.86089e-19 $X=4.21 $Y=0.585
+ $X2=0 $Y2=0
cc_373 N_A_369_392#_c_488_n N_VPWR_M1018_d 0.00600649f $X=3.18 $Y=1.885 $X2=0
+ $Y2=0
cc_374 N_A_369_392#_M1012_g N_VPWR_c_771_n 0.00333926f $X=3.27 $Y=2.46 $X2=0
+ $Y2=0
cc_375 N_A_369_392#_M1012_g N_VPWR_c_758_n 0.00427637f $X=3.27 $Y=2.46 $X2=0
+ $Y2=0
cc_376 N_A_369_392#_c_488_n A_588_392# 0.00381401f $X=3.18 $Y=1.885 $X2=-0.19
+ $Y2=-0.245
cc_377 N_A_369_392#_c_479_n N_VGND_c_864_n 0.0189626f $X=3.485 $Y=0.42 $X2=0
+ $Y2=0
cc_378 N_A_369_392#_c_484_n N_VGND_c_864_n 0.0183503f $X=3.345 $Y=1.47 $X2=0
+ $Y2=0
cc_379 N_A_369_392#_c_480_n N_VGND_c_865_n 0.0133466f $X=4.21 $Y=0.42 $X2=0
+ $Y2=0
cc_380 N_A_369_392#_c_481_n N_VGND_c_865_n 0.00191229f $X=4.21 $Y=0.42 $X2=0
+ $Y2=0
cc_381 N_A_369_392#_c_479_n N_VGND_c_871_n 0.0121867f $X=3.485 $Y=0.42 $X2=0
+ $Y2=0
cc_382 N_A_369_392#_c_480_n N_VGND_c_871_n 0.0589947f $X=4.21 $Y=0.42 $X2=0
+ $Y2=0
cc_383 N_A_369_392#_c_481_n N_VGND_c_871_n 0.00783549f $X=4.21 $Y=0.42 $X2=0
+ $Y2=0
cc_384 N_A_369_392#_c_479_n N_VGND_c_878_n 0.00660921f $X=3.485 $Y=0.42 $X2=0
+ $Y2=0
cc_385 N_A_369_392#_c_480_n N_VGND_c_878_n 0.0337644f $X=4.21 $Y=0.42 $X2=0
+ $Y2=0
cc_386 N_A_369_392#_c_481_n N_VGND_c_878_n 0.011167f $X=4.21 $Y=0.42 $X2=0 $Y2=0
cc_387 N_A_369_392#_c_484_n A_658_79# 0.00191955f $X=3.345 $Y=1.47 $X2=-0.19
+ $Y2=-0.245
cc_388 N_A_842_405#_M1007_g N_A_672_392#_M1014_g 0.00639596f $X=4.3 $Y=2.725
+ $X2=0 $Y2=0
cc_389 N_A_842_405#_M1006_g N_A_672_392#_M1014_g 0.0281932f $X=4.69 $Y=0.905
+ $X2=0 $Y2=0
cc_390 N_A_842_405#_c_598_n N_A_672_392#_M1014_g 0.0195051f $X=5.25 $Y=2.19
+ $X2=0 $Y2=0
cc_391 N_A_842_405#_c_599_n N_A_672_392#_M1014_g 0.00697018f $X=5.415 $Y=2.355
+ $X2=0 $Y2=0
cc_392 N_A_842_405#_c_600_n N_A_672_392#_M1014_g 0.0169626f $X=5.415 $Y=2.79
+ $X2=0 $Y2=0
cc_393 N_A_842_405#_c_601_n N_A_672_392#_M1014_g 0.00555164f $X=5.59 $Y=1.795
+ $X2=0 $Y2=0
cc_394 N_A_842_405#_M1006_g N_A_672_392#_M1011_g 0.0137357f $X=4.69 $Y=0.905
+ $X2=0 $Y2=0
cc_395 N_A_842_405#_c_590_n N_A_672_392#_M1011_g 0.00180139f $X=5.415 $Y=0.52
+ $X2=0 $Y2=0
cc_396 N_A_842_405#_c_591_n N_A_672_392#_M1011_g 0.00353515f $X=5.59 $Y=1.295
+ $X2=0 $Y2=0
cc_397 N_A_842_405#_M1006_g N_A_672_392#_c_686_n 0.0251514f $X=4.69 $Y=0.905
+ $X2=0 $Y2=0
cc_398 N_A_842_405#_c_588_n N_A_672_392#_c_686_n 3.60437e-19 $X=6.11 $Y=1.46
+ $X2=0 $Y2=0
cc_399 N_A_842_405#_c_598_n N_A_672_392#_c_686_n 0.00911219f $X=5.25 $Y=2.19
+ $X2=0 $Y2=0
cc_400 N_A_842_405#_c_599_n N_A_672_392#_c_686_n 0.0070682f $X=5.415 $Y=2.355
+ $X2=0 $Y2=0
cc_401 N_A_842_405#_c_591_n N_A_672_392#_c_686_n 0.0069888f $X=5.59 $Y=1.295
+ $X2=0 $Y2=0
cc_402 N_A_842_405#_c_593_n N_A_672_392#_c_686_n 0.0281337f $X=5.59 $Y=1.46
+ $X2=0 $Y2=0
cc_403 N_A_842_405#_M1006_g N_A_672_392#_c_687_n 0.00134353f $X=4.69 $Y=0.905
+ $X2=0 $Y2=0
cc_404 N_A_842_405#_M1006_g N_A_672_392#_c_689_n 0.0166985f $X=4.69 $Y=0.905
+ $X2=0 $Y2=0
cc_405 N_A_842_405#_c_588_n N_A_672_392#_c_689_n 0.0182244f $X=6.11 $Y=1.46
+ $X2=0 $Y2=0
cc_406 N_A_842_405#_c_598_n N_A_672_392#_c_689_n 3.97081e-19 $X=5.25 $Y=2.19
+ $X2=0 $Y2=0
cc_407 N_A_842_405#_c_599_n N_A_672_392#_c_689_n 4.3531e-19 $X=5.415 $Y=2.355
+ $X2=0 $Y2=0
cc_408 N_A_842_405#_c_593_n N_A_672_392#_c_689_n 0.00127754f $X=5.59 $Y=1.46
+ $X2=0 $Y2=0
cc_409 N_A_842_405#_c_598_n N_VPWR_M1007_d 0.00913472f $X=5.25 $Y=2.19 $X2=0
+ $Y2=0
cc_410 N_A_842_405#_M1005_g N_VPWR_c_761_n 0.00678238f $X=6.2 $Y=2.4 $X2=0 $Y2=0
cc_411 N_A_842_405#_c_588_n N_VPWR_c_761_n 0.00489956f $X=6.11 $Y=1.46 $X2=0
+ $Y2=0
cc_412 N_A_842_405#_c_599_n N_VPWR_c_761_n 0.0355476f $X=5.415 $Y=2.355 $X2=0
+ $Y2=0
cc_413 N_A_842_405#_c_600_n N_VPWR_c_761_n 0.0345914f $X=5.415 $Y=2.79 $X2=0
+ $Y2=0
cc_414 N_A_842_405#_c_641_p N_VPWR_c_761_n 0.0162042f $X=6.08 $Y=1.46 $X2=0
+ $Y2=0
cc_415 N_A_842_405#_M1019_g N_VPWR_c_763_n 0.00684991f $X=6.695 $Y=2.4 $X2=0
+ $Y2=0
cc_416 N_A_842_405#_c_600_n N_VPWR_c_766_n 0.0132154f $X=5.415 $Y=2.79 $X2=0
+ $Y2=0
cc_417 N_A_842_405#_M1005_g N_VPWR_c_769_n 0.00523177f $X=6.2 $Y=2.4 $X2=0 $Y2=0
cc_418 N_A_842_405#_M1019_g N_VPWR_c_769_n 0.00523177f $X=6.695 $Y=2.4 $X2=0
+ $Y2=0
cc_419 N_A_842_405#_M1007_g N_VPWR_c_771_n 0.00558361f $X=4.3 $Y=2.725 $X2=0
+ $Y2=0
cc_420 N_A_842_405#_M1007_g N_VPWR_c_772_n 0.00874065f $X=4.3 $Y=2.725 $X2=0
+ $Y2=0
cc_421 N_A_842_405#_c_598_n N_VPWR_c_772_n 0.0383579f $X=5.25 $Y=2.19 $X2=0
+ $Y2=0
cc_422 N_A_842_405#_c_600_n N_VPWR_c_772_n 0.0132969f $X=5.415 $Y=2.79 $X2=0
+ $Y2=0
cc_423 N_A_842_405#_c_602_n N_VPWR_c_772_n 0.00856791f $X=4.69 $Y=2.19 $X2=0
+ $Y2=0
cc_424 N_A_842_405#_M1007_g N_VPWR_c_758_n 0.00537853f $X=4.3 $Y=2.725 $X2=0
+ $Y2=0
cc_425 N_A_842_405#_M1005_g N_VPWR_c_758_n 0.00990289f $X=6.2 $Y=2.4 $X2=0 $Y2=0
cc_426 N_A_842_405#_M1019_g N_VPWR_c_758_n 0.00988898f $X=6.695 $Y=2.4 $X2=0
+ $Y2=0
cc_427 N_A_842_405#_c_600_n N_VPWR_c_758_n 0.0119049f $X=5.415 $Y=2.79 $X2=0
+ $Y2=0
cc_428 N_A_842_405#_M1000_g N_Q_c_841_n 5.5543e-19 $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_429 N_A_842_405#_M1010_g N_Q_c_841_n 0.00487958f $X=6.68 $Y=0.74 $X2=0 $Y2=0
cc_430 N_A_842_405#_c_589_n N_Q_c_842_n 0.00276508f $X=6.68 $Y=1.46 $X2=0 $Y2=0
cc_431 N_A_842_405#_M1005_g Q 0.022085f $X=6.2 $Y=2.4 $X2=0 $Y2=0
cc_432 N_A_842_405#_M1019_g Q 0.022085f $X=6.695 $Y=2.4 $X2=0 $Y2=0
cc_433 N_A_842_405#_c_589_n Q 0.00136087f $X=6.68 $Y=1.46 $X2=0 $Y2=0
cc_434 N_A_842_405#_M1005_g N_Q_c_843_n 0.00512371f $X=6.2 $Y=2.4 $X2=0 $Y2=0
cc_435 N_A_842_405#_M1000_g N_Q_c_843_n 0.00369108f $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_436 N_A_842_405#_M1019_g N_Q_c_843_n 0.00544497f $X=6.695 $Y=2.4 $X2=0 $Y2=0
cc_437 N_A_842_405#_c_589_n N_Q_c_843_n 0.0273845f $X=6.68 $Y=1.46 $X2=0 $Y2=0
cc_438 N_A_842_405#_c_641_p N_Q_c_843_n 0.0249855f $X=6.08 $Y=1.46 $X2=0 $Y2=0
cc_439 N_A_842_405#_M1006_g N_VGND_c_865_n 0.00480566f $X=4.69 $Y=0.905 $X2=0
+ $Y2=0
cc_440 N_A_842_405#_c_590_n N_VGND_c_865_n 0.0229496f $X=5.415 $Y=0.52 $X2=0
+ $Y2=0
cc_441 N_A_842_405#_M1000_g N_VGND_c_866_n 0.014912f $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_442 N_A_842_405#_M1010_g N_VGND_c_866_n 5.38476e-19 $X=6.68 $Y=0.74 $X2=0
+ $Y2=0
cc_443 N_A_842_405#_c_588_n N_VGND_c_866_n 0.006266f $X=6.11 $Y=1.46 $X2=0 $Y2=0
cc_444 N_A_842_405#_c_590_n N_VGND_c_866_n 0.0346502f $X=5.415 $Y=0.52 $X2=0
+ $Y2=0
cc_445 N_A_842_405#_c_641_p N_VGND_c_866_n 0.0245638f $X=6.08 $Y=1.46 $X2=0
+ $Y2=0
cc_446 N_A_842_405#_c_592_n N_VGND_c_866_n 0.0138526f $X=5.502 $Y=1.125 $X2=0
+ $Y2=0
cc_447 N_A_842_405#_M1010_g N_VGND_c_868_n 0.00553267f $X=6.68 $Y=0.74 $X2=0
+ $Y2=0
cc_448 N_A_842_405#_c_589_n N_VGND_c_868_n 0.00120202f $X=6.68 $Y=1.46 $X2=0
+ $Y2=0
cc_449 N_A_842_405#_M1006_g N_VGND_c_871_n 0.00380268f $X=4.69 $Y=0.905 $X2=0
+ $Y2=0
cc_450 N_A_842_405#_c_590_n N_VGND_c_872_n 0.0108483f $X=5.415 $Y=0.52 $X2=0
+ $Y2=0
cc_451 N_A_842_405#_M1000_g N_VGND_c_873_n 0.00383152f $X=6.19 $Y=0.74 $X2=0
+ $Y2=0
cc_452 N_A_842_405#_M1010_g N_VGND_c_873_n 0.00460063f $X=6.68 $Y=0.74 $X2=0
+ $Y2=0
cc_453 N_A_842_405#_M1006_g N_VGND_c_878_n 0.0045051f $X=4.69 $Y=0.905 $X2=0
+ $Y2=0
cc_454 N_A_842_405#_M1000_g N_VGND_c_878_n 0.00758109f $X=6.19 $Y=0.74 $X2=0
+ $Y2=0
cc_455 N_A_842_405#_M1010_g N_VGND_c_878_n 0.0091141f $X=6.68 $Y=0.74 $X2=0
+ $Y2=0
cc_456 N_A_842_405#_c_590_n N_VGND_c_878_n 0.00913189f $X=5.415 $Y=0.52 $X2=0
+ $Y2=0
cc_457 N_A_672_392#_M1014_g N_VPWR_c_761_n 0.0046118f $X=5.19 $Y=2.375 $X2=0
+ $Y2=0
cc_458 N_A_672_392#_M1014_g N_VPWR_c_766_n 0.00640648f $X=5.19 $Y=2.375 $X2=0
+ $Y2=0
cc_459 N_A_672_392#_M1014_g N_VPWR_c_772_n 0.00451287f $X=5.19 $Y=2.375 $X2=0
+ $Y2=0
cc_460 N_A_672_392#_M1014_g N_VPWR_c_758_n 0.00645424f $X=5.19 $Y=2.375 $X2=0
+ $Y2=0
cc_461 N_A_672_392#_M1011_g N_VGND_c_865_n 0.014975f $X=5.2 $Y=0.745 $X2=0 $Y2=0
cc_462 N_A_672_392#_c_686_n N_VGND_c_865_n 0.0253469f $X=4.99 $Y=1.23 $X2=0
+ $Y2=0
cc_463 N_A_672_392#_c_689_n N_VGND_c_865_n 5.31358e-19 $X=5.17 $Y=1.46 $X2=0
+ $Y2=0
cc_464 N_A_672_392#_M1011_g N_VGND_c_866_n 0.0039491f $X=5.2 $Y=0.745 $X2=0
+ $Y2=0
cc_465 N_A_672_392#_M1011_g N_VGND_c_872_n 0.00379792f $X=5.2 $Y=0.745 $X2=0
+ $Y2=0
cc_466 N_A_672_392#_M1011_g N_VGND_c_878_n 0.00457201f $X=5.2 $Y=0.745 $X2=0
+ $Y2=0
cc_467 N_VPWR_c_769_n Q 0.01003f $X=6.835 $Y=3.33 $X2=0 $Y2=0
cc_468 N_VPWR_c_758_n Q 0.0127021f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_469 N_VPWR_c_761_n N_Q_c_843_n 0.00256271f $X=5.975 $Y=1.985 $X2=0 $Y2=0
cc_470 N_VPWR_c_763_n N_Q_c_843_n 0.00112461f $X=6.92 $Y=1.985 $X2=0 $Y2=0
cc_471 N_Q_c_841_n N_VGND_c_866_n 0.0285797f $X=6.41 $Y=0.515 $X2=0 $Y2=0
cc_472 N_Q_c_841_n N_VGND_c_868_n 0.0313502f $X=6.41 $Y=0.515 $X2=0 $Y2=0
cc_473 N_Q_c_841_n N_VGND_c_873_n 0.0117353f $X=6.41 $Y=0.515 $X2=0 $Y2=0
cc_474 N_Q_c_841_n N_VGND_c_878_n 0.00971347f $X=6.41 $Y=0.515 $X2=0 $Y2=0

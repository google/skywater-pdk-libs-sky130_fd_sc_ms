* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_163_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X1 VPWR a_247_368# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X2 VGND a_247_368# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_54_74# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_54_74# B1 a_247_368# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 X a_247_368# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 X a_247_368# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 a_163_368# A2 a_247_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X8 a_247_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X9 VGND A2 a_54_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__dlclkp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__dlclkp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN GATE
    ANTENNAGATEAREA  0.276000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.450000 1.335000 1.780000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.805000 0.440000 7.135000 2.980000 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.553200 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 4.550000 1.445000 5.220000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.680000 0.085000 ;
        RECT 0.545000  0.085000 0.880000 0.600000 ;
        RECT 2.920000  0.755000 3.535000 1.005000 ;
        RECT 3.340000  0.085000 3.535000 0.755000 ;
        RECT 4.765000  0.085000 5.095000 1.275000 ;
        RECT 6.305000  0.085000 6.635000 0.770000 ;
        RECT 7.315000  0.085000 7.565000 1.220000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 7.680000 3.415000 ;
        RECT 0.685000 2.290000 1.075000 3.245000 ;
        RECT 2.945000 2.650000 3.485000 3.245000 ;
        RECT 4.715000 2.075000 5.045000 3.245000 ;
        RECT 5.730000 1.950000 6.635000 3.245000 ;
        RECT 7.315000 1.820000 7.565000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 0.350000 0.365000 0.770000 ;
      RECT 0.095000 0.770000 1.220000 0.940000 ;
      RECT 0.095000 0.940000 0.265000 1.820000 ;
      RECT 0.095000 1.820000 0.445000 2.980000 ;
      RECT 0.435000 1.110000 1.560000 1.280000 ;
      RECT 0.435000 1.280000 0.785000 1.550000 ;
      RECT 0.615000 1.550000 0.785000 1.950000 ;
      RECT 0.615000 1.950000 1.705000 2.120000 ;
      RECT 1.050000 0.255000 3.160000 0.425000 ;
      RECT 1.050000 0.425000 1.220000 0.770000 ;
      RECT 1.390000 0.620000 2.245000 0.950000 ;
      RECT 1.390000 0.950000 1.560000 1.110000 ;
      RECT 1.535000 2.120000 1.705000 2.550000 ;
      RECT 1.535000 2.550000 2.405000 2.880000 ;
      RECT 1.730000 1.120000 2.045000 1.450000 ;
      RECT 1.875000 1.450000 2.045000 2.050000 ;
      RECT 1.875000 2.050000 3.325000 2.220000 ;
      RECT 2.225000 2.220000 2.555000 2.380000 ;
      RECT 2.255000 1.215000 4.035000 1.385000 ;
      RECT 2.255000 1.385000 2.585000 1.840000 ;
      RECT 2.830000 0.425000 3.160000 0.585000 ;
      RECT 3.155000 1.555000 3.485000 1.885000 ;
      RECT 3.155000 1.885000 3.325000 2.050000 ;
      RECT 3.655000 1.385000 3.825000 2.100000 ;
      RECT 3.655000 2.100000 3.985000 2.980000 ;
      RECT 3.705000 0.605000 4.035000 1.215000 ;
      RECT 3.995000 1.555000 4.380000 1.885000 ;
      RECT 4.210000 0.575000 4.595000 1.275000 ;
      RECT 4.210000 1.275000 4.380000 1.555000 ;
      RECT 4.210000 1.885000 4.380000 2.075000 ;
      RECT 4.210000 2.075000 4.545000 2.955000 ;
      RECT 5.215000 1.950000 5.560000 2.955000 ;
      RECT 5.390000 0.940000 6.305000 1.610000 ;
      RECT 5.390000 1.610000 5.560000 1.950000 ;
      RECT 5.555000 0.575000 5.885000 0.940000 ;
  END
END sky130_fd_sc_ms__dlclkp_2

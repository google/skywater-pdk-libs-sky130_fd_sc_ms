* File: sky130_fd_sc_ms__nor2b_1.pxi.spice
* Created: Fri Aug 28 17:47:21 2020
* 
x_PM_SKY130_FD_SC_MS__NOR2B_1%B_N N_B_N_M1003_g N_B_N_c_43_n N_B_N_M1004_g
+ N_B_N_c_44_n N_B_N_c_45_n B_N PM_SKY130_FD_SC_MS__NOR2B_1%B_N
x_PM_SKY130_FD_SC_MS__NOR2B_1%A N_A_M1000_g N_A_M1005_g A N_A_c_75_n N_A_c_76_n
+ PM_SKY130_FD_SC_MS__NOR2B_1%A
x_PM_SKY130_FD_SC_MS__NOR2B_1%A_27_112# N_A_27_112#_M1004_s N_A_27_112#_M1003_s
+ N_A_27_112#_M1001_g N_A_27_112#_M1002_g N_A_27_112#_c_119_n
+ N_A_27_112#_c_114_n N_A_27_112#_c_110_n N_A_27_112#_c_116_n
+ N_A_27_112#_c_117_n N_A_27_112#_c_111_n N_A_27_112#_c_112_n
+ PM_SKY130_FD_SC_MS__NOR2B_1%A_27_112#
x_PM_SKY130_FD_SC_MS__NOR2B_1%VPWR N_VPWR_M1003_d N_VPWR_c_179_n VPWR
+ N_VPWR_c_180_n N_VPWR_c_181_n N_VPWR_c_178_n N_VPWR_c_183_n
+ PM_SKY130_FD_SC_MS__NOR2B_1%VPWR
x_PM_SKY130_FD_SC_MS__NOR2B_1%Y N_Y_M1005_d N_Y_M1001_d N_Y_c_203_n N_Y_c_204_n
+ N_Y_c_205_n Y Y Y N_Y_c_208_n N_Y_c_206_n Y PM_SKY130_FD_SC_MS__NOR2B_1%Y
x_PM_SKY130_FD_SC_MS__NOR2B_1%VGND N_VGND_M1004_d N_VGND_M1002_d N_VGND_c_236_n
+ N_VGND_c_237_n N_VGND_c_238_n N_VGND_c_239_n N_VGND_c_240_n VGND
+ N_VGND_c_241_n N_VGND_c_242_n PM_SKY130_FD_SC_MS__NOR2B_1%VGND
cc_1 VNB N_B_N_c_43_n 0.0233618f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.22
cc_2 VNB N_B_N_c_44_n 0.0628724f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.385
cc_3 VNB N_B_N_c_45_n 0.0198916f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.22
cc_4 VNB B_N 0.017759f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_5 VNB N_A_M1000_g 0.00668999f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.26
cc_6 VNB A 0.00407508f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.385
cc_7 VNB N_A_c_75_n 0.0370951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_c_76_n 0.0201157f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.385
cc_9 VNB N_A_27_112#_M1001_g 5.03068e-19 $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.22
cc_10 VNB N_A_27_112#_M1002_g 0.0253088f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.385
cc_11 VNB N_A_27_112#_c_110_n 0.00853715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_112#_c_111_n 0.0111198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_112#_c_112_n 0.0342437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_VPWR_c_178_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_Y_c_203_n 0.00208979f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.22
cc_16 VNB N_Y_c_204_n 0.012465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_205_n 0.00221952f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.385
cc_18 VNB N_Y_c_206_n 0.0242534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_236_n 0.0131348f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.22
cc_20 VNB N_VGND_c_237_n 0.0129133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_238_n 0.011907f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.385
cc_22 VNB N_VGND_c_239_n 0.0302402f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.295
cc_23 VNB N_VGND_c_240_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_241_n 0.0193208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_242_n 0.178959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VPB N_B_N_M1003_g 0.0263115f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=2.26
cc_27 VPB N_B_N_c_45_n 0.00288981f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.22
cc_28 VPB N_A_M1000_g 0.0238494f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=2.26
cc_29 VPB N_A_27_112#_M1001_g 0.026483f $X=-0.19 $Y=1.66 $X2=0.615 $Y2=1.22
cc_30 VPB N_A_27_112#_c_114_n 0.0346733f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_31 VPB N_A_27_112#_c_110_n 0.00202686f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB N_A_27_112#_c_116_n 0.0141291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_33 VPB N_A_27_112#_c_117_n 0.0101533f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_A_27_112#_c_111_n 5.62371e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_179_n 0.0169832f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.835
cc_36 VPB N_VPWR_c_180_n 0.0300706f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=1.385
cc_37 VPB N_VPWR_c_181_n 0.0349999f $X=-0.19 $Y=1.66 $X2=0.275 $Y2=1.385
cc_38 VPB N_VPWR_c_178_n 0.0795025f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_183_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB Y 0.0448941f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_Y_c_208_n 0.0129651f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_Y_c_206_n 0.0078509f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 N_B_N_c_45_n N_A_M1000_g 0.0197372f $X=0.615 $Y=1.22 $X2=0 $Y2=0
cc_44 N_B_N_c_43_n A 3.04755e-19 $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_45 N_B_N_c_45_n A 8.64176e-19 $X=0.615 $Y=1.22 $X2=0 $Y2=0
cc_46 N_B_N_c_45_n N_A_c_75_n 0.0166901f $X=0.615 $Y=1.22 $X2=0 $Y2=0
cc_47 N_B_N_c_43_n N_A_c_76_n 0.0094315f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_48 N_B_N_c_43_n N_A_27_112#_c_119_n 0.00851666f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_49 N_B_N_c_44_n N_A_27_112#_c_119_n 0.00741677f $X=0.615 $Y=1.385 $X2=0 $Y2=0
cc_50 B_N N_A_27_112#_c_119_n 0.0152451f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_51 N_B_N_M1003_g N_A_27_112#_c_114_n 0.0167241f $X=0.705 $Y=2.26 $X2=0 $Y2=0
cc_52 N_B_N_M1003_g N_A_27_112#_c_110_n 7.94248e-19 $X=0.705 $Y=2.26 $X2=0 $Y2=0
cc_53 N_B_N_c_43_n N_A_27_112#_c_110_n 0.00809053f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_54 N_B_N_c_44_n N_A_27_112#_c_110_n 0.0046103f $X=0.615 $Y=1.385 $X2=0 $Y2=0
cc_55 N_B_N_c_45_n N_A_27_112#_c_110_n 0.0134498f $X=0.615 $Y=1.22 $X2=0 $Y2=0
cc_56 B_N N_A_27_112#_c_110_n 0.026737f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_57 N_B_N_M1003_g N_A_27_112#_c_116_n 0.00374172f $X=0.705 $Y=2.26 $X2=0 $Y2=0
cc_58 N_B_N_M1003_g N_A_27_112#_c_117_n 0.0119883f $X=0.705 $Y=2.26 $X2=0 $Y2=0
cc_59 N_B_N_c_44_n N_A_27_112#_c_117_n 0.00858089f $X=0.615 $Y=1.385 $X2=0 $Y2=0
cc_60 B_N N_A_27_112#_c_117_n 0.0105909f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_61 N_B_N_M1003_g N_VPWR_c_179_n 0.00919593f $X=0.705 $Y=2.26 $X2=0 $Y2=0
cc_62 N_B_N_M1003_g N_VPWR_c_180_n 0.00465228f $X=0.705 $Y=2.26 $X2=0 $Y2=0
cc_63 N_B_N_M1003_g N_VPWR_c_178_n 0.00555093f $X=0.705 $Y=2.26 $X2=0 $Y2=0
cc_64 N_B_N_c_43_n N_VGND_c_236_n 0.00905753f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_65 N_B_N_c_43_n N_VGND_c_239_n 0.00360585f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_66 N_B_N_c_43_n N_VGND_c_242_n 0.00487769f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_67 N_A_M1000_g N_A_27_112#_M1001_g 0.0462713f $X=1.315 $Y=2.4 $X2=0 $Y2=0
cc_68 A N_A_27_112#_M1002_g 7.63572e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_69 N_A_c_76_n N_A_27_112#_M1002_g 0.0219036f $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_70 N_A_M1000_g N_A_27_112#_c_114_n 4.84573e-19 $X=1.315 $Y=2.4 $X2=0 $Y2=0
cc_71 N_A_M1000_g N_A_27_112#_c_110_n 0.00158717f $X=1.315 $Y=2.4 $X2=0 $Y2=0
cc_72 A N_A_27_112#_c_110_n 0.0199505f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_73 N_A_c_75_n N_A_27_112#_c_110_n 0.00164547f $X=1.2 $Y=1.385 $X2=0 $Y2=0
cc_74 N_A_c_76_n N_A_27_112#_c_110_n 6.54906e-19 $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_75 N_A_M1000_g N_A_27_112#_c_116_n 0.0180507f $X=1.315 $Y=2.4 $X2=0 $Y2=0
cc_76 A N_A_27_112#_c_116_n 0.0244703f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_77 N_A_c_75_n N_A_27_112#_c_116_n 0.00133235f $X=1.2 $Y=1.385 $X2=0 $Y2=0
cc_78 A N_A_27_112#_c_111_n 0.0187161f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_79 N_A_c_75_n N_A_27_112#_c_111_n 0.00565605f $X=1.2 $Y=1.385 $X2=0 $Y2=0
cc_80 A N_A_27_112#_c_112_n 2.21841e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_81 N_A_c_75_n N_A_27_112#_c_112_n 0.0462713f $X=1.2 $Y=1.385 $X2=0 $Y2=0
cc_82 N_A_M1000_g N_VPWR_c_179_n 0.0238204f $X=1.315 $Y=2.4 $X2=0 $Y2=0
cc_83 N_A_M1000_g N_VPWR_c_181_n 0.00460063f $X=1.315 $Y=2.4 $X2=0 $Y2=0
cc_84 N_A_M1000_g N_VPWR_c_178_n 0.00908371f $X=1.315 $Y=2.4 $X2=0 $Y2=0
cc_85 N_A_c_76_n N_Y_c_203_n 0.00516456f $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_86 N_A_c_76_n N_Y_c_205_n 0.00443842f $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_87 A N_VGND_c_236_n 0.0185651f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_88 N_A_c_75_n N_VGND_c_236_n 0.00139293f $X=1.2 $Y=1.385 $X2=0 $Y2=0
cc_89 N_A_c_76_n N_VGND_c_236_n 0.0139704f $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_90 N_A_c_76_n N_VGND_c_241_n 0.00383152f $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_91 N_A_c_76_n N_VGND_c_242_n 0.00758292f $X=1.22 $Y=1.22 $X2=0 $Y2=0
cc_92 N_A_27_112#_c_116_n N_VPWR_M1003_d 0.00558587f $X=1.535 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_93 N_A_27_112#_M1001_g N_VPWR_c_179_n 0.0032432f $X=1.735 $Y=2.4 $X2=0 $Y2=0
cc_94 N_A_27_112#_c_114_n N_VPWR_c_179_n 0.0339227f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_95 N_A_27_112#_c_116_n N_VPWR_c_179_n 0.0218557f $X=1.535 $Y=1.805 $X2=0
+ $Y2=0
cc_96 N_A_27_112#_c_114_n N_VPWR_c_180_n 0.0066444f $X=0.48 $Y=1.985 $X2=0 $Y2=0
cc_97 N_A_27_112#_M1001_g N_VPWR_c_181_n 0.00553757f $X=1.735 $Y=2.4 $X2=0 $Y2=0
cc_98 N_A_27_112#_M1001_g N_VPWR_c_178_n 0.0109376f $X=1.735 $Y=2.4 $X2=0 $Y2=0
cc_99 N_A_27_112#_c_114_n N_VPWR_c_178_n 0.00995531f $X=0.48 $Y=1.985 $X2=0
+ $Y2=0
cc_100 N_A_27_112#_c_116_n A_281_368# 0.0027472f $X=1.535 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_101 N_A_27_112#_c_111_n A_281_368# 0.00234086f $X=1.81 $Y=1.485 $X2=-0.19
+ $Y2=-0.245
cc_102 N_A_27_112#_M1002_g N_Y_c_203_n 0.0130905f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_103 N_A_27_112#_M1002_g N_Y_c_204_n 0.0127588f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_104 N_A_27_112#_c_111_n N_Y_c_204_n 0.0138485f $X=1.81 $Y=1.485 $X2=0 $Y2=0
cc_105 N_A_27_112#_c_112_n N_Y_c_204_n 4.58216e-19 $X=1.81 $Y=1.485 $X2=0 $Y2=0
cc_106 N_A_27_112#_M1002_g N_Y_c_205_n 0.00116669f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_107 N_A_27_112#_c_111_n N_Y_c_205_n 0.0221208f $X=1.81 $Y=1.485 $X2=0 $Y2=0
cc_108 N_A_27_112#_c_112_n N_Y_c_205_n 8.9933e-19 $X=1.81 $Y=1.485 $X2=0 $Y2=0
cc_109 N_A_27_112#_M1001_g N_Y_c_208_n 0.00207194f $X=1.735 $Y=2.4 $X2=0 $Y2=0
cc_110 N_A_27_112#_c_111_n N_Y_c_208_n 0.0121675f $X=1.81 $Y=1.485 $X2=0 $Y2=0
cc_111 N_A_27_112#_c_112_n N_Y_c_208_n 7.80347e-19 $X=1.81 $Y=1.485 $X2=0 $Y2=0
cc_112 N_A_27_112#_M1001_g N_Y_c_206_n 0.00318862f $X=1.735 $Y=2.4 $X2=0 $Y2=0
cc_113 N_A_27_112#_M1002_g N_Y_c_206_n 0.00539566f $X=1.835 $Y=0.74 $X2=0 $Y2=0
cc_114 N_A_27_112#_c_111_n N_Y_c_206_n 0.0318104f $X=1.81 $Y=1.485 $X2=0 $Y2=0
cc_115 N_A_27_112#_c_112_n N_Y_c_206_n 0.00232633f $X=1.81 $Y=1.485 $X2=0 $Y2=0
cc_116 N_A_27_112#_M1002_g N_VGND_c_236_n 6.08003e-19 $X=1.835 $Y=0.74 $X2=0
+ $Y2=0
cc_117 N_A_27_112#_c_119_n N_VGND_c_236_n 0.02666f $X=0.61 $Y=0.845 $X2=0 $Y2=0
cc_118 N_A_27_112#_M1002_g N_VGND_c_238_n 0.00521557f $X=1.835 $Y=0.74 $X2=0
+ $Y2=0
cc_119 N_A_27_112#_c_119_n N_VGND_c_239_n 0.00820401f $X=0.61 $Y=0.845 $X2=0
+ $Y2=0
cc_120 N_A_27_112#_M1002_g N_VGND_c_241_n 0.00434272f $X=1.835 $Y=0.74 $X2=0
+ $Y2=0
cc_121 N_A_27_112#_M1002_g N_VGND_c_242_n 0.00824687f $X=1.835 $Y=0.74 $X2=0
+ $Y2=0
cc_122 N_A_27_112#_c_119_n N_VGND_c_242_n 0.0148718f $X=0.61 $Y=0.845 $X2=0
+ $Y2=0
cc_123 N_VPWR_c_179_n Y 0.0121179f $X=1.09 $Y=2.145 $X2=0 $Y2=0
cc_124 N_VPWR_c_181_n Y 0.019544f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_125 N_VPWR_c_178_n Y 0.0161768f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_126 N_Y_c_204_n N_VGND_M1002_d 0.00568412f $X=2.145 $Y=1.065 $X2=0 $Y2=0
cc_127 N_Y_c_203_n N_VGND_c_236_n 0.0350754f $X=1.62 $Y=0.515 $X2=0 $Y2=0
cc_128 N_Y_c_205_n N_VGND_c_236_n 0.00181371f $X=1.785 $Y=1.065 $X2=0 $Y2=0
cc_129 N_Y_c_203_n N_VGND_c_238_n 0.0173103f $X=1.62 $Y=0.515 $X2=0 $Y2=0
cc_130 N_Y_c_204_n N_VGND_c_238_n 0.0220189f $X=2.145 $Y=1.065 $X2=0 $Y2=0
cc_131 N_Y_c_203_n N_VGND_c_241_n 0.0109942f $X=1.62 $Y=0.515 $X2=0 $Y2=0
cc_132 N_Y_c_203_n N_VGND_c_242_n 0.00904371f $X=1.62 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__a21boi_4.spice
* Created: Wed Sep  2 11:51:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a21boi_4.pex.spice"
.subckt sky130_fd_sc_ms__a21boi_4  VNB VPB A1 A2 B1_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1_N	B1_N
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1003 N_A_46_74#_M1003_d N_A1_M1003_g N_Y_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1005 N_A_46_74#_M1005_d N_A1_M1005_g N_Y_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1006 N_A_46_74#_M1005_d N_A1_M1006_g N_Y_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1015 N_A_46_74#_M1015_d N_A1_M1015_g N_Y_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1002 N_A_46_74#_M1015_d N_A2_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1011 N_A_46_74#_M1011_d N_A2_M1011_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1012 N_A_46_74#_M1011_d N_A2_M1012_g N_VGND_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1023 N_A_46_74#_M1023_d N_A2_M1023_g N_VGND_M1012_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_A_803_323#_M1000_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1013_d N_A_803_323#_M1013_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1013_d N_A_803_323#_M1021_g N_Y_M1021_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1024 N_VGND_M1024_d N_A_803_323#_M1024_g N_Y_M1021_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1004 N_A_803_323#_M1004_d N_B1_N_M1004_g N_VGND_M1024_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g N_A_31_368#_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90005.1 A=0.2016 P=2.6 MULT=1
MM1009 N_VPWR_M1008_d N_A1_M1009_g N_A_31_368#_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90004.7 A=0.2016 P=2.6 MULT=1
MM1010 N_VPWR_M1010_d N_A1_M1010_g N_A_31_368#_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90004.2 A=0.2016 P=2.6 MULT=1
MM1014 N_VPWR_M1010_d N_A1_M1014_g N_A_31_368#_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90003.8 A=0.2016 P=2.6 MULT=1
MM1016 N_VPWR_M1016_d N_A2_M1016_g N_A_31_368#_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90003.3 A=0.2016 P=2.6 MULT=1
MM1018 N_VPWR_M1016_d N_A2_M1018_g N_A_31_368#_M1018_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.4
+ SB=90002.9 A=0.2016 P=2.6 MULT=1
MM1020 N_VPWR_M1020_d N_A2_M1020_g N_A_31_368#_M1018_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.9
+ SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1022 N_VPWR_M1020_d N_A2_M1022_g N_A_31_368#_M1022_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.3
+ SB=90002 A=0.2016 P=2.6 MULT=1
MM1001 N_Y_M1001_d N_A_803_323#_M1001_g N_A_31_368#_M1022_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90003.8 SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1007 N_Y_M1001_d N_A_803_323#_M1007_g N_A_31_368#_M1007_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90004.2 SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1025 N_Y_M1025_d N_A_803_323#_M1025_g N_A_31_368#_M1007_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90004.7 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1026 N_Y_M1025_d N_A_803_323#_M1026_g N_A_31_368#_M1026_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90005.1 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1017 N_A_803_323#_M1017_d N_B1_N_M1017_g N_VPWR_M1017_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1134 AS=0.2184 PD=1.11 PS=2.2 NRD=0 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.6 A=0.1512 P=2.04 MULT=1
MM1019 N_A_803_323#_M1017_d N_B1_N_M1019_g N_VPWR_M1019_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1134 AS=0.2184 PD=1.11 PS=2.2 NRD=0 NRS=0 M=1 R=4.66667 SA=90000.6
+ SB=90000.2 A=0.1512 P=2.04 MULT=1
DX27_noxref VNB VPB NWDIODE A=14.9916 P=19.84
c_59 VNB 0 1.93315e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__a21boi_4.pxi.spice"
*
.ends
*
*

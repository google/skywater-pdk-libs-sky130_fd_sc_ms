* File: sky130_fd_sc_ms__dfrtp_2.pex.spice
* Created: Wed Sep  2 12:03:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DFRTP_2%D 2 5 9 11 12 13 18 19 22
c31 5 0 1.98761e-19 $X=0.495 $Y=2.845
r32 22 24 40.9207 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.845
+ $X2=0.402 $Y2=2.01
r33 22 23 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.845 $X2=0.385 $Y2=1.845
r34 18 20 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.165
+ $X2=0.402 $Y2=1
r35 18 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.165 $X2=0.385 $Y2=1.165
r36 13 23 5.91795 $w=3.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.31 $Y=2.035
+ $X2=0.31 $Y2=1.845
r37 12 23 5.60648 $w=3.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.31 $Y=1.665
+ $X2=0.31 $Y2=1.845
r38 11 12 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.31 $Y=1.295
+ $X2=0.31 $Y2=1.665
r39 11 19 4.04912 $w=3.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.31 $Y=1.295
+ $X2=0.31 $Y2=1.165
r40 9 20 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.51 $Y=0.6 $X2=0.51
+ $Y2=1
r41 5 24 324.573 $w=1.8e-07 $l=8.35e-07 $layer=POLY_cond $X=0.495 $Y=2.845
+ $X2=0.495 $Y2=2.01
r42 2 22 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=0.402 $Y=1.828
+ $X2=0.402 $Y2=1.845
r43 1 18 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=0.402 $Y=1.182
+ $X2=0.402 $Y2=1.165
r44 1 2 102.129 $w=3.65e-07 $l=6.46e-07 $layer=POLY_cond $X=0.402 $Y=1.182
+ $X2=0.402 $Y2=1.828
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_2%CLK 3 6 8 11 13
c45 11 0 6.1174e-20 $X=1.91 $Y=1.61
c46 8 0 1.39258e-19 $X=2.16 $Y=1.665
r47 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.91 $Y=1.61
+ $X2=1.91 $Y2=1.775
r48 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.91 $Y=1.61
+ $X2=1.91 $Y2=1.445
r49 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.91
+ $Y=1.61 $X2=1.91 $Y2=1.61
r50 8 12 6.67396 $w=4.57e-07 $l=2.5e-07 $layer=LI1_cond $X=2.16 $Y=1.55 $X2=1.91
+ $Y2=1.55
r51 6 14 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.925 $Y=2.495
+ $X2=1.925 $Y2=1.775
r52 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.89 $Y=0.965 $X2=1.89
+ $Y2=1.445
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_2%A_493_387# 1 2 7 9 11 13 15 17 19 20 21 24
+ 28 29 31 33 36 39 40 41 44 48 49 57 63 66 76
c197 44 0 1.33493e-19 $X=7.12 $Y=2.14
c198 31 0 1.39258e-19 $X=3.08 $Y=1.77
c199 29 0 7.88206e-20 $X=4.27 $Y=0.415
c200 21 0 4.38853e-20 $X=6.355 $Y=1.27
c201 15 0 8.97095e-20 $X=4.01 $Y=0.9
c202 7 0 8.96654e-20 $X=3.405 $Y=1.935
r203 65 66 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=7.12 $Y=1.18
+ $X2=7.37 $Y2=1.18
r204 63 72 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.88 $Y=1.18 $X2=6.88
+ $Y2=1.27
r205 62 65 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=6.88 $Y=1.18
+ $X2=7.12 $Y2=1.18
r206 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.88
+ $Y=1.18 $X2=6.88 $Y2=1.18
r207 57 59 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.355 $Y=0.415
+ $X2=4.355 $Y2=0.7
r208 52 53 7.89897 $w=5.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=0.725
+ $X2=2.775 $Y2=0.81
r209 49 52 6.99593 $w=5.28e-07 $l=3.1e-07 $layer=LI1_cond $X=2.775 $Y=0.415
+ $X2=2.775 $Y2=0.725
r210 48 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.37 $Y=1.015
+ $X2=7.37 $Y2=1.18
r211 47 48 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.37 $Y=0.425
+ $X2=7.37 $Y2=1.015
r212 45 76 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=7.12 $Y=2.14
+ $X2=7.315 $Y2=2.14
r213 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.12
+ $Y=2.14 $X2=7.12 $Y2=2.14
r214 42 65 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.12 $Y=1.345
+ $X2=7.12 $Y2=1.18
r215 42 44 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=7.12 $Y=1.345
+ $X2=7.12 $Y2=2.14
r216 40 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.285 $Y=0.34
+ $X2=7.37 $Y2=0.425
r217 40 41 104.385 $w=1.68e-07 $l=1.6e-06 $layer=LI1_cond $X=7.285 $Y=0.34
+ $X2=5.685 $Y2=0.34
r218 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.6 $Y=0.425
+ $X2=5.685 $Y2=0.34
r219 38 39 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.6 $Y=0.425
+ $X2=5.6 $Y2=0.615
r220 37 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.44 $Y=0.7
+ $X2=4.355 $Y2=0.7
r221 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.515 $Y=0.7
+ $X2=5.6 $Y2=0.615
r222 36 37 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=5.515 $Y=0.7
+ $X2=4.44 $Y2=0.7
r223 34 68 13.2256 $w=3.28e-07 $l=9e-08 $layer=POLY_cond $X=3.33 $Y=1.77
+ $X2=3.33 $Y2=1.68
r224 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.33
+ $Y=1.77 $X2=3.33 $Y2=1.77
r225 31 56 11.1806 $w=3.71e-07 $l=5.54527e-07 $layer=LI1_cond $X=3.08 $Y=1.77
+ $X2=2.67 $Y2=2.11
r226 31 33 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.08 $Y=1.77
+ $X2=3.33 $Y2=1.77
r227 30 49 7.52407 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=3.04 $Y=0.415
+ $X2=2.775 $Y2=0.415
r228 29 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.27 $Y=0.415
+ $X2=4.355 $Y2=0.415
r229 29 30 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=4.27 $Y=0.415
+ $X2=3.04 $Y2=0.415
r230 28 31 9.04258 $w=3.71e-07 $l=2.18746e-07 $layer=LI1_cond $X=2.955 $Y=1.605
+ $X2=3.08 $Y2=1.77
r231 28 53 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=2.955 $Y=1.605
+ $X2=2.955 $Y2=0.81
r232 22 76 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.315 $Y=2.305
+ $X2=7.315 $Y2=2.14
r233 22 24 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=7.315 $Y=2.305
+ $X2=7.315 $Y2=2.675
r234 20 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.715 $Y=1.27
+ $X2=6.88 $Y2=1.27
r235 20 21 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=6.715 $Y=1.27
+ $X2=6.355 $Y2=1.27
r236 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.28 $Y=1.195
+ $X2=6.355 $Y2=1.27
r237 17 19 146.207 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=6.28 $Y=1.195
+ $X2=6.28 $Y2=0.74
r238 13 26 70.1453 $w=1.97e-07 $l=3.01247e-07 $layer=POLY_cond $X=4.01 $Y=1.405
+ $X2=3.955 $Y2=1.68
r239 13 15 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.01 $Y=1.405
+ $X2=4.01 $Y2=0.9
r240 12 68 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.495 $Y=1.68
+ $X2=3.33 $Y2=1.68
r241 11 26 9.2281 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=3.825 $Y=1.68
+ $X2=3.955 $Y2=1.68
r242 11 12 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.825 $Y=1.68
+ $X2=3.495 $Y2=1.68
r243 7 34 33.9886 $w=3.28e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.405 $Y=1.935
+ $X2=3.33 $Y2=1.77
r244 7 9 229.339 $w=1.8e-07 $l=5.9e-07 $layer=POLY_cond $X=3.405 $Y=1.935
+ $X2=3.405 $Y2=2.525
r245 2 56 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.935 $X2=2.6 $Y2=2.11
r246 1 52 182 $w=1.7e-07 $l=1.94422e-07 $layer=licon1_NDIFF $count=1 $X=2.535
+ $Y=0.595 $X2=2.675 $Y2=0.725
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_2%A_837_359# 1 2 9 13 17 18 20 21 24 30 32 33
c85 21 0 1.95601e-19 $X=4.445 $Y=1.04
c86 17 0 4.03239e-20 $X=4.36 $Y=1.96
c87 13 0 1.23255e-19 $X=4.4 $Y=0.9
r88 30 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.18 $Y=2.02
+ $X2=6.18 $Y2=1.855
r89 26 32 3.70735 $w=2.5e-07 $l=1.21589e-07 $layer=LI1_cond $X=6.1 $Y=1.13
+ $X2=6.02 $Y2=1.042
r90 26 33 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=6.1 $Y=1.13 $X2=6.1
+ $Y2=1.855
r91 22 32 3.70735 $w=2.5e-07 $l=8.7e-08 $layer=LI1_cond $X=6.02 $Y=0.955
+ $X2=6.02 $Y2=1.042
r92 22 24 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=6.02 $Y=0.955
+ $X2=6.02 $Y2=0.86
r93 20 32 2.76166 $w=1.7e-07 $l=1.65997e-07 $layer=LI1_cond $X=5.855 $Y=1.04
+ $X2=6.02 $Y2=1.042
r94 20 21 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=5.855 $Y=1.04
+ $X2=4.445 $Y2=1.04
r95 18 36 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=4.355 $Y=1.96
+ $X2=4.355 $Y2=2.125
r96 18 35 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=4.355 $Y=1.96
+ $X2=4.355 $Y2=1.795
r97 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.36
+ $Y=1.96 $X2=4.36 $Y2=1.96
r98 15 21 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=4.357 $Y=1.125
+ $X2=4.445 $Y2=1.04
r99 15 17 52.9195 $w=1.73e-07 $l=8.35e-07 $layer=LI1_cond $X=4.357 $Y=1.125
+ $X2=4.357 $Y2=1.96
r100 13 35 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=4.4 $Y=0.9 $X2=4.4
+ $Y2=1.795
r101 9 36 155.484 $w=1.8e-07 $l=4e-07 $layer=POLY_cond $X=4.275 $Y=2.525
+ $X2=4.275 $Y2=2.125
r102 2 30 300 $w=1.7e-07 $l=3.65992e-07 $layer=licon1_PDIFF $count=2 $X=5.995
+ $Y=1.735 $X2=6.18 $Y2=2.02
r103 1 24 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=5.88
+ $Y=0.37 $X2=6.02 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_2%RESET_B 4 6 9 11 12 16 18 21 25 29 33 35 36
+ 37 38 41 43 46 49 50 53 60 64 65
c210 49 0 1.04983e-19 $X=1.12 $Y=1.305
c211 43 0 3.83476e-20 $X=7.92 $Y=2.035
c212 37 0 4.38853e-20 $X=7.775 $Y=2.035
c213 33 0 4.03239e-20 $X=4.88 $Y=1.26
c214 11 0 1.93401e-20 $X=4.715 $Y=0.18
r215 64 67 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.23 $Y=2.11
+ $X2=8.23 $Y2=2.275
r216 64 66 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.23 $Y=2.11
+ $X2=8.23 $Y2=1.945
r217 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.23
+ $Y=2.11 $X2=8.23 $Y2=2.11
r218 58 60 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=4.895 $Y=1.96
+ $X2=5.12 $Y2=1.96
r219 56 58 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.88 $Y=1.96
+ $X2=4.895 $Y2=1.96
r220 53 55 41.3282 $w=4.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.985
+ $X2=1.055 $Y2=2.15
r221 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.12
+ $Y=1.985 $X2=1.12 $Y2=1.985
r222 50 54 27.9879 $w=2.78e-07 $l=6.8e-07 $layer=LI1_cond $X=1.145 $Y=1.305
+ $X2=1.145 $Y2=1.985
r223 49 51 47.2161 $w=4.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.305
+ $X2=1.055 $Y2=1.14
r224 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.12
+ $Y=1.305 $X2=1.12 $Y2=1.305
r225 46 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.035
+ $X2=1.2 $Y2=2.035
r226 44 65 10.0636 $w=3.53e-07 $l=3.1e-07 $layer=LI1_cond $X=7.92 $Y=2.097
+ $X2=8.23 $Y2=2.097
r227 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r228 41 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.12
+ $Y=1.96 $X2=5.12 $Y2=1.96
r229 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=2.035
+ $X2=5.04 $Y2=2.035
r230 38 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=2.035
+ $X2=5.04 $Y2=2.035
r231 37 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r232 37 38 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=5.185 $Y2=2.035
r233 36 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=2.035
+ $X2=1.2 $Y2=2.035
r234 35 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=5.04 $Y2=2.035
r235 35 36 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=1.345 $Y2=2.035
r236 31 33 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.79 $Y=1.26 $X2=4.88
+ $Y2=1.26
r237 29 66 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=8.24 $Y=0.615
+ $X2=8.24 $Y2=1.945
r238 25 67 155.484 $w=1.8e-07 $l=4e-07 $layer=POLY_cond $X=8.235 $Y=2.675
+ $X2=8.235 $Y2=2.275
r239 19 58 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.895 $Y=2.125
+ $X2=4.895 $Y2=1.96
r240 19 21 155.484 $w=1.8e-07 $l=4e-07 $layer=POLY_cond $X=4.895 $Y=2.125
+ $X2=4.895 $Y2=2.525
r241 18 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.88 $Y=1.795
+ $X2=4.88 $Y2=1.96
r242 17 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.88 $Y=1.335
+ $X2=4.88 $Y2=1.26
r243 17 18 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=4.88 $Y=1.335
+ $X2=4.88 $Y2=1.795
r244 14 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.79 $Y=1.185
+ $X2=4.79 $Y2=1.26
r245 14 16 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.79 $Y=1.185
+ $X2=4.79 $Y2=0.9
r246 13 16 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=4.79 $Y=0.255
+ $X2=4.79 $Y2=0.9
r247 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.715 $Y=0.18
+ $X2=4.79 $Y2=0.255
r248 11 12 1917.74 $w=1.5e-07 $l=3.74e-06 $layer=POLY_cond $X=4.715 $Y=0.18
+ $X2=0.975 $Y2=0.18
r249 9 55 270.153 $w=1.8e-07 $l=6.95e-07 $layer=POLY_cond $X=0.945 $Y=2.845
+ $X2=0.945 $Y2=2.15
r250 6 53 7.8587 $w=4.6e-07 $l=6.5e-08 $layer=POLY_cond $X=1.055 $Y=1.92
+ $X2=1.055 $Y2=1.985
r251 5 49 7.8587 $w=4.6e-07 $l=6.5e-08 $layer=POLY_cond $X=1.055 $Y=1.37
+ $X2=1.055 $Y2=1.305
r252 5 6 66.4967 $w=4.6e-07 $l=5.5e-07 $layer=POLY_cond $X=1.055 $Y=1.37
+ $X2=1.055 $Y2=1.92
r253 4 51 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=0.9 $Y=0.6 $X2=0.9
+ $Y2=1.14
r254 1 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.9 $Y=0.255
+ $X2=0.975 $Y2=0.18
r255 1 4 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=0.9 $Y=0.255 $X2=0.9
+ $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_2%A_699_463# 1 2 3 12 16 18 19 21 22 23 25 26
+ 28 33 41 43
c120 41 0 1.23255e-19 $X=4.015 $Y=0.867
c121 26 0 1.21261e-19 $X=4.785 $Y=1.435
r122 39 41 6.41867 $w=3.93e-07 $l=2.2e-07 $layer=LI1_cond $X=3.795 $Y=0.867
+ $X2=4.015 $Y2=0.867
r123 36 37 9.72464 $w=4.83e-07 $l=3.85e-07 $layer=LI1_cond $X=3.63 $Y=2.577
+ $X2=4.015 $Y2=2.577
r124 31 43 4.18896 $w=2.17e-07 $l=9.0802e-08 $layer=LI1_cond $X=4.785 $Y=2.422
+ $X2=4.7 $Y2=2.41
r125 31 33 18.1242 $w=2.03e-07 $l=3.35e-07 $layer=LI1_cond $X=4.785 $Y=2.422
+ $X2=5.12 $Y2=2.422
r126 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.52
+ $Y=1.41 $X2=5.52 $Y2=1.41
r127 26 28 30.2516 $w=2.78e-07 $l=7.35e-07 $layer=LI1_cond $X=4.785 $Y=1.435
+ $X2=5.52 $Y2=1.435
r128 25 43 2.24312 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.7 $Y=2.295
+ $X2=4.7 $Y2=2.41
r129 24 26 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=4.7 $Y=1.575
+ $X2=4.785 $Y2=1.435
r130 24 25 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=4.7 $Y=1.575
+ $X2=4.7 $Y2=2.295
r131 23 37 9.29934 $w=4.83e-07 $l=3.0736e-07 $layer=LI1_cond $X=4.25 $Y=2.41
+ $X2=4.015 $Y2=2.577
r132 22 43 4.18896 $w=2.17e-07 $l=8.5e-08 $layer=LI1_cond $X=4.615 $Y=2.41
+ $X2=4.7 $Y2=2.41
r133 22 23 18.2888 $w=2.28e-07 $l=3.65e-07 $layer=LI1_cond $X=4.615 $Y=2.41
+ $X2=4.25 $Y2=2.41
r134 21 37 6.94006 $w=1.7e-07 $l=2.82e-07 $layer=LI1_cond $X=4.015 $Y=2.295
+ $X2=4.015 $Y2=2.577
r135 20 41 5.70203 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=4.015 $Y=1.065
+ $X2=4.015 $Y2=0.867
r136 20 21 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=4.015 $Y=1.065
+ $X2=4.015 $Y2=2.295
r137 18 29 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.73 $Y=1.41
+ $X2=5.52 $Y2=1.41
r138 18 19 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.73 $Y=1.41
+ $X2=5.73 $Y2=1.245
r139 14 19 34.7346 $w=1.65e-07 $l=4.08228e-07 $layer=POLY_cond $X=5.905 $Y=1.575
+ $X2=5.73 $Y2=1.245
r140 14 16 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=5.905 $Y=1.575
+ $X2=5.905 $Y2=2.235
r141 10 19 34.7346 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=5.805 $Y=1.245
+ $X2=5.73 $Y2=1.245
r142 10 12 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.805 $Y=1.245
+ $X2=5.805 $Y2=0.74
r143 3 33 600 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=4.985
+ $Y=2.315 $X2=5.12 $Y2=2.44
r144 2 36 600 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_PDIFF $count=1 $X=3.495
+ $Y=2.315 $X2=3.63 $Y2=2.61
r145 1 39 182 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.69 $X2=3.795 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_2%A_306_119# 1 2 9 11 13 15 16 17 18 19 20 22
+ 25 27 32 33 34 37 39 42 45 46 49 50 54
c178 50 0 1.04983e-19 $X=1.647 $Y=1.065
c179 49 0 8.96654e-20 $X=2.572 $Y=1.423
c180 33 0 3.77492e-20 $X=7.255 $Y=1.66
c181 11 0 7.88206e-20 $X=2.46 $Y=1.41
r182 58 62 34.8734 $w=3.87e-07 $l=2.8e-07 $layer=POLY_cond $X=2.6 $Y=1.48
+ $X2=2.88 $Y2=1.48
r183 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.6
+ $Y=1.61 $X2=2.6 $Y2=1.61
r184 51 54 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.54 $Y=2.11 $X2=1.7
+ $Y2=2.11
r185 49 57 9.3627 $w=2.55e-07 $l=1.87e-07 $layer=LI1_cond $X=2.572 $Y=1.423
+ $X2=2.572 $Y2=1.61
r186 48 49 12.3379 $w=2.53e-07 $l=2.73e-07 $layer=LI1_cond $X=2.572 $Y=1.15
+ $X2=2.572 $Y2=1.423
r187 47 50 3.15366 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.84 $Y=1.065
+ $X2=1.647 $Y2=1.065
r188 46 48 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=2.445 $Y=1.065
+ $X2=2.572 $Y2=1.15
r189 46 47 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.445 $Y=1.065
+ $X2=1.84 $Y2=1.065
r190 45 51 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=1.945
+ $X2=1.54 $Y2=2.11
r191 44 50 3.37808 $w=2.77e-07 $l=1.43332e-07 $layer=LI1_cond $X=1.54 $Y=1.15
+ $X2=1.647 $Y2=1.065
r192 44 45 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=1.54 $Y=1.15
+ $X2=1.54 $Y2=1.945
r193 40 50 3.37808 $w=2.77e-07 $l=8.5e-08 $layer=LI1_cond $X=1.647 $Y=0.98
+ $X2=1.647 $Y2=1.065
r194 40 42 7.63306 $w=3.83e-07 $l=2.55e-07 $layer=LI1_cond $X=1.647 $Y=0.98
+ $X2=1.647 $Y2=0.725
r195 35 37 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=7.33 $Y=1.585
+ $X2=7.33 $Y2=0.615
r196 33 35 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.255 $Y=1.66
+ $X2=7.33 $Y2=1.585
r197 33 34 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=7.255 $Y=1.66
+ $X2=6.5 $Y2=1.66
r198 30 32 297.363 $w=1.8e-07 $l=7.65e-07 $layer=POLY_cond $X=6.41 $Y=3.075
+ $X2=6.41 $Y2=2.31
r199 29 34 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.41 $Y=1.735
+ $X2=6.5 $Y2=1.66
r200 29 32 223.508 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.41 $Y=1.735
+ $X2=6.41 $Y2=2.31
r201 28 39 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.945 $Y=3.15
+ $X2=3.855 $Y2=3.15
r202 27 30 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.32 $Y=3.15
+ $X2=6.41 $Y2=3.075
r203 27 28 1217.82 $w=1.5e-07 $l=2.375e-06 $layer=POLY_cond $X=6.32 $Y=3.15
+ $X2=3.945 $Y2=3.15
r204 23 39 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.855 $Y=3.075
+ $X2=3.855 $Y2=3.15
r205 23 25 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=3.855 $Y=3.075
+ $X2=3.855 $Y2=2.525
r206 20 22 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.51 $Y=1.185
+ $X2=3.51 $Y2=0.9
r207 19 62 33.8265 $w=3.87e-07 $l=2.73542e-07 $layer=POLY_cond $X=3.04 $Y=1.275
+ $X2=2.88 $Y2=1.48
r208 18 20 27.2212 $w=1.8e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.435 $Y=1.275
+ $X2=3.51 $Y2=1.185
r209 18 19 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.435 $Y=1.275
+ $X2=3.04 $Y2=1.275
r210 16 39 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.765 $Y=3.15
+ $X2=3.855 $Y2=3.15
r211 16 17 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.765 $Y=3.15
+ $X2=2.955 $Y2=3.15
r212 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.88 $Y=3.075
+ $X2=2.955 $Y2=3.15
r213 14 62 25.0561 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=2.88 $Y=1.775
+ $X2=2.88 $Y2=1.48
r214 14 15 666.596 $w=1.5e-07 $l=1.3e-06 $layer=POLY_cond $X=2.88 $Y=1.775
+ $X2=2.88 $Y2=3.075
r215 11 58 17.4367 $w=3.87e-07 $l=1.4e-07 $layer=POLY_cond $X=2.46 $Y=1.48
+ $X2=2.6 $Y2=1.48
r216 11 59 10.5866 $w=3.87e-07 $l=8.5e-08 $layer=POLY_cond $X=2.46 $Y=1.48
+ $X2=2.375 $Y2=1.48
r217 11 13 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.46 $Y=1.41
+ $X2=2.46 $Y2=0.965
r218 7 59 20.6767 $w=1.8e-07 $l=2.95e-07 $layer=POLY_cond $X=2.375 $Y=1.775
+ $X2=2.375 $Y2=1.48
r219 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.375 $Y=1.775
+ $X2=2.375 $Y2=2.495
r220 2 54 600 $w=1.7e-07 $l=2.3103e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=1.935 $X2=1.7 $Y2=2.11
r221 1 42 91 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_NDIFF $count=2 $X=1.53
+ $Y=0.595 $X2=1.675 $Y2=0.725
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_2%A_1525_212# 1 2 9 13 15 17 18 20 26 29 30 31
+ 32 35 37 38 42
c114 38 0 1.33493e-19 $X=7.79 $Y=1.225
c115 35 0 4.37308e-20 $X=9.29 $Y=2.105
c116 20 0 4.77539e-20 $X=8.715 $Y=2.61
c117 13 0 3.83476e-20 $X=7.735 $Y=2.065
r118 38 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.79 $Y=1.225
+ $X2=7.79 $Y2=1.39
r119 38 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.79 $Y=1.225
+ $X2=7.79 $Y2=1.06
r120 37 40 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.79 $Y=1.225 $X2=7.79
+ $Y2=1.305
r121 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.79
+ $Y=1.225 $X2=7.79 $Y2=1.225
r122 34 35 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=9.29 $Y=1.39
+ $X2=9.29 $Y2=2.105
r123 33 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.01 $Y=1.305
+ $X2=8.845 $Y2=1.305
r124 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.205 $Y=1.305
+ $X2=9.29 $Y2=1.39
r125 32 33 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=9.205 $Y=1.305
+ $X2=9.01 $Y2=1.305
r126 30 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.205 $Y=2.19
+ $X2=9.29 $Y2=2.105
r127 30 31 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=9.205 $Y=2.19
+ $X2=8.885 $Y2=2.19
r128 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.8 $Y=2.275
+ $X2=8.885 $Y2=2.19
r129 28 29 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=8.8 $Y=2.275
+ $X2=8.8 $Y2=2.445
r130 24 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.845 $Y=1.22
+ $X2=8.845 $Y2=1.305
r131 24 26 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=8.845 $Y=1.22
+ $X2=8.845 $Y2=0.615
r132 20 29 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.715 $Y=2.61
+ $X2=8.8 $Y2=2.445
r133 20 22 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=8.715 $Y=2.61
+ $X2=8.59 $Y2=2.61
r134 19 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.955 $Y=1.305
+ $X2=7.79 $Y2=1.305
r135 18 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.68 $Y=1.305
+ $X2=8.845 $Y2=1.305
r136 18 19 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=8.68 $Y=1.305
+ $X2=7.955 $Y2=1.305
r137 17 45 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=7.72 $Y=1.975
+ $X2=7.72 $Y2=1.39
r138 13 17 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=7.735 $Y=2.065
+ $X2=7.735 $Y2=1.975
r139 13 15 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=7.735 $Y=2.065
+ $X2=7.735 $Y2=2.675
r140 9 44 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=7.72 $Y=0.615
+ $X2=7.72 $Y2=1.06
r141 2 22 600 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_PDIFF $count=1 $X=8.325
+ $Y=2.465 $X2=8.59 $Y2=2.61
r142 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.705
+ $Y=0.405 $X2=8.845 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_2%A_1271_74# 1 2 9 13 15 16 19 23 25 26 27 29
+ 32 34 35 39 40 41 46 48
c140 39 0 3.77492e-20 $X=7.54 $Y=2.475
c141 16 0 4.77539e-20 $X=9.035 $Y=1.63
c142 13 0 1.34198e-19 $X=8.945 $Y=2.675
r143 52 56 13.0505 $w=2.77e-07 $l=7.5e-08 $layer=POLY_cond $X=8.87 $Y=1.722
+ $X2=8.945 $Y2=1.722
r144 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.87
+ $Y=1.725 $X2=8.87 $Y2=1.725
r145 48 51 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=8.87 $Y=1.645 $X2=8.87
+ $Y2=1.725
r146 44 46 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=6.44 $Y=1.6 $X2=6.6
+ $Y2=1.6
r147 40 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.705 $Y=1.645
+ $X2=8.87 $Y2=1.645
r148 40 41 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=8.705 $Y=1.645
+ $X2=7.625 $Y2=1.645
r149 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.54 $Y=1.73
+ $X2=7.625 $Y2=1.645
r150 38 39 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=7.54 $Y=1.73
+ $X2=7.54 $Y2=2.475
r151 35 37 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=6.685 $Y=2.64
+ $X2=7.09 $Y2=2.64
r152 34 39 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.455 $Y=2.64
+ $X2=7.54 $Y2=2.475
r153 34 37 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=7.455 $Y=2.64
+ $X2=7.09 $Y2=2.64
r154 30 43 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.525 $Y=0.72
+ $X2=6.44 $Y2=0.72
r155 30 32 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=6.525 $Y=0.72
+ $X2=6.95 $Y2=0.72
r156 29 35 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.6 $Y=2.475
+ $X2=6.685 $Y2=2.64
r157 28 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.6 $Y=1.685
+ $X2=6.6 $Y2=1.6
r158 28 29 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=6.6 $Y=1.685
+ $X2=6.6 $Y2=2.475
r159 27 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.44 $Y=1.515
+ $X2=6.44 $Y2=1.6
r160 26 43 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.44 $Y=0.845
+ $X2=6.44 $Y2=0.72
r161 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.44 $Y=0.845
+ $X2=6.44 $Y2=1.515
r162 21 25 18.8402 $w=1.65e-07 $l=9.60469e-08 $layer=POLY_cond $X=9.61 $Y=1.555
+ $X2=9.562 $Y2=1.63
r163 21 23 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=9.61 $Y=1.555
+ $X2=9.61 $Y2=0.74
r164 17 25 18.8402 $w=1.65e-07 $l=8.95824e-08 $layer=POLY_cond $X=9.53 $Y=1.705
+ $X2=9.562 $Y2=1.63
r165 17 19 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=9.53 $Y=1.705
+ $X2=9.53 $Y2=2.465
r166 16 56 25.7246 $w=2.77e-07 $l=1.29399e-07 $layer=POLY_cond $X=9.035 $Y=1.63
+ $X2=8.945 $Y2=1.722
r167 15 25 6.66866 $w=1.5e-07 $l=1.22e-07 $layer=POLY_cond $X=9.44 $Y=1.63
+ $X2=9.562 $Y2=1.63
r168 15 16 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=9.44 $Y=1.63
+ $X2=9.035 $Y2=1.63
r169 11 56 12.8788 $w=1.8e-07 $l=1.68e-07 $layer=POLY_cond $X=8.945 $Y=1.89
+ $X2=8.945 $Y2=1.722
r170 11 13 305.137 $w=1.8e-07 $l=7.85e-07 $layer=POLY_cond $X=8.945 $Y=1.89
+ $X2=8.945 $Y2=2.675
r171 7 52 41.7617 $w=2.77e-07 $l=3.12538e-07 $layer=POLY_cond $X=8.63 $Y=1.555
+ $X2=8.87 $Y2=1.722
r172 7 9 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=8.63 $Y=1.555 $X2=8.63
+ $Y2=0.615
r173 2 37 300 $w=1.7e-07 $l=1.08563e-06 $layer=licon1_PDIFF $count=2 $X=6.5
+ $Y=1.81 $X2=7.09 $Y2=2.64
r174 1 43 182 $w=1.7e-07 $l=3.83732e-07 $layer=licon1_NDIFF $count=1 $X=6.355
+ $Y=0.37 $X2=6.52 $Y2=0.68
r175 1 32 182 $w=1.7e-07 $l=7.33809e-07 $layer=licon1_NDIFF $count=1 $X=6.355
+ $Y=0.37 $X2=6.95 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_2%A_1924_409# 1 2 7 11 15 17 21 25 27 28 31 35
+ 39 44 47
c67 47 0 4.37308e-20 $X=10.09 $Y=1.375
c68 31 0 1.34198e-19 $X=9.755 $Y=2.195
r69 45 47 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=10.09 $Y=1.465
+ $X2=10.09 $Y2=1.375
r70 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.09
+ $Y=1.465 $X2=10.09 $Y2=1.465
r71 42 44 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=9.825 $Y=1.465
+ $X2=10.09 $Y2=1.465
r72 40 42 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=9.79 $Y=1.465
+ $X2=9.825 $Y2=1.465
r73 37 40 2.13598 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=9.79 $Y=1.63
+ $X2=9.79 $Y2=1.465
r74 37 39 17.7299 $w=2.58e-07 $l=4e-07 $layer=LI1_cond $X=9.79 $Y=1.63 $X2=9.79
+ $Y2=2.03
r75 33 42 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.825 $Y=1.3
+ $X2=9.825 $Y2=1.465
r76 33 35 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=9.825 $Y=1.3
+ $X2=9.825 $Y2=0.515
r77 31 39 6.31279 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.755 $Y=2.195
+ $X2=9.755 $Y2=2.03
r78 23 28 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=11.03 $Y=1.3
+ $X2=11.015 $Y2=1.375
r79 23 25 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.03 $Y=1.3
+ $X2=11.03 $Y2=0.74
r80 19 28 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=11.015 $Y=1.45
+ $X2=11.015 $Y2=1.375
r81 19 21 369.274 $w=1.8e-07 $l=9.5e-07 $layer=POLY_cond $X=11.015 $Y=1.45
+ $X2=11.015 $Y2=2.4
r82 18 27 13.2179 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=10.675 $Y=1.375
+ $X2=10.575 $Y2=1.375
r83 17 28 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=10.925 $Y=1.375
+ $X2=11.015 $Y2=1.375
r84 17 18 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=10.925 $Y=1.375
+ $X2=10.675 $Y2=1.375
r85 13 27 10.9219 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=10.6 $Y=1.3
+ $X2=10.575 $Y2=1.375
r86 13 15 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=10.6 $Y=1.3 $X2=10.6
+ $Y2=0.74
r87 9 27 10.9219 $w=1.8e-07 $l=7.98436e-08 $layer=POLY_cond $X=10.565 $Y=1.45
+ $X2=10.575 $Y2=1.375
r88 9 11 369.274 $w=1.8e-07 $l=9.5e-07 $layer=POLY_cond $X=10.565 $Y=1.45
+ $X2=10.565 $Y2=2.4
r89 8 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.255 $Y=1.375
+ $X2=10.09 $Y2=1.375
r90 7 27 13.2179 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=10.475 $Y=1.375
+ $X2=10.575 $Y2=1.375
r91 7 8 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=10.475 $Y=1.375
+ $X2=10.255 $Y2=1.375
r92 2 31 300 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=2 $X=9.62
+ $Y=2.045 $X2=9.755 $Y2=2.195
r93 1 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.685
+ $Y=0.37 $X2=9.825 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_2%VPWR 1 2 3 4 5 6 7 8 9 28 30 34 38 42 44 48
+ 54 58 62 66 68 73 74 75 77 82 87 95 107 111 120 123 126 129 132 135 139
r152 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r153 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r154 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r155 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r156 127 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r157 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r158 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r159 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r160 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r161 115 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r162 115 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=10.32 $Y2=3.33
r163 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r164 112 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.48 $Y=3.33
+ $X2=10.315 $Y2=3.33
r165 112 114 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=10.48 $Y=3.33
+ $X2=10.8 $Y2=3.33
r166 111 138 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=11.155 $Y=3.33
+ $X2=11.337 $Y2=3.33
r167 111 114 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=11.155 $Y=3.33
+ $X2=10.8 $Y2=3.33
r168 110 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r169 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r170 107 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.15 $Y=3.33
+ $X2=10.315 $Y2=3.33
r171 107 109 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.15 $Y=3.33
+ $X2=9.84 $Y2=3.33
r172 106 110 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.84 $Y2=3.33
r173 106 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=7.92 $Y2=3.33
r174 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r175 103 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.125 $Y=3.33
+ $X2=7.96 $Y2=3.33
r176 103 105 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=8.125 $Y=3.33
+ $X2=8.88 $Y2=3.33
r177 102 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r178 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r179 99 102 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=7.44 $Y2=3.33
r180 98 101 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6 $Y=3.33
+ $X2=7.44 $Y2=3.33
r181 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r182 96 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=5.68 $Y2=3.33
r183 96 98 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.845 $Y=3.33
+ $X2=6 $Y2=3.33
r184 95 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.795 $Y=3.33
+ $X2=7.96 $Y2=3.33
r185 95 101 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.795 $Y=3.33
+ $X2=7.44 $Y2=3.33
r186 94 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r187 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r188 91 94 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r189 91 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r190 90 93 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r191 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r192 88 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=2.15 $Y2=3.33
r193 88 90 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.315 $Y=3.33
+ $X2=2.64 $Y2=3.33
r194 87 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.42 $Y=3.33
+ $X2=4.585 $Y2=3.33
r195 87 93 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.42 $Y=3.33
+ $X2=4.08 $Y2=3.33
r196 86 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r197 86 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r198 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r199 83 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.17 $Y2=3.33
r200 83 85 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.68 $Y2=3.33
r201 82 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=2.15 $Y2=3.33
r202 82 85 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.985 $Y=3.33
+ $X2=1.68 $Y2=3.33
r203 81 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r204 81 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r205 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r206 78 117 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.217 $Y2=3.33
r207 78 80 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.72 $Y2=3.33
r208 77 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.17 $Y2=3.33
r209 77 80 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.72 $Y2=3.33
r210 75 99 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=6 $Y2=3.33
r211 75 130 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=3.33
+ $X2=5.52 $Y2=3.33
r212 73 105 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=9.09 $Y=3.33
+ $X2=8.88 $Y2=3.33
r213 73 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.09 $Y=3.33
+ $X2=9.255 $Y2=3.33
r214 72 109 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=9.42 $Y=3.33
+ $X2=9.84 $Y2=3.33
r215 72 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.42 $Y=3.33
+ $X2=9.255 $Y2=3.33
r216 68 71 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=11.28 $Y=1.985
+ $X2=11.28 $Y2=2.815
r217 66 138 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=11.28 $Y=3.245
+ $X2=11.337 $Y2=3.33
r218 66 71 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.28 $Y=3.245
+ $X2=11.28 $Y2=2.815
r219 62 65 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=10.315 $Y=1.985
+ $X2=10.315 $Y2=2.815
r220 60 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.315 $Y=3.245
+ $X2=10.315 $Y2=3.33
r221 60 65 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.315 $Y=3.245
+ $X2=10.315 $Y2=2.815
r222 56 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.255 $Y=3.245
+ $X2=9.255 $Y2=3.33
r223 56 58 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=9.255 $Y=3.245
+ $X2=9.255 $Y2=2.675
r224 52 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.96 $Y=3.245
+ $X2=7.96 $Y2=3.33
r225 52 54 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=7.96 $Y=3.245
+ $X2=7.96 $Y2=2.675
r226 48 51 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.68 $Y=1.91
+ $X2=5.68 $Y2=2.59
r227 46 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.68 $Y=3.245
+ $X2=5.68 $Y2=3.33
r228 46 51 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=5.68 $Y=3.245
+ $X2=5.68 $Y2=2.59
r229 45 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.75 $Y=3.33
+ $X2=4.585 $Y2=3.33
r230 44 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.515 $Y=3.33
+ $X2=5.68 $Y2=3.33
r231 44 45 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=5.515 $Y=3.33
+ $X2=4.75 $Y2=3.33
r232 40 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.585 $Y=3.245
+ $X2=4.585 $Y2=3.33
r233 40 42 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.585 $Y=3.245
+ $X2=4.585 $Y2=2.78
r234 36 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=3.245
+ $X2=2.15 $Y2=3.33
r235 36 38 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.15 $Y=3.245
+ $X2=2.15 $Y2=2.88
r236 32 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=3.33
r237 32 34 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=2.88
r238 28 117 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.217 $Y2=3.33
r239 28 30 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=0.27 $Y=3.245 $X2=0.27
+ $Y2=2.845
r240 9 71 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=11.105
+ $Y=1.84 $X2=11.24 $Y2=2.815
r241 9 68 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=11.105
+ $Y=1.84 $X2=11.24 $Y2=1.985
r242 8 65 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=10.17
+ $Y=1.84 $X2=10.315 $Y2=2.815
r243 8 62 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.17
+ $Y=1.84 $X2=10.315 $Y2=1.985
r244 7 58 600 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_PDIFF $count=1 $X=9.035
+ $Y=2.465 $X2=9.255 $Y2=2.675
r245 6 54 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=7.825
+ $Y=2.465 $X2=7.96 $Y2=2.675
r246 5 51 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.535
+ $Y=1.735 $X2=5.68 $Y2=2.59
r247 5 48 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.535
+ $Y=1.735 $X2=5.68 $Y2=1.91
r248 4 42 600 $w=1.7e-07 $l=5.6438e-07 $layer=licon1_PDIFF $count=1 $X=4.365
+ $Y=2.315 $X2=4.585 $Y2=2.78
r249 3 38 600 $w=1.7e-07 $l=1.01025e-06 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.935 $X2=2.15 $Y2=2.88
r250 2 34 600 $w=1.7e-07 $l=3.05123e-07 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=2.635 $X2=1.17 $Y2=2.88
r251 1 30 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.635 $X2=0.27 $Y2=2.845
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_2%A_30_78# 1 2 3 4 13 17 20 24 27 29 30 32 34
+ 38 41 42 46
c120 41 0 6.1174e-20 $X=3.015 $Y=2.585
c121 17 0 1.98761e-19 $X=0.72 $Y=2.845
r122 40 42 4.73325 $w=2.78e-07 $l=1.15e-07 $layer=LI1_cond $X=3.175 $Y=2.585
+ $X2=3.29 $Y2=2.585
r123 40 41 8.05131 $w=2.78e-07 $l=1.6e-07 $layer=LI1_cond $X=3.175 $Y=2.585
+ $X2=3.015 $Y2=2.585
r124 34 36 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.295 $Y=0.6
+ $X2=0.295 $Y2=0.745
r125 31 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.675 $Y=1.405
+ $X2=3.675 $Y2=1.32
r126 31 32 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.675 $Y=1.405
+ $X2=3.675 $Y2=2.105
r127 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.59 $Y=2.19
+ $X2=3.675 $Y2=2.105
r128 29 30 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.59 $Y=2.19
+ $X2=3.375 $Y2=2.19
r129 25 46 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.335 $Y=1.32
+ $X2=3.675 $Y2=1.32
r130 25 27 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.335 $Y=1.235
+ $X2=3.335 $Y2=0.9
r131 24 42 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.29 $Y=2.445
+ $X2=3.29 $Y2=2.585
r132 23 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.29 $Y=2.275
+ $X2=3.375 $Y2=2.19
r133 23 24 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.29 $Y=2.275
+ $X2=3.29 $Y2=2.445
r134 22 38 1.44141 $w=1.8e-07 $l=2.07364e-07 $layer=LI1_cond $X=0.835 $Y=2.535
+ $X2=0.635 $Y2=2.52
r135 22 41 134.323 $w=1.78e-07 $l=2.18e-06 $layer=LI1_cond $X=0.835 $Y=2.535
+ $X2=3.015 $Y2=2.535
r136 20 38 5.04926 $w=1.85e-07 $l=1.47817e-07 $layer=LI1_cond $X=0.75 $Y=2.445
+ $X2=0.635 $Y2=2.52
r137 19 20 105.364 $w=1.68e-07 $l=1.615e-06 $layer=LI1_cond $X=0.75 $Y=0.83
+ $X2=0.75 $Y2=2.445
r138 15 38 5.04926 $w=1.85e-07 $l=1.46714e-07 $layer=LI1_cond $X=0.735 $Y=2.625
+ $X2=0.635 $Y2=2.52
r139 15 17 12.2 $w=1.98e-07 $l=2.2e-07 $layer=LI1_cond $X=0.735 $Y=2.625
+ $X2=0.735 $Y2=2.845
r140 14 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.46 $Y=0.745
+ $X2=0.295 $Y2=0.745
r141 13 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.665 $Y=0.745
+ $X2=0.75 $Y2=0.83
r142 13 14 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.665 $Y=0.745
+ $X2=0.46 $Y2=0.745
r143 4 40 600 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=2.315 $X2=3.175 $Y2=2.535
r144 3 17 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.635 $X2=0.72 $Y2=2.845
r145 2 27 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.15
+ $Y=0.69 $X2=3.295 $Y2=0.9
r146 1 34 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.39 $X2=0.295 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_2%Q 1 2 7 8 9 10 11 12 13
r20 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.815 $Y=2.405
+ $X2=10.815 $Y2=2.775
r21 11 12 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=10.815 $Y=1.985
+ $X2=10.815 $Y2=2.405
r22 10 11 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=10.815 $Y=1.665
+ $X2=10.815 $Y2=1.985
r23 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.815 $Y=1.295
+ $X2=10.815 $Y2=1.665
r24 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.815 $Y=0.925
+ $X2=10.815 $Y2=1.295
r25 7 8 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=10.815 $Y=0.515
+ $X2=10.815 $Y2=0.925
r26 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.655
+ $Y=1.84 $X2=10.79 $Y2=2.815
r27 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.655
+ $Y=1.84 $X2=10.79 $Y2=1.985
r28 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.675
+ $Y=0.37 $X2=10.815 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_2%VGND 1 2 3 4 5 6 7 24 28 32 36 40 42 44 47
+ 48 49 55 59 67 75 80 85 91 101 104 107 111
r118 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r119 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r120 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r121 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r122 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r123 89 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r124 89 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r125 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r126 86 107 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.47 $Y=0
+ $X2=10.345 $Y2=0
r127 86 88 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=10.47 $Y=0 $X2=10.8
+ $Y2=0
r128 85 110 4.01803 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=11.16 $Y=0
+ $X2=11.34 $Y2=0
r129 85 88 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=11.16 $Y=0 $X2=10.8
+ $Y2=0
r130 84 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r131 84 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=9.36 $Y2=0
r132 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r133 81 104 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.48 $Y=0
+ $X2=9.355 $Y2=0
r134 81 83 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=9.48 $Y=0 $X2=9.84
+ $Y2=0
r135 80 107 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.22 $Y=0
+ $X2=10.345 $Y2=0
r136 80 83 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=10.22 $Y=0 $X2=9.84
+ $Y2=0
r137 79 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r138 79 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=7.92 $Y2=0
r139 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r140 76 101 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=8.19 $Y=0 $X2=7.98
+ $Y2=0
r141 76 78 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.19 $Y=0 $X2=8.88
+ $Y2=0
r142 75 104 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.23 $Y=0
+ $X2=9.355 $Y2=0
r143 75 78 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=9.23 $Y=0 $X2=8.88
+ $Y2=0
r144 74 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r145 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r146 71 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r147 70 73 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=7.44
+ $Y2=0
r148 70 71 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r149 68 70 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.345 $Y=0
+ $X2=5.52 $Y2=0
r150 67 101 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=7.77 $Y=0 $X2=7.98
+ $Y2=0
r151 67 73 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.77 $Y=0 $X2=7.44
+ $Y2=0
r152 66 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r153 65 66 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r154 63 66 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.56 $Y2=0
r155 63 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r156 62 65 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r157 62 63 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r158 60 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.175
+ $Y2=0
r159 60 62 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.64
+ $Y2=0
r160 59 98 7.59257 $w=4.23e-07 $l=2.8e-07 $layer=LI1_cond $X=5.132 $Y=0
+ $X2=5.132 $Y2=0.28
r161 59 68 6.14847 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=5.132 $Y=0
+ $X2=5.345 $Y2=0
r162 59 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r163 59 65 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.92 $Y=0 $X2=4.56
+ $Y2=0
r164 58 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r165 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r166 55 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=2.175
+ $Y2=0
r167 55 57 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=1.68
+ $Y2=0
r168 53 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r169 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r170 49 74 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=7.44 $Y2=0
r171 49 71 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.76 $Y=0
+ $X2=5.52 $Y2=0
r172 47 52 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=0.72
+ $Y2=0
r173 47 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=1.155
+ $Y2=0
r174 46 57 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.68
+ $Y2=0
r175 46 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.155
+ $Y2=0
r176 42 110 3.12513 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=11.285 $Y=0.085
+ $X2=11.34 $Y2=0
r177 42 44 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.285 $Y=0.085
+ $X2=11.285 $Y2=0.515
r178 38 107 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.345 $Y=0.085
+ $X2=10.345 $Y2=0
r179 38 40 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.345 $Y=0.085
+ $X2=10.345 $Y2=0.515
r180 34 104 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.355 $Y=0.085
+ $X2=9.355 $Y2=0
r181 34 36 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.355 $Y=0.085
+ $X2=9.355 $Y2=0.515
r182 30 101 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=7.98 $Y=0.085
+ $X2=7.98 $Y2=0
r183 30 32 12.7592 $w=4.18e-07 $l=4.65e-07 $layer=LI1_cond $X=7.98 $Y=0.085
+ $X2=7.98 $Y2=0.55
r184 26 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.175 $Y=0.085
+ $X2=2.175 $Y2=0
r185 26 28 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=2.175 $Y=0.085
+ $X2=2.175 $Y2=0.725
r186 22 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0
r187 22 24 23.5098 $w=2.48e-07 $l=5.1e-07 $layer=LI1_cond $X=1.155 $Y=0.085
+ $X2=1.155 $Y2=0.595
r188 7 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.105
+ $Y=0.37 $X2=11.245 $Y2=0.515
r189 6 40 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=10.24
+ $Y=0.37 $X2=10.385 $Y2=0.515
r190 5 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.255
+ $Y=0.37 $X2=9.395 $Y2=0.515
r191 4 32 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=7.795
+ $Y=0.405 $X2=7.98 $Y2=0.55
r192 3 98 182 $w=1.7e-07 $l=5.2607e-07 $layer=licon1_NDIFF $count=1 $X=4.865
+ $Y=0.69 $X2=5.13 $Y2=0.28
r193 2 28 182 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_NDIFF $count=1 $X=1.965
+ $Y=0.595 $X2=2.175 $Y2=0.725
r194 1 24 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=0.975
+ $Y=0.39 $X2=1.115 $Y2=0.595
.ends


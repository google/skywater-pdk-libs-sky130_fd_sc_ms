* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 VGND A2 a_245_94# VNB nlowvt w=640000u l=150000u
+  ad=4.931e+11p pd=4.19e+06u as=4.032e+11p ps=3.82e+06u
M1001 a_245_94# B2 a_456_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.576e+11p ps=3.99e+06u
M1002 a_83_264# A2 a_267_392# VPB pshort w=1e+06u l=180000u
+  ad=6.7e+11p pd=5.34e+06u as=2.4e+11p ps=2.48e+06u
M1003 a_245_94# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND a_83_264# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1005 VPWR B1 a_465_392# VPB pshort w=1e+06u l=180000u
+  ad=1.42e+12p pd=7.02e+06u as=3.9e+11p ps=2.78e+06u
M1006 a_83_264# C1 a_456_74# VNB nlowvt w=640000u l=150000u
+  ad=2.944e+11p pd=2.2e+06u as=0p ps=0u
M1007 VPWR a_83_264# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1008 a_456_74# B1 a_245_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_83_264# C1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_267_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_465_392# B2 a_83_264# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and3_1 A B C VGND VNB VPB VPWR X
M1000 X a_27_398# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=1.00785e+12p ps=6.04e+06u
M1001 a_121_136# A a_27_398# VNB nlowvt w=640000u l=150000u
+  ad=2.624e+11p pd=2.1e+06u as=1.824e+11p ps=1.85e+06u
M1002 a_233_136# B a_121_136# VNB nlowvt w=640000u l=150000u
+  ad=2.22e+11p pd=2.09e+06u as=0p ps=0u
M1003 a_27_398# B VPWR VPB pshort w=840000u l=180000u
+  ad=4.62e+11p pd=4.46e+06u as=0p ps=0u
M1004 VGND C a_233_136# VNB nlowvt w=640000u l=150000u
+  ad=3.107e+11p pd=2.34e+06u as=0p ps=0u
M1005 VPWR C a_27_398# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A a_27_398# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_27_398# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
.ends

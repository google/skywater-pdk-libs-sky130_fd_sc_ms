* File: sky130_fd_sc_ms__dfrtp_4.spice
* Created: Wed Sep  2 12:03:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dfrtp_4.pex.spice"
.subckt sky130_fd_sc_ms__dfrtp_4  VNB VPB D CLK RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* CLK	CLK
* D	D
* VPB	VPB
* VNB	VNB
MM1017 A_124_78# N_D_M1017_g N_A_37_78#_M1017_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_RESET_B_M1005_g A_124_78# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0504 PD=1.37 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_CLK_M1001_g N_A_303_395#_M1001_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.13745 AS=0.245475 PD=1.115 PS=2.15 NRD=7.296 NRS=7.296 M=1
+ R=4.93333 SA=75000.3 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1002 N_A_497_395#_M1002_d N_A_303_395#_M1002_g N_VGND_M1001_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2262 AS=0.13745 PD=2.14 PS=1.115 NRD=4.044 NRS=7.296 M=1
+ R=4.93333 SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_702_463#_M1000_d N_A_303_395#_M1000_g N_A_37_78#_M1000_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1113 PD=0.77 PS=1.37 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.6 A=0.063 P=1.14 MULT=1
MM1036 A_812_138# N_A_497_395#_M1036_g N_A_702_463#_M1000_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75004.1 A=0.063 P=1.14 MULT=1
MM1024 A_890_138# N_A_834_355#_M1024_g A_812_138# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75003.7 A=0.063 P=1.14 MULT=1
MM1033 N_VGND_M1033_d N_RESET_B_M1033_g A_890_138# VNB NLOWVT L=0.15 W=0.42
+ AD=0.221767 AS=0.0504 PD=1.26 PS=0.66 NRD=135.144 NRS=18.564 M=1 R=2.8
+ SA=75001.5 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1011 N_A_834_355#_M1011_d N_A_702_463#_M1011_g N_VGND_M1033_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.47175 AS=0.390733 PD=2.015 PS=2.22 NRD=0 NRS=76.704 M=1
+ R=4.93333 SA=75001.6 SB=75002.9 A=0.111 P=1.78 MULT=1
MM1004 N_A_1353_392#_M1004_d N_A_497_395#_M1004_g N_A_834_355#_M1011_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.292172 AS=0.47175 PD=2.09241 PS=2.015 NRD=0
+ NRS=11.34 M=1 R=4.93333 SA=75003 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1037 A_1647_81# N_A_303_395#_M1037_g N_A_1353_392#_M1004_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.165828 PD=0.66 PS=1.18759 NRD=18.564 NRS=49.992 M=1
+ R=2.8 SA=75003.7 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_A_1678_395#_M1022_g A_1647_81# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0756 AS=0.0504 PD=0.78 PS=0.66 NRD=7.14 NRS=18.564 M=1 R=2.8 SA=75004.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1030 A_1827_81# N_RESET_B_M1030_g N_VGND_M1022_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0756 PD=0.66 PS=0.78 NRD=18.564 NRS=15.708 M=1 R=2.8 SA=75004.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1031 N_A_1678_395#_M1031_d N_A_1353_392#_M1031_g A_1827_81# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75005
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 N_A_2013_409#_M1018_d N_A_1353_392#_M1018_g N_VGND_M1018_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.2627 PD=2.05 PS=2.19 NRD=0 NRS=11.34 M=1
+ R=4.93333 SA=75000.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A_2013_409#_M1003_g N_Q_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.13875 PD=2.05 PS=1.115 NRD=0 NRS=7.296 M=1 R=4.93333 SA=75000.2
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1023 N_VGND_M1023_d N_A_2013_409#_M1023_g N_Q_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.13875 PD=1.09 PS=1.115 NRD=0 NRS=8.1 M=1 R=4.93333 SA=75000.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1032 N_VGND_M1023_d N_A_2013_409#_M1032_g N_Q_M1032_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1038 N_VGND_M1038_d N_A_2013_409#_M1038_g N_Q_M1032_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2035 AS=0.1036 PD=2.03 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1034 N_A_37_78#_M1034_d N_D_M1034_g N_VPWR_M1034_s VPB PSHORT L=0.18 W=0.42
+ AD=0.0567 AS=0.1155 PD=0.69 PS=1.39 NRD=0 NRS=0 M=1 R=2.33333 SA=90000.2
+ SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1035 N_VPWR_M1035_d N_RESET_B_M1035_g N_A_37_78#_M1034_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1134 AS=0.0567 PD=1.38 PS=0.69 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1010_d N_CLK_M1010_g N_A_303_395#_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.332375 PD=1.39 PS=2.92 NRD=0 NRS=13.1793 M=1 R=6.22222
+ SA=90000.2 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1013 N_A_497_395#_M1013_d N_A_303_395#_M1013_g N_VPWR_M1010_d VPB PSHORT
+ L=0.18 W=1.12 AD=0.3024 AS=0.1512 PD=2.78 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.7 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1014 N_A_702_463#_M1014_d N_A_497_395#_M1014_g N_A_37_78#_M1014_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0567 AS=0.1155 PD=0.69 PS=1.39 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90001.6 A=0.0756 P=1.2 MULT=1
MM1019 A_792_463# N_A_303_395#_M1019_g N_A_702_463#_M1014_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0441 AS=0.0567 PD=0.63 PS=0.69 NRD=23.443 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1006 N_VPWR_M1006_d N_A_834_355#_M1006_g A_792_463# VPB PSHORT L=0.18 W=0.42
+ AD=0.1232 AS=0.0441 PD=1.085 PS=0.63 NRD=111.778 NRS=23.443 M=1 R=2.33333
+ SA=90001 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1016 N_A_702_463#_M1016_d N_RESET_B_M1016_g N_VPWR_M1006_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1155 AS=0.1232 PD=1.39 PS=1.085 NRD=0 NRS=111.778 M=1 R=2.33333
+ SA=90001.6 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1015 N_A_834_355#_M1015_d N_A_702_463#_M1015_g N_VPWR_M1015_s VPB PSHORT
+ L=0.18 W=1 AD=0.135 AS=0.2695 PD=1.27 PS=2.65 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90003.2 A=0.18 P=2.36 MULT=1
MM1020 N_A_1353_392#_M1020_d N_A_303_395#_M1020_g N_A_834_355#_M1015_d VPB
+ PSHORT L=0.18 W=1 AD=0.458521 AS=0.135 PD=3.10563 PS=1.27 NRD=66.98 NRS=0 M=1
+ R=5.55556 SA=90000.6 SB=90002.8 A=0.18 P=2.36 MULT=1
MM1007 A_1630_493# N_A_497_395#_M1007_g N_A_1353_392#_M1020_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.192579 PD=0.66 PS=1.30437 NRD=30.4759 NRS=0 M=1
+ R=2.33333 SA=90002 SB=90005 A=0.0756 P=1.2 MULT=1
MM1012 N_VPWR_M1012_d N_A_1678_395#_M1012_g A_1630_493# VPB PSHORT L=0.18 W=0.42
+ AD=0.0756 AS=0.0504 PD=0.78 PS=0.66 NRD=16.4101 NRS=30.4759 M=1 R=2.33333
+ SA=90002.4 SB=90004.6 A=0.0756 P=1.2 MULT=1
MM1026 N_A_1678_395#_M1026_d N_RESET_B_M1026_g N_VPWR_M1012_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0567 AS=0.0756 PD=0.69 PS=0.78 NRD=0 NRS=21.0987 M=1 R=2.33333
+ SA=90003 SB=90004 A=0.0756 P=1.2 MULT=1
MM1027 N_VPWR_M1027_d N_A_1353_392#_M1027_g N_A_1678_395#_M1026_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.0805 AS=0.0567 PD=0.776667 PS=0.69 NRD=16.4101 NRS=0 M=1
+ R=2.33333 SA=90003.4 SB=90003.6 A=0.0756 P=1.2 MULT=1
MM1008 N_VPWR_M1027_d N_A_1353_392#_M1008_g N_A_2013_409#_M1008_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.161 AS=0.1134 PD=1.55333 PS=1.11 NRD=2.3443 NRS=0 M=1
+ R=4.66667 SA=90002.1 SB=90003.1 A=0.1512 P=2.04 MULT=1
MM1025 N_VPWR_M1025_d N_A_1353_392#_M1025_g N_A_2013_409#_M1008_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.147 AS=0.1134 PD=1.23857 PS=1.11 NRD=10.5395 NRS=0 M=1
+ R=4.66667 SA=90002.5 SB=90002.6 A=0.1512 P=2.04 MULT=1
MM1009 N_Q_M1009_d N_A_2013_409#_M1009_g N_VPWR_M1025_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1764 AS=0.196 PD=1.435 PS=1.65143 NRD=7.0329 NRS=0 M=1 R=6.22222
+ SA=90002.3 SB=90002.1 A=0.2016 P=2.6 MULT=1
MM1021 N_Q_M1009_d N_A_2013_409#_M1021_g N_VPWR_M1021_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1764 AS=0.4172 PD=1.435 PS=1.865 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.8
+ SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1028 N_Q_M1028_d N_A_2013_409#_M1028_g N_VPWR_M1021_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.4172 PD=1.39 PS=1.865 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.7
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1029 N_Q_M1028_d N_A_2013_409#_M1029_g N_VPWR_M1029_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90004.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX39_noxref VNB VPB NWDIODE A=25.5078 P=31.6
c_1942 A_1630_493# 0 9.99956e-20 $X=8.15 $Y=2.465
*
.include "sky130_fd_sc_ms__dfrtp_4.pxi.spice"
*
.ends
*
*

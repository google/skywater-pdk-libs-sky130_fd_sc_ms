* File: sky130_fd_sc_ms__a21boi_2.pex.spice
* Created: Wed Sep  2 11:51:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A21BOI_2%B1_N 3 7 9 10 11
c33 11 0 1.32054e-19 $X=0.24 $Y=1.665
r34 11 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.31
+ $Y=1.615 $X2=0.31 $Y2=1.615
r35 9 14 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=0.495 $Y=1.615
+ $X2=0.31 $Y2=1.615
r36 9 10 3.90195 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=0.495 $Y=1.615
+ $X2=0.61 $Y2=1.615
r37 5 10 34.7346 $w=1.65e-07 $l=1.83916e-07 $layer=POLY_cond $X=0.65 $Y=1.45
+ $X2=0.61 $Y2=1.615
r38 5 7 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.65 $Y=1.45 $X2=0.65
+ $Y2=0.79
r39 1 10 34.7346 $w=1.65e-07 $l=1.77059e-07 $layer=POLY_cond $X=0.585 $Y=1.78
+ $X2=0.61 $Y2=1.615
r40 1 3 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=0.585 $Y=1.78
+ $X2=0.585 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A21BOI_2%A_62_94# 1 2 9 11 13 16 18 19 20 22 25 27
+ 28 31 33 35 37
c80 37 0 1.97879e-19 $X=0.81 $Y=1.94
c81 20 0 3.38845e-19 $X=2.005 $Y=1.765
c82 19 0 1.32054e-19 $X=1.645 $Y=1.69
r83 44 45 1.98082 $w=3.65e-07 $l=1.5e-08 $layer=POLY_cond $X=1.555 $Y=1.542
+ $X2=1.57 $Y2=1.542
r84 41 44 42.9178 $w=3.65e-07 $l=3.25e-07 $layer=POLY_cond $X=1.23 $Y=1.542
+ $X2=1.555 $Y2=1.542
r85 41 42 11.8849 $w=3.65e-07 $l=9e-08 $layer=POLY_cond $X=1.23 $Y=1.542
+ $X2=1.14 $Y2=1.542
r86 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.23
+ $Y=1.485 $X2=1.23 $Y2=1.485
r87 35 40 9.27913 $w=4.26e-07 $l=2.80624e-07 $layer=LI1_cond $X=0.89 $Y=1.65
+ $X2=1.1 $Y2=1.485
r88 35 37 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.89 $Y=1.65
+ $X2=0.89 $Y2=1.94
r89 31 37 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.81 $Y=2.105
+ $X2=0.81 $Y2=1.94
r90 31 33 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.81 $Y=2.105
+ $X2=0.81 $Y2=2.815
r91 27 40 8.30516 $w=4.26e-07 $l=4.15421e-07 $layer=LI1_cond $X=0.805 $Y=1.195
+ $X2=1.1 $Y2=1.485
r92 27 28 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.805 $Y=1.195
+ $X2=0.52 $Y2=1.195
r93 23 28 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.395 $Y=1.11
+ $X2=0.52 $Y2=1.195
r94 23 25 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.395 $Y=1.11
+ $X2=0.395 $Y2=0.615
r95 20 22 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=2.005 $Y=1.765
+ $X2=2.005 $Y2=2.4
r96 19 45 27.0958 $w=3.65e-07 $l=1.8167e-07 $layer=POLY_cond $X=1.645 $Y=1.69
+ $X2=1.57 $Y2=1.542
r97 18 20 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.915 $Y=1.69
+ $X2=2.005 $Y2=1.765
r98 18 19 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.915 $Y=1.69
+ $X2=1.645 $Y2=1.69
r99 14 45 23.6381 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1.57 $Y=1.32
+ $X2=1.57 $Y2=1.542
r100 14 16 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.57 $Y=1.32
+ $X2=1.57 $Y2=0.74
r101 11 44 19.2931 $w=1.8e-07 $l=2.23e-07 $layer=POLY_cond $X=1.555 $Y=1.765
+ $X2=1.555 $Y2=1.542
r102 11 13 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=1.555 $Y=1.765
+ $X2=1.555 $Y2=2.4
r103 7 42 23.6381 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=1.14 $Y=1.32
+ $X2=1.14 $Y2=1.542
r104 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.14 $Y=1.32 $X2=1.14
+ $Y2=0.74
r105 2 33 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.675
+ $Y=1.96 $X2=0.81 $Y2=2.815
r106 2 31 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.675
+ $Y=1.96 $X2=0.81 $Y2=2.105
r107 1 25 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.31
+ $Y=0.47 $X2=0.435 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__A21BOI_2%A1 3 7 11 15 17 23 24
c58 15 0 2.70769e-20 $X=2.95 $Y=0.74
r59 24 25 6.75701 $w=3.21e-07 $l=4.5e-08 $layer=POLY_cond $X=2.905 $Y=1.485
+ $X2=2.95 $Y2=1.485
r60 22 24 38.2897 $w=3.21e-07 $l=2.55e-07 $layer=POLY_cond $X=2.65 $Y=1.485
+ $X2=2.905 $Y2=1.485
r61 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.65
+ $Y=1.485 $X2=2.65 $Y2=1.485
r62 20 22 19.5202 $w=3.21e-07 $l=1.3e-07 $layer=POLY_cond $X=2.52 $Y=1.485
+ $X2=2.65 $Y2=1.485
r63 19 20 9.76012 $w=3.21e-07 $l=6.5e-08 $layer=POLY_cond $X=2.455 $Y=1.485
+ $X2=2.52 $Y2=1.485
r64 17 23 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=2.65 $Y=1.665
+ $X2=2.65 $Y2=1.485
r65 13 25 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.32
+ $X2=2.95 $Y2=1.485
r66 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.95 $Y=1.32
+ $X2=2.95 $Y2=0.74
r67 9 24 16.2883 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.905 $Y=1.65
+ $X2=2.905 $Y2=1.485
r68 9 11 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=2.905 $Y=1.65
+ $X2=2.905 $Y2=2.4
r69 5 20 20.5661 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.52 $Y=1.32
+ $X2=2.52 $Y2=1.485
r70 5 7 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.52 $Y=1.32 $X2=2.52
+ $Y2=0.74
r71 1 19 16.2883 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.455 $Y=1.65
+ $X2=2.455 $Y2=1.485
r72 1 3 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=2.455 $Y=1.65
+ $X2=2.455 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A21BOI_2%A2 3 5 7 8 10 13 15 24
c44 5 0 1.6164e-19 $X=3.38 $Y=1.22
r45 23 24 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.81 $Y=1.385
+ $X2=3.825 $Y2=1.385
r46 21 23 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=3.43 $Y=1.385
+ $X2=3.81 $Y2=1.385
r47 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.43
+ $Y=1.385 $X2=3.43 $Y2=1.385
r48 19 21 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=3.38 $Y=1.385 $X2=3.43
+ $Y2=1.385
r49 17 19 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=3.355 $Y=1.385
+ $X2=3.38 $Y2=1.385
r50 15 22 5.92571 $w=3.5e-07 $l=1.7e-07 $layer=LI1_cond $X=3.6 $Y=1.365 $X2=3.43
+ $Y2=1.365
r51 11 24 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.825 $Y=1.55
+ $X2=3.825 $Y2=1.385
r52 11 13 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.825 $Y=1.55
+ $X2=3.825 $Y2=2.4
r53 8 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.81 $Y=1.22
+ $X2=3.81 $Y2=1.385
r54 8 10 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.81 $Y=1.22 $X2=3.81
+ $Y2=0.74
r55 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.38 $Y=1.22
+ $X2=3.38 $Y2=1.385
r56 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.38 $Y=1.22 $X2=3.38
+ $Y2=0.74
r57 1 17 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.355 $Y=1.55
+ $X2=3.355 $Y2=1.385
r58 1 3 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.355 $Y=1.55
+ $X2=3.355 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A21BOI_2%VPWR 1 2 3 10 12 18 22 26 28 36 43 44 50 53
c53 18 0 1.88192e-19 $X=2.68 $Y=2.375
r54 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r55 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r57 44 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r58 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r59 41 53 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.765 $Y=3.33
+ $X2=3.59 $Y2=3.33
r60 41 43 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.765 $Y=3.33
+ $X2=4.08 $Y2=3.33
r61 40 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r62 40 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r64 37 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=2.68 $Y2=3.33
r65 37 39 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=3.12 $Y2=3.33
r66 36 53 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.415 $Y=3.33
+ $X2=3.59 $Y2=3.33
r67 36 39 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.415 $Y=3.33
+ $X2=3.12 $Y2=3.33
r68 32 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r69 31 34 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r70 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r71 29 47 3.92346 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r72 29 31 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r73 28 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.515 $Y=3.33
+ $X2=2.68 $Y2=3.33
r74 28 34 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.515 $Y=3.33
+ $X2=2.16 $Y2=3.33
r75 26 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r76 26 32 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=0.72 $Y2=3.33
r77 26 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r78 22 25 22.3903 $w=3.48e-07 $l=6.8e-07 $layer=LI1_cond $X=3.59 $Y=2.145
+ $X2=3.59 $Y2=2.825
r79 20 53 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.59 $Y=3.245
+ $X2=3.59 $Y2=3.33
r80 20 25 13.8293 $w=3.48e-07 $l=4.2e-07 $layer=LI1_cond $X=3.59 $Y=3.245
+ $X2=3.59 $Y2=2.825
r81 16 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=3.245
+ $X2=2.68 $Y2=3.33
r82 16 18 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=2.68 $Y=3.245
+ $X2=2.68 $Y2=2.375
r83 12 15 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=0.32 $Y=2.115 $X2=0.32
+ $Y2=2.815
r84 10 47 3.2197 $w=2.5e-07 $l=1.33918e-07 $layer=LI1_cond $X=0.32 $Y=3.245
+ $X2=0.222 $Y2=3.33
r85 10 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.32 $Y=3.245
+ $X2=0.32 $Y2=2.815
r86 3 25 400 $w=1.7e-07 $l=1.05501e-06 $layer=licon1_PDIFF $count=1 $X=3.445
+ $Y=1.84 $X2=3.59 $Y2=2.825
r87 3 22 400 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_PDIFF $count=1 $X=3.445
+ $Y=1.84 $X2=3.59 $Y2=2.145
r88 2 18 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=2.545
+ $Y=1.84 $X2=2.68 $Y2=2.375
r89 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.235
+ $Y=1.96 $X2=0.36 $Y2=2.815
r90 1 12 400 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=0.235
+ $Y=1.96 $X2=0.36 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__A21BOI_2%A_241_368# 1 2 3 4 15 19 20 21 25 29 31 35
+ 41
c59 21 0 1.50652e-19 $X=2.215 $Y=2.12
r60 41 44 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.13 $Y=1.805
+ $X2=3.13 $Y2=1.985
r61 35 37 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=4.09 $Y=1.985
+ $X2=4.09 $Y2=2.815
r62 33 35 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=4.09 $Y=1.89
+ $X2=4.09 $Y2=1.985
r63 32 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=1.805
+ $X2=3.13 $Y2=1.805
r64 31 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.965 $Y=1.805
+ $X2=4.09 $Y2=1.89
r65 31 32 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=3.965 $Y=1.805
+ $X2=3.215 $Y2=1.805
r66 27 44 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.13 $Y=2.12
+ $X2=3.13 $Y2=1.985
r67 27 29 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.13 $Y=2.12
+ $X2=3.13 $Y2=2.4
r68 26 40 3.60116 $w=1.7e-07 $l=1.28452e-07 $layer=LI1_cond $X=2.315 $Y=2.035
+ $X2=2.215 $Y2=1.97
r69 25 44 0.716491 $w=1.7e-07 $l=1.07121e-07 $layer=LI1_cond $X=3.045 $Y=2.035
+ $X2=3.13 $Y2=1.985
r70 25 26 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.045 $Y=2.035
+ $X2=2.315 $Y2=2.035
r71 22 24 28.0045 $w=1.98e-07 $l=5.05e-07 $layer=LI1_cond $X=2.215 $Y=2.905
+ $X2=2.215 $Y2=2.4
r72 21 40 3.27378 $w=2e-07 $l=1.5e-07 $layer=LI1_cond $X=2.215 $Y=2.12 $X2=2.215
+ $Y2=1.97
r73 21 24 15.5273 $w=1.98e-07 $l=2.8e-07 $layer=LI1_cond $X=2.215 $Y=2.12
+ $X2=2.215 $Y2=2.4
r74 19 22 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.115 $Y=2.99
+ $X2=2.215 $Y2=2.905
r75 19 20 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.115 $Y=2.99
+ $X2=1.415 $Y2=2.99
r76 15 18 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=1.29 $Y=1.985
+ $X2=1.29 $Y2=2.815
r77 13 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.29 $Y=2.905
+ $X2=1.415 $Y2=2.99
r78 13 18 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.29 $Y=2.905 $X2=1.29
+ $Y2=2.815
r79 4 37 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.915
+ $Y=1.84 $X2=4.05 $Y2=2.815
r80 4 35 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.915
+ $Y=1.84 $X2=4.05 $Y2=1.985
r81 3 44 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.995
+ $Y=1.84 $X2=3.13 $Y2=1.985
r82 3 29 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=2.995
+ $Y=1.84 $X2=3.13 $Y2=2.4
r83 2 40 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.095
+ $Y=1.84 $X2=2.23 $Y2=1.985
r84 2 24 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=2.095
+ $Y=1.84 $X2=2.23 $Y2=2.4
r85 1 18 400 $w=1.7e-07 $l=1.03562e-06 $layer=licon1_PDIFF $count=1 $X=1.205
+ $Y=1.84 $X2=1.33 $Y2=2.815
r86 1 15 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.205
+ $Y=1.84 $X2=1.33 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__A21BOI_2%Y 1 2 3 12 15 18 22 25 29 32 35
c56 22 0 2.70769e-20 $X=2.57 $Y=1.065
r57 31 32 8.78489 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.78 $Y=1.195
+ $X2=1.615 $Y2=1.195
r58 29 35 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.16 $Y=1.195
+ $X2=2.275 $Y2=1.195
r59 29 31 10.1844 $w=4.28e-07 $l=3.8e-07 $layer=LI1_cond $X=2.16 $Y=1.195
+ $X2=1.78 $Y2=1.195
r60 25 27 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.735 $Y=0.91
+ $X2=2.735 $Y2=1.065
r61 22 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.57 $Y=1.065
+ $X2=2.735 $Y2=1.065
r62 22 35 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.57 $Y=1.065
+ $X2=2.275 $Y2=1.065
r63 18 20 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=1.78 $Y=1.965
+ $X2=1.78 $Y2=2.65
r64 16 31 2.28972 $w=3.3e-07 $l=2.15e-07 $layer=LI1_cond $X=1.78 $Y=1.41
+ $X2=1.78 $Y2=1.195
r65 16 18 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=1.78 $Y=1.41
+ $X2=1.78 $Y2=1.965
r66 15 32 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.44 $Y=1.065
+ $X2=1.615 $Y2=1.065
r67 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.355 $Y=0.98
+ $X2=1.44 $Y2=1.065
r68 10 12 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=1.355 $Y=0.98
+ $X2=1.355 $Y2=0.515
r69 3 20 400 $w=1.7e-07 $l=8.749e-07 $layer=licon1_PDIFF $count=1 $X=1.645
+ $Y=1.84 $X2=1.78 $Y2=2.65
r70 3 18 400 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=1.645
+ $Y=1.84 $X2=1.78 $Y2=1.965
r71 2 25 182 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_NDIFF $count=1 $X=2.595
+ $Y=0.37 $X2=2.735 $Y2=0.91
r72 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.215
+ $Y=0.37 $X2=1.355 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A21BOI_2%VGND 1 2 3 12 16 20 24 26 27 28 34 44 45 48
+ 51
r59 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r60 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r61 45 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r62 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r63 42 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.595
+ $Y2=0
r64 42 44 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=4.08
+ $Y2=0
r65 41 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r66 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r67 37 40 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r68 35 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.95 $Y=0 $X2=1.785
+ $Y2=0
r69 35 37 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.95 $Y=0 $X2=2.16
+ $Y2=0
r70 34 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.43 $Y=0 $X2=3.595
+ $Y2=0
r71 34 40 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.43 $Y=0 $X2=3.12
+ $Y2=0
r72 32 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r73 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r74 28 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r75 28 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r76 28 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r77 26 31 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=0.76 $Y=0 $X2=0.72
+ $Y2=0
r78 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.76 $Y=0 $X2=0.925
+ $Y2=0
r79 22 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=0.085
+ $X2=3.595 $Y2=0
r80 22 24 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.595 $Y=0.085
+ $X2=3.595 $Y2=0.55
r81 18 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=0.085
+ $X2=1.785 $Y2=0
r82 18 20 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=1.785 $Y=0.085
+ $X2=1.785 $Y2=0.645
r83 17 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.09 $Y=0 $X2=0.925
+ $Y2=0
r84 16 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.62 $Y=0 $X2=1.785
+ $Y2=0
r85 16 17 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.62 $Y=0 $X2=1.09
+ $Y2=0
r86 12 14 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.925 $Y=0.515
+ $X2=0.925 $Y2=0.855
r87 10 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.925 $Y=0.085
+ $X2=0.925 $Y2=0
r88 10 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.925 $Y=0.085
+ $X2=0.925 $Y2=0.515
r89 3 24 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.455 $Y=0.37
+ $X2=3.595 $Y2=0.55
r90 2 20 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.645
+ $Y=0.37 $X2=1.785 $Y2=0.645
r91 1 14 182 $w=1.7e-07 $l=4.74579e-07 $layer=licon1_NDIFF $count=1 $X=0.725
+ $Y=0.47 $X2=0.925 $Y2=0.855
r92 1 12 182 $w=1.7e-07 $l=2.21359e-07 $layer=licon1_NDIFF $count=1 $X=0.725
+ $Y=0.47 $X2=0.925 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A21BOI_2%A_436_74# 1 2 3 10 14 15 16 18 20
c33 14 0 1.6164e-19 $X=3.165 $Y=0.6
r34 18 27 3.13866 $w=2.5e-07 $l=1.45e-07 $layer=LI1_cond $X=4.065 $Y=0.84
+ $X2=4.065 $Y2=0.985
r35 18 20 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=4.065 $Y=0.84
+ $X2=4.065 $Y2=0.515
r36 17 25 3.40825 $w=1.7e-07 $l=9.44722e-08 $layer=LI1_cond $X=3.25 $Y=0.925
+ $X2=3.165 $Y2=0.945
r37 16 27 4.0045 $w=1.7e-07 $l=1.52069e-07 $layer=LI1_cond $X=3.94 $Y=0.925
+ $X2=4.065 $Y2=0.985
r38 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.94 $Y=0.925
+ $X2=3.25 $Y2=0.925
r39 15 25 3.40825 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.165 $Y=0.84
+ $X2=3.165 $Y2=0.945
r40 14 23 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.165 $Y=0.6
+ $X2=3.165 $Y2=0.475
r41 14 15 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.165 $Y=0.6
+ $X2=3.165 $Y2=0.84
r42 10 23 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.475
+ $X2=3.165 $Y2=0.475
r43 10 12 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=3.08 $Y=0.475
+ $X2=2.305 $Y2=0.475
r44 3 27 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.37 $X2=4.025 $Y2=0.965
r45 3 20 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.37 $X2=4.025 $Y2=0.515
r46 2 25 182 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_NDIFF $count=1 $X=3.025
+ $Y=0.37 $X2=3.165 $Y2=0.885
r47 2 23 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.025
+ $Y=0.37 $X2=3.165 $Y2=0.515
r48 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.18
+ $Y=0.37 $X2=2.305 $Y2=0.515
.ends


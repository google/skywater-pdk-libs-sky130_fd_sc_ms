* File: sky130_fd_sc_ms__clkbuf_16.spice
* Created: Wed Sep  2 12:00:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__clkbuf_16.pex.spice"
.subckt sky130_fd_sc_ms__clkbuf_16  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_A_114_74#_M1000_d N_A_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75008.8
+ A=0.063 P=1.14 MULT=1
MM1024 N_A_114_74#_M1000_d N_A_M1024_g N_VGND_M1024_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.063 PD=0.7 PS=0.72 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75008.4
+ A=0.063 P=1.14 MULT=1
MM1032 N_A_114_74#_M1032_d N_A_M1032_g N_VGND_M1024_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.063 PD=0.7 PS=0.72 NRD=0 NRS=5.712 M=1 R=2.8 SA=75001.1
+ SB=75007.9 A=0.063 P=1.14 MULT=1
MM1033 N_A_114_74#_M1032_d N_A_M1033_g N_VGND_M1033_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0735 PD=0.7 PS=0.77 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75007.5
+ A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1033_s N_A_114_74#_M1001_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8 SA=75002
+ SB=75007 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_114_74#_M1002_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.4 SB=75006.6
+ A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1002_d N_A_114_74#_M1008_g N_X_M1008_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.9 SB=75006.1
+ A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_114_74#_M1010_g N_X_M1008_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75003.3 SB=75005.7
+ A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1010_d N_A_114_74#_M1012_g N_X_M1012_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75003.7 SB=75005.3
+ A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_A_114_74#_M1014_g N_X_M1012_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75004.2 SB=75004.9
+ A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1014_d N_A_114_74#_M1015_g N_X_M1015_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8 SA=75004.7
+ SB=75004.4 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_114_74#_M1016_g N_X_M1015_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75005.1 SB=75003.9
+ A=0.063 P=1.14 MULT=1
MM1018 N_VGND_M1016_d N_A_114_74#_M1018_g N_X_M1018_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8 SA=75005.6
+ SB=75003.4 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_114_74#_M1019_g N_X_M1018_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75006 SB=75003
+ A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1019_d N_A_114_74#_M1020_g N_X_M1020_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8 SA=75006.5
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_A_114_74#_M1021_g N_X_M1020_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75007 SB=75002.1
+ A=0.063 P=1.14 MULT=1
MM1028 N_VGND_M1021_d N_A_114_74#_M1028_g N_X_M1028_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8 SA=75007.5
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_A_114_74#_M1029_g N_X_M1028_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75007.9 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1034 N_VGND_M1029_d N_A_114_74#_M1034_g N_X_M1034_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.0588 PD=0.77 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8 SA=75008.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1037 N_VGND_M1037_d N_A_114_74#_M1037_g N_X_M1034_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75008.8 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1003 N_A_114_74#_M1003_d N_A_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90008.8 A=0.2016 P=2.6 MULT=1
MM1004 N_A_114_74#_M1003_d N_A_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90008.3 A=0.2016 P=2.6 MULT=1
MM1006 N_A_114_74#_M1006_d N_A_M1006_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90007.9 A=0.2016 P=2.6 MULT=1
MM1007 N_A_114_74#_M1006_d N_A_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1568 PD=1.39 PS=1.4 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90007.4 A=0.2016 P=2.6 MULT=1
MM1005 N_X_M1005_d N_A_114_74#_M1005_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1568 PD=1.39 PS=1.4 NRD=0 NRS=0.8668 M=1 R=6.22222 SA=90002
+ SB=90007 A=0.2016 P=2.6 MULT=1
MM1009 N_X_M1005_d N_A_114_74#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.4
+ SB=90006.5 A=0.2016 P=2.6 MULT=1
MM1011 N_X_M1011_d N_A_114_74#_M1011_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.9
+ SB=90006.1 A=0.2016 P=2.6 MULT=1
MM1013 N_X_M1011_d N_A_114_74#_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.3
+ SB=90005.6 A=0.2016 P=2.6 MULT=1
MM1017 N_X_M1017_d N_A_114_74#_M1017_g N_VPWR_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.8
+ SB=90005.2 A=0.2016 P=2.6 MULT=1
MM1022 N_X_M1017_d N_A_114_74#_M1022_g N_VPWR_M1022_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.2
+ SB=90004.7 A=0.2016 P=2.6 MULT=1
MM1023 N_X_M1023_d N_A_114_74#_M1023_g N_VPWR_M1022_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.7
+ SB=90004.3 A=0.2016 P=2.6 MULT=1
MM1025 N_X_M1023_d N_A_114_74#_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90005.1
+ SB=90003.8 A=0.2016 P=2.6 MULT=1
MM1026 N_X_M1026_d N_A_114_74#_M1026_g N_VPWR_M1025_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90005.6
+ SB=90003.4 A=0.2016 P=2.6 MULT=1
MM1027 N_X_M1026_d N_A_114_74#_M1027_g N_VPWR_M1027_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90006
+ SB=90002.9 A=0.2016 P=2.6 MULT=1
MM1030 N_X_M1030_d N_A_114_74#_M1030_g N_VPWR_M1027_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90006.5
+ SB=90002.5 A=0.2016 P=2.6 MULT=1
MM1031 N_X_M1030_d N_A_114_74#_M1031_g N_VPWR_M1031_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90006.9
+ SB=90002 A=0.2016 P=2.6 MULT=1
MM1035 N_X_M1035_d N_A_114_74#_M1035_g N_VPWR_M1031_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90007.4
+ SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1036 N_X_M1035_d N_A_114_74#_M1036_g N_VPWR_M1036_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1624 PD=1.39 PS=1.41 NRD=0 NRS=0 M=1 R=6.22222 SA=90007.8
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1038 N_X_M1038_d N_A_114_74#_M1038_g N_VPWR_M1036_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1624 PD=1.39 PS=1.41 NRD=0 NRS=2.6201 M=1 R=6.22222 SA=90008.3
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1039 N_X_M1038_d N_A_114_74#_M1039_g N_VPWR_M1039_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90008.8
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX40_noxref VNB VPB NWDIODE A=18.5628 P=23.68
*
.include "sky130_fd_sc_ms__clkbuf_16.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__o22ai_1.pxi.spice
* Created: Wed Sep  2 12:23:49 2020
* 
x_PM_SKY130_FD_SC_MS__O22AI_1%B1 N_B1_c_48_n N_B1_M1006_g N_B1_M1005_g B1
+ N_B1_c_51_n PM_SKY130_FD_SC_MS__O22AI_1%B1
x_PM_SKY130_FD_SC_MS__O22AI_1%B2 N_B2_M1000_g N_B2_M1003_g B2 N_B2_c_77_n
+ N_B2_c_78_n PM_SKY130_FD_SC_MS__O22AI_1%B2
x_PM_SKY130_FD_SC_MS__O22AI_1%A2 N_A2_M1007_g N_A2_M1002_g A2 N_A2_c_108_n
+ N_A2_c_109_n PM_SKY130_FD_SC_MS__O22AI_1%A2
x_PM_SKY130_FD_SC_MS__O22AI_1%A1 N_A1_M1001_g N_A1_M1004_g N_A1_c_148_n A1 A1
+ N_A1_c_150_n PM_SKY130_FD_SC_MS__O22AI_1%A1
x_PM_SKY130_FD_SC_MS__O22AI_1%VPWR N_VPWR_M1005_s N_VPWR_M1001_d N_VPWR_c_179_n
+ N_VPWR_c_180_n N_VPWR_c_181_n N_VPWR_c_182_n N_VPWR_c_183_n N_VPWR_c_184_n
+ VPWR N_VPWR_c_178_n PM_SKY130_FD_SC_MS__O22AI_1%VPWR
x_PM_SKY130_FD_SC_MS__O22AI_1%Y N_Y_M1006_d N_Y_M1000_d N_Y_c_206_n Y Y
+ N_Y_c_208_n N_Y_c_207_n PM_SKY130_FD_SC_MS__O22AI_1%Y
x_PM_SKY130_FD_SC_MS__O22AI_1%A_27_74# N_A_27_74#_M1006_s N_A_27_74#_M1003_d
+ N_A_27_74#_M1004_d N_A_27_74#_c_237_n N_A_27_74#_c_238_n N_A_27_74#_c_239_n
+ N_A_27_74#_c_251_n N_A_27_74#_c_240_n N_A_27_74#_c_241_n N_A_27_74#_c_242_n
+ PM_SKY130_FD_SC_MS__O22AI_1%A_27_74#
x_PM_SKY130_FD_SC_MS__O22AI_1%VGND N_VGND_M1002_d N_VGND_c_278_n N_VGND_c_279_n
+ N_VGND_c_280_n VGND N_VGND_c_281_n N_VGND_c_282_n
+ PM_SKY130_FD_SC_MS__O22AI_1%VGND
cc_1 VNB N_B1_c_48_n 0.0245603f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_2 VNB N_B1_M1005_g 0.00857766f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.4
cc_3 VNB B1 0.00820169f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_B1_c_51_n 0.0715868f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.385
cc_5 VNB N_B2_M1003_g 0.0285891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_B2_c_77_n 0.0253507f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_7 VNB N_B2_c_78_n 0.00694829f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.385
cc_8 VNB N_A2_M1002_g 0.0268957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A2_c_108_n 0.0269875f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_10 VNB N_A2_c_109_n 0.00181735f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.385
cc_11 VNB N_A1_M1001_g 0.00172115f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_12 VNB N_A1_M1004_g 0.0317431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_c_148_n 0.0182188f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_14 VNB A1 0.0177202f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_15 VNB N_A1_c_150_n 0.0481093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_178_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_206_n 0.00809472f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_18 VNB N_Y_c_207_n 0.00612152f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_c_237_n 0.0200157f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_20 VNB N_A_27_74#_c_238_n 0.00778015f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.55
cc_21 VNB N_A_27_74#_c_239_n 0.00972033f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.295
cc_22 VNB N_A_27_74#_c_240_n 0.0168726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_74#_c_241_n 0.00894964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_74#_c_242_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_278_n 0.0095417f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.4
cc_26 VNB N_VGND_c_279_n 0.0477009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_280_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_28 VNB N_VGND_c_281_n 0.0221746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_282_n 0.188569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VPB N_B1_M1005_g 0.0272611f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=2.4
cc_31 VPB N_B2_M1000_g 0.0225007f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_32 VPB N_B2_c_77_n 0.0055692f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.385
cc_33 VPB N_B2_c_78_n 0.0023831f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.385
cc_34 VPB N_A2_M1007_g 0.0242106f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_35 VPB N_A2_c_108_n 0.00566891f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.385
cc_36 VPB N_A2_c_109_n 0.00637181f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.385
cc_37 VPB N_A1_M1001_g 0.0282233f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_38 VPB A1 0.0182295f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.385
cc_39 VPB N_VPWR_c_179_n 0.0125099f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_180_n 0.0594498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_181_n 0.0484149f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.295
cc_42 VPB N_VPWR_c_182_n 0.0115308f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_183_n 0.0498476f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_184_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_178_n 0.076907f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_Y_c_208_n 0.00542649f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.385
cc_47 VPB N_Y_c_207_n 0.00129681f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 N_B1_M1005_g N_B2_M1000_g 0.0454889f $X=0.635 $Y=2.4 $X2=0 $Y2=0
cc_49 N_B1_c_48_n N_B2_M1003_g 0.0175332f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_50 N_B1_c_51_n N_B2_c_77_n 0.0467209f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_51 N_B1_c_51_n N_B2_c_78_n 4.20038e-19 $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_52 N_B1_M1005_g N_VPWR_c_180_n 0.030275f $X=0.635 $Y=2.4 $X2=0 $Y2=0
cc_53 B1 N_VPWR_c_180_n 0.0192059f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_54 N_B1_c_51_n N_VPWR_c_180_n 0.00281221f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_55 N_B1_M1005_g N_VPWR_c_183_n 0.00441589f $X=0.635 $Y=2.4 $X2=0 $Y2=0
cc_56 N_B1_M1005_g N_VPWR_c_178_n 0.00730287f $X=0.635 $Y=2.4 $X2=0 $Y2=0
cc_57 N_B1_c_48_n N_Y_c_206_n 0.0041759f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_58 N_B1_c_51_n N_Y_c_206_n 3.73516e-19 $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_59 N_B1_M1005_g N_Y_c_208_n 0.0285831f $X=0.635 $Y=2.4 $X2=0 $Y2=0
cc_60 N_B1_c_48_n N_Y_c_207_n 0.00431169f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_61 N_B1_M1005_g N_Y_c_207_n 0.0167133f $X=0.635 $Y=2.4 $X2=0 $Y2=0
cc_62 B1 N_Y_c_207_n 0.0260309f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_63 N_B1_c_51_n N_Y_c_207_n 0.00663293f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_64 N_B1_c_48_n N_A_27_74#_c_237_n 0.0118446f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_65 B1 N_A_27_74#_c_237_n 0.0261036f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_66 N_B1_c_51_n N_A_27_74#_c_237_n 0.00199342f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_67 N_B1_c_48_n N_A_27_74#_c_238_n 0.0116366f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_68 N_B1_c_48_n N_A_27_74#_c_239_n 0.00167496f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_69 N_B1_c_48_n N_VGND_c_279_n 0.00286814f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_70 N_B1_c_48_n N_VGND_c_282_n 0.00361864f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_71 N_B2_M1000_g N_A2_M1007_g 0.0279268f $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_72 N_B2_M1003_g N_A2_M1002_g 0.0250863f $X=1.22 $Y=0.74 $X2=0 $Y2=0
cc_73 N_B2_c_77_n N_A2_c_108_n 0.0175474f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_74 N_B2_c_78_n N_A2_c_108_n 0.00274004f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_75 N_B2_c_77_n N_A2_c_109_n 4.06701e-19 $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_76 N_B2_c_78_n N_A2_c_109_n 0.0281717f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_77 N_B2_M1000_g N_VPWR_c_183_n 0.00349816f $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_78 N_B2_M1000_g N_VPWR_c_178_n 0.00430348f $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_79 N_B2_M1003_g N_Y_c_206_n 0.00587202f $X=1.22 $Y=0.74 $X2=0 $Y2=0
cc_80 N_B2_c_77_n N_Y_c_206_n 7.12446e-19 $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_81 N_B2_c_78_n N_Y_c_206_n 0.00676358f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_82 N_B2_M1000_g N_Y_c_208_n 0.0325006f $X=1.055 $Y=2.4 $X2=0 $Y2=0
cc_83 N_B2_c_77_n N_Y_c_208_n 7.69767e-19 $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_84 N_B2_c_78_n N_Y_c_208_n 0.027039f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_85 N_B2_M1003_g N_Y_c_207_n 0.00318696f $X=1.22 $Y=0.74 $X2=0 $Y2=0
cc_86 N_B2_c_77_n N_Y_c_207_n 0.0049319f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_87 N_B2_c_78_n N_Y_c_207_n 0.0324255f $X=1.13 $Y=1.515 $X2=0 $Y2=0
cc_88 N_B2_M1003_g N_A_27_74#_c_238_n 0.0157492f $X=1.22 $Y=0.74 $X2=0 $Y2=0
cc_89 N_B2_M1003_g N_A_27_74#_c_241_n 0.00100357f $X=1.22 $Y=0.74 $X2=0 $Y2=0
cc_90 N_B2_M1003_g N_VGND_c_279_n 0.00286838f $X=1.22 $Y=0.74 $X2=0 $Y2=0
cc_91 N_B2_M1003_g N_VGND_c_282_n 0.0035893f $X=1.22 $Y=0.74 $X2=0 $Y2=0
cc_92 N_A2_M1007_g N_A1_M1001_g 0.0426063f $X=1.625 $Y=2.4 $X2=0 $Y2=0
cc_93 N_A2_c_109_n N_A1_M1001_g 3.30229e-19 $X=1.7 $Y=1.515 $X2=0 $Y2=0
cc_94 N_A2_M1002_g N_A1_M1004_g 0.0250949f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_95 N_A2_M1002_g N_A1_c_148_n 0.00181425f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_96 N_A2_c_108_n N_A1_c_148_n 0.0174347f $X=1.7 $Y=1.515 $X2=0 $Y2=0
cc_97 N_A2_c_109_n N_A1_c_148_n 3.69555e-19 $X=1.7 $Y=1.515 $X2=0 $Y2=0
cc_98 N_A2_M1007_g A1 3.07828e-19 $X=1.625 $Y=2.4 $X2=0 $Y2=0
cc_99 N_A2_M1002_g A1 0.00123883f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_100 N_A2_c_108_n A1 0.00216744f $X=1.7 $Y=1.515 $X2=0 $Y2=0
cc_101 N_A2_c_109_n A1 0.0350655f $X=1.7 $Y=1.515 $X2=0 $Y2=0
cc_102 N_A2_M1007_g N_VPWR_c_181_n 0.00518719f $X=1.625 $Y=2.4 $X2=0 $Y2=0
cc_103 N_A2_M1007_g N_VPWR_c_183_n 0.00537895f $X=1.625 $Y=2.4 $X2=0 $Y2=0
cc_104 N_A2_M1007_g N_VPWR_c_178_n 0.0104067f $X=1.625 $Y=2.4 $X2=0 $Y2=0
cc_105 N_A2_M1007_g N_Y_c_208_n 0.0380253f $X=1.625 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A2_c_109_n N_Y_c_208_n 0.00106339f $X=1.7 $Y=1.515 $X2=0 $Y2=0
cc_107 N_A2_M1002_g N_A_27_74#_c_238_n 0.00272067f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_108 N_A2_M1002_g N_A_27_74#_c_251_n 0.00730256f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_109 N_A2_M1002_g N_A_27_74#_c_240_n 0.0120407f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_110 N_A2_c_108_n N_A_27_74#_c_240_n 4.60538e-19 $X=1.7 $Y=1.515 $X2=0 $Y2=0
cc_111 N_A2_c_109_n N_A_27_74#_c_240_n 0.0118018f $X=1.7 $Y=1.515 $X2=0 $Y2=0
cc_112 N_A2_M1002_g N_A_27_74#_c_241_n 0.00102901f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_113 N_A2_c_108_n N_A_27_74#_c_241_n 8.26843e-19 $X=1.7 $Y=1.515 $X2=0 $Y2=0
cc_114 N_A2_c_109_n N_A_27_74#_c_241_n 0.00940645f $X=1.7 $Y=1.515 $X2=0 $Y2=0
cc_115 N_A2_M1002_g N_A_27_74#_c_242_n 6.18925e-19 $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A2_M1002_g N_VGND_c_278_n 0.00522681f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_117 N_A2_M1002_g N_VGND_c_279_n 0.00432337f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_118 N_A2_M1002_g N_VGND_c_282_n 0.00817838f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_119 N_A1_M1001_g N_VPWR_c_181_n 0.0274317f $X=2.195 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A1_c_148_n N_VPWR_c_181_n 0.00151573f $X=2.235 $Y=1.465 $X2=0 $Y2=0
cc_121 A1 N_VPWR_c_181_n 0.0264613f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_122 N_A1_M1001_g N_VPWR_c_183_n 0.00460063f $X=2.195 $Y=2.4 $X2=0 $Y2=0
cc_123 N_A1_M1001_g N_VPWR_c_178_n 0.00909693f $X=2.195 $Y=2.4 $X2=0 $Y2=0
cc_124 N_A1_M1001_g N_Y_c_208_n 0.00452194f $X=2.195 $Y=2.4 $X2=0 $Y2=0
cc_125 N_A1_M1004_g N_A_27_74#_c_251_n 5.91875e-19 $X=2.29 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A1_M1004_g N_A_27_74#_c_240_n 0.0129307f $X=2.29 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A1_c_148_n N_A_27_74#_c_240_n 0.00289965f $X=2.235 $Y=1.465 $X2=0 $Y2=0
cc_128 A1 N_A_27_74#_c_240_n 0.0509938f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_129 N_A1_c_150_n N_A_27_74#_c_240_n 0.00708493f $X=2.61 $Y=1.465 $X2=0 $Y2=0
cc_130 N_A1_M1004_g N_A_27_74#_c_242_n 0.00981823f $X=2.29 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A1_M1004_g N_VGND_c_278_n 0.00592235f $X=2.29 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A1_M1004_g N_VGND_c_281_n 0.00434272f $X=2.29 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A1_M1004_g N_VGND_c_282_n 0.00825253f $X=2.29 $Y=0.74 $X2=0 $Y2=0
cc_134 N_VPWR_c_183_n N_Y_c_208_n 0.0402719f $X=2.255 $Y=3.33 $X2=0 $Y2=0
cc_135 N_VPWR_c_178_n N_Y_c_208_n 0.0326649f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_136 N_VPWR_c_180_n N_Y_c_207_n 0.0945274f $X=0.29 $Y=1.985 $X2=0 $Y2=0
cc_137 A_145_368# N_Y_c_208_n 0.00509749f $X=0.725 $Y=1.84 $X2=1.335 $Y2=2.115
cc_138 A_145_368# N_Y_c_207_n 6.959e-19 $X=0.725 $Y=1.84 $X2=1.087 $Y2=1.95
cc_139 N_Y_M1006_d N_A_27_74#_c_238_n 0.00691776f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_140 N_Y_c_206_n N_A_27_74#_c_238_n 0.0331049f $X=0.855 $Y=0.84 $X2=0 $Y2=0
cc_141 N_Y_c_206_n N_A_27_74#_c_241_n 0.00568934f $X=0.855 $Y=0.84 $X2=0 $Y2=0
cc_142 N_A_27_74#_c_240_n N_VGND_M1002_d 0.00374767f $X=2.34 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_143 N_A_27_74#_c_238_n N_VGND_c_278_n 0.0094172f $X=1.34 $Y=0.4 $X2=0 $Y2=0
cc_144 N_A_27_74#_c_240_n N_VGND_c_278_n 0.0248957f $X=2.34 $Y=1.045 $X2=0 $Y2=0
cc_145 N_A_27_74#_c_242_n N_VGND_c_278_n 0.0173003f $X=2.505 $Y=0.515 $X2=0
+ $Y2=0
cc_146 N_A_27_74#_c_238_n N_VGND_c_279_n 0.0581922f $X=1.34 $Y=0.4 $X2=0 $Y2=0
cc_147 N_A_27_74#_c_239_n N_VGND_c_279_n 0.0170692f $X=0.445 $Y=0.4 $X2=0 $Y2=0
cc_148 N_A_27_74#_c_242_n N_VGND_c_281_n 0.0145639f $X=2.505 $Y=0.515 $X2=0
+ $Y2=0
cc_149 N_A_27_74#_c_238_n N_VGND_c_282_n 0.0434237f $X=1.34 $Y=0.4 $X2=0 $Y2=0
cc_150 N_A_27_74#_c_239_n N_VGND_c_282_n 0.0123284f $X=0.445 $Y=0.4 $X2=0 $Y2=0
cc_151 N_A_27_74#_c_242_n N_VGND_c_282_n 0.0119984f $X=2.505 $Y=0.515 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__o31ai_1.pxi.spice
* Created: Fri Aug 28 18:02:49 2020
* 
x_PM_SKY130_FD_SC_MS__O31AI_1%A1 N_A1_c_46_n N_A1_M1005_g N_A1_M1003_g A1
+ N_A1_c_49_n PM_SKY130_FD_SC_MS__O31AI_1%A1
x_PM_SKY130_FD_SC_MS__O31AI_1%A2 N_A2_M1006_g N_A2_M1000_g A2 A2 A2 A2
+ N_A2_c_71_n N_A2_c_72_n PM_SKY130_FD_SC_MS__O31AI_1%A2
x_PM_SKY130_FD_SC_MS__O31AI_1%A3 N_A3_M1007_g N_A3_M1001_g A3 N_A3_c_111_n
+ PM_SKY130_FD_SC_MS__O31AI_1%A3
x_PM_SKY130_FD_SC_MS__O31AI_1%B1 N_B1_M1002_g N_B1_M1004_g B1 N_B1_c_145_n
+ N_B1_c_146_n PM_SKY130_FD_SC_MS__O31AI_1%B1
x_PM_SKY130_FD_SC_MS__O31AI_1%VPWR N_VPWR_M1003_s N_VPWR_M1004_d N_VPWR_c_170_n
+ N_VPWR_c_171_n N_VPWR_c_172_n N_VPWR_c_173_n VPWR N_VPWR_c_174_n
+ N_VPWR_c_169_n PM_SKY130_FD_SC_MS__O31AI_1%VPWR
x_PM_SKY130_FD_SC_MS__O31AI_1%Y N_Y_M1002_d N_Y_M1007_d N_Y_c_200_n N_Y_c_201_n
+ N_Y_c_202_n Y Y N_Y_c_204_n N_Y_c_203_n PM_SKY130_FD_SC_MS__O31AI_1%Y
x_PM_SKY130_FD_SC_MS__O31AI_1%VGND N_VGND_M1005_s N_VGND_M1006_d N_VGND_c_242_n
+ N_VGND_c_243_n VGND N_VGND_c_244_n N_VGND_c_245_n N_VGND_c_246_n
+ N_VGND_c_247_n PM_SKY130_FD_SC_MS__O31AI_1%VGND
x_PM_SKY130_FD_SC_MS__O31AI_1%A_114_74# N_A_114_74#_M1005_d N_A_114_74#_M1001_d
+ N_A_114_74#_c_282_n N_A_114_74#_c_278_n N_A_114_74#_c_279_n
+ N_A_114_74#_c_280_n PM_SKY130_FD_SC_MS__O31AI_1%A_114_74#
cc_1 VNB N_A1_c_46_n 0.0213825f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_2 VNB N_A1_M1003_g 0.00857766f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=2.4
cc_3 VNB A1 0.0103026f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A1_c_49_n 0.0599265f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.385
cc_5 VNB N_A2_M1006_g 0.0235915f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_6 VNB N_A2_M1000_g 0.00139203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A2_c_71_n 0.0329091f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_8 VNB N_A2_c_72_n 0.00639141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A3_M1001_g 0.026895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB A3 0.0037708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A3_c_111_n 0.0356322f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.385
cc_12 VNB N_B1_M1002_g 0.0302921f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_13 VNB N_B1_M1004_g 0.0015157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B1_c_145_n 0.0597714f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_15 VNB N_B1_c_146_n 0.00461578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_169_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_200_n 0.0150819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_201_n 3.20099e-19 $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_19 VNB N_Y_c_202_n 0.0262708f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.385
cc_20 VNB N_Y_c_203_n 0.00868892f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_242_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_243_n 0.0337878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_244_n 0.0319663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_245_n 0.179964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_246_n 0.0164203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_247_n 0.0228461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_114_74#_c_278_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_28 VNB N_A_114_74#_c_279_n 0.00231275f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.385
cc_29 VNB N_A_114_74#_c_280_n 0.002553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VPB N_A1_M1003_g 0.0273807f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=2.4
cc_31 VPB N_A2_M1000_g 0.0224514f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB N_A2_c_72_n 0.00114345f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_33 VPB N_A3_M1007_g 0.0257107f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_34 VPB A3 0.00680374f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_A3_c_111_n 0.0134181f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.385
cc_36 VPB N_B1_M1004_g 0.0293495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_37 VPB N_B1_c_146_n 0.00926033f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_170_n 0.0111306f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_171_n 0.0563955f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_172_n 0.0127942f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.385
cc_41 VPB N_VPWR_c_173_n 0.0484147f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.295
cc_42 VPB N_VPWR_c_174_n 0.0537421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_169_n 0.0655869f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_Y_c_204_n 0.00669049f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_Y_c_203_n 0.00117058f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 N_A1_c_46_n N_A2_M1006_g 0.0106343f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_47 A1 N_A2_M1006_g 5.69588e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_48 N_A1_M1003_g N_A2_M1000_g 0.0463449f $X=0.52 $Y=2.4 $X2=0 $Y2=0
cc_49 N_A1_c_49_n N_A2_c_71_n 0.0569792f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_50 N_A1_M1003_g N_A2_c_72_n 0.038071f $X=0.52 $Y=2.4 $X2=0 $Y2=0
cc_51 A1 N_A2_c_72_n 0.0200321f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_52 N_A1_c_49_n N_A2_c_72_n 0.00472914f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_53 N_A1_M1003_g N_VPWR_c_171_n 0.00684253f $X=0.52 $Y=2.4 $X2=0 $Y2=0
cc_54 A1 N_VPWR_c_171_n 0.0149782f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_55 N_A1_c_49_n N_VPWR_c_171_n 0.00185549f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_56 N_A1_M1003_g N_VPWR_c_174_n 0.00549539f $X=0.52 $Y=2.4 $X2=0 $Y2=0
cc_57 N_A1_M1003_g N_VPWR_c_169_n 0.0107381f $X=0.52 $Y=2.4 $X2=0 $Y2=0
cc_58 N_A1_c_46_n N_VGND_c_243_n 0.0130745f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_59 A1 N_VGND_c_243_n 0.025255f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_60 N_A1_c_49_n N_VGND_c_243_n 0.00199898f $X=0.495 $Y=1.385 $X2=0 $Y2=0
cc_61 N_A1_c_46_n N_VGND_c_245_n 0.00757637f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_62 N_A1_c_46_n N_VGND_c_246_n 0.00383152f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_63 N_A1_c_46_n N_A_114_74#_c_278_n 8.89831e-19 $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_64 N_A2_c_71_n N_A3_M1001_g 5.59819e-19 $X=1.015 $Y=1.465 $X2=0 $Y2=0
cc_65 N_A2_M1000_g N_A3_c_111_n 0.0428901f $X=0.94 $Y=2.4 $X2=0 $Y2=0
cc_66 N_A2_c_71_n N_A3_c_111_n 0.00845062f $X=1.015 $Y=1.465 $X2=0 $Y2=0
cc_67 N_A2_c_72_n N_A3_c_111_n 0.00455628f $X=1.015 $Y=1.465 $X2=0 $Y2=0
cc_68 N_A2_c_72_n N_VPWR_c_171_n 0.0355557f $X=1.015 $Y=1.465 $X2=0 $Y2=0
cc_69 N_A2_M1000_g N_VPWR_c_174_n 0.00363952f $X=0.94 $Y=2.4 $X2=0 $Y2=0
cc_70 N_A2_c_72_n N_VPWR_c_174_n 0.0153197f $X=1.015 $Y=1.465 $X2=0 $Y2=0
cc_71 N_A2_M1000_g N_VPWR_c_169_n 0.00445545f $X=0.94 $Y=2.4 $X2=0 $Y2=0
cc_72 N_A2_c_72_n N_VPWR_c_169_n 0.0190617f $X=1.015 $Y=1.465 $X2=0 $Y2=0
cc_73 N_A2_c_72_n A_122_368# 0.00175001f $X=1.015 $Y=1.465 $X2=-0.19 $Y2=-0.245
cc_74 N_A2_c_72_n A_206_368# 0.0106388f $X=1.015 $Y=1.465 $X2=-0.19 $Y2=-0.245
cc_75 N_A2_M1006_g N_Y_c_201_n 0.00330111f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_76 N_A2_M1000_g N_Y_c_204_n 0.00217055f $X=0.94 $Y=2.4 $X2=0 $Y2=0
cc_77 N_A2_M1006_g N_Y_c_203_n 0.00477786f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_78 N_A2_M1000_g N_Y_c_203_n 0.00365144f $X=0.94 $Y=2.4 $X2=0 $Y2=0
cc_79 N_A2_c_71_n N_Y_c_203_n 0.00267004f $X=1.015 $Y=1.465 $X2=0 $Y2=0
cc_80 N_A2_c_72_n N_Y_c_203_n 0.135014f $X=1.015 $Y=1.465 $X2=0 $Y2=0
cc_81 N_A2_M1006_g N_VGND_c_243_n 5.69788e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_82 N_A2_M1006_g N_VGND_c_245_n 0.00404728f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_83 N_A2_M1006_g N_VGND_c_246_n 0.00320194f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_84 N_A2_M1006_g N_VGND_c_247_n 0.00531017f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_85 N_A2_M1006_g N_A_114_74#_c_282_n 0.0122762f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_86 N_A2_c_71_n N_A_114_74#_c_282_n 7.85402e-19 $X=1.015 $Y=1.465 $X2=0 $Y2=0
cc_87 N_A2_c_72_n N_A_114_74#_c_282_n 0.008902f $X=1.015 $Y=1.465 $X2=0 $Y2=0
cc_88 N_A2_M1006_g N_A_114_74#_c_278_n 0.010161f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_89 N_A2_M1006_g N_A_114_74#_c_279_n 0.0107236f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_90 N_A2_c_72_n N_A_114_74#_c_279_n 0.0230199f $X=1.015 $Y=1.465 $X2=0 $Y2=0
cc_91 N_A3_M1001_g N_B1_M1002_g 0.0316207f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_92 N_A3_M1007_g N_B1_M1004_g 0.0071017f $X=1.51 $Y=2.4 $X2=0 $Y2=0
cc_93 A3 N_B1_M1004_g 0.0047681f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_94 A3 N_B1_c_145_n 0.00748727f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_95 N_A3_c_111_n N_B1_c_145_n 0.0181891f $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_96 N_A3_M1001_g N_B1_c_146_n 2.15196e-19 $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_97 A3 N_B1_c_146_n 0.0343232f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_98 N_A3_M1007_g N_VPWR_c_174_n 0.00349816f $X=1.51 $Y=2.4 $X2=0 $Y2=0
cc_99 N_A3_M1007_g N_VPWR_c_169_n 0.00433306f $X=1.51 $Y=2.4 $X2=0 $Y2=0
cc_100 N_A3_M1001_g N_Y_c_200_n 0.0125598f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_101 A3 N_Y_c_200_n 0.0374035f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_102 N_A3_c_111_n N_Y_c_200_n 0.00890833f $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_103 N_A3_M1007_g N_Y_c_204_n 0.0310236f $X=1.51 $Y=2.4 $X2=0 $Y2=0
cc_104 A3 N_Y_c_204_n 0.0464791f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_105 N_A3_c_111_n N_Y_c_204_n 0.00410852f $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_106 N_A3_M1007_g N_Y_c_203_n 0.0115939f $X=1.51 $Y=2.4 $X2=0 $Y2=0
cc_107 N_A3_M1001_g N_Y_c_203_n 0.00612746f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_108 A3 N_Y_c_203_n 0.0332669f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_109 N_A3_c_111_n N_Y_c_203_n 0.00720293f $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_110 N_A3_M1001_g N_VGND_c_244_n 0.00320194f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_111 N_A3_M1001_g N_VGND_c_245_n 0.00404912f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_112 N_A3_M1001_g N_VGND_c_247_n 0.00703231f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_113 N_A3_M1001_g N_A_114_74#_c_282_n 0.0108636f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_114 N_A3_M1001_g N_A_114_74#_c_280_n 0.0106282f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_115 N_B1_M1004_g N_VPWR_c_173_n 0.0217046f $X=2.35 $Y=2.4 $X2=0 $Y2=0
cc_116 N_B1_c_145_n N_VPWR_c_173_n 0.00150147f $X=2.61 $Y=1.465 $X2=0 $Y2=0
cc_117 N_B1_c_146_n N_VPWR_c_173_n 0.0239693f $X=2.61 $Y=1.465 $X2=0 $Y2=0
cc_118 N_B1_M1004_g N_VPWR_c_174_n 0.00460063f $X=2.35 $Y=2.4 $X2=0 $Y2=0
cc_119 N_B1_M1004_g N_VPWR_c_169_n 0.00911329f $X=2.35 $Y=2.4 $X2=0 $Y2=0
cc_120 N_B1_M1002_g N_Y_c_200_n 0.0174305f $X=2.335 $Y=0.74 $X2=0 $Y2=0
cc_121 N_B1_c_145_n N_Y_c_200_n 0.00405369f $X=2.61 $Y=1.465 $X2=0 $Y2=0
cc_122 N_B1_c_146_n N_Y_c_200_n 0.0277433f $X=2.61 $Y=1.465 $X2=0 $Y2=0
cc_123 N_B1_M1002_g N_Y_c_202_n 0.00164953f $X=2.335 $Y=0.74 $X2=0 $Y2=0
cc_124 N_B1_M1004_g N_Y_c_204_n 2.67293e-19 $X=2.35 $Y=2.4 $X2=0 $Y2=0
cc_125 N_B1_M1002_g N_VGND_c_244_n 0.00456932f $X=2.335 $Y=0.74 $X2=0 $Y2=0
cc_126 N_B1_M1002_g N_VGND_c_245_n 0.00894956f $X=2.335 $Y=0.74 $X2=0 $Y2=0
cc_127 N_B1_M1002_g N_A_114_74#_c_280_n 0.004688f $X=2.335 $Y=0.74 $X2=0 $Y2=0
cc_128 N_VPWR_c_173_n N_Y_c_204_n 0.0377637f $X=2.575 $Y=2.115 $X2=0 $Y2=0
cc_129 N_VPWR_c_174_n N_Y_c_204_n 0.0386391f $X=2.41 $Y=3.33 $X2=0 $Y2=0
cc_130 N_VPWR_c_169_n N_Y_c_204_n 0.0315593f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_131 A_206_368# N_Y_c_204_n 0.00978205f $X=1.03 $Y=1.84 $X2=1.015 $Y2=1.3
cc_132 A_206_368# N_Y_c_203_n 9.66534e-19 $X=1.03 $Y=1.84 $X2=1.015 $Y2=1.63
cc_133 N_Y_c_200_n N_VGND_M1006_d 0.00337116f $X=2.435 $Y=1.045 $X2=0 $Y2=0
cc_134 N_Y_c_201_n N_VGND_M1006_d 0.00548721f $X=1.52 $Y=1.045 $X2=0 $Y2=0
cc_135 N_Y_c_202_n N_VGND_c_244_n 0.0146357f $X=2.6 $Y=0.515 $X2=0 $Y2=0
cc_136 N_Y_c_202_n N_VGND_c_245_n 0.0121141f $X=2.6 $Y=0.515 $X2=0 $Y2=0
cc_137 N_Y_c_200_n N_A_114_74#_M1001_d 0.00197722f $X=2.435 $Y=1.045 $X2=0 $Y2=0
cc_138 N_Y_c_200_n N_A_114_74#_c_282_n 0.0253598f $X=2.435 $Y=1.045 $X2=0 $Y2=0
cc_139 N_Y_c_201_n N_A_114_74#_c_282_n 0.013831f $X=1.52 $Y=1.045 $X2=0 $Y2=0
cc_140 N_Y_c_201_n N_A_114_74#_c_279_n 0.0062517f $X=1.52 $Y=1.045 $X2=0 $Y2=0
cc_141 N_Y_c_200_n N_A_114_74#_c_280_n 0.016668f $X=2.435 $Y=1.045 $X2=0 $Y2=0
cc_142 N_Y_c_202_n N_A_114_74#_c_280_n 0.0173003f $X=2.6 $Y=0.515 $X2=0 $Y2=0
cc_143 N_VGND_M1006_d N_A_114_74#_c_282_n 0.023923f $X=1 $Y=0.37 $X2=0 $Y2=0
cc_144 N_VGND_c_244_n N_A_114_74#_c_282_n 0.00266409f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_145 N_VGND_c_245_n N_A_114_74#_c_282_n 0.0123863f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_146 N_VGND_c_246_n N_A_114_74#_c_282_n 0.00266409f $X=1.055 $Y=0.182 $X2=0
+ $Y2=0
cc_147 N_VGND_c_247_n N_A_114_74#_c_282_n 0.0525207f $X=1.755 $Y=0.182 $X2=0
+ $Y2=0
cc_148 N_VGND_c_243_n N_A_114_74#_c_278_n 0.0243832f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_149 N_VGND_c_245_n N_A_114_74#_c_278_n 0.00904371f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_150 N_VGND_c_246_n N_A_114_74#_c_278_n 0.0109942f $X=1.055 $Y=0.182 $X2=0
+ $Y2=0
cc_151 N_VGND_c_247_n N_A_114_74#_c_278_n 0.00426994f $X=1.755 $Y=0.182 $X2=0
+ $Y2=0
cc_152 N_VGND_c_244_n N_A_114_74#_c_280_n 0.0141059f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_153 N_VGND_c_245_n N_A_114_74#_c_280_n 0.0118064f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_154 N_VGND_c_247_n N_A_114_74#_c_280_n 0.00441839f $X=1.755 $Y=0.182 $X2=0
+ $Y2=0

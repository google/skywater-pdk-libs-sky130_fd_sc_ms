* File: sky130_fd_sc_ms__o32ai_2.pxi.spice
* Created: Fri Aug 28 18:04:16 2020
* 
x_PM_SKY130_FD_SC_MS__O32AI_2%B2 N_B2_M1002_g N_B2_M1015_g N_B2_M1016_g
+ N_B2_M1003_g B2 B2 B2 N_B2_c_100_n PM_SKY130_FD_SC_MS__O32AI_2%B2
x_PM_SKY130_FD_SC_MS__O32AI_2%B1 N_B1_M1004_g N_B1_M1011_g N_B1_M1005_g
+ N_B1_M1013_g B1 N_B1_c_144_n N_B1_c_145_n PM_SKY130_FD_SC_MS__O32AI_2%B1
x_PM_SKY130_FD_SC_MS__O32AI_2%A3 N_A3_M1008_g N_A3_M1017_g N_A3_M1009_g
+ N_A3_M1019_g A3 A3 N_A3_c_199_n PM_SKY130_FD_SC_MS__O32AI_2%A3
x_PM_SKY130_FD_SC_MS__O32AI_2%A2 N_A2_M1014_g N_A2_M1000_g N_A2_M1001_g
+ N_A2_M1018_g A2 A2 N_A2_c_258_n PM_SKY130_FD_SC_MS__O32AI_2%A2
x_PM_SKY130_FD_SC_MS__O32AI_2%A1 N_A1_M1007_g N_A1_M1006_g N_A1_M1010_g
+ N_A1_M1012_g N_A1_c_306_n A1 A1 A1 A1 N_A1_c_308_n N_A1_c_309_n
+ PM_SKY130_FD_SC_MS__O32AI_2%A1
x_PM_SKY130_FD_SC_MS__O32AI_2%A_27_368# N_A_27_368#_M1002_s N_A_27_368#_M1003_s
+ N_A_27_368#_M1005_s N_A_27_368#_c_351_n N_A_27_368#_c_352_n
+ N_A_27_368#_c_353_n N_A_27_368#_c_366_p N_A_27_368#_c_359_n
+ N_A_27_368#_c_354_n PM_SKY130_FD_SC_MS__O32AI_2%A_27_368#
x_PM_SKY130_FD_SC_MS__O32AI_2%Y N_Y_M1015_d N_Y_M1011_s N_Y_M1002_d N_Y_M1017_d
+ N_Y_c_390_n N_Y_c_382_n N_Y_c_383_n N_Y_c_387_n N_Y_c_413_n N_Y_c_384_n
+ N_Y_c_401_n N_Y_c_385_n Y Y N_Y_c_388_n N_Y_c_386_n
+ PM_SKY130_FD_SC_MS__O32AI_2%Y
x_PM_SKY130_FD_SC_MS__O32AI_2%VPWR N_VPWR_M1004_d N_VPWR_M1006_d N_VPWR_M1010_d
+ N_VPWR_c_469_n N_VPWR_c_470_n N_VPWR_c_471_n N_VPWR_c_472_n VPWR
+ N_VPWR_c_473_n N_VPWR_c_474_n N_VPWR_c_475_n N_VPWR_c_476_n N_VPWR_c_477_n
+ N_VPWR_c_468_n PM_SKY130_FD_SC_MS__O32AI_2%VPWR
x_PM_SKY130_FD_SC_MS__O32AI_2%A_499_368# N_A_499_368#_M1017_s
+ N_A_499_368#_M1019_s N_A_499_368#_M1001_s N_A_499_368#_c_532_n
+ N_A_499_368#_c_533_n N_A_499_368#_c_534_n N_A_499_368#_c_541_n
+ N_A_499_368#_c_535_n N_A_499_368#_c_536_n N_A_499_368#_c_537_n
+ PM_SKY130_FD_SC_MS__O32AI_2%A_499_368#
x_PM_SKY130_FD_SC_MS__O32AI_2%A_771_368# N_A_771_368#_M1000_d
+ N_A_771_368#_M1006_s N_A_771_368#_c_566_n N_A_771_368#_c_576_n
+ N_A_771_368#_c_567_n N_A_771_368#_c_570_n
+ PM_SKY130_FD_SC_MS__O32AI_2%A_771_368#
x_PM_SKY130_FD_SC_MS__O32AI_2%A_27_74# N_A_27_74#_M1015_s N_A_27_74#_M1016_s
+ N_A_27_74#_M1013_d N_A_27_74#_M1009_s N_A_27_74#_M1018_s N_A_27_74#_M1012_d
+ N_A_27_74#_c_592_n N_A_27_74#_c_593_n N_A_27_74#_c_594_n N_A_27_74#_c_609_n
+ N_A_27_74#_c_595_n N_A_27_74#_c_615_n N_A_27_74#_c_616_n N_A_27_74#_c_619_n
+ N_A_27_74#_c_620_n N_A_27_74#_c_596_n N_A_27_74#_c_597_n N_A_27_74#_c_598_n
+ N_A_27_74#_c_599_n N_A_27_74#_c_600_n N_A_27_74#_c_601_n N_A_27_74#_c_602_n
+ N_A_27_74#_c_603_n PM_SKY130_FD_SC_MS__O32AI_2%A_27_74#
x_PM_SKY130_FD_SC_MS__O32AI_2%VGND N_VGND_M1008_d N_VGND_M1014_d N_VGND_M1007_s
+ N_VGND_c_683_n N_VGND_c_684_n N_VGND_c_685_n VGND N_VGND_c_686_n
+ N_VGND_c_687_n N_VGND_c_688_n N_VGND_c_689_n N_VGND_c_690_n N_VGND_c_691_n
+ PM_SKY130_FD_SC_MS__O32AI_2%VGND
cc_1 VNB N_B2_M1015_g 0.0312487f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_B2_M1016_g 0.0234839f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_3 VNB B2 0.0183784f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_4 VNB N_B2_c_100_n 0.0436935f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.515
cc_5 VNB N_B1_M1011_g 0.0244803f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_6 VNB N_B1_M1013_g 0.0244812f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_7 VNB N_B1_c_144_n 0.0015808f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_8 VNB N_B1_c_145_n 0.0402406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A3_M1008_g 0.0281248f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_10 VNB N_A3_M1009_g 0.0287756f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_11 VNB A3 0.00626365f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_12 VNB N_A3_c_199_n 0.0602501f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.515
cc_13 VNB N_A2_M1014_g 0.0246043f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_14 VNB N_A2_M1018_g 0.0247047f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_15 VNB A2 0.00438466f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_16 VNB N_A2_c_258_n 0.0353344f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.515
cc_17 VNB N_A1_M1007_g 0.0305737f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_18 VNB N_A1_M1012_g 0.0393239f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_19 VNB N_A1_c_306_n 0.00935177f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_20 VNB A1 0.0203068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_c_308_n 0.0219884f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.515
cc_22 VNB N_A1_c_309_n 0.0398575f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_23 VNB N_Y_c_382_n 0.00349006f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_24 VNB N_Y_c_383_n 0.00229732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_384_n 0.0091475f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.515
cc_26 VNB N_Y_c_385_n 0.0033895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_386_n 0.00357335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_468_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_74#_c_592_n 0.0288468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_74#_c_593_n 0.0026914f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_31 VNB N_A_27_74#_c_594_n 0.00931596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_74#_c_595_n 0.00501991f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.515
cc_33 VNB N_A_27_74#_c_596_n 0.00291303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_27_74#_c_597_n 0.00565856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_74#_c_598_n 0.00280814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_27_74#_c_599_n 0.017779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_27_74#_c_600_n 0.0277086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_27_74#_c_601_n 0.00220635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_74#_c_602_n 0.00280429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_27_74#_c_603_n 0.00725128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_683_n 0.00582196f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_684_n 0.0181004f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_43 VNB N_VGND_c_685_n 0.00616254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_686_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.565
cc_45 VNB N_VGND_c_687_n 0.334788f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_46 VNB N_VGND_c_688_n 0.060757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_689_n 0.0195534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_690_n 0.018682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_691_n 0.0300631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VPB N_B2_M1002_g 0.0252952f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_51 VPB N_B2_M1003_g 0.0197873f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_52 VPB B2 0.0145149f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_53 VPB N_B2_c_100_n 0.00734846f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.515
cc_54 VPB N_B1_M1004_g 0.0202002f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_55 VPB N_B1_M1005_g 0.0251433f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_56 VPB N_B1_c_144_n 0.00251564f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.515
cc_57 VPB N_B1_c_145_n 0.00464585f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A3_M1017_g 0.0243179f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_59 VPB N_A3_M1019_g 0.0206154f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_60 VPB A3 0.0085226f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_61 VPB N_A3_c_199_n 0.0173781f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.515
cc_62 VPB N_A2_M1000_g 0.0197858f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_63 VPB N_A2_M1001_g 0.0244741f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_64 VPB A2 0.00676776f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_65 VPB N_A2_c_258_n 0.00458006f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.515
cc_66 VPB N_A1_M1006_g 0.0246944f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_67 VPB N_A1_M1010_g 0.0247049f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_68 VPB N_A1_c_306_n 0.0048851f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_69 VPB A1 0.0198762f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A1_c_308_n 0.0129865f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.515
cc_71 VPB N_A1_c_309_n 0.00463455f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_72 VPB N_A_27_368#_c_351_n 0.0354954f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_27_368#_c_352_n 0.00473643f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_27_368#_c_353_n 0.00929469f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_75 VPB N_A_27_368#_c_354_n 0.00891286f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.515
cc_76 VPB N_Y_c_387_n 0.0120361f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_Y_c_388_n 0.00411182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_Y_c_386_n 0.00115453f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_469_n 0.00554449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_470_n 0.0157535f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_471_n 0.0107598f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_82 VPB N_VPWR_c_472_n 0.0495391f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_473_n 0.0375062f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.515
cc_84 VPB N_VPWR_c_474_n 0.076072f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_475_n 0.0197695f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_476_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_477_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_468_n 0.092217f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_499_368#_c_532_n 0.00553942f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_499_368#_c_533_n 0.0026202f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_91 VPB N_A_499_368#_c_534_n 0.00446997f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_92 VPB N_A_499_368#_c_535_n 0.00643559f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_499_368#_c_536_n 0.00571534f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.515
cc_94 VPB N_A_499_368#_c_537_n 0.00123754f $X=-0.19 $Y=1.66 $X2=0.835 $Y2=1.515
cc_95 VPB N_A_771_368#_c_566_n 0.011775f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.35
cc_96 VPB N_A_771_368#_c_567_n 0.00235902f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.68
cc_97 N_B2_M1003_g N_B1_M1004_g 0.0251003f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_98 N_B2_M1016_g N_B1_M1011_g 0.0301413f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_99 B2 N_B1_c_144_n 0.0340851f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_100 N_B2_c_100_n N_B1_c_144_n 2.75325e-19 $X=0.955 $Y=1.515 $X2=0 $Y2=0
cc_101 B2 N_B1_c_145_n 0.00443562f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_102 N_B2_c_100_n N_B1_c_145_n 0.0251003f $X=0.955 $Y=1.515 $X2=0 $Y2=0
cc_103 B2 N_A_27_368#_c_351_n 0.0208754f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_104 N_B2_M1002_g N_A_27_368#_c_352_n 0.01495f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_105 N_B2_M1003_g N_A_27_368#_c_352_n 0.0137017f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_106 N_B2_M1015_g N_Y_c_390_n 0.00516364f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_107 N_B2_M1016_g N_Y_c_390_n 0.00668237f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_108 N_B2_M1016_g N_Y_c_382_n 0.00933793f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_109 B2 N_Y_c_382_n 0.0344043f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_110 N_B2_c_100_n N_Y_c_382_n 0.00118622f $X=0.955 $Y=1.515 $X2=0 $Y2=0
cc_111 N_B2_M1015_g N_Y_c_383_n 0.00605998f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_112 N_B2_M1016_g N_Y_c_383_n 0.00277595f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_113 B2 N_Y_c_383_n 0.0277268f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_114 N_B2_c_100_n N_Y_c_383_n 0.00241236f $X=0.955 $Y=1.515 $X2=0 $Y2=0
cc_115 N_B2_M1003_g N_Y_c_387_n 0.0128923f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_116 B2 N_Y_c_387_n 0.0282763f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_117 N_B2_M1002_g N_Y_c_401_n 0.0114036f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_118 N_B2_M1003_g N_Y_c_401_n 0.0105298f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_119 B2 N_Y_c_401_n 0.0235495f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_120 N_B2_c_100_n N_Y_c_401_n 5.53716e-19 $X=0.955 $Y=1.515 $X2=0 $Y2=0
cc_121 N_B2_M1002_g N_VPWR_c_473_n 0.00333926f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_122 N_B2_M1003_g N_VPWR_c_473_n 0.00333926f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_123 N_B2_M1002_g N_VPWR_c_468_n 0.00426429f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_124 N_B2_M1003_g N_VPWR_c_468_n 0.00422798f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_125 N_B2_M1015_g N_A_27_74#_c_592_n 0.00159289f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_126 B2 N_A_27_74#_c_592_n 0.0178256f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_127 N_B2_c_100_n N_A_27_74#_c_592_n 7.71522e-19 $X=0.955 $Y=1.515 $X2=0 $Y2=0
cc_128 N_B2_M1015_g N_A_27_74#_c_593_n 0.0132764f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_129 N_B2_M1016_g N_A_27_74#_c_593_n 0.0111757f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_130 N_B2_M1015_g N_VGND_c_687_n 0.00357086f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_131 N_B2_M1016_g N_VGND_c_687_n 0.0035414f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_132 N_B2_M1015_g N_VGND_c_688_n 0.00278271f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_133 N_B2_M1016_g N_VGND_c_688_n 0.00278271f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_134 N_B1_M1013_g N_A3_M1008_g 0.0178748f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_135 N_B1_c_144_n A3 0.0288593f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_136 N_B1_c_145_n A3 0.00634473f $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_137 N_B1_c_144_n N_A3_c_199_n 2.25325e-19 $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_138 N_B1_c_145_n N_A3_c_199_n 0.0226324f $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_139 N_B1_M1004_g N_A_27_368#_c_352_n 0.00101073f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_140 N_B1_M1004_g N_A_27_368#_c_359_n 0.0140196f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_141 N_B1_M1005_g N_A_27_368#_c_359_n 0.0126573f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_142 N_B1_M1004_g N_A_27_368#_c_354_n 5.87944e-19 $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_143 N_B1_M1005_g N_A_27_368#_c_354_n 0.00913184f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_144 N_B1_M1011_g N_Y_c_390_n 5.09814e-19 $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_145 N_B1_M1011_g N_Y_c_382_n 0.0170272f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_146 N_B1_c_144_n N_Y_c_382_n 0.00445816f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_147 N_B1_c_145_n N_Y_c_382_n 0.00145272f $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_148 N_B1_M1004_g N_Y_c_387_n 0.0167852f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_149 N_B1_M1005_g N_Y_c_387_n 0.0177843f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_150 N_B1_c_144_n N_Y_c_387_n 0.0217013f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_151 N_B1_c_145_n N_Y_c_387_n 4.89526e-19 $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_152 N_B1_M1013_g N_Y_c_413_n 0.0064205f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_153 N_B1_M1013_g N_Y_c_384_n 0.0129057f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_154 N_B1_M1004_g N_Y_c_401_n 7.43219e-19 $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_155 N_B1_M1013_g N_Y_c_385_n 0.00404963f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_156 N_B1_c_144_n N_Y_c_385_n 0.0228889f $X=1.65 $Y=1.515 $X2=0 $Y2=0
cc_157 N_B1_c_145_n N_Y_c_385_n 0.00131074f $X=1.855 $Y=1.515 $X2=0 $Y2=0
cc_158 N_B1_M1004_g N_VPWR_c_469_n 0.00769625f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_159 N_B1_M1005_g N_VPWR_c_469_n 0.002979f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_160 N_B1_M1004_g N_VPWR_c_473_n 0.00460063f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_161 N_B1_M1005_g N_VPWR_c_474_n 0.005209f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_162 N_B1_M1004_g N_VPWR_c_468_n 0.00908665f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_163 N_B1_M1005_g N_VPWR_c_468_n 0.00987399f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_164 N_B1_M1005_g N_A_499_368#_c_534_n 0.00292778f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_165 N_B1_M1011_g N_A_27_74#_c_609_n 0.00668986f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_166 N_B1_M1013_g N_A_27_74#_c_609_n 5.09814e-19 $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_167 N_B1_M1011_g N_A_27_74#_c_595_n 0.00831967f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_168 N_B1_M1013_g N_A_27_74#_c_595_n 0.011569f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_169 N_B1_M1011_g N_A_27_74#_c_601_n 0.00288559f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_170 N_B1_M1011_g N_VGND_c_687_n 0.00354796f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_171 N_B1_M1013_g N_VGND_c_687_n 0.00354798f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_172 N_B1_M1011_g N_VGND_c_688_n 0.00278247f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_173 N_B1_M1013_g N_VGND_c_688_n 0.00278271f $X=1.925 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A3_M1009_g N_A2_M1014_g 0.0150421f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A3_M1019_g N_A2_M1000_g 0.0122378f $X=3.315 $Y=2.4 $X2=0 $Y2=0
cc_176 N_A3_c_199_n A2 0.0053632f $X=3.255 $Y=1.515 $X2=0 $Y2=0
cc_177 N_A3_c_199_n N_A2_c_258_n 0.02728f $X=3.255 $Y=1.515 $X2=0 $Y2=0
cc_178 N_A3_M1017_g N_Y_c_387_n 0.0204188f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_179 A3 N_Y_c_387_n 0.0555676f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_180 N_A3_c_199_n N_Y_c_387_n 0.0021247f $X=3.255 $Y=1.515 $X2=0 $Y2=0
cc_181 N_A3_M1008_g N_Y_c_413_n 8.78205e-19 $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A3_M1008_g N_Y_c_384_n 0.0121505f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_183 N_A3_M1009_g N_Y_c_384_n 0.00213938f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_184 A3 N_Y_c_384_n 0.0552068f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_185 N_A3_c_199_n N_Y_c_384_n 0.0106593f $X=3.255 $Y=1.515 $X2=0 $Y2=0
cc_186 N_A3_M1017_g Y 0.0157053f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A3_M1019_g Y 0.00996565f $X=3.315 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A3_M1017_g N_Y_c_388_n 0.00697813f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_189 N_A3_M1019_g N_Y_c_388_n 0.00622698f $X=3.315 $Y=2.4 $X2=0 $Y2=0
cc_190 N_A3_c_199_n N_Y_c_388_n 0.00199936f $X=3.255 $Y=1.515 $X2=0 $Y2=0
cc_191 N_A3_M1008_g N_Y_c_386_n 0.00299821f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A3_M1017_g N_Y_c_386_n 0.00375683f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_193 N_A3_M1009_g N_Y_c_386_n 0.00459856f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A3_M1019_g N_Y_c_386_n 0.00172226f $X=3.315 $Y=2.4 $X2=0 $Y2=0
cc_195 A3 N_Y_c_386_n 0.0331353f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_196 N_A3_c_199_n N_Y_c_386_n 0.0195181f $X=3.255 $Y=1.515 $X2=0 $Y2=0
cc_197 N_A3_M1017_g N_VPWR_c_474_n 0.00333926f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_198 N_A3_M1019_g N_VPWR_c_474_n 0.00333926f $X=3.315 $Y=2.4 $X2=0 $Y2=0
cc_199 N_A3_M1017_g N_VPWR_c_468_n 0.0042782f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_200 N_A3_M1019_g N_VPWR_c_468_n 0.00422798f $X=3.315 $Y=2.4 $X2=0 $Y2=0
cc_201 N_A3_M1017_g N_A_499_368#_c_533_n 0.0149887f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_202 N_A3_M1019_g N_A_499_368#_c_533_n 0.0139961f $X=3.315 $Y=2.4 $X2=0 $Y2=0
cc_203 N_A3_M1008_g N_A_27_74#_c_595_n 0.00401363f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_204 N_A3_M1008_g N_A_27_74#_c_615_n 0.00816247f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_205 N_A3_M1008_g N_A_27_74#_c_616_n 0.00998617f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A3_M1009_g N_A_27_74#_c_616_n 0.0143601f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A3_c_199_n N_A_27_74#_c_616_n 9.64261e-19 $X=3.255 $Y=1.515 $X2=0 $Y2=0
cc_208 N_A3_M1008_g N_A_27_74#_c_619_n 0.00134994f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_209 N_A3_M1009_g N_A_27_74#_c_620_n 0.00728117f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_210 N_A3_M1009_g N_A_27_74#_c_597_n 0.00424559f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A3_c_199_n N_A_27_74#_c_597_n 0.00299651f $X=3.255 $Y=1.515 $X2=0 $Y2=0
cc_212 N_A3_M1009_g N_A_27_74#_c_602_n 0.0111563f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A3_M1009_g N_VGND_c_683_n 6.70813e-19 $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A3_M1009_g N_VGND_c_684_n 0.00324657f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A3_M1008_g N_VGND_c_687_n 0.00413263f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A3_M1009_g N_VGND_c_687_n 0.00413208f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A3_M1008_g N_VGND_c_688_n 0.00321293f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A3_M1008_g N_VGND_c_689_n 0.00303822f $X=2.425 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A3_M1009_g N_VGND_c_689_n 0.00514433f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A2_M1018_g N_A1_M1007_g 0.0155173f $X=4.23 $Y=0.74 $X2=0 $Y2=0
cc_221 A2 N_A1_c_306_n 2.78011e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_222 N_A2_c_258_n N_A1_c_306_n 0.0155173f $X=4.23 $Y=1.515 $X2=0 $Y2=0
cc_223 A2 A1 0.0285909f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_224 N_A2_c_258_n A1 0.00549615f $X=4.23 $Y=1.515 $X2=0 $Y2=0
cc_225 N_A2_M1000_g N_Y_c_388_n 8.03043e-19 $X=3.765 $Y=2.4 $X2=0 $Y2=0
cc_226 A2 N_Y_c_386_n 0.0190657f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_227 N_A2_c_258_n N_Y_c_386_n 2.34445e-19 $X=4.23 $Y=1.515 $X2=0 $Y2=0
cc_228 N_A2_M1001_g N_VPWR_c_470_n 0.00196089f $X=4.215 $Y=2.4 $X2=0 $Y2=0
cc_229 N_A2_M1000_g N_VPWR_c_474_n 0.00333926f $X=3.765 $Y=2.4 $X2=0 $Y2=0
cc_230 N_A2_M1001_g N_VPWR_c_474_n 0.00333896f $X=4.215 $Y=2.4 $X2=0 $Y2=0
cc_231 N_A2_M1000_g N_VPWR_c_468_n 0.00422798f $X=3.765 $Y=2.4 $X2=0 $Y2=0
cc_232 N_A2_M1001_g N_VPWR_c_468_n 0.00427818f $X=4.215 $Y=2.4 $X2=0 $Y2=0
cc_233 A2 N_A_499_368#_c_541_n 0.012018f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_234 N_A2_M1000_g N_A_499_368#_c_535_n 0.0139518f $X=3.765 $Y=2.4 $X2=0 $Y2=0
cc_235 N_A2_M1001_g N_A_499_368#_c_535_n 0.014552f $X=4.215 $Y=2.4 $X2=0 $Y2=0
cc_236 N_A2_M1000_g N_A_499_368#_c_536_n 6.1567e-19 $X=3.765 $Y=2.4 $X2=0 $Y2=0
cc_237 N_A2_M1001_g N_A_499_368#_c_536_n 0.00912569f $X=4.215 $Y=2.4 $X2=0 $Y2=0
cc_238 N_A2_M1001_g N_A_771_368#_c_566_n 0.0197388f $X=4.215 $Y=2.4 $X2=0 $Y2=0
cc_239 A2 N_A_771_368#_c_566_n 0.00724026f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_240 N_A2_M1000_g N_A_771_368#_c_570_n 0.0107104f $X=3.765 $Y=2.4 $X2=0 $Y2=0
cc_241 A2 N_A_771_368#_c_570_n 0.0189743f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_242 N_A2_c_258_n N_A_771_368#_c_570_n 5.54777e-19 $X=4.23 $Y=1.515 $X2=0
+ $Y2=0
cc_243 N_A2_M1014_g N_A_27_74#_c_596_n 0.0151193f $X=3.75 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A2_M1018_g N_A_27_74#_c_596_n 0.0166108f $X=4.23 $Y=0.74 $X2=0 $Y2=0
cc_245 A2 N_A_27_74#_c_596_n 0.0423811f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_246 N_A2_c_258_n N_A_27_74#_c_596_n 0.00359948f $X=4.23 $Y=1.515 $X2=0 $Y2=0
cc_247 A2 N_A_27_74#_c_597_n 0.0135252f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_248 N_A2_M1018_g N_A_27_74#_c_598_n 4.71232e-19 $X=4.23 $Y=0.74 $X2=0 $Y2=0
cc_249 N_A2_M1014_g N_A_27_74#_c_602_n 0.00349724f $X=3.75 $Y=0.74 $X2=0 $Y2=0
cc_250 N_A2_M1018_g N_A_27_74#_c_603_n 8.63921e-19 $X=4.23 $Y=0.74 $X2=0 $Y2=0
cc_251 N_A2_M1014_g N_VGND_c_683_n 0.00955922f $X=3.75 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A2_M1018_g N_VGND_c_683_n 0.00230425f $X=4.23 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A2_M1014_g N_VGND_c_684_n 0.00398535f $X=3.75 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A2_M1014_g N_VGND_c_687_n 0.00788205f $X=3.75 $Y=0.74 $X2=0 $Y2=0
cc_255 N_A2_M1018_g N_VGND_c_687_n 0.00908353f $X=4.23 $Y=0.74 $X2=0 $Y2=0
cc_256 N_A2_M1018_g N_VGND_c_690_n 0.00461464f $X=4.23 $Y=0.74 $X2=0 $Y2=0
cc_257 N_A1_M1006_g N_VPWR_c_470_n 0.00534567f $X=5.275 $Y=2.4 $X2=0 $Y2=0
cc_258 N_A1_M1010_g N_VPWR_c_472_n 0.00501904f $X=5.73 $Y=2.4 $X2=0 $Y2=0
cc_259 A1 N_VPWR_c_472_n 0.0213263f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_260 N_A1_M1006_g N_VPWR_c_475_n 0.005209f $X=5.275 $Y=2.4 $X2=0 $Y2=0
cc_261 N_A1_M1010_g N_VPWR_c_475_n 0.005209f $X=5.73 $Y=2.4 $X2=0 $Y2=0
cc_262 N_A1_M1006_g N_VPWR_c_468_n 0.00986778f $X=5.275 $Y=2.4 $X2=0 $Y2=0
cc_263 N_A1_M1010_g N_VPWR_c_468_n 0.00986076f $X=5.73 $Y=2.4 $X2=0 $Y2=0
cc_264 N_A1_M1006_g N_A_771_368#_c_566_n 0.0150541f $X=5.275 $Y=2.4 $X2=0 $Y2=0
cc_265 N_A1_c_306_n N_A_771_368#_c_566_n 0.00300836f $X=4.76 $Y=1.515 $X2=0
+ $Y2=0
cc_266 A1 N_A_771_368#_c_566_n 0.0681406f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_267 N_A1_M1006_g N_A_771_368#_c_576_n 8.84614e-19 $X=5.275 $Y=2.4 $X2=0 $Y2=0
cc_268 N_A1_M1010_g N_A_771_368#_c_576_n 0.0025567f $X=5.73 $Y=2.4 $X2=0 $Y2=0
cc_269 A1 N_A_771_368#_c_576_n 0.0239914f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_270 N_A1_c_309_n N_A_771_368#_c_576_n 5.85598e-19 $X=5.745 $Y=1.515 $X2=0
+ $Y2=0
cc_271 N_A1_M1006_g N_A_771_368#_c_567_n 0.016262f $X=5.275 $Y=2.4 $X2=0 $Y2=0
cc_272 N_A1_M1010_g N_A_771_368#_c_567_n 0.0114458f $X=5.73 $Y=2.4 $X2=0 $Y2=0
cc_273 N_A1_M1007_g N_A_27_74#_c_598_n 0.0148256f $X=4.685 $Y=0.74 $X2=0 $Y2=0
cc_274 N_A1_M1007_g N_A_27_74#_c_599_n 0.0131906f $X=4.685 $Y=0.74 $X2=0 $Y2=0
cc_275 N_A1_M1012_g N_A_27_74#_c_599_n 0.0153378f $X=5.745 $Y=0.74 $X2=0 $Y2=0
cc_276 A1 N_A_27_74#_c_599_n 0.116536f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_277 N_A1_c_308_n N_A_27_74#_c_599_n 0.0175287f $X=5.185 $Y=1.515 $X2=0 $Y2=0
cc_278 N_A1_M1012_g N_A_27_74#_c_600_n 0.0155483f $X=5.745 $Y=0.74 $X2=0 $Y2=0
cc_279 N_A1_M1007_g N_A_27_74#_c_603_n 0.0016171f $X=4.685 $Y=0.74 $X2=0 $Y2=0
cc_280 A1 N_A_27_74#_c_603_n 0.0169123f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_281 N_A1_M1012_g N_VGND_c_686_n 0.00434272f $X=5.745 $Y=0.74 $X2=0 $Y2=0
cc_282 N_A1_M1007_g N_VGND_c_687_n 0.00825362f $X=4.685 $Y=0.74 $X2=0 $Y2=0
cc_283 N_A1_M1012_g N_VGND_c_687_n 0.00828694f $X=5.745 $Y=0.74 $X2=0 $Y2=0
cc_284 N_A1_M1007_g N_VGND_c_690_n 0.00434272f $X=4.685 $Y=0.74 $X2=0 $Y2=0
cc_285 N_A1_M1007_g N_VGND_c_691_n 0.00539931f $X=4.685 $Y=0.74 $X2=0 $Y2=0
cc_286 N_A1_M1012_g N_VGND_c_691_n 0.00705014f $X=5.745 $Y=0.74 $X2=0 $Y2=0
cc_287 N_A_27_368#_c_352_n N_Y_M1002_d 0.00165831f $X=1.095 $Y=2.99 $X2=0 $Y2=0
cc_288 N_A_27_368#_M1003_s N_Y_c_387_n 0.00332066f $X=1.045 $Y=1.84 $X2=0 $Y2=0
cc_289 N_A_27_368#_M1005_s N_Y_c_387_n 0.00685921f $X=1.945 $Y=1.84 $X2=0 $Y2=0
cc_290 N_A_27_368#_c_366_p N_Y_c_387_n 0.0126919f $X=1.18 $Y=2.46 $X2=0 $Y2=0
cc_291 N_A_27_368#_c_359_n N_Y_c_387_n 0.0336305f $X=1.915 $Y=2.375 $X2=0 $Y2=0
cc_292 N_A_27_368#_c_354_n N_Y_c_387_n 0.0221016f $X=2.08 $Y=2.455 $X2=0 $Y2=0
cc_293 N_A_27_368#_c_352_n N_Y_c_401_n 0.0159318f $X=1.095 $Y=2.99 $X2=0 $Y2=0
cc_294 N_A_27_368#_c_359_n N_VPWR_M1004_d 0.00324075f $X=1.915 $Y=2.375
+ $X2=-0.19 $Y2=1.66
cc_295 N_A_27_368#_c_352_n N_VPWR_c_469_n 0.010126f $X=1.095 $Y=2.99 $X2=0 $Y2=0
cc_296 N_A_27_368#_c_359_n N_VPWR_c_469_n 0.0148589f $X=1.915 $Y=2.375 $X2=0
+ $Y2=0
cc_297 N_A_27_368#_c_354_n N_VPWR_c_469_n 0.0122069f $X=2.08 $Y=2.455 $X2=0
+ $Y2=0
cc_298 N_A_27_368#_c_352_n N_VPWR_c_473_n 0.0581059f $X=1.095 $Y=2.99 $X2=0
+ $Y2=0
cc_299 N_A_27_368#_c_353_n N_VPWR_c_473_n 0.0179217f $X=0.365 $Y=2.99 $X2=0
+ $Y2=0
cc_300 N_A_27_368#_c_354_n N_VPWR_c_474_n 0.0145644f $X=2.08 $Y=2.455 $X2=0
+ $Y2=0
cc_301 N_A_27_368#_c_352_n N_VPWR_c_468_n 0.0324093f $X=1.095 $Y=2.99 $X2=0
+ $Y2=0
cc_302 N_A_27_368#_c_353_n N_VPWR_c_468_n 0.00971942f $X=0.365 $Y=2.99 $X2=0
+ $Y2=0
cc_303 N_A_27_368#_c_354_n N_VPWR_c_468_n 0.0119803f $X=2.08 $Y=2.455 $X2=0
+ $Y2=0
cc_304 N_A_27_368#_c_354_n N_A_499_368#_c_532_n 0.0412426f $X=2.08 $Y=2.455
+ $X2=0 $Y2=0
cc_305 N_A_27_368#_c_354_n N_A_499_368#_c_534_n 0.00536542f $X=2.08 $Y=2.455
+ $X2=0 $Y2=0
cc_306 N_Y_c_387_n N_VPWR_M1004_d 0.00314436f $X=2.925 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_307 N_Y_c_387_n N_A_499_368#_M1017_s 0.0052384f $X=2.925 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_308 N_Y_c_387_n N_A_499_368#_c_532_n 0.0197477f $X=2.925 $Y=2.035 $X2=0 $Y2=0
cc_309 N_Y_M1017_d N_A_499_368#_c_533_n 0.00165831f $X=2.955 $Y=1.84 $X2=0 $Y2=0
cc_310 Y N_A_499_368#_c_533_n 0.0159318f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_311 N_Y_c_382_n N_A_27_74#_M1016_s 0.0025999f $X=1.545 $Y=1.095 $X2=0 $Y2=0
cc_312 N_Y_c_384_n N_A_27_74#_M1013_d 0.00250873f $X=2.925 $Y=1.095 $X2=0 $Y2=0
cc_313 N_Y_c_383_n N_A_27_74#_c_592_n 0.00555794f $X=0.875 $Y=1.095 $X2=0 $Y2=0
cc_314 N_Y_M1015_d N_A_27_74#_c_593_n 0.00182874f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_315 N_Y_c_390_n N_A_27_74#_c_593_n 0.0146462f $X=0.71 $Y=0.775 $X2=0 $Y2=0
cc_316 N_Y_c_382_n N_A_27_74#_c_593_n 0.00304353f $X=1.545 $Y=1.095 $X2=0 $Y2=0
cc_317 N_Y_c_382_n N_A_27_74#_c_609_n 0.0194125f $X=1.545 $Y=1.095 $X2=0 $Y2=0
cc_318 N_Y_M1011_s N_A_27_74#_c_595_n 0.0025999f $X=1.5 $Y=0.37 $X2=0 $Y2=0
cc_319 N_Y_c_382_n N_A_27_74#_c_595_n 0.00304353f $X=1.545 $Y=1.095 $X2=0 $Y2=0
cc_320 N_Y_c_413_n N_A_27_74#_c_595_n 0.0180071f $X=1.71 $Y=0.775 $X2=0 $Y2=0
cc_321 N_Y_c_384_n N_A_27_74#_c_595_n 0.00304353f $X=2.925 $Y=1.095 $X2=0 $Y2=0
cc_322 N_Y_c_384_n N_A_27_74#_c_616_n 0.0489623f $X=2.925 $Y=1.095 $X2=0 $Y2=0
cc_323 N_Y_c_384_n N_A_27_74#_c_619_n 0.0208474f $X=2.925 $Y=1.095 $X2=0 $Y2=0
cc_324 N_Y_c_384_n N_A_27_74#_c_597_n 0.0127334f $X=2.925 $Y=1.095 $X2=0 $Y2=0
cc_325 N_Y_c_384_n N_VGND_M1008_d 0.00894066f $X=2.925 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_326 N_VPWR_c_474_n N_A_499_368#_c_533_n 0.0459191f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_327 N_VPWR_c_468_n N_A_499_368#_c_533_n 0.0258001f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_328 N_VPWR_c_474_n N_A_499_368#_c_534_n 0.0179217f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_329 N_VPWR_c_468_n N_A_499_368#_c_534_n 0.00971942f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_330 N_VPWR_c_470_n N_A_499_368#_c_535_n 0.0121617f $X=5 $Y=2.455 $X2=0 $Y2=0
cc_331 N_VPWR_c_474_n N_A_499_368#_c_535_n 0.0644071f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_332 N_VPWR_c_468_n N_A_499_368#_c_535_n 0.0356218f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_333 N_VPWR_c_470_n N_A_499_368#_c_536_n 0.0414289f $X=5 $Y=2.455 $X2=0 $Y2=0
cc_334 N_VPWR_c_474_n N_A_499_368#_c_537_n 0.0121867f $X=4.835 $Y=3.33 $X2=0
+ $Y2=0
cc_335 N_VPWR_c_468_n N_A_499_368#_c_537_n 0.00660921f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_336 N_VPWR_M1006_d N_A_771_368#_c_566_n 0.00666938f $X=4.855 $Y=1.84 $X2=0
+ $Y2=0
cc_337 N_VPWR_c_470_n N_A_771_368#_c_566_n 0.0238156f $X=5 $Y=2.455 $X2=0 $Y2=0
cc_338 N_VPWR_c_470_n N_A_771_368#_c_567_n 0.0267406f $X=5 $Y=2.455 $X2=0 $Y2=0
cc_339 N_VPWR_c_472_n N_A_771_368#_c_567_n 0.0290413f $X=5.955 $Y=2.115 $X2=0
+ $Y2=0
cc_340 N_VPWR_c_475_n N_A_771_368#_c_567_n 0.0146854f $X=5.87 $Y=3.33 $X2=0
+ $Y2=0
cc_341 N_VPWR_c_468_n N_A_771_368#_c_567_n 0.012019f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_342 N_A_499_368#_c_535_n N_A_771_368#_M1000_d 0.00165831f $X=4.275 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_343 N_A_499_368#_M1001_s N_A_771_368#_c_566_n 0.00795918f $X=4.305 $Y=1.84
+ $X2=0 $Y2=0
cc_344 N_A_499_368#_c_536_n N_A_771_368#_c_566_n 0.0219147f $X=4.44 $Y=2.455
+ $X2=0 $Y2=0
cc_345 N_A_499_368#_c_535_n N_A_771_368#_c_570_n 0.0139027f $X=4.275 $Y=2.99
+ $X2=0 $Y2=0
cc_346 N_A_27_74#_c_616_n N_VGND_M1008_d 0.0150186f $X=3.305 $Y=0.755 $X2=-0.19
+ $Y2=-0.245
cc_347 N_A_27_74#_c_596_n N_VGND_M1014_d 0.00251619f $X=4.305 $Y=1.095 $X2=0
+ $Y2=0
cc_348 N_A_27_74#_c_599_n N_VGND_M1007_s 0.0122066f $X=5.795 $Y=1.095 $X2=0
+ $Y2=0
cc_349 N_A_27_74#_c_596_n N_VGND_c_683_n 0.0162019f $X=4.305 $Y=1.095 $X2=0
+ $Y2=0
cc_350 N_A_27_74#_c_598_n N_VGND_c_683_n 0.0169744f $X=4.47 $Y=0.515 $X2=0 $Y2=0
cc_351 N_A_27_74#_c_602_n N_VGND_c_683_n 0.0176756f $X=3.47 $Y=0.515 $X2=0 $Y2=0
cc_352 N_A_27_74#_c_616_n N_VGND_c_684_n 0.0023667f $X=3.305 $Y=0.755 $X2=0
+ $Y2=0
cc_353 N_A_27_74#_c_602_n N_VGND_c_684_n 0.0145639f $X=3.47 $Y=0.515 $X2=0 $Y2=0
cc_354 N_A_27_74#_c_600_n N_VGND_c_686_n 0.0145639f $X=5.96 $Y=0.515 $X2=0 $Y2=0
cc_355 N_A_27_74#_c_593_n N_VGND_c_687_n 0.0241933f $X=1.045 $Y=0.34 $X2=0 $Y2=0
cc_356 N_A_27_74#_c_594_n N_VGND_c_687_n 0.00971942f $X=0.365 $Y=0.34 $X2=0
+ $Y2=0
cc_357 N_A_27_74#_c_595_n N_VGND_c_687_n 0.0365966f $X=2.045 $Y=0.34 $X2=0 $Y2=0
cc_358 N_A_27_74#_c_616_n N_VGND_c_687_n 0.0111582f $X=3.305 $Y=0.755 $X2=0
+ $Y2=0
cc_359 N_A_27_74#_c_598_n N_VGND_c_687_n 0.0119984f $X=4.47 $Y=0.515 $X2=0 $Y2=0
cc_360 N_A_27_74#_c_600_n N_VGND_c_687_n 0.0119984f $X=5.96 $Y=0.515 $X2=0 $Y2=0
cc_361 N_A_27_74#_c_601_n N_VGND_c_687_n 0.0126568f $X=1.21 $Y=0.34 $X2=0 $Y2=0
cc_362 N_A_27_74#_c_602_n N_VGND_c_687_n 0.0119984f $X=3.47 $Y=0.515 $X2=0 $Y2=0
cc_363 N_A_27_74#_c_593_n N_VGND_c_688_n 0.0428729f $X=1.045 $Y=0.34 $X2=0 $Y2=0
cc_364 N_A_27_74#_c_594_n N_VGND_c_688_n 0.0179217f $X=0.365 $Y=0.34 $X2=0 $Y2=0
cc_365 N_A_27_74#_c_595_n N_VGND_c_688_n 0.0656076f $X=2.045 $Y=0.34 $X2=0 $Y2=0
cc_366 N_A_27_74#_c_616_n N_VGND_c_688_n 0.00236055f $X=3.305 $Y=0.755 $X2=0
+ $Y2=0
cc_367 N_A_27_74#_c_601_n N_VGND_c_688_n 0.0232598f $X=1.21 $Y=0.34 $X2=0 $Y2=0
cc_368 N_A_27_74#_c_595_n N_VGND_c_689_n 0.0118583f $X=2.045 $Y=0.34 $X2=0 $Y2=0
cc_369 N_A_27_74#_c_616_n N_VGND_c_689_n 0.0433812f $X=3.305 $Y=0.755 $X2=0
+ $Y2=0
cc_370 N_A_27_74#_c_602_n N_VGND_c_689_n 0.00619249f $X=3.47 $Y=0.515 $X2=0
+ $Y2=0
cc_371 N_A_27_74#_c_598_n N_VGND_c_690_n 0.0145639f $X=4.47 $Y=0.515 $X2=0 $Y2=0
cc_372 N_A_27_74#_c_598_n N_VGND_c_691_n 0.0180018f $X=4.47 $Y=0.515 $X2=0 $Y2=0
cc_373 N_A_27_74#_c_599_n N_VGND_c_691_n 0.0561308f $X=5.795 $Y=1.095 $X2=0
+ $Y2=0
cc_374 N_A_27_74#_c_600_n N_VGND_c_691_n 0.0180018f $X=5.96 $Y=0.515 $X2=0 $Y2=0

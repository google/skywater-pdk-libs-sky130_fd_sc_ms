* File: sky130_fd_sc_ms__o21ai_1.pex.spice
* Created: Wed Sep  2 12:21:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O21AI_1%A1 1 3 6 8 12 15
r30 14 15 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=0.495 $Y=1.385
+ $X2=0.735 $Y2=1.385
r31 11 14 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=0.39 $Y=1.385
+ $X2=0.495 $Y2=1.385
r32 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.39
+ $Y=1.385 $X2=0.39 $Y2=1.385
r33 8 12 4.67207 $w=3.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.24 $Y=1.365
+ $X2=0.39 $Y2=1.365
r34 4 15 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.735 $Y=1.55
+ $X2=0.735 $Y2=1.385
r35 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.735 $Y=1.55
+ $X2=0.735 $Y2=2.4
r36 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.22
+ $X2=0.495 $Y2=1.385
r37 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=1.22 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O21AI_1%A2 3 7 9 15 16
r35 14 16 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=1.23 $Y=1.515
+ $X2=1.405 $Y2=1.515
r36 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.23
+ $Y=1.515 $X2=1.23 $Y2=1.515
r37 11 14 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.155 $Y=1.515
+ $X2=1.23 $Y2=1.515
r38 9 15 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.23 $Y=1.665
+ $X2=1.23 $Y2=1.515
r39 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.35
+ $X2=1.405 $Y2=1.515
r40 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.405 $Y=1.35
+ $X2=1.405 $Y2=0.74
r41 1 11 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=1.68
+ $X2=1.155 $Y2=1.515
r42 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.155 $Y=1.68
+ $X2=1.155 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O21AI_1%B1 3 7 9 10 14
r28 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=1.515
+ $X2=1.885 $Y2=1.68
r29 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=1.515
+ $X2=1.885 $Y2=1.35
r30 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.885
+ $Y=1.515 $X2=1.885 $Y2=1.515
r31 10 15 7.37028 $w=4.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=1.885 $Y2=1.565
r32 9 15 5.4942 $w=4.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.885 $Y2=1.565
r33 7 16 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.835 $Y=0.74
+ $X2=1.835 $Y2=1.35
r34 3 17 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.81 $Y=2.4 $X2=1.81
+ $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O21AI_1%VPWR 1 2 9 13 15 20 21 22 27 36
r25 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r26 33 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r27 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r28 29 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r29 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r30 27 35 4.57341 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=1.87 $Y=3.33
+ $X2=2.135 $Y2=3.33
r31 27 32 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.87 $Y=3.33
+ $X2=1.68 $Y2=3.33
r32 26 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r33 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r34 22 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r35 22 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r36 20 25 4.66471 $w=1.7e-07 $l=6.5e-08 $layer=LI1_cond $X=0.305 $Y=3.33
+ $X2=0.24 $Y2=3.33
r37 20 21 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.305 $Y=3.33
+ $X2=0.43 $Y2=3.33
r38 19 29 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 19 21 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.43 $Y2=3.33
r40 15 18 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=2.035 $Y=2.115
+ $X2=2.035 $Y2=2.815
r41 13 35 3.19276 $w=3.3e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.035 $Y=3.245
+ $X2=2.135 $Y2=3.33
r42 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.035 $Y=3.245
+ $X2=2.035 $Y2=2.815
r43 9 12 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.43 $Y=1.985
+ $X2=0.43 $Y2=2.815
r44 7 21 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.43 $Y=3.245
+ $X2=0.43 $Y2=3.33
r45 7 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.43 $Y=3.245 $X2=0.43
+ $Y2=2.815
r46 2 18 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.9
+ $Y=1.84 $X2=2.035 $Y2=2.815
r47 2 15 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.9
+ $Y=1.84 $X2=2.035 $Y2=2.115
r48 1 12 400 $w=1.7e-07 $l=1.08167e-06 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.84 $X2=0.47 $Y2=2.815
r49 1 9 400 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.84 $X2=0.47 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__O21AI_1%Y 1 2 9 10 13 15 16 20 21
r40 20 21 11.5563 $w=8.18e-07 $l=1.65e-07 $layer=LI1_cond $X=1.135 $Y=2.115
+ $X2=1.135 $Y2=1.95
r41 16 27 0.583453 $w=8.18e-07 $l=4e-08 $layer=LI1_cond $X=1.135 $Y=2.775
+ $X2=1.135 $Y2=2.815
r42 15 16 5.39694 $w=8.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.135 $Y=2.405
+ $X2=1.135 $Y2=2.775
r43 15 20 4.23003 $w=8.18e-07 $l=2.9e-07 $layer=LI1_cond $X=1.135 $Y=2.405
+ $X2=1.135 $Y2=2.115
r44 11 13 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.12 $Y=1.01
+ $X2=2.12 $Y2=0.515
r45 9 11 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.955 $Y=1.095
+ $X2=2.12 $Y2=1.01
r46 9 10 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=1.955 $Y=1.095
+ $X2=0.895 $Y2=1.095
r47 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.81 $Y=1.18
+ $X2=0.895 $Y2=1.095
r48 7 21 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.81 $Y=1.18 $X2=0.81
+ $Y2=1.95
r49 2 27 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.245
+ $Y=1.84 $X2=1.38 $Y2=2.815
r50 2 20 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.245
+ $Y=1.84 $X2=1.38 $Y2=2.115
r51 1 13 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.91
+ $Y=0.37 $X2=2.12 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O21AI_1%A_27_74# 1 2 9 11 12 13
r31 13 15 0.6 $w=3.05e-07 $l=1.5e-08 $layer=LI1_cond $X=1.632 $Y=0.67 $X2=1.632
+ $Y2=0.655
r32 11 13 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=1.48 $Y=0.755
+ $X2=1.632 $Y2=0.67
r33 11 12 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=1.48 $Y=0.755
+ $X2=0.445 $Y2=0.755
r34 7 12 7.55824 $w=1.7e-07 $l=2.16365e-07 $layer=LI1_cond $X=0.267 $Y=0.67
+ $X2=0.445 $Y2=0.755
r35 7 9 5.85668 $w=3.03e-07 $l=1.55e-07 $layer=LI1_cond $X=0.267 $Y=0.67
+ $X2=0.267 $Y2=0.515
r36 2 15 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=1.48
+ $Y=0.37 $X2=1.62 $Y2=0.655
r37 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O21AI_1%VGND 1 4 13 14 19 25
r29 23 25 8.62718 $w=5.83e-07 $l=9.5e-08 $layer=LI1_cond $X=1.2 $Y=0.207
+ $X2=1.295 $Y2=0.207
r30 21 23 1.4312 $w=5.83e-07 $l=7e-08 $layer=LI1_cond $X=1.13 $Y=0.207 $X2=1.2
+ $Y2=0.207
r31 17 21 8.38277 $w=5.83e-07 $l=4.1e-07 $layer=LI1_cond $X=0.72 $Y=0.207
+ $X2=1.13 $Y2=0.207
r32 17 19 9.0361 $w=5.83e-07 $l=1.15e-07 $layer=LI1_cond $X=0.72 $Y=0.207
+ $X2=0.605 $Y2=0.207
r33 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r34 13 25 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=1.295
+ $Y2=0
r35 13 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r36 9 18 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r37 8 19 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=0.605
+ $Y2=0
r38 8 9 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r39 4 14 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r40 4 18 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r41 4 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r42 1 21 91 $w=1.7e-07 $l=5.77235e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=1.13 $Y2=0.335
.ends


* File: sky130_fd_sc_ms__sedfxbp_2.pxi.spice
* Created: Fri Aug 28 18:15:51 2020
* 
x_PM_SKY130_FD_SC_MS__SEDFXBP_2%D N_D_M1027_g N_D_M1001_g D D N_D_c_344_n
+ N_D_c_345_n N_D_c_346_n N_D_c_350_n PM_SKY130_FD_SC_MS__SEDFXBP_2%D
x_PM_SKY130_FD_SC_MS__SEDFXBP_2%A_183_290# N_A_183_290#_M1020_s
+ N_A_183_290#_M1013_s N_A_183_290#_M1003_g N_A_183_290#_M1021_g
+ N_A_183_290#_c_392_n N_A_183_290#_c_384_n N_A_183_290#_c_385_n
+ N_A_183_290#_c_386_n N_A_183_290#_c_387_n N_A_183_290#_c_394_n
+ N_A_183_290#_c_395_n N_A_183_290#_c_388_n N_A_183_290#_c_396_n
+ N_A_183_290#_c_397_n N_A_183_290#_c_389_n N_A_183_290#_c_390_n
+ N_A_183_290#_c_400_n PM_SKY130_FD_SC_MS__SEDFXBP_2%A_183_290#
x_PM_SKY130_FD_SC_MS__SEDFXBP_2%DE N_DE_M1042_g N_DE_c_493_n N_DE_c_494_n
+ N_DE_c_495_n N_DE_c_501_n N_DE_c_496_n N_DE_M1020_g N_DE_c_502_n N_DE_M1013_g
+ N_DE_c_503_n N_DE_c_504_n N_DE_c_505_n N_DE_M1045_g N_DE_c_497_n DE
+ N_DE_c_499_n N_DE_c_500_n PM_SKY130_FD_SC_MS__SEDFXBP_2%DE
x_PM_SKY130_FD_SC_MS__SEDFXBP_2%A_575_87# N_A_575_87#_M1012_d
+ N_A_575_87#_M1044_d N_A_575_87#_M1005_g N_A_575_87#_M1024_g
+ N_A_575_87#_c_582_n N_A_575_87#_M1022_g N_A_575_87#_c_583_n
+ N_A_575_87#_c_584_n N_A_575_87#_M1006_g N_A_575_87#_M1023_g
+ N_A_575_87#_M1002_g N_A_575_87#_M1041_g N_A_575_87#_M1046_g
+ N_A_575_87#_c_605_n N_A_575_87#_c_606_n N_A_575_87#_c_589_n
+ N_A_575_87#_c_608_n N_A_575_87#_c_590_n N_A_575_87#_c_591_n
+ N_A_575_87#_c_717_p N_A_575_87#_c_592_n N_A_575_87#_c_593_n
+ N_A_575_87#_c_594_n N_A_575_87#_c_595_n N_A_575_87#_c_618_n
+ N_A_575_87#_c_596_n N_A_575_87#_c_597_n N_A_575_87#_c_598_n
+ N_A_575_87#_c_599_n N_A_575_87#_c_600_n
+ PM_SKY130_FD_SC_MS__SEDFXBP_2%A_575_87#
x_PM_SKY130_FD_SC_MS__SEDFXBP_2%A_661_87# N_A_661_87#_M1037_s
+ N_A_661_87#_M1014_s N_A_661_87#_c_868_n N_A_661_87#_M1009_g
+ N_A_661_87#_c_869_n N_A_661_87#_c_870_n N_A_661_87#_M1040_g
+ N_A_661_87#_c_871_n N_A_661_87#_c_878_n N_A_661_87#_c_872_n
+ N_A_661_87#_c_888_n N_A_661_87#_c_879_n N_A_661_87#_c_873_n
+ N_A_661_87#_c_880_n N_A_661_87#_c_874_n N_A_661_87#_c_881_n
+ N_A_661_87#_c_875_n N_A_661_87#_c_883_n N_A_661_87#_c_884_n
+ N_A_661_87#_c_876_n PM_SKY130_FD_SC_MS__SEDFXBP_2%A_661_87#
x_PM_SKY130_FD_SC_MS__SEDFXBP_2%SCD N_SCD_M1031_g N_SCD_M1017_g SCD
+ N_SCD_c_979_n PM_SKY130_FD_SC_MS__SEDFXBP_2%SCD
x_PM_SKY130_FD_SC_MS__SEDFXBP_2%SCE N_SCE_c_1024_n N_SCE_M1028_g N_SCE_c_1025_n
+ N_SCE_c_1026_n N_SCE_M1014_g N_SCE_M1037_g N_SCE_c_1019_n N_SCE_c_1020_n
+ N_SCE_M1033_g SCE N_SCE_c_1022_n N_SCE_c_1023_n
+ PM_SKY130_FD_SC_MS__SEDFXBP_2%SCE
x_PM_SKY130_FD_SC_MS__SEDFXBP_2%CLK N_CLK_M1000_g N_CLK_M1029_g CLK
+ N_CLK_c_1094_n N_CLK_c_1095_n PM_SKY130_FD_SC_MS__SEDFXBP_2%CLK
x_PM_SKY130_FD_SC_MS__SEDFXBP_2%A_1586_74# N_A_1586_74#_M1004_d
+ N_A_1586_74#_M1008_d N_A_1586_74#_M1015_g N_A_1586_74#_c_1131_n
+ N_A_1586_74#_M1038_g N_A_1586_74#_M1010_g N_A_1586_74#_M1030_g
+ N_A_1586_74#_c_1134_n N_A_1586_74#_c_1135_n N_A_1586_74#_c_1136_n
+ N_A_1586_74#_c_1157_n N_A_1586_74#_c_1137_n N_A_1586_74#_c_1138_n
+ N_A_1586_74#_c_1139_n N_A_1586_74#_c_1140_n N_A_1586_74#_c_1141_n
+ N_A_1586_74#_c_1237_p N_A_1586_74#_c_1142_n N_A_1586_74#_c_1143_n
+ N_A_1586_74#_c_1144_n N_A_1586_74#_c_1145_n N_A_1586_74#_c_1146_n
+ N_A_1586_74#_c_1147_n N_A_1586_74#_c_1148_n N_A_1586_74#_c_1149_n
+ N_A_1586_74#_c_1159_n N_A_1586_74#_c_1150_n N_A_1586_74#_c_1161_n
+ N_A_1586_74#_c_1151_n N_A_1586_74#_c_1275_p N_A_1586_74#_c_1152_n
+ N_A_1586_74#_c_1153_n N_A_1586_74#_c_1154_n
+ PM_SKY130_FD_SC_MS__SEDFXBP_2%A_1586_74#
x_PM_SKY130_FD_SC_MS__SEDFXBP_2%A_1377_368# N_A_1377_368#_M1029_d
+ N_A_1377_368#_M1000_d N_A_1377_368#_M1004_g N_A_1377_368#_c_1364_n
+ N_A_1377_368#_c_1378_n N_A_1377_368#_M1008_g N_A_1377_368#_c_1365_n
+ N_A_1377_368#_M1035_g N_A_1377_368#_c_1367_n N_A_1377_368#_M1019_g
+ N_A_1377_368#_M1034_g N_A_1377_368#_M1011_g N_A_1377_368#_c_1369_n
+ N_A_1377_368#_c_1370_n N_A_1377_368#_c_1385_n N_A_1377_368#_c_1386_n
+ N_A_1377_368#_c_1387_n N_A_1377_368#_c_1371_n N_A_1377_368#_c_1372_n
+ N_A_1377_368#_c_1389_n N_A_1377_368#_c_1373_n N_A_1377_368#_c_1390_n
+ N_A_1377_368#_c_1391_n N_A_1377_368#_c_1374_n N_A_1377_368#_c_1375_n
+ N_A_1377_368#_c_1376_n N_A_1377_368#_c_1395_n
+ PM_SKY130_FD_SC_MS__SEDFXBP_2%A_1377_368#
x_PM_SKY130_FD_SC_MS__SEDFXBP_2%A_2013_71# N_A_2013_71#_M1018_d
+ N_A_2013_71#_M1032_d N_A_2013_71#_M1025_g N_A_2013_71#_M1016_g
+ N_A_2013_71#_c_1556_n N_A_2013_71#_M1043_g N_A_2013_71#_c_1558_n
+ N_A_2013_71#_M1007_g N_A_2013_71#_c_1559_n N_A_2013_71#_c_1569_n
+ N_A_2013_71#_c_1560_n N_A_2013_71#_c_1561_n N_A_2013_71#_c_1562_n
+ N_A_2013_71#_c_1563_n N_A_2013_71#_c_1564_n N_A_2013_71#_c_1565_n
+ N_A_2013_71#_c_1566_n PM_SKY130_FD_SC_MS__SEDFXBP_2%A_2013_71#
x_PM_SKY130_FD_SC_MS__SEDFXBP_2%A_1784_97# N_A_1784_97#_M1035_d
+ N_A_1784_97#_M1015_d N_A_1784_97#_M1032_g N_A_1784_97#_M1018_g
+ N_A_1784_97#_c_1668_n N_A_1784_97#_c_1671_n N_A_1784_97#_c_1672_n
+ N_A_1784_97#_c_1673_n N_A_1784_97#_c_1674_n N_A_1784_97#_c_1675_n
+ N_A_1784_97#_c_1669_n PM_SKY130_FD_SC_MS__SEDFXBP_2%A_1784_97#
x_PM_SKY130_FD_SC_MS__SEDFXBP_2%A_2489_74# N_A_2489_74#_M1010_d
+ N_A_2489_74#_M1034_d N_A_2489_74#_M1044_g N_A_2489_74#_M1012_g
+ N_A_2489_74#_c_1757_n N_A_2489_74#_M1036_g N_A_2489_74#_M1026_g
+ N_A_2489_74#_M1039_g N_A_2489_74#_M1047_g N_A_2489_74#_c_1762_n
+ N_A_2489_74#_c_1833_n N_A_2489_74#_c_1763_n N_A_2489_74#_c_1764_n
+ N_A_2489_74#_c_1772_n N_A_2489_74#_c_1773_n N_A_2489_74#_c_1774_n
+ N_A_2489_74#_c_1765_n N_A_2489_74#_c_1766_n N_A_2489_74#_c_1767_n
+ N_A_2489_74#_c_1768_n N_A_2489_74#_c_1776_n
+ PM_SKY130_FD_SC_MS__SEDFXBP_2%A_2489_74#
x_PM_SKY130_FD_SC_MS__SEDFXBP_2%A_32_74# N_A_32_74#_M1001_s N_A_32_74#_M1005_d
+ N_A_32_74#_M1027_s N_A_32_74#_M1024_d N_A_32_74#_c_1907_n N_A_32_74#_c_1913_n
+ N_A_32_74#_c_1914_n N_A_32_74#_c_1915_n N_A_32_74#_c_1916_n
+ N_A_32_74#_c_1917_n N_A_32_74#_c_1956_n N_A_32_74#_c_1918_n
+ N_A_32_74#_c_1919_n N_A_32_74#_c_1908_n N_A_32_74#_c_1909_n
+ N_A_32_74#_c_1910_n N_A_32_74#_c_1921_n N_A_32_74#_c_1911_n
+ N_A_32_74#_c_1922_n PM_SKY130_FD_SC_MS__SEDFXBP_2%A_32_74#
x_PM_SKY130_FD_SC_MS__SEDFXBP_2%VPWR N_VPWR_M1003_d N_VPWR_M1013_d
+ N_VPWR_M1014_d N_VPWR_M1000_s N_VPWR_M1008_s N_VPWR_M1016_d N_VPWR_M1043_s
+ N_VPWR_M1006_d N_VPWR_M1036_s N_VPWR_M1039_s N_VPWR_M1046_d N_VPWR_c_2024_n
+ N_VPWR_c_2025_n N_VPWR_c_2026_n N_VPWR_c_2027_n N_VPWR_c_2028_n
+ N_VPWR_c_2029_n N_VPWR_c_2030_n N_VPWR_c_2031_n N_VPWR_c_2032_n
+ N_VPWR_c_2033_n N_VPWR_c_2034_n N_VPWR_c_2035_n N_VPWR_c_2036_n
+ N_VPWR_c_2037_n N_VPWR_c_2038_n N_VPWR_c_2039_n VPWR N_VPWR_c_2040_n
+ N_VPWR_c_2041_n N_VPWR_c_2042_n N_VPWR_c_2043_n N_VPWR_c_2044_n
+ N_VPWR_c_2045_n N_VPWR_c_2046_n N_VPWR_c_2047_n N_VPWR_c_2048_n
+ N_VPWR_c_2049_n N_VPWR_c_2050_n N_VPWR_c_2051_n N_VPWR_c_2052_n
+ N_VPWR_c_2053_n N_VPWR_c_2054_n N_VPWR_c_2055_n N_VPWR_c_2056_n
+ N_VPWR_c_2023_n PM_SKY130_FD_SC_MS__SEDFXBP_2%VPWR
x_PM_SKY130_FD_SC_MS__SEDFXBP_2%A_691_113# N_A_691_113#_M1009_d
+ N_A_691_113#_M1033_d N_A_691_113#_M1035_s N_A_691_113#_M1028_d
+ N_A_691_113#_M1040_d N_A_691_113#_M1015_s N_A_691_113#_c_2231_n
+ N_A_691_113#_c_2294_n N_A_691_113#_c_2232_n N_A_691_113#_c_2243_n
+ N_A_691_113#_c_2259_n N_A_691_113#_c_2233_n N_A_691_113#_c_2234_n
+ N_A_691_113#_c_2223_n N_A_691_113#_c_2224_n N_A_691_113#_c_2236_n
+ N_A_691_113#_c_2237_n N_A_691_113#_c_2238_n N_A_691_113#_c_2225_n
+ N_A_691_113#_c_2226_n N_A_691_113#_c_2252_n N_A_691_113#_c_2227_n
+ N_A_691_113#_c_2239_n N_A_691_113#_c_2240_n N_A_691_113#_c_2228_n
+ N_A_691_113#_c_2229_n N_A_691_113#_c_2230_n N_A_691_113#_c_2390_n
+ N_A_691_113#_c_2329_n PM_SKY130_FD_SC_MS__SEDFXBP_2%A_691_113#
x_PM_SKY130_FD_SC_MS__SEDFXBP_2%Q N_Q_M1026_d N_Q_M1036_d Q Q Q Q Q
+ PM_SKY130_FD_SC_MS__SEDFXBP_2%Q
x_PM_SKY130_FD_SC_MS__SEDFXBP_2%Q_N N_Q_N_M1023_d N_Q_N_M1002_s N_Q_N_c_2428_n
+ N_Q_N_c_2429_n Q_N Q_N Q_N Q_N Q_N Q_N Q_N PM_SKY130_FD_SC_MS__SEDFXBP_2%Q_N
x_PM_SKY130_FD_SC_MS__SEDFXBP_2%VGND N_VGND_M1042_d N_VGND_M1020_d
+ N_VGND_M1037_d N_VGND_M1029_s N_VGND_M1004_s N_VGND_M1025_d N_VGND_M1007_s
+ N_VGND_M1022_d N_VGND_M1026_s N_VGND_M1047_s N_VGND_M1041_s N_VGND_c_2461_n
+ N_VGND_c_2462_n N_VGND_c_2463_n N_VGND_c_2464_n N_VGND_c_2465_n
+ N_VGND_c_2466_n N_VGND_c_2467_n N_VGND_c_2468_n N_VGND_c_2469_n
+ N_VGND_c_2470_n N_VGND_c_2471_n N_VGND_c_2472_n N_VGND_c_2473_n
+ N_VGND_c_2474_n N_VGND_c_2475_n N_VGND_c_2476_n N_VGND_c_2477_n
+ N_VGND_c_2478_n N_VGND_c_2479_n N_VGND_c_2480_n N_VGND_c_2481_n VGND
+ N_VGND_c_2482_n N_VGND_c_2483_n N_VGND_c_2484_n N_VGND_c_2485_n
+ N_VGND_c_2486_n N_VGND_c_2487_n N_VGND_c_2488_n N_VGND_c_2489_n
+ N_VGND_c_2490_n N_VGND_c_2491_n N_VGND_c_2492_n N_VGND_c_2493_n
+ N_VGND_c_2494_n N_VGND_c_2495_n N_VGND_c_2496_n
+ PM_SKY130_FD_SC_MS__SEDFXBP_2%VGND
cc_1 VNB N_D_M1001_g 0.0264128f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.58
cc_2 VNB N_D_c_344_n 0.0166671f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_3 VNB N_D_c_345_n 0.0120671f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_4 VNB N_D_c_346_n 0.0398527f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.825
cc_5 VNB N_A_183_290#_M1021_g 0.0449705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_183_290#_c_384_n 0.00295485f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.825
cc_7 VNB N_A_183_290#_c_385_n 0.0231869f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.825
cc_8 VNB N_A_183_290#_c_386_n 0.0073121f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.99
cc_9 VNB N_A_183_290#_c_387_n 4.59932e-19 $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.145
cc_10 VNB N_A_183_290#_c_388_n 0.00999719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_183_290#_c_389_n 0.00268811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_183_290#_c_390_n 0.0162115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_DE_M1042_g 0.0299417f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.64
cc_14 VNB N_DE_c_493_n 0.0304597f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.98
cc_15 VNB N_DE_c_494_n 0.00725655f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.58
cc_16 VNB N_DE_c_495_n 0.0266857f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_17 VNB N_DE_c_496_n 0.0179672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_DE_c_497_n 0.00950241f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB DE 0.0038178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_DE_c_499_n 0.0165295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_DE_c_500_n 0.0196098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_575_87#_M1005_g 0.0399729f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_23 VNB N_A_575_87#_c_582_n 0.0170882f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.825
cc_24 VNB N_A_575_87#_c_583_n 0.0400986f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_25 VNB N_A_575_87#_c_584_n 0.00716283f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.825
cc_26 VNB N_A_575_87#_M1023_g 0.0215195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_575_87#_M1002_g 0.0013098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_575_87#_M1041_g 0.023699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_575_87#_M1046_g 0.00169511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_575_87#_c_589_n 5.3143e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_575_87#_c_590_n 0.00811762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_575_87#_c_591_n 0.00364338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_575_87#_c_592_n 9.39012e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_575_87#_c_593_n 0.00301273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_575_87#_c_594_n 0.01027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_575_87#_c_595_n 0.0465057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_575_87#_c_596_n 2.4907e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_575_87#_c_597_n 0.00101108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_575_87#_c_598_n 0.01914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_575_87#_c_599_n 0.0335071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_575_87#_c_600_n 0.0425155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_661_87#_c_868_n 0.0164494f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.58
cc_43 VNB N_A_661_87#_c_869_n 0.0374808f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.98
cc_44 VNB N_A_661_87#_c_870_n 0.00865069f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_45 VNB N_A_661_87#_c_871_n 0.00880625f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_46 VNB N_A_661_87#_c_872_n 0.00219983f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.825
cc_47 VNB N_A_661_87#_c_873_n 0.00716145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_661_87#_c_874_n 0.0680445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_661_87#_c_875_n 0.0346451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_661_87#_c_876_n 0.032224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_SCD_M1031_g 0.00875717f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.64
cc_52 VNB N_SCD_M1017_g 0.0175076f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.58
cc_53 VNB SCD 0.0142331f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_54 VNB N_SCD_c_979_n 0.0311734f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_55 VNB N_SCE_M1014_g 0.00875383f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_56 VNB N_SCE_M1037_g 0.0334855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_SCE_c_1019_n 0.0681329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_SCE_c_1020_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.825
cc_59 VNB N_SCE_M1033_g 0.0359126f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_60 VNB N_SCE_c_1022_n 0.027336f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.145
cc_61 VNB N_SCE_c_1023_n 0.0059654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_CLK_M1000_g 0.00709984f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.64
cc_63 VNB CLK 0.00807833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_CLK_c_1094_n 0.037862f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_65 VNB N_CLK_c_1095_n 0.0212689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1586_74#_c_1131_n 0.0185214f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_67 VNB N_A_1586_74#_M1010_g 0.035432f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_68 VNB N_A_1586_74#_M1030_g 0.00537699f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.825
cc_69 VNB N_A_1586_74#_c_1134_n 0.00958186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1586_74#_c_1135_n 0.0189124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1586_74#_c_1136_n 0.00279267f $X=-0.19 $Y=-0.245 $X2=0.63
+ $Y2=1.665
cc_72 VNB N_A_1586_74#_c_1137_n 0.017477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1586_74#_c_1138_n 5.87492e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1586_74#_c_1139_n 0.0022144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1586_74#_c_1140_n 0.0434353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1586_74#_c_1141_n 0.0082121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1586_74#_c_1142_n 0.00904398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1586_74#_c_1143_n 0.00203028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1586_74#_c_1144_n 0.00953978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1586_74#_c_1145_n 0.00466954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1586_74#_c_1146_n 0.00313816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1586_74#_c_1147_n 0.00318285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1586_74#_c_1148_n 0.00302573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1586_74#_c_1149_n 0.0116019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1586_74#_c_1150_n 0.00571213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1586_74#_c_1151_n 0.00123754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1586_74#_c_1152_n 0.00280784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1586_74#_c_1153_n 0.0296806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1586_74#_c_1154_n 0.0174662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1377_368#_M1004_g 0.0392551f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_91 VNB N_A_1377_368#_c_1364_n 0.00338077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1377_368#_c_1365_n 0.0154568f $X=-0.19 $Y=-0.245 $X2=0.54
+ $Y2=1.145
cc_93 VNB N_A_1377_368#_M1035_g 0.053968f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.99
cc_94 VNB N_A_1377_368#_c_1367_n 0.0309731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1377_368#_M1011_g 0.0511607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1377_368#_c_1369_n 0.00656975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1377_368#_c_1370_n 0.00119395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1377_368#_c_1371_n 0.0123224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1377_368#_c_1372_n 0.010047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1377_368#_c_1373_n 0.00894163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1377_368#_c_1374_n 0.00381838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1377_368#_c_1375_n 0.0151412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1377_368#_c_1376_n 0.033009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_2013_71#_M1025_g 0.030024f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_105 VNB N_A_2013_71#_M1016_g 0.00884039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_2013_71#_c_1556_n 0.0300468f $X=-0.19 $Y=-0.245 $X2=0.54
+ $Y2=1.145
cc_107 VNB N_A_2013_71#_M1043_g 0.0086274f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.825
cc_108 VNB N_A_2013_71#_c_1558_n 0.0198235f $X=-0.19 $Y=-0.245 $X2=0.54
+ $Y2=1.825
cc_109 VNB N_A_2013_71#_c_1559_n 0.00999316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_2013_71#_c_1560_n 0.00548308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_2013_71#_c_1561_n 0.00253632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_2013_71#_c_1562_n 0.00496828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_2013_71#_c_1563_n 0.00184523f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_2013_71#_c_1564_n 0.0564399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_2013_71#_c_1565_n 0.00274233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_2013_71#_c_1566_n 0.0364327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_1784_97#_M1018_g 0.0420339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_1784_97#_c_1668_n 0.013135f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_119 VNB N_A_1784_97#_c_1669_n 0.0192949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_2489_74#_M1044_g 0.00206851f $X=-0.19 $Y=-0.245 $X2=0.54
+ $Y2=1.145
cc_121 VNB N_A_2489_74#_M1012_g 0.0257653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_2489_74#_c_1757_n 0.0701032f $X=-0.19 $Y=-0.245 $X2=0.54
+ $Y2=1.825
cc_123 VNB N_A_2489_74#_M1036_g 0.00151236f $X=-0.19 $Y=-0.245 $X2=0.54
+ $Y2=1.825
cc_124 VNB N_A_2489_74#_M1026_g 0.022963f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.145
cc_125 VNB N_A_2489_74#_M1039_g 0.00139073f $X=-0.19 $Y=-0.245 $X2=0.63
+ $Y2=1.665
cc_126 VNB N_A_2489_74#_M1047_g 0.0208419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_A_2489_74#_c_1762_n 0.0346105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_2489_74#_c_1763_n 0.00286498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_A_2489_74#_c_1764_n 0.00321929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_A_2489_74#_c_1765_n 0.00525878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_A_2489_74#_c_1766_n 0.00283454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_A_2489_74#_c_1767_n 0.0083479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_A_2489_74#_c_1768_n 0.0288173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_A_32_74#_c_1907_n 0.0434942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_A_32_74#_c_1908_n 0.00382371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_A_32_74#_c_1909_n 0.00641878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_A_32_74#_c_1910_n 0.0138478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_A_32_74#_c_1911_n 0.00433514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VPWR_c_2023_n 0.720949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_A_691_113#_c_2223_n 0.0105451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_A_691_113#_c_2224_n 0.0100696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_A_691_113#_c_2225_n 0.0104521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_A_691_113#_c_2226_n 0.00181722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_A_691_113#_c_2227_n 0.0173316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_A_691_113#_c_2228_n 0.00973194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_A_691_113#_c_2229_n 0.00794098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_A_691_113#_c_2230_n 0.0192996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB Q 0.00240191f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.58
cc_149 VNB N_Q_N_c_2428_n 0.0132008f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=0.58
cc_150 VNB N_Q_N_c_2429_n 0.0239423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB Q_N 0.00239713f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.145
cc_152 VNB N_VGND_c_2461_n 0.0193314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2462_n 0.0301467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2463_n 0.0105113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2464_n 0.0172622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2465_n 0.00978559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_2466_n 0.0106328f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2467_n 0.00590394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_2468_n 0.0119255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_2469_n 0.00982717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_VGND_c_2470_n 0.00206318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VNB N_VGND_c_2471_n 0.0206041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_VGND_c_2472_n 0.0192796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VNB N_VGND_c_2473_n 0.0192531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_VGND_c_2474_n 0.00984545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_VGND_c_2475_n 0.0124653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_VGND_c_2476_n 0.0280494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_VGND_c_2477_n 0.023012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_169 VNB N_VGND_c_2478_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_170 VNB N_VGND_c_2479_n 0.0220562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_VGND_c_2480_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_172 VNB N_VGND_c_2481_n 0.0403351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_173 VNB N_VGND_c_2482_n 0.032665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_174 VNB N_VGND_c_2483_n 0.0688863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_175 VNB N_VGND_c_2484_n 0.0331395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_176 VNB N_VGND_c_2485_n 0.0636008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_177 VNB N_VGND_c_2486_n 0.0296519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_178 VNB N_VGND_c_2487_n 0.019013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_179 VNB N_VGND_c_2488_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_180 VNB N_VGND_c_2489_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_181 VNB N_VGND_c_2490_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_182 VNB N_VGND_c_2491_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_183 VNB N_VGND_c_2492_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_184 VNB N_VGND_c_2493_n 0.0112842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_185 VNB N_VGND_c_2494_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_186 VNB N_VGND_c_2495_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_187 VNB N_VGND_c_2496_n 0.938824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_188 VPB N_D_M1027_g 0.0364358f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=2.64
cc_189 VPB N_D_c_345_n 0.00461728f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.145
cc_190 VPB N_D_c_346_n 0.0112765f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_191 VPB N_D_c_350_n 0.0156268f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.99
cc_192 VPB N_A_183_290#_M1003_g 0.0284703f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.145
cc_193 VPB N_A_183_290#_c_392_n 0.0239716f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.145
cc_194 VPB N_A_183_290#_c_385_n 0.020582f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_195 VPB N_A_183_290#_c_394_n 0.0113728f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_183_290#_c_395_n 0.00225372f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.295
cc_197 VPB N_A_183_290#_c_396_n 0.0026814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_183_290#_c_397_n 0.0123271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_183_290#_c_389_n 0.00274132f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_183_290#_c_390_n 0.0179737f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_183_290#_c_400_n 0.00136575f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_DE_c_501_n 0.0193526f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_203 VPB N_DE_c_502_n 0.0183667f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.145
cc_204 VPB N_DE_c_503_n 0.0399818f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_205 VPB N_DE_c_504_n 0.0299518f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_206 VPB N_DE_c_505_n 0.0161934f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_207 VPB DE 0.0020259f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_DE_c_499_n 0.0123229f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_575_87#_M1024_g 0.0420777f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_575_87#_M1006_g 0.0235439f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.99
cc_211 VPB N_A_575_87#_M1002_g 0.0220571f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_575_87#_M1046_g 0.0257045f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_A_575_87#_c_605_n 0.0059015f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_575_87#_c_606_n 0.0303245f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_575_87#_c_589_n 0.015414f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_575_87#_c_608_n 0.00860613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_575_87#_c_592_n 0.00293318f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_575_87#_c_595_n 0.0554236f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_575_87#_c_596_n 0.00131138f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_575_87#_c_597_n 0.00129194f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_575_87#_c_598_n 0.0226993f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_575_87#_c_599_n 0.0226425f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_661_87#_M1040_g 0.0249271f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_661_87#_c_878_n 0.0278493f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_225 VPB N_A_661_87#_c_879_n 0.00433316f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.665
cc_226 VPB N_A_661_87#_c_880_n 0.0208166f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_661_87#_c_881_n 0.00321747f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_A_661_87#_c_875_n 0.0418704f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_661_87#_c_883_n 0.00982317f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_661_87#_c_884_n 0.00242577f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_661_87#_c_876_n 0.0173302f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_SCD_M1031_g 0.048286f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=2.64
cc_233 VPB N_SCE_c_1024_n 0.0204383f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.99
cc_234 VPB N_SCE_c_1025_n 0.0742449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_SCE_c_1026_n 0.0134074f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=0.98
cc_236 VPB N_SCE_M1014_g 0.0454819f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.145
cc_237 VPB N_CLK_M1000_g 0.0301874f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=2.64
cc_238 VPB N_A_1586_74#_M1015_g 0.0305862f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.145
cc_239 VPB N_A_1586_74#_M1030_g 0.0596692f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_240 VPB N_A_1586_74#_c_1157_n 0.00485351f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_A_1586_74#_c_1148_n 0.00648383f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_A_1586_74#_c_1159_n 0.0050371f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_A_1586_74#_c_1150_n 0.00177748f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_A_1586_74#_c_1161_n 0.0497984f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_A_1586_74#_c_1154_n 0.0189353f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_A_1377_368#_c_1364_n 0.00340931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_A_1377_368#_c_1378_n 0.0253459f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_248 VPB N_A_1377_368#_c_1365_n 0.0166204f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.145
cc_249 VPB N_A_1377_368#_c_1367_n 0.0173878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_A_1377_368#_M1019_g 0.0239851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_A_1377_368#_M1034_g 0.0286145f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_A_1377_368#_c_1369_n 0.00143274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_A_1377_368#_c_1370_n 0.00298346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_A_1377_368#_c_1385_n 0.00395733f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_A_1377_368#_c_1386_n 0.0121562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_A_1377_368#_c_1387_n 0.00260289f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_A_1377_368#_c_1372_n 0.00680749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_A_1377_368#_c_1389_n 0.0403178f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_A_1377_368#_c_1390_n 0.00755953f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_A_1377_368#_c_1391_n 0.0301553f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_A_1377_368#_c_1374_n 0.00210725f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_A_1377_368#_c_1375_n 0.0157621f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_A_1377_368#_c_1376_n 0.0123378f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_A_1377_368#_c_1395_n 0.0180856f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_A_2013_71#_M1016_g 0.0649216f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_A_2013_71#_M1043_g 0.0385568f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_267 VPB N_A_2013_71#_c_1569_n 0.00602683f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_A_2013_71#_c_1561_n 0.00900558f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_A_1784_97#_M1032_g 0.0250206f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.145
cc_270 VPB N_A_1784_97#_c_1671_n 0.0162618f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_271 VPB N_A_1784_97#_c_1672_n 0.00117381f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.145
cc_272 VPB N_A_1784_97#_c_1673_n 0.00454891f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.295
cc_273 VPB N_A_1784_97#_c_1674_n 0.00721179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_A_1784_97#_c_1675_n 0.0017703f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.825
cc_275 VPB N_A_1784_97#_c_1669_n 0.0195927f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_A_2489_74#_M1044_g 0.0282104f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.145
cc_277 VPB N_A_2489_74#_M1036_g 0.0239827f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_278 VPB N_A_2489_74#_M1039_g 0.0213437f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.665
cc_279 VPB N_A_2489_74#_c_1772_n 0.00586333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_280 VPB N_A_2489_74#_c_1773_n 0.0110034f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_281 VPB N_A_2489_74#_c_1774_n 0.0015169f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_A_2489_74#_c_1766_n 0.0014512f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_283 VPB N_A_2489_74#_c_1776_n 0.0043814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_284 VPB N_A_32_74#_c_1907_n 0.0303354f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_285 VPB N_A_32_74#_c_1913_n 0.0260862f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.145
cc_286 VPB N_A_32_74#_c_1914_n 0.0153562f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_287 VPB N_A_32_74#_c_1915_n 0.00991141f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.99
cc_288 VPB N_A_32_74#_c_1916_n 0.00911955f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.145
cc_289 VPB N_A_32_74#_c_1917_n 0.00348146f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_290 VPB N_A_32_74#_c_1918_n 0.00680986f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.665
cc_291 VPB N_A_32_74#_c_1919_n 9.33339e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_292 VPB N_A_32_74#_c_1909_n 0.0122383f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_293 VPB N_A_32_74#_c_1921_n 0.0139437f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_294 VPB N_A_32_74#_c_1922_n 0.00404895f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_295 VPB N_VPWR_c_2024_n 0.00585142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_296 VPB N_VPWR_c_2025_n 0.00572224f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_297 VPB N_VPWR_c_2026_n 0.00806049f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_298 VPB N_VPWR_c_2027_n 0.00734079f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_299 VPB N_VPWR_c_2028_n 0.0218871f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_300 VPB N_VPWR_c_2029_n 0.0114049f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_301 VPB N_VPWR_c_2030_n 0.016189f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_302 VPB N_VPWR_c_2031_n 0.00864425f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_303 VPB N_VPWR_c_2032_n 0.0089741f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_304 VPB N_VPWR_c_2033_n 0.00261791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_305 VPB N_VPWR_c_2034_n 0.0119967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_306 VPB N_VPWR_c_2035_n 0.0403893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_307 VPB N_VPWR_c_2036_n 0.0342477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_308 VPB N_VPWR_c_2037_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_309 VPB N_VPWR_c_2038_n 0.0242802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_310 VPB N_VPWR_c_2039_n 0.00632182f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_311 VPB N_VPWR_c_2040_n 0.0324541f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_312 VPB N_VPWR_c_2041_n 0.0296421f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_313 VPB N_VPWR_c_2042_n 0.0590043f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_314 VPB N_VPWR_c_2043_n 0.0335097f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_315 VPB N_VPWR_c_2044_n 0.059622f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_316 VPB N_VPWR_c_2045_n 0.0636904f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_317 VPB N_VPWR_c_2046_n 0.0203698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_318 VPB N_VPWR_c_2047_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_319 VPB N_VPWR_c_2048_n 0.01587f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_320 VPB N_VPWR_c_2049_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_321 VPB N_VPWR_c_2050_n 0.00466629f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_322 VPB N_VPWR_c_2051_n 0.00516749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_323 VPB N_VPWR_c_2052_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_324 VPB N_VPWR_c_2053_n 0.00613689f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_325 VPB N_VPWR_c_2054_n 0.0101667f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_326 VPB N_VPWR_c_2055_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_327 VPB N_VPWR_c_2056_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_328 VPB N_VPWR_c_2023_n 0.203348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_329 VPB N_A_691_113#_c_2231_n 0.00173654f $X=-0.19 $Y=1.66 $X2=0.54 $Y2=1.825
cc_330 VPB N_A_691_113#_c_2232_n 0.0114257f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.295
cc_331 VPB N_A_691_113#_c_2233_n 0.00777695f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.825
cc_332 VPB N_A_691_113#_c_2234_n 0.00122302f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_333 VPB N_A_691_113#_c_2224_n 0.0091361f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_334 VPB N_A_691_113#_c_2236_n 0.020222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_335 VPB N_A_691_113#_c_2237_n 0.0201404f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_336 VPB N_A_691_113#_c_2238_n 0.00161506f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_337 VPB N_A_691_113#_c_2239_n 0.00985592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_338 VPB N_A_691_113#_c_2240_n 0.00716663f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_339 VPB N_A_691_113#_c_2229_n 0.0099146f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_340 VPB N_Q_N_c_2429_n 0.0183485f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_341 VPB Q_N 0.00281594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_342 N_D_M1027_g N_A_183_290#_c_392_n 0.0593694f $X=0.585 $Y=2.64 $X2=0 $Y2=0
cc_343 N_D_c_350_n N_A_183_290#_c_392_n 0.0169614f $X=0.54 $Y=1.99 $X2=0 $Y2=0
cc_344 N_D_c_345_n N_A_183_290#_c_384_n 0.0545333f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_345 N_D_c_346_n N_A_183_290#_c_384_n 0.00133474f $X=0.54 $Y=1.825 $X2=0 $Y2=0
cc_346 N_D_c_345_n N_A_183_290#_c_385_n 0.00384651f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_347 N_D_c_346_n N_A_183_290#_c_385_n 0.0169614f $X=0.54 $Y=1.825 $X2=0 $Y2=0
cc_348 N_D_c_345_n N_A_183_290#_c_387_n 0.0148197f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_349 N_D_c_346_n N_A_183_290#_c_387_n 4.03978e-19 $X=0.54 $Y=1.825 $X2=0 $Y2=0
cc_350 N_D_M1027_g N_A_183_290#_c_395_n 6.9419e-19 $X=0.585 $Y=2.64 $X2=0 $Y2=0
cc_351 N_D_c_345_n N_A_183_290#_c_395_n 0.00341199f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_352 N_D_M1001_g N_DE_M1042_g 0.025244f $X=0.63 $Y=0.58 $X2=0 $Y2=0
cc_353 N_D_c_345_n N_DE_M1042_g 0.00420913f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_354 N_D_c_344_n N_DE_c_494_n 0.025244f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_355 N_D_M1027_g N_A_32_74#_c_1907_n 0.00969435f $X=0.585 $Y=2.64 $X2=0 $Y2=0
cc_356 N_D_M1001_g N_A_32_74#_c_1907_n 0.00669921f $X=0.63 $Y=0.58 $X2=0 $Y2=0
cc_357 N_D_c_344_n N_A_32_74#_c_1907_n 0.0239763f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_358 N_D_c_345_n N_A_32_74#_c_1907_n 0.0771054f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_359 N_D_M1027_g N_A_32_74#_c_1913_n 0.0104235f $X=0.585 $Y=2.64 $X2=0 $Y2=0
cc_360 N_D_M1027_g N_A_32_74#_c_1914_n 0.013196f $X=0.585 $Y=2.64 $X2=0 $Y2=0
cc_361 N_D_c_345_n N_A_32_74#_c_1914_n 0.0161175f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_362 N_D_M1001_g N_A_32_74#_c_1910_n 0.0058515f $X=0.63 $Y=0.58 $X2=0 $Y2=0
cc_363 N_D_c_344_n N_A_32_74#_c_1910_n 0.00276862f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_364 N_D_c_345_n N_A_32_74#_c_1910_n 0.00757623f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_365 N_D_M1027_g N_A_32_74#_c_1921_n 0.00166609f $X=0.585 $Y=2.64 $X2=0 $Y2=0
cc_366 N_D_c_345_n N_A_32_74#_c_1921_n 0.00562948f $X=0.54 $Y=1.145 $X2=0 $Y2=0
cc_367 N_D_c_350_n N_A_32_74#_c_1921_n 0.00263932f $X=0.54 $Y=1.99 $X2=0 $Y2=0
cc_368 N_D_M1027_g N_VPWR_c_2024_n 0.00153898f $X=0.585 $Y=2.64 $X2=0 $Y2=0
cc_369 N_D_M1027_g N_VPWR_c_2040_n 0.005209f $X=0.585 $Y=2.64 $X2=0 $Y2=0
cc_370 N_D_M1027_g N_VPWR_c_2023_n 0.0098717f $X=0.585 $Y=2.64 $X2=0 $Y2=0
cc_371 N_D_M1001_g N_VGND_c_2461_n 0.00218592f $X=0.63 $Y=0.58 $X2=0 $Y2=0
cc_372 N_D_M1001_g N_VGND_c_2482_n 0.004347f $X=0.63 $Y=0.58 $X2=0 $Y2=0
cc_373 N_D_M1001_g N_VGND_c_2496_n 0.00822933f $X=0.63 $Y=0.58 $X2=0 $Y2=0
cc_374 N_A_183_290#_c_388_n N_DE_M1042_g 0.00659112f $X=1.845 $Y=0.775 $X2=0
+ $Y2=0
cc_375 N_A_183_290#_c_386_n N_DE_c_493_n 0.0130203f $X=1.68 $Y=1.195 $X2=0 $Y2=0
cc_376 N_A_183_290#_c_387_n N_DE_c_493_n 0.00791665f $X=1.335 $Y=1.195 $X2=0
+ $Y2=0
cc_377 N_A_183_290#_c_385_n N_DE_c_494_n 0.0226593f $X=1.17 $Y=1.615 $X2=0 $Y2=0
cc_378 N_A_183_290#_c_387_n N_DE_c_494_n 0.00629125f $X=1.335 $Y=1.195 $X2=0
+ $Y2=0
cc_379 N_A_183_290#_c_386_n N_DE_c_495_n 0.00690186f $X=1.68 $Y=1.195 $X2=0
+ $Y2=0
cc_380 N_A_183_290#_c_388_n N_DE_c_495_n 0.00596863f $X=1.845 $Y=0.775 $X2=0
+ $Y2=0
cc_381 N_A_183_290#_c_384_n N_DE_c_501_n 9.54411e-19 $X=1.17 $Y=1.615 $X2=0
+ $Y2=0
cc_382 N_A_183_290#_c_385_n N_DE_c_501_n 0.00491474f $X=1.17 $Y=1.615 $X2=0
+ $Y2=0
cc_383 N_A_183_290#_c_394_n N_DE_c_501_n 0.00391046f $X=1.825 $Y=2.035 $X2=0
+ $Y2=0
cc_384 N_A_183_290#_c_389_n N_DE_c_501_n 0.00303743f $X=2.47 $Y=1.68 $X2=0 $Y2=0
cc_385 N_A_183_290#_c_400_n N_DE_c_501_n 0.00539719f $X=1.91 $Y=2.035 $X2=0
+ $Y2=0
cc_386 N_A_183_290#_M1021_g N_DE_c_496_n 0.0184318f $X=2.56 $Y=0.775 $X2=0 $Y2=0
cc_387 N_A_183_290#_c_388_n N_DE_c_496_n 0.00860606f $X=1.845 $Y=0.775 $X2=0
+ $Y2=0
cc_388 N_A_183_290#_c_396_n N_DE_c_502_n 0.00332874f $X=1.91 $Y=2.51 $X2=0 $Y2=0
cc_389 N_A_183_290#_c_397_n N_DE_c_503_n 0.0105094f $X=2.305 $Y=2.035 $X2=0
+ $Y2=0
cc_390 N_A_183_290#_c_390_n N_DE_c_503_n 0.0181303f $X=2.47 $Y=1.68 $X2=0 $Y2=0
cc_391 N_A_183_290#_M1003_g N_DE_c_504_n 0.00302257f $X=1.005 $Y=2.64 $X2=0
+ $Y2=0
cc_392 N_A_183_290#_c_392_n N_DE_c_504_n 0.00491474f $X=1.125 $Y=2.12 $X2=0
+ $Y2=0
cc_393 N_A_183_290#_c_394_n N_DE_c_504_n 0.00339243f $X=1.825 $Y=2.035 $X2=0
+ $Y2=0
cc_394 N_A_183_290#_c_396_n N_DE_c_504_n 0.0148926f $X=1.91 $Y=2.51 $X2=0 $Y2=0
cc_395 N_A_183_290#_c_397_n N_DE_c_504_n 0.0126169f $X=2.305 $Y=2.035 $X2=0
+ $Y2=0
cc_396 N_A_183_290#_c_400_n N_DE_c_504_n 0.00209363f $X=1.91 $Y=2.035 $X2=0
+ $Y2=0
cc_397 N_A_183_290#_c_386_n N_DE_c_497_n 0.00525481f $X=1.68 $Y=1.195 $X2=0
+ $Y2=0
cc_398 N_A_183_290#_c_388_n N_DE_c_497_n 0.00353956f $X=1.845 $Y=0.775 $X2=0
+ $Y2=0
cc_399 N_A_183_290#_M1021_g DE 3.21021e-19 $X=2.56 $Y=0.775 $X2=0 $Y2=0
cc_400 N_A_183_290#_c_384_n DE 0.020843f $X=1.17 $Y=1.615 $X2=0 $Y2=0
cc_401 N_A_183_290#_c_385_n DE 0.00206473f $X=1.17 $Y=1.615 $X2=0 $Y2=0
cc_402 N_A_183_290#_c_386_n DE 0.0270293f $X=1.68 $Y=1.195 $X2=0 $Y2=0
cc_403 N_A_183_290#_c_394_n DE 0.019286f $X=1.825 $Y=2.035 $X2=0 $Y2=0
cc_404 N_A_183_290#_c_389_n DE 0.00999033f $X=2.47 $Y=1.68 $X2=0 $Y2=0
cc_405 N_A_183_290#_c_390_n DE 0.00111448f $X=2.47 $Y=1.68 $X2=0 $Y2=0
cc_406 N_A_183_290#_c_400_n DE 0.00638598f $X=1.91 $Y=2.035 $X2=0 $Y2=0
cc_407 N_A_183_290#_M1021_g N_DE_c_499_n 9.94929e-19 $X=2.56 $Y=0.775 $X2=0
+ $Y2=0
cc_408 N_A_183_290#_c_384_n N_DE_c_499_n 4.11485e-19 $X=1.17 $Y=1.615 $X2=0
+ $Y2=0
cc_409 N_A_183_290#_c_385_n N_DE_c_499_n 0.0179198f $X=1.17 $Y=1.615 $X2=0 $Y2=0
cc_410 N_A_183_290#_c_386_n N_DE_c_499_n 0.00127783f $X=1.68 $Y=1.195 $X2=0
+ $Y2=0
cc_411 N_A_183_290#_c_394_n N_DE_c_499_n 0.00462669f $X=1.825 $Y=2.035 $X2=0
+ $Y2=0
cc_412 N_A_183_290#_c_389_n N_DE_c_499_n 7.04955e-19 $X=2.47 $Y=1.68 $X2=0 $Y2=0
cc_413 N_A_183_290#_c_390_n N_DE_c_499_n 0.00950624f $X=2.47 $Y=1.68 $X2=0 $Y2=0
cc_414 N_A_183_290#_c_384_n N_DE_c_500_n 0.00581511f $X=1.17 $Y=1.615 $X2=0
+ $Y2=0
cc_415 N_A_183_290#_c_386_n N_DE_c_500_n 0.00597544f $X=1.68 $Y=1.195 $X2=0
+ $Y2=0
cc_416 N_A_183_290#_M1021_g N_A_575_87#_M1005_g 0.0369397f $X=2.56 $Y=0.775
+ $X2=0 $Y2=0
cc_417 N_A_183_290#_c_397_n N_A_575_87#_M1024_g 0.00421101f $X=2.305 $Y=2.035
+ $X2=0 $Y2=0
cc_418 N_A_183_290#_c_389_n N_A_575_87#_M1024_g 0.00283945f $X=2.47 $Y=1.68
+ $X2=0 $Y2=0
cc_419 N_A_183_290#_c_389_n N_A_575_87#_c_618_n 0.00127953f $X=2.47 $Y=1.68
+ $X2=0 $Y2=0
cc_420 N_A_183_290#_c_389_n N_A_575_87#_c_597_n 0.0172952f $X=2.47 $Y=1.68 $X2=0
+ $Y2=0
cc_421 N_A_183_290#_c_390_n N_A_575_87#_c_597_n 0.00120934f $X=2.47 $Y=1.68
+ $X2=0 $Y2=0
cc_422 N_A_183_290#_c_389_n N_A_575_87#_c_598_n 4.18224e-19 $X=2.47 $Y=1.68
+ $X2=0 $Y2=0
cc_423 N_A_183_290#_c_390_n N_A_575_87#_c_598_n 0.0369397f $X=2.47 $Y=1.68 $X2=0
+ $Y2=0
cc_424 N_A_183_290#_M1003_g N_A_32_74#_c_1913_n 0.00180084f $X=1.005 $Y=2.64
+ $X2=0 $Y2=0
cc_425 N_A_183_290#_M1003_g N_A_32_74#_c_1914_n 0.0204717f $X=1.005 $Y=2.64
+ $X2=0 $Y2=0
cc_426 N_A_183_290#_c_392_n N_A_32_74#_c_1914_n 0.00167134f $X=1.125 $Y=2.12
+ $X2=0 $Y2=0
cc_427 N_A_183_290#_c_394_n N_A_32_74#_c_1914_n 0.0255781f $X=1.825 $Y=2.035
+ $X2=0 $Y2=0
cc_428 N_A_183_290#_c_395_n N_A_32_74#_c_1914_n 0.0260356f $X=1.335 $Y=2.035
+ $X2=0 $Y2=0
cc_429 N_A_183_290#_c_396_n N_A_32_74#_c_1914_n 0.0141581f $X=1.91 $Y=2.51 $X2=0
+ $Y2=0
cc_430 N_A_183_290#_M1003_g N_A_32_74#_c_1915_n 0.00441379f $X=1.005 $Y=2.64
+ $X2=0 $Y2=0
cc_431 N_A_183_290#_c_396_n N_A_32_74#_c_1915_n 0.0203027f $X=1.91 $Y=2.51 $X2=0
+ $Y2=0
cc_432 N_A_183_290#_M1013_s N_A_32_74#_c_1916_n 0.00292485f $X=1.765 $Y=2.31
+ $X2=0 $Y2=0
cc_433 N_A_183_290#_c_396_n N_A_32_74#_c_1916_n 0.0123303f $X=1.91 $Y=2.51 $X2=0
+ $Y2=0
cc_434 N_A_183_290#_M1003_g N_A_32_74#_c_1917_n 6.68791e-19 $X=1.005 $Y=2.64
+ $X2=0 $Y2=0
cc_435 N_A_183_290#_c_397_n N_A_32_74#_c_1918_n 0.0237119f $X=2.305 $Y=2.035
+ $X2=0 $Y2=0
cc_436 N_A_183_290#_c_396_n N_A_32_74#_c_1919_n 0.00787895f $X=1.91 $Y=2.51
+ $X2=0 $Y2=0
cc_437 N_A_183_290#_c_397_n N_A_32_74#_c_1919_n 0.0136117f $X=2.305 $Y=2.035
+ $X2=0 $Y2=0
cc_438 N_A_183_290#_M1021_g N_A_32_74#_c_1908_n 0.00214472f $X=2.56 $Y=0.775
+ $X2=0 $Y2=0
cc_439 N_A_183_290#_M1021_g N_A_32_74#_c_1911_n 8.2814e-19 $X=2.56 $Y=0.775
+ $X2=0 $Y2=0
cc_440 N_A_183_290#_M1003_g N_VPWR_c_2024_n 0.0119286f $X=1.005 $Y=2.64 $X2=0
+ $Y2=0
cc_441 N_A_183_290#_M1003_g N_VPWR_c_2040_n 0.00460063f $X=1.005 $Y=2.64 $X2=0
+ $Y2=0
cc_442 N_A_183_290#_M1003_g N_VPWR_c_2023_n 0.00908371f $X=1.005 $Y=2.64 $X2=0
+ $Y2=0
cc_443 N_A_183_290#_c_385_n N_VGND_c_2461_n 2.63289e-19 $X=1.17 $Y=1.615 $X2=0
+ $Y2=0
cc_444 N_A_183_290#_c_386_n N_VGND_c_2461_n 0.00336712f $X=1.68 $Y=1.195 $X2=0
+ $Y2=0
cc_445 N_A_183_290#_c_387_n N_VGND_c_2461_n 0.0152311f $X=1.335 $Y=1.195 $X2=0
+ $Y2=0
cc_446 N_A_183_290#_c_388_n N_VGND_c_2461_n 0.0156036f $X=1.845 $Y=0.775 $X2=0
+ $Y2=0
cc_447 N_A_183_290#_M1021_g N_VGND_c_2462_n 0.0129344f $X=2.56 $Y=0.775 $X2=0
+ $Y2=0
cc_448 N_A_183_290#_c_388_n N_VGND_c_2462_n 0.0188413f $X=1.845 $Y=0.775 $X2=0
+ $Y2=0
cc_449 N_A_183_290#_c_389_n N_VGND_c_2462_n 0.00772803f $X=2.47 $Y=1.68 $X2=0
+ $Y2=0
cc_450 N_A_183_290#_c_390_n N_VGND_c_2462_n 0.0011905f $X=2.47 $Y=1.68 $X2=0
+ $Y2=0
cc_451 N_A_183_290#_c_388_n N_VGND_c_2477_n 0.00805126f $X=1.845 $Y=0.775 $X2=0
+ $Y2=0
cc_452 N_A_183_290#_M1021_g N_VGND_c_2483_n 0.00372658f $X=2.56 $Y=0.775 $X2=0
+ $Y2=0
cc_453 N_A_183_290#_M1021_g N_VGND_c_2496_n 0.00408518f $X=2.56 $Y=0.775 $X2=0
+ $Y2=0
cc_454 N_A_183_290#_c_388_n N_VGND_c_2496_n 0.0106012f $X=1.845 $Y=0.775 $X2=0
+ $Y2=0
cc_455 N_DE_c_503_n N_A_575_87#_M1024_g 0.0627553f $X=2.725 $Y=2.16 $X2=0 $Y2=0
cc_456 N_DE_c_503_n N_A_575_87#_c_598_n 0.00182507f $X=2.725 $Y=2.16 $X2=0 $Y2=0
cc_457 N_DE_c_502_n N_A_32_74#_c_1915_n 0.00342304f $X=2.135 $Y=2.235 $X2=0
+ $Y2=0
cc_458 N_DE_c_502_n N_A_32_74#_c_1916_n 0.0145926f $X=2.135 $Y=2.235 $X2=0 $Y2=0
cc_459 N_DE_c_504_n N_A_32_74#_c_1916_n 0.00219605f $X=2.225 $Y=2.16 $X2=0 $Y2=0
cc_460 N_DE_c_505_n N_A_32_74#_c_1916_n 4.3999e-19 $X=2.815 $Y=2.235 $X2=0 $Y2=0
cc_461 N_DE_c_502_n N_A_32_74#_c_1956_n 0.0122347f $X=2.135 $Y=2.235 $X2=0 $Y2=0
cc_462 N_DE_c_505_n N_A_32_74#_c_1956_n 0.00288039f $X=2.815 $Y=2.235 $X2=0
+ $Y2=0
cc_463 N_DE_c_503_n N_A_32_74#_c_1918_n 0.00657284f $X=2.725 $Y=2.16 $X2=0 $Y2=0
cc_464 N_DE_c_505_n N_A_32_74#_c_1918_n 0.0205385f $X=2.815 $Y=2.235 $X2=0 $Y2=0
cc_465 N_DE_c_502_n N_A_32_74#_c_1919_n 0.00630877f $X=2.135 $Y=2.235 $X2=0
+ $Y2=0
cc_466 N_DE_c_503_n N_A_32_74#_c_1919_n 4.60303e-19 $X=2.725 $Y=2.16 $X2=0 $Y2=0
cc_467 N_DE_M1042_g N_A_32_74#_c_1910_n 8.70603e-19 $X=1.02 $Y=0.58 $X2=0 $Y2=0
cc_468 N_DE_c_505_n N_A_32_74#_c_1922_n 0.00175158f $X=2.815 $Y=2.235 $X2=0
+ $Y2=0
cc_469 N_DE_c_502_n N_VPWR_c_2025_n 0.00145184f $X=2.135 $Y=2.235 $X2=0 $Y2=0
cc_470 N_DE_c_505_n N_VPWR_c_2025_n 0.0107317f $X=2.815 $Y=2.235 $X2=0 $Y2=0
cc_471 N_DE_c_502_n N_VPWR_c_2041_n 0.00468793f $X=2.135 $Y=2.235 $X2=0 $Y2=0
cc_472 N_DE_c_505_n N_VPWR_c_2042_n 0.00569568f $X=2.815 $Y=2.235 $X2=0 $Y2=0
cc_473 N_DE_c_502_n N_VPWR_c_2023_n 0.00651205f $X=2.135 $Y=2.235 $X2=0 $Y2=0
cc_474 N_DE_c_505_n N_VPWR_c_2023_n 0.00546289f $X=2.815 $Y=2.235 $X2=0 $Y2=0
cc_475 N_DE_M1042_g N_VGND_c_2461_n 0.0143553f $X=1.02 $Y=0.58 $X2=0 $Y2=0
cc_476 N_DE_c_493_n N_VGND_c_2461_n 0.00425745f $X=1.575 $Y=1.135 $X2=0 $Y2=0
cc_477 N_DE_c_496_n N_VGND_c_2461_n 0.00322863f $X=2.06 $Y=1.06 $X2=0 $Y2=0
cc_478 N_DE_c_496_n N_VGND_c_2462_n 0.00564371f $X=2.06 $Y=1.06 $X2=0 $Y2=0
cc_479 N_DE_c_496_n N_VGND_c_2477_n 0.00430863f $X=2.06 $Y=1.06 $X2=0 $Y2=0
cc_480 N_DE_M1042_g N_VGND_c_2482_n 0.00383152f $X=1.02 $Y=0.58 $X2=0 $Y2=0
cc_481 N_DE_M1042_g N_VGND_c_2496_n 0.0075725f $X=1.02 $Y=0.58 $X2=0 $Y2=0
cc_482 N_DE_c_496_n N_VGND_c_2496_n 0.00486331f $X=2.06 $Y=1.06 $X2=0 $Y2=0
cc_483 N_A_575_87#_M1005_g N_A_661_87#_c_868_n 0.0180128f $X=2.95 $Y=0.775 $X2=0
+ $Y2=0
cc_484 N_A_575_87#_c_595_n N_A_661_87#_c_869_n 0.00616126f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_485 N_A_575_87#_c_595_n N_A_661_87#_c_888_n 0.0186276f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_486 N_A_575_87#_c_595_n N_A_661_87#_c_873_n 0.00389277f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_487 N_A_575_87#_c_595_n N_A_661_87#_c_880_n 0.0516509f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_488 N_A_575_87#_c_595_n N_A_661_87#_c_881_n 0.00884701f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_489 N_A_575_87#_c_595_n N_A_661_87#_c_875_n 0.00594097f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_490 N_A_575_87#_c_598_n N_A_661_87#_c_875_n 0.00551319f $X=3.205 $Y=1.68
+ $X2=0 $Y2=0
cc_491 N_A_575_87#_c_595_n N_A_661_87#_c_883_n 0.00183705f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_492 N_A_575_87#_c_595_n N_A_661_87#_c_884_n 0.0192345f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_493 N_A_575_87#_c_595_n N_A_661_87#_c_876_n 0.00382946f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_494 N_A_575_87#_c_595_n N_SCD_M1031_g 0.00279625f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_495 N_A_575_87#_c_595_n SCD 0.0135615f $X=14.975 $Y=1.665 $X2=0 $Y2=0
cc_496 N_A_575_87#_c_595_n N_SCD_c_979_n 0.00380723f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_497 N_A_575_87#_M1024_g N_SCE_c_1024_n 0.0115875f $X=3.205 $Y=2.63 $X2=-0.19
+ $Y2=-0.245
cc_498 N_A_575_87#_c_595_n N_SCE_c_1024_n 0.00357925f $X=14.975 $Y=1.665
+ $X2=-0.19 $Y2=-0.245
cc_499 N_A_575_87#_c_595_n N_SCE_M1014_g 0.00267168f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_500 N_A_575_87#_c_595_n N_SCE_M1033_g 5.5049e-19 $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_501 N_A_575_87#_c_595_n N_SCE_c_1022_n 0.0043941f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_502 N_A_575_87#_c_595_n N_SCE_c_1023_n 0.0115832f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_503 N_A_575_87#_c_595_n N_CLK_M1000_g 0.00765274f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_504 N_A_575_87#_c_595_n CLK 0.012981f $X=14.975 $Y=1.665 $X2=0 $Y2=0
cc_505 N_A_575_87#_M1006_g N_A_1586_74#_M1030_g 0.0369612f $X=13.705 $Y=2.75
+ $X2=0 $Y2=0
cc_506 N_A_575_87#_c_605_n N_A_1586_74#_M1030_g 0.00104682f $X=14.475 $Y=2.217
+ $X2=0 $Y2=0
cc_507 N_A_575_87#_c_606_n N_A_1586_74#_M1030_g 0.0199166f $X=13.75 $Y=2.215
+ $X2=0 $Y2=0
cc_508 N_A_575_87#_c_595_n N_A_1586_74#_M1030_g 0.00305397f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_509 N_A_575_87#_c_599_n N_A_1586_74#_M1030_g 0.0151002f $X=13.75 $Y=2.05
+ $X2=0 $Y2=0
cc_510 N_A_575_87#_c_595_n N_A_1586_74#_c_1134_n 0.00221507f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_511 N_A_575_87#_c_595_n N_A_1586_74#_c_1157_n 0.0119622f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_512 N_A_575_87#_c_595_n N_A_1586_74#_c_1139_n 0.0070403f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_513 N_A_575_87#_c_595_n N_A_1586_74#_c_1140_n 7.16649e-19 $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_514 N_A_575_87#_c_595_n N_A_1586_74#_c_1141_n 0.00501141f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_515 N_A_575_87#_c_595_n N_A_1586_74#_c_1145_n 0.00603531f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_516 N_A_575_87#_c_595_n N_A_1586_74#_c_1146_n 3.66988e-19 $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_517 N_A_575_87#_c_595_n N_A_1586_74#_c_1148_n 0.0387409f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_518 N_A_575_87#_c_595_n N_A_1586_74#_c_1149_n 0.0165713f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_519 N_A_575_87#_c_595_n N_A_1586_74#_c_1159_n 0.00818568f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_520 N_A_575_87#_c_595_n N_A_1586_74#_c_1150_n 0.0201078f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_521 N_A_575_87#_c_595_n N_A_1586_74#_c_1161_n 0.00102983f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_522 N_A_575_87#_c_584_n N_A_1586_74#_c_1152_n 0.00221728f $X=13.345 $Y=0.94
+ $X2=0 $Y2=0
cc_523 N_A_575_87#_c_595_n N_A_1586_74#_c_1152_n 0.00886866f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_524 N_A_575_87#_c_599_n N_A_1586_74#_c_1152_n 9.53696e-19 $X=13.75 $Y=2.05
+ $X2=0 $Y2=0
cc_525 N_A_575_87#_c_584_n N_A_1586_74#_c_1153_n 0.0204808f $X=13.345 $Y=0.94
+ $X2=0 $Y2=0
cc_526 N_A_575_87#_c_595_n N_A_1586_74#_c_1153_n 0.00391026f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_527 N_A_575_87#_c_599_n N_A_1586_74#_c_1153_n 0.0173096f $X=13.75 $Y=2.05
+ $X2=0 $Y2=0
cc_528 N_A_575_87#_c_595_n N_A_1586_74#_c_1154_n 0.00371475f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_529 N_A_575_87#_c_595_n N_A_1377_368#_c_1364_n 2.73502e-19 $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_530 N_A_575_87#_c_595_n N_A_1377_368#_c_1365_n 0.00365728f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_531 N_A_575_87#_c_595_n N_A_1377_368#_c_1367_n 0.0122449f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_532 N_A_575_87#_c_582_n N_A_1377_368#_M1011_g 0.0417021f $X=13.27 $Y=0.865
+ $X2=0 $Y2=0
cc_533 N_A_575_87#_c_595_n N_A_1377_368#_c_1369_n 0.00240871f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_534 N_A_575_87#_c_595_n N_A_1377_368#_c_1370_n 0.00496775f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_535 N_A_575_87#_c_595_n N_A_1377_368#_c_1385_n 0.0146173f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_536 N_A_575_87#_c_595_n N_A_1377_368#_c_1387_n 0.0015259f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_537 N_A_575_87#_c_595_n N_A_1377_368#_c_1371_n 0.00629485f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_538 N_A_575_87#_c_595_n N_A_1377_368#_c_1372_n 0.0400993f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_539 N_A_575_87#_c_595_n N_A_1377_368#_c_1390_n 0.00208407f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_540 N_A_575_87#_c_595_n N_A_1377_368#_c_1374_n 0.030391f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_541 N_A_575_87#_c_595_n N_A_1377_368#_c_1375_n 6.94548e-19 $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_542 N_A_575_87#_c_595_n N_A_1377_368#_c_1376_n 0.0100197f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_543 N_A_575_87#_c_595_n N_A_2013_71#_M1016_g 0.00298149f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_544 N_A_575_87#_c_595_n N_A_2013_71#_c_1556_n 0.00463613f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_545 N_A_575_87#_c_595_n N_A_2013_71#_M1043_g 0.0128298f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_546 N_A_575_87#_c_595_n N_A_2013_71#_c_1559_n 0.0112107f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_547 N_A_575_87#_c_595_n N_A_2013_71#_c_1569_n 0.0117181f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_548 N_A_575_87#_c_595_n N_A_2013_71#_c_1561_n 0.0215524f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_549 N_A_575_87#_c_595_n N_A_2013_71#_c_1562_n 0.00903406f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_550 N_A_575_87#_c_595_n N_A_2013_71#_c_1563_n 0.0240966f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_551 N_A_575_87#_c_595_n N_A_2013_71#_c_1564_n 0.00849763f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_552 N_A_575_87#_c_595_n N_A_2013_71#_c_1565_n 0.00853542f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_553 N_A_575_87#_c_595_n N_A_1784_97#_c_1668_n 0.0141202f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_554 N_A_575_87#_c_595_n N_A_1784_97#_c_1671_n 0.0600244f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_555 N_A_575_87#_c_595_n N_A_1784_97#_c_1672_n 0.00882231f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_556 N_A_575_87#_c_595_n N_A_1784_97#_c_1675_n 0.0224528f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_557 N_A_575_87#_c_595_n N_A_1784_97#_c_1669_n 0.00373529f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_558 N_A_575_87#_M1006_g N_A_2489_74#_M1044_g 0.0133737f $X=13.705 $Y=2.75
+ $X2=0 $Y2=0
cc_559 N_A_575_87#_c_605_n N_A_2489_74#_M1044_g 0.0199941f $X=14.475 $Y=2.217
+ $X2=0 $Y2=0
cc_560 N_A_575_87#_c_589_n N_A_2489_74#_M1044_g 0.017091f $X=14.655 $Y=2.49
+ $X2=0 $Y2=0
cc_561 N_A_575_87#_c_608_n N_A_2489_74#_M1044_g 0.00869081f $X=14.64 $Y=2.815
+ $X2=0 $Y2=0
cc_562 N_A_575_87#_c_595_n N_A_2489_74#_M1044_g 0.00446587f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_563 N_A_575_87#_c_599_n N_A_2489_74#_M1044_g 0.0216668f $X=13.75 $Y=2.05
+ $X2=0 $Y2=0
cc_564 N_A_575_87#_c_583_n N_A_2489_74#_M1012_g 0.00727204f $X=13.765 $Y=0.94
+ $X2=0 $Y2=0
cc_565 N_A_575_87#_c_590_n N_A_2489_74#_M1012_g 0.00834476f $X=14.67 $Y=0.515
+ $X2=0 $Y2=0
cc_566 N_A_575_87#_c_591_n N_A_2489_74#_M1012_g 0.00600966f $X=14.75 $Y=1.55
+ $X2=0 $Y2=0
cc_567 N_A_575_87#_c_593_n N_A_2489_74#_M1012_g 0.00284604f $X=14.67 $Y=1.13
+ $X2=0 $Y2=0
cc_568 N_A_575_87#_c_589_n N_A_2489_74#_c_1757_n 0.0323203f $X=14.655 $Y=2.49
+ $X2=0 $Y2=0
cc_569 N_A_575_87#_c_591_n N_A_2489_74#_c_1757_n 0.0185398f $X=14.75 $Y=1.55
+ $X2=0 $Y2=0
cc_570 N_A_575_87#_c_593_n N_A_2489_74#_c_1757_n 0.00135743f $X=14.67 $Y=1.13
+ $X2=0 $Y2=0
cc_571 N_A_575_87#_c_595_n N_A_2489_74#_c_1757_n 0.00233301f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_572 N_A_575_87#_c_596_n N_A_2489_74#_c_1757_n 0.00658771f $X=15.12 $Y=1.665
+ $X2=0 $Y2=0
cc_573 N_A_575_87#_c_589_n N_A_2489_74#_M1036_g 0.0199041f $X=14.655 $Y=2.49
+ $X2=0 $Y2=0
cc_574 N_A_575_87#_c_608_n N_A_2489_74#_M1036_g 0.00422206f $X=14.64 $Y=2.815
+ $X2=0 $Y2=0
cc_575 N_A_575_87#_c_717_p N_A_2489_74#_M1036_g 0.0197773f $X=15.995 $Y=2.405
+ $X2=0 $Y2=0
cc_576 N_A_575_87#_c_596_n N_A_2489_74#_M1036_g 0.0043528f $X=15.12 $Y=1.665
+ $X2=0 $Y2=0
cc_577 N_A_575_87#_c_590_n N_A_2489_74#_M1026_g 0.00393219f $X=14.67 $Y=0.515
+ $X2=0 $Y2=0
cc_578 N_A_575_87#_M1002_g N_A_2489_74#_M1039_g 0.0439104f $X=16.325 $Y=2.4
+ $X2=0 $Y2=0
cc_579 N_A_575_87#_c_717_p N_A_2489_74#_M1039_g 0.0169107f $X=15.995 $Y=2.405
+ $X2=0 $Y2=0
cc_580 N_A_575_87#_c_592_n N_A_2489_74#_M1039_g 0.00367985f $X=16.09 $Y=2.32
+ $X2=0 $Y2=0
cc_581 N_A_575_87#_M1023_g N_A_2489_74#_M1047_g 0.0151259f $X=16.305 $Y=0.74
+ $X2=0 $Y2=0
cc_582 N_A_575_87#_c_717_p N_A_2489_74#_c_1762_n 2.28684e-19 $X=15.995 $Y=2.405
+ $X2=0 $Y2=0
cc_583 N_A_575_87#_c_594_n N_A_2489_74#_c_1762_n 0.00326102f $X=16.395 $Y=1.465
+ $X2=0 $Y2=0
cc_584 N_A_575_87#_c_600_n N_A_2489_74#_c_1762_n 0.0161842f $X=16.735 $Y=1.467
+ $X2=0 $Y2=0
cc_585 N_A_575_87#_c_582_n N_A_2489_74#_c_1764_n 0.00739677f $X=13.27 $Y=0.865
+ $X2=0 $Y2=0
cc_586 N_A_575_87#_c_583_n N_A_2489_74#_c_1764_n 0.0200523f $X=13.765 $Y=0.94
+ $X2=0 $Y2=0
cc_587 N_A_575_87#_c_584_n N_A_2489_74#_c_1764_n 0.00284537f $X=13.345 $Y=0.94
+ $X2=0 $Y2=0
cc_588 N_A_575_87#_M1006_g N_A_2489_74#_c_1772_n 8.29366e-19 $X=13.705 $Y=2.75
+ $X2=0 $Y2=0
cc_589 N_A_575_87#_c_605_n N_A_2489_74#_c_1772_n 0.017493f $X=14.475 $Y=2.217
+ $X2=0 $Y2=0
cc_590 N_A_575_87#_c_606_n N_A_2489_74#_c_1772_n 4.19728e-19 $X=13.75 $Y=2.215
+ $X2=0 $Y2=0
cc_591 N_A_575_87#_c_599_n N_A_2489_74#_c_1772_n 8.72783e-19 $X=13.75 $Y=2.05
+ $X2=0 $Y2=0
cc_592 N_A_575_87#_c_605_n N_A_2489_74#_c_1773_n 0.00772483f $X=14.475 $Y=2.217
+ $X2=0 $Y2=0
cc_593 N_A_575_87#_c_606_n N_A_2489_74#_c_1773_n 0.00279764f $X=13.75 $Y=2.215
+ $X2=0 $Y2=0
cc_594 N_A_575_87#_c_595_n N_A_2489_74#_c_1773_n 0.0191403f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_595 N_A_575_87#_c_599_n N_A_2489_74#_c_1773_n 3.91756e-19 $X=13.75 $Y=2.05
+ $X2=0 $Y2=0
cc_596 N_A_575_87#_c_595_n N_A_2489_74#_c_1774_n 0.0108527f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_597 N_A_575_87#_c_583_n N_A_2489_74#_c_1765_n 0.00639798f $X=13.765 $Y=0.94
+ $X2=0 $Y2=0
cc_598 N_A_575_87#_c_593_n N_A_2489_74#_c_1765_n 2.36907e-19 $X=14.67 $Y=1.13
+ $X2=0 $Y2=0
cc_599 N_A_575_87#_c_599_n N_A_2489_74#_c_1765_n 0.00974521f $X=13.75 $Y=2.05
+ $X2=0 $Y2=0
cc_600 N_A_575_87#_c_605_n N_A_2489_74#_c_1766_n 0.0128991f $X=14.475 $Y=2.217
+ $X2=0 $Y2=0
cc_601 N_A_575_87#_c_606_n N_A_2489_74#_c_1766_n 0.00189071f $X=13.75 $Y=2.215
+ $X2=0 $Y2=0
cc_602 N_A_575_87#_c_589_n N_A_2489_74#_c_1766_n 0.00223908f $X=14.655 $Y=2.49
+ $X2=0 $Y2=0
cc_603 N_A_575_87#_c_595_n N_A_2489_74#_c_1766_n 0.0191046f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_604 N_A_575_87#_c_599_n N_A_2489_74#_c_1766_n 0.0154352f $X=13.75 $Y=2.05
+ $X2=0 $Y2=0
cc_605 N_A_575_87#_c_605_n N_A_2489_74#_c_1767_n 0.0134002f $X=14.475 $Y=2.217
+ $X2=0 $Y2=0
cc_606 N_A_575_87#_c_589_n N_A_2489_74#_c_1767_n 0.00717225f $X=14.655 $Y=2.49
+ $X2=0 $Y2=0
cc_607 N_A_575_87#_c_591_n N_A_2489_74#_c_1767_n 0.0188124f $X=14.75 $Y=1.55
+ $X2=0 $Y2=0
cc_608 N_A_575_87#_c_595_n N_A_2489_74#_c_1767_n 0.0309319f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_609 N_A_575_87#_c_599_n N_A_2489_74#_c_1767_n 0.00891743f $X=13.75 $Y=2.05
+ $X2=0 $Y2=0
cc_610 N_A_575_87#_c_605_n N_A_2489_74#_c_1768_n 0.00188686f $X=14.475 $Y=2.217
+ $X2=0 $Y2=0
cc_611 N_A_575_87#_c_595_n N_A_2489_74#_c_1768_n 0.002332f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_612 N_A_575_87#_c_599_n N_A_2489_74#_c_1768_n 0.0172806f $X=13.75 $Y=2.05
+ $X2=0 $Y2=0
cc_613 N_A_575_87#_M1006_g N_A_2489_74#_c_1776_n 0.00185499f $X=13.705 $Y=2.75
+ $X2=0 $Y2=0
cc_614 N_A_575_87#_M1024_g N_A_32_74#_c_1918_n 0.0135821f $X=3.205 $Y=2.63 $X2=0
+ $Y2=0
cc_615 N_A_575_87#_c_618_n N_A_32_74#_c_1918_n 0.00294718f $X=3.265 $Y=1.665
+ $X2=0 $Y2=0
cc_616 N_A_575_87#_c_597_n N_A_32_74#_c_1918_n 0.010147f $X=3.04 $Y=1.68 $X2=0
+ $Y2=0
cc_617 N_A_575_87#_c_598_n N_A_32_74#_c_1918_n 0.00428552f $X=3.205 $Y=1.68
+ $X2=0 $Y2=0
cc_618 N_A_575_87#_M1005_g N_A_32_74#_c_1908_n 0.0139535f $X=2.95 $Y=0.775 $X2=0
+ $Y2=0
cc_619 N_A_575_87#_M1005_g N_A_32_74#_c_1909_n 0.00479218f $X=2.95 $Y=0.775
+ $X2=0 $Y2=0
cc_620 N_A_575_87#_c_595_n N_A_32_74#_c_1909_n 0.0165546f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_621 N_A_575_87#_c_618_n N_A_32_74#_c_1909_n 0.00240104f $X=3.265 $Y=1.665
+ $X2=0 $Y2=0
cc_622 N_A_575_87#_c_597_n N_A_32_74#_c_1909_n 0.0226176f $X=3.04 $Y=1.68 $X2=0
+ $Y2=0
cc_623 N_A_575_87#_c_598_n N_A_32_74#_c_1909_n 0.0173097f $X=3.205 $Y=1.68 $X2=0
+ $Y2=0
cc_624 N_A_575_87#_M1005_g N_A_32_74#_c_1911_n 0.00700496f $X=2.95 $Y=0.775
+ $X2=0 $Y2=0
cc_625 N_A_575_87#_c_595_n N_A_32_74#_c_1911_n 0.00516988f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_626 N_A_575_87#_c_618_n N_A_32_74#_c_1911_n 0.00394327f $X=3.265 $Y=1.665
+ $X2=0 $Y2=0
cc_627 N_A_575_87#_c_597_n N_A_32_74#_c_1911_n 0.0139741f $X=3.04 $Y=1.68 $X2=0
+ $Y2=0
cc_628 N_A_575_87#_c_598_n N_A_32_74#_c_1911_n 0.00812585f $X=3.205 $Y=1.68
+ $X2=0 $Y2=0
cc_629 N_A_575_87#_M1024_g N_A_32_74#_c_1922_n 0.0110121f $X=3.205 $Y=2.63 $X2=0
+ $Y2=0
cc_630 N_A_575_87#_c_595_n N_A_32_74#_c_1922_n 0.0037917f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_631 N_A_575_87#_c_605_n N_VPWR_M1006_d 0.00618258f $X=14.475 $Y=2.217 $X2=0
+ $Y2=0
cc_632 N_A_575_87#_c_589_n N_VPWR_M1036_s 0.0122256f $X=14.655 $Y=2.49 $X2=0
+ $Y2=0
cc_633 N_A_575_87#_c_717_p N_VPWR_M1036_s 0.00140071f $X=15.995 $Y=2.405 $X2=0
+ $Y2=0
cc_634 N_A_575_87#_c_717_p N_VPWR_M1039_s 0.00199514f $X=15.995 $Y=2.405 $X2=0
+ $Y2=0
cc_635 N_A_575_87#_c_592_n N_VPWR_M1039_s 0.00292416f $X=16.09 $Y=2.32 $X2=0
+ $Y2=0
cc_636 N_A_575_87#_M1024_g N_VPWR_c_2025_n 0.00146487f $X=3.205 $Y=2.63 $X2=0
+ $Y2=0
cc_637 N_A_575_87#_M1006_g N_VPWR_c_2031_n 0.0165816f $X=13.705 $Y=2.75 $X2=0
+ $Y2=0
cc_638 N_A_575_87#_c_605_n N_VPWR_c_2031_n 0.0283078f $X=14.475 $Y=2.217 $X2=0
+ $Y2=0
cc_639 N_A_575_87#_c_606_n N_VPWR_c_2031_n 0.00284999f $X=13.75 $Y=2.215 $X2=0
+ $Y2=0
cc_640 N_A_575_87#_c_608_n N_VPWR_c_2031_n 0.0133999f $X=14.64 $Y=2.815 $X2=0
+ $Y2=0
cc_641 N_A_575_87#_c_589_n N_VPWR_c_2032_n 0.0175754f $X=14.655 $Y=2.49 $X2=0
+ $Y2=0
cc_642 N_A_575_87#_c_608_n N_VPWR_c_2032_n 0.0239304f $X=14.64 $Y=2.815 $X2=0
+ $Y2=0
cc_643 N_A_575_87#_c_717_p N_VPWR_c_2032_n 0.00550577f $X=15.995 $Y=2.405 $X2=0
+ $Y2=0
cc_644 N_A_575_87#_M1002_g N_VPWR_c_2033_n 0.00894733f $X=16.325 $Y=2.4 $X2=0
+ $Y2=0
cc_645 N_A_575_87#_M1046_g N_VPWR_c_2033_n 3.30472e-19 $X=16.775 $Y=2.4 $X2=0
+ $Y2=0
cc_646 N_A_575_87#_c_717_p N_VPWR_c_2033_n 0.015845f $X=15.995 $Y=2.405 $X2=0
+ $Y2=0
cc_647 N_A_575_87#_M1002_g N_VPWR_c_2035_n 4.70425e-19 $X=16.325 $Y=2.4 $X2=0
+ $Y2=0
cc_648 N_A_575_87#_M1046_g N_VPWR_c_2035_n 0.0176187f $X=16.775 $Y=2.4 $X2=0
+ $Y2=0
cc_649 N_A_575_87#_M1024_g N_VPWR_c_2042_n 0.00653037f $X=3.205 $Y=2.63 $X2=0
+ $Y2=0
cc_650 N_A_575_87#_M1006_g N_VPWR_c_2045_n 0.00460063f $X=13.705 $Y=2.75 $X2=0
+ $Y2=0
cc_651 N_A_575_87#_c_608_n N_VPWR_c_2046_n 0.0158876f $X=14.64 $Y=2.815 $X2=0
+ $Y2=0
cc_652 N_A_575_87#_M1002_g N_VPWR_c_2048_n 0.00460063f $X=16.325 $Y=2.4 $X2=0
+ $Y2=0
cc_653 N_A_575_87#_M1046_g N_VPWR_c_2048_n 0.00460063f $X=16.775 $Y=2.4 $X2=0
+ $Y2=0
cc_654 N_A_575_87#_M1024_g N_VPWR_c_2023_n 0.00651205f $X=3.205 $Y=2.63 $X2=0
+ $Y2=0
cc_655 N_A_575_87#_M1006_g N_VPWR_c_2023_n 0.00908371f $X=13.705 $Y=2.75 $X2=0
+ $Y2=0
cc_656 N_A_575_87#_M1002_g N_VPWR_c_2023_n 0.00908554f $X=16.325 $Y=2.4 $X2=0
+ $Y2=0
cc_657 N_A_575_87#_M1046_g N_VPWR_c_2023_n 0.00908554f $X=16.775 $Y=2.4 $X2=0
+ $Y2=0
cc_658 N_A_575_87#_c_589_n N_VPWR_c_2023_n 0.00864971f $X=14.655 $Y=2.49 $X2=0
+ $Y2=0
cc_659 N_A_575_87#_c_608_n N_VPWR_c_2023_n 0.0130823f $X=14.64 $Y=2.815 $X2=0
+ $Y2=0
cc_660 N_A_575_87#_c_717_p N_VPWR_c_2023_n 0.0188721f $X=15.995 $Y=2.405 $X2=0
+ $Y2=0
cc_661 N_A_575_87#_c_595_n N_A_691_113#_c_2231_n 0.00288899f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_662 N_A_575_87#_M1024_g N_A_691_113#_c_2243_n 5.18417e-19 $X=3.205 $Y=2.63
+ $X2=0 $Y2=0
cc_663 N_A_575_87#_c_595_n N_A_691_113#_c_2233_n 0.00528828f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_664 N_A_575_87#_c_595_n N_A_691_113#_c_2234_n 0.00109913f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_665 N_A_575_87#_c_595_n N_A_691_113#_c_2224_n 0.0202067f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_666 N_A_575_87#_c_595_n N_A_691_113#_c_2236_n 0.0197345f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_667 N_A_575_87#_c_595_n N_A_691_113#_c_2237_n 0.00764576f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_668 N_A_575_87#_c_595_n N_A_691_113#_c_2238_n 0.013888f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_669 N_A_575_87#_c_595_n N_A_691_113#_c_2225_n 0.0347249f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_670 N_A_575_87#_c_595_n N_A_691_113#_c_2226_n 0.00439964f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_671 N_A_575_87#_c_595_n N_A_691_113#_c_2252_n 0.00274217f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_672 N_A_575_87#_c_595_n N_A_691_113#_c_2228_n 0.00579027f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_673 N_A_575_87#_M1005_g N_A_691_113#_c_2229_n 5.8879e-19 $X=2.95 $Y=0.775
+ $X2=0 $Y2=0
cc_674 N_A_575_87#_c_595_n N_A_691_113#_c_2229_n 0.0183113f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_675 N_A_575_87#_c_595_n N_A_691_113#_c_2230_n 0.00878755f $X=14.975 $Y=1.665
+ $X2=0 $Y2=0
cc_676 N_A_575_87#_c_717_p N_Q_M1036_d 0.00473092f $X=15.995 $Y=2.405 $X2=0
+ $Y2=0
cc_677 N_A_575_87#_M1023_g Q 0.0010619f $X=16.305 $Y=0.74 $X2=0 $Y2=0
cc_678 N_A_575_87#_c_589_n Q 0.0328163f $X=14.655 $Y=2.49 $X2=0 $Y2=0
cc_679 N_A_575_87#_c_591_n Q 0.0104168f $X=14.75 $Y=1.55 $X2=0 $Y2=0
cc_680 N_A_575_87#_c_717_p Q 0.0177876f $X=15.995 $Y=2.405 $X2=0 $Y2=0
cc_681 N_A_575_87#_c_592_n Q 0.0272185f $X=16.09 $Y=2.32 $X2=0 $Y2=0
cc_682 N_A_575_87#_c_594_n Q 0.0274627f $X=16.395 $Y=1.465 $X2=0 $Y2=0
cc_683 N_A_575_87#_c_596_n Q 0.00675851f $X=15.12 $Y=1.665 $X2=0 $Y2=0
cc_684 N_A_575_87#_c_600_n Q 2.32068e-19 $X=16.735 $Y=1.467 $X2=0 $Y2=0
cc_685 N_A_575_87#_M1023_g N_Q_N_c_2428_n 0.00237533f $X=16.305 $Y=0.74 $X2=0
+ $Y2=0
cc_686 N_A_575_87#_M1041_g N_Q_N_c_2428_n 0.0132482f $X=16.735 $Y=0.74 $X2=0
+ $Y2=0
cc_687 N_A_575_87#_c_594_n N_Q_N_c_2428_n 0.0115705f $X=16.395 $Y=1.465 $X2=0
+ $Y2=0
cc_688 N_A_575_87#_c_600_n N_Q_N_c_2428_n 0.00294111f $X=16.735 $Y=1.467 $X2=0
+ $Y2=0
cc_689 N_A_575_87#_M1023_g N_Q_N_c_2429_n 9.68429e-19 $X=16.305 $Y=0.74 $X2=0
+ $Y2=0
cc_690 N_A_575_87#_M1002_g N_Q_N_c_2429_n 3.50236e-19 $X=16.325 $Y=2.4 $X2=0
+ $Y2=0
cc_691 N_A_575_87#_M1041_g N_Q_N_c_2429_n 0.00816363f $X=16.735 $Y=0.74 $X2=0
+ $Y2=0
cc_692 N_A_575_87#_M1046_g N_Q_N_c_2429_n 0.0231607f $X=16.775 $Y=2.4 $X2=0
+ $Y2=0
cc_693 N_A_575_87#_c_592_n N_Q_N_c_2429_n 0.00784387f $X=16.09 $Y=2.32 $X2=0
+ $Y2=0
cc_694 N_A_575_87#_c_594_n N_Q_N_c_2429_n 0.0303249f $X=16.395 $Y=1.465 $X2=0
+ $Y2=0
cc_695 N_A_575_87#_c_600_n N_Q_N_c_2429_n 0.0207727f $X=16.735 $Y=1.467 $X2=0
+ $Y2=0
cc_696 N_A_575_87#_M1023_g Q_N 0.00756419f $X=16.305 $Y=0.74 $X2=0 $Y2=0
cc_697 N_A_575_87#_M1041_g Q_N 0.0133151f $X=16.735 $Y=0.74 $X2=0 $Y2=0
cc_698 N_A_575_87#_M1002_g Q_N 0.00395201f $X=16.325 $Y=2.4 $X2=0 $Y2=0
cc_699 N_A_575_87#_M1046_g Q_N 0.00395201f $X=16.775 $Y=2.4 $X2=0 $Y2=0
cc_700 N_A_575_87#_M1005_g N_VGND_c_2462_n 0.0018473f $X=2.95 $Y=0.775 $X2=0
+ $Y2=0
cc_701 N_A_575_87#_c_595_n N_VGND_c_2463_n 0.00383642f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_702 N_A_575_87#_c_595_n N_VGND_c_2465_n 0.00319228f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_703 N_A_575_87#_c_583_n N_VGND_c_2468_n 0.00216966f $X=13.765 $Y=0.94 $X2=0
+ $Y2=0
cc_704 N_A_575_87#_c_582_n N_VGND_c_2469_n 0.0105517f $X=13.27 $Y=0.865 $X2=0
+ $Y2=0
cc_705 N_A_575_87#_c_583_n N_VGND_c_2469_n 0.00310568f $X=13.765 $Y=0.94 $X2=0
+ $Y2=0
cc_706 N_A_575_87#_c_583_n N_VGND_c_2470_n 0.00246324f $X=13.765 $Y=0.94 $X2=0
+ $Y2=0
cc_707 N_A_575_87#_c_590_n N_VGND_c_2470_n 0.0198374f $X=14.67 $Y=0.515 $X2=0
+ $Y2=0
cc_708 N_A_575_87#_c_595_n N_VGND_c_2470_n 0.00126635f $X=14.975 $Y=1.665 $X2=0
+ $Y2=0
cc_709 N_A_575_87#_c_590_n N_VGND_c_2471_n 0.0145639f $X=14.67 $Y=0.515 $X2=0
+ $Y2=0
cc_710 N_A_575_87#_c_589_n N_VGND_c_2472_n 0.00440301f $X=14.655 $Y=2.49 $X2=0
+ $Y2=0
cc_711 N_A_575_87#_c_590_n N_VGND_c_2472_n 0.0514703f $X=14.67 $Y=0.515 $X2=0
+ $Y2=0
cc_712 N_A_575_87#_c_596_n N_VGND_c_2472_n 0.00254943f $X=15.12 $Y=1.665 $X2=0
+ $Y2=0
cc_713 N_A_575_87#_M1023_g N_VGND_c_2474_n 0.00315608f $X=16.305 $Y=0.74 $X2=0
+ $Y2=0
cc_714 N_A_575_87#_c_594_n N_VGND_c_2474_n 0.0148775f $X=16.395 $Y=1.465 $X2=0
+ $Y2=0
cc_715 N_A_575_87#_M1041_g N_VGND_c_2476_n 0.00611725f $X=16.735 $Y=0.74 $X2=0
+ $Y2=0
cc_716 N_A_575_87#_c_582_n N_VGND_c_2481_n 0.00383152f $X=13.27 $Y=0.865 $X2=0
+ $Y2=0
cc_717 N_A_575_87#_M1005_g N_VGND_c_2483_n 0.00430863f $X=2.95 $Y=0.775 $X2=0
+ $Y2=0
cc_718 N_A_575_87#_M1023_g N_VGND_c_2487_n 0.00434272f $X=16.305 $Y=0.74 $X2=0
+ $Y2=0
cc_719 N_A_575_87#_M1041_g N_VGND_c_2487_n 0.00434272f $X=16.735 $Y=0.74 $X2=0
+ $Y2=0
cc_720 N_A_575_87#_c_590_n N_VGND_c_2493_n 0.0103109f $X=14.67 $Y=0.515 $X2=0
+ $Y2=0
cc_721 N_A_575_87#_M1005_g N_VGND_c_2496_n 0.00486331f $X=2.95 $Y=0.775 $X2=0
+ $Y2=0
cc_722 N_A_575_87#_c_582_n N_VGND_c_2496_n 0.00367447f $X=13.27 $Y=0.865 $X2=0
+ $Y2=0
cc_723 N_A_575_87#_M1023_g N_VGND_c_2496_n 0.00820382f $X=16.305 $Y=0.74 $X2=0
+ $Y2=0
cc_724 N_A_575_87#_M1041_g N_VGND_c_2496_n 0.00823877f $X=16.735 $Y=0.74 $X2=0
+ $Y2=0
cc_725 N_A_575_87#_c_590_n N_VGND_c_2496_n 0.0119984f $X=14.67 $Y=0.515 $X2=0
+ $Y2=0
cc_726 N_A_661_87#_c_878_n N_SCD_M1031_g 0.044978f $X=5.915 $Y=2.085 $X2=0 $Y2=0
cc_727 N_A_661_87#_c_880_n N_SCD_M1031_g 0.0128834f $X=5.805 $Y=1.765 $X2=0
+ $Y2=0
cc_728 N_A_661_87#_c_884_n N_SCD_M1031_g 0.00130006f $X=5.97 $Y=1.58 $X2=0 $Y2=0
cc_729 N_A_661_87#_c_880_n SCD 0.0330694f $X=5.805 $Y=1.765 $X2=0 $Y2=0
cc_730 N_A_661_87#_c_884_n SCD 0.00650547f $X=5.97 $Y=1.58 $X2=0 $Y2=0
cc_731 N_A_661_87#_c_876_n SCD 8.85081e-19 $X=5.97 $Y=1.58 $X2=0 $Y2=0
cc_732 N_A_661_87#_c_880_n N_SCD_c_979_n 0.00329296f $X=5.805 $Y=1.765 $X2=0
+ $Y2=0
cc_733 N_A_661_87#_c_884_n N_SCD_c_979_n 0.00122864f $X=5.97 $Y=1.58 $X2=0 $Y2=0
cc_734 N_A_661_87#_c_876_n N_SCD_c_979_n 0.044978f $X=5.97 $Y=1.58 $X2=0 $Y2=0
cc_735 N_A_661_87#_c_879_n N_SCE_c_1024_n 3.18939e-19 $X=4.22 $Y=2.245 $X2=-0.19
+ $Y2=-0.245
cc_736 N_A_661_87#_c_883_n N_SCE_c_1024_n 0.00107892f $X=4.44 $Y=2.49 $X2=-0.19
+ $Y2=-0.245
cc_737 N_A_661_87#_c_883_n N_SCE_c_1025_n 0.00207399f $X=4.44 $Y=2.49 $X2=0
+ $Y2=0
cc_738 N_A_661_87#_c_879_n N_SCE_M1014_g 0.00588825f $X=4.22 $Y=2.245 $X2=0
+ $Y2=0
cc_739 N_A_661_87#_c_880_n N_SCE_M1014_g 0.0153221f $X=5.805 $Y=1.765 $X2=0
+ $Y2=0
cc_740 N_A_661_87#_c_881_n N_SCE_M1014_g 0.00200108f $X=4.18 $Y=1.765 $X2=0
+ $Y2=0
cc_741 N_A_661_87#_c_875_n N_SCE_M1014_g 0.0241622f $X=4.18 $Y=1.89 $X2=0 $Y2=0
cc_742 N_A_661_87#_c_883_n N_SCE_M1014_g 0.00374935f $X=4.44 $Y=2.49 $X2=0 $Y2=0
cc_743 N_A_661_87#_c_872_n N_SCE_M1037_g 8.75597e-19 $X=4.18 $Y=1.01 $X2=0 $Y2=0
cc_744 N_A_661_87#_c_888_n N_SCE_M1037_g 8.91698e-19 $X=4.18 $Y=1.21 $X2=0 $Y2=0
cc_745 N_A_661_87#_c_873_n N_SCE_M1037_g 0.00549146f $X=4.625 $Y=0.805 $X2=0
+ $Y2=0
cc_746 N_A_661_87#_c_874_n N_SCE_M1037_g 0.0176733f $X=4.18 $Y=0.53 $X2=0 $Y2=0
cc_747 N_A_661_87#_c_880_n N_SCE_M1033_g 7.90301e-19 $X=5.805 $Y=1.765 $X2=0
+ $Y2=0
cc_748 N_A_661_87#_c_876_n N_SCE_M1033_g 0.0100355f $X=5.97 $Y=1.58 $X2=0 $Y2=0
cc_749 N_A_661_87#_c_871_n N_SCE_c_1022_n 0.0241622f $X=4.18 $Y=1.135 $X2=0
+ $Y2=0
cc_750 N_A_661_87#_c_888_n N_SCE_c_1022_n 9.78573e-19 $X=4.18 $Y=1.21 $X2=0
+ $Y2=0
cc_751 N_A_661_87#_c_873_n N_SCE_c_1022_n 0.00467945f $X=4.625 $Y=0.805 $X2=0
+ $Y2=0
cc_752 N_A_661_87#_c_880_n N_SCE_c_1022_n 0.00388395f $X=5.805 $Y=1.765 $X2=0
+ $Y2=0
cc_753 N_A_661_87#_c_871_n N_SCE_c_1023_n 0.00222389f $X=4.18 $Y=1.135 $X2=0
+ $Y2=0
cc_754 N_A_661_87#_c_888_n N_SCE_c_1023_n 0.0261395f $X=4.18 $Y=1.21 $X2=0 $Y2=0
cc_755 N_A_661_87#_c_873_n N_SCE_c_1023_n 0.0223339f $X=4.625 $Y=0.805 $X2=0
+ $Y2=0
cc_756 N_A_661_87#_c_880_n N_SCE_c_1023_n 0.0283146f $X=5.805 $Y=1.765 $X2=0
+ $Y2=0
cc_757 N_A_661_87#_c_878_n N_CLK_M1000_g 0.00512042f $X=5.915 $Y=2.085 $X2=0
+ $Y2=0
cc_758 N_A_661_87#_c_876_n N_CLK_c_1094_n 0.00512042f $X=5.97 $Y=1.58 $X2=0
+ $Y2=0
cc_759 N_A_661_87#_c_868_n N_A_32_74#_c_1908_n 0.00745701f $X=3.38 $Y=1.06 $X2=0
+ $Y2=0
cc_760 N_A_661_87#_c_870_n N_A_32_74#_c_1908_n 0.00424876f $X=3.455 $Y=1.135
+ $X2=0 $Y2=0
cc_761 N_A_661_87#_c_870_n N_A_32_74#_c_1909_n 9.15581e-19 $X=3.455 $Y=1.135
+ $X2=0 $Y2=0
cc_762 N_A_661_87#_c_869_n N_A_32_74#_c_1911_n 0.00486125f $X=4.015 $Y=1.135
+ $X2=0 $Y2=0
cc_763 N_A_661_87#_c_870_n N_A_32_74#_c_1911_n 0.00908768f $X=3.455 $Y=1.135
+ $X2=0 $Y2=0
cc_764 N_A_661_87#_M1040_g N_VPWR_c_2026_n 0.00146667f $X=5.785 $Y=2.585 $X2=0
+ $Y2=0
cc_765 N_A_661_87#_M1040_g N_VPWR_c_2027_n 0.00290007f $X=5.785 $Y=2.585 $X2=0
+ $Y2=0
cc_766 N_A_661_87#_M1040_g N_VPWR_c_2036_n 0.00615629f $X=5.785 $Y=2.585 $X2=0
+ $Y2=0
cc_767 N_A_661_87#_M1040_g N_VPWR_c_2023_n 0.00634024f $X=5.785 $Y=2.585 $X2=0
+ $Y2=0
cc_768 N_A_661_87#_c_883_n N_A_691_113#_c_2231_n 0.0362005f $X=4.44 $Y=2.49
+ $X2=0 $Y2=0
cc_769 N_A_661_87#_c_883_n N_A_691_113#_c_2232_n 0.0295498f $X=4.44 $Y=2.49
+ $X2=0 $Y2=0
cc_770 N_A_661_87#_c_883_n N_A_691_113#_c_2259_n 0.0232576f $X=4.44 $Y=2.49
+ $X2=0 $Y2=0
cc_771 N_A_661_87#_M1040_g N_A_691_113#_c_2233_n 0.0133138f $X=5.785 $Y=2.585
+ $X2=0 $Y2=0
cc_772 N_A_661_87#_c_880_n N_A_691_113#_c_2233_n 0.0308201f $X=5.805 $Y=1.765
+ $X2=0 $Y2=0
cc_773 N_A_661_87#_c_884_n N_A_691_113#_c_2233_n 0.00284364f $X=5.97 $Y=1.58
+ $X2=0 $Y2=0
cc_774 N_A_661_87#_c_880_n N_A_691_113#_c_2234_n 0.00599699f $X=5.805 $Y=1.765
+ $X2=0 $Y2=0
cc_775 N_A_661_87#_c_883_n N_A_691_113#_c_2234_n 0.0142675f $X=4.44 $Y=2.49
+ $X2=0 $Y2=0
cc_776 N_A_661_87#_M1040_g N_A_691_113#_c_2224_n 0.00448935f $X=5.785 $Y=2.585
+ $X2=0 $Y2=0
cc_777 N_A_661_87#_c_884_n N_A_691_113#_c_2224_n 0.0481738f $X=5.97 $Y=1.58
+ $X2=0 $Y2=0
cc_778 N_A_661_87#_c_876_n N_A_691_113#_c_2224_n 0.00638291f $X=5.97 $Y=1.58
+ $X2=0 $Y2=0
cc_779 N_A_661_87#_M1040_g N_A_691_113#_c_2237_n 0.011321f $X=5.785 $Y=2.585
+ $X2=0 $Y2=0
cc_780 N_A_661_87#_c_878_n N_A_691_113#_c_2237_n 0.0020149f $X=5.915 $Y=2.085
+ $X2=0 $Y2=0
cc_781 N_A_661_87#_c_884_n N_A_691_113#_c_2237_n 0.024676f $X=5.97 $Y=1.58 $X2=0
+ $Y2=0
cc_782 N_A_661_87#_c_868_n N_A_691_113#_c_2228_n 0.00364479f $X=3.38 $Y=1.06
+ $X2=0 $Y2=0
cc_783 N_A_661_87#_c_869_n N_A_691_113#_c_2228_n 0.00746942f $X=4.015 $Y=1.135
+ $X2=0 $Y2=0
cc_784 N_A_661_87#_c_872_n N_A_691_113#_c_2228_n 0.0390571f $X=4.18 $Y=1.01
+ $X2=0 $Y2=0
cc_785 N_A_661_87#_c_874_n N_A_691_113#_c_2228_n 0.00543315f $X=4.18 $Y=0.53
+ $X2=0 $Y2=0
cc_786 N_A_661_87#_c_868_n N_A_691_113#_c_2229_n 4.83295e-19 $X=3.38 $Y=1.06
+ $X2=0 $Y2=0
cc_787 N_A_661_87#_c_869_n N_A_691_113#_c_2229_n 0.0150982f $X=4.015 $Y=1.135
+ $X2=0 $Y2=0
cc_788 N_A_661_87#_c_888_n N_A_691_113#_c_2229_n 0.0753924f $X=4.18 $Y=1.21
+ $X2=0 $Y2=0
cc_789 N_A_661_87#_c_879_n N_A_691_113#_c_2229_n 0.0109072f $X=4.22 $Y=2.245
+ $X2=0 $Y2=0
cc_790 N_A_661_87#_c_875_n N_A_691_113#_c_2229_n 0.013121f $X=4.18 $Y=1.89 $X2=0
+ $Y2=0
cc_791 N_A_661_87#_c_883_n N_A_691_113#_c_2229_n 0.00268191f $X=4.44 $Y=2.49
+ $X2=0 $Y2=0
cc_792 N_A_661_87#_c_884_n N_A_691_113#_c_2230_n 0.0235691f $X=5.97 $Y=1.58
+ $X2=0 $Y2=0
cc_793 N_A_661_87#_c_876_n N_A_691_113#_c_2230_n 0.00784966f $X=5.97 $Y=1.58
+ $X2=0 $Y2=0
cc_794 N_A_661_87#_c_872_n N_VGND_c_2463_n 0.00663031f $X=4.18 $Y=1.01 $X2=0
+ $Y2=0
cc_795 N_A_661_87#_c_873_n N_VGND_c_2463_n 0.0177281f $X=4.625 $Y=0.805 $X2=0
+ $Y2=0
cc_796 N_A_661_87#_c_880_n N_VGND_c_2463_n 0.00247704f $X=5.805 $Y=1.765 $X2=0
+ $Y2=0
cc_797 N_A_661_87#_c_868_n N_VGND_c_2483_n 0.00430863f $X=3.38 $Y=1.06 $X2=0
+ $Y2=0
cc_798 N_A_661_87#_c_872_n N_VGND_c_2483_n 0.00979148f $X=4.18 $Y=1.01 $X2=0
+ $Y2=0
cc_799 N_A_661_87#_c_873_n N_VGND_c_2483_n 0.00989191f $X=4.625 $Y=0.805 $X2=0
+ $Y2=0
cc_800 N_A_661_87#_c_874_n N_VGND_c_2483_n 0.0036882f $X=4.18 $Y=0.53 $X2=0
+ $Y2=0
cc_801 N_A_661_87#_c_868_n N_VGND_c_2496_n 0.00486331f $X=3.38 $Y=1.06 $X2=0
+ $Y2=0
cc_802 N_A_661_87#_c_872_n N_VGND_c_2496_n 0.00893856f $X=4.18 $Y=1.01 $X2=0
+ $Y2=0
cc_803 N_A_661_87#_c_873_n N_VGND_c_2496_n 0.0145109f $X=4.625 $Y=0.805 $X2=0
+ $Y2=0
cc_804 N_A_661_87#_c_874_n N_VGND_c_2496_n 0.00270334f $X=4.18 $Y=0.53 $X2=0
+ $Y2=0
cc_805 N_SCD_M1031_g N_SCE_M1014_g 0.0313259f $X=5.365 $Y=2.585 $X2=0 $Y2=0
cc_806 N_SCD_M1017_g N_SCE_M1037_g 0.013329f $X=5.38 $Y=0.835 $X2=0 $Y2=0
cc_807 N_SCD_M1017_g N_SCE_c_1019_n 0.00907339f $X=5.38 $Y=0.835 $X2=0 $Y2=0
cc_808 N_SCD_M1017_g N_SCE_M1033_g 0.0345301f $X=5.38 $Y=0.835 $X2=0 $Y2=0
cc_809 SCD N_SCE_c_1022_n 4.12687e-19 $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_810 N_SCD_c_979_n N_SCE_c_1022_n 0.0214313f $X=5.29 $Y=1.345 $X2=0 $Y2=0
cc_811 SCD N_SCE_c_1023_n 0.0221522f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_812 N_SCD_c_979_n N_SCE_c_1023_n 4.13447e-19 $X=5.29 $Y=1.345 $X2=0 $Y2=0
cc_813 N_SCD_M1031_g N_VPWR_c_2026_n 0.0109071f $X=5.365 $Y=2.585 $X2=0 $Y2=0
cc_814 N_SCD_M1031_g N_VPWR_c_2036_n 0.00536686f $X=5.365 $Y=2.585 $X2=0 $Y2=0
cc_815 N_SCD_M1031_g N_VPWR_c_2023_n 0.00531876f $X=5.365 $Y=2.585 $X2=0 $Y2=0
cc_816 N_SCD_M1031_g N_A_691_113#_c_2232_n 3.50727e-19 $X=5.365 $Y=2.585 $X2=0
+ $Y2=0
cc_817 N_SCD_M1031_g N_A_691_113#_c_2259_n 0.00280416f $X=5.365 $Y=2.585 $X2=0
+ $Y2=0
cc_818 N_SCD_M1031_g N_A_691_113#_c_2233_n 0.0182826f $X=5.365 $Y=2.585 $X2=0
+ $Y2=0
cc_819 N_SCD_M1017_g N_A_691_113#_c_2223_n 0.00156538f $X=5.38 $Y=0.835 $X2=0
+ $Y2=0
cc_820 SCD N_A_691_113#_c_2224_n 0.00535427f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_821 N_SCD_M1031_g N_A_691_113#_c_2237_n 0.00174746f $X=5.365 $Y=2.585 $X2=0
+ $Y2=0
cc_822 N_SCD_M1017_g N_A_691_113#_c_2230_n 5.99886e-19 $X=5.38 $Y=0.835 $X2=0
+ $Y2=0
cc_823 SCD N_A_691_113#_c_2230_n 0.00671568f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_824 N_SCD_c_979_n N_A_691_113#_c_2230_n 4.02826e-19 $X=5.29 $Y=1.345 $X2=0
+ $Y2=0
cc_825 N_SCD_M1017_g N_VGND_c_2463_n 0.0036597f $X=5.38 $Y=0.835 $X2=0 $Y2=0
cc_826 SCD N_VGND_c_2463_n 0.0114218f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_827 N_SCD_c_979_n N_VGND_c_2463_n 0.00375077f $X=5.29 $Y=1.345 $X2=0 $Y2=0
cc_828 N_SCD_M1017_g N_VGND_c_2496_n 9.49986e-19 $X=5.38 $Y=0.835 $X2=0 $Y2=0
cc_829 N_SCE_c_1024_n N_A_32_74#_c_1909_n 8.29346e-19 $X=3.655 $Y=3.025 $X2=0
+ $Y2=0
cc_830 N_SCE_c_1025_n N_VPWR_c_2026_n 0.00271219f $X=4.585 $Y=3.1 $X2=0 $Y2=0
cc_831 N_SCE_M1014_g N_VPWR_c_2026_n 0.00160643f $X=4.675 $Y=2.585 $X2=0 $Y2=0
cc_832 N_SCE_c_1026_n N_VPWR_c_2042_n 0.0258782f $X=3.745 $Y=3.1 $X2=0 $Y2=0
cc_833 N_SCE_c_1025_n N_VPWR_c_2023_n 0.0261661f $X=4.585 $Y=3.1 $X2=0 $Y2=0
cc_834 N_SCE_c_1026_n N_VPWR_c_2023_n 0.011582f $X=3.745 $Y=3.1 $X2=0 $Y2=0
cc_835 N_SCE_c_1024_n N_A_691_113#_c_2231_n 0.00175302f $X=3.655 $Y=3.025 $X2=0
+ $Y2=0
cc_836 N_SCE_M1014_g N_A_691_113#_c_2231_n 0.00438085f $X=4.675 $Y=2.585 $X2=0
+ $Y2=0
cc_837 N_SCE_c_1024_n N_A_691_113#_c_2294_n 0.00545621f $X=3.655 $Y=3.025 $X2=0
+ $Y2=0
cc_838 N_SCE_c_1025_n N_A_691_113#_c_2232_n 0.0191584f $X=4.585 $Y=3.1 $X2=0
+ $Y2=0
cc_839 N_SCE_M1014_g N_A_691_113#_c_2232_n 0.0109005f $X=4.675 $Y=2.585 $X2=0
+ $Y2=0
cc_840 N_SCE_c_1024_n N_A_691_113#_c_2243_n 0.00361732f $X=3.655 $Y=3.025 $X2=0
+ $Y2=0
cc_841 N_SCE_c_1025_n N_A_691_113#_c_2243_n 0.00577343f $X=4.585 $Y=3.1 $X2=0
+ $Y2=0
cc_842 N_SCE_c_1026_n N_A_691_113#_c_2243_n 0.00125602f $X=3.745 $Y=3.1 $X2=0
+ $Y2=0
cc_843 N_SCE_M1014_g N_A_691_113#_c_2259_n 0.0169951f $X=4.675 $Y=2.585 $X2=0
+ $Y2=0
cc_844 N_SCE_M1014_g N_A_691_113#_c_2234_n 0.00712881f $X=4.675 $Y=2.585 $X2=0
+ $Y2=0
cc_845 N_SCE_M1033_g N_A_691_113#_c_2223_n 0.0109232f $X=5.77 $Y=0.835 $X2=0
+ $Y2=0
cc_846 N_SCE_c_1024_n N_A_691_113#_c_2229_n 0.00380768f $X=3.655 $Y=3.025 $X2=0
+ $Y2=0
cc_847 N_SCE_M1033_g N_A_691_113#_c_2230_n 0.00377254f $X=5.77 $Y=0.835 $X2=0
+ $Y2=0
cc_848 N_SCE_M1037_g N_VGND_c_2463_n 0.0126683f $X=4.84 $Y=0.835 $X2=0 $Y2=0
cc_849 N_SCE_c_1019_n N_VGND_c_2463_n 0.0244098f $X=5.695 $Y=0.18 $X2=0 $Y2=0
cc_850 N_SCE_M1033_g N_VGND_c_2463_n 0.00789535f $X=5.77 $Y=0.835 $X2=0 $Y2=0
cc_851 N_SCE_c_1019_n N_VGND_c_2464_n 0.0109961f $X=5.695 $Y=0.18 $X2=0 $Y2=0
cc_852 N_SCE_M1033_g N_VGND_c_2464_n 6.60132e-19 $X=5.77 $Y=0.835 $X2=0 $Y2=0
cc_853 N_SCE_c_1020_n N_VGND_c_2483_n 0.00729633f $X=4.915 $Y=0.18 $X2=0 $Y2=0
cc_854 N_SCE_c_1019_n N_VGND_c_2484_n 0.0201823f $X=5.695 $Y=0.18 $X2=0 $Y2=0
cc_855 N_SCE_c_1019_n N_VGND_c_2496_n 0.0326416f $X=5.695 $Y=0.18 $X2=0 $Y2=0
cc_856 N_SCE_c_1020_n N_VGND_c_2496_n 0.0106185f $X=4.915 $Y=0.18 $X2=0 $Y2=0
cc_857 N_CLK_M1000_g N_A_1377_368#_c_1385_n 0.00662111f $X=6.795 $Y=2.4 $X2=0
+ $Y2=0
cc_858 CLK N_A_1377_368#_c_1385_n 0.00655916f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_859 N_CLK_c_1094_n N_A_1377_368#_c_1385_n 0.00102013f $X=6.87 $Y=1.385 $X2=0
+ $Y2=0
cc_860 CLK N_A_1377_368#_c_1371_n 0.00829649f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_861 N_CLK_c_1094_n N_A_1377_368#_c_1371_n 5.12853e-19 $X=6.87 $Y=1.385 $X2=0
+ $Y2=0
cc_862 N_CLK_c_1095_n N_A_1377_368#_c_1371_n 0.0115578f $X=6.87 $Y=1.22 $X2=0
+ $Y2=0
cc_863 N_CLK_M1000_g N_A_1377_368#_c_1372_n 0.00489956f $X=6.795 $Y=2.4 $X2=0
+ $Y2=0
cc_864 CLK N_A_1377_368#_c_1373_n 0.0298284f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_865 N_CLK_c_1094_n N_A_1377_368#_c_1373_n 0.00200244f $X=6.87 $Y=1.385 $X2=0
+ $Y2=0
cc_866 N_CLK_c_1095_n N_A_1377_368#_c_1373_n 0.00389062f $X=6.87 $Y=1.22 $X2=0
+ $Y2=0
cc_867 N_CLK_M1000_g N_A_1377_368#_c_1376_n 0.0107805f $X=6.795 $Y=2.4 $X2=0
+ $Y2=0
cc_868 CLK N_A_1377_368#_c_1376_n 2.18476e-19 $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_869 N_CLK_c_1094_n N_A_1377_368#_c_1376_n 0.00348307f $X=6.87 $Y=1.385 $X2=0
+ $Y2=0
cc_870 N_CLK_M1000_g N_VPWR_c_2027_n 0.0221646f $X=6.795 $Y=2.4 $X2=0 $Y2=0
cc_871 N_CLK_M1000_g N_VPWR_c_2043_n 0.00460063f $X=6.795 $Y=2.4 $X2=0 $Y2=0
cc_872 N_CLK_M1000_g N_VPWR_c_2023_n 0.00468499f $X=6.795 $Y=2.4 $X2=0 $Y2=0
cc_873 N_CLK_c_1095_n N_A_691_113#_c_2223_n 0.00440404f $X=6.87 $Y=1.22 $X2=0
+ $Y2=0
cc_874 CLK N_A_691_113#_c_2224_n 0.0174202f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_875 N_CLK_c_1094_n N_A_691_113#_c_2224_n 0.0172136f $X=6.87 $Y=1.385 $X2=0
+ $Y2=0
cc_876 N_CLK_M1000_g N_A_691_113#_c_2236_n 0.0188567f $X=6.795 $Y=2.4 $X2=0
+ $Y2=0
cc_877 N_CLK_M1000_g N_A_691_113#_c_2237_n 0.00700241f $X=6.795 $Y=2.4 $X2=0
+ $Y2=0
cc_878 CLK N_A_691_113#_c_2230_n 0.0054797f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_879 N_CLK_c_1094_n N_A_691_113#_c_2230_n 8.76987e-19 $X=6.87 $Y=1.385 $X2=0
+ $Y2=0
cc_880 N_CLK_c_1095_n N_A_691_113#_c_2230_n 0.00334486f $X=6.87 $Y=1.22 $X2=0
+ $Y2=0
cc_881 CLK N_VGND_c_2464_n 0.00209233f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_882 N_CLK_c_1094_n N_VGND_c_2464_n 2.21134e-19 $X=6.87 $Y=1.385 $X2=0 $Y2=0
cc_883 N_CLK_c_1095_n N_VGND_c_2464_n 0.0157427f $X=6.87 $Y=1.22 $X2=0 $Y2=0
cc_884 N_CLK_c_1095_n N_VGND_c_2465_n 0.00305448f $X=6.87 $Y=1.22 $X2=0 $Y2=0
cc_885 N_CLK_c_1095_n N_VGND_c_2479_n 0.00434272f $X=6.87 $Y=1.22 $X2=0 $Y2=0
cc_886 N_CLK_c_1095_n N_VGND_c_2496_n 0.00830058f $X=6.87 $Y=1.22 $X2=0 $Y2=0
cc_887 N_A_1586_74#_c_1134_n N_A_1377_368#_M1004_g 0.00979223f $X=8.07 $Y=0.515
+ $X2=0 $Y2=0
cc_888 N_A_1586_74#_c_1136_n N_A_1377_368#_M1004_g 0.00474255f $X=8.235 $Y=0.34
+ $X2=0 $Y2=0
cc_889 N_A_1586_74#_c_1134_n N_A_1377_368#_c_1364_n 0.00127711f $X=8.07 $Y=0.515
+ $X2=0 $Y2=0
cc_890 N_A_1586_74#_c_1157_n N_A_1377_368#_c_1378_n 0.00485867f $X=8.725 $Y=1.98
+ $X2=0 $Y2=0
cc_891 N_A_1586_74#_c_1159_n N_A_1377_368#_c_1378_n 4.73056e-19 $X=8.89 $Y=1.98
+ $X2=0 $Y2=0
cc_892 N_A_1586_74#_c_1150_n N_A_1377_368#_c_1378_n 0.00186049f $X=8.89 $Y=1.82
+ $X2=0 $Y2=0
cc_893 N_A_1586_74#_c_1161_n N_A_1377_368#_c_1378_n 0.00530826f $X=8.89 $Y=2.14
+ $X2=0 $Y2=0
cc_894 N_A_1586_74#_c_1157_n N_A_1377_368#_c_1365_n 0.00704839f $X=8.725 $Y=1.98
+ $X2=0 $Y2=0
cc_895 N_A_1586_74#_c_1159_n N_A_1377_368#_c_1365_n 0.00441444f $X=8.89 $Y=1.98
+ $X2=0 $Y2=0
cc_896 N_A_1586_74#_c_1161_n N_A_1377_368#_c_1365_n 0.0186888f $X=8.89 $Y=2.14
+ $X2=0 $Y2=0
cc_897 N_A_1586_74#_c_1131_n N_A_1377_368#_M1035_g 0.013497f $X=9.525 $Y=1.015
+ $X2=0 $Y2=0
cc_898 N_A_1586_74#_c_1134_n N_A_1377_368#_M1035_g 0.00327787f $X=8.07 $Y=0.515
+ $X2=0 $Y2=0
cc_899 N_A_1586_74#_c_1135_n N_A_1377_368#_M1035_g 0.00929412f $X=8.885 $Y=0.34
+ $X2=0 $Y2=0
cc_900 N_A_1586_74#_c_1150_n N_A_1377_368#_M1035_g 0.0298706f $X=8.89 $Y=1.82
+ $X2=0 $Y2=0
cc_901 N_A_1586_74#_c_1151_n N_A_1377_368#_M1035_g 0.00206916f $X=8.97 $Y=0.34
+ $X2=0 $Y2=0
cc_902 N_A_1586_74#_c_1139_n N_A_1377_368#_c_1367_n 4.9149e-19 $X=9.69 $Y=1.18
+ $X2=0 $Y2=0
cc_903 N_A_1586_74#_c_1140_n N_A_1377_368#_c_1367_n 0.0139692f $X=9.69 $Y=1.18
+ $X2=0 $Y2=0
cc_904 N_A_1586_74#_c_1150_n N_A_1377_368#_c_1367_n 0.0076216f $X=8.89 $Y=1.82
+ $X2=0 $Y2=0
cc_905 N_A_1586_74#_c_1161_n N_A_1377_368#_c_1367_n 0.00716403f $X=8.89 $Y=2.14
+ $X2=0 $Y2=0
cc_906 N_A_1586_74#_M1015_g N_A_1377_368#_M1019_g 0.0160665f $X=9.195 $Y=2.75
+ $X2=0 $Y2=0
cc_907 N_A_1586_74#_M1030_g N_A_1377_368#_M1034_g 0.0352231f $X=13.285 $Y=2.75
+ $X2=0 $Y2=0
cc_908 N_A_1586_74#_M1010_g N_A_1377_368#_M1011_g 0.0293304f $X=12.37 $Y=0.69
+ $X2=0 $Y2=0
cc_909 N_A_1586_74#_c_1148_n N_A_1377_368#_M1011_g 8.82425e-19 $X=12.26 $Y=1.635
+ $X2=0 $Y2=0
cc_910 N_A_1586_74#_c_1149_n N_A_1377_368#_M1011_g 0.0114972f $X=13.195 $Y=1.215
+ $X2=0 $Y2=0
cc_911 N_A_1586_74#_c_1152_n N_A_1377_368#_M1011_g 0.00153298f $X=13.36 $Y=1.215
+ $X2=0 $Y2=0
cc_912 N_A_1586_74#_c_1153_n N_A_1377_368#_M1011_g 0.0135859f $X=13.36 $Y=1.39
+ $X2=0 $Y2=0
cc_913 N_A_1586_74#_c_1150_n N_A_1377_368#_c_1370_n 0.00342855f $X=8.89 $Y=1.82
+ $X2=0 $Y2=0
cc_914 N_A_1586_74#_c_1148_n N_A_1377_368#_c_1386_n 0.00881567f $X=12.26
+ $Y=1.635 $X2=0 $Y2=0
cc_915 N_A_1586_74#_c_1154_n N_A_1377_368#_c_1386_n 0.00321743f $X=12.37
+ $Y=1.635 $X2=0 $Y2=0
cc_916 N_A_1586_74#_M1030_g N_A_1377_368#_c_1387_n 6.09453e-19 $X=13.285 $Y=2.75
+ $X2=0 $Y2=0
cc_917 N_A_1586_74#_c_1140_n N_A_1377_368#_c_1391_n 0.00184475f $X=9.69 $Y=1.18
+ $X2=0 $Y2=0
cc_918 N_A_1586_74#_c_1161_n N_A_1377_368#_c_1391_n 0.0107199f $X=8.89 $Y=2.14
+ $X2=0 $Y2=0
cc_919 N_A_1586_74#_c_1148_n N_A_1377_368#_c_1374_n 0.0248923f $X=12.26 $Y=1.635
+ $X2=0 $Y2=0
cc_920 N_A_1586_74#_c_1149_n N_A_1377_368#_c_1374_n 0.0303637f $X=13.195
+ $Y=1.215 $X2=0 $Y2=0
cc_921 N_A_1586_74#_c_1152_n N_A_1377_368#_c_1374_n 0.00481086f $X=13.36
+ $Y=1.215 $X2=0 $Y2=0
cc_922 N_A_1586_74#_c_1153_n N_A_1377_368#_c_1374_n 0.00193886f $X=13.36 $Y=1.39
+ $X2=0 $Y2=0
cc_923 N_A_1586_74#_c_1154_n N_A_1377_368#_c_1374_n 0.00195577f $X=12.37
+ $Y=1.635 $X2=0 $Y2=0
cc_924 N_A_1586_74#_c_1148_n N_A_1377_368#_c_1375_n 3.6914e-19 $X=12.26 $Y=1.635
+ $X2=0 $Y2=0
cc_925 N_A_1586_74#_c_1149_n N_A_1377_368#_c_1375_n 0.00460699f $X=13.195
+ $Y=1.215 $X2=0 $Y2=0
cc_926 N_A_1586_74#_c_1153_n N_A_1377_368#_c_1375_n 0.0213123f $X=13.36 $Y=1.39
+ $X2=0 $Y2=0
cc_927 N_A_1586_74#_c_1154_n N_A_1377_368#_c_1375_n 0.021367f $X=12.37 $Y=1.635
+ $X2=0 $Y2=0
cc_928 N_A_1586_74#_c_1150_n N_A_1377_368#_c_1395_n 4.63241e-19 $X=8.89 $Y=1.82
+ $X2=0 $Y2=0
cc_929 N_A_1586_74#_c_1161_n N_A_1377_368#_c_1395_n 0.00326764f $X=8.89 $Y=2.14
+ $X2=0 $Y2=0
cc_930 N_A_1586_74#_c_1142_n N_A_2013_71#_M1018_d 0.00350583f $X=11.37 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_931 N_A_1586_74#_c_1131_n N_A_2013_71#_M1025_g 0.013612f $X=9.525 $Y=1.015
+ $X2=0 $Y2=0
cc_932 N_A_1586_74#_c_1137_n N_A_2013_71#_M1025_g 7.07453e-19 $X=9.565 $Y=0.34
+ $X2=0 $Y2=0
cc_933 N_A_1586_74#_c_1138_n N_A_2013_71#_M1025_g 0.00524926f $X=9.65 $Y=0.85
+ $X2=0 $Y2=0
cc_934 N_A_1586_74#_c_1139_n N_A_2013_71#_M1025_g 0.00166923f $X=9.69 $Y=1.18
+ $X2=0 $Y2=0
cc_935 N_A_1586_74#_c_1140_n N_A_2013_71#_M1025_g 0.0210021f $X=9.69 $Y=1.18
+ $X2=0 $Y2=0
cc_936 N_A_1586_74#_c_1141_n N_A_2013_71#_M1025_g 0.0138659f $X=10.69 $Y=0.935
+ $X2=0 $Y2=0
cc_937 N_A_1586_74#_c_1237_p N_A_2013_71#_M1025_g 0.00308709f $X=10.775 $Y=0.85
+ $X2=0 $Y2=0
cc_938 N_A_1586_74#_M1010_g N_A_2013_71#_c_1556_n 0.0056233f $X=12.37 $Y=0.69
+ $X2=0 $Y2=0
cc_939 N_A_1586_74#_c_1147_n N_A_2013_71#_c_1556_n 0.00681315f $X=12.23 $Y=1.3
+ $X2=0 $Y2=0
cc_940 N_A_1586_74#_c_1148_n N_A_2013_71#_c_1556_n 0.00612673f $X=12.26 $Y=1.635
+ $X2=0 $Y2=0
cc_941 N_A_1586_74#_c_1154_n N_A_2013_71#_c_1556_n 0.021065f $X=12.37 $Y=1.635
+ $X2=0 $Y2=0
cc_942 N_A_1586_74#_M1010_g N_A_2013_71#_c_1558_n 0.0605761f $X=12.37 $Y=0.69
+ $X2=0 $Y2=0
cc_943 N_A_1586_74#_c_1142_n N_A_2013_71#_c_1558_n 6.63977e-19 $X=11.37 $Y=0.34
+ $X2=0 $Y2=0
cc_944 N_A_1586_74#_c_1144_n N_A_2013_71#_c_1558_n 0.004173f $X=11.455 $Y=0.85
+ $X2=0 $Y2=0
cc_945 N_A_1586_74#_c_1145_n N_A_2013_71#_c_1558_n 0.0123107f $X=12.08 $Y=0.935
+ $X2=0 $Y2=0
cc_946 N_A_1586_74#_c_1147_n N_A_2013_71#_c_1558_n 0.0052319f $X=12.23 $Y=1.3
+ $X2=0 $Y2=0
cc_947 N_A_1586_74#_c_1141_n N_A_2013_71#_c_1559_n 0.035239f $X=10.69 $Y=0.935
+ $X2=0 $Y2=0
cc_948 N_A_1586_74#_c_1141_n N_A_2013_71#_c_1560_n 0.00750114f $X=10.69 $Y=0.935
+ $X2=0 $Y2=0
cc_949 N_A_1586_74#_c_1142_n N_A_2013_71#_c_1560_n 0.0127109f $X=11.37 $Y=0.34
+ $X2=0 $Y2=0
cc_950 N_A_1586_74#_c_1144_n N_A_2013_71#_c_1560_n 0.0188234f $X=11.455 $Y=0.85
+ $X2=0 $Y2=0
cc_951 N_A_1586_74#_c_1146_n N_A_2013_71#_c_1560_n 0.0141448f $X=11.54 $Y=0.935
+ $X2=0 $Y2=0
cc_952 N_A_1586_74#_c_1146_n N_A_2013_71#_c_1562_n 0.00130064f $X=11.54 $Y=0.935
+ $X2=0 $Y2=0
cc_953 N_A_1586_74#_M1010_g N_A_2013_71#_c_1563_n 2.44748e-19 $X=12.37 $Y=0.69
+ $X2=0 $Y2=0
cc_954 N_A_1586_74#_c_1145_n N_A_2013_71#_c_1563_n 0.0251569f $X=12.08 $Y=0.935
+ $X2=0 $Y2=0
cc_955 N_A_1586_74#_c_1146_n N_A_2013_71#_c_1563_n 0.01265f $X=11.54 $Y=0.935
+ $X2=0 $Y2=0
cc_956 N_A_1586_74#_c_1147_n N_A_2013_71#_c_1563_n 0.00844044f $X=12.23 $Y=1.3
+ $X2=0 $Y2=0
cc_957 N_A_1586_74#_c_1148_n N_A_2013_71#_c_1563_n 0.0163961f $X=12.26 $Y=1.635
+ $X2=0 $Y2=0
cc_958 N_A_1586_74#_c_1142_n N_A_2013_71#_c_1564_n 0.00351137f $X=11.37 $Y=0.34
+ $X2=0 $Y2=0
cc_959 N_A_1586_74#_c_1145_n N_A_2013_71#_c_1564_n 0.0113034f $X=12.08 $Y=0.935
+ $X2=0 $Y2=0
cc_960 N_A_1586_74#_c_1146_n N_A_2013_71#_c_1564_n 0.00455524f $X=11.54 $Y=0.935
+ $X2=0 $Y2=0
cc_961 N_A_1586_74#_c_1139_n N_A_2013_71#_c_1565_n 0.00972664f $X=9.69 $Y=1.18
+ $X2=0 $Y2=0
cc_962 N_A_1586_74#_c_1140_n N_A_2013_71#_c_1565_n 5.60957e-19 $X=9.69 $Y=1.18
+ $X2=0 $Y2=0
cc_963 N_A_1586_74#_c_1141_n N_A_2013_71#_c_1565_n 0.0235913f $X=10.69 $Y=0.935
+ $X2=0 $Y2=0
cc_964 N_A_1586_74#_c_1141_n N_A_2013_71#_c_1566_n 0.00125903f $X=10.69 $Y=0.935
+ $X2=0 $Y2=0
cc_965 N_A_1586_74#_c_1150_n N_A_1784_97#_M1035_d 0.0043242f $X=8.89 $Y=1.82
+ $X2=-0.19 $Y2=-0.245
cc_966 N_A_1586_74#_c_1141_n N_A_1784_97#_M1018_g 0.00576525f $X=10.69 $Y=0.935
+ $X2=0 $Y2=0
cc_967 N_A_1586_74#_c_1237_p N_A_1784_97#_M1018_g 0.0116034f $X=10.775 $Y=0.85
+ $X2=0 $Y2=0
cc_968 N_A_1586_74#_c_1142_n N_A_1784_97#_M1018_g 0.0112842f $X=11.37 $Y=0.34
+ $X2=0 $Y2=0
cc_969 N_A_1586_74#_c_1143_n N_A_1784_97#_M1018_g 0.00332344f $X=10.86 $Y=0.34
+ $X2=0 $Y2=0
cc_970 N_A_1586_74#_c_1144_n N_A_1784_97#_M1018_g 0.00327684f $X=11.455 $Y=0.85
+ $X2=0 $Y2=0
cc_971 N_A_1586_74#_c_1131_n N_A_1784_97#_c_1668_n 0.00497183f $X=9.525 $Y=1.015
+ $X2=0 $Y2=0
cc_972 N_A_1586_74#_c_1137_n N_A_1784_97#_c_1668_n 0.012971f $X=9.565 $Y=0.34
+ $X2=0 $Y2=0
cc_973 N_A_1586_74#_c_1139_n N_A_1784_97#_c_1668_n 0.0241468f $X=9.69 $Y=1.18
+ $X2=0 $Y2=0
cc_974 N_A_1586_74#_c_1150_n N_A_1784_97#_c_1668_n 0.0805264f $X=8.89 $Y=1.82
+ $X2=0 $Y2=0
cc_975 N_A_1586_74#_c_1275_p N_A_1784_97#_c_1668_n 0.0114261f $X=9.71 $Y=0.935
+ $X2=0 $Y2=0
cc_976 N_A_1586_74#_c_1139_n N_A_1784_97#_c_1671_n 0.0087019f $X=9.69 $Y=1.18
+ $X2=0 $Y2=0
cc_977 N_A_1586_74#_c_1140_n N_A_1784_97#_c_1671_n 0.00188502f $X=9.69 $Y=1.18
+ $X2=0 $Y2=0
cc_978 N_A_1586_74#_c_1141_n N_A_1784_97#_c_1671_n 0.00312506f $X=10.69 $Y=0.935
+ $X2=0 $Y2=0
cc_979 N_A_1586_74#_c_1150_n N_A_1784_97#_c_1672_n 0.0136362f $X=8.89 $Y=1.82
+ $X2=0 $Y2=0
cc_980 N_A_1586_74#_M1015_g N_A_1784_97#_c_1673_n 0.0074834f $X=9.195 $Y=2.75
+ $X2=0 $Y2=0
cc_981 N_A_1586_74#_M1015_g N_A_1784_97#_c_1674_n 0.00959071f $X=9.195 $Y=2.75
+ $X2=0 $Y2=0
cc_982 N_A_1586_74#_c_1159_n N_A_1784_97#_c_1674_n 0.0333201f $X=8.89 $Y=1.98
+ $X2=0 $Y2=0
cc_983 N_A_1586_74#_c_1161_n N_A_1784_97#_c_1674_n 0.00616979f $X=8.89 $Y=2.14
+ $X2=0 $Y2=0
cc_984 N_A_1586_74#_M1010_g N_A_2489_74#_c_1833_n 0.00274767f $X=12.37 $Y=0.69
+ $X2=0 $Y2=0
cc_985 N_A_1586_74#_c_1149_n N_A_2489_74#_c_1833_n 0.0224089f $X=13.195 $Y=1.215
+ $X2=0 $Y2=0
cc_986 N_A_1586_74#_M1010_g N_A_2489_74#_c_1763_n 0.00726238f $X=12.37 $Y=0.69
+ $X2=0 $Y2=0
cc_987 N_A_1586_74#_c_1149_n N_A_2489_74#_c_1764_n 0.0298078f $X=13.195 $Y=1.215
+ $X2=0 $Y2=0
cc_988 N_A_1586_74#_c_1152_n N_A_2489_74#_c_1764_n 0.0233024f $X=13.36 $Y=1.215
+ $X2=0 $Y2=0
cc_989 N_A_1586_74#_c_1153_n N_A_2489_74#_c_1764_n 3.05108e-19 $X=13.36 $Y=1.39
+ $X2=0 $Y2=0
cc_990 N_A_1586_74#_M1030_g N_A_2489_74#_c_1772_n 0.0190596f $X=13.285 $Y=2.75
+ $X2=0 $Y2=0
cc_991 N_A_1586_74#_M1030_g N_A_2489_74#_c_1773_n 0.00549922f $X=13.285 $Y=2.75
+ $X2=0 $Y2=0
cc_992 N_A_1586_74#_c_1152_n N_A_2489_74#_c_1773_n 0.0129484f $X=13.36 $Y=1.215
+ $X2=0 $Y2=0
cc_993 N_A_1586_74#_c_1153_n N_A_2489_74#_c_1773_n 0.00334366f $X=13.36 $Y=1.39
+ $X2=0 $Y2=0
cc_994 N_A_1586_74#_M1030_g N_A_2489_74#_c_1774_n 0.00374558f $X=13.285 $Y=2.75
+ $X2=0 $Y2=0
cc_995 N_A_1586_74#_c_1149_n N_A_2489_74#_c_1774_n 0.00104657f $X=13.195
+ $Y=1.215 $X2=0 $Y2=0
cc_996 N_A_1586_74#_c_1152_n N_A_2489_74#_c_1774_n 0.00824827f $X=13.36 $Y=1.215
+ $X2=0 $Y2=0
cc_997 N_A_1586_74#_c_1152_n N_A_2489_74#_c_1765_n 0.0315436f $X=13.36 $Y=1.215
+ $X2=0 $Y2=0
cc_998 N_A_1586_74#_c_1153_n N_A_2489_74#_c_1765_n 0.00202138f $X=13.36 $Y=1.39
+ $X2=0 $Y2=0
cc_999 N_A_1586_74#_M1030_g N_A_2489_74#_c_1766_n 0.00242749f $X=13.285 $Y=2.75
+ $X2=0 $Y2=0
cc_1000 N_A_1586_74#_M1030_g N_A_2489_74#_c_1776_n 0.0184909f $X=13.285 $Y=2.75
+ $X2=0 $Y2=0
cc_1001 N_A_1586_74#_M1030_g N_VPWR_c_2031_n 0.00143219f $X=13.285 $Y=2.75 $X2=0
+ $Y2=0
cc_1002 N_A_1586_74#_M1015_g N_VPWR_c_2044_n 0.0048691f $X=9.195 $Y=2.75 $X2=0
+ $Y2=0
cc_1003 N_A_1586_74#_M1030_g N_VPWR_c_2045_n 0.00406584f $X=13.285 $Y=2.75 $X2=0
+ $Y2=0
cc_1004 N_A_1586_74#_M1015_g N_VPWR_c_2023_n 0.00878547f $X=9.195 $Y=2.75 $X2=0
+ $Y2=0
cc_1005 N_A_1586_74#_M1030_g N_VPWR_c_2023_n 0.00612649f $X=13.285 $Y=2.75 $X2=0
+ $Y2=0
cc_1006 N_A_1586_74#_c_1157_n N_A_691_113#_c_2238_n 0.013384f $X=8.725 $Y=1.98
+ $X2=0 $Y2=0
cc_1007 N_A_1586_74#_c_1159_n N_A_691_113#_c_2238_n 0.00206609f $X=8.89 $Y=1.98
+ $X2=0 $Y2=0
cc_1008 N_A_1586_74#_c_1134_n N_A_691_113#_c_2225_n 0.00680159f $X=8.07 $Y=0.515
+ $X2=0 $Y2=0
cc_1009 N_A_1586_74#_c_1157_n N_A_691_113#_c_2225_n 0.0305951f $X=8.725 $Y=1.98
+ $X2=0 $Y2=0
cc_1010 N_A_1586_74#_c_1150_n N_A_691_113#_c_2225_n 0.0128117f $X=8.89 $Y=1.82
+ $X2=0 $Y2=0
cc_1011 N_A_1586_74#_c_1134_n N_A_691_113#_c_2226_n 0.00798758f $X=8.07 $Y=0.515
+ $X2=0 $Y2=0
cc_1012 N_A_1586_74#_c_1157_n N_A_691_113#_c_2252_n 0.0020452f $X=8.725 $Y=1.98
+ $X2=0 $Y2=0
cc_1013 N_A_1586_74#_c_1134_n N_A_691_113#_c_2227_n 0.0353265f $X=8.07 $Y=0.515
+ $X2=0 $Y2=0
cc_1014 N_A_1586_74#_c_1135_n N_A_691_113#_c_2227_n 0.0191962f $X=8.885 $Y=0.34
+ $X2=0 $Y2=0
cc_1015 N_A_1586_74#_c_1150_n N_A_691_113#_c_2227_n 0.0528515f $X=8.89 $Y=1.82
+ $X2=0 $Y2=0
cc_1016 N_A_1586_74#_M1008_d N_A_691_113#_c_2239_n 0.00421794f $X=8.275 $Y=1.84
+ $X2=0 $Y2=0
cc_1017 N_A_1586_74#_M1015_g N_A_691_113#_c_2239_n 0.00172768f $X=9.195 $Y=2.75
+ $X2=0 $Y2=0
cc_1018 N_A_1586_74#_c_1157_n N_A_691_113#_c_2239_n 0.0124469f $X=8.725 $Y=1.98
+ $X2=0 $Y2=0
cc_1019 N_A_1586_74#_c_1159_n N_A_691_113#_c_2239_n 0.0270109f $X=8.89 $Y=1.98
+ $X2=0 $Y2=0
cc_1020 N_A_1586_74#_c_1161_n N_A_691_113#_c_2239_n 0.00245339f $X=8.89 $Y=2.14
+ $X2=0 $Y2=0
cc_1021 N_A_1586_74#_M1015_g N_A_691_113#_c_2240_n 7.6107e-19 $X=9.195 $Y=2.75
+ $X2=0 $Y2=0
cc_1022 N_A_1586_74#_M1008_d N_A_691_113#_c_2329_n 0.00738599f $X=8.275 $Y=1.84
+ $X2=0 $Y2=0
cc_1023 N_A_1586_74#_M1015_g N_A_691_113#_c_2329_n 0.0036778f $X=9.195 $Y=2.75
+ $X2=0 $Y2=0
cc_1024 N_A_1586_74#_c_1157_n N_A_691_113#_c_2329_n 0.0103555f $X=8.725 $Y=1.98
+ $X2=0 $Y2=0
cc_1025 N_A_1586_74#_c_1141_n N_VGND_M1025_d 0.00719284f $X=10.69 $Y=0.935 $X2=0
+ $Y2=0
cc_1026 N_A_1586_74#_c_1237_p N_VGND_M1025_d 0.00493253f $X=10.775 $Y=0.85 $X2=0
+ $Y2=0
cc_1027 N_A_1586_74#_c_1143_n N_VGND_M1025_d 5.37788e-19 $X=10.86 $Y=0.34 $X2=0
+ $Y2=0
cc_1028 N_A_1586_74#_c_1145_n N_VGND_M1007_s 0.00391333f $X=12.08 $Y=0.935 $X2=0
+ $Y2=0
cc_1029 N_A_1586_74#_c_1134_n N_VGND_c_2465_n 0.0259189f $X=8.07 $Y=0.515 $X2=0
+ $Y2=0
cc_1030 N_A_1586_74#_c_1136_n N_VGND_c_2465_n 0.010974f $X=8.235 $Y=0.34 $X2=0
+ $Y2=0
cc_1031 N_A_1586_74#_c_1137_n N_VGND_c_2466_n 0.00662337f $X=9.565 $Y=0.34 $X2=0
+ $Y2=0
cc_1032 N_A_1586_74#_c_1138_n N_VGND_c_2466_n 0.00506803f $X=9.65 $Y=0.85 $X2=0
+ $Y2=0
cc_1033 N_A_1586_74#_c_1141_n N_VGND_c_2466_n 0.0196718f $X=10.69 $Y=0.935 $X2=0
+ $Y2=0
cc_1034 N_A_1586_74#_c_1237_p N_VGND_c_2466_n 0.0190358f $X=10.775 $Y=0.85 $X2=0
+ $Y2=0
cc_1035 N_A_1586_74#_c_1143_n N_VGND_c_2466_n 0.0145685f $X=10.86 $Y=0.34 $X2=0
+ $Y2=0
cc_1036 N_A_1586_74#_M1010_g N_VGND_c_2467_n 0.00147043f $X=12.37 $Y=0.69 $X2=0
+ $Y2=0
cc_1037 N_A_1586_74#_c_1142_n N_VGND_c_2467_n 0.0146661f $X=11.37 $Y=0.34 $X2=0
+ $Y2=0
cc_1038 N_A_1586_74#_c_1144_n N_VGND_c_2467_n 0.0193741f $X=11.455 $Y=0.85 $X2=0
+ $Y2=0
cc_1039 N_A_1586_74#_c_1145_n N_VGND_c_2467_n 0.015048f $X=12.08 $Y=0.935 $X2=0
+ $Y2=0
cc_1040 N_A_1586_74#_M1010_g N_VGND_c_2481_n 0.00434272f $X=12.37 $Y=0.69 $X2=0
+ $Y2=0
cc_1041 N_A_1586_74#_c_1131_n N_VGND_c_2485_n 7.53287e-19 $X=9.525 $Y=1.015
+ $X2=0 $Y2=0
cc_1042 N_A_1586_74#_c_1135_n N_VGND_c_2485_n 0.0418136f $X=8.885 $Y=0.34 $X2=0
+ $Y2=0
cc_1043 N_A_1586_74#_c_1136_n N_VGND_c_2485_n 0.0235688f $X=8.235 $Y=0.34 $X2=0
+ $Y2=0
cc_1044 N_A_1586_74#_c_1137_n N_VGND_c_2485_n 0.0449818f $X=9.565 $Y=0.34 $X2=0
+ $Y2=0
cc_1045 N_A_1586_74#_c_1151_n N_VGND_c_2485_n 0.0121867f $X=8.97 $Y=0.34 $X2=0
+ $Y2=0
cc_1046 N_A_1586_74#_c_1142_n N_VGND_c_2486_n 0.0446499f $X=11.37 $Y=0.34 $X2=0
+ $Y2=0
cc_1047 N_A_1586_74#_c_1143_n N_VGND_c_2486_n 0.0120637f $X=10.86 $Y=0.34 $X2=0
+ $Y2=0
cc_1048 N_A_1586_74#_M1010_g N_VGND_c_2496_n 0.00821463f $X=12.37 $Y=0.69 $X2=0
+ $Y2=0
cc_1049 N_A_1586_74#_c_1135_n N_VGND_c_2496_n 0.0244305f $X=8.885 $Y=0.34 $X2=0
+ $Y2=0
cc_1050 N_A_1586_74#_c_1136_n N_VGND_c_2496_n 0.0127152f $X=8.235 $Y=0.34 $X2=0
+ $Y2=0
cc_1051 N_A_1586_74#_c_1137_n N_VGND_c_2496_n 0.025776f $X=9.565 $Y=0.34 $X2=0
+ $Y2=0
cc_1052 N_A_1586_74#_c_1141_n N_VGND_c_2496_n 0.0203559f $X=10.69 $Y=0.935 $X2=0
+ $Y2=0
cc_1053 N_A_1586_74#_c_1142_n N_VGND_c_2496_n 0.0252533f $X=11.37 $Y=0.34 $X2=0
+ $Y2=0
cc_1054 N_A_1586_74#_c_1143_n N_VGND_c_2496_n 0.00644906f $X=10.86 $Y=0.34 $X2=0
+ $Y2=0
cc_1055 N_A_1586_74#_c_1145_n N_VGND_c_2496_n 0.00988673f $X=12.08 $Y=0.935
+ $X2=0 $Y2=0
cc_1056 N_A_1586_74#_c_1147_n N_VGND_c_2496_n 0.00660638f $X=12.23 $Y=1.3 $X2=0
+ $Y2=0
cc_1057 N_A_1586_74#_c_1151_n N_VGND_c_2496_n 0.00660921f $X=8.97 $Y=0.34 $X2=0
+ $Y2=0
cc_1058 N_A_1586_74#_c_1275_p N_VGND_c_2496_n 0.00454674f $X=9.71 $Y=0.935 $X2=0
+ $Y2=0
cc_1059 N_A_1586_74#_c_1138_n A_1920_97# 0.00506914f $X=9.65 $Y=0.85 $X2=-0.19
+ $Y2=-0.245
cc_1060 N_A_1586_74#_c_1141_n A_1920_97# 0.00308187f $X=10.69 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_1061 N_A_1586_74#_c_1275_p A_1920_97# 0.00274383f $X=9.71 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_1062 N_A_1586_74#_c_1147_n A_2417_74# 0.00229931f $X=12.23 $Y=1.3 $X2=-0.19
+ $Y2=-0.245
cc_1063 N_A_1377_368#_c_1386_n N_A_2013_71#_M1032_d 0.0073881f $X=12.55 $Y=2.475
+ $X2=0 $Y2=0
cc_1064 N_A_1377_368#_c_1367_n N_A_2013_71#_M1016_g 0.014422f $X=9.525 $Y=1.66
+ $X2=0 $Y2=0
cc_1065 N_A_1377_368#_M1019_g N_A_2013_71#_M1016_g 0.0261968f $X=9.645 $Y=2.75
+ $X2=0 $Y2=0
cc_1066 N_A_1377_368#_c_1386_n N_A_2013_71#_M1016_g 0.0155462f $X=12.55 $Y=2.475
+ $X2=0 $Y2=0
cc_1067 N_A_1377_368#_c_1390_n N_A_2013_71#_M1016_g 0.00865029f $X=9.69 $Y=2.195
+ $X2=0 $Y2=0
cc_1068 N_A_1377_368#_c_1391_n N_A_2013_71#_M1016_g 0.0196783f $X=9.69 $Y=2.195
+ $X2=0 $Y2=0
cc_1069 N_A_1377_368#_c_1386_n N_A_2013_71#_M1043_g 0.0228105f $X=12.55 $Y=2.475
+ $X2=0 $Y2=0
cc_1070 N_A_1377_368#_c_1387_n N_A_2013_71#_M1043_g 0.0123694f $X=12.635 $Y=2.39
+ $X2=0 $Y2=0
cc_1071 N_A_1377_368#_c_1386_n N_A_2013_71#_c_1569_n 0.0432049f $X=12.55
+ $Y=2.475 $X2=0 $Y2=0
cc_1072 N_A_1377_368#_c_1386_n N_A_1784_97#_M1032_g 0.0173005f $X=12.55 $Y=2.475
+ $X2=0 $Y2=0
cc_1073 N_A_1377_368#_M1035_g N_A_1784_97#_c_1668_n 0.00328193f $X=8.845
+ $Y=0.695 $X2=0 $Y2=0
cc_1074 N_A_1377_368#_c_1367_n N_A_1784_97#_c_1668_n 0.00874168f $X=9.525
+ $Y=1.66 $X2=0 $Y2=0
cc_1075 N_A_1377_368#_c_1367_n N_A_1784_97#_c_1671_n 0.00645603f $X=9.525
+ $Y=1.66 $X2=0 $Y2=0
cc_1076 N_A_1377_368#_c_1386_n N_A_1784_97#_c_1671_n 0.0208227f $X=12.55
+ $Y=2.475 $X2=0 $Y2=0
cc_1077 N_A_1377_368#_c_1390_n N_A_1784_97#_c_1671_n 0.025582f $X=9.69 $Y=2.195
+ $X2=0 $Y2=0
cc_1078 N_A_1377_368#_c_1391_n N_A_1784_97#_c_1671_n 7.5533e-19 $X=9.69 $Y=2.195
+ $X2=0 $Y2=0
cc_1079 N_A_1377_368#_c_1395_n N_A_1784_97#_c_1671_n 0.00862473f $X=9.69 $Y=2.03
+ $X2=0 $Y2=0
cc_1080 N_A_1377_368#_c_1367_n N_A_1784_97#_c_1672_n 0.00465441f $X=9.525
+ $Y=1.66 $X2=0 $Y2=0
cc_1081 N_A_1377_368#_M1019_g N_A_1784_97#_c_1673_n 0.0104187f $X=9.645 $Y=2.75
+ $X2=0 $Y2=0
cc_1082 N_A_1377_368#_c_1390_n N_A_1784_97#_c_1673_n 0.00304136f $X=9.69
+ $Y=2.195 $X2=0 $Y2=0
cc_1083 N_A_1377_368#_c_1391_n N_A_1784_97#_c_1673_n 9.93333e-19 $X=9.69
+ $Y=2.195 $X2=0 $Y2=0
cc_1084 N_A_1377_368#_M1019_g N_A_1784_97#_c_1674_n 0.00131924f $X=9.645 $Y=2.75
+ $X2=0 $Y2=0
cc_1085 N_A_1377_368#_c_1390_n N_A_1784_97#_c_1674_n 0.0334054f $X=9.69 $Y=2.195
+ $X2=0 $Y2=0
cc_1086 N_A_1377_368#_c_1395_n N_A_1784_97#_c_1674_n 0.00778971f $X=9.69 $Y=2.03
+ $X2=0 $Y2=0
cc_1087 N_A_1377_368#_c_1386_n N_A_1784_97#_c_1675_n 0.00420338f $X=12.55
+ $Y=2.475 $X2=0 $Y2=0
cc_1088 N_A_1377_368#_M1011_g N_A_2489_74#_c_1763_n 0.00236994f $X=12.88 $Y=0.58
+ $X2=0 $Y2=0
cc_1089 N_A_1377_368#_M1011_g N_A_2489_74#_c_1764_n 0.0118688f $X=12.88 $Y=0.58
+ $X2=0 $Y2=0
cc_1090 N_A_1377_368#_M1034_g N_A_2489_74#_c_1772_n 0.00452582f $X=12.75 $Y=2.46
+ $X2=0 $Y2=0
cc_1091 N_A_1377_368#_c_1386_n N_A_2489_74#_c_1772_n 0.00510983f $X=12.55
+ $Y=2.475 $X2=0 $Y2=0
cc_1092 N_A_1377_368#_c_1387_n N_A_2489_74#_c_1772_n 0.0178812f $X=12.635
+ $Y=2.39 $X2=0 $Y2=0
cc_1093 N_A_1377_368#_M1034_g N_A_2489_74#_c_1774_n 7.04126e-19 $X=12.75 $Y=2.46
+ $X2=0 $Y2=0
cc_1094 N_A_1377_368#_c_1387_n N_A_2489_74#_c_1774_n 0.00332661f $X=12.635
+ $Y=2.39 $X2=0 $Y2=0
cc_1095 N_A_1377_368#_c_1374_n N_A_2489_74#_c_1774_n 0.00682912f $X=12.82
+ $Y=1.635 $X2=0 $Y2=0
cc_1096 N_A_1377_368#_c_1375_n N_A_2489_74#_c_1774_n 2.83747e-19 $X=12.82
+ $Y=1.635 $X2=0 $Y2=0
cc_1097 N_A_1377_368#_M1034_g N_A_2489_74#_c_1776_n 8.13469e-19 $X=12.75 $Y=2.46
+ $X2=0 $Y2=0
cc_1098 N_A_1377_368#_c_1386_n N_VPWR_M1016_d 0.00625831f $X=12.55 $Y=2.475
+ $X2=0 $Y2=0
cc_1099 N_A_1377_368#_c_1386_n N_VPWR_M1043_s 0.0154325f $X=12.55 $Y=2.475 $X2=0
+ $Y2=0
cc_1100 N_A_1377_368#_c_1378_n N_VPWR_c_2028_n 0.0229156f $X=8.185 $Y=1.735
+ $X2=0 $Y2=0
cc_1101 N_A_1377_368#_M1019_g N_VPWR_c_2029_n 0.00126439f $X=9.645 $Y=2.75 $X2=0
+ $Y2=0
cc_1102 N_A_1377_368#_c_1386_n N_VPWR_c_2029_n 0.021216f $X=12.55 $Y=2.475 $X2=0
+ $Y2=0
cc_1103 N_A_1377_368#_c_1386_n N_VPWR_c_2030_n 0.0259191f $X=12.55 $Y=2.475
+ $X2=0 $Y2=0
cc_1104 N_A_1377_368#_c_1378_n N_VPWR_c_2044_n 0.00460063f $X=8.185 $Y=1.735
+ $X2=0 $Y2=0
cc_1105 N_A_1377_368#_M1019_g N_VPWR_c_2044_n 0.005209f $X=9.645 $Y=2.75 $X2=0
+ $Y2=0
cc_1106 N_A_1377_368#_M1034_g N_VPWR_c_2045_n 0.00553757f $X=12.75 $Y=2.46 $X2=0
+ $Y2=0
cc_1107 N_A_1377_368#_c_1378_n N_VPWR_c_2023_n 0.00468499f $X=8.185 $Y=1.735
+ $X2=0 $Y2=0
cc_1108 N_A_1377_368#_M1019_g N_VPWR_c_2023_n 0.00984127f $X=9.645 $Y=2.75 $X2=0
+ $Y2=0
cc_1109 N_A_1377_368#_M1034_g N_VPWR_c_2023_n 0.00910759f $X=12.75 $Y=2.46 $X2=0
+ $Y2=0
cc_1110 N_A_1377_368#_c_1386_n N_VPWR_c_2023_n 0.0781996f $X=12.55 $Y=2.475
+ $X2=0 $Y2=0
cc_1111 N_A_1377_368#_c_1390_n N_VPWR_c_2023_n 0.00695798f $X=9.69 $Y=2.195
+ $X2=0 $Y2=0
cc_1112 N_A_1377_368#_c_1385_n N_A_691_113#_c_2224_n 0.0127786f $X=7.215 $Y=1.98
+ $X2=0 $Y2=0
cc_1113 N_A_1377_368#_M1000_d N_A_691_113#_c_2236_n 0.00778164f $X=6.885 $Y=1.84
+ $X2=0 $Y2=0
cc_1114 N_A_1377_368#_c_1385_n N_A_691_113#_c_2236_n 0.0224655f $X=7.215 $Y=1.98
+ $X2=0 $Y2=0
cc_1115 N_A_1377_368#_c_1372_n N_A_691_113#_c_2236_n 0.0346f $X=7.49 $Y=1.635
+ $X2=0 $Y2=0
cc_1116 N_A_1377_368#_c_1389_n N_A_691_113#_c_2236_n 0.00229113f $X=7.49
+ $Y=1.635 $X2=0 $Y2=0
cc_1117 N_A_1377_368#_c_1376_n N_A_691_113#_c_2236_n 0.00305541f $X=7.93
+ $Y=1.602 $X2=0 $Y2=0
cc_1118 N_A_1377_368#_c_1364_n N_A_691_113#_c_2238_n 0.00501137f $X=8.095
+ $Y=1.66 $X2=0 $Y2=0
cc_1119 N_A_1377_368#_c_1378_n N_A_691_113#_c_2238_n 0.00812288f $X=8.185
+ $Y=1.735 $X2=0 $Y2=0
cc_1120 N_A_1377_368#_c_1372_n N_A_691_113#_c_2238_n 0.0264305f $X=7.49 $Y=1.635
+ $X2=0 $Y2=0
cc_1121 N_A_1377_368#_c_1389_n N_A_691_113#_c_2238_n 0.00314109f $X=7.49
+ $Y=1.635 $X2=0 $Y2=0
cc_1122 N_A_1377_368#_c_1376_n N_A_691_113#_c_2238_n 0.00171162f $X=7.93
+ $Y=1.602 $X2=0 $Y2=0
cc_1123 N_A_1377_368#_c_1364_n N_A_691_113#_c_2225_n 7.62721e-19 $X=8.095
+ $Y=1.66 $X2=0 $Y2=0
cc_1124 N_A_1377_368#_c_1365_n N_A_691_113#_c_2225_n 0.0133058f $X=8.77 $Y=1.66
+ $X2=0 $Y2=0
cc_1125 N_A_1377_368#_M1035_g N_A_691_113#_c_2225_n 0.00239961f $X=8.845
+ $Y=0.695 $X2=0 $Y2=0
cc_1126 N_A_1377_368#_c_1369_n N_A_691_113#_c_2225_n 0.00725359f $X=8.185
+ $Y=1.66 $X2=0 $Y2=0
cc_1127 N_A_1377_368#_c_1364_n N_A_691_113#_c_2226_n 0.00178115f $X=8.095
+ $Y=1.66 $X2=0 $Y2=0
cc_1128 N_A_1377_368#_c_1372_n N_A_691_113#_c_2226_n 0.00922738f $X=7.49
+ $Y=1.635 $X2=0 $Y2=0
cc_1129 N_A_1377_368#_c_1376_n N_A_691_113#_c_2226_n 0.00619128f $X=7.93
+ $Y=1.602 $X2=0 $Y2=0
cc_1130 N_A_1377_368#_c_1378_n N_A_691_113#_c_2252_n 0.0177608f $X=8.185
+ $Y=1.735 $X2=0 $Y2=0
cc_1131 N_A_1377_368#_M1004_g N_A_691_113#_c_2227_n 0.00963337f $X=7.855 $Y=0.74
+ $X2=0 $Y2=0
cc_1132 N_A_1377_368#_M1035_g N_A_691_113#_c_2227_n 0.0127542f $X=8.845 $Y=0.695
+ $X2=0 $Y2=0
cc_1133 N_A_1377_368#_c_1378_n N_A_691_113#_c_2240_n 0.00826897f $X=8.185
+ $Y=1.735 $X2=0 $Y2=0
cc_1134 N_A_1377_368#_c_1386_n A_1947_508# 0.00154876f $X=12.55 $Y=2.475
+ $X2=-0.19 $Y2=-0.245
cc_1135 N_A_1377_368#_c_1390_n A_1947_508# 0.00298282f $X=9.69 $Y=2.195
+ $X2=-0.19 $Y2=-0.245
cc_1136 N_A_1377_368#_c_1386_n A_2377_392# 0.0319474f $X=12.55 $Y=2.475
+ $X2=-0.19 $Y2=-0.245
cc_1137 N_A_1377_368#_c_1387_n A_2377_392# 0.00757088f $X=12.635 $Y=2.39
+ $X2=-0.19 $Y2=-0.245
cc_1138 N_A_1377_368#_c_1371_n N_VGND_c_2464_n 0.023367f $X=7.08 $Y=0.515 $X2=0
+ $Y2=0
cc_1139 N_A_1377_368#_M1004_g N_VGND_c_2465_n 0.00467695f $X=7.855 $Y=0.74 $X2=0
+ $Y2=0
cc_1140 N_A_1377_368#_c_1371_n N_VGND_c_2465_n 0.0618465f $X=7.08 $Y=0.515 $X2=0
+ $Y2=0
cc_1141 N_A_1377_368#_c_1372_n N_VGND_c_2465_n 0.00440058f $X=7.49 $Y=1.635
+ $X2=0 $Y2=0
cc_1142 N_A_1377_368#_c_1376_n N_VGND_c_2465_n 0.00353088f $X=7.93 $Y=1.602
+ $X2=0 $Y2=0
cc_1143 N_A_1377_368#_M1011_g N_VGND_c_2469_n 0.00128745f $X=12.88 $Y=0.58 $X2=0
+ $Y2=0
cc_1144 N_A_1377_368#_c_1371_n N_VGND_c_2479_n 0.0207821f $X=7.08 $Y=0.515 $X2=0
+ $Y2=0
cc_1145 N_A_1377_368#_M1011_g N_VGND_c_2481_n 0.00461464f $X=12.88 $Y=0.58 $X2=0
+ $Y2=0
cc_1146 N_A_1377_368#_M1004_g N_VGND_c_2485_n 0.00430908f $X=7.855 $Y=0.74 $X2=0
+ $Y2=0
cc_1147 N_A_1377_368#_M1035_g N_VGND_c_2485_n 7.53287e-19 $X=8.845 $Y=0.695
+ $X2=0 $Y2=0
cc_1148 N_A_1377_368#_M1004_g N_VGND_c_2496_n 0.0082568f $X=7.855 $Y=0.74 $X2=0
+ $Y2=0
cc_1149 N_A_1377_368#_M1011_g N_VGND_c_2496_n 0.00447595f $X=12.88 $Y=0.58 $X2=0
+ $Y2=0
cc_1150 N_A_1377_368#_c_1371_n N_VGND_c_2496_n 0.0171578f $X=7.08 $Y=0.515 $X2=0
+ $Y2=0
cc_1151 N_A_2013_71#_c_1569_n N_A_1784_97#_M1032_g 0.00449958f $X=11.215
+ $Y=2.135 $X2=0 $Y2=0
cc_1152 N_A_2013_71#_c_1561_n N_A_1784_97#_M1032_g 0.00439318f $X=11.3 $Y=2.05
+ $X2=0 $Y2=0
cc_1153 N_A_2013_71#_M1025_g N_A_1784_97#_M1018_g 0.0125129f $X=10.14 $Y=0.695
+ $X2=0 $Y2=0
cc_1154 N_A_2013_71#_c_1559_n N_A_1784_97#_M1018_g 0.0144178f $X=11.03 $Y=1.275
+ $X2=0 $Y2=0
cc_1155 N_A_2013_71#_c_1560_n N_A_1784_97#_M1018_g 0.00603479f $X=11.115
+ $Y=0.805 $X2=0 $Y2=0
cc_1156 N_A_2013_71#_c_1562_n N_A_1784_97#_M1018_g 0.0010369f $X=11.385 $Y=1.355
+ $X2=0 $Y2=0
cc_1157 N_A_2013_71#_c_1564_n N_A_1784_97#_M1018_g 0.0214312f $X=11.72 $Y=1.355
+ $X2=0 $Y2=0
cc_1158 N_A_2013_71#_c_1565_n N_A_1784_97#_M1018_g 8.94976e-19 $X=10.23 $Y=1.275
+ $X2=0 $Y2=0
cc_1159 N_A_2013_71#_c_1566_n N_A_1784_97#_M1018_g 0.00852329f $X=10.23 $Y=1.355
+ $X2=0 $Y2=0
cc_1160 N_A_2013_71#_M1025_g N_A_1784_97#_c_1668_n 0.00400396f $X=10.14 $Y=0.695
+ $X2=0 $Y2=0
cc_1161 N_A_2013_71#_M1016_g N_A_1784_97#_c_1668_n 4.86365e-19 $X=10.155 $Y=2.75
+ $X2=0 $Y2=0
cc_1162 N_A_2013_71#_c_1565_n N_A_1784_97#_c_1668_n 0.00461219f $X=10.23
+ $Y=1.275 $X2=0 $Y2=0
cc_1163 N_A_2013_71#_M1016_g N_A_1784_97#_c_1671_n 0.0137448f $X=10.155 $Y=2.75
+ $X2=0 $Y2=0
cc_1164 N_A_2013_71#_c_1559_n N_A_1784_97#_c_1671_n 0.00704001f $X=11.03
+ $Y=1.275 $X2=0 $Y2=0
cc_1165 N_A_2013_71#_c_1565_n N_A_1784_97#_c_1671_n 0.0208348f $X=10.23 $Y=1.275
+ $X2=0 $Y2=0
cc_1166 N_A_2013_71#_c_1566_n N_A_1784_97#_c_1671_n 9.81093e-19 $X=10.23
+ $Y=1.355 $X2=0 $Y2=0
cc_1167 N_A_2013_71#_M1016_g N_A_1784_97#_c_1673_n 0.00157631f $X=10.155 $Y=2.75
+ $X2=0 $Y2=0
cc_1168 N_A_2013_71#_M1016_g N_A_1784_97#_c_1675_n 0.001345f $X=10.155 $Y=2.75
+ $X2=0 $Y2=0
cc_1169 N_A_2013_71#_c_1559_n N_A_1784_97#_c_1675_n 0.0224081f $X=11.03 $Y=1.275
+ $X2=0 $Y2=0
cc_1170 N_A_2013_71#_c_1569_n N_A_1784_97#_c_1675_n 0.0101481f $X=11.215
+ $Y=2.135 $X2=0 $Y2=0
cc_1171 N_A_2013_71#_c_1561_n N_A_1784_97#_c_1675_n 0.0158264f $X=11.3 $Y=2.05
+ $X2=0 $Y2=0
cc_1172 N_A_2013_71#_M1016_g N_A_1784_97#_c_1669_n 0.0442614f $X=10.155 $Y=2.75
+ $X2=0 $Y2=0
cc_1173 N_A_2013_71#_c_1559_n N_A_1784_97#_c_1669_n 0.00573884f $X=11.03
+ $Y=1.275 $X2=0 $Y2=0
cc_1174 N_A_2013_71#_c_1569_n N_A_1784_97#_c_1669_n 0.00222911f $X=11.215
+ $Y=2.135 $X2=0 $Y2=0
cc_1175 N_A_2013_71#_c_1561_n N_A_1784_97#_c_1669_n 0.00605217f $X=11.3 $Y=2.05
+ $X2=0 $Y2=0
cc_1176 N_A_2013_71#_c_1566_n N_A_1784_97#_c_1669_n 0.00132858f $X=10.23
+ $Y=1.355 $X2=0 $Y2=0
cc_1177 N_A_2013_71#_c_1558_n N_A_2489_74#_c_1833_n 4.65641e-19 $X=12.01 $Y=1.11
+ $X2=0 $Y2=0
cc_1178 N_A_2013_71#_c_1558_n N_A_2489_74#_c_1763_n 0.00134647f $X=12.01 $Y=1.11
+ $X2=0 $Y2=0
cc_1179 N_A_2013_71#_c_1569_n N_VPWR_M1043_s 0.00348329f $X=11.215 $Y=2.135
+ $X2=0 $Y2=0
cc_1180 N_A_2013_71#_c_1561_n N_VPWR_M1043_s 0.00138186f $X=11.3 $Y=2.05 $X2=0
+ $Y2=0
cc_1181 N_A_2013_71#_M1016_g N_VPWR_c_2029_n 0.0103698f $X=10.155 $Y=2.75 $X2=0
+ $Y2=0
cc_1182 N_A_2013_71#_M1043_g N_VPWR_c_2030_n 0.0101031f $X=11.795 $Y=2.46 $X2=0
+ $Y2=0
cc_1183 N_A_2013_71#_M1016_g N_VPWR_c_2044_n 0.00490827f $X=10.155 $Y=2.75 $X2=0
+ $Y2=0
cc_1184 N_A_2013_71#_M1043_g N_VPWR_c_2045_n 0.00553757f $X=11.795 $Y=2.46 $X2=0
+ $Y2=0
cc_1185 N_A_2013_71#_M1016_g N_VPWR_c_2023_n 0.00473297f $X=10.155 $Y=2.75 $X2=0
+ $Y2=0
cc_1186 N_A_2013_71#_M1043_g N_VPWR_c_2023_n 0.00544364f $X=11.795 $Y=2.46 $X2=0
+ $Y2=0
cc_1187 N_A_2013_71#_M1025_g N_VGND_c_2466_n 0.00364778f $X=10.14 $Y=0.695 $X2=0
+ $Y2=0
cc_1188 N_A_2013_71#_c_1558_n N_VGND_c_2467_n 0.010393f $X=12.01 $Y=1.11 $X2=0
+ $Y2=0
cc_1189 N_A_2013_71#_c_1558_n N_VGND_c_2481_n 0.00383152f $X=12.01 $Y=1.11 $X2=0
+ $Y2=0
cc_1190 N_A_2013_71#_M1025_g N_VGND_c_2485_n 0.00497279f $X=10.14 $Y=0.695 $X2=0
+ $Y2=0
cc_1191 N_A_2013_71#_M1025_g N_VGND_c_2496_n 0.00509887f $X=10.14 $Y=0.695 $X2=0
+ $Y2=0
cc_1192 N_A_2013_71#_c_1558_n N_VGND_c_2496_n 0.0038545f $X=12.01 $Y=1.11 $X2=0
+ $Y2=0
cc_1193 N_A_1784_97#_M1032_g N_VPWR_c_2029_n 0.0042229f $X=10.7 $Y=2.41 $X2=0
+ $Y2=0
cc_1194 N_A_1784_97#_c_1673_n N_VPWR_c_2029_n 0.00626404f $X=9.42 $Y=2.755 $X2=0
+ $Y2=0
cc_1195 N_A_1784_97#_M1032_g N_VPWR_c_2030_n 0.0059693f $X=10.7 $Y=2.41 $X2=0
+ $Y2=0
cc_1196 N_A_1784_97#_M1032_g N_VPWR_c_2038_n 0.00585197f $X=10.7 $Y=2.41 $X2=0
+ $Y2=0
cc_1197 N_A_1784_97#_c_1673_n N_VPWR_c_2044_n 0.0154692f $X=9.42 $Y=2.755 $X2=0
+ $Y2=0
cc_1198 N_A_1784_97#_M1032_g N_VPWR_c_2023_n 0.00606454f $X=10.7 $Y=2.41 $X2=0
+ $Y2=0
cc_1199 N_A_1784_97#_c_1673_n N_VPWR_c_2023_n 0.0127033f $X=9.42 $Y=2.755 $X2=0
+ $Y2=0
cc_1200 N_A_1784_97#_c_1674_n N_A_691_113#_c_2239_n 0.0089467f $X=9.405 $Y=2.53
+ $X2=0 $Y2=0
cc_1201 N_A_1784_97#_c_1673_n N_A_691_113#_c_2240_n 0.0133064f $X=9.42 $Y=2.755
+ $X2=0 $Y2=0
cc_1202 N_A_1784_97#_M1018_g N_VGND_c_2466_n 0.00193352f $X=10.9 $Y=0.69 $X2=0
+ $Y2=0
cc_1203 N_A_1784_97#_M1018_g N_VGND_c_2486_n 0.00278237f $X=10.9 $Y=0.69 $X2=0
+ $Y2=0
cc_1204 N_A_1784_97#_M1018_g N_VGND_c_2496_n 0.00363424f $X=10.9 $Y=0.69 $X2=0
+ $Y2=0
cc_1205 N_A_2489_74#_M1044_g N_VPWR_c_2031_n 0.00649758f $X=14.415 $Y=2.4 $X2=0
+ $Y2=0
cc_1206 N_A_2489_74#_c_1776_n N_VPWR_c_2031_n 0.0121551f $X=13.24 $Y=2.75 $X2=0
+ $Y2=0
cc_1207 N_A_2489_74#_M1044_g N_VPWR_c_2032_n 0.00333672f $X=14.415 $Y=2.4 $X2=0
+ $Y2=0
cc_1208 N_A_2489_74#_M1036_g N_VPWR_c_2032_n 0.0118211f $X=15.425 $Y=2.4 $X2=0
+ $Y2=0
cc_1209 N_A_2489_74#_M1039_g N_VPWR_c_2032_n 0.00125818f $X=15.875 $Y=2.4 $X2=0
+ $Y2=0
cc_1210 N_A_2489_74#_M1036_g N_VPWR_c_2033_n 0.00125818f $X=15.425 $Y=2.4 $X2=0
+ $Y2=0
cc_1211 N_A_2489_74#_M1039_g N_VPWR_c_2033_n 0.0106899f $X=15.875 $Y=2.4 $X2=0
+ $Y2=0
cc_1212 N_A_2489_74#_c_1776_n N_VPWR_c_2045_n 0.018423f $X=13.24 $Y=2.75 $X2=0
+ $Y2=0
cc_1213 N_A_2489_74#_M1044_g N_VPWR_c_2046_n 0.005209f $X=14.415 $Y=2.4 $X2=0
+ $Y2=0
cc_1214 N_A_2489_74#_M1036_g N_VPWR_c_2047_n 0.00460063f $X=15.425 $Y=2.4 $X2=0
+ $Y2=0
cc_1215 N_A_2489_74#_M1039_g N_VPWR_c_2047_n 0.00460063f $X=15.875 $Y=2.4 $X2=0
+ $Y2=0
cc_1216 N_A_2489_74#_M1044_g N_VPWR_c_2023_n 0.00988813f $X=14.415 $Y=2.4 $X2=0
+ $Y2=0
cc_1217 N_A_2489_74#_M1036_g N_VPWR_c_2023_n 0.0046086f $X=15.425 $Y=2.4 $X2=0
+ $Y2=0
cc_1218 N_A_2489_74#_M1039_g N_VPWR_c_2023_n 0.0046086f $X=15.875 $Y=2.4 $X2=0
+ $Y2=0
cc_1219 N_A_2489_74#_c_1776_n N_VPWR_c_2023_n 0.0152212f $X=13.24 $Y=2.75 $X2=0
+ $Y2=0
cc_1220 N_A_2489_74#_M1036_g Q 0.00988085f $X=15.425 $Y=2.4 $X2=0 $Y2=0
cc_1221 N_A_2489_74#_M1026_g Q 0.016221f $X=15.445 $Y=0.74 $X2=0 $Y2=0
cc_1222 N_A_2489_74#_M1039_g Q 0.00910089f $X=15.875 $Y=2.4 $X2=0 $Y2=0
cc_1223 N_A_2489_74#_M1047_g Q 0.0145925f $X=15.875 $Y=0.74 $X2=0 $Y2=0
cc_1224 N_A_2489_74#_c_1762_n Q 0.0264058f $X=15.875 $Y=1.465 $X2=0 $Y2=0
cc_1225 N_A_2489_74#_c_1764_n N_VGND_M1022_d 0.00511003f $X=13.695 $Y=0.855
+ $X2=0 $Y2=0
cc_1226 N_A_2489_74#_c_1763_n N_VGND_c_2467_n 0.010811f $X=12.585 $Y=0.515 $X2=0
+ $Y2=0
cc_1227 N_A_2489_74#_c_1764_n N_VGND_c_2468_n 0.0147778f $X=13.695 $Y=0.855
+ $X2=0 $Y2=0
cc_1228 N_A_2489_74#_c_1763_n N_VGND_c_2469_n 0.00419512f $X=12.585 $Y=0.515
+ $X2=0 $Y2=0
cc_1229 N_A_2489_74#_c_1764_n N_VGND_c_2469_n 0.024775f $X=13.695 $Y=0.855 $X2=0
+ $Y2=0
cc_1230 N_A_2489_74#_M1012_g N_VGND_c_2470_n 0.00106276f $X=14.455 $Y=0.74 $X2=0
+ $Y2=0
cc_1231 N_A_2489_74#_c_1764_n N_VGND_c_2470_n 0.0125741f $X=13.695 $Y=0.855
+ $X2=0 $Y2=0
cc_1232 N_A_2489_74#_c_1765_n N_VGND_c_2470_n 0.011522f $X=13.78 $Y=1.3 $X2=0
+ $Y2=0
cc_1233 N_A_2489_74#_c_1767_n N_VGND_c_2470_n 0.0210027f $X=14.33 $Y=1.465 $X2=0
+ $Y2=0
cc_1234 N_A_2489_74#_c_1768_n N_VGND_c_2470_n 0.00395268f $X=14.33 $Y=1.465
+ $X2=0 $Y2=0
cc_1235 N_A_2489_74#_M1012_g N_VGND_c_2471_n 0.00434272f $X=14.455 $Y=0.74 $X2=0
+ $Y2=0
cc_1236 N_A_2489_74#_M1012_g N_VGND_c_2472_n 0.00413259f $X=14.455 $Y=0.74 $X2=0
+ $Y2=0
cc_1237 N_A_2489_74#_c_1757_n N_VGND_c_2472_n 0.006711f $X=15.335 $Y=1.465 $X2=0
+ $Y2=0
cc_1238 N_A_2489_74#_M1026_g N_VGND_c_2472_n 0.00646793f $X=15.445 $Y=0.74 $X2=0
+ $Y2=0
cc_1239 N_A_2489_74#_M1026_g N_VGND_c_2473_n 0.00422942f $X=15.445 $Y=0.74 $X2=0
+ $Y2=0
cc_1240 N_A_2489_74#_M1047_g N_VGND_c_2473_n 0.00434272f $X=15.875 $Y=0.74 $X2=0
+ $Y2=0
cc_1241 N_A_2489_74#_M1047_g N_VGND_c_2474_n 0.00313962f $X=15.875 $Y=0.74 $X2=0
+ $Y2=0
cc_1242 N_A_2489_74#_c_1763_n N_VGND_c_2481_n 0.014415f $X=12.585 $Y=0.515 $X2=0
+ $Y2=0
cc_1243 N_A_2489_74#_M1012_g N_VGND_c_2493_n 0.005596f $X=14.455 $Y=0.74 $X2=0
+ $Y2=0
cc_1244 N_A_2489_74#_M1012_g N_VGND_c_2496_n 0.00830035f $X=14.455 $Y=0.74 $X2=0
+ $Y2=0
cc_1245 N_A_2489_74#_M1026_g N_VGND_c_2496_n 0.00788596f $X=15.445 $Y=0.74 $X2=0
+ $Y2=0
cc_1246 N_A_2489_74#_M1047_g N_VGND_c_2496_n 0.00820382f $X=15.875 $Y=0.74 $X2=0
+ $Y2=0
cc_1247 N_A_2489_74#_c_1763_n N_VGND_c_2496_n 0.0119404f $X=12.585 $Y=0.515
+ $X2=0 $Y2=0
cc_1248 N_A_2489_74#_c_1764_n N_VGND_c_2496_n 0.0209551f $X=13.695 $Y=0.855
+ $X2=0 $Y2=0
cc_1249 N_A_2489_74#_c_1764_n A_2591_74# 0.0023798f $X=13.695 $Y=0.855 $X2=-0.19
+ $Y2=-0.245
cc_1250 N_A_32_74#_c_1914_n A_135_464# 0.0048076f $X=1.485 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_1251 N_A_32_74#_c_1914_n N_VPWR_M1003_d 0.00481895f $X=1.485 $Y=2.375
+ $X2=-0.19 $Y2=-0.245
cc_1252 N_A_32_74#_c_1916_n N_VPWR_M1013_d 4.26874e-19 $X=2.165 $Y=2.99 $X2=0
+ $Y2=0
cc_1253 N_A_32_74#_c_1956_n N_VPWR_M1013_d 0.00485499f $X=2.25 $Y=2.905 $X2=0
+ $Y2=0
cc_1254 N_A_32_74#_c_1918_n N_VPWR_M1013_d 0.00936314f $X=3.265 $Y=2.375 $X2=0
+ $Y2=0
cc_1255 N_A_32_74#_c_1913_n N_VPWR_c_2024_n 0.0101945f $X=0.36 $Y=2.465 $X2=0
+ $Y2=0
cc_1256 N_A_32_74#_c_1914_n N_VPWR_c_2024_n 0.015347f $X=1.485 $Y=2.375 $X2=0
+ $Y2=0
cc_1257 N_A_32_74#_c_1915_n N_VPWR_c_2024_n 0.0208966f $X=1.57 $Y=2.905 $X2=0
+ $Y2=0
cc_1258 N_A_32_74#_c_1917_n N_VPWR_c_2024_n 0.0146661f $X=1.655 $Y=2.99 $X2=0
+ $Y2=0
cc_1259 N_A_32_74#_c_1916_n N_VPWR_c_2025_n 0.0146f $X=2.165 $Y=2.99 $X2=0 $Y2=0
cc_1260 N_A_32_74#_c_1956_n N_VPWR_c_2025_n 0.0205315f $X=2.25 $Y=2.905 $X2=0
+ $Y2=0
cc_1261 N_A_32_74#_c_1918_n N_VPWR_c_2025_n 0.015347f $X=3.265 $Y=2.375 $X2=0
+ $Y2=0
cc_1262 N_A_32_74#_c_1922_n N_VPWR_c_2025_n 0.0100543f $X=3.43 $Y=2.455 $X2=0
+ $Y2=0
cc_1263 N_A_32_74#_c_1913_n N_VPWR_c_2040_n 0.0194699f $X=0.36 $Y=2.465 $X2=0
+ $Y2=0
cc_1264 N_A_32_74#_c_1916_n N_VPWR_c_2041_n 0.0444245f $X=2.165 $Y=2.99 $X2=0
+ $Y2=0
cc_1265 N_A_32_74#_c_1917_n N_VPWR_c_2041_n 0.0121867f $X=1.655 $Y=2.99 $X2=0
+ $Y2=0
cc_1266 N_A_32_74#_c_1922_n N_VPWR_c_2042_n 0.0118405f $X=3.43 $Y=2.455 $X2=0
+ $Y2=0
cc_1267 N_A_32_74#_c_1913_n N_VPWR_c_2023_n 0.0160419f $X=0.36 $Y=2.465 $X2=0
+ $Y2=0
cc_1268 N_A_32_74#_c_1916_n N_VPWR_c_2023_n 0.0256732f $X=2.165 $Y=2.99 $X2=0
+ $Y2=0
cc_1269 N_A_32_74#_c_1917_n N_VPWR_c_2023_n 0.00660921f $X=1.655 $Y=2.99 $X2=0
+ $Y2=0
cc_1270 N_A_32_74#_c_1922_n N_VPWR_c_2023_n 0.0101813f $X=3.43 $Y=2.455 $X2=0
+ $Y2=0
cc_1271 N_A_32_74#_c_1918_n A_581_462# 0.00366293f $X=3.265 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_1272 N_A_32_74#_c_1922_n N_A_691_113#_c_2231_n 0.00699176f $X=3.43 $Y=2.455
+ $X2=0 $Y2=0
cc_1273 N_A_32_74#_c_1922_n N_A_691_113#_c_2243_n 0.00351236f $X=3.43 $Y=2.455
+ $X2=0 $Y2=0
cc_1274 N_A_32_74#_c_1908_n N_A_691_113#_c_2228_n 0.0188786f $X=3.165 $Y=0.775
+ $X2=0 $Y2=0
cc_1275 N_A_32_74#_c_1911_n N_A_691_113#_c_2228_n 0.00333703f $X=3.46 $Y=1.26
+ $X2=0 $Y2=0
cc_1276 N_A_32_74#_c_1908_n N_A_691_113#_c_2229_n 0.00645754f $X=3.165 $Y=0.775
+ $X2=0 $Y2=0
cc_1277 N_A_32_74#_c_1909_n N_A_691_113#_c_2229_n 0.0697173f $X=3.46 $Y=2.29
+ $X2=0 $Y2=0
cc_1278 N_A_32_74#_c_1911_n N_A_691_113#_c_2229_n 0.0136555f $X=3.46 $Y=1.26
+ $X2=0 $Y2=0
cc_1279 N_A_32_74#_c_1910_n N_VGND_c_2461_n 0.0100909f $X=0.415 $Y=0.585 $X2=0
+ $Y2=0
cc_1280 N_A_32_74#_c_1908_n N_VGND_c_2462_n 0.0145731f $X=3.165 $Y=0.775 $X2=0
+ $Y2=0
cc_1281 N_A_32_74#_c_1910_n N_VGND_c_2482_n 0.0149954f $X=0.415 $Y=0.585 $X2=0
+ $Y2=0
cc_1282 N_A_32_74#_c_1908_n N_VGND_c_2483_n 0.00794834f $X=3.165 $Y=0.775 $X2=0
+ $Y2=0
cc_1283 N_A_32_74#_c_1908_n N_VGND_c_2496_n 0.0105391f $X=3.165 $Y=0.775 $X2=0
+ $Y2=0
cc_1284 N_A_32_74#_c_1910_n N_VGND_c_2496_n 0.0168506f $X=0.415 $Y=0.585 $X2=0
+ $Y2=0
cc_1285 N_VPWR_c_2026_n N_A_691_113#_c_2232_n 0.0148242f $X=5.13 $Y=2.76 $X2=0
+ $Y2=0
cc_1286 N_VPWR_c_2042_n N_A_691_113#_c_2232_n 0.0567624f $X=5.035 $Y=3.33 $X2=0
+ $Y2=0
cc_1287 N_VPWR_c_2023_n N_A_691_113#_c_2232_n 0.0303734f $X=17.04 $Y=3.33 $X2=0
+ $Y2=0
cc_1288 N_VPWR_c_2042_n N_A_691_113#_c_2243_n 0.0170104f $X=5.035 $Y=3.33 $X2=0
+ $Y2=0
cc_1289 N_VPWR_c_2023_n N_A_691_113#_c_2243_n 0.00854122f $X=17.04 $Y=3.33 $X2=0
+ $Y2=0
cc_1290 N_VPWR_M1014_d N_A_691_113#_c_2259_n 0.00523858f $X=4.765 $Y=2.265 $X2=0
+ $Y2=0
cc_1291 N_VPWR_c_2026_n N_A_691_113#_c_2259_n 0.0232873f $X=5.13 $Y=2.76 $X2=0
+ $Y2=0
cc_1292 N_VPWR_M1014_d N_A_691_113#_c_2233_n 0.00974124f $X=4.765 $Y=2.265 $X2=0
+ $Y2=0
cc_1293 N_VPWR_c_2026_n N_A_691_113#_c_2233_n 0.0169742f $X=5.13 $Y=2.76 $X2=0
+ $Y2=0
cc_1294 N_VPWR_M1000_s N_A_691_113#_c_2224_n 0.00609051f $X=6.425 $Y=1.84 $X2=0
+ $Y2=0
cc_1295 N_VPWR_M1000_s N_A_691_113#_c_2236_n 0.00575729f $X=6.425 $Y=1.84 $X2=0
+ $Y2=0
cc_1296 N_VPWR_M1008_s N_A_691_113#_c_2236_n 0.00250916f $X=7.815 $Y=1.84 $X2=0
+ $Y2=0
cc_1297 N_VPWR_c_2027_n N_A_691_113#_c_2236_n 0.0150227f $X=6.57 $Y=2.815 $X2=0
+ $Y2=0
cc_1298 N_VPWR_c_2028_n N_A_691_113#_c_2236_n 0.00870407f $X=7.96 $Y=2.815 $X2=0
+ $Y2=0
cc_1299 N_VPWR_c_2023_n N_A_691_113#_c_2236_n 0.0367797f $X=17.04 $Y=3.33 $X2=0
+ $Y2=0
cc_1300 N_VPWR_M1000_s N_A_691_113#_c_2237_n 0.00258383f $X=6.425 $Y=1.84 $X2=0
+ $Y2=0
cc_1301 N_VPWR_c_2026_n N_A_691_113#_c_2237_n 0.00972016f $X=5.13 $Y=2.76 $X2=0
+ $Y2=0
cc_1302 N_VPWR_c_2027_n N_A_691_113#_c_2237_n 0.0217987f $X=6.57 $Y=2.815 $X2=0
+ $Y2=0
cc_1303 N_VPWR_c_2036_n N_A_691_113#_c_2237_n 0.0166983f $X=6.485 $Y=3.33 $X2=0
+ $Y2=0
cc_1304 N_VPWR_c_2023_n N_A_691_113#_c_2237_n 0.022982f $X=17.04 $Y=3.33 $X2=0
+ $Y2=0
cc_1305 N_VPWR_M1008_s N_A_691_113#_c_2238_n 0.011134f $X=7.815 $Y=1.84 $X2=0
+ $Y2=0
cc_1306 N_VPWR_c_2028_n N_A_691_113#_c_2252_n 0.00212051f $X=7.96 $Y=2.815 $X2=0
+ $Y2=0
cc_1307 N_VPWR_c_2023_n N_A_691_113#_c_2252_n 0.00492308f $X=17.04 $Y=3.33 $X2=0
+ $Y2=0
cc_1308 N_VPWR_c_2044_n N_A_691_113#_c_2239_n 0.00557176f $X=10.225 $Y=3.33
+ $X2=0 $Y2=0
cc_1309 N_VPWR_c_2023_n N_A_691_113#_c_2239_n 0.00937585f $X=17.04 $Y=3.33 $X2=0
+ $Y2=0
cc_1310 N_VPWR_c_2044_n N_A_691_113#_c_2240_n 0.0108228f $X=10.225 $Y=3.33 $X2=0
+ $Y2=0
cc_1311 N_VPWR_c_2023_n N_A_691_113#_c_2240_n 0.00906589f $X=17.04 $Y=3.33 $X2=0
+ $Y2=0
cc_1312 N_VPWR_M1008_s N_A_691_113#_c_2390_n 0.00153606f $X=7.815 $Y=1.84 $X2=0
+ $Y2=0
cc_1313 N_VPWR_c_2028_n N_A_691_113#_c_2390_n 0.0116705f $X=7.96 $Y=2.815 $X2=0
+ $Y2=0
cc_1314 N_VPWR_c_2023_n N_A_691_113#_c_2390_n 6.0606e-19 $X=17.04 $Y=3.33 $X2=0
+ $Y2=0
cc_1315 N_VPWR_c_2044_n N_A_691_113#_c_2329_n 0.00251491f $X=10.225 $Y=3.33
+ $X2=0 $Y2=0
cc_1316 N_VPWR_c_2023_n N_A_691_113#_c_2329_n 0.00477661f $X=17.04 $Y=3.33 $X2=0
+ $Y2=0
cc_1317 N_VPWR_M1046_d N_Q_N_c_2429_n 0.00311223f $X=16.865 $Y=1.84 $X2=0 $Y2=0
cc_1318 N_VPWR_c_2035_n N_Q_N_c_2429_n 0.0219147f $X=17 $Y=2.25 $X2=0 $Y2=0
cc_1319 N_VPWR_c_2033_n Q_N 0.015063f $X=16.1 $Y=2.78 $X2=0 $Y2=0
cc_1320 N_VPWR_c_2035_n Q_N 0.034387f $X=17 $Y=2.25 $X2=0 $Y2=0
cc_1321 N_VPWR_c_2048_n Q_N 0.0115612f $X=16.835 $Y=3.33 $X2=0 $Y2=0
cc_1322 N_VPWR_c_2023_n Q_N 0.00856962f $X=17.04 $Y=3.33 $X2=0 $Y2=0
cc_1323 N_A_691_113#_c_2233_n A_1091_453# 0.0048076f $X=5.845 $Y=2.34 $X2=-0.19
+ $Y2=-0.245
cc_1324 N_A_691_113#_c_2230_n N_VGND_M1029_s 7.58458e-19 $X=6.39 $Y=1.175 $X2=0
+ $Y2=0
cc_1325 N_A_691_113#_c_2223_n N_VGND_c_2463_n 0.00634222f $X=5.985 $Y=0.835
+ $X2=0 $Y2=0
cc_1326 N_A_691_113#_c_2223_n N_VGND_c_2464_n 0.0192622f $X=5.985 $Y=0.835 $X2=0
+ $Y2=0
cc_1327 N_A_691_113#_c_2230_n N_VGND_c_2464_n 0.00485909f $X=6.39 $Y=1.175 $X2=0
+ $Y2=0
cc_1328 N_A_691_113#_c_2228_n N_VGND_c_2483_n 0.00932016f $X=3.665 $Y=0.775
+ $X2=0 $Y2=0
cc_1329 N_A_691_113#_c_2223_n N_VGND_c_2484_n 0.00684598f $X=5.985 $Y=0.835
+ $X2=0 $Y2=0
cc_1330 N_A_691_113#_c_2223_n N_VGND_c_2496_n 0.00989908f $X=5.985 $Y=0.835
+ $X2=0 $Y2=0
cc_1331 N_A_691_113#_c_2228_n N_VGND_c_2496_n 0.0122951f $X=3.665 $Y=0.775 $X2=0
+ $Y2=0
cc_1332 Q N_VGND_c_2472_n 0.0309174f $X=15.515 $Y=0.47 $X2=0 $Y2=0
cc_1333 Q N_VGND_c_2473_n 0.0149085f $X=15.515 $Y=0.47 $X2=0 $Y2=0
cc_1334 Q N_VGND_c_2474_n 0.0294574f $X=15.515 $Y=0.47 $X2=0 $Y2=0
cc_1335 Q N_VGND_c_2496_n 0.0122037f $X=15.515 $Y=0.47 $X2=0 $Y2=0
cc_1336 N_Q_N_c_2428_n N_VGND_M1041_s 0.00328964f $X=16.932 $Y=1.13 $X2=0 $Y2=0
cc_1337 N_Q_N_c_2428_n N_VGND_c_2474_n 0.00741094f $X=16.932 $Y=1.13 $X2=0 $Y2=0
cc_1338 Q_N N_VGND_c_2474_n 0.0225498f $X=16.475 $Y=0.47 $X2=0 $Y2=0
cc_1339 N_Q_N_c_2428_n N_VGND_c_2476_n 0.0201545f $X=16.932 $Y=1.13 $X2=0 $Y2=0
cc_1340 Q_N N_VGND_c_2476_n 0.0172723f $X=16.475 $Y=0.47 $X2=0 $Y2=0
cc_1341 Q_N N_VGND_c_2487_n 0.014379f $X=16.475 $Y=0.47 $X2=0 $Y2=0
cc_1342 Q_N N_VGND_c_2496_n 0.0118382f $X=16.475 $Y=0.47 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__clkinv_4.pex.spice
* Created: Fri Aug 28 17:20:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__CLKINV_4%A 3 6 9 13 17 21 25 29 33 37 41 43 44 45 46
+ 47 54 68
r107 67 68 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.805 $Y=1.515
+ $X2=2.82 $Y2=1.515
r108 65 67 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=2.39 $Y=1.515
+ $X2=2.805 $Y2=1.515
r109 65 66 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.39
+ $Y=1.515 $X2=2.39 $Y2=1.515
r110 63 65 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.365 $Y=1.515
+ $X2=2.39 $Y2=1.515
r111 62 63 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=2.355 $Y=1.515
+ $X2=2.365 $Y2=1.515
r112 61 62 87.4306 $w=3.3e-07 $l=5e-07 $layer=POLY_cond $X=1.855 $Y=1.515
+ $X2=2.355 $Y2=1.515
r113 60 61 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=1.795 $Y=1.515
+ $X2=1.855 $Y2=1.515
r114 59 60 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=1.405 $Y=1.515
+ $X2=1.795 $Y2=1.515
r115 57 59 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=1.03 $Y=1.515
+ $X2=1.405 $Y2=1.515
r116 57 58 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=1.03
+ $Y=1.515 $X2=1.03 $Y2=1.515
r117 55 57 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.955 $Y=1.515
+ $X2=1.03 $Y2=1.515
r118 53 55 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.94 $Y=1.515
+ $X2=0.955 $Y2=1.515
r119 53 54 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.94 $Y=1.515
+ $X2=0.865 $Y2=1.515
r120 47 66 6.70025 $w=4.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.39 $Y2=1.565
r121 46 66 6.16423 $w=4.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.39 $Y2=1.565
r122 45 46 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=2.16 $Y2=1.565
r123 44 45 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.68 $Y2=1.565
r124 44 58 4.55617 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.03 $Y2=1.565
r125 43 58 8.30831 $w=4.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.03 $Y2=1.565
r126 39 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.82 $Y=1.35
+ $X2=2.82 $Y2=1.515
r127 39 41 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.82 $Y=1.35
+ $X2=2.82 $Y2=0.61
r128 35 67 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.805 $Y=1.68
+ $X2=2.805 $Y2=1.515
r129 35 37 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.805 $Y=1.68
+ $X2=2.805 $Y2=2.4
r130 31 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.365 $Y=1.35
+ $X2=2.365 $Y2=1.515
r131 31 33 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.365 $Y=1.35
+ $X2=2.365 $Y2=0.61
r132 27 62 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.355 $Y=1.68
+ $X2=2.355 $Y2=1.515
r133 27 29 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.355 $Y=1.68
+ $X2=2.355 $Y2=2.4
r134 23 61 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.68
+ $X2=1.855 $Y2=1.515
r135 23 25 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.855 $Y=1.68
+ $X2=1.855 $Y2=2.4
r136 19 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.795 $Y=1.35
+ $X2=1.795 $Y2=1.515
r137 19 21 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.795 $Y=1.35
+ $X2=1.795 $Y2=0.61
r138 15 59 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.68
+ $X2=1.405 $Y2=1.515
r139 15 17 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.405 $Y=1.68
+ $X2=1.405 $Y2=2.4
r140 11 55 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.68
+ $X2=0.955 $Y2=1.515
r141 11 13 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.955 $Y=1.68
+ $X2=0.955 $Y2=2.4
r142 7 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.94 $Y=1.35
+ $X2=0.94 $Y2=1.515
r143 7 9 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.94 $Y=1.35 $X2=0.94
+ $Y2=0.61
r144 6 54 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.595 $Y=1.605
+ $X2=0.865 $Y2=1.605
r145 1 6 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=0.505 $Y=1.68
+ $X2=0.595 $Y2=1.605
r146 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.505 $Y=1.68
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__CLKINV_4%VPWR 1 2 3 4 13 15 19 23 25 27 30 31 32 38
+ 42 51 55
r53 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 46 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 46 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r58 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 43 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.12 $Y2=3.33
r60 43 45 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 42 54 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=3.137 $Y2=3.33
r62 42 45 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 38 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=2.12 $Y2=3.33
r64 38 40 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 37 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r66 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r67 34 48 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r68 34 36 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r69 32 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r70 32 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r71 32 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r72 30 36 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.72 $Y2=3.33
r73 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.18 $Y2=3.33
r74 29 40 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.68 $Y2=3.33
r75 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.18 $Y2=3.33
r76 25 54 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.137 $Y2=3.33
r77 25 27 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.08 $Y2=2.455
r78 21 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=3.245
+ $X2=2.12 $Y2=3.33
r79 21 23 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=2.12 $Y=3.245
+ $X2=2.12 $Y2=2.455
r80 17 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r81 17 19 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.455
r82 13 48 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r83 13 15 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.455
r84 4 27 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=2.895
+ $Y=1.84 $X2=3.08 $Y2=2.455
r85 3 23 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.945
+ $Y=1.84 $X2=2.08 $Y2=2.455
r86 2 19 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.045
+ $Y=1.84 $X2=1.18 $Y2=2.455
r87 1 15 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__CLKINV_4%Y 1 2 3 4 5 17 19 22 24 25 28 30 32 36 40
+ 42 44 52 53 55 56 58 61
r107 60 61 32.8196 $w=2.28e-07 $l=6.55e-07 $layer=LI1_cond $X=3.12 $Y=1.95
+ $X2=3.12 $Y2=1.295
r108 59 61 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=1.18
+ $X2=3.12 $Y2=1.295
r109 51 53 10.9648 $w=7.23e-07 $l=1.65e-07 $layer=LI1_cond $X=1.58 $Y=0.817
+ $X2=1.745 $Y2=0.817
r110 51 52 17.9763 $w=7.23e-07 $l=5.9e-07 $layer=LI1_cond $X=1.58 $Y=0.817
+ $X2=0.99 $Y2=0.817
r111 46 49 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.35 $Y=2.035
+ $X2=0.73 $Y2=2.035
r112 45 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=2.035
+ $X2=2.58 $Y2=2.035
r113 44 60 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.005 $Y=2.035
+ $X2=3.12 $Y2=1.95
r114 44 45 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.005 $Y=2.035
+ $X2=2.745 $Y2=2.035
r115 43 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=1.095
+ $X2=2.58 $Y2=1.095
r116 42 59 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.005 $Y=1.095
+ $X2=3.12 $Y2=1.18
r117 42 43 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.005 $Y=1.095
+ $X2=2.745 $Y2=1.095
r118 38 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=2.12
+ $X2=2.58 $Y2=2.035
r119 38 40 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.58 $Y=2.12
+ $X2=2.58 $Y2=2.815
r120 34 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=1.01
+ $X2=2.58 $Y2=1.095
r121 34 36 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=2.58 $Y=1.01 $X2=2.58
+ $Y2=0.61
r122 33 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=2.035
+ $X2=1.63 $Y2=2.035
r123 32 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=2.035
+ $X2=2.58 $Y2=2.035
r124 32 33 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.415 $Y=2.035
+ $X2=1.795 $Y2=2.035
r125 30 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=1.095
+ $X2=2.58 $Y2=1.095
r126 30 53 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.415 $Y=1.095
+ $X2=1.745 $Y2=1.095
r127 26 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=2.12
+ $X2=1.63 $Y2=2.035
r128 26 28 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.63 $Y=2.12
+ $X2=1.63 $Y2=2.815
r129 25 49 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=2.035
+ $X2=0.73 $Y2=2.035
r130 24 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=2.035
+ $X2=1.63 $Y2=2.035
r131 24 25 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.465 $Y=2.035
+ $X2=0.895 $Y2=2.035
r132 22 49 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.73 $Y=2.815
+ $X2=0.73 $Y2=2.12
r133 19 52 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=0.435 $Y=1.095
+ $X2=0.99 $Y2=1.095
r134 17 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.35 $Y=1.95
+ $X2=0.35 $Y2=2.035
r135 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.35 $Y=1.18
+ $X2=0.435 $Y2=1.095
r136 16 17 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.35 $Y=1.18
+ $X2=0.35 $Y2=1.95
r137 5 58 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=2.445
+ $Y=1.84 $X2=2.58 $Y2=2.035
r138 5 40 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.445
+ $Y=1.84 $X2=2.58 $Y2=2.815
r139 4 55 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.84 $X2=1.63 $Y2=2.035
r140 4 28 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=1.84 $X2=1.63 $Y2=2.815
r141 3 49 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.035
r142 3 22 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.815
r143 2 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.44
+ $Y=0.4 $X2=2.58 $Y2=0.61
r144 1 51 91 $w=1.7e-07 $l=6.65977e-07 $layer=licon1_NDIFF $count=2 $X=1.015
+ $Y=0.4 $X2=1.58 $Y2=0.62
.ends

.subckt PM_SKY130_FD_SC_MS__CLKINV_4%VGND 1 2 3 12 14 16 18 20 25 31 38 42
r31 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r32 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r33 32 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r34 31 36 9.12071 $w=7.29e-07 $l=5.45e-07 $layer=LI1_cond $X=0.41 $Y=0 $X2=0.41
+ $Y2=0.545
r35 31 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r36 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r37 29 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r38 29 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r39 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r40 26 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.08
+ $Y2=0
r41 26 28 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.64
+ $Y2=0
r42 25 41 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=3.137
+ $Y2=0
r43 25 28 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=2.64
+ $Y2=0
r44 21 31 9.58964 $w=1.7e-07 $l=4.1e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=0.41
+ $Y2=0
r45 21 23 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=1.68
+ $Y2=0
r46 20 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.915 $Y=0 $X2=2.08
+ $Y2=0
r47 20 23 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.915 $Y=0 $X2=1.68
+ $Y2=0
r48 18 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r49 18 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r50 18 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r51 14 41 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.137 $Y2=0
r52 14 16 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0.61
r53 10 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=0.085
+ $X2=2.08 $Y2=0
r54 10 12 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=2.08 $Y=0.085
+ $X2=2.08 $Y2=0.61
r55 3 16 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.4 $X2=3.08 $Y2=0.61
r56 2 12 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=1.87
+ $Y=0.4 $X2=2.08 $Y2=0.61
r57 1 36 91 $w=1.7e-07 $l=5.88048e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.4 $X2=0.655 $Y2=0.545
.ends


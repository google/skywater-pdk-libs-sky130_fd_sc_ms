* File: sky130_fd_sc_ms__clkbuf_2.pex.spice
* Created: Fri Aug 28 17:17:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__CLKBUF_2%A_43_192# 1 2 9 13 17 21 25 29 30 31 34 37
+ 38 40 44 49
c79 30 0 1.09492e-19 $X=1.535 $Y=2.405
r80 48 49 1.5971 $w=6.7e-07 $l=2e-08 $layer=POLY_cond $X=0.925 $Y=1.295
+ $X2=0.945 $Y2=1.295
r81 47 48 34.3377 $w=6.7e-07 $l=4.3e-07 $layer=POLY_cond $X=0.495 $Y=1.295
+ $X2=0.925 $Y2=1.295
r82 40 42 10.5918 $w=3.58e-07 $l=2.3e-07 $layer=LI1_cond $X=1.655 $Y=0.58
+ $X2=1.655 $Y2=0.81
r83 37 44 3.91525 $w=2.35e-07 $l=1.12916e-07 $layer=LI1_cond $X=1.75 $Y=2.32
+ $X2=1.685 $Y2=2.405
r84 37 42 98.5134 $w=1.68e-07 $l=1.51e-06 $layer=LI1_cond $X=1.75 $Y=2.32
+ $X2=1.75 $Y2=0.81
r85 32 44 3.91525 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.685 $Y=2.49
+ $X2=1.685 $Y2=2.405
r86 32 34 12.4848 $w=2.98e-07 $l=3.25e-07 $layer=LI1_cond $X=1.685 $Y=2.49
+ $X2=1.685 $Y2=2.815
r87 30 44 2.53056 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.535 $Y=2.405
+ $X2=1.685 $Y2=2.405
r88 30 31 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=1.535 $Y=2.405
+ $X2=0.385 $Y2=2.405
r89 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.3 $Y=2.32
+ $X2=0.385 $Y2=2.405
r90 29 38 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.3 $Y=2.32 $X2=0.3
+ $Y2=1.63
r91 26 47 9.18334 $w=6.7e-07 $l=1.15e-07 $layer=POLY_cond $X=0.38 $Y=1.295
+ $X2=0.495 $Y2=1.295
r92 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.38
+ $Y=1.125 $X2=0.38 $Y2=1.125
r93 23 38 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.38 $Y=1.465
+ $X2=0.38 $Y2=1.63
r94 23 25 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.38 $Y=1.465
+ $X2=0.38 $Y2=1.125
r95 19 49 34.2182 $w=1.8e-07 $l=3.35e-07 $layer=POLY_cond $X=0.945 $Y=1.63
+ $X2=0.945 $Y2=1.295
r96 19 21 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.945 $Y=1.63
+ $X2=0.945 $Y2=2.4
r97 15 48 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.925 $Y=0.96
+ $X2=0.925 $Y2=1.295
r98 15 17 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=0.925 $Y=0.96
+ $X2=0.925 $Y2=0.58
r99 11 47 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.495 $Y=0.96
+ $X2=0.495 $Y2=1.295
r100 11 13 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=0.495 $Y=0.96
+ $X2=0.495 $Y2=0.58
r101 7 47 34.2182 $w=1.8e-07 $l=3.35e-07 $layer=POLY_cond $X=0.495 $Y=1.63
+ $X2=0.495 $Y2=1.295
r102 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.495 $Y=1.63
+ $X2=0.495 $Y2=2.4
r103 2 44 600 $w=1.7e-07 $l=6.33364e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.84 $X2=1.63 $Y2=2.405
r104 2 34 600 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=1.84 $X2=1.63 $Y2=2.815
r105 1 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.37 $X2=1.64 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__CLKBUF_2%A 3 7 11 12 13 14 15 20 21
c38 12 0 1.09492e-19 $X=1.41 $Y=1.68
r39 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.41
+ $Y=1.175 $X2=1.41 $Y2=1.175
r40 14 15 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.29 $Y=1.665
+ $X2=1.29 $Y2=2.035
r41 13 14 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.29 $Y=1.295
+ $X2=1.29 $Y2=1.665
r42 13 21 3.373 $w=4.08e-07 $l=1.2e-07 $layer=LI1_cond $X=1.29 $Y=1.295 $X2=1.29
+ $Y2=1.175
r43 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.41 $Y=1.515
+ $X2=1.41 $Y2=1.175
r44 11 12 35.4289 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.515
+ $X2=1.41 $Y2=1.68
r45 10 20 38.3209 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.01
+ $X2=1.41 $Y2=1.175
r46 7 10 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.425 $Y=0.58
+ $X2=1.425 $Y2=1.01
r47 3 12 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.395 $Y=2.4
+ $X2=1.395 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__CLKBUF_2%VPWR 1 2 7 9 13 15 17 24 25 31
r31 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r32 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 25 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r34 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r35 22 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.17 $Y2=3.33
r36 22 24 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.68 $Y2=3.33
r37 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r38 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 18 28 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.217 $Y2=3.33
r40 18 20 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.17 $Y2=3.33
r42 17 20 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 15 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.2 $Y2=3.33
r44 15 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 11 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=3.33
r46 11 13 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=2.78
r47 7 28 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.217 $Y2=3.33
r48 7 9 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.27 $Y=3.245 $X2=0.27
+ $Y2=2.78
r49 2 13 600 $w=1.7e-07 $l=1.00524e-06 $layer=licon1_PDIFF $count=1 $X=1.035
+ $Y=1.84 $X2=1.17 $Y2=2.78
r50 1 9 600 $w=1.7e-07 $l=1.00524e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_MS__CLKBUF_2%X 1 2 10 11 13
r28 13 19 10.8446 $w=3.38e-07 $l=2.35e-07 $layer=LI1_cond $X=0.715 $Y=0.555
+ $X2=0.715 $Y2=0.79
r29 11 19 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=0.8 $Y=1.82 $X2=0.8
+ $Y2=0.79
r30 10 11 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.72 $Y=1.985
+ $X2=0.72 $Y2=1.82
r31 2 10 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.84 $X2=0.72 $Y2=1.985
r32 1 13 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_MS__CLKBUF_2%VGND 1 2 7 9 13 15 17 24 25 31
r27 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r28 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r29 25 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r30 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r31 22 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.18
+ $Y2=0
r32 22 24 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.68
+ $Y2=0
r33 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r34 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r35 18 28 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r36 18 20 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.72
+ $Y2=0
r37 17 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.18
+ $Y2=0
r38 17 20 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=0.72
+ $Y2=0
r39 15 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r40 15 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r41 11 31 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.18 $Y2=0
r42 11 13 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.18 $Y2=0.58
r43 7 28 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r44 7 9 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.57
r45 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1 $Y=0.37
+ $X2=1.14 $Y2=0.58
r46 1 9 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.57
.ends


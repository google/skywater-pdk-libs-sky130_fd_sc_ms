# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__dlrbp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__dlrbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.233700 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.450000 0.805000 1.780000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.150000 0.350000 6.480000 0.960000 ;
        RECT 6.150000 0.960000 7.075000 1.130000 ;
        RECT 6.295000 1.800000 7.075000 1.970000 ;
        RECT 6.295000 1.970000 6.465000 2.980000 ;
        RECT 6.845000 1.130000 7.075000 1.800000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.225000 1.820000 8.585000 2.980000 ;
        RECT 8.245000 0.350000 8.585000 1.130000 ;
        RECT 8.415000 1.130000 8.585000 1.820000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.435000 1.180000 5.785000 1.550000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.262200 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.975000 1.180000 1.285000 1.550000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.120000 0.085000 ;
        RECT 0.625000  0.085000 0.955000 1.010000 ;
        RECT 2.305000  0.085000 2.640000 0.410000 ;
        RECT 4.230000  0.085000 4.560000 1.060000 ;
        RECT 5.610000  0.085000 5.940000 1.010000 ;
        RECT 6.650000  0.085000 6.980000 0.790000 ;
        RECT 7.745000  0.085000 8.075000 1.130000 ;
        RECT 8.755000  0.085000 9.005000 1.130000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
        RECT 8.315000 -0.085000 8.485000 0.085000 ;
        RECT 8.795000 -0.085000 8.965000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 9.120000 3.415000 ;
        RECT 0.650000 2.700000 0.980000 3.245000 ;
        RECT 2.330000 2.700000 2.695000 3.245000 ;
        RECT 4.425000 2.650000 5.065000 3.245000 ;
        RECT 5.735000 2.060000 6.065000 3.245000 ;
        RECT 6.665000 2.140000 6.995000 3.245000 ;
        RECT 7.725000 1.820000 8.055000 3.245000 ;
        RECT 8.755000 1.820000 9.005000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
        RECT 8.315000 3.245000 8.485000 3.415000 ;
        RECT 8.795000 3.245000 8.965000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.540000 0.445000 1.130000 ;
      RECT 0.085000 1.130000 0.255000 1.950000 ;
      RECT 0.085000 1.950000 0.445000 2.360000 ;
      RECT 0.085000 2.360000 2.805000 2.530000 ;
      RECT 0.085000 2.530000 0.445000 2.820000 ;
      RECT 1.125000 0.350000 1.625000 0.580000 ;
      RECT 1.125000 0.580000 2.980000 0.750000 ;
      RECT 1.125000 0.750000 1.625000 1.010000 ;
      RECT 1.185000 1.940000 1.625000 2.190000 ;
      RECT 1.455000 1.010000 1.625000 1.340000 ;
      RECT 1.455000 1.340000 1.865000 1.670000 ;
      RECT 1.455000 1.670000 1.625000 1.940000 ;
      RECT 1.795000 0.920000 2.205000 1.130000 ;
      RECT 1.795000 1.130000 3.385000 1.170000 ;
      RECT 1.795000 1.940000 2.205000 2.190000 ;
      RECT 2.035000 1.170000 3.385000 1.300000 ;
      RECT 2.035000 1.300000 2.205000 1.940000 ;
      RECT 2.485000 1.470000 2.805000 2.360000 ;
      RECT 2.810000 0.255000 3.895000 0.510000 ;
      RECT 2.810000 0.510000 2.980000 0.580000 ;
      RECT 2.975000 1.300000 3.385000 1.480000 ;
      RECT 2.975000 1.480000 3.145000 2.905000 ;
      RECT 2.975000 2.905000 4.035000 3.075000 ;
      RECT 3.180000 0.790000 3.740000 0.960000 ;
      RECT 3.315000 1.650000 4.925000 1.820000 ;
      RECT 3.315000 1.820000 3.485000 2.735000 ;
      RECT 3.570000 0.960000 3.740000 1.650000 ;
      RECT 3.705000 2.050000 4.035000 2.905000 ;
      RECT 4.245000 1.990000 5.565000 2.320000 ;
      RECT 4.605000 1.350000 4.925000 1.650000 ;
      RECT 4.790000 0.350000 5.265000 1.130000 ;
      RECT 5.095000 1.130000 5.265000 1.720000 ;
      RECT 5.095000 1.720000 6.125000 1.890000 ;
      RECT 5.095000 1.890000 5.565000 1.990000 ;
      RECT 5.235000 2.320000 5.565000 2.980000 ;
      RECT 5.955000 1.300000 6.650000 1.630000 ;
      RECT 5.955000 1.630000 6.125000 1.720000 ;
      RECT 7.245000 0.450000 7.575000 1.130000 ;
      RECT 7.245000 1.130000 7.555000 1.300000 ;
      RECT 7.245000 1.300000 8.245000 1.630000 ;
      RECT 7.245000 1.630000 7.555000 2.860000 ;
  END
END sky130_fd_sc_ms__dlrbp_2

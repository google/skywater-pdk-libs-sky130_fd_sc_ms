* File: sky130_fd_sc_ms__or3b_1.pxi.spice
* Created: Wed Sep  2 12:28:30 2020
* 
x_PM_SKY130_FD_SC_MS__OR3B_1%C_N N_C_N_c_75_n N_C_N_M1008_g N_C_N_M1007_g
+ N_C_N_c_77_n C_N C_N N_C_N_c_78_n N_C_N_c_79_n PM_SKY130_FD_SC_MS__OR3B_1%C_N
x_PM_SKY130_FD_SC_MS__OR3B_1%A_127_74# N_A_127_74#_M1007_d N_A_127_74#_M1008_d
+ N_A_127_74#_c_108_n N_A_127_74#_c_109_n N_A_127_74#_c_117_n
+ N_A_127_74#_c_118_n N_A_127_74#_M1004_g N_A_127_74#_c_119_n
+ N_A_127_74#_M1009_g N_A_127_74#_c_111_n N_A_127_74#_c_120_n
+ N_A_127_74#_c_112_n N_A_127_74#_c_113_n N_A_127_74#_c_121_n
+ N_A_127_74#_c_114_n N_A_127_74#_c_115_n N_A_127_74#_c_116_n
+ N_A_127_74#_c_123_n PM_SKY130_FD_SC_MS__OR3B_1%A_127_74#
x_PM_SKY130_FD_SC_MS__OR3B_1%B N_B_M1000_g N_B_c_169_n N_B_M1001_g B B B B
+ N_B_c_171_n PM_SKY130_FD_SC_MS__OR3B_1%B
x_PM_SKY130_FD_SC_MS__OR3B_1%A N_A_M1002_g N_A_M1005_g A N_A_c_210_n N_A_c_211_n
+ PM_SKY130_FD_SC_MS__OR3B_1%A
x_PM_SKY130_FD_SC_MS__OR3B_1%A_239_74# N_A_239_74#_M1004_s N_A_239_74#_M1000_d
+ N_A_239_74#_M1009_s N_A_239_74#_M1003_g N_A_239_74#_M1006_g
+ N_A_239_74#_c_245_n N_A_239_74#_c_246_n N_A_239_74#_c_247_n
+ N_A_239_74#_c_248_n N_A_239_74#_c_249_n N_A_239_74#_c_250_n
+ N_A_239_74#_c_251_n N_A_239_74#_c_252_n N_A_239_74#_c_253_n
+ N_A_239_74#_c_254_n PM_SKY130_FD_SC_MS__OR3B_1%A_239_74#
x_PM_SKY130_FD_SC_MS__OR3B_1%VPWR N_VPWR_M1008_s N_VPWR_M1005_d N_VPWR_c_336_n
+ N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n N_VPWR_c_340_n VPWR
+ N_VPWR_c_341_n N_VPWR_c_335_n PM_SKY130_FD_SC_MS__OR3B_1%VPWR
x_PM_SKY130_FD_SC_MS__OR3B_1%X N_X_M1006_d N_X_M1003_d N_X_c_375_n N_X_c_376_n
+ N_X_c_372_n X X X PM_SKY130_FD_SC_MS__OR3B_1%X
x_PM_SKY130_FD_SC_MS__OR3B_1%VGND N_VGND_M1007_s N_VGND_M1004_d N_VGND_M1002_d
+ N_VGND_c_397_n N_VGND_c_398_n N_VGND_c_399_n N_VGND_c_400_n VGND
+ N_VGND_c_401_n N_VGND_c_402_n N_VGND_c_403_n N_VGND_c_404_n N_VGND_c_405_n
+ N_VGND_c_406_n PM_SKY130_FD_SC_MS__OR3B_1%VGND
cc_1 VNB N_C_N_c_75_n 0.0260596f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.6
cc_2 VNB N_C_N_M1007_g 0.0316419f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.645
cc_3 VNB N_C_N_c_77_n 0.00507655f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.78
cc_4 VNB N_C_N_c_78_n 0.0218412f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=1.275
cc_5 VNB N_C_N_c_79_n 0.0261056f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=1.275
cc_6 VNB N_A_127_74#_c_108_n 0.0232951f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.11
cc_7 VNB N_A_127_74#_c_109_n 0.0163801f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=0.645
cc_8 VNB N_A_127_74#_M1004_g 0.0337631f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_9 VNB N_A_127_74#_c_111_n 0.00648012f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.295
cc_10 VNB N_A_127_74#_c_112_n 0.00141058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_127_74#_c_113_n 0.00714418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_127_74#_c_114_n 0.0109289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_127_74#_c_115_n 0.0189698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_127_74#_c_116_n 0.00472452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_M1000_g 0.0276545f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.78
cc_16 VNB N_B_c_169_n 0.0404634f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.54
cc_17 VNB N_B_M1001_g 0.00319841f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.11
cc_18 VNB N_B_c_171_n 0.00612656f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.11
cc_19 VNB N_A_M1002_g 0.0365472f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.78
cc_20 VNB N_A_M1005_g 0.00157694f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.11
cc_21 VNB N_A_c_210_n 0.0329279f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_22 VNB N_A_c_211_n 0.00235452f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_23 VNB N_A_239_74#_M1003_g 0.0019512f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_24 VNB N_A_239_74#_M1006_g 0.0301771f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.275
cc_25 VNB N_A_239_74#_c_245_n 0.0071094f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.275
cc_26 VNB N_A_239_74#_c_246_n 0.0101214f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.665
cc_27 VNB N_A_239_74#_c_247_n 0.00821763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_239_74#_c_248_n 0.00280782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_239_74#_c_249_n 0.00833839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_239_74#_c_250_n 0.00380922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_239_74#_c_251_n 0.00406482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_239_74#_c_252_n 0.00983809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_239_74#_c_253_n 0.00276147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_239_74#_c_254_n 0.0344827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VPWR_c_335_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_X_c_372_n 0.0247788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB X 0.0265914f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.275
cc_38 VNB X 0.0139041f $X=-0.19 $Y=-0.245 $X2=0.44 $Y2=1.275
cc_39 VNB N_VGND_c_397_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_398_n 0.0379781f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_41 VNB N_VGND_c_399_n 0.00900728f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.275
cc_42 VNB N_VGND_c_400_n 0.0114492f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.275
cc_43 VNB N_VGND_c_401_n 0.0339528f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.665
cc_44 VNB N_VGND_c_402_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_403_n 0.0189171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_404_n 0.232138f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_405_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_406_n 0.0105791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VPB N_C_N_M1008_g 0.0478973f $X=-0.19 $Y=1.66 $X2=0.545 $Y2=2.54
cc_50 VPB N_C_N_c_77_n 0.0152909f $X=-0.19 $Y=1.66 $X2=0.455 $Y2=1.78
cc_51 VPB N_C_N_c_79_n 0.00895383f $X=-0.19 $Y=1.66 $X2=0.44 $Y2=1.275
cc_52 VPB N_A_127_74#_c_117_n 0.0477998f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.645
cc_53 VPB N_A_127_74#_c_118_n 0.0163801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_127_74#_c_119_n 0.0215139f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_127_74#_c_120_n 0.0212506f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_127_74#_c_121_n 0.0047323f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_127_74#_c_115_n 0.0031572f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_127_74#_c_123_n 0.012278f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_B_M1001_g 0.0285357f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=1.11
cc_60 VPB N_B_c_171_n 0.00211217f $X=-0.19 $Y=1.66 $X2=0.455 $Y2=1.11
cc_61 VPB N_A_M1005_g 0.0309676f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=1.11
cc_62 VPB N_A_c_211_n 0.00438681f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_63 VPB N_A_239_74#_M1003_g 0.0307264f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_64 VPB N_A_239_74#_c_246_n 0.0194148f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.665
cc_65 VPB N_VPWR_c_336_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=1.11
cc_66 VPB N_VPWR_c_337_n 0.0498598f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.645
cc_67 VPB N_VPWR_c_338_n 0.0100179f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_68 VPB N_VPWR_c_339_n 0.0658301f $X=-0.19 $Y=1.66 $X2=0.44 $Y2=1.275
cc_69 VPB N_VPWR_c_340_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.455 $Y2=1.11
cc_70 VPB N_VPWR_c_341_n 0.0223986f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_335_n 0.0896543f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_X_c_375_n 0.0462568f $X=-0.19 $Y=1.66 $X2=0.56 $Y2=0.645
cc_73 VPB N_X_c_376_n 0.0194191f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_X_c_372_n 0.00789123f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 N_C_N_c_78_n N_A_127_74#_c_109_n 0.0116947f $X=0.44 $Y=1.275 $X2=0 $Y2=0
cc_76 N_C_N_c_79_n N_A_127_74#_c_109_n 5.66699e-19 $X=0.44 $Y=1.275 $X2=0 $Y2=0
cc_77 N_C_N_c_77_n N_A_127_74#_c_118_n 0.0116947f $X=0.455 $Y=1.78 $X2=0 $Y2=0
cc_78 N_C_N_M1007_g N_A_127_74#_c_111_n 0.00659399f $X=0.56 $Y=0.645 $X2=0 $Y2=0
cc_79 N_C_N_M1008_g N_A_127_74#_c_120_n 0.0149079f $X=0.545 $Y=2.54 $X2=0 $Y2=0
cc_80 N_C_N_c_75_n N_A_127_74#_c_112_n 0.00380448f $X=0.455 $Y=1.6 $X2=0 $Y2=0
cc_81 N_C_N_M1007_g N_A_127_74#_c_113_n 0.00470727f $X=0.56 $Y=0.645 $X2=0 $Y2=0
cc_82 N_C_N_M1008_g N_A_127_74#_c_121_n 0.00380448f $X=0.545 $Y=2.54 $X2=0 $Y2=0
cc_83 N_C_N_c_78_n N_A_127_74#_c_114_n 0.00380448f $X=0.44 $Y=1.275 $X2=0 $Y2=0
cc_84 N_C_N_c_75_n N_A_127_74#_c_115_n 0.0116947f $X=0.455 $Y=1.6 $X2=0 $Y2=0
cc_85 N_C_N_M1007_g N_A_127_74#_c_116_n 0.00380448f $X=0.56 $Y=0.645 $X2=0 $Y2=0
cc_86 N_C_N_c_79_n N_A_127_74#_c_116_n 0.0548703f $X=0.44 $Y=1.275 $X2=0 $Y2=0
cc_87 N_C_N_c_77_n N_A_127_74#_c_123_n 0.00380448f $X=0.455 $Y=1.78 $X2=0 $Y2=0
cc_88 N_C_N_M1007_g N_A_239_74#_c_245_n 0.00109764f $X=0.56 $Y=0.645 $X2=0 $Y2=0
cc_89 N_C_N_M1007_g N_A_239_74#_c_251_n 0.00111956f $X=0.56 $Y=0.645 $X2=0 $Y2=0
cc_90 N_C_N_M1008_g N_VPWR_c_337_n 0.00925233f $X=0.545 $Y=2.54 $X2=0 $Y2=0
cc_91 N_C_N_c_77_n N_VPWR_c_337_n 0.00122656f $X=0.455 $Y=1.78 $X2=0 $Y2=0
cc_92 N_C_N_c_79_n N_VPWR_c_337_n 0.0183299f $X=0.44 $Y=1.275 $X2=0 $Y2=0
cc_93 N_C_N_M1008_g N_VPWR_c_339_n 0.0053223f $X=0.545 $Y=2.54 $X2=0 $Y2=0
cc_94 N_C_N_M1008_g N_VPWR_c_335_n 0.0102706f $X=0.545 $Y=2.54 $X2=0 $Y2=0
cc_95 N_C_N_M1007_g N_VGND_c_398_n 0.0162837f $X=0.56 $Y=0.645 $X2=0 $Y2=0
cc_96 N_C_N_c_78_n N_VGND_c_398_n 0.00132308f $X=0.44 $Y=1.275 $X2=0 $Y2=0
cc_97 N_C_N_c_79_n N_VGND_c_398_n 0.0289964f $X=0.44 $Y=1.275 $X2=0 $Y2=0
cc_98 N_C_N_M1007_g N_VGND_c_401_n 0.00439937f $X=0.56 $Y=0.645 $X2=0 $Y2=0
cc_99 N_C_N_M1007_g N_VGND_c_404_n 0.00847151f $X=0.56 $Y=0.645 $X2=0 $Y2=0
cc_100 N_A_127_74#_M1004_g N_B_M1000_g 0.0210899f $X=1.555 $Y=0.645 $X2=0 $Y2=0
cc_101 N_A_127_74#_M1004_g N_B_c_169_n 0.00720842f $X=1.555 $Y=0.645 $X2=0 $Y2=0
cc_102 N_A_127_74#_c_115_n N_B_c_169_n 6.62475e-19 $X=1.04 $Y=1.375 $X2=0 $Y2=0
cc_103 N_A_127_74#_c_117_n N_B_M1001_g 0.069654f $X=1.675 $Y=1.805 $X2=0 $Y2=0
cc_104 N_A_127_74#_c_117_n N_B_c_171_n 0.00919075f $X=1.675 $Y=1.805 $X2=0 $Y2=0
cc_105 N_A_127_74#_M1004_g N_A_239_74#_c_245_n 0.00929209f $X=1.555 $Y=0.645
+ $X2=0 $Y2=0
cc_106 N_A_127_74#_c_111_n N_A_239_74#_c_245_n 0.0336418f $X=0.78 $Y=0.645 $X2=0
+ $Y2=0
cc_107 N_A_127_74#_c_108_n N_A_239_74#_c_246_n 0.0127495f $X=1.48 $Y=1.285 $X2=0
+ $Y2=0
cc_108 N_A_127_74#_c_117_n N_A_239_74#_c_246_n 0.020889f $X=1.675 $Y=1.805 $X2=0
+ $Y2=0
cc_109 N_A_127_74#_M1004_g N_A_239_74#_c_246_n 0.00721297f $X=1.555 $Y=0.645
+ $X2=0 $Y2=0
cc_110 N_A_127_74#_c_119_n N_A_239_74#_c_246_n 0.0158808f $X=1.765 $Y=1.88 $X2=0
+ $Y2=0
cc_111 N_A_127_74#_c_121_n N_A_239_74#_c_246_n 0.0477325f $X=0.78 $Y=2.1 $X2=0
+ $Y2=0
cc_112 N_A_127_74#_c_114_n N_A_239_74#_c_246_n 0.0526809f $X=1.04 $Y=1.375 $X2=0
+ $Y2=0
cc_113 N_A_127_74#_c_115_n N_A_239_74#_c_246_n 0.00351858f $X=1.04 $Y=1.375
+ $X2=0 $Y2=0
cc_114 N_A_127_74#_c_116_n N_A_239_74#_c_246_n 0.00789174f $X=0.99 $Y=1.21 $X2=0
+ $Y2=0
cc_115 N_A_127_74#_M1004_g N_A_239_74#_c_248_n 5.97046e-19 $X=1.555 $Y=0.645
+ $X2=0 $Y2=0
cc_116 N_A_127_74#_c_109_n N_A_239_74#_c_251_n 0.00702615f $X=1.205 $Y=1.285
+ $X2=0 $Y2=0
cc_117 N_A_127_74#_M1004_g N_A_239_74#_c_251_n 0.0119206f $X=1.555 $Y=0.645
+ $X2=0 $Y2=0
cc_118 N_A_127_74#_c_113_n N_A_239_74#_c_251_n 0.0122227f $X=0.78 $Y=0.94 $X2=0
+ $Y2=0
cc_119 N_A_127_74#_c_114_n N_A_239_74#_c_251_n 0.00237099f $X=1.04 $Y=1.375
+ $X2=0 $Y2=0
cc_120 N_A_127_74#_c_120_n N_VPWR_c_337_n 0.0345631f $X=0.78 $Y=2.265 $X2=0
+ $Y2=0
cc_121 N_A_127_74#_c_119_n N_VPWR_c_339_n 0.00516426f $X=1.765 $Y=1.88 $X2=0
+ $Y2=0
cc_122 N_A_127_74#_c_120_n N_VPWR_c_339_n 0.0145789f $X=0.78 $Y=2.265 $X2=0
+ $Y2=0
cc_123 N_A_127_74#_c_119_n N_VPWR_c_335_n 0.00653145f $X=1.765 $Y=1.88 $X2=0
+ $Y2=0
cc_124 N_A_127_74#_c_120_n N_VPWR_c_335_n 0.0120225f $X=0.78 $Y=2.265 $X2=0
+ $Y2=0
cc_125 N_A_127_74#_c_111_n N_VGND_c_398_n 0.0236817f $X=0.78 $Y=0.645 $X2=0
+ $Y2=0
cc_126 N_A_127_74#_M1004_g N_VGND_c_399_n 0.00525427f $X=1.555 $Y=0.645 $X2=0
+ $Y2=0
cc_127 N_A_127_74#_M1004_g N_VGND_c_401_n 0.00434272f $X=1.555 $Y=0.645 $X2=0
+ $Y2=0
cc_128 N_A_127_74#_c_111_n N_VGND_c_401_n 0.0145071f $X=0.78 $Y=0.645 $X2=0
+ $Y2=0
cc_129 N_A_127_74#_M1004_g N_VGND_c_404_n 0.00452955f $X=1.555 $Y=0.645 $X2=0
+ $Y2=0
cc_130 N_A_127_74#_c_111_n N_VGND_c_404_n 0.0119944f $X=0.78 $Y=0.645 $X2=0
+ $Y2=0
cc_131 N_B_M1000_g N_A_M1002_g 0.0220773f $X=2.125 $Y=0.645 $X2=0 $Y2=0
cc_132 N_B_c_169_n N_A_M1002_g 0.0148343f $X=2.185 $Y=1.61 $X2=0 $Y2=0
cc_133 N_B_c_171_n N_A_M1002_g 0.00384055f $X=2.08 $Y=1.355 $X2=0 $Y2=0
cc_134 N_B_M1001_g N_A_M1005_g 0.0395829f $X=2.185 $Y=2.455 $X2=0 $Y2=0
cc_135 N_B_c_169_n N_A_c_210_n 0.0395829f $X=2.185 $Y=1.61 $X2=0 $Y2=0
cc_136 N_B_c_171_n N_A_c_210_n 0.00559495f $X=2.08 $Y=1.355 $X2=0 $Y2=0
cc_137 N_B_c_169_n N_A_c_211_n 0.00112073f $X=2.185 $Y=1.61 $X2=0 $Y2=0
cc_138 N_B_c_171_n N_A_c_211_n 0.0284132f $X=2.08 $Y=1.355 $X2=0 $Y2=0
cc_139 N_B_M1000_g N_A_239_74#_c_245_n 5.97046e-19 $X=2.125 $Y=0.645 $X2=0 $Y2=0
cc_140 N_B_M1000_g N_A_239_74#_c_246_n 0.00341621f $X=2.125 $Y=0.645 $X2=0 $Y2=0
cc_141 N_B_c_169_n N_A_239_74#_c_246_n 0.00491731f $X=2.185 $Y=1.61 $X2=0 $Y2=0
cc_142 N_B_M1001_g N_A_239_74#_c_246_n 0.0012981f $X=2.185 $Y=2.455 $X2=0 $Y2=0
cc_143 N_B_c_171_n N_A_239_74#_c_246_n 0.115003f $X=2.08 $Y=1.355 $X2=0 $Y2=0
cc_144 N_B_M1000_g N_A_239_74#_c_247_n 0.00920125f $X=2.125 $Y=0.645 $X2=0 $Y2=0
cc_145 N_B_c_169_n N_A_239_74#_c_247_n 9.4463e-19 $X=2.185 $Y=1.61 $X2=0 $Y2=0
cc_146 N_B_c_171_n N_A_239_74#_c_247_n 0.0201966f $X=2.08 $Y=1.355 $X2=0 $Y2=0
cc_147 N_B_M1000_g N_A_239_74#_c_248_n 0.00831927f $X=2.125 $Y=0.645 $X2=0 $Y2=0
cc_148 N_B_M1000_g N_A_239_74#_c_252_n 0.00293078f $X=2.125 $Y=0.645 $X2=0 $Y2=0
cc_149 N_B_c_169_n N_A_239_74#_c_252_n 4.61596e-19 $X=2.185 $Y=1.61 $X2=0 $Y2=0
cc_150 N_B_c_171_n N_A_239_74#_c_252_n 0.00883544f $X=2.08 $Y=1.355 $X2=0 $Y2=0
cc_151 N_B_c_171_n N_VPWR_c_338_n 0.015575f $X=2.08 $Y=1.355 $X2=0 $Y2=0
cc_152 N_B_M1001_g N_VPWR_c_339_n 0.00361543f $X=2.185 $Y=2.455 $X2=0 $Y2=0
cc_153 N_B_c_171_n N_VPWR_c_339_n 0.0102024f $X=2.08 $Y=1.355 $X2=0 $Y2=0
cc_154 N_B_M1001_g N_VPWR_c_335_n 0.00653145f $X=2.185 $Y=2.455 $X2=0 $Y2=0
cc_155 N_B_c_171_n N_VPWR_c_335_n 0.0115903f $X=2.08 $Y=1.355 $X2=0 $Y2=0
cc_156 N_B_c_171_n A_371_391# 0.0101478f $X=2.08 $Y=1.355 $X2=-0.19 $Y2=-0.245
cc_157 N_B_M1000_g N_VGND_c_399_n 0.00387235f $X=2.125 $Y=0.645 $X2=0 $Y2=0
cc_158 N_B_M1000_g N_VGND_c_402_n 0.00434272f $X=2.125 $Y=0.645 $X2=0 $Y2=0
cc_159 N_B_M1000_g N_VGND_c_404_n 0.00448578f $X=2.125 $Y=0.645 $X2=0 $Y2=0
cc_160 N_A_M1005_g N_A_239_74#_M1003_g 0.0218657f $X=2.605 $Y=2.455 $X2=0 $Y2=0
cc_161 N_A_c_211_n N_A_239_74#_M1003_g 0.00337622f $X=2.68 $Y=1.465 $X2=0 $Y2=0
cc_162 N_A_M1002_g N_A_239_74#_M1006_g 0.0141364f $X=2.59 $Y=0.645 $X2=0 $Y2=0
cc_163 N_A_M1002_g N_A_239_74#_c_248_n 6.3123e-19 $X=2.59 $Y=0.645 $X2=0 $Y2=0
cc_164 N_A_M1002_g N_A_239_74#_c_249_n 0.0138558f $X=2.59 $Y=0.645 $X2=0 $Y2=0
cc_165 N_A_c_210_n N_A_239_74#_c_249_n 0.00113397f $X=2.68 $Y=1.465 $X2=0 $Y2=0
cc_166 N_A_c_211_n N_A_239_74#_c_249_n 0.0169506f $X=2.68 $Y=1.465 $X2=0 $Y2=0
cc_167 N_A_M1002_g N_A_239_74#_c_250_n 0.00504171f $X=2.59 $Y=0.645 $X2=0 $Y2=0
cc_168 N_A_c_210_n N_A_239_74#_c_253_n 0.00201625f $X=2.68 $Y=1.465 $X2=0 $Y2=0
cc_169 N_A_c_211_n N_A_239_74#_c_253_n 0.0224088f $X=2.68 $Y=1.465 $X2=0 $Y2=0
cc_170 N_A_c_210_n N_A_239_74#_c_254_n 0.0175372f $X=2.68 $Y=1.465 $X2=0 $Y2=0
cc_171 N_A_c_211_n N_A_239_74#_c_254_n 3.95231e-19 $X=2.68 $Y=1.465 $X2=0 $Y2=0
cc_172 N_A_M1005_g N_VPWR_c_338_n 0.00981917f $X=2.605 $Y=2.455 $X2=0 $Y2=0
cc_173 N_A_c_210_n N_VPWR_c_338_n 5.13337e-19 $X=2.68 $Y=1.465 $X2=0 $Y2=0
cc_174 N_A_c_211_n N_VPWR_c_338_n 0.00836062f $X=2.68 $Y=1.465 $X2=0 $Y2=0
cc_175 N_A_M1005_g N_VPWR_c_339_n 0.005489f $X=2.605 $Y=2.455 $X2=0 $Y2=0
cc_176 N_A_M1005_g N_VPWR_c_335_n 0.00653145f $X=2.605 $Y=2.455 $X2=0 $Y2=0
cc_177 N_A_M1005_g N_X_c_376_n 7.81367e-19 $X=2.605 $Y=2.455 $X2=0 $Y2=0
cc_178 N_A_M1002_g N_VGND_c_400_n 0.00526056f $X=2.59 $Y=0.645 $X2=0 $Y2=0
cc_179 N_A_M1002_g N_VGND_c_402_n 0.00461464f $X=2.59 $Y=0.645 $X2=0 $Y2=0
cc_180 N_A_M1002_g N_VGND_c_404_n 0.00467888f $X=2.59 $Y=0.645 $X2=0 $Y2=0
cc_181 N_A_239_74#_M1003_g N_VPWR_c_338_n 0.00355945f $X=3.19 $Y=2.4 $X2=0 $Y2=0
cc_182 N_A_239_74#_c_246_n N_VPWR_c_339_n 0.0142618f $X=1.54 $Y=2.1 $X2=0 $Y2=0
cc_183 N_A_239_74#_M1003_g N_VPWR_c_341_n 0.005209f $X=3.19 $Y=2.4 $X2=0 $Y2=0
cc_184 N_A_239_74#_M1003_g N_VPWR_c_335_n 0.00990877f $X=3.19 $Y=2.4 $X2=0 $Y2=0
cc_185 N_A_239_74#_c_246_n N_VPWR_c_335_n 0.0119375f $X=1.54 $Y=2.1 $X2=0 $Y2=0
cc_186 N_A_239_74#_M1003_g N_X_c_375_n 0.0121628f $X=3.19 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A_239_74#_M1003_g N_X_c_376_n 0.00512884f $X=3.19 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A_239_74#_c_253_n N_X_c_376_n 0.0125883f $X=3.25 $Y=1.465 $X2=0 $Y2=0
cc_189 N_A_239_74#_c_254_n N_X_c_376_n 0.00387134f $X=3.25 $Y=1.465 $X2=0 $Y2=0
cc_190 N_A_239_74#_M1003_g N_X_c_372_n 0.00422132f $X=3.19 $Y=2.4 $X2=0 $Y2=0
cc_191 N_A_239_74#_M1006_g N_X_c_372_n 0.0100339f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A_239_74#_c_250_n N_X_c_372_n 0.00535893f $X=3.14 $Y=1.3 $X2=0 $Y2=0
cc_193 N_A_239_74#_c_253_n N_X_c_372_n 0.0249377f $X=3.25 $Y=1.465 $X2=0 $Y2=0
cc_194 N_A_239_74#_M1006_g X 0.0138808f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_195 N_A_239_74#_M1006_g X 0.00282902f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A_239_74#_c_250_n X 0.00489765f $X=3.14 $Y=1.3 $X2=0 $Y2=0
cc_197 N_A_239_74#_c_253_n X 0.00151667f $X=3.25 $Y=1.465 $X2=0 $Y2=0
cc_198 N_A_239_74#_c_247_n N_VGND_M1004_d 0.00324086f $X=2.175 $Y=0.935 $X2=0
+ $Y2=0
cc_199 N_A_239_74#_c_249_n N_VGND_M1002_d 0.00894604f $X=3.055 $Y=0.935 $X2=0
+ $Y2=0
cc_200 N_A_239_74#_c_250_n N_VGND_M1002_d 0.00201508f $X=3.14 $Y=1.3 $X2=0 $Y2=0
cc_201 N_A_239_74#_c_245_n N_VGND_c_399_n 0.0131729f $X=1.34 $Y=0.645 $X2=0
+ $Y2=0
cc_202 N_A_239_74#_c_247_n N_VGND_c_399_n 0.0229024f $X=2.175 $Y=0.935 $X2=0
+ $Y2=0
cc_203 N_A_239_74#_c_248_n N_VGND_c_399_n 0.0131729f $X=2.34 $Y=0.645 $X2=0
+ $Y2=0
cc_204 N_A_239_74#_c_251_n N_VGND_c_399_n 0.00158528f $X=1.44 $Y=0.935 $X2=0
+ $Y2=0
cc_205 N_A_239_74#_M1006_g N_VGND_c_400_n 0.00646208f $X=3.345 $Y=0.74 $X2=0
+ $Y2=0
cc_206 N_A_239_74#_c_248_n N_VGND_c_400_n 0.00164437f $X=2.34 $Y=0.645 $X2=0
+ $Y2=0
cc_207 N_A_239_74#_c_249_n N_VGND_c_400_n 0.0400007f $X=3.055 $Y=0.935 $X2=0
+ $Y2=0
cc_208 N_A_239_74#_c_254_n N_VGND_c_400_n 4.27896e-19 $X=3.25 $Y=1.465 $X2=0
+ $Y2=0
cc_209 N_A_239_74#_c_245_n N_VGND_c_401_n 0.0145543f $X=1.34 $Y=0.645 $X2=0
+ $Y2=0
cc_210 N_A_239_74#_c_248_n N_VGND_c_402_n 0.0145482f $X=2.34 $Y=0.645 $X2=0
+ $Y2=0
cc_211 N_A_239_74#_M1006_g N_VGND_c_403_n 0.00434272f $X=3.345 $Y=0.74 $X2=0
+ $Y2=0
cc_212 N_A_239_74#_M1006_g N_VGND_c_404_n 0.00826108f $X=3.345 $Y=0.74 $X2=0
+ $Y2=0
cc_213 N_A_239_74#_c_245_n N_VGND_c_404_n 0.0119947f $X=1.34 $Y=0.645 $X2=0
+ $Y2=0
cc_214 N_A_239_74#_c_247_n N_VGND_c_404_n 0.00589553f $X=2.175 $Y=0.935 $X2=0
+ $Y2=0
cc_215 N_A_239_74#_c_248_n N_VGND_c_404_n 0.0119922f $X=2.34 $Y=0.645 $X2=0
+ $Y2=0
cc_216 N_A_239_74#_c_249_n N_VGND_c_404_n 0.00654887f $X=3.055 $Y=0.935 $X2=0
+ $Y2=0
cc_217 N_A_239_74#_c_251_n N_VGND_c_404_n 0.00582685f $X=1.44 $Y=0.935 $X2=0
+ $Y2=0
cc_218 N_VPWR_c_341_n N_X_c_375_n 0.0223576f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_219 N_VPWR_c_335_n N_X_c_375_n 0.0184376f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_220 N_VPWR_c_338_n N_X_c_376_n 0.0419968f $X=2.915 $Y=2.115 $X2=0 $Y2=0
cc_221 X N_VGND_c_400_n 0.0134023f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_222 X N_VGND_c_403_n 0.0159025f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_223 X N_VGND_c_404_n 0.0131064f $X=3.515 $Y=0.47 $X2=0 $Y2=0

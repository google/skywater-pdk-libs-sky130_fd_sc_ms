* NGSPICE file created from sky130_fd_sc_ms__and3b_4.ext - technology: sky130A

.subckt sky130_fd_sc_ms__and3b_4 A_N B C VGND VNB VPB VPWR X
M1000 VPWR A_N a_27_74# VPB pshort w=1e+06u l=180000u
+  ad=2.3986e+12p pd=1.727e+07u as=2.8e+11p ps=2.56e+06u
M1001 VPWR a_301_368# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=6.048e+11p ps=5.56e+06u
M1002 a_239_98# a_27_74# a_301_368# VNB nlowvt w=640000u l=150000u
+  ad=5.44e+11p pd=5.54e+06u as=1.792e+11p ps=1.84e+06u
M1003 a_498_98# C VGND VNB nlowvt w=640000u l=150000u
+  ad=4.032e+11p pd=3.82e+06u as=1.063e+12p ps=1.005e+07u
M1004 VGND a_301_368# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.662e+11p ps=4.22e+06u
M1005 a_301_368# C VPWR VPB pshort w=1e+06u l=180000u
+  ad=8.1e+11p pd=7.62e+06u as=0p ps=0u
M1006 VPWR C a_301_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_301_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_301_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND C a_498_98# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_239_98# B a_498_98# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_498_98# B a_239_98# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_301_368# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_301_368# a_27_74# a_239_98# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_301_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_301_368# B VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_301_368# a_27_74# VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_301_368# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A_N a_27_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1019 VPWR B a_301_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_27_74# a_301_368# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_301_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__nor2_2.pxi.spice
* Created: Wed Sep  2 12:15:18 2020
* 
x_PM_SKY130_FD_SC_MS__NOR2_2%B N_B_M1002_g N_B_M1001_g N_B_c_41_n N_B_c_46_n
+ N_B_M1003_g N_B_c_42_n N_B_c_43_n N_B_c_48_n B PM_SKY130_FD_SC_MS__NOR2_2%B
x_PM_SKY130_FD_SC_MS__NOR2_2%A N_A_c_79_n N_A_M1000_g N_A_c_80_n N_A_c_81_n
+ N_A_M1004_g N_A_M1005_g A A A N_A_c_86_n N_A_c_87_n N_A_c_88_n
+ PM_SKY130_FD_SC_MS__NOR2_2%A
x_PM_SKY130_FD_SC_MS__NOR2_2%A_35_368# N_A_35_368#_M1002_s N_A_35_368#_M1003_s
+ N_A_35_368#_M1005_s N_A_35_368#_c_125_n N_A_35_368#_c_126_n
+ N_A_35_368#_c_127_n N_A_35_368#_c_128_n N_A_35_368#_c_129_n
+ N_A_35_368#_c_130_n PM_SKY130_FD_SC_MS__NOR2_2%A_35_368#
x_PM_SKY130_FD_SC_MS__NOR2_2%Y N_Y_M1001_d N_Y_M1002_d N_Y_c_162_n Y Y Y
+ PM_SKY130_FD_SC_MS__NOR2_2%Y
x_PM_SKY130_FD_SC_MS__NOR2_2%VPWR N_VPWR_M1004_d N_VPWR_c_186_n N_VPWR_c_187_n
+ N_VPWR_c_188_n VPWR N_VPWR_c_189_n N_VPWR_c_185_n
+ PM_SKY130_FD_SC_MS__NOR2_2%VPWR
x_PM_SKY130_FD_SC_MS__NOR2_2%VGND N_VGND_M1001_s N_VGND_M1000_d N_VGND_c_211_n
+ N_VGND_c_212_n N_VGND_c_213_n VGND N_VGND_c_214_n N_VGND_c_215_n
+ N_VGND_c_216_n N_VGND_c_217_n PM_SKY130_FD_SC_MS__NOR2_2%VGND
cc_1 VNB N_B_c_41_n 0.0140858f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.69
cc_2 VNB N_B_c_42_n 0.0737008f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.385
cc_3 VNB N_B_c_43_n 0.0196224f $X=-0.19 $Y=-0.245 $X2=0.547 $Y2=1.22
cc_4 VNB B 0.0105321f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_5 VNB N_A_c_79_n 0.0173873f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.765
cc_6 VNB N_A_c_80_n 0.0177118f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.22
cc_7 VNB N_A_c_81_n 0.00722892f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.74
cc_8 VNB N_A_M1004_g 0.00408765f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.69
cc_9 VNB N_A_M1005_g 0.00454286f $X=-0.19 $Y=-0.245 $X2=0.547 $Y2=1.385
cc_10 VNB A 0.0193805f $X=-0.19 $Y=-0.245 $X2=0.547 $Y2=1.69
cc_11 VNB A 0.0201373f $X=-0.19 $Y=-0.245 $X2=0.547 $Y2=1.765
cc_12 VNB N_A_c_86_n 0.0955767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_c_87_n 0.0779857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_c_88_n 0.0251329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_Y_c_162_n 0.00598888f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.765
cc_16 VNB N_VPWR_c_185_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_211_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.69
cc_18 VNB N_VGND_c_212_n 0.0370023f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=1.765
cc_19 VNB N_VGND_c_213_n 0.0207786f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.385
cc_20 VNB N_VGND_c_214_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_21 VNB N_VGND_c_215_n 0.0282826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_216_n 0.174237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_217_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VPB N_B_c_41_n 0.00956914f $X=-0.19 $Y=1.66 $X2=0.905 $Y2=1.69
cc_25 VPB N_B_c_46_n 0.015741f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.765
cc_26 VPB N_B_c_42_n 0.00778644f $X=-0.19 $Y=1.66 $X2=0.455 $Y2=1.385
cc_27 VPB N_B_c_48_n 0.0195853f $X=-0.19 $Y=1.66 $X2=0.547 $Y2=1.765
cc_28 VPB N_A_M1004_g 0.0216644f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.69
cc_29 VPB N_A_M1005_g 0.0300699f $X=-0.19 $Y=1.66 $X2=0.547 $Y2=1.385
cc_30 VPB N_A_35_368#_c_125_n 0.0419632f $X=-0.19 $Y=1.66 $X2=0.547 $Y2=1.385
cc_31 VPB N_A_35_368#_c_126_n 0.00473643f $X=-0.19 $Y=1.66 $X2=0.547 $Y2=1.765
cc_32 VPB N_A_35_368#_c_127_n 0.00929469f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_33 VPB N_A_35_368#_c_128_n 0.0179802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_A_35_368#_c_129_n 0.00250101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_A_35_368#_c_130_n 0.0419012f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_186_n 0.00554449f $X=-0.19 $Y=1.66 $X2=0.565 $Y2=0.74
cc_37 VPB N_VPWR_c_187_n 0.038779f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=1.765
cc_38 VPB N_VPWR_c_188_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0.995 $Y2=2.4
cc_39 VPB N_VPWR_c_189_n 0.0201062f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.385
cc_40 VPB N_VPWR_c_185_n 0.05906f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 N_B_c_43_n N_A_c_79_n 0.00920383f $X=0.547 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_42 N_B_c_41_n N_A_c_81_n 0.0101464f $X=0.905 $Y=1.69 $X2=0 $Y2=0
cc_43 N_B_c_42_n N_A_c_81_n 0.00920383f $X=0.455 $Y=1.385 $X2=0 $Y2=0
cc_44 N_B_c_41_n N_A_M1004_g 0.0189209f $X=0.905 $Y=1.69 $X2=0 $Y2=0
cc_45 N_B_c_42_n N_A_c_87_n 0.00301438f $X=0.455 $Y=1.385 $X2=0 $Y2=0
cc_46 N_B_c_42_n N_A_35_368#_c_125_n 0.00185549f $X=0.455 $Y=1.385 $X2=0 $Y2=0
cc_47 N_B_c_48_n N_A_35_368#_c_125_n 0.00147311f $X=0.547 $Y=1.765 $X2=0 $Y2=0
cc_48 B N_A_35_368#_c_125_n 0.0149782f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_49 N_B_c_46_n N_A_35_368#_c_126_n 0.0133958f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_50 N_B_c_48_n N_A_35_368#_c_126_n 0.01495f $X=0.547 $Y=1.765 $X2=0 $Y2=0
cc_51 N_B_c_46_n N_A_35_368#_c_129_n 5.56095e-19 $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_52 N_B_c_41_n N_Y_c_162_n 0.0160525f $X=0.905 $Y=1.69 $X2=0 $Y2=0
cc_53 N_B_c_46_n N_Y_c_162_n 0.00132992f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_54 N_B_c_42_n N_Y_c_162_n 0.0209871f $X=0.455 $Y=1.385 $X2=0 $Y2=0
cc_55 N_B_c_43_n N_Y_c_162_n 0.01725f $X=0.547 $Y=1.22 $X2=0 $Y2=0
cc_56 N_B_c_48_n N_Y_c_162_n 0.00291398f $X=0.547 $Y=1.765 $X2=0 $Y2=0
cc_57 B N_Y_c_162_n 0.0278923f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_58 N_B_c_46_n Y 0.00230765f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_59 N_B_c_48_n Y 0.00281784f $X=0.547 $Y=1.765 $X2=0 $Y2=0
cc_60 N_B_c_46_n Y 0.0119971f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_61 N_B_c_48_n Y 0.0119915f $X=0.547 $Y=1.765 $X2=0 $Y2=0
cc_62 N_B_c_46_n N_VPWR_c_187_n 0.00333926f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_63 N_B_c_48_n N_VPWR_c_187_n 0.00333926f $X=0.547 $Y=1.765 $X2=0 $Y2=0
cc_64 N_B_c_46_n N_VPWR_c_185_n 0.00422798f $X=0.995 $Y=1.765 $X2=0 $Y2=0
cc_65 N_B_c_48_n N_VPWR_c_185_n 0.0042656f $X=0.547 $Y=1.765 $X2=0 $Y2=0
cc_66 N_B_c_42_n N_VGND_c_212_n 0.0022982f $X=0.455 $Y=1.385 $X2=0 $Y2=0
cc_67 N_B_c_43_n N_VGND_c_212_n 0.0161039f $X=0.547 $Y=1.22 $X2=0 $Y2=0
cc_68 B N_VGND_c_212_n 0.0283463f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_69 N_B_c_43_n N_VGND_c_214_n 0.00434272f $X=0.547 $Y=1.22 $X2=0 $Y2=0
cc_70 N_B_c_43_n N_VGND_c_216_n 0.00824032f $X=0.547 $Y=1.22 $X2=0 $Y2=0
cc_71 N_A_M1004_g N_A_35_368#_c_126_n 0.00101073f $X=1.445 $Y=2.4 $X2=0 $Y2=0
cc_72 N_A_c_80_n N_A_35_368#_c_128_n 8.34335e-19 $X=1.355 $Y=1.26 $X2=0 $Y2=0
cc_73 N_A_M1004_g N_A_35_368#_c_128_n 0.0185489f $X=1.445 $Y=2.4 $X2=0 $Y2=0
cc_74 N_A_M1005_g N_A_35_368#_c_128_n 0.0150781f $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_75 A N_A_35_368#_c_128_n 0.0350052f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_76 N_A_c_87_n N_A_35_368#_c_128_n 0.00458538f $X=1.97 $Y=1.44 $X2=0 $Y2=0
cc_77 N_A_c_80_n N_A_35_368#_c_129_n 0.00332308f $X=1.355 $Y=1.26 $X2=0 $Y2=0
cc_78 N_A_M1004_g N_A_35_368#_c_130_n 7.90488e-19 $X=1.445 $Y=2.4 $X2=0 $Y2=0
cc_79 N_A_M1005_g N_A_35_368#_c_130_n 0.0153871f $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_80 N_A_c_79_n N_Y_c_162_n 0.0126271f $X=0.995 $Y=1.185 $X2=0 $Y2=0
cc_81 N_A_c_81_n N_Y_c_162_n 0.00958281f $X=1.07 $Y=1.26 $X2=0 $Y2=0
cc_82 N_A_M1004_g N_Y_c_162_n 8.54645e-19 $X=1.445 $Y=2.4 $X2=0 $Y2=0
cc_83 N_A_c_87_n N_Y_c_162_n 0.0062569f $X=1.97 $Y=1.44 $X2=0 $Y2=0
cc_84 N_A_M1004_g N_VPWR_c_186_n 0.0150892f $X=1.445 $Y=2.4 $X2=0 $Y2=0
cc_85 N_A_M1005_g N_VPWR_c_186_n 0.00360149f $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_86 N_A_M1004_g N_VPWR_c_187_n 0.00460063f $X=1.445 $Y=2.4 $X2=0 $Y2=0
cc_87 N_A_M1005_g N_VPWR_c_189_n 0.005209f $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_88 N_A_M1004_g N_VPWR_c_185_n 0.00908665f $X=1.445 $Y=2.4 $X2=0 $Y2=0
cc_89 N_A_M1005_g N_VPWR_c_185_n 0.00986008f $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_90 N_A_c_79_n N_VGND_c_213_n 0.0184907f $X=0.995 $Y=1.185 $X2=0 $Y2=0
cc_91 N_A_c_80_n N_VGND_c_213_n 0.00955654f $X=1.355 $Y=1.26 $X2=0 $Y2=0
cc_92 A N_VGND_c_213_n 0.0211138f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_93 N_A_c_86_n N_VGND_c_213_n 0.0118488f $X=1.97 $Y=0.42 $X2=0 $Y2=0
cc_94 N_A_c_88_n N_VGND_c_213_n 0.0193455f $X=2.04 $Y=0.675 $X2=0 $Y2=0
cc_95 N_A_c_79_n N_VGND_c_214_n 0.00434272f $X=0.995 $Y=1.185 $X2=0 $Y2=0
cc_96 N_A_c_86_n N_VGND_c_215_n 0.00214182f $X=1.97 $Y=0.42 $X2=0 $Y2=0
cc_97 N_A_c_88_n N_VGND_c_215_n 0.0270748f $X=2.04 $Y=0.675 $X2=0 $Y2=0
cc_98 N_A_c_79_n N_VGND_c_216_n 0.00825157f $X=0.995 $Y=1.185 $X2=0 $Y2=0
cc_99 N_A_c_88_n N_VGND_c_216_n 0.0175158f $X=2.04 $Y=0.675 $X2=0 $Y2=0
cc_100 N_A_35_368#_c_126_n N_Y_M1002_d 0.00165831f $X=1.135 $Y=2.99 $X2=0 $Y2=0
cc_101 N_A_35_368#_c_129_n N_Y_c_162_n 0.00860227f $X=1.305 $Y=1.86 $X2=0 $Y2=0
cc_102 N_A_35_368#_c_125_n Y 0.030926f $X=0.32 $Y=1.985 $X2=0 $Y2=0
cc_103 N_A_35_368#_c_126_n Y 0.0166444f $X=1.135 $Y=2.99 $X2=0 $Y2=0
cc_104 N_A_35_368#_c_128_n N_VPWR_M1004_d 0.00165831f $X=1.955 $Y=1.86 $X2=-0.19
+ $Y2=1.66
cc_105 N_A_35_368#_c_126_n N_VPWR_c_186_n 0.010126f $X=1.135 $Y=2.99 $X2=0 $Y2=0
cc_106 N_A_35_368#_c_128_n N_VPWR_c_186_n 0.0148589f $X=1.955 $Y=1.86 $X2=0
+ $Y2=0
cc_107 N_A_35_368#_c_130_n N_VPWR_c_186_n 0.0291737f $X=2.12 $Y=1.985 $X2=0
+ $Y2=0
cc_108 N_A_35_368#_c_126_n N_VPWR_c_187_n 0.0581059f $X=1.135 $Y=2.99 $X2=0
+ $Y2=0
cc_109 N_A_35_368#_c_127_n N_VPWR_c_187_n 0.0179217f $X=0.405 $Y=2.99 $X2=0
+ $Y2=0
cc_110 N_A_35_368#_c_130_n N_VPWR_c_189_n 0.014549f $X=2.12 $Y=1.985 $X2=0 $Y2=0
cc_111 N_A_35_368#_c_126_n N_VPWR_c_185_n 0.0324093f $X=1.135 $Y=2.99 $X2=0
+ $Y2=0
cc_112 N_A_35_368#_c_127_n N_VPWR_c_185_n 0.00971942f $X=0.405 $Y=2.99 $X2=0
+ $Y2=0
cc_113 N_A_35_368#_c_130_n N_VPWR_c_185_n 0.0119743f $X=2.12 $Y=1.985 $X2=0
+ $Y2=0
cc_114 N_A_35_368#_c_128_n N_VGND_c_213_n 0.00422276f $X=1.955 $Y=1.86 $X2=0
+ $Y2=0
cc_115 N_A_35_368#_c_129_n N_VGND_c_213_n 0.00618439f $X=1.305 $Y=1.86 $X2=0
+ $Y2=0
cc_116 N_Y_c_162_n N_VGND_c_212_n 0.0255553f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_117 N_Y_c_162_n N_VGND_c_213_n 0.0308485f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_118 N_Y_c_162_n N_VGND_c_214_n 0.0144922f $X=0.78 $Y=0.515 $X2=0 $Y2=0
cc_119 N_Y_c_162_n N_VGND_c_216_n 0.0118826f $X=0.78 $Y=0.515 $X2=0 $Y2=0

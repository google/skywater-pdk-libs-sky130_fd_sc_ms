* File: sky130_fd_sc_ms__o211a_1.pex.spice
* Created: Fri Aug 28 17:52:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O211A_1%A_83_264# 1 2 3 12 16 19 22 23 24 25 28 31
+ 32 33 34 36 38 41 42 44 46
c110 44 0 1.43802e-19 $X=2.56 $Y=2.105
c111 23 0 1.605e-19 $X=1.01 $Y=1.97
r112 46 47 13.5953 $w=3.41e-07 $l=3.8e-07 $layer=LI1_cond $X=3.947 $Y=0.855
+ $X2=3.947 $Y2=1.235
r113 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.93
+ $Y=1.485 $X2=0.93 $Y2=1.485
r114 36 49 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=2.14 $X2=4.04
+ $Y2=2.055
r115 36 38 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.04 $Y=2.14
+ $X2=4.04 $Y2=2.815
r116 35 44 4.30018 $w=1.7e-07 $l=2.27376e-07 $layer=LI1_cond $X=2.835 $Y=2.055
+ $X2=2.615 $Y2=2.04
r117 34 49 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=2.055
+ $X2=4.04 $Y2=2.055
r118 34 35 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=3.875 $Y=2.055
+ $X2=2.835 $Y2=2.055
r119 32 47 4.81864 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=3.76 $Y=1.235
+ $X2=3.947 $Y2=1.235
r120 32 33 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=3.76 $Y=1.235
+ $X2=2.835 $Y2=1.235
r121 31 44 1.96316 $w=1.7e-07 $l=1.78115e-07 $layer=LI1_cond $X=2.75 $Y=1.94
+ $X2=2.615 $Y2=2.04
r122 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.75 $Y=1.32
+ $X2=2.835 $Y2=1.235
r123 30 31 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.75 $Y=1.32
+ $X2=2.75 $Y2=1.94
r124 26 44 1.96316 $w=3.3e-07 $l=1.24499e-07 $layer=LI1_cond $X=2.56 $Y=2.14
+ $X2=2.615 $Y2=2.04
r125 26 28 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.56 $Y=2.14
+ $X2=2.56 $Y2=2.815
r126 24 44 4.30018 $w=1.7e-07 $l=2.27376e-07 $layer=LI1_cond $X=2.395 $Y=2.055
+ $X2=2.615 $Y2=2.04
r127 24 25 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=2.395 $Y=2.055
+ $X2=1.095 $Y2=2.055
r128 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.01 $Y=1.97
+ $X2=1.095 $Y2=2.055
r129 22 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.01 $Y=1.65
+ $X2=1.01 $Y2=1.485
r130 22 23 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.01 $Y=1.65
+ $X2=1.01 $Y2=1.97
r131 18 42 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=0.595 $Y=1.485
+ $X2=0.93 $Y2=1.485
r132 18 19 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.595 $Y=1.485
+ $X2=0.505 $Y2=1.485
r133 14 19 34.7346 $w=1.65e-07 $l=1.69926e-07 $layer=POLY_cond $X=0.495 $Y=1.32
+ $X2=0.505 $Y2=1.485
r134 14 16 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.495 $Y=1.32
+ $X2=0.495 $Y2=0.74
r135 10 19 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.65
+ $X2=0.505 $Y2=1.485
r136 10 12 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=0.505 $Y=1.65
+ $X2=0.505 $Y2=2.4
r137 3 49 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=1.96 $X2=4.04 $Y2=2.135
r138 3 38 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=1.96 $X2=4.04 $Y2=2.815
r139 2 44 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.425
+ $Y=1.96 $X2=2.56 $Y2=2.105
r140 2 28 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.425
+ $Y=1.96 $X2=2.56 $Y2=2.815
r141 1 46 91 $w=1.7e-07 $l=2.5807e-07 $layer=licon1_NDIFF $count=2 $X=3.785
+ $Y=0.68 $X2=3.97 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_1%A1 3 7 9 15 16
c38 7 0 1.43802e-19 $X=1.915 $Y=2.46
r39 14 16 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.635
+ $X2=1.915 $Y2=1.635
r40 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.84
+ $Y=1.635 $X2=1.84 $Y2=1.635
r41 11 14 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.69 $Y=1.635
+ $X2=1.84 $Y2=1.635
r42 9 15 0.535558 $w=6.68e-07 $l=3e-08 $layer=LI1_cond $X=1.67 $Y=1.665 $X2=1.67
+ $Y2=1.635
r43 5 16 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.8
+ $X2=1.915 $Y2=1.635
r44 5 7 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.915 $Y=1.8 $X2=1.915
+ $Y2=2.46
r45 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.47
+ $X2=1.69 $Y2=1.635
r46 1 3 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.69 $Y=1.47 $X2=1.69
+ $Y2=1
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_1%A2 1 3 8 10 11 12 19
r38 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.49
+ $Y=0.405 $X2=2.49 $Y2=0.405
r39 16 19 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=2.35 $Y=0.405
+ $X2=2.49 $Y2=0.405
r40 11 12 14.3681 $w=3.83e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=0.447
+ $X2=3.6 $Y2=0.447
r41 10 11 14.3681 $w=3.83e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=0.447
+ $X2=3.12 $Y2=0.447
r42 10 20 4.49004 $w=3.83e-07 $l=1.5e-07 $layer=LI1_cond $X=2.64 $Y=0.447
+ $X2=2.49 $Y2=0.447
r43 8 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.35 $Y=1 $X2=2.35
+ $Y2=1.41
r44 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.35 $Y=0.57
+ $X2=2.35 $Y2=0.405
r45 5 8 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.35 $Y=0.57 $X2=2.35
+ $Y2=1
r46 1 9 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.335 $Y=1.5 $X2=2.335
+ $Y2=1.41
r47 1 3 373.161 $w=1.8e-07 $l=9.6e-07 $layer=POLY_cond $X=2.335 $Y=1.5 $X2=2.335
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_1%B1 3 7 9 16
r36 14 16 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=3.17 $Y=1.635
+ $X2=3.235 $Y2=1.635
r37 11 14 67.3216 $w=3.3e-07 $l=3.85e-07 $layer=POLY_cond $X=2.785 $Y=1.635
+ $X2=3.17 $Y2=1.635
r38 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.17
+ $Y=1.635 $X2=3.17 $Y2=1.635
r39 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.235 $Y=1.47
+ $X2=3.235 $Y2=1.635
r40 5 7 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=3.235 $Y=1.47 $X2=3.235
+ $Y2=1
r41 1 11 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.785 $Y=1.8
+ $X2=2.785 $Y2=1.635
r42 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.785 $Y=1.8 $X2=2.785
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_1%C1 3 7 9 12
r30 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.8 $Y=1.635
+ $X2=3.8 $Y2=1.8
r31 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.8 $Y=1.635
+ $X2=3.8 $Y2=1.47
r32 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.8
+ $Y=1.635 $X2=3.8 $Y2=1.635
r33 9 13 10.4092 $w=3.08e-07 $l=2.8e-07 $layer=LI1_cond $X=4.08 $Y=1.645 $X2=3.8
+ $Y2=1.645
r34 7 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.815 $Y=2.46
+ $X2=3.815 $Y2=1.8
r35 3 14 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=3.71 $Y=1 $X2=3.71
+ $Y2=1.47
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_1%X 1 2 9 13 14 15 16 23 32
r25 21 23 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=0.265 $Y=2 $X2=0.265
+ $Y2=2.035
r26 15 16 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.265 $Y=2.405
+ $X2=0.265 $Y2=2.775
r27 14 21 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.265 $Y=1.975
+ $X2=0.265 $Y2=2
r28 14 32 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=0.265 $Y=1.975
+ $X2=0.265 $Y2=1.82
r29 14 15 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=0.265 $Y=2.06
+ $X2=0.265 $Y2=2.405
r30 14 23 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.265 $Y=2.06
+ $X2=0.265 $Y2=2.035
r31 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.17 $Y=1.13 $X2=0.17
+ $Y2=1.82
r32 7 13 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.265 $Y=0.95
+ $X2=0.265 $Y2=1.13
r33 7 9 13.9254 $w=3.58e-07 $l=4.35e-07 $layer=LI1_cond $X=0.265 $Y=0.95
+ $X2=0.265 $Y2=0.515
r34 2 14 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r35 2 16 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r36 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_1%VPWR 1 2 9 11 18 25 26 31 39 41
r42 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r43 38 39 13.4207 $w=1.103e-06 $l=1.65e-07 $layer=LI1_cond $X=1.69 $Y=2.862
+ $X2=1.855 $Y2=2.862
r44 35 38 0.110407 $w=1.103e-06 $l=1e-08 $layer=LI1_cond $X=1.68 $Y=2.862
+ $X2=1.69 $Y2=2.862
r45 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 33 35 9.93665 $w=1.103e-06 $l=9e-07 $layer=LI1_cond $X=0.78 $Y=2.862
+ $X2=1.68 $Y2=2.862
r47 30 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 29 33 0.662443 $w=1.103e-06 $l=6e-08 $layer=LI1_cond $X=0.72 $Y=2.862
+ $X2=0.78 $Y2=2.862
r49 29 31 12.7583 $w=1.103e-06 $l=1.05e-07 $layer=LI1_cond $X=0.72 $Y=2.862
+ $X2=0.615 $Y2=2.862
r50 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 26 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r52 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r53 23 41 14.7259 $w=1.7e-07 $l=4.05e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=3.3 $Y2=3.33
r54 23 25 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=4.08 $Y2=3.33
r55 22 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r56 21 39 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=1.855 $Y2=3.33
r57 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r58 18 41 14.7259 $w=1.7e-07 $l=4.05e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=3.3 $Y2=3.33
r59 18 21 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=2.64 $Y2=3.33
r60 16 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 15 31 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=0.615 $Y2=3.33
r62 15 16 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r63 11 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r64 11 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 7 41 3.15573 $w=8.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=3.245 $X2=3.3
+ $Y2=3.33
r66 7 9 12.5514 $w=8.08e-07 $l=8.5e-07 $layer=LI1_cond $X=3.3 $Y=3.245 $X2=3.3
+ $Y2=2.395
r67 2 9 150 $w=1.7e-07 $l=8.55278e-07 $layer=licon1_PDIFF $count=4 $X=2.875
+ $Y=1.96 $X2=3.54 $Y2=2.395
r68 1 38 200 $w=1.7e-07 $l=1.34415e-06 $layer=licon1_PDIFF $count=3 $X=0.595
+ $Y=1.84 $X2=1.69 $Y2=2.395
r69 1 33 200 $w=1.7e-07 $l=6.40859e-07 $layer=licon1_PDIFF $count=3 $X=0.595
+ $Y=1.84 $X2=0.78 $Y2=2.395
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_1%VGND 1 2 9 13 16 17 18 20 33 34 37
r39 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r41 30 33 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r42 28 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r43 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r44 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r45 25 27 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.68
+ $Y2=0
r46 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r47 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r49 20 22 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r50 18 34 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r51 18 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r52 18 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r53 16 27 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=0 $X2=1.68
+ $Y2=0
r54 16 17 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.765 $Y=0 $X2=1.96
+ $Y2=0
r55 15 30 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.155 $Y=0 $X2=2.16
+ $Y2=0
r56 15 17 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.155 $Y=0 $X2=1.96
+ $Y2=0
r57 11 17 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0
r58 11 13 22.3101 $w=3.88e-07 $l=7.55e-07 $layer=LI1_cond $X=1.96 $Y=0.085
+ $X2=1.96 $Y2=0.84
r59 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0
r60 7 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.78 $Y=0.085 $X2=0.78
+ $Y2=0.515
r61 2 13 182 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_NDIFF $count=1 $X=1.765
+ $Y=0.68 $X2=1.96 $Y2=0.84
r62 1 9 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O211A_1%A_257_136# 1 2 9 11 12 14 15 17
r38 15 17 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.495 $Y=0.895
+ $X2=3.02 $Y2=0.895
r39 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.41 $Y=0.98
+ $X2=2.495 $Y2=0.895
r40 13 14 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.41 $Y=0.98 $X2=2.41
+ $Y2=1.13
r41 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.325 $Y=1.215
+ $X2=2.41 $Y2=1.13
r42 11 12 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.325 $Y=1.215
+ $X2=1.595 $Y2=1.215
r43 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.43 $Y=1.13
+ $X2=1.595 $Y2=1.215
r44 7 9 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.43 $Y=1.13 $X2=1.43
+ $Y2=0.825
r45 2 17 91 $w=1.7e-07 $l=6.94226e-07 $layer=licon1_NDIFF $count=2 $X=2.425
+ $Y=0.68 $X2=3.02 $Y2=0.895
r46 1 9 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=1.285
+ $Y=0.68 $X2=1.475 $Y2=0.825
.ends


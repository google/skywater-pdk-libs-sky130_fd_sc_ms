* File: sky130_fd_sc_ms__a21bo_4.pex.spice
* Created: Fri Aug 28 16:58:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A21BO_4%B1_N 3 8 11 13 19
c31 3 0 1.05294e-19 $X=0.495 $Y=2.46
r32 16 19 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.46 $Y=0.34
+ $X2=0.665 $Y2=0.34
r33 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.46
+ $Y=0.34 $X2=0.46 $Y2=0.34
r34 13 17 8.25846 $w=3.25e-07 $l=2.2e-07 $layer=LI1_cond $X=0.24 $Y=0.462
+ $X2=0.46 $Y2=0.462
r35 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.665 $Y=1.33
+ $X2=0.665 $Y2=1.405
r36 6 8 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.665 $Y=1.33
+ $X2=0.665 $Y2=0.935
r37 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.665 $Y=0.505
+ $X2=0.665 $Y2=0.34
r38 5 8 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.665 $Y=0.505
+ $X2=0.665 $Y2=0.935
r39 1 11 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.495 $Y=1.405
+ $X2=0.665 $Y2=1.405
r40 1 3 380.935 $w=1.8e-07 $l=9.8e-07 $layer=POLY_cond $X=0.495 $Y=1.48
+ $X2=0.495 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_4%A_184_338# 1 2 3 10 12 13 15 18 20 22 25 27
+ 29 32 34 36 37 44 45 49 53 55 56 59 61
c149 59 0 1.44963e-19 $X=4.95 $Y=0.76
c150 34 0 1.44963e-19 $X=2.545 $Y=1.35
c151 20 0 1.47805e-19 $X=1.685 $Y=1.35
r152 67 68 35.3563 $w=3.34e-07 $l=2.45e-07 $layer=POLY_cond $X=1.01 $Y=1.565
+ $X2=1.255 $Y2=1.565
r153 57 59 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=4.91 $Y=1.11
+ $X2=4.91 $Y2=0.76
r154 55 57 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.785 $Y=1.195
+ $X2=4.91 $Y2=1.11
r155 55 56 69.4813 $w=1.68e-07 $l=1.065e-06 $layer=LI1_cond $X=4.785 $Y=1.195
+ $X2=3.72 $Y2=1.195
r156 51 56 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.595 $Y=1.195
+ $X2=3.72 $Y2=1.195
r157 51 53 38.4916 $w=2.48e-07 $l=8.35e-07 $layer=LI1_cond $X=3.595 $Y=1.28
+ $X2=3.595 $Y2=2.115
r158 47 51 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.25 $Y=1.195
+ $X2=3.595 $Y2=1.195
r159 47 49 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=3.25 $Y=1.11
+ $X2=3.25 $Y2=0.76
r160 46 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=1.195
+ $X2=2.67 $Y2=1.195
r161 45 47 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=1.195
+ $X2=3.25 $Y2=1.195
r162 45 46 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.085 $Y=1.195
+ $X2=2.755 $Y2=1.195
r163 44 76 15.8743 $w=3.34e-07 $l=1.1e-07 $layer=POLY_cond $X=2.435 $Y=1.565
+ $X2=2.545 $Y2=1.565
r164 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.435
+ $Y=1.515 $X2=2.435 $Y2=1.515
r165 40 70 10.1018 $w=3.34e-07 $l=7e-08 $layer=POLY_cond $X=1.755 $Y=1.565
+ $X2=1.685 $Y2=1.565
r166 39 43 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.755 $Y=1.515
+ $X2=2.435 $Y2=1.515
r167 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.755
+ $Y=1.515 $X2=1.755 $Y2=1.515
r168 37 61 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.67 $Y=1.515
+ $X2=2.67 $Y2=1.195
r169 37 43 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.585 $Y=1.515
+ $X2=2.435 $Y2=1.515
r170 34 76 21.5099 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=2.545 $Y=1.35
+ $X2=2.545 $Y2=1.565
r171 34 36 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.545 $Y=1.35
+ $X2=2.545 $Y2=0.87
r172 30 44 10.8234 $w=3.34e-07 $l=7.5e-08 $layer=POLY_cond $X=2.36 $Y=1.565
+ $X2=2.435 $Y2=1.565
r173 30 73 35.3563 $w=3.34e-07 $l=2.45e-07 $layer=POLY_cond $X=2.36 $Y=1.565
+ $X2=2.115 $Y2=1.565
r174 30 32 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.36 $Y=1.68
+ $X2=2.36 $Y2=2.4
r175 27 73 21.5099 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=2.115 $Y=1.35
+ $X2=2.115 $Y2=1.565
r176 27 29 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.115 $Y=1.35
+ $X2=2.115 $Y2=0.87
r177 23 73 29.5838 $w=3.34e-07 $l=2.05e-07 $layer=POLY_cond $X=1.91 $Y=1.565
+ $X2=2.115 $Y2=1.565
r178 23 40 22.3683 $w=3.34e-07 $l=1.55e-07 $layer=POLY_cond $X=1.91 $Y=1.565
+ $X2=1.755 $Y2=1.565
r179 23 25 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.91 $Y=1.68
+ $X2=1.91 $Y2=2.4
r180 20 70 21.5099 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.685 $Y=1.35
+ $X2=1.685 $Y2=1.565
r181 20 22 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.685 $Y=1.35
+ $X2=1.685 $Y2=0.87
r182 16 70 32.4701 $w=3.34e-07 $l=2.25e-07 $layer=POLY_cond $X=1.46 $Y=1.565
+ $X2=1.685 $Y2=1.565
r183 16 68 29.5838 $w=3.34e-07 $l=2.05e-07 $layer=POLY_cond $X=1.46 $Y=1.565
+ $X2=1.255 $Y2=1.565
r184 16 18 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.46 $Y=1.68
+ $X2=1.46 $Y2=2.4
r185 13 68 21.5099 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.255 $Y=1.35
+ $X2=1.255 $Y2=1.565
r186 13 15 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.255 $Y=1.35
+ $X2=1.255 $Y2=0.87
r187 10 67 17.2128 $w=1.8e-07 $l=2.15e-07 $layer=POLY_cond $X=1.01 $Y=1.78
+ $X2=1.01 $Y2=1.565
r188 10 12 166.022 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=1.01 $Y=1.78
+ $X2=1.01 $Y2=2.4
r189 3 53 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=3.42
+ $Y=1.96 $X2=3.555 $Y2=2.115
r190 2 59 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.81
+ $Y=0.615 $X2=4.95 $Y2=0.76
r191 1 49 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.11
+ $Y=0.615 $X2=3.25 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_4%A_29_392# 1 2 9 13 15 17 21 26 29 31 34 35
+ 36 39 45 47
c106 21 0 3.47333e-19 $X=3.78 $Y=2.46
r107 42 45 4.76873 $w=4.33e-07 $l=1.8e-07 $layer=LI1_cond $X=0.27 $Y=1.057
+ $X2=0.45 $Y2=1.057
r108 40 50 41.1708 $w=2.4e-07 $l=2.05e-07 $layer=POLY_cond $X=3.125 $Y=1.615
+ $X2=3.33 $Y2=1.615
r109 40 48 18.075 $w=2.4e-07 $l=9e-08 $layer=POLY_cond $X=3.125 $Y=1.615
+ $X2=3.035 $Y2=1.615
r110 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.125
+ $Y=1.615 $X2=3.125 $Y2=1.615
r111 37 39 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=3.125 $Y=1.85
+ $X2=3.125 $Y2=1.615
r112 35 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.96 $Y=1.935
+ $X2=3.125 $Y2=1.85
r113 35 36 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.96 $Y=1.935
+ $X2=2.64 $Y2=1.935
r114 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.555 $Y=2.02
+ $X2=2.64 $Y2=1.935
r115 33 34 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.555 $Y=2.02
+ $X2=2.555 $Y2=2.27
r116 32 47 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.435 $Y=2.355
+ $X2=0.27 $Y2=2.355
r117 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.47 $Y=2.355
+ $X2=2.555 $Y2=2.27
r118 31 32 132.765 $w=1.68e-07 $l=2.035e-06 $layer=LI1_cond $X=2.47 $Y=2.355
+ $X2=0.435 $Y2=2.355
r119 27 47 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=2.44
+ $X2=0.27 $Y2=2.355
r120 27 29 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=0.27 $Y=2.44
+ $X2=0.27 $Y2=2.815
r121 24 47 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=2.27
+ $X2=0.27 $Y2=2.355
r122 24 26 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.27 $Y=2.27
+ $X2=0.27 $Y2=2.105
r123 23 42 2.35727 $w=3.3e-07 $l=2.18e-07 $layer=LI1_cond $X=0.27 $Y=1.275
+ $X2=0.27 $Y2=1.057
r124 23 26 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.27 $Y=1.275
+ $X2=0.27 $Y2=2.105
r125 19 21 334.29 $w=1.8e-07 $l=8.6e-07 $layer=POLY_cond $X=3.78 $Y=1.6 $X2=3.78
+ $Y2=2.46
r126 15 19 63.2625 $w=2.4e-07 $l=3.82721e-07 $layer=POLY_cond $X=3.465 $Y=1.45
+ $X2=3.78 $Y2=1.6
r127 15 50 27.1125 $w=2.4e-07 $l=2.22486e-07 $layer=POLY_cond $X=3.465 $Y=1.45
+ $X2=3.33 $Y2=1.615
r128 15 17 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=3.465 $Y=1.45
+ $X2=3.465 $Y2=0.935
r129 11 50 9.57678 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.33 $Y=1.78
+ $X2=3.33 $Y2=1.615
r130 11 13 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=3.33 $Y=1.78
+ $X2=3.33 $Y2=2.46
r131 7 48 13.7767 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.035 $Y=1.45
+ $X2=3.035 $Y2=1.615
r132 7 9 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=3.035 $Y=1.45
+ $X2=3.035 $Y2=0.935
r133 2 29 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.96 $X2=0.27 $Y2=2.815
r134 2 26 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.96 $X2=0.27 $Y2=2.105
r135 1 45 182 $w=1.7e-07 $l=4.98598e-07 $layer=licon1_NDIFF $count=1 $X=0.325
+ $Y=0.615 $X2=0.45 $Y2=1.055
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_4%A1 3 7 11 15 17 18 26
c44 15 0 1.44963e-19 $X=5.165 $Y=0.935
r45 26 27 5.20679 $w=3.24e-07 $l=3.5e-08 $layer=POLY_cond $X=5.13 $Y=1.615
+ $X2=5.165 $Y2=1.615
r46 24 26 55.787 $w=3.24e-07 $l=3.75e-07 $layer=POLY_cond $X=4.755 $Y=1.615
+ $X2=5.13 $Y2=1.615
r47 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.755
+ $Y=1.615 $X2=4.755 $Y2=1.615
r48 22 24 2.97531 $w=3.24e-07 $l=2e-08 $layer=POLY_cond $X=4.735 $Y=1.615
+ $X2=4.755 $Y2=1.615
r49 21 22 8.1821 $w=3.24e-07 $l=5.5e-08 $layer=POLY_cond $X=4.68 $Y=1.615
+ $X2=4.735 $Y2=1.615
r50 18 25 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=5.04 $Y=1.615
+ $X2=4.755 $Y2=1.615
r51 17 25 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=4.56 $Y=1.615
+ $X2=4.755 $Y2=1.615
r52 13 27 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.165 $Y=1.45
+ $X2=5.165 $Y2=1.615
r53 13 15 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=5.165 $Y=1.45
+ $X2=5.165 $Y2=0.935
r54 9 26 16.5046 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.13 $Y=1.78
+ $X2=5.13 $Y2=1.615
r55 9 11 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=5.13 $Y=1.78 $X2=5.13
+ $Y2=2.46
r56 5 22 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.735 $Y=1.45
+ $X2=4.735 $Y2=1.615
r57 5 7 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=4.735 $Y=1.45
+ $X2=4.735 $Y2=0.935
r58 1 21 16.5046 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.68 $Y=1.78
+ $X2=4.68 $Y2=1.615
r59 1 3 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=4.68 $Y=1.78 $X2=4.68
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_4%A2 1 3 8 9 11 13 18 21 23 27
r66 26 28 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=4.127 $Y=0.34
+ $X2=4.127 $Y2=0.505
r67 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.1
+ $Y=0.34 $X2=4.1 $Y2=0.34
r68 23 26 20.2238 $w=3.85e-07 $l=1.4e-07 $layer=POLY_cond $X=4.127 $Y=0.2
+ $X2=4.127 $Y2=0.34
r69 21 27 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=4.1 $Y=0.555
+ $X2=4.1 $Y2=0.34
r70 18 20 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.595 $Y=0.935
+ $X2=5.595 $Y2=1.33
r71 15 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.595 $Y=0.275
+ $X2=5.595 $Y2=0.935
r72 11 20 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.58 $Y=1.42 $X2=5.58
+ $Y2=1.33
r73 11 13 404.258 $w=1.8e-07 $l=1.04e-06 $layer=POLY_cond $X=5.58 $Y=1.42
+ $X2=5.58 $Y2=2.46
r74 10 23 24.9301 $w=1.5e-07 $l=1.93e-07 $layer=POLY_cond $X=4.32 $Y=0.2
+ $X2=4.127 $Y2=0.2
r75 9 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.52 $Y=0.2
+ $X2=5.595 $Y2=0.275
r76 9 10 615.319 $w=1.5e-07 $l=1.2e-06 $layer=POLY_cond $X=5.52 $Y=0.2 $X2=4.32
+ $Y2=0.2
r77 8 19 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=4.245 $Y=0.935
+ $X2=4.245 $Y2=1.33
r78 8 28 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.245 $Y=0.935
+ $X2=4.245 $Y2=0.505
r79 1 19 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.23 $Y=1.42 $X2=4.23
+ $Y2=1.33
r80 1 3 404.258 $w=1.8e-07 $l=1.04e-06 $layer=POLY_cond $X=4.23 $Y=1.42 $X2=4.23
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_4%VPWR 1 2 3 4 5 18 22 26 30 34 37 38 40 41 42
+ 44 49 54 70 71 74 77 80
c87 30 0 1.87992e-19 $X=4.455 $Y=2.455
r88 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r89 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r90 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r91 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r92 68 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r93 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r94 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r95 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r96 61 64 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=3.33 $X2=4.08
+ $Y2=3.33
r97 59 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=3.33
+ $X2=2.585 $Y2=3.33
r98 59 61 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.75 $Y=3.33 $X2=3.12
+ $Y2=3.33
r99 58 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r100 58 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r101 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r102 55 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.85 $Y=3.33
+ $X2=1.685 $Y2=3.33
r103 55 57 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.85 $Y=3.33
+ $X2=2.16 $Y2=3.33
r104 54 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.42 $Y=3.33
+ $X2=2.585 $Y2=3.33
r105 54 57 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.42 $Y=3.33
+ $X2=2.16 $Y2=3.33
r106 53 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r107 53 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r108 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r109 50 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=3.33
+ $X2=0.785 $Y2=3.33
r110 50 52 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.95 $Y=3.33
+ $X2=1.2 $Y2=3.33
r111 49 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=3.33
+ $X2=1.685 $Y2=3.33
r112 49 52 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.52 $Y=3.33 $X2=1.2
+ $Y2=3.33
r113 47 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r114 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r115 44 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=3.33
+ $X2=0.785 $Y2=3.33
r116 44 46 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.62 $Y=3.33
+ $X2=0.24 $Y2=3.33
r117 42 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r118 42 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r119 42 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r120 40 67 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.27 $Y=3.33
+ $X2=5.04 $Y2=3.33
r121 40 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.27 $Y=3.33
+ $X2=5.395 $Y2=3.33
r122 39 70 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r123 39 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=5.395 $Y2=3.33
r124 37 64 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.29 $Y=3.33
+ $X2=4.08 $Y2=3.33
r125 37 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.29 $Y=3.33
+ $X2=4.415 $Y2=3.33
r126 36 67 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=4.54 $Y=3.33 $X2=5.04
+ $Y2=3.33
r127 36 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.54 $Y=3.33
+ $X2=4.415 $Y2=3.33
r128 32 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=3.245
+ $X2=5.395 $Y2=3.33
r129 32 34 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=5.395 $Y=3.245
+ $X2=5.395 $Y2=2.455
r130 28 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.415 $Y=3.245
+ $X2=4.415 $Y2=3.33
r131 28 30 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=4.415 $Y=3.245
+ $X2=4.415 $Y2=2.455
r132 24 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=3.245
+ $X2=2.585 $Y2=3.33
r133 24 26 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=2.585 $Y=3.245
+ $X2=2.585 $Y2=2.775
r134 20 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.685 $Y=3.245
+ $X2=1.685 $Y2=3.33
r135 20 22 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=1.685 $Y=3.245
+ $X2=1.685 $Y2=2.775
r136 16 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=3.245
+ $X2=0.785 $Y2=3.33
r137 16 18 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.785 $Y=3.245
+ $X2=0.785 $Y2=2.775
r138 5 34 300 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=2 $X=5.22
+ $Y=1.96 $X2=5.355 $Y2=2.455
r139 4 30 300 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=2 $X=4.32
+ $Y=1.96 $X2=4.455 $Y2=2.455
r140 3 26 600 $w=1.7e-07 $l=1.00022e-06 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.84 $X2=2.585 $Y2=2.775
r141 2 22 600 $w=1.7e-07 $l=1.00022e-06 $layer=licon1_PDIFF $count=1 $X=1.55
+ $Y=1.84 $X2=1.685 $Y2=2.775
r142 1 18 600 $w=1.7e-07 $l=9.09519e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.96 $X2=0.785 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_4%X 1 2 3 4 15 18 21 23 27 29 30 31 32
c54 27 0 1.44963e-19 $X=2.33 $Y=0.645
c55 18 0 1.05294e-19 $X=1.335 $Y=1.51
c56 15 0 1.47805e-19 $X=1.47 $Y=0.645
r57 32 38 10.4403 $w=5.88e-07 $l=5.15e-07 $layer=LI1_cond $X=0.72 $Y=1.805
+ $X2=1.235 $Y2=1.805
r58 30 38 0.304088 $w=5.88e-07 $l=1.5e-08 $layer=LI1_cond $X=1.25 $Y=1.805
+ $X2=1.235 $Y2=1.805
r59 30 31 2.31106 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=1.805
+ $X2=1.335 $Y2=1.805
r60 25 27 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=2.29 $Y=1.01
+ $X2=2.29 $Y2=0.645
r61 24 29 2.57001 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.555 $Y=1.095
+ $X2=1.402 $Y2=1.095
r62 23 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.165 $Y=1.095
+ $X2=2.29 $Y2=1.01
r63 23 24 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.165 $Y=1.095
+ $X2=1.555 $Y2=1.095
r64 19 31 2.31106 $w=4.2e-07 $l=2.08207e-07 $layer=LI1_cond $X=1.42 $Y=1.975
+ $X2=1.335 $Y2=1.805
r65 19 21 32.9599 $w=2.48e-07 $l=7.15e-07 $layer=LI1_cond $X=1.42 $Y=1.975
+ $X2=2.135 $Y2=1.975
r66 18 31 4.73016 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=1.335 $Y=1.51
+ $X2=1.335 $Y2=1.805
r67 17 29 3.87901 $w=2.37e-07 $l=1.13666e-07 $layer=LI1_cond $X=1.335 $Y=1.18
+ $X2=1.402 $Y2=1.095
r68 17 18 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.335 $Y=1.18
+ $X2=1.335 $Y2=1.51
r69 13 29 3.87901 $w=2.37e-07 $l=8.5e-08 $layer=LI1_cond $X=1.402 $Y=1.01
+ $X2=1.402 $Y2=1.095
r70 13 15 13.7915 $w=3.03e-07 $l=3.65e-07 $layer=LI1_cond $X=1.402 $Y=1.01
+ $X2=1.402 $Y2=0.645
r71 4 21 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2 $Y=1.84
+ $X2=2.135 $Y2=2.015
r72 3 38 600 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=1 $X=1.1
+ $Y=1.84 $X2=1.235 $Y2=2
r73 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.19
+ $Y=0.5 $X2=2.33 $Y2=0.645
r74 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.33
+ $Y=0.5 $X2=1.47 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_4%A_596_392# 1 2 3 4 15 17 18 19 23 27 29 31
+ 33 38
c66 19 0 1.59341e-19 $X=4.005 $Y=2.12
r67 31 40 2.9222 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=5.845 $Y=2.12 $X2=5.845
+ $Y2=2.03
r68 31 33 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=5.845 $Y=2.12
+ $X2=5.845 $Y2=2.815
r69 30 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.07 $Y=2.035
+ $X2=4.905 $Y2=2.035
r70 29 40 4.22096 $w=1.7e-07 $l=1.27475e-07 $layer=LI1_cond $X=5.72 $Y=2.035
+ $X2=5.845 $Y2=2.03
r71 29 30 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.72 $Y=2.035
+ $X2=5.07 $Y2=2.035
r72 25 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.905 $Y=2.12
+ $X2=4.905 $Y2=2.035
r73 25 27 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.905 $Y=2.12
+ $X2=4.905 $Y2=2.815
r74 24 36 3.40825 $w=1.7e-07 $l=8.74643e-08 $layer=LI1_cond $X=4.09 $Y=2.035
+ $X2=4.005 $Y2=2.03
r75 23 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.74 $Y=2.035
+ $X2=4.905 $Y2=2.035
r76 23 24 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.74 $Y=2.035
+ $X2=4.09 $Y2=2.035
r77 20 22 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.005 $Y=2.905
+ $X2=4.005 $Y2=2.815
r78 19 36 3.40825 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=4.005 $Y=2.12 $X2=4.005
+ $Y2=2.03
r79 19 22 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.005 $Y=2.12
+ $X2=4.005 $Y2=2.815
r80 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.92 $Y=2.99
+ $X2=4.005 $Y2=2.905
r81 17 18 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.92 $Y=2.99
+ $X2=3.27 $Y2=2.99
r82 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.105 $Y=2.905
+ $X2=3.27 $Y2=2.99
r83 13 15 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=3.105 $Y=2.905
+ $X2=3.105 $Y2=2.355
r84 4 40 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.67
+ $Y=1.96 $X2=5.805 $Y2=2.105
r85 4 33 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=5.67
+ $Y=1.96 $X2=5.805 $Y2=2.815
r86 3 38 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=4.77
+ $Y=1.96 $X2=4.905 $Y2=2.115
r87 3 27 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.77
+ $Y=1.96 $X2=4.905 $Y2=2.815
r88 2 36 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.87
+ $Y=1.96 $X2=4.005 $Y2=2.105
r89 2 22 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.87
+ $Y=1.96 $X2=4.005 $Y2=2.815
r90 1 15 300 $w=1.7e-07 $l=4.53211e-07 $layer=licon1_PDIFF $count=2 $X=2.98
+ $Y=1.96 $X2=3.105 $Y2=2.355
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_4%VGND 1 2 3 4 5 18 24 26 30 32 36 38 40 43 44
+ 45 46 47 56 65 68 72
r87 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r88 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r89 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r90 63 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r91 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r92 60 63 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.52
+ $Y2=0
r93 60 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r94 59 62 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.52
+ $Y2=0
r95 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r96 57 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.765 $Y=0 $X2=3.68
+ $Y2=0
r97 57 59 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.765 $Y=0 $X2=4.08
+ $Y2=0
r98 56 71 3.87298 $w=1.7e-07 $l=2.57e-07 $layer=LI1_cond $X=5.725 $Y=0 $X2=5.982
+ $Y2=0
r99 56 62 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.725 $Y=0 $X2=5.52
+ $Y2=0
r100 55 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r101 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r102 51 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r103 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r104 47 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r105 47 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r106 45 54 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.735 $Y=0 $X2=1.68
+ $Y2=0
r107 45 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.735 $Y=0 $X2=1.86
+ $Y2=0
r108 43 50 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.72
+ $Y2=0
r109 43 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.92
+ $Y2=0
r110 42 54 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.045 $Y=0
+ $X2=1.68 $Y2=0
r111 42 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=0.92
+ $Y2=0
r112 38 71 3.27018 $w=2.5e-07 $l=1.69245e-07 $layer=LI1_cond $X=5.85 $Y=0.085
+ $X2=5.982 $Y2=0
r113 38 40 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.85 $Y=0.085
+ $X2=5.85 $Y2=0.76
r114 34 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.68 $Y=0.085
+ $X2=3.68 $Y2=0
r115 34 36 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.68 $Y=0.085
+ $X2=3.68 $Y2=0.775
r116 33 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.845 $Y=0 $X2=2.72
+ $Y2=0
r117 32 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=0 $X2=3.68
+ $Y2=0
r118 32 33 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=3.595 $Y=0
+ $X2=2.845 $Y2=0
r119 28 65 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.72 $Y=0.085
+ $X2=2.72 $Y2=0
r120 28 30 31.8074 $w=2.48e-07 $l=6.9e-07 $layer=LI1_cond $X=2.72 $Y=0.085
+ $X2=2.72 $Y2=0.775
r121 27 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.985 $Y=0 $X2=1.86
+ $Y2=0
r122 26 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.595 $Y=0 $X2=2.72
+ $Y2=0
r123 26 27 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.595 $Y=0
+ $X2=1.985 $Y2=0
r124 22 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.86 $Y=0.085
+ $X2=1.86 $Y2=0
r125 22 24 26.5062 $w=2.48e-07 $l=5.75e-07 $layer=LI1_cond $X=1.86 $Y=0.085
+ $X2=1.86 $Y2=0.66
r126 18 20 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=0.92 $Y=0.645
+ $X2=0.92 $Y2=1.11
r127 16 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.92 $Y=0.085
+ $X2=0.92 $Y2=0
r128 16 18 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=0.92 $Y=0.085
+ $X2=0.92 $Y2=0.645
r129 5 40 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.67
+ $Y=0.615 $X2=5.81 $Y2=0.76
r130 4 36 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=3.54
+ $Y=0.615 $X2=3.68 $Y2=0.775
r131 3 30 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.62
+ $Y=0.5 $X2=2.76 $Y2=0.775
r132 2 24 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=1.76
+ $Y=0.5 $X2=1.9 $Y2=0.66
r133 1 20 182 $w=1.7e-07 $l=5.94916e-07 $layer=licon1_NDIFF $count=1 $X=0.74
+ $Y=0.615 $X2=0.96 $Y2=1.11
r134 1 18 182 $w=1.7e-07 $l=2.34521e-07 $layer=licon1_NDIFF $count=1 $X=0.74
+ $Y=0.615 $X2=0.96 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__A21BO_4%A_864_123# 1 2 9 11 12 15
r32 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.38 $Y=0.425
+ $X2=5.38 $Y2=0.76
r33 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.215 $Y=0.34
+ $X2=5.38 $Y2=0.425
r34 11 12 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.215 $Y=0.34
+ $X2=4.605 $Y2=0.34
r35 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.52 $Y=0.425
+ $X2=4.605 $Y2=0.34
r36 7 9 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.52 $Y=0.425 $X2=4.52
+ $Y2=0.765
r37 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.24
+ $Y=0.615 $X2=5.38 $Y2=0.76
r38 1 9 182 $w=1.7e-07 $l=2.64575e-07 $layer=licon1_NDIFF $count=1 $X=4.32
+ $Y=0.615 $X2=4.52 $Y2=0.765
.ends


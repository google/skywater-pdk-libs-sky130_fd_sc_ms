* File: sky130_fd_sc_ms__sedfxtp_1.spice
* Created: Fri Aug 28 18:16:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sedfxtp_1.pex.spice"
.subckt sky130_fd_sc_ms__sedfxtp_1  VNB VPB D DE SCD SCE CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCE	SCE
* SCD	SCD
* DE	DE
* D	D
* VPB	VPB
* VNB	VNB
MM1010 A_143_74# N_D_M1010_g N_A_27_74#_M1010_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1806 PD=0.66 PS=1.7 NRD=18.564 NRS=21.42 M=1 R=2.8 SA=75000.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_DE_M1002_g A_143_74# VNB NLOWVT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.7 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_DE_M1007_g N_A_159_404#_M1007_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1008 A_505_111# N_A_159_404#_M1008_g N_VGND_M1007_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1039 N_A_27_74#_M1039_d N_A_547_301#_M1039_g A_505_111# VNB NLOWVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1022 N_A_669_111#_M1022_d N_A_639_85#_M1022_g N_A_27_74#_M1039_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1491 AS=0.0588 PD=1.55 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1040 N_VGND_M1040_d N_SCE_M1040_g N_A_639_85#_M1040_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1176 PD=0.7 PS=1.4 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1031 A_1026_125# N_SCD_M1031_g N_VGND_M1040_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1028 N_A_669_111#_M1028_d N_SCE_M1028_g A_1026_125# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1176 AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_A_1295_74#_M1011_d N_CLK_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2072 AS=0.2109 PD=2.04 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1004 N_A_1492_74#_M1004_d N_A_1295_74#_M1004_g N_VGND_M1004_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2072 AS=0.2109 PD=2.04 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1023 N_A_1688_97#_M1023_d N_A_1295_74#_M1023_g N_A_669_111#_M1023_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1176 PD=0.95 PS=1.4 NRD=71.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1032 A_1824_97# N_A_1492_74#_M1032_g N_A_1688_97#_M1023_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0903 AS=0.1113 PD=0.85 PS=0.95 NRD=45.708 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_A_1910_71#_M1029_g A_1824_97# VNB NLOWVT L=0.15 W=0.42
+ AD=0.135232 AS=0.0903 PD=0.986604 PS=0.85 NRD=22.848 NRS=45.708 M=1 R=2.8
+ SA=75001.5 SB=75001 A=0.063 P=1.14 MULT=1
MM1033 N_A_1910_71#_M1033_d N_A_1688_97#_M1033_g N_VGND_M1029_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.206068 PD=1.85 PS=1.5034 NRD=0 NRS=46.872 M=1
+ R=4.26667 SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1016 A_2313_74# N_A_1910_71#_M1016_g N_VGND_M1016_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1824 PD=0.85 PS=1.85 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1018 N_A_2385_74#_M1018_d N_A_1492_74#_M1018_g A_2313_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.129147 AS=0.0672 PD=1.20755 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667
+ SA=75000.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1035 A_2487_74# N_A_1295_74#_M1035_g N_A_2385_74#_M1018_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0847528 PD=0.66 PS=0.792453 NRD=18.564 NRS=23.568 M=1
+ R=2.8 SA=75001.1 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1036 N_VGND_M1036_d N_A_547_301#_M1036_g A_2487_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.20475 AS=0.0504 PD=1.395 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.5
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1013 N_A_547_301#_M1013_d N_A_2385_74#_M1013_g N_VGND_M1036_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1197 AS=0.20475 PD=1.41 PS=1.395 NRD=0 NRS=19.992 M=1 R=2.8
+ SA=75002.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_2385_74#_M1003_g N_Q_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1024 A_117_464# N_D_M1024_g N_A_27_74#_M1024_s VPB PSHORT L=0.18 W=0.64
+ AD=0.0672 AS=0.1728 PD=0.85 PS=1.82 NRD=15.3857 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1038 N_VPWR_M1038_d N_A_159_404#_M1038_g A_117_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.1792 AS=0.0672 PD=1.84 PS=0.85 NRD=0 NRS=15.3857 M=1 R=3.55556 SA=90000.6
+ SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1021 N_VPWR_M1021_d N_DE_M1021_g N_A_159_404#_M1021_s VPB PSHORT L=0.18 W=0.64
+ AD=0.16 AS=0.1792 PD=1.14 PS=1.84 NRD=69.2455 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90001.7 A=0.1152 P=1.64 MULT=1
MM1001 A_557_463# N_DE_M1001_g N_VPWR_M1021_d VPB PSHORT L=0.18 W=0.64 AD=0.0672
+ AS=0.16 PD=0.85 PS=1.14 NRD=15.3857 NRS=0 M=1 R=3.55556 SA=90000.9 SB=90001
+ A=0.1152 P=1.64 MULT=1
MM1015 N_A_27_74#_M1015_d N_A_547_301#_M1015_g A_557_463# VPB PSHORT L=0.18
+ W=0.64 AD=0.0864 AS=0.0672 PD=0.91 PS=0.85 NRD=0 NRS=15.3857 M=1 R=3.55556
+ SA=90001.3 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1019 N_A_669_111#_M1019_d N_SCE_M1019_g N_A_27_74#_M1015_d VPB PSHORT L=0.18
+ W=0.64 AD=0.1664 AS=0.0864 PD=1.8 PS=0.91 NRD=0 NRS=0 M=1 R=3.55556 SA=90001.7
+ SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1014 N_VPWR_M1014_d N_SCE_M1014_g N_A_639_85#_M1014_s VPB PSHORT L=0.18 W=0.64
+ AD=0.16 AS=0.1696 PD=1.14 PS=1.81 NRD=69.2455 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90001.2 A=0.1152 P=1.64 MULT=1
MM1005 A_1056_455# N_SCD_M1005_g N_VPWR_M1014_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0672 AS=0.16 PD=0.85 PS=1.14 NRD=15.3857 NRS=0 M=1 R=3.55556 SA=90000.9
+ SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1020 N_A_669_111#_M1020_d N_A_639_85#_M1020_g A_1056_455# VPB PSHORT L=0.18
+ W=0.64 AD=0.1664 AS=0.0672 PD=1.8 PS=0.85 NRD=0 NRS=15.3857 M=1 R=3.55556
+ SA=90001.2 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1006 N_A_1295_74#_M1006_d N_CLK_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18
+ W=1.12 AD=0.2912 AS=0.2912 PD=2.76 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1017 N_A_1492_74#_M1017_d N_A_1295_74#_M1017_g N_VPWR_M1017_s VPB PSHORT
+ L=0.18 W=1.12 AD=0.2912 AS=0.2912 PD=2.76 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1026 N_A_1688_97#_M1026_d N_A_1492_74#_M1026_g N_A_669_111#_M1026_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0672 AS=0.1113 PD=0.74 PS=1.37 NRD=21.0987 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90001.5 A=0.0756 P=1.2 MULT=1
MM1027 A_1893_508# N_A_1295_74#_M1027_g N_A_1688_97#_M1026_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0525 AS=0.0672 PD=0.67 PS=0.74 NRD=32.8202 NRS=0 M=1 R=2.33333
+ SA=90000.7 SB=90001 A=0.0756 P=1.2 MULT=1
MM1030 N_VPWR_M1030_d N_A_1910_71#_M1030_g A_1893_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.0901833 AS=0.0525 PD=0.873333 PS=0.67 NRD=0 NRS=32.8202 M=1 R=2.33333
+ SA=90001.1 SB=90000.5 A=0.0756 P=1.2 MULT=1
MM1009 N_A_1910_71#_M1009_d N_A_1688_97#_M1009_g N_VPWR_M1030_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2184 AS=0.180367 PD=2.2 PS=1.74667 NRD=0 NRS=16.4101 M=1
+ R=4.66667 SA=90000.7 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1041 A_2277_392# N_A_1910_71#_M1041_g N_VPWR_M1041_s VPB PSHORT L=0.18 W=1
+ AD=0.3775 AS=0.26 PD=1.755 PS=2.52 NRD=63.5128 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.8 A=0.18 P=2.36 MULT=1
MM1012 N_A_2385_74#_M1012_d N_A_1295_74#_M1012_g A_2277_392# VPB PSHORT L=0.18
+ W=1 AD=0.219366 AS=0.3775 PD=1.90845 PS=1.755 NRD=0 NRS=63.5128 M=1 R=5.55556
+ SA=90001.1 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1025 A_2571_508# N_A_1492_74#_M1025_g N_A_2385_74#_M1012_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0921338 PD=0.66 PS=0.801549 NRD=30.4759 NRS=38.6908 M=1
+ R=2.33333 SA=90001.6 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1037 N_VPWR_M1037_d N_A_547_301#_M1037_g A_2571_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.109992 AS=0.0504 PD=0.92717 PS=0.66 NRD=65.6601 NRS=30.4759 M=1 R=2.33333
+ SA=90002.1 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1034 N_A_547_301#_M1034_d N_A_2385_74#_M1034_g N_VPWR_M1037_d VPB PSHORT
+ L=0.18 W=0.64 AD=0.1664 AS=0.167608 PD=1.8 PS=1.41283 NRD=0 NRS=33.8446 M=1
+ R=3.55556 SA=90001.9 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1000 N_VPWR_M1000_d N_A_2385_74#_M1000_g N_Q_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3024 AS=0.2912 PD=2.78 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX42_noxref VNB VPB NWDIODE A=29.34 P=35.32
c_171 VNB 0 2.70131e-19 $X=0 $Y=0
c_324 VPB 0 8.71884e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__sedfxtp_1.pxi.spice"
*
.ends
*
*

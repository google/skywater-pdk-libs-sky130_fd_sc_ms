* File: sky130_fd_sc_ms__dlxtn_4.pxi.spice
* Created: Fri Aug 28 17:29:51 2020
* 
x_PM_SKY130_FD_SC_MS__DLXTN_4%D N_D_M1010_g N_D_M1011_g D N_D_c_158_n
+ N_D_c_159_n PM_SKY130_FD_SC_MS__DLXTN_4%D
x_PM_SKY130_FD_SC_MS__DLXTN_4%GATE_N N_GATE_N_M1006_g N_GATE_N_M1016_g GATE_N
+ N_GATE_N_c_186_n PM_SKY130_FD_SC_MS__DLXTN_4%GATE_N
x_PM_SKY130_FD_SC_MS__DLXTN_4%A_232_114# N_A_232_114#_M1016_d
+ N_A_232_114#_M1006_d N_A_232_114#_M1020_g N_A_232_114#_c_224_n
+ N_A_232_114#_M1005_g N_A_232_114#_c_225_n N_A_232_114#_M1001_g
+ N_A_232_114#_c_226_n N_A_232_114#_M1000_g N_A_232_114#_c_227_n
+ N_A_232_114#_c_228_n N_A_232_114#_c_229_n N_A_232_114#_c_230_n
+ N_A_232_114#_c_238_n N_A_232_114#_c_239_n N_A_232_114#_c_240_n
+ N_A_232_114#_c_241_n N_A_232_114#_c_242_n N_A_232_114#_c_243_n
+ N_A_232_114#_c_231_n N_A_232_114#_c_232_n N_A_232_114#_c_233_n
+ N_A_232_114#_c_234_n N_A_232_114#_c_235_n
+ PM_SKY130_FD_SC_MS__DLXTN_4%A_232_114#
x_PM_SKY130_FD_SC_MS__DLXTN_4%A_27_115# N_A_27_115#_M1010_s N_A_27_115#_M1011_s
+ N_A_27_115#_M1021_g N_A_27_115#_c_370_n N_A_27_115#_M1002_g
+ N_A_27_115#_c_380_n N_A_27_115#_c_371_n N_A_27_115#_c_398_n
+ N_A_27_115#_c_372_n N_A_27_115#_c_373_n N_A_27_115#_c_374_n
+ N_A_27_115#_c_375_n N_A_27_115#_c_376_n N_A_27_115#_c_382_n
+ N_A_27_115#_c_377_n N_A_27_115#_c_378_n PM_SKY130_FD_SC_MS__DLXTN_4%A_27_115#
x_PM_SKY130_FD_SC_MS__DLXTN_4%A_369_392# N_A_369_392#_M1005_s
+ N_A_369_392#_M1020_s N_A_369_392#_M1009_g N_A_369_392#_c_479_n
+ N_A_369_392#_M1008_g N_A_369_392#_c_480_n N_A_369_392#_c_488_n
+ N_A_369_392#_c_481_n N_A_369_392#_c_482_n N_A_369_392#_c_489_n
+ N_A_369_392#_c_483_n N_A_369_392#_c_484_n N_A_369_392#_c_485_n
+ N_A_369_392#_c_486_n PM_SKY130_FD_SC_MS__DLXTN_4%A_369_392#
x_PM_SKY130_FD_SC_MS__DLXTN_4%A_840_395# N_A_840_395#_M1007_s
+ N_A_840_395#_M1004_d N_A_840_395#_M1014_g N_A_840_395#_M1003_g
+ N_A_840_395#_M1013_g N_A_840_395#_M1012_g N_A_840_395#_c_576_n
+ N_A_840_395#_M1015_g N_A_840_395#_M1017_g N_A_840_395#_M1023_g
+ N_A_840_395#_M1018_g N_A_840_395#_M1025_g N_A_840_395#_M1019_g
+ N_A_840_395#_c_595_n N_A_840_395#_c_596_n N_A_840_395#_c_583_n
+ N_A_840_395#_c_584_n N_A_840_395#_c_597_n N_A_840_395#_c_585_n
+ N_A_840_395#_c_586_n N_A_840_395#_c_598_n N_A_840_395#_c_587_n
+ N_A_840_395#_c_632_p N_A_840_395#_c_588_n
+ PM_SKY130_FD_SC_MS__DLXTN_4%A_840_395#
x_PM_SKY130_FD_SC_MS__DLXTN_4%A_678_392# N_A_678_392#_M1001_d
+ N_A_678_392#_M1009_d N_A_678_392#_M1004_g N_A_678_392#_M1007_g
+ N_A_678_392#_M1024_g N_A_678_392#_M1022_g N_A_678_392#_c_729_n
+ N_A_678_392#_c_730_n N_A_678_392#_c_731_n N_A_678_392#_c_732_n
+ N_A_678_392#_c_733_n N_A_678_392#_c_738_n N_A_678_392#_c_734_n
+ N_A_678_392#_c_735_n PM_SKY130_FD_SC_MS__DLXTN_4%A_678_392#
x_PM_SKY130_FD_SC_MS__DLXTN_4%VPWR N_VPWR_M1011_d N_VPWR_M1020_d N_VPWR_M1014_d
+ N_VPWR_M1022_s N_VPWR_M1017_s N_VPWR_M1019_s N_VPWR_c_831_n N_VPWR_c_832_n
+ N_VPWR_c_833_n N_VPWR_c_834_n N_VPWR_c_835_n N_VPWR_c_836_n VPWR
+ N_VPWR_c_837_n N_VPWR_c_838_n N_VPWR_c_839_n N_VPWR_c_840_n N_VPWR_c_841_n
+ N_VPWR_c_842_n N_VPWR_c_843_n N_VPWR_c_844_n N_VPWR_c_845_n N_VPWR_c_846_n
+ N_VPWR_c_847_n N_VPWR_c_830_n PM_SKY130_FD_SC_MS__DLXTN_4%VPWR
x_PM_SKY130_FD_SC_MS__DLXTN_4%Q N_Q_M1013_d N_Q_M1023_d N_Q_M1012_d N_Q_M1018_d
+ N_Q_c_932_n N_Q_c_939_n N_Q_c_940_n N_Q_c_933_n N_Q_c_934_n N_Q_c_935_n
+ N_Q_c_941_n N_Q_c_936_n N_Q_c_937_n Q Q Q N_Q_c_944_n
+ PM_SKY130_FD_SC_MS__DLXTN_4%Q
x_PM_SKY130_FD_SC_MS__DLXTN_4%VGND N_VGND_M1010_d N_VGND_M1005_d N_VGND_M1003_d
+ N_VGND_M1024_d N_VGND_M1015_s N_VGND_M1025_s N_VGND_c_1005_n N_VGND_c_1006_n
+ N_VGND_c_1007_n N_VGND_c_1008_n N_VGND_c_1009_n N_VGND_c_1010_n
+ N_VGND_c_1011_n N_VGND_c_1012_n N_VGND_c_1013_n VGND N_VGND_c_1014_n
+ N_VGND_c_1015_n N_VGND_c_1016_n N_VGND_c_1017_n N_VGND_c_1018_n
+ N_VGND_c_1019_n N_VGND_c_1020_n N_VGND_c_1021_n N_VGND_c_1022_n
+ N_VGND_c_1023_n PM_SKY130_FD_SC_MS__DLXTN_4%VGND
cc_1 VNB N_D_M1010_g 0.0301791f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.85
cc_2 VNB N_D_M1011_g 0.00201979f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.54
cc_3 VNB N_D_c_158_n 0.00385705f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_4 VNB N_D_c_159_n 0.060667f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.465
cc_5 VNB N_GATE_N_M1016_g 0.0248735f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.54
cc_6 VNB GATE_N 0.00210952f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_GATE_N_c_186_n 0.0147706f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_8 VNB N_A_232_114#_c_224_n 0.0184509f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_9 VNB N_A_232_114#_c_225_n 0.0146603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_232_114#_c_226_n 0.010741f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_11 VNB N_A_232_114#_c_227_n 0.0315798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_232_114#_c_228_n 0.0078699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_232_114#_c_229_n 0.00995015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_232_114#_c_230_n 0.00246166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_232_114#_c_231_n 0.0390372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_232_114#_c_232_n 5.47787e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_232_114#_c_233_n 0.00385597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_232_114#_c_234_n 0.0373933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_232_114#_c_235_n 0.0699058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_115#_M1021_g 0.00682663f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_21 VNB N_A_27_115#_c_370_n 0.0158604f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_22 VNB N_A_27_115#_c_371_n 0.00858581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_115#_c_372_n 0.0302799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_115#_c_373_n 0.00508052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_115#_c_374_n 0.023918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_115#_c_375_n 0.00292455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_115#_c_376_n 0.00224314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_115#_c_377_n 0.00833773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_115#_c_378_n 0.061162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_369_392#_c_479_n 0.0203856f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_31 VNB N_A_369_392#_c_480_n 4.52811e-19 $X=-0.19 $Y=-0.245 $X2=0.525
+ $Y2=1.465
cc_32 VNB N_A_369_392#_c_481_n 0.00222566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_369_392#_c_482_n 0.00678992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_369_392#_c_483_n 0.00365986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_369_392#_c_484_n 0.0210765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_369_392#_c_485_n 0.00796467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_369_392#_c_486_n 0.0480288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_840_395#_M1003_g 0.0448479f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_39 VNB N_A_840_395#_M1013_g 0.0247252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_840_395#_M1012_g 5.39107e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_840_395#_c_576_n 0.0204821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_840_395#_M1015_g 0.0223921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_840_395#_M1017_g 5.05799e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_840_395#_M1023_g 0.0217972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_840_395#_M1018_g 4.78571e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_840_395#_M1025_g 0.0243109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_840_395#_M1019_g 5.20689e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_840_395#_c_583_n 0.00214537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_840_395#_c_584_n 0.00197273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_840_395#_c_585_n 0.0115825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_840_395#_c_586_n 0.0105365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_840_395#_c_587_n 0.00409951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_840_395#_c_588_n 0.0571456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_678_392#_M1007_g 0.0272194f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_55 VNB N_A_678_392#_M1024_g 0.0240565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_678_392#_c_729_n 0.0071265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_678_392#_c_730_n 2.95717e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_678_392#_c_731_n 0.0027358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_678_392#_c_732_n 0.00356499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_678_392#_c_733_n 0.00933825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_678_392#_c_734_n 0.00418601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_678_392#_c_735_n 0.0430674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VPWR_c_830_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_Q_c_932_n 0.00299103f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.465
cc_65 VNB N_Q_c_933_n 0.00315465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_Q_c_934_n 0.00244574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_Q_c_935_n 0.00253236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_Q_c_936_n 0.00875216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_Q_c_937_n 0.00219521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB Q 0.0258321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1005_n 0.0163672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1006_n 0.00988336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1007_n 0.0147111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1008_n 0.0061968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1009_n 0.00333063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1010_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1011_n 0.0296685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1012_n 0.0175031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1013_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1014_n 0.0195521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1015_n 0.0440818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1016_n 0.0436262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1017_n 0.0194943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1018_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1019_n 0.00631593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1020_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1021_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1022_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1023_n 0.453881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VPB N_D_M1011_g 0.0515638f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=2.54
cc_91 VPB N_D_c_158_n 0.00761464f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_92 VPB N_GATE_N_M1006_g 0.0363533f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.85
cc_93 VPB GATE_N 0.002419f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_94 VPB N_GATE_N_c_186_n 0.0155942f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_95 VPB N_A_232_114#_M1020_g 0.0277937f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_96 VPB N_A_232_114#_M1000_g 0.0578592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_A_232_114#_c_238_n 0.00668201f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_A_232_114#_c_239_n 0.00497786f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB N_A_232_114#_c_240_n 0.00204029f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_A_232_114#_c_241_n 0.00750386f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_A_232_114#_c_242_n 0.0301725f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A_232_114#_c_243_n 0.00691911f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB N_A_232_114#_c_232_n 0.00367977f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_232_114#_c_233_n 0.00174569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_232_114#_c_234_n 0.0181944f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_232_114#_c_235_n 0.0284749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_27_115#_M1021_g 0.031074f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_108 VPB N_A_27_115#_c_380_n 0.0358457f $X=-0.19 $Y=1.66 $X2=0.525 $Y2=1.465
cc_109 VPB N_A_27_115#_c_371_n 0.00559717f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_27_115#_c_382_n 0.0150907f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_369_392#_M1009_g 0.0209105f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_112 VPB N_A_369_392#_c_488_n 0.0203997f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_113 VPB N_A_369_392#_c_489_n 0.00695488f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_369_392#_c_483_n 0.00195856f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_369_392#_c_484_n 0.0136685f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_840_395#_M1014_g 0.0314297f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_117 VPB N_A_840_395#_M1003_g 0.00568598f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_118 VPB N_A_840_395#_M1012_g 0.0235404f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_840_395#_M1017_g 0.0225465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_840_395#_M1018_g 0.0216049f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_840_395#_M1019_g 0.0246711f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_840_395#_c_595_n 0.00525346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_840_395#_c_596_n 0.072084f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_840_395#_c_597_n 0.00171094f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_840_395#_c_598_n 0.00951883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_678_392#_M1004_g 0.0356434f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_127 VPB N_A_678_392#_M1022_g 0.0333267f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_678_392#_c_738_n 0.00162764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_678_392#_c_734_n 0.00325512f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_678_392#_c_735_n 0.0089239f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_831_n 0.00969617f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_832_n 0.0141076f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_833_n 0.00536824f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_834_n 0.00274039f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_835_n 0.0119967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_836_n 0.0340169f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_837_n 0.0197879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_838_n 0.0402815f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_839_n 0.0185359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_840_n 0.0183588f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_841_n 0.0159778f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_842_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_843_n 0.00862826f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_844_n 0.0377769f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_845_n 0.024389f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_846_n 0.00615051f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_847_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_830_n 0.0800364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_Q_c_939_n 0.00251554f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_Q_c_940_n 0.0029897f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_Q_c_941_n 0.00233077f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB Q 0.0085109f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB Q 0.0177184f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_Q_c_944_n 0.00254338f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 N_D_M1011_g N_GATE_N_M1006_g 0.0121914f $X=0.525 $Y=2.54 $X2=0 $Y2=0
cc_156 N_D_M1010_g N_GATE_N_M1016_g 0.0187327f $X=0.495 $Y=0.85 $X2=0 $Y2=0
cc_157 N_D_c_159_n N_GATE_N_M1016_g 0.00470907f $X=0.525 $Y=1.465 $X2=0 $Y2=0
cc_158 N_D_c_159_n N_GATE_N_c_186_n 0.0121914f $X=0.525 $Y=1.465 $X2=0 $Y2=0
cc_159 N_D_M1011_g N_A_232_114#_c_242_n 6.18071e-19 $X=0.525 $Y=2.54 $X2=0 $Y2=0
cc_160 N_D_M1011_g N_A_27_115#_c_380_n 0.0154244f $X=0.525 $Y=2.54 $X2=0 $Y2=0
cc_161 N_D_M1010_g N_A_27_115#_c_371_n 0.00436712f $X=0.495 $Y=0.85 $X2=0 $Y2=0
cc_162 N_D_c_158_n N_A_27_115#_c_371_n 0.036032f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_163 N_D_c_159_n N_A_27_115#_c_371_n 0.00955881f $X=0.525 $Y=1.465 $X2=0 $Y2=0
cc_164 N_D_M1010_g N_A_27_115#_c_372_n 0.0278868f $X=0.495 $Y=0.85 $X2=0 $Y2=0
cc_165 N_D_c_158_n N_A_27_115#_c_372_n 0.0279826f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_166 N_D_c_159_n N_A_27_115#_c_372_n 0.00435879f $X=0.525 $Y=1.465 $X2=0 $Y2=0
cc_167 N_D_M1010_g N_A_27_115#_c_373_n 7.68306e-19 $X=0.495 $Y=0.85 $X2=0 $Y2=0
cc_168 N_D_M1011_g N_A_27_115#_c_382_n 0.0220014f $X=0.525 $Y=2.54 $X2=0 $Y2=0
cc_169 N_D_c_158_n N_A_27_115#_c_382_n 0.0260287f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_170 N_D_c_159_n N_A_27_115#_c_382_n 0.00146215f $X=0.525 $Y=1.465 $X2=0 $Y2=0
cc_171 N_D_M1011_g N_VPWR_c_831_n 0.00343717f $X=0.525 $Y=2.54 $X2=0 $Y2=0
cc_172 N_D_M1011_g N_VPWR_c_837_n 0.005209f $X=0.525 $Y=2.54 $X2=0 $Y2=0
cc_173 N_D_M1011_g N_VPWR_c_830_n 0.00986386f $X=0.525 $Y=2.54 $X2=0 $Y2=0
cc_174 N_D_M1010_g N_VGND_c_1005_n 0.00130869f $X=0.495 $Y=0.85 $X2=0 $Y2=0
cc_175 N_D_M1010_g N_VGND_c_1014_n 0.00341528f $X=0.495 $Y=0.85 $X2=0 $Y2=0
cc_176 N_D_M1010_g N_VGND_c_1023_n 0.0048347f $X=0.495 $Y=0.85 $X2=0 $Y2=0
cc_177 N_GATE_N_M1016_g N_A_232_114#_c_228_n 0.00566256f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_178 GATE_N N_A_232_114#_c_228_n 0.0141427f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_179 N_GATE_N_c_186_n N_A_232_114#_c_228_n 0.00355095f $X=1.15 $Y=1.665 $X2=0
+ $Y2=0
cc_180 N_GATE_N_M1016_g N_A_232_114#_c_229_n 0.00371584f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_181 N_GATE_N_M1016_g N_A_232_114#_c_230_n 0.00359662f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_182 GATE_N N_A_232_114#_c_230_n 0.0260997f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_183 N_GATE_N_c_186_n N_A_232_114#_c_230_n 0.00135088f $X=1.15 $Y=1.665 $X2=0
+ $Y2=0
cc_184 N_GATE_N_M1006_g N_A_232_114#_c_238_n 2.35278e-19 $X=1.075 $Y=2.54 $X2=0
+ $Y2=0
cc_185 N_GATE_N_M1006_g N_A_232_114#_c_242_n 0.0170103f $X=1.075 $Y=2.54 $X2=0
+ $Y2=0
cc_186 GATE_N N_A_232_114#_c_242_n 0.0105591f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_187 N_GATE_N_c_186_n N_A_232_114#_c_242_n 0.00330449f $X=1.15 $Y=1.665 $X2=0
+ $Y2=0
cc_188 N_GATE_N_M1006_g N_A_232_114#_c_243_n 0.00801264f $X=1.075 $Y=2.54 $X2=0
+ $Y2=0
cc_189 N_GATE_N_M1016_g N_A_232_114#_c_231_n 0.0155068f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_190 GATE_N N_A_232_114#_c_235_n 2.97788e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_191 N_GATE_N_c_186_n N_A_232_114#_c_235_n 0.0149176f $X=1.15 $Y=1.665 $X2=0
+ $Y2=0
cc_192 N_GATE_N_M1006_g N_A_27_115#_c_380_n 6.00788e-19 $X=1.075 $Y=2.54 $X2=0
+ $Y2=0
cc_193 N_GATE_N_M1016_g N_A_27_115#_c_371_n 0.00516253f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_194 GATE_N N_A_27_115#_c_371_n 0.022773f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_195 N_GATE_N_c_186_n N_A_27_115#_c_371_n 0.00370129f $X=1.15 $Y=1.665 $X2=0
+ $Y2=0
cc_196 N_GATE_N_M1016_g N_A_27_115#_c_398_n 0.0140794f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_197 GATE_N N_A_27_115#_c_398_n 0.00313461f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_198 N_GATE_N_M1016_g N_A_27_115#_c_372_n 0.00639387f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_199 N_GATE_N_M1016_g N_A_27_115#_c_373_n 0.00773574f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_200 N_GATE_N_M1006_g N_A_27_115#_c_382_n 0.004281f $X=1.075 $Y=2.54 $X2=0
+ $Y2=0
cc_201 N_GATE_N_M1006_g N_VPWR_c_831_n 0.00343717f $X=1.075 $Y=2.54 $X2=0 $Y2=0
cc_202 N_GATE_N_M1006_g N_VPWR_c_838_n 0.005209f $X=1.075 $Y=2.54 $X2=0 $Y2=0
cc_203 N_GATE_N_M1006_g N_VPWR_c_830_n 0.00987709f $X=1.075 $Y=2.54 $X2=0 $Y2=0
cc_204 N_GATE_N_M1016_g N_VGND_c_1005_n 5.5317e-19 $X=1.085 $Y=0.94 $X2=0 $Y2=0
cc_205 N_GATE_N_M1016_g N_VGND_c_1015_n 0.00318127f $X=1.085 $Y=0.94 $X2=0 $Y2=0
cc_206 N_GATE_N_M1016_g N_VGND_c_1023_n 0.00438121f $X=1.085 $Y=0.94 $X2=0 $Y2=0
cc_207 N_A_232_114#_c_238_n N_A_27_115#_M1021_g 0.01509f $X=2.99 $Y=2.475 $X2=0
+ $Y2=0
cc_208 N_A_232_114#_c_240_n N_A_27_115#_M1021_g 0.0011759f $X=3.16 $Y=2.99 $X2=0
+ $Y2=0
cc_209 N_A_232_114#_c_235_n N_A_27_115#_M1021_g 0.0342524f $X=2.215 $Y=1.477
+ $X2=0 $Y2=0
cc_210 N_A_232_114#_c_224_n N_A_27_115#_c_370_n 0.00442933f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_211 N_A_232_114#_c_225_n N_A_27_115#_c_370_n 0.0227686f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_212 N_A_232_114#_c_242_n N_A_27_115#_c_380_n 0.00419744f $X=1.3 $Y=2.265
+ $X2=0 $Y2=0
cc_213 N_A_232_114#_c_228_n N_A_27_115#_c_371_n 0.00915345f $X=1.485 $Y=1.165
+ $X2=0 $Y2=0
cc_214 N_A_232_114#_M1016_d N_A_27_115#_c_398_n 0.00613024f $X=1.16 $Y=0.57
+ $X2=0 $Y2=0
cc_215 N_A_232_114#_c_228_n N_A_27_115#_c_398_n 0.00997713f $X=1.485 $Y=1.165
+ $X2=0 $Y2=0
cc_216 N_A_232_114#_c_229_n N_A_27_115#_c_398_n 0.00618319f $X=1.685 $Y=1.33
+ $X2=0 $Y2=0
cc_217 N_A_232_114#_c_231_n N_A_27_115#_c_398_n 2.54774e-19 $X=1.72 $Y=0.925
+ $X2=0 $Y2=0
cc_218 N_A_232_114#_c_228_n N_A_27_115#_c_372_n 0.00659465f $X=1.485 $Y=1.165
+ $X2=0 $Y2=0
cc_219 N_A_232_114#_M1016_d N_A_27_115#_c_373_n 0.00339584f $X=1.16 $Y=0.57
+ $X2=0 $Y2=0
cc_220 N_A_232_114#_c_224_n N_A_27_115#_c_374_n 0.0157054f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_221 N_A_232_114#_c_228_n N_A_27_115#_c_374_n 0.00552911f $X=1.485 $Y=1.165
+ $X2=0 $Y2=0
cc_222 N_A_232_114#_c_229_n N_A_27_115#_c_374_n 0.0169889f $X=1.685 $Y=1.33
+ $X2=0 $Y2=0
cc_223 N_A_232_114#_c_231_n N_A_27_115#_c_374_n 0.00199179f $X=1.72 $Y=0.925
+ $X2=0 $Y2=0
cc_224 N_A_232_114#_c_224_n N_A_27_115#_c_376_n 0.00730669f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_225 N_A_232_114#_c_242_n N_A_27_115#_c_382_n 9.83406e-19 $X=1.3 $Y=2.265
+ $X2=0 $Y2=0
cc_226 N_A_232_114#_c_235_n N_A_27_115#_c_377_n 0.00293022f $X=2.215 $Y=1.477
+ $X2=0 $Y2=0
cc_227 N_A_232_114#_c_224_n N_A_27_115#_c_378_n 0.00242956f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_228 N_A_232_114#_c_227_n N_A_27_115#_c_378_n 0.0227686f $X=3.855 $Y=1.185
+ $X2=0 $Y2=0
cc_229 N_A_232_114#_c_235_n N_A_27_115#_c_378_n 0.0131368f $X=2.215 $Y=1.477
+ $X2=0 $Y2=0
cc_230 N_A_232_114#_c_238_n N_A_369_392#_M1020_s 0.00732034f $X=2.99 $Y=2.475
+ $X2=0 $Y2=0
cc_231 N_A_232_114#_M1000_g N_A_369_392#_M1009_g 0.0265964f $X=3.87 $Y=2.75
+ $X2=0 $Y2=0
cc_232 N_A_232_114#_c_239_n N_A_369_392#_M1009_g 0.0146467f $X=4.05 $Y=2.99
+ $X2=0 $Y2=0
cc_233 N_A_232_114#_c_225_n N_A_369_392#_c_479_n 0.00527673f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_234 N_A_232_114#_c_227_n N_A_369_392#_c_479_n 0.00161375f $X=3.855 $Y=1.185
+ $X2=0 $Y2=0
cc_235 N_A_232_114#_c_233_n N_A_369_392#_c_479_n 2.45027e-19 $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_236 N_A_232_114#_c_234_n N_A_369_392#_c_479_n 0.00312708f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_237 N_A_232_114#_c_224_n N_A_369_392#_c_480_n 0.00940637f $X=2.355 $Y=1.185
+ $X2=0 $Y2=0
cc_238 N_A_232_114#_c_229_n N_A_369_392#_c_480_n 0.044954f $X=1.685 $Y=1.33
+ $X2=0 $Y2=0
cc_239 N_A_232_114#_c_230_n N_A_369_392#_c_480_n 0.0289818f $X=1.685 $Y=1.57
+ $X2=0 $Y2=0
cc_240 N_A_232_114#_c_231_n N_A_369_392#_c_480_n 0.00156461f $X=1.72 $Y=0.925
+ $X2=0 $Y2=0
cc_241 N_A_232_114#_c_235_n N_A_369_392#_c_480_n 0.0278331f $X=2.215 $Y=1.477
+ $X2=0 $Y2=0
cc_242 N_A_232_114#_c_238_n N_A_369_392#_c_488_n 0.0256967f $X=2.99 $Y=2.475
+ $X2=0 $Y2=0
cc_243 N_A_232_114#_c_235_n N_A_369_392#_c_488_n 0.00411697f $X=2.215 $Y=1.477
+ $X2=0 $Y2=0
cc_244 N_A_232_114#_c_225_n N_A_369_392#_c_482_n 0.0173976f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_245 N_A_232_114#_c_227_n N_A_369_392#_c_482_n 6.03378e-19 $X=3.855 $Y=1.185
+ $X2=0 $Y2=0
cc_246 N_A_232_114#_M1020_g N_A_369_392#_c_489_n 0.0197697f $X=2.215 $Y=2.38
+ $X2=0 $Y2=0
cc_247 N_A_232_114#_c_238_n N_A_369_392#_c_489_n 0.0286499f $X=2.99 $Y=2.475
+ $X2=0 $Y2=0
cc_248 N_A_232_114#_c_243_n N_A_369_392#_c_489_n 0.0311122f $X=1.395 $Y=2.1
+ $X2=0 $Y2=0
cc_249 N_A_232_114#_c_232_n N_A_369_392#_c_489_n 0.00896259f $X=1.72 $Y=1.605
+ $X2=0 $Y2=0
cc_250 N_A_232_114#_c_235_n N_A_369_392#_c_489_n 0.0121398f $X=2.215 $Y=1.477
+ $X2=0 $Y2=0
cc_251 N_A_232_114#_M1000_g N_A_369_392#_c_483_n 2.90398e-19 $X=3.87 $Y=2.75
+ $X2=0 $Y2=0
cc_252 N_A_232_114#_c_234_n N_A_369_392#_c_483_n 3.62762e-19 $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_253 N_A_232_114#_c_227_n N_A_369_392#_c_484_n 6.79409e-19 $X=3.855 $Y=1.185
+ $X2=0 $Y2=0
cc_254 N_A_232_114#_c_234_n N_A_369_392#_c_484_n 0.0173938f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_255 N_A_232_114#_c_225_n N_A_369_392#_c_485_n 0.00376963f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_256 N_A_232_114#_c_226_n N_A_369_392#_c_485_n 0.00118688f $X=3.855 $Y=1.405
+ $X2=0 $Y2=0
cc_257 N_A_232_114#_c_225_n N_A_369_392#_c_486_n 0.00586767f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_258 N_A_232_114#_c_239_n N_A_840_395#_M1014_g 0.003725f $X=4.05 $Y=2.99 $X2=0
+ $Y2=0
cc_259 N_A_232_114#_c_241_n N_A_840_395#_M1014_g 0.0188065f $X=4.135 $Y=2.905
+ $X2=0 $Y2=0
cc_260 N_A_232_114#_c_241_n N_A_840_395#_M1003_g 6.0243e-19 $X=4.135 $Y=2.905
+ $X2=0 $Y2=0
cc_261 N_A_232_114#_c_233_n N_A_840_395#_M1003_g 7.74691e-19 $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_262 N_A_232_114#_c_234_n N_A_840_395#_M1003_g 0.0136936f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_263 N_A_232_114#_c_241_n N_A_840_395#_c_595_n 0.0249855f $X=4.135 $Y=2.905
+ $X2=0 $Y2=0
cc_264 N_A_232_114#_M1000_g N_A_840_395#_c_596_n 0.0587776f $X=3.87 $Y=2.75
+ $X2=0 $Y2=0
cc_265 N_A_232_114#_c_241_n N_A_840_395#_c_596_n 0.0113486f $X=4.135 $Y=2.905
+ $X2=0 $Y2=0
cc_266 N_A_232_114#_c_233_n N_A_840_395#_c_596_n 0.00120658f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_267 N_A_232_114#_c_234_n N_A_840_395#_c_596_n 0.0101853f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_268 N_A_232_114#_c_239_n N_A_678_392#_M1009_d 0.0030236f $X=4.05 $Y=2.99
+ $X2=0 $Y2=0
cc_269 N_A_232_114#_c_227_n N_A_678_392#_c_729_n 0.00249179f $X=3.855 $Y=1.185
+ $X2=0 $Y2=0
cc_270 N_A_232_114#_c_233_n N_A_678_392#_c_729_n 0.0154026f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_271 N_A_232_114#_c_234_n N_A_678_392#_c_729_n 0.00598369f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_272 N_A_232_114#_c_225_n N_A_678_392#_c_730_n 0.00514497f $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_273 N_A_232_114#_c_227_n N_A_678_392#_c_730_n 0.00126393f $X=3.855 $Y=1.185
+ $X2=0 $Y2=0
cc_274 N_A_232_114#_c_227_n N_A_678_392#_c_731_n 0.00254147f $X=3.855 $Y=1.185
+ $X2=0 $Y2=0
cc_275 N_A_232_114#_c_226_n N_A_678_392#_c_732_n 0.00128751f $X=3.855 $Y=1.405
+ $X2=0 $Y2=0
cc_276 N_A_232_114#_c_233_n N_A_678_392#_c_732_n 0.0206617f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_277 N_A_232_114#_c_234_n N_A_678_392#_c_732_n 0.00196022f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_278 N_A_232_114#_M1000_g N_A_678_392#_c_738_n 0.0223877f $X=3.87 $Y=2.75
+ $X2=0 $Y2=0
cc_279 N_A_232_114#_c_239_n N_A_678_392#_c_738_n 0.0300777f $X=4.05 $Y=2.99
+ $X2=0 $Y2=0
cc_280 N_A_232_114#_c_241_n N_A_678_392#_c_738_n 0.0494986f $X=4.135 $Y=2.905
+ $X2=0 $Y2=0
cc_281 N_A_232_114#_c_225_n N_A_678_392#_c_734_n 6.76373e-19 $X=3.605 $Y=1.11
+ $X2=0 $Y2=0
cc_282 N_A_232_114#_c_226_n N_A_678_392#_c_734_n 0.00615882f $X=3.855 $Y=1.405
+ $X2=0 $Y2=0
cc_283 N_A_232_114#_M1000_g N_A_678_392#_c_734_n 0.00750246f $X=3.87 $Y=2.75
+ $X2=0 $Y2=0
cc_284 N_A_232_114#_c_227_n N_A_678_392#_c_734_n 0.0117959f $X=3.855 $Y=1.185
+ $X2=0 $Y2=0
cc_285 N_A_232_114#_c_233_n N_A_678_392#_c_734_n 0.0494986f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_286 N_A_232_114#_c_234_n N_A_678_392#_c_734_n 0.00971643f $X=4.215 $Y=1.57
+ $X2=0 $Y2=0
cc_287 N_A_232_114#_c_238_n N_VPWR_M1020_d 0.0117295f $X=2.99 $Y=2.475 $X2=0
+ $Y2=0
cc_288 N_A_232_114#_c_242_n N_VPWR_c_831_n 0.0285454f $X=1.3 $Y=2.265 $X2=0
+ $Y2=0
cc_289 N_A_232_114#_M1020_g N_VPWR_c_832_n 0.00458264f $X=2.215 $Y=2.38 $X2=0
+ $Y2=0
cc_290 N_A_232_114#_c_238_n N_VPWR_c_832_n 0.0314893f $X=2.99 $Y=2.475 $X2=0
+ $Y2=0
cc_291 N_A_232_114#_c_240_n N_VPWR_c_832_n 0.0120576f $X=3.16 $Y=2.99 $X2=0
+ $Y2=0
cc_292 N_A_232_114#_M1020_g N_VPWR_c_838_n 0.00562877f $X=2.215 $Y=2.38 $X2=0
+ $Y2=0
cc_293 N_A_232_114#_c_242_n N_VPWR_c_838_n 0.0230269f $X=1.3 $Y=2.265 $X2=0
+ $Y2=0
cc_294 N_A_232_114#_M1000_g N_VPWR_c_844_n 0.00333926f $X=3.87 $Y=2.75 $X2=0
+ $Y2=0
cc_295 N_A_232_114#_c_239_n N_VPWR_c_844_n 0.0682836f $X=4.05 $Y=2.99 $X2=0
+ $Y2=0
cc_296 N_A_232_114#_c_240_n N_VPWR_c_844_n 0.0121935f $X=3.16 $Y=2.99 $X2=0
+ $Y2=0
cc_297 N_A_232_114#_c_239_n N_VPWR_c_845_n 0.0125322f $X=4.05 $Y=2.99 $X2=0
+ $Y2=0
cc_298 N_A_232_114#_M1020_g N_VPWR_c_830_n 0.00595788f $X=2.215 $Y=2.38 $X2=0
+ $Y2=0
cc_299 N_A_232_114#_M1000_g N_VPWR_c_830_n 0.00423643f $X=3.87 $Y=2.75 $X2=0
+ $Y2=0
cc_300 N_A_232_114#_c_238_n N_VPWR_c_830_n 0.0321309f $X=2.99 $Y=2.475 $X2=0
+ $Y2=0
cc_301 N_A_232_114#_c_239_n N_VPWR_c_830_n 0.0383253f $X=4.05 $Y=2.99 $X2=0
+ $Y2=0
cc_302 N_A_232_114#_c_240_n N_VPWR_c_830_n 0.00661049f $X=3.16 $Y=2.99 $X2=0
+ $Y2=0
cc_303 N_A_232_114#_c_242_n N_VPWR_c_830_n 0.0189916f $X=1.3 $Y=2.265 $X2=0
+ $Y2=0
cc_304 N_A_232_114#_c_238_n A_594_392# 0.00241277f $X=2.99 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_305 N_A_232_114#_c_239_n A_792_508# 0.00122098f $X=4.05 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_306 N_A_232_114#_c_241_n A_792_508# 0.00347384f $X=4.135 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_307 N_A_232_114#_c_224_n N_VGND_c_1006_n 0.00195643f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_308 N_A_232_114#_c_225_n N_VGND_c_1006_n 3.35588e-19 $X=3.605 $Y=1.11 $X2=0
+ $Y2=0
cc_309 N_A_232_114#_c_224_n N_VGND_c_1015_n 0.00278271f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_310 N_A_232_114#_c_225_n N_VGND_c_1016_n 9.44495e-19 $X=3.605 $Y=1.11 $X2=0
+ $Y2=0
cc_311 N_A_232_114#_c_224_n N_VGND_c_1023_n 0.00363426f $X=2.355 $Y=1.185 $X2=0
+ $Y2=0
cc_312 N_A_27_115#_c_374_n N_A_369_392#_M1005_s 0.00441657f $X=2.475 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_313 N_A_27_115#_M1021_g N_A_369_392#_c_480_n 9.39281e-19 $X=2.88 $Y=2.46
+ $X2=0 $Y2=0
cc_314 N_A_27_115#_c_374_n N_A_369_392#_c_480_n 0.0144209f $X=2.475 $Y=0.34
+ $X2=0 $Y2=0
cc_315 N_A_27_115#_c_376_n N_A_369_392#_c_480_n 0.0265397f $X=2.56 $Y=1.22 $X2=0
+ $Y2=0
cc_316 N_A_27_115#_c_377_n N_A_369_392#_c_480_n 0.0265613f $X=2.835 $Y=1.385
+ $X2=0 $Y2=0
cc_317 N_A_27_115#_c_378_n N_A_369_392#_c_480_n 2.87669e-19 $X=2.88 $Y=1.33
+ $X2=0 $Y2=0
cc_318 N_A_27_115#_M1021_g N_A_369_392#_c_488_n 0.0143931f $X=2.88 $Y=2.46 $X2=0
+ $Y2=0
cc_319 N_A_27_115#_c_377_n N_A_369_392#_c_488_n 0.0395884f $X=2.835 $Y=1.385
+ $X2=0 $Y2=0
cc_320 N_A_27_115#_c_378_n N_A_369_392#_c_488_n 0.00785784f $X=2.88 $Y=1.33
+ $X2=0 $Y2=0
cc_321 N_A_27_115#_c_370_n N_A_369_392#_c_481_n 0.00147103f $X=3.215 $Y=1.11
+ $X2=0 $Y2=0
cc_322 N_A_27_115#_M1021_g N_A_369_392#_c_489_n 0.00160177f $X=2.88 $Y=2.46
+ $X2=0 $Y2=0
cc_323 N_A_27_115#_M1021_g N_A_369_392#_c_483_n 0.00123314f $X=2.88 $Y=2.46
+ $X2=0 $Y2=0
cc_324 N_A_27_115#_c_377_n N_A_369_392#_c_483_n 0.00521207f $X=2.835 $Y=1.385
+ $X2=0 $Y2=0
cc_325 N_A_27_115#_c_378_n N_A_369_392#_c_483_n 7.06729e-19 $X=2.88 $Y=1.33
+ $X2=0 $Y2=0
cc_326 N_A_27_115#_M1021_g N_A_369_392#_c_484_n 0.0803546f $X=2.88 $Y=2.46 $X2=0
+ $Y2=0
cc_327 N_A_27_115#_c_377_n N_A_369_392#_c_484_n 2.74972e-19 $X=2.835 $Y=1.385
+ $X2=0 $Y2=0
cc_328 N_A_27_115#_c_378_n N_A_369_392#_c_484_n 0.0104185f $X=2.88 $Y=1.33 $X2=0
+ $Y2=0
cc_329 N_A_27_115#_c_370_n N_A_369_392#_c_485_n 0.00497566f $X=3.215 $Y=1.11
+ $X2=0 $Y2=0
cc_330 N_A_27_115#_c_376_n N_A_369_392#_c_485_n 0.00474149f $X=2.56 $Y=1.22
+ $X2=0 $Y2=0
cc_331 N_A_27_115#_c_377_n N_A_369_392#_c_485_n 0.0122394f $X=2.835 $Y=1.385
+ $X2=0 $Y2=0
cc_332 N_A_27_115#_c_378_n N_A_369_392#_c_485_n 0.00129573f $X=2.88 $Y=1.33
+ $X2=0 $Y2=0
cc_333 N_A_27_115#_M1021_g N_A_678_392#_c_738_n 0.00176441f $X=2.88 $Y=2.46
+ $X2=0 $Y2=0
cc_334 N_A_27_115#_c_380_n N_VPWR_c_831_n 0.0266809f $X=0.3 $Y=2.265 $X2=0 $Y2=0
cc_335 N_A_27_115#_c_382_n N_VPWR_c_831_n 0.0114941f $X=0.71 $Y=2.035 $X2=0
+ $Y2=0
cc_336 N_A_27_115#_M1021_g N_VPWR_c_832_n 0.0118711f $X=2.88 $Y=2.46 $X2=0 $Y2=0
cc_337 N_A_27_115#_c_380_n N_VPWR_c_837_n 0.014549f $X=0.3 $Y=2.265 $X2=0 $Y2=0
cc_338 N_A_27_115#_M1021_g N_VPWR_c_844_n 0.00460063f $X=2.88 $Y=2.46 $X2=0
+ $Y2=0
cc_339 N_A_27_115#_M1021_g N_VPWR_c_830_n 0.00443063f $X=2.88 $Y=2.46 $X2=0
+ $Y2=0
cc_340 N_A_27_115#_c_380_n N_VPWR_c_830_n 0.0119743f $X=0.3 $Y=2.265 $X2=0 $Y2=0
cc_341 N_A_27_115#_c_371_n N_VGND_M1010_d 0.00236148f $X=0.71 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_342 N_A_27_115#_c_398_n N_VGND_M1010_d 0.007918f $X=1.145 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_343 N_A_27_115#_c_372_n N_VGND_M1010_d 0.00690665f $X=0.795 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_344 N_A_27_115#_c_374_n N_VGND_M1005_d 6.47853e-19 $X=2.475 $Y=0.34 $X2=0
+ $Y2=0
cc_345 N_A_27_115#_c_376_n N_VGND_M1005_d 0.0110808f $X=2.56 $Y=1.22 $X2=0 $Y2=0
cc_346 N_A_27_115#_c_398_n N_VGND_c_1005_n 0.0121815f $X=1.145 $Y=0.745 $X2=0
+ $Y2=0
cc_347 N_A_27_115#_c_372_n N_VGND_c_1005_n 0.0143324f $X=0.795 $Y=0.745 $X2=0
+ $Y2=0
cc_348 N_A_27_115#_c_373_n N_VGND_c_1005_n 0.0045384f $X=1.23 $Y=0.66 $X2=0
+ $Y2=0
cc_349 N_A_27_115#_c_375_n N_VGND_c_1005_n 0.0139003f $X=1.315 $Y=0.34 $X2=0
+ $Y2=0
cc_350 N_A_27_115#_c_370_n N_VGND_c_1006_n 0.0092719f $X=3.215 $Y=1.11 $X2=0
+ $Y2=0
cc_351 N_A_27_115#_c_374_n N_VGND_c_1006_n 0.0148948f $X=2.475 $Y=0.34 $X2=0
+ $Y2=0
cc_352 N_A_27_115#_c_376_n N_VGND_c_1006_n 0.0477502f $X=2.56 $Y=1.22 $X2=0
+ $Y2=0
cc_353 N_A_27_115#_c_377_n N_VGND_c_1006_n 0.0155155f $X=2.835 $Y=1.385 $X2=0
+ $Y2=0
cc_354 N_A_27_115#_c_378_n N_VGND_c_1006_n 0.00987931f $X=2.88 $Y=1.33 $X2=0
+ $Y2=0
cc_355 N_A_27_115#_c_372_n N_VGND_c_1014_n 0.0103718f $X=0.795 $Y=0.745 $X2=0
+ $Y2=0
cc_356 N_A_27_115#_c_398_n N_VGND_c_1015_n 0.00257035f $X=1.145 $Y=0.745 $X2=0
+ $Y2=0
cc_357 N_A_27_115#_c_374_n N_VGND_c_1015_n 0.086417f $X=2.475 $Y=0.34 $X2=0
+ $Y2=0
cc_358 N_A_27_115#_c_375_n N_VGND_c_1015_n 0.0120335f $X=1.315 $Y=0.34 $X2=0
+ $Y2=0
cc_359 N_A_27_115#_c_370_n N_VGND_c_1016_n 0.00539704f $X=3.215 $Y=1.11 $X2=0
+ $Y2=0
cc_360 N_A_27_115#_c_370_n N_VGND_c_1023_n 0.0052351f $X=3.215 $Y=1.11 $X2=0
+ $Y2=0
cc_361 N_A_27_115#_c_398_n N_VGND_c_1023_n 0.00589268f $X=1.145 $Y=0.745 $X2=0
+ $Y2=0
cc_362 N_A_27_115#_c_372_n N_VGND_c_1023_n 0.0164998f $X=0.795 $Y=0.745 $X2=0
+ $Y2=0
cc_363 N_A_27_115#_c_374_n N_VGND_c_1023_n 0.049532f $X=2.475 $Y=0.34 $X2=0
+ $Y2=0
cc_364 N_A_27_115#_c_375_n N_VGND_c_1023_n 0.00658039f $X=1.315 $Y=0.34 $X2=0
+ $Y2=0
cc_365 N_A_369_392#_c_486_n N_A_840_395#_M1003_g 0.0424929f $X=4.4 $Y=0.34 $X2=0
+ $Y2=0
cc_366 N_A_369_392#_c_482_n N_A_678_392#_M1001_d 0.00252704f $X=4.28 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_367 N_A_369_392#_c_486_n N_A_678_392#_M1007_g 0.00207621f $X=4.4 $Y=0.34
+ $X2=0 $Y2=0
cc_368 N_A_369_392#_c_479_n N_A_678_392#_c_729_n 0.0151004f $X=4.4 $Y=0.505
+ $X2=0 $Y2=0
cc_369 N_A_369_392#_c_482_n N_A_678_392#_c_729_n 0.0316369f $X=4.28 $Y=0.34
+ $X2=0 $Y2=0
cc_370 N_A_369_392#_c_486_n N_A_678_392#_c_729_n 0.00447421f $X=4.4 $Y=0.34
+ $X2=0 $Y2=0
cc_371 N_A_369_392#_c_482_n N_A_678_392#_c_730_n 0.0105171f $X=4.28 $Y=0.34
+ $X2=0 $Y2=0
cc_372 N_A_369_392#_c_485_n N_A_678_392#_c_730_n 0.0146188f $X=3.375 $Y=1.47
+ $X2=0 $Y2=0
cc_373 N_A_369_392#_c_479_n N_A_678_392#_c_731_n 0.0012686f $X=4.4 $Y=0.505
+ $X2=0 $Y2=0
cc_374 N_A_369_392#_M1009_g N_A_678_392#_c_738_n 0.0112988f $X=3.3 $Y=2.46 $X2=0
+ $Y2=0
cc_375 N_A_369_392#_c_483_n N_A_678_392#_c_738_n 0.0133577f $X=3.375 $Y=1.635
+ $X2=0 $Y2=0
cc_376 N_A_369_392#_c_484_n N_A_678_392#_c_738_n 7.89148e-19 $X=3.375 $Y=1.635
+ $X2=0 $Y2=0
cc_377 N_A_369_392#_M1009_g N_A_678_392#_c_734_n 0.00320718f $X=3.3 $Y=2.46
+ $X2=0 $Y2=0
cc_378 N_A_369_392#_c_479_n N_A_678_392#_c_734_n 6.66919e-19 $X=4.4 $Y=0.505
+ $X2=0 $Y2=0
cc_379 N_A_369_392#_c_483_n N_A_678_392#_c_734_n 0.031936f $X=3.375 $Y=1.635
+ $X2=0 $Y2=0
cc_380 N_A_369_392#_c_484_n N_A_678_392#_c_734_n 0.00187211f $X=3.375 $Y=1.635
+ $X2=0 $Y2=0
cc_381 N_A_369_392#_c_485_n N_A_678_392#_c_734_n 0.0250348f $X=3.375 $Y=1.47
+ $X2=0 $Y2=0
cc_382 N_A_369_392#_M1009_g N_VPWR_c_832_n 2.60877e-19 $X=3.3 $Y=2.46 $X2=0
+ $Y2=0
cc_383 N_A_369_392#_M1009_g N_VPWR_c_844_n 0.00333926f $X=3.3 $Y=2.46 $X2=0
+ $Y2=0
cc_384 N_A_369_392#_M1009_g N_VPWR_c_830_n 0.00423643f $X=3.3 $Y=2.46 $X2=0
+ $Y2=0
cc_385 N_A_369_392#_c_488_n N_VGND_c_1006_n 0.00457271f $X=3.21 $Y=1.805 $X2=0
+ $Y2=0
cc_386 N_A_369_392#_c_481_n N_VGND_c_1006_n 0.0159466f $X=3.485 $Y=0.38 $X2=0
+ $Y2=0
cc_387 N_A_369_392#_c_485_n N_VGND_c_1006_n 0.0209764f $X=3.375 $Y=1.47 $X2=0
+ $Y2=0
cc_388 N_A_369_392#_c_482_n N_VGND_c_1007_n 0.0098708f $X=4.28 $Y=0.34 $X2=0
+ $Y2=0
cc_389 N_A_369_392#_c_486_n N_VGND_c_1007_n 0.00431935f $X=4.4 $Y=0.34 $X2=0
+ $Y2=0
cc_390 N_A_369_392#_c_481_n N_VGND_c_1016_n 0.0121867f $X=3.485 $Y=0.38 $X2=0
+ $Y2=0
cc_391 N_A_369_392#_c_482_n N_VGND_c_1016_n 0.062486f $X=4.28 $Y=0.34 $X2=0
+ $Y2=0
cc_392 N_A_369_392#_c_486_n N_VGND_c_1016_n 0.00730902f $X=4.4 $Y=0.34 $X2=0
+ $Y2=0
cc_393 N_A_369_392#_c_481_n N_VGND_c_1023_n 0.00660921f $X=3.485 $Y=0.38 $X2=0
+ $Y2=0
cc_394 N_A_369_392#_c_482_n N_VGND_c_1023_n 0.0348893f $X=4.28 $Y=0.34 $X2=0
+ $Y2=0
cc_395 N_A_369_392#_c_486_n N_VGND_c_1023_n 0.0113113f $X=4.4 $Y=0.34 $X2=0
+ $Y2=0
cc_396 N_A_369_392#_c_485_n A_658_79# 0.00247748f $X=3.375 $Y=1.47 $X2=-0.19
+ $Y2=-0.245
cc_397 N_A_840_395#_c_595_n N_A_678_392#_M1004_g 0.0237588f $X=5.315 $Y=2.14
+ $X2=0 $Y2=0
cc_398 N_A_840_395#_c_596_n N_A_678_392#_M1004_g 0.0193515f $X=4.555 $Y=2.14
+ $X2=0 $Y2=0
cc_399 N_A_840_395#_c_598_n N_A_678_392#_M1004_g 0.00608885f $X=5.48 $Y=2.265
+ $X2=0 $Y2=0
cc_400 N_A_840_395#_M1003_g N_A_678_392#_M1007_g 0.0178603f $X=4.76 $Y=0.825
+ $X2=0 $Y2=0
cc_401 N_A_840_395#_c_583_n N_A_678_392#_M1007_g 0.00687953f $X=5.485 $Y=0.54
+ $X2=0 $Y2=0
cc_402 N_A_840_395#_c_584_n N_A_678_392#_M1007_g 9.92594e-19 $X=5.745 $Y=1.32
+ $X2=0 $Y2=0
cc_403 N_A_840_395#_c_587_n N_A_678_392#_M1007_g 0.00431125f $X=5.745 $Y=1.065
+ $X2=0 $Y2=0
cc_404 N_A_840_395#_M1013_g N_A_678_392#_M1024_g 0.0239087f $X=6.215 $Y=0.74
+ $X2=0 $Y2=0
cc_405 N_A_840_395#_c_584_n N_A_678_392#_M1024_g 0.00552835f $X=5.745 $Y=1.32
+ $X2=0 $Y2=0
cc_406 N_A_840_395#_c_587_n N_A_678_392#_M1024_g 0.0120291f $X=5.745 $Y=1.065
+ $X2=0 $Y2=0
cc_407 N_A_840_395#_c_597_n N_A_678_392#_M1022_g 0.00253684f $X=5.745 $Y=1.82
+ $X2=0 $Y2=0
cc_408 N_A_840_395#_c_598_n N_A_678_392#_M1022_g 0.0303956f $X=5.48 $Y=2.265
+ $X2=0 $Y2=0
cc_409 N_A_840_395#_M1003_g N_A_678_392#_c_729_n 0.00733517f $X=4.76 $Y=0.825
+ $X2=0 $Y2=0
cc_410 N_A_840_395#_M1003_g N_A_678_392#_c_731_n 0.00826027f $X=4.76 $Y=0.825
+ $X2=0 $Y2=0
cc_411 N_A_840_395#_c_587_n N_A_678_392#_c_731_n 0.00244264f $X=5.745 $Y=1.065
+ $X2=0 $Y2=0
cc_412 N_A_840_395#_M1003_g N_A_678_392#_c_732_n 0.00512512f $X=4.76 $Y=0.825
+ $X2=0 $Y2=0
cc_413 N_A_840_395#_c_595_n N_A_678_392#_c_732_n 0.00868744f $X=5.315 $Y=2.14
+ $X2=0 $Y2=0
cc_414 N_A_840_395#_c_596_n N_A_678_392#_c_732_n 0.0034639f $X=4.555 $Y=2.14
+ $X2=0 $Y2=0
cc_415 N_A_840_395#_M1003_g N_A_678_392#_c_733_n 0.0152674f $X=4.76 $Y=0.825
+ $X2=0 $Y2=0
cc_416 N_A_840_395#_c_595_n N_A_678_392#_c_733_n 0.0294526f $X=5.315 $Y=2.14
+ $X2=0 $Y2=0
cc_417 N_A_840_395#_c_598_n N_A_678_392#_c_733_n 0.01476f $X=5.48 $Y=2.265 $X2=0
+ $Y2=0
cc_418 N_A_840_395#_c_587_n N_A_678_392#_c_733_n 0.0126845f $X=5.745 $Y=1.065
+ $X2=0 $Y2=0
cc_419 N_A_840_395#_c_632_p N_A_678_392#_c_733_n 0.0277655f $X=5.745 $Y=1.485
+ $X2=0 $Y2=0
cc_420 N_A_840_395#_M1014_g N_A_678_392#_c_738_n 3.23029e-19 $X=4.29 $Y=2.75
+ $X2=0 $Y2=0
cc_421 N_A_840_395#_c_596_n N_A_678_392#_c_734_n 3.23029e-19 $X=4.555 $Y=2.14
+ $X2=0 $Y2=0
cc_422 N_A_840_395#_M1003_g N_A_678_392#_c_735_n 0.0186005f $X=4.76 $Y=0.825
+ $X2=0 $Y2=0
cc_423 N_A_840_395#_M1012_g N_A_678_392#_c_735_n 0.0243781f $X=6.23 $Y=2.4 $X2=0
+ $Y2=0
cc_424 N_A_840_395#_c_597_n N_A_678_392#_c_735_n 0.00389059f $X=5.745 $Y=1.82
+ $X2=0 $Y2=0
cc_425 N_A_840_395#_c_585_n N_A_678_392#_c_735_n 0.0110379f $X=6.305 $Y=1.485
+ $X2=0 $Y2=0
cc_426 N_A_840_395#_c_598_n N_A_678_392#_c_735_n 0.00393379f $X=5.48 $Y=2.265
+ $X2=0 $Y2=0
cc_427 N_A_840_395#_c_587_n N_A_678_392#_c_735_n 0.00257842f $X=5.745 $Y=1.065
+ $X2=0 $Y2=0
cc_428 N_A_840_395#_c_632_p N_A_678_392#_c_735_n 0.0142276f $X=5.745 $Y=1.485
+ $X2=0 $Y2=0
cc_429 N_A_840_395#_c_595_n N_VPWR_M1014_d 0.00265897f $X=5.315 $Y=2.14 $X2=0
+ $Y2=0
cc_430 N_A_840_395#_M1012_g N_VPWR_c_833_n 0.0161012f $X=6.23 $Y=2.4 $X2=0 $Y2=0
cc_431 N_A_840_395#_M1017_g N_VPWR_c_833_n 4.98184e-19 $X=6.755 $Y=2.4 $X2=0
+ $Y2=0
cc_432 N_A_840_395#_c_586_n N_VPWR_c_833_n 0.0103183f $X=7.325 $Y=1.485 $X2=0
+ $Y2=0
cc_433 N_A_840_395#_c_598_n N_VPWR_c_833_n 0.0613366f $X=5.48 $Y=2.265 $X2=0
+ $Y2=0
cc_434 N_A_840_395#_M1012_g N_VPWR_c_834_n 5.54949e-19 $X=6.23 $Y=2.4 $X2=0
+ $Y2=0
cc_435 N_A_840_395#_M1017_g N_VPWR_c_834_n 0.0159367f $X=6.755 $Y=2.4 $X2=0
+ $Y2=0
cc_436 N_A_840_395#_M1018_g N_VPWR_c_834_n 0.0156265f $X=7.205 $Y=2.4 $X2=0
+ $Y2=0
cc_437 N_A_840_395#_M1019_g N_VPWR_c_834_n 5.45866e-19 $X=7.655 $Y=2.4 $X2=0
+ $Y2=0
cc_438 N_A_840_395#_M1018_g N_VPWR_c_836_n 5.02386e-19 $X=7.205 $Y=2.4 $X2=0
+ $Y2=0
cc_439 N_A_840_395#_M1019_g N_VPWR_c_836_n 0.0134762f $X=7.655 $Y=2.4 $X2=0
+ $Y2=0
cc_440 N_A_840_395#_c_598_n N_VPWR_c_839_n 0.0146088f $X=5.48 $Y=2.265 $X2=0
+ $Y2=0
cc_441 N_A_840_395#_M1012_g N_VPWR_c_840_n 0.00532442f $X=6.23 $Y=2.4 $X2=0
+ $Y2=0
cc_442 N_A_840_395#_M1017_g N_VPWR_c_840_n 0.00460063f $X=6.755 $Y=2.4 $X2=0
+ $Y2=0
cc_443 N_A_840_395#_M1018_g N_VPWR_c_841_n 0.00460063f $X=7.205 $Y=2.4 $X2=0
+ $Y2=0
cc_444 N_A_840_395#_M1019_g N_VPWR_c_841_n 0.00460063f $X=7.655 $Y=2.4 $X2=0
+ $Y2=0
cc_445 N_A_840_395#_M1014_g N_VPWR_c_844_n 0.00529312f $X=4.29 $Y=2.75 $X2=0
+ $Y2=0
cc_446 N_A_840_395#_M1014_g N_VPWR_c_845_n 0.00380629f $X=4.29 $Y=2.75 $X2=0
+ $Y2=0
cc_447 N_A_840_395#_c_595_n N_VPWR_c_845_n 0.0381205f $X=5.315 $Y=2.14 $X2=0
+ $Y2=0
cc_448 N_A_840_395#_c_596_n N_VPWR_c_845_n 0.00854028f $X=4.555 $Y=2.14 $X2=0
+ $Y2=0
cc_449 N_A_840_395#_c_598_n N_VPWR_c_845_n 0.0171801f $X=5.48 $Y=2.265 $X2=0
+ $Y2=0
cc_450 N_A_840_395#_M1014_g N_VPWR_c_830_n 0.0101857f $X=4.29 $Y=2.75 $X2=0
+ $Y2=0
cc_451 N_A_840_395#_M1012_g N_VPWR_c_830_n 0.0104134f $X=6.23 $Y=2.4 $X2=0 $Y2=0
cc_452 N_A_840_395#_M1017_g N_VPWR_c_830_n 0.0090927f $X=6.755 $Y=2.4 $X2=0
+ $Y2=0
cc_453 N_A_840_395#_M1018_g N_VPWR_c_830_n 0.00908554f $X=7.205 $Y=2.4 $X2=0
+ $Y2=0
cc_454 N_A_840_395#_M1019_g N_VPWR_c_830_n 0.00908554f $X=7.655 $Y=2.4 $X2=0
+ $Y2=0
cc_455 N_A_840_395#_c_598_n N_VPWR_c_830_n 0.0120707f $X=5.48 $Y=2.265 $X2=0
+ $Y2=0
cc_456 N_A_840_395#_M1013_g N_Q_c_932_n 0.00944159f $X=6.215 $Y=0.74 $X2=0 $Y2=0
cc_457 N_A_840_395#_M1015_g N_Q_c_932_n 0.00350623f $X=6.735 $Y=0.74 $X2=0 $Y2=0
cc_458 N_A_840_395#_M1012_g N_Q_c_939_n 0.00311328f $X=6.23 $Y=2.4 $X2=0 $Y2=0
cc_459 N_A_840_395#_c_576_n N_Q_c_939_n 0.0038635f $X=6.66 $Y=1.485 $X2=0 $Y2=0
cc_460 N_A_840_395#_c_586_n N_Q_c_939_n 0.0277729f $X=7.325 $Y=1.485 $X2=0 $Y2=0
cc_461 N_A_840_395#_c_598_n N_Q_c_939_n 0.00672843f $X=5.48 $Y=2.265 $X2=0 $Y2=0
cc_462 N_A_840_395#_M1012_g N_Q_c_940_n 0.015337f $X=6.23 $Y=2.4 $X2=0 $Y2=0
cc_463 N_A_840_395#_M1017_g N_Q_c_940_n 4.61969e-19 $X=6.755 $Y=2.4 $X2=0 $Y2=0
cc_464 N_A_840_395#_c_598_n N_Q_c_940_n 0.00428293f $X=5.48 $Y=2.265 $X2=0 $Y2=0
cc_465 N_A_840_395#_M1015_g N_Q_c_933_n 0.0148325f $X=6.735 $Y=0.74 $X2=0 $Y2=0
cc_466 N_A_840_395#_M1023_g N_Q_c_933_n 0.0127898f $X=7.165 $Y=0.74 $X2=0 $Y2=0
cc_467 N_A_840_395#_c_586_n N_Q_c_933_n 0.049875f $X=7.325 $Y=1.485 $X2=0 $Y2=0
cc_468 N_A_840_395#_c_588_n N_Q_c_933_n 0.00237995f $X=7.64 $Y=1.485 $X2=0 $Y2=0
cc_469 N_A_840_395#_M1013_g N_Q_c_934_n 0.00366127f $X=6.215 $Y=0.74 $X2=0 $Y2=0
cc_470 N_A_840_395#_c_576_n N_Q_c_934_n 0.0045445f $X=6.66 $Y=1.485 $X2=0 $Y2=0
cc_471 N_A_840_395#_c_586_n N_Q_c_934_n 0.0293689f $X=7.325 $Y=1.485 $X2=0 $Y2=0
cc_472 N_A_840_395#_c_587_n N_Q_c_934_n 0.00593633f $X=5.745 $Y=1.065 $X2=0
+ $Y2=0
cc_473 N_A_840_395#_M1023_g N_Q_c_935_n 4.44219e-19 $X=7.165 $Y=0.74 $X2=0 $Y2=0
cc_474 N_A_840_395#_M1025_g N_Q_c_935_n 4.74419e-19 $X=7.64 $Y=0.74 $X2=0 $Y2=0
cc_475 N_A_840_395#_M1018_g N_Q_c_941_n 3.8104e-19 $X=7.205 $Y=2.4 $X2=0 $Y2=0
cc_476 N_A_840_395#_M1019_g N_Q_c_941_n 3.8104e-19 $X=7.655 $Y=2.4 $X2=0 $Y2=0
cc_477 N_A_840_395#_M1025_g N_Q_c_936_n 0.0171604f $X=7.64 $Y=0.74 $X2=0 $Y2=0
cc_478 N_A_840_395#_c_588_n N_Q_c_936_n 7.81529e-19 $X=7.64 $Y=1.485 $X2=0 $Y2=0
cc_479 N_A_840_395#_c_586_n N_Q_c_937_n 0.016446f $X=7.325 $Y=1.485 $X2=0 $Y2=0
cc_480 N_A_840_395#_c_588_n N_Q_c_937_n 0.0035948f $X=7.64 $Y=1.485 $X2=0 $Y2=0
cc_481 N_A_840_395#_M1025_g Q 0.0112315f $X=7.64 $Y=0.74 $X2=0 $Y2=0
cc_482 N_A_840_395#_c_586_n Q 0.0168437f $X=7.325 $Y=1.485 $X2=0 $Y2=0
cc_483 N_A_840_395#_c_588_n Q 0.0127563f $X=7.64 $Y=1.485 $X2=0 $Y2=0
cc_484 N_A_840_395#_M1019_g Q 0.0248508f $X=7.655 $Y=2.4 $X2=0 $Y2=0
cc_485 N_A_840_395#_c_588_n Q 0.00205041f $X=7.64 $Y=1.485 $X2=0 $Y2=0
cc_486 N_A_840_395#_M1017_g N_Q_c_944_n 0.0145261f $X=6.755 $Y=2.4 $X2=0 $Y2=0
cc_487 N_A_840_395#_M1018_g N_Q_c_944_n 0.01448f $X=7.205 $Y=2.4 $X2=0 $Y2=0
cc_488 N_A_840_395#_c_586_n N_Q_c_944_n 0.0627487f $X=7.325 $Y=1.485 $X2=0 $Y2=0
cc_489 N_A_840_395#_c_588_n N_Q_c_944_n 0.00211635f $X=7.64 $Y=1.485 $X2=0 $Y2=0
cc_490 N_A_840_395#_M1003_g N_VGND_c_1007_n 0.00349542f $X=4.76 $Y=0.825 $X2=0
+ $Y2=0
cc_491 N_A_840_395#_c_583_n N_VGND_c_1007_n 0.0215088f $X=5.485 $Y=0.54 $X2=0
+ $Y2=0
cc_492 N_A_840_395#_c_587_n N_VGND_c_1007_n 0.00358005f $X=5.745 $Y=1.065 $X2=0
+ $Y2=0
cc_493 N_A_840_395#_M1013_g N_VGND_c_1008_n 0.00739063f $X=6.215 $Y=0.74 $X2=0
+ $Y2=0
cc_494 N_A_840_395#_c_583_n N_VGND_c_1008_n 0.0163189f $X=5.485 $Y=0.54 $X2=0
+ $Y2=0
cc_495 N_A_840_395#_c_586_n N_VGND_c_1008_n 0.00973029f $X=7.325 $Y=1.485 $X2=0
+ $Y2=0
cc_496 N_A_840_395#_c_587_n N_VGND_c_1008_n 0.00182821f $X=5.745 $Y=1.065 $X2=0
+ $Y2=0
cc_497 N_A_840_395#_M1013_g N_VGND_c_1009_n 6.65972e-19 $X=6.215 $Y=0.74 $X2=0
+ $Y2=0
cc_498 N_A_840_395#_M1015_g N_VGND_c_1009_n 0.0099317f $X=6.735 $Y=0.74 $X2=0
+ $Y2=0
cc_499 N_A_840_395#_M1023_g N_VGND_c_1009_n 0.00988667f $X=7.165 $Y=0.74 $X2=0
+ $Y2=0
cc_500 N_A_840_395#_M1025_g N_VGND_c_1009_n 4.5982e-19 $X=7.64 $Y=0.74 $X2=0
+ $Y2=0
cc_501 N_A_840_395#_M1025_g N_VGND_c_1011_n 0.00497413f $X=7.64 $Y=0.74 $X2=0
+ $Y2=0
cc_502 N_A_840_395#_c_583_n N_VGND_c_1012_n 0.00990263f $X=5.485 $Y=0.54 $X2=0
+ $Y2=0
cc_503 N_A_840_395#_M1003_g N_VGND_c_1016_n 0.00399533f $X=4.76 $Y=0.825 $X2=0
+ $Y2=0
cc_504 N_A_840_395#_M1013_g N_VGND_c_1017_n 0.00434272f $X=6.215 $Y=0.74 $X2=0
+ $Y2=0
cc_505 N_A_840_395#_M1015_g N_VGND_c_1017_n 0.00383152f $X=6.735 $Y=0.74 $X2=0
+ $Y2=0
cc_506 N_A_840_395#_M1023_g N_VGND_c_1018_n 0.00383152f $X=7.165 $Y=0.74 $X2=0
+ $Y2=0
cc_507 N_A_840_395#_M1025_g N_VGND_c_1018_n 0.00460063f $X=7.64 $Y=0.74 $X2=0
+ $Y2=0
cc_508 N_A_840_395#_M1003_g N_VGND_c_1023_n 0.00472204f $X=4.76 $Y=0.825 $X2=0
+ $Y2=0
cc_509 N_A_840_395#_M1013_g N_VGND_c_1023_n 0.00826226f $X=6.215 $Y=0.74 $X2=0
+ $Y2=0
cc_510 N_A_840_395#_M1015_g N_VGND_c_1023_n 0.00758371f $X=6.735 $Y=0.74 $X2=0
+ $Y2=0
cc_511 N_A_840_395#_M1023_g N_VGND_c_1023_n 0.00757973f $X=7.165 $Y=0.74 $X2=0
+ $Y2=0
cc_512 N_A_840_395#_M1025_g N_VGND_c_1023_n 0.00911274f $X=7.64 $Y=0.74 $X2=0
+ $Y2=0
cc_513 N_A_840_395#_c_583_n N_VGND_c_1023_n 0.0089622f $X=5.485 $Y=0.54 $X2=0
+ $Y2=0
cc_514 N_A_678_392#_M1022_g N_VPWR_c_833_n 0.00259356f $X=5.725 $Y=2.54 $X2=0
+ $Y2=0
cc_515 N_A_678_392#_M1004_g N_VPWR_c_839_n 0.0050621f $X=5.22 $Y=2.54 $X2=0
+ $Y2=0
cc_516 N_A_678_392#_M1022_g N_VPWR_c_839_n 0.00542159f $X=5.725 $Y=2.54 $X2=0
+ $Y2=0
cc_517 N_A_678_392#_M1004_g N_VPWR_c_845_n 0.010146f $X=5.22 $Y=2.54 $X2=0 $Y2=0
cc_518 N_A_678_392#_M1022_g N_VPWR_c_845_n 4.36892e-19 $X=5.725 $Y=2.54 $X2=0
+ $Y2=0
cc_519 N_A_678_392#_M1004_g N_VPWR_c_830_n 0.00994771f $X=5.22 $Y=2.54 $X2=0
+ $Y2=0
cc_520 N_A_678_392#_M1022_g N_VPWR_c_830_n 0.0105566f $X=5.725 $Y=2.54 $X2=0
+ $Y2=0
cc_521 N_A_678_392#_M1024_g N_Q_c_932_n 9.40157e-19 $X=5.7 $Y=0.715 $X2=0 $Y2=0
cc_522 N_A_678_392#_M1022_g N_Q_c_940_n 6.15093e-19 $X=5.725 $Y=2.54 $X2=0 $Y2=0
cc_523 N_A_678_392#_M1007_g N_VGND_c_1007_n 0.00607982f $X=5.27 $Y=0.715 $X2=0
+ $Y2=0
cc_524 N_A_678_392#_c_729_n N_VGND_c_1007_n 0.0146621f $X=4.55 $Y=0.89 $X2=0
+ $Y2=0
cc_525 N_A_678_392#_c_733_n N_VGND_c_1007_n 0.0160858f $X=5.325 $Y=1.485 $X2=0
+ $Y2=0
cc_526 N_A_678_392#_M1007_g N_VGND_c_1008_n 4.73318e-19 $X=5.27 $Y=0.715 $X2=0
+ $Y2=0
cc_527 N_A_678_392#_M1024_g N_VGND_c_1008_n 0.00930995f $X=5.7 $Y=0.715 $X2=0
+ $Y2=0
cc_528 N_A_678_392#_M1007_g N_VGND_c_1012_n 0.00534051f $X=5.27 $Y=0.715 $X2=0
+ $Y2=0
cc_529 N_A_678_392#_M1024_g N_VGND_c_1012_n 0.00465077f $X=5.7 $Y=0.715 $X2=0
+ $Y2=0
cc_530 N_A_678_392#_c_729_n N_VGND_c_1016_n 0.00333424f $X=4.55 $Y=0.89 $X2=0
+ $Y2=0
cc_531 N_A_678_392#_M1007_g N_VGND_c_1023_n 0.00537853f $X=5.27 $Y=0.715 $X2=0
+ $Y2=0
cc_532 N_A_678_392#_M1024_g N_VGND_c_1023_n 0.00451796f $X=5.7 $Y=0.715 $X2=0
+ $Y2=0
cc_533 N_A_678_392#_c_729_n N_VGND_c_1023_n 0.00882318f $X=4.55 $Y=0.89 $X2=0
+ $Y2=0
cc_534 N_A_678_392#_c_729_n A_895_123# 0.00190356f $X=4.55 $Y=0.89 $X2=-0.19
+ $Y2=-0.245
cc_535 N_VPWR_c_833_n N_Q_c_940_n 0.0615367f $X=5.98 $Y=2.325 $X2=0 $Y2=0
cc_536 N_VPWR_c_834_n N_Q_c_940_n 0.0315588f $X=6.98 $Y=2.265 $X2=0 $Y2=0
cc_537 N_VPWR_c_840_n N_Q_c_940_n 0.0146237f $X=6.815 $Y=3.33 $X2=0 $Y2=0
cc_538 N_VPWR_c_830_n N_Q_c_940_n 0.0120948f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_539 N_VPWR_c_834_n N_Q_c_941_n 0.0315168f $X=6.98 $Y=2.265 $X2=0 $Y2=0
cc_540 N_VPWR_c_836_n N_Q_c_941_n 0.0255132f $X=7.88 $Y=2.405 $X2=0 $Y2=0
cc_541 N_VPWR_c_841_n N_Q_c_941_n 0.0101736f $X=7.715 $Y=3.33 $X2=0 $Y2=0
cc_542 N_VPWR_c_830_n N_Q_c_941_n 0.0084208f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_543 N_VPWR_M1019_s Q 0.00412975f $X=7.745 $Y=1.84 $X2=0 $Y2=0
cc_544 N_VPWR_c_836_n Q 0.0221071f $X=7.88 $Y=2.405 $X2=0 $Y2=0
cc_545 N_VPWR_M1017_s N_Q_c_944_n 0.00165831f $X=6.845 $Y=1.84 $X2=0 $Y2=0
cc_546 N_VPWR_c_834_n N_Q_c_944_n 0.0170259f $X=6.98 $Y=2.265 $X2=0 $Y2=0
cc_547 N_Q_c_933_n N_VGND_M1015_s 0.00176461f $X=7.295 $Y=1.065 $X2=0 $Y2=0
cc_548 N_Q_c_936_n N_VGND_M1025_s 0.00371016f $X=7.805 $Y=1.065 $X2=0 $Y2=0
cc_549 N_Q_c_932_n N_VGND_c_1008_n 0.0336294f $X=6.44 $Y=0.515 $X2=0 $Y2=0
cc_550 N_Q_c_932_n N_VGND_c_1009_n 0.0180579f $X=6.44 $Y=0.515 $X2=0 $Y2=0
cc_551 N_Q_c_933_n N_VGND_c_1009_n 0.0170777f $X=7.295 $Y=1.065 $X2=0 $Y2=0
cc_552 N_Q_c_935_n N_VGND_c_1009_n 0.017215f $X=7.38 $Y=0.515 $X2=0 $Y2=0
cc_553 N_Q_c_935_n N_VGND_c_1011_n 0.0175659f $X=7.38 $Y=0.515 $X2=0 $Y2=0
cc_554 N_Q_c_936_n N_VGND_c_1011_n 0.0234209f $X=7.805 $Y=1.065 $X2=0 $Y2=0
cc_555 N_Q_c_932_n N_VGND_c_1017_n 0.0154563f $X=6.44 $Y=0.515 $X2=0 $Y2=0
cc_556 N_Q_c_935_n N_VGND_c_1018_n 0.011066f $X=7.38 $Y=0.515 $X2=0 $Y2=0
cc_557 N_Q_c_932_n N_VGND_c_1023_n 0.012737f $X=6.44 $Y=0.515 $X2=0 $Y2=0
cc_558 N_Q_c_935_n N_VGND_c_1023_n 0.00915947f $X=7.38 $Y=0.515 $X2=0 $Y2=0

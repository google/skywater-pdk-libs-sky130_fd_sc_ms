* File: sky130_fd_sc_ms__sedfxtp_2.spice
* Created: Wed Sep  2 12:32:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sedfxtp_2.pex.spice"
.subckt sky130_fd_sc_ms__sedfxtp_2  VNB VPB D DE SCD SCE CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCE	SCE
* SCD	SCD
* DE	DE
* D	D
* VPB	VPB
* VNB	VNB
MM1012 A_138_74# N_D_M1012_g N_A_40_464#_M1012_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1039 N_VGND_M1039_d N_DE_M1039_g A_138_74# VNB NLOWVT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_DE_M1021_g N_A_180_290#_M1021_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1023 A_500_113# N_A_180_290#_M1023_g N_VGND_M1021_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1036 N_A_40_464#_M1036_d N_A_548_87#_M1036_g A_500_113# VNB NLOWVT L=0.15
+ W=0.42 AD=0.08925 AS=0.0504 PD=0.845 PS=0.66 NRD=19.992 NRS=18.564 M=1 R=2.8
+ SA=75001 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1037 N_A_693_113#_M1037_d N_A_663_87#_M1037_g N_A_40_464#_M1036_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1491 AS=0.08925 PD=1.55 PS=0.845 NRD=19.992 NRS=21.42 M=1
+ R=2.8 SA=75001.6 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1040 N_VGND_M1040_d N_SCE_M1040_g N_A_663_87#_M1040_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 A_1068_125# N_SCD_M1003_g N_VGND_M1040_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0735 PD=0.63 PS=0.77 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_A_693_113#_M1008_d N_SCE_M1008_g A_1068_125# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_1340_74#_M1004_d N_CLK_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.2183 PD=2.05 PS=2.07 NRD=0 NRS=0.804 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1035 N_A_1538_74#_M1035_d N_A_1340_74#_M1035_g N_VGND_M1035_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1020 N_A_1736_97#_M1020_d N_A_1340_74#_M1020_g N_A_693_113#_M1020_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1197 PD=0.95 PS=1.41 NRD=71.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1027 A_1872_97# N_A_1538_74#_M1027_g N_A_1736_97#_M1020_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.11235 AS=0.1113 PD=0.955 PS=0.95 NRD=60.708 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_A_1979_71#_M1029_g A_1872_97# VNB NLOWVT L=0.15 W=0.42
+ AD=0.139472 AS=0.11235 PD=1.00245 PS=0.955 NRD=25.704 NRS=60.708 M=1 R=2.8
+ SA=75001.6 SB=75001 A=0.063 P=1.14 MULT=1
MM1028 N_A_1979_71#_M1028_d N_A_1736_97#_M1028_g N_VGND_M1029_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.212528 PD=1.85 PS=1.52755 NRD=0 NRS=48.744 M=1
+ R=4.26667 SA=75001.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1043 A_2402_74# N_A_1979_71#_M1043_g N_VGND_M1043_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1824 PD=0.85 PS=1.85 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1001 N_A_2474_74#_M1001_d N_A_1538_74#_M1001_g A_2402_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.115623 AS=0.0672 PD=1.16528 PS=0.85 NRD=8.436 NRS=9.372 M=1
+ R=4.26667 SA=75000.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1031 A_2569_74# N_A_1340_74#_M1031_g N_A_2474_74#_M1001_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0758774 PD=0.66 PS=0.764717 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75001 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1032 N_VGND_M1032_d N_A_548_87#_M1032_g A_2569_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.20055 AS=0.0504 PD=1.375 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1033 N_A_548_87#_M1033_d N_A_2474_74#_M1033_g N_VGND_M1032_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.20055 PD=1.41 PS=1.375 NRD=0 NRS=19.992 M=1 R=2.8
+ SA=75002.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 N_Q_M1017_d N_A_2474_74#_M1017_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.3
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1041 N_Q_M1017_d N_A_2474_74#_M1041_g N_VGND_M1041_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.7
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1018 A_132_464# N_D_M1018_g N_A_40_464#_M1018_s VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.1792 PD=0.88 PS=1.84 NRD=19.9955 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1038 N_VPWR_M1038_d N_A_180_290#_M1038_g A_132_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.1792 AS=0.0768 PD=1.84 PS=0.88 NRD=0 NRS=19.9955 M=1 R=3.55556 SA=90000.6
+ SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1005 N_VPWR_M1005_d N_DE_M1005_g N_A_180_290#_M1005_s VPB PSHORT L=0.18 W=0.64
+ AD=0.16 AS=0.1792 PD=1.14 PS=1.84 NRD=69.2455 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90001.7 A=0.1152 P=1.64 MULT=1
MM1030 A_578_463# N_DE_M1030_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=0.64 AD=0.0672
+ AS=0.16 PD=0.85 PS=1.14 NRD=15.3857 NRS=0 M=1 R=3.55556 SA=90000.9 SB=90001
+ A=0.1152 P=1.64 MULT=1
MM1016 N_A_40_464#_M1016_d N_A_548_87#_M1016_g A_578_463# VPB PSHORT L=0.18
+ W=0.64 AD=0.0864 AS=0.0672 PD=0.91 PS=0.85 NRD=0 NRS=15.3857 M=1 R=3.55556
+ SA=90001.3 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1019 N_A_693_113#_M1019_d N_SCE_M1019_g N_A_40_464#_M1016_d VPB PSHORT L=0.18
+ W=0.64 AD=0.176 AS=0.0864 PD=1.83 PS=0.91 NRD=0 NRS=0 M=1 R=3.55556 SA=90001.7
+ SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1006 N_VPWR_M1006_d N_SCE_M1006_g N_A_663_87#_M1006_s VPB PSHORT L=0.18 W=0.64
+ AD=0.16 AS=0.176 PD=1.14 PS=1.83 NRD=69.2455 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90001.3 A=0.1152 P=1.64 MULT=1
MM1026 A_1082_455# N_SCD_M1026_g N_VPWR_M1006_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.16 PD=0.88 PS=1.14 NRD=19.9955 NRS=0 M=1 R=3.55556 SA=90000.9
+ SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1002 N_A_693_113#_M1002_d N_A_663_87#_M1002_g A_1082_455# VPB PSHORT L=0.18
+ W=0.64 AD=0.1792 AS=0.0768 PD=1.84 PS=0.88 NRD=0 NRS=19.9955 M=1 R=3.55556
+ SA=90001.3 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1034 N_A_1340_74#_M1034_d N_CLK_M1034_g N_VPWR_M1034_s VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.3192 PD=2.8 PS=2.81 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1013 N_A_1538_74#_M1013_d N_A_1340_74#_M1013_g N_VPWR_M1013_s VPB PSHORT
+ L=0.18 W=1.12 AD=0.3136 AS=0.3136 PD=2.8 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1007 N_A_1736_97#_M1007_d N_A_1538_74#_M1007_g N_A_693_113#_M1007_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0567 AS=0.1176 PD=0.69 PS=1.4 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90001.6 A=0.0756 P=1.2 MULT=1
MM1011 A_1939_508# N_A_1340_74#_M1011_g N_A_1736_97#_M1007_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0777 AS=0.0567 PD=0.79 PS=0.69 NRD=60.9715 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1024 N_VPWR_M1024_d N_A_1979_71#_M1024_g A_1939_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.0922833 AS=0.0777 PD=0.883333 PS=0.79 NRD=0 NRS=60.9715 M=1 R=2.33333
+ SA=90001.2 SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1014 N_A_1979_71#_M1014_d N_A_1736_97#_M1014_g N_VPWR_M1024_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2352 AS=0.184567 PD=2.24 PS=1.76667 NRD=0 NRS=19.9167 M=1
+ R=4.66667 SA=90000.7 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1022 A_2360_392# N_A_1979_71#_M1022_g N_VPWR_M1022_s VPB PSHORT L=0.18 W=1
+ AD=0.39 AS=0.29 PD=1.78 PS=2.58 NRD=65.9753 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.8 A=0.18 P=2.36 MULT=1
MM1042 N_A_2474_74#_M1042_d N_A_1340_74#_M1042_g A_2360_392# VPB PSHORT L=0.18
+ W=1 AD=0.208592 AS=0.39 PD=1.91549 PS=1.78 NRD=16.7253 NRS=65.9753 M=1
+ R=5.55556 SA=90001.2 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1000 A_2660_508# N_A_1538_74#_M1000_g N_A_2474_74#_M1042_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0876085 PD=0.66 PS=0.804507 NRD=30.4759 NRS=0 M=1
+ R=2.33333 SA=90001.7 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1015 N_VPWR_M1015_d N_A_548_87#_M1015_g A_2660_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.109992 AS=0.0504 PD=0.92717 PS=0.66 NRD=46.886 NRS=30.4759 M=1 R=2.33333
+ SA=90002.1 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1009 N_A_548_87#_M1009_d N_A_2474_74#_M1009_g N_VPWR_M1015_d VPB PSHORT L=0.18
+ W=0.64 AD=0.1792 AS=0.167608 PD=1.84 PS=1.41283 NRD=0 NRS=46.1571 M=1
+ R=3.55556 SA=90001.9 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1010 N_Q_M1010_d N_A_2474_74#_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1596 AS=0.3136 PD=1.405 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1025 N_Q_M1010_d N_A_2474_74#_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1596 AS=0.3136 PD=1.405 PS=2.8 NRD=0.8668 NRS=0 M=1 R=6.22222 SA=90000.7
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX44_noxref VNB VPB NWDIODE A=31.0841 P=37.16
c_176 VNB 0 3.03176e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__sedfxtp_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__a41o_2.pex.spice
* Created: Wed Sep  2 11:56:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A41O_2%A4 3 5 7 8 15
r27 14 15 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.505 $Y=1.385
+ $X2=0.53 $Y2=1.385
r28 11 14 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.29 $Y=1.385
+ $X2=0.505 $Y2=1.385
r29 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.385 $X2=0.29 $Y2=1.385
r30 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.29 $Y=1.295 $X2=0.29
+ $Y2=1.385
r31 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.22
+ $X2=0.53 $Y2=1.385
r32 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.53 $Y=1.22 $X2=0.53
+ $Y2=0.74
r33 1 14 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.55
+ $X2=0.505 $Y2=1.385
r34 1 3 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=0.505 $Y=1.55
+ $X2=0.505 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__A41O_2%A3 3 6 8 9 10 15 17
c36 6 0 5.73195e-21 $X=1.055 $Y=2.46
r37 15 18 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.01 $Y=1.385
+ $X2=1.01 $Y2=1.55
r38 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.01 $Y=1.385
+ $X2=1.01 $Y2=1.22
r39 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.01
+ $Y=1.385 $X2=1.01 $Y2=1.385
r40 10 16 2.29036 $w=4.68e-07 $l=9e-08 $layer=LI1_cond $X=1.08 $Y=1.295 $X2=1.08
+ $Y2=1.385
r41 9 10 9.41594 $w=4.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.08 $Y=0.925
+ $X2=1.08 $Y2=1.295
r42 8 9 9.41594 $w=4.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.08 $Y=0.555 $X2=1.08
+ $Y2=0.925
r43 6 18 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=1.055 $Y=2.46
+ $X2=1.055 $Y2=1.55
r44 3 17 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.92 $Y=0.74 $X2=0.92
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__A41O_2%A2 3 6 8 9 10 15 17
c36 6 0 1.00085e-19 $X=1.505 $Y=2.46
r37 15 18 39.9775 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.615 $Y=1.385
+ $X2=1.615 $Y2=1.55
r38 15 17 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.615 $Y=1.385
+ $X2=1.615 $Y2=1.22
r39 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.385 $X2=1.65 $Y2=1.385
r40 10 16 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.65 $Y=1.295 $X2=1.65
+ $Y2=1.385
r41 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.65 $Y=0.925
+ $X2=1.65 $Y2=1.295
r42 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.65 $Y=0.555 $X2=1.65
+ $Y2=0.925
r43 6 18 353.726 $w=1.8e-07 $l=9.1e-07 $layer=POLY_cond $X=1.505 $Y=2.46
+ $X2=1.505 $Y2=1.55
r44 3 17 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.49 $Y=0.74 $X2=1.49
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__A41O_2%A1 3 7 9 12
r40 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.19 $Y=1.615
+ $X2=2.19 $Y2=1.78
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.19 $Y=1.615
+ $X2=2.19 $Y2=1.45
r42 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.19
+ $Y=1.615 $X2=2.19 $Y2=1.615
r43 7 15 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=2.235 $Y=2.46
+ $X2=2.235 $Y2=1.78
r44 3 14 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.13 $Y=0.74 $X2=2.13
+ $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_MS__A41O_2%B1 3 7 9 12 13
c37 13 0 1.06575e-19 $X=2.76 $Y=1.615
r38 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.76 $Y=1.615
+ $X2=2.76 $Y2=1.78
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.76 $Y=1.615
+ $X2=2.76 $Y2=1.45
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.76
+ $Y=1.615 $X2=2.76 $Y2=1.615
r41 9 13 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.64 $Y=1.615 $X2=2.76
+ $Y2=1.615
r42 7 15 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=2.685 $Y=2.46
+ $X2=2.685 $Y2=1.78
r43 3 14 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.67 $Y=0.74 $X2=2.67
+ $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_MS__A41O_2%A_441_74# 1 2 7 9 12 14 16 19 21 22 25 29 31
+ 32 35 41 45 46 48
c84 21 0 1.06575e-19 $X=3.325 $Y=1.385
c85 14 0 1.91222e-19 $X=3.81 $Y=1.22
r86 45 47 1.20266 $w=4.68e-07 $l=5e-09 $layer=LI1_cond $X=3.03 $Y=2.115 $X2=3.03
+ $Y2=2.12
r87 45 46 9.33757 $w=4.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.03 $Y=2.115
+ $X2=3.03 $Y2=1.95
r88 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.68
+ $Y=1.385 $X2=3.68 $Y2=1.385
r89 39 48 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.265 $Y=1.33
+ $X2=3.18 $Y2=1.33
r90 39 41 10.8696 $w=4.38e-07 $l=4.15e-07 $layer=LI1_cond $X=3.265 $Y=1.33
+ $X2=3.68 $Y2=1.33
r91 37 48 3.51065 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=3.18 $Y=1.55 $X2=3.18
+ $Y2=1.33
r92 37 46 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.18 $Y=1.55 $X2=3.18
+ $Y2=1.95
r93 35 47 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.96 $Y=2.815
+ $X2=2.96 $Y2=2.12
r94 31 48 3.10218 $w=3.05e-07 $l=1.72337e-07 $layer=LI1_cond $X=3.095 $Y=1.195
+ $X2=3.18 $Y2=1.33
r95 31 32 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.095 $Y=1.195
+ $X2=2.56 $Y2=1.195
r96 27 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.395 $Y=1.11
+ $X2=2.56 $Y2=1.195
r97 27 29 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=2.395 $Y=1.11
+ $X2=2.395 $Y2=0.515
r98 24 25 76.0647 $w=3.3e-07 $l=4.35e-07 $layer=POLY_cond $X=3.81 $Y=1.385
+ $X2=4.245 $Y2=1.385
r99 23 24 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.795 $Y=1.385
+ $X2=3.81 $Y2=1.385
r100 22 42 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=3.705 $Y=1.385
+ $X2=3.68 $Y2=1.385
r101 22 23 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.705 $Y=1.385
+ $X2=3.795 $Y2=1.385
r102 21 42 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=3.325 $Y=1.385
+ $X2=3.68 $Y2=1.385
r103 17 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.245 $Y=1.55
+ $X2=4.245 $Y2=1.385
r104 17 19 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=4.245 $Y=1.55
+ $X2=4.245 $Y2=2.4
r105 14 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.81 $Y=1.22
+ $X2=3.81 $Y2=1.385
r106 14 16 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.81 $Y=1.22
+ $X2=3.81 $Y2=0.74
r107 10 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.795 $Y=1.55
+ $X2=3.795 $Y2=1.385
r108 10 12 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.795 $Y=1.55
+ $X2=3.795 $Y2=2.4
r109 7 21 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.25 $Y=1.22
+ $X2=3.325 $Y2=1.385
r110 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.25 $Y=1.22 $X2=3.25
+ $Y2=0.74
r111 2 45 400 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.96 $X2=2.96 $Y2=2.115
r112 2 35 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=2.775
+ $Y=1.96 $X2=2.96 $Y2=2.815
r113 1 29 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=2.205
+ $Y=0.37 $X2=2.395 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A41O_2%A_27_392# 1 2 3 12 16 17 20 22 24 26 28
c57 22 0 5.73195e-21 $X=2.295 $Y=2.035
c58 16 0 1.00085e-19 $X=1.115 $Y=1.805
r59 30 32 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=1.28 $Y=2.035 $X2=1.28
+ $Y2=2.105
r60 28 30 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.28 $Y=1.805
+ $X2=1.28 $Y2=2.035
r61 24 34 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.46 $Y=2.12 $X2=2.46
+ $Y2=2.035
r62 24 26 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.46 $Y=2.12
+ $X2=2.46 $Y2=2.815
r63 23 30 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=2.035
+ $X2=1.28 $Y2=2.035
r64 22 34 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=2.035
+ $X2=2.46 $Y2=2.035
r65 22 23 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=2.295 $Y=2.035
+ $X2=1.445 $Y2=2.035
r66 18 32 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.28 $Y=2.12
+ $X2=1.28 $Y2=2.105
r67 18 20 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.28 $Y=2.12
+ $X2=1.28 $Y2=2.815
r68 16 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=1.805
+ $X2=1.28 $Y2=1.805
r69 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=1.805
+ $X2=0.445 $Y2=1.805
r70 12 14 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.28 $Y=2.105
+ $X2=0.28 $Y2=2.815
r71 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.89
+ $X2=0.445 $Y2=1.805
r72 10 12 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=0.28 $Y=1.89
+ $X2=0.28 $Y2=2.105
r73 3 34 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.96 $X2=2.46 $Y2=2.115
r74 3 26 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.96 $X2=2.46 $Y2=2.815
r75 2 32 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.96 $X2=1.28 $Y2=2.105
r76 2 20 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.96 $X2=1.28 $Y2=2.815
r77 1 14 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r78 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_MS__A41O_2%VPWR 1 2 3 4 15 19 23 27 29 31 35 37 42 50 56
+ 59 62 66
r55 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r56 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r57 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 57 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r59 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 54 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r61 54 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r62 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r63 51 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=3.33
+ $X2=3.52 $Y2=3.33
r64 51 53 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.685 $Y=3.33
+ $X2=4.08 $Y2=3.33
r65 50 65 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=4.355 $Y=3.33
+ $X2=4.577 $Y2=3.33
r66 50 53 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.355 $Y=3.33
+ $X2=4.08 $Y2=3.33
r67 49 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r68 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r69 46 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 45 48 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r71 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r72 43 59 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=2.125 $Y=3.33
+ $X2=1.87 $Y2=3.33
r73 43 45 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.125 $Y=3.33
+ $X2=2.16 $Y2=3.33
r74 42 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.355 $Y=3.33
+ $X2=3.52 $Y2=3.33
r75 42 48 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.355 $Y=3.33
+ $X2=3.12 $Y2=3.33
r76 40 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r77 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r78 37 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r79 37 39 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r80 35 49 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=3.12 $Y2=3.33
r81 35 46 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r82 31 34 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.52 $Y=1.985
+ $X2=4.52 $Y2=2.815
r83 29 65 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.52 $Y=3.245
+ $X2=4.577 $Y2=3.33
r84 29 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.52 $Y=3.245
+ $X2=4.52 $Y2=2.815
r85 25 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.52 $Y=3.245
+ $X2=3.52 $Y2=3.33
r86 25 27 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=3.52 $Y=3.245
+ $X2=3.52 $Y2=2.38
r87 21 59 2.12513 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.87 $Y=3.245
+ $X2=1.87 $Y2=3.33
r88 21 23 20.4037 $w=5.08e-07 $l=8.7e-07 $layer=LI1_cond $X=1.87 $Y=3.245
+ $X2=1.87 $Y2=2.375
r89 20 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r90 19 59 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.615 $Y=3.33
+ $X2=1.87 $Y2=3.33
r91 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.615 $Y=3.33
+ $X2=0.945 $Y2=3.33
r92 15 18 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.78 $Y=2.145
+ $X2=0.78 $Y2=2.825
r93 13 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r94 13 18 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.825
r95 4 34 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=4.335
+ $Y=1.84 $X2=4.52 $Y2=2.815
r96 4 31 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=4.335
+ $Y=1.84 $X2=4.52 $Y2=1.985
r97 3 27 300 $w=1.7e-07 $l=6.08194e-07 $layer=licon1_PDIFF $count=2 $X=3.375
+ $Y=1.84 $X2=3.52 $Y2=2.38
r98 2 23 300 $w=1.7e-07 $l=5.35117e-07 $layer=licon1_PDIFF $count=2 $X=1.595
+ $Y=1.96 $X2=1.87 $Y2=2.375
r99 1 18 400 $w=1.7e-07 $l=9.53021e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.96 $X2=0.78 $Y2=2.825
r100 1 15 400 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.96 $X2=0.78 $Y2=2.145
.ends

.subckt PM_SKY130_FD_SC_MS__A41O_2%X 1 2 7 11 13 17 20 21
c36 21 0 1.91222e-19 $X=3.6 $Y=0.555
r37 17 21 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.55 $Y=0.77
+ $X2=3.55 $Y2=0.495
r38 17 19 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=0.77 $X2=3.55
+ $Y2=0.855
r39 15 20 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=4.1 $Y=0.94 $X2=4.1
+ $Y2=1.82
r40 11 20 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.02 $Y=1.985
+ $X2=4.02 $Y2=1.82
r41 11 13 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=4.02 $Y=1.985
+ $X2=4.02 $Y2=2.815
r42 8 19 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.715 $Y=0.855
+ $X2=3.55 $Y2=0.855
r43 7 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.015 $Y=0.855
+ $X2=4.1 $Y2=0.94
r44 7 8 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.015 $Y=0.855 $X2=3.715
+ $Y2=0.855
r45 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.885
+ $Y=1.84 $X2=4.02 $Y2=2.815
r46 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.885
+ $Y=1.84 $X2=4.02 $Y2=1.985
r47 1 21 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=3.325
+ $Y=0.37 $X2=3.55 $Y2=0.495
r48 1 19 182 $w=1.7e-07 $l=5.86813e-07 $layer=licon1_NDIFF $count=1 $X=3.325
+ $Y=0.37 $X2=3.55 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_MS__A41O_2%VGND 1 2 3 10 12 16 19 20 21 30 41 44
r50 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r51 41 43 0.787097 $w=6.2e-07 $l=4e-08 $layer=LI1_cond $X=4.52 $Y=0.257 $X2=4.56
+ $Y2=0.257
r52 39 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r53 38 41 8.65806 $w=6.2e-07 $l=4.4e-07 $layer=LI1_cond $X=4.08 $Y=0.257
+ $X2=4.52 $Y2=0.257
r54 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r55 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r56 33 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r57 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r58 30 38 11.0826 $w=6.2e-07 $l=3.40828e-07 $layer=LI1_cond $X=3.885 $Y=0
+ $X2=4.08 $Y2=0.257
r59 30 32 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.885 $Y=0 $X2=3.6
+ $Y2=0
r60 29 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r61 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r62 26 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r63 25 28 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.64
+ $Y2=0
r64 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r65 23 35 4.65971 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=0.48 $Y=0 $X2=0.24
+ $Y2=0
r66 23 25 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.48 $Y=0 $X2=0.72
+ $Y2=0
r67 21 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r68 21 26 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=0.72
+ $Y2=0
r69 19 28 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.79 $Y=0 $X2=2.64
+ $Y2=0
r70 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.79 $Y=0 $X2=2.955
+ $Y2=0
r71 18 32 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r72 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=2.955
+ $Y2=0
r73 14 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.955 $Y=0.085
+ $X2=2.955 $Y2=0
r74 14 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.955 $Y=0.085
+ $X2=2.955 $Y2=0.515
r75 10 35 3.10647 $w=3.3e-07 $l=1.16619e-07 $layer=LI1_cond $X=0.315 $Y=0.085
+ $X2=0.24 $Y2=0
r76 10 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.315 $Y=0.085
+ $X2=0.315 $Y2=0.515
r77 3 41 91 $w=1.7e-07 $l=7.03776e-07 $layer=licon1_NDIFF $count=2 $X=3.885
+ $Y=0.37 $X2=4.52 $Y2=0.515
r78 2 16 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=2.745
+ $Y=0.37 $X2=2.955 $Y2=0.515
r79 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.17
+ $Y=0.37 $X2=0.315 $Y2=0.515
.ends


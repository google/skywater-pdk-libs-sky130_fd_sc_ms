* File: sky130_fd_sc_ms__buf_1.pex.spice
* Created: Fri Aug 28 17:15:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__BUF_1%A 3 7 9 10 11 12
c37 10 0 7.3311e-20 $X=0.77 $Y=1.45
c38 3 0 1.25263e-20 $X=0.845 $Y=0.835
r39 12 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.745
+ $Y=1.615 $X2=0.745 $Y2=1.615
r40 11 12 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.72 $Y2=1.615
r41 9 16 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.77 $Y=1.615
+ $X2=0.745 $Y2=1.615
r42 9 10 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.77 $Y=1.615
+ $X2=0.77 $Y2=1.45
r43 5 10 34.7346 $w=1.65e-07 $l=5.53173e-07 $layer=POLY_cond $X=0.86 $Y=1.96
+ $X2=0.77 $Y2=1.45
r44 5 7 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=0.86 $Y=1.96 $X2=0.86
+ $Y2=2.54
r45 1 10 34.7346 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=0.845 $Y=1.45
+ $X2=0.77 $Y2=1.45
r46 1 3 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=0.845 $Y=1.45
+ $X2=0.845 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__BUF_1%A_27_164# 1 2 9 13 17 19 21 22 23 24 30 34
r62 34 37 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.465
+ $X2=1.33 $Y2=1.63
r63 34 36 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.33 $Y=1.465
+ $X2=1.33 $Y2=1.3
r64 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.465 $X2=1.325 $Y2=1.465
r65 29 30 9.39634 $w=4.78e-07 $l=1.65e-07 $layer=LI1_cond $X=0.63 $Y=1.04
+ $X2=0.795 $Y2=1.04
r66 26 29 8.72141 $w=4.78e-07 $l=3.5e-07 $layer=LI1_cond $X=0.28 $Y=1.04
+ $X2=0.63 $Y2=1.04
r67 23 33 9.01297 $w=2.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=1.215 $Y=1.63
+ $X2=1.31 $Y2=1.465
r68 23 24 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.215 $Y=1.63
+ $X2=1.215 $Y2=1.95
r69 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.13 $Y=2.035
+ $X2=1.215 $Y2=1.95
r70 21 22 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.13 $Y=2.035
+ $X2=0.8 $Y2=2.035
r71 19 33 11.3586 $w=2.9e-07 $l=3.48569e-07 $layer=LI1_cond $X=1.13 $Y=1.195
+ $X2=1.31 $Y2=1.465
r72 19 30 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.13 $Y=1.195
+ $X2=0.795 $Y2=1.195
r73 15 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.635 $Y=2.12
+ $X2=0.8 $Y2=2.035
r74 15 17 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.635 $Y=2.12
+ $X2=0.635 $Y2=2.265
r75 13 36 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.425 $Y=0.74
+ $X2=1.425 $Y2=1.3
r76 9 37 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.41 $Y=2.4 $X2=1.41
+ $Y2=1.63
r77 2 17 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.49
+ $Y=2.12 $X2=0.635 $Y2=2.265
r78 1 29 182 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.82 $X2=0.63 $Y2=0.965
r79 1 26 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.82 $X2=0.28 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_MS__BUF_1%VPWR 1 6 8 10 17 18 21
r22 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r23 18 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r24 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r25 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.3 $Y=3.33
+ $X2=1.135 $Y2=3.33
r26 15 17 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.3 $Y=3.33 $X2=1.68
+ $Y2=3.33
r27 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r28 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=1.135 $Y2=3.33
r29 10 12 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=0.72 $Y2=3.33
r30 8 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.2 $Y2=3.33
r31 8 13 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r32 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=3.245
+ $X2=1.135 $Y2=3.33
r33 4 6 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.135 $Y=3.245
+ $X2=1.135 $Y2=2.455
r34 1 6 300 $w=1.7e-07 $l=4.17373e-07 $layer=licon1_PDIFF $count=2 $X=0.95
+ $Y=2.12 $X2=1.135 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__BUF_1%X 1 2 9 13 14 15 16 23 32
c25 14 0 7.3311e-20 $X=1.595 $Y=1.95
c26 13 0 1.25263e-20 $X=1.652 $Y=1.13
r27 21 23 1.12043 $w=3.58e-07 $l=3.5e-08 $layer=LI1_cond $X=1.65 $Y=2 $X2=1.65
+ $Y2=2.035
r28 15 16 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.65 $Y=2.405
+ $X2=1.65 $Y2=2.775
r29 14 21 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=1.65 $Y=1.975
+ $X2=1.65 $Y2=2
r30 14 32 8.1909 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=1.65 $Y=1.975
+ $X2=1.65 $Y2=1.82
r31 14 15 11.0442 $w=3.58e-07 $l=3.45e-07 $layer=LI1_cond $X=1.65 $Y=2.06
+ $X2=1.65 $Y2=2.405
r32 14 23 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=1.65 $Y=2.06
+ $X2=1.65 $Y2=2.035
r33 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.745 $Y=1.13
+ $X2=1.745 $Y2=1.82
r34 7 13 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=1.652 $Y=0.953
+ $X2=1.652 $Y2=1.13
r35 7 9 14.2189 $w=3.53e-07 $l=4.38e-07 $layer=LI1_cond $X=1.652 $Y=0.953
+ $X2=1.652 $Y2=0.515
r36 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.84 $X2=1.635 $Y2=1.985
r37 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.84 $X2=1.635 $Y2=2.815
r38 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.5 $Y=0.37
+ $X2=1.64 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__BUF_1%VGND 1 6 8 10 17 18 21
r19 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r20 18 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r21 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r22 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.14
+ $Y2=0
r23 15 17 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.68
+ $Y2=0
r24 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r25 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.14
+ $Y2=0
r26 10 12 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=0.72
+ $Y2=0
r27 8 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r28 8 13 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r29 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.085 $X2=1.14
+ $Y2=0
r30 4 6 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.14 $Y=0.085 $X2=1.14
+ $Y2=0.515
r31 1 6 91 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=2 $X=0.92
+ $Y=0.56 $X2=1.14 $Y2=0.515
.ends


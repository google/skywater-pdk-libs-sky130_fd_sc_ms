* File: sky130_fd_sc_ms__xor3_1.pxi.spice
* Created: Wed Sep  2 12:34:19 2020
* 
x_PM_SKY130_FD_SC_MS__XOR3_1%A_84_108# N_A_84_108#_M1000_d N_A_84_108#_M1020_d
+ N_A_84_108#_M1002_d N_A_84_108#_M1010_d N_A_84_108#_M1019_g
+ N_A_84_108#_M1005_g N_A_84_108#_c_189_n N_A_84_108#_c_190_n
+ N_A_84_108#_c_197_n N_A_84_108#_c_198_n N_A_84_108#_c_199_n
+ N_A_84_108#_c_191_n N_A_84_108#_c_201_n N_A_84_108#_c_202_n
+ N_A_84_108#_c_203_n N_A_84_108#_c_204_n N_A_84_108#_c_205_n
+ N_A_84_108#_c_192_n N_A_84_108#_c_193_n PM_SKY130_FD_SC_MS__XOR3_1%A_84_108#
x_PM_SKY130_FD_SC_MS__XOR3_1%A N_A_M1002_g N_A_c_302_n N_A_M1000_g A N_A_c_304_n
+ PM_SKY130_FD_SC_MS__XOR3_1%A
x_PM_SKY130_FD_SC_MS__XOR3_1%A_452_288# N_A_452_288#_M1011_s
+ N_A_452_288#_M1021_s N_A_452_288#_M1008_g N_A_452_288#_M1006_g
+ N_A_452_288#_c_340_n N_A_452_288#_c_341_n N_A_452_288#_M1010_g
+ N_A_452_288#_M1020_g N_A_452_288#_c_344_n N_A_452_288#_c_345_n
+ N_A_452_288#_c_346_n N_A_452_288#_c_347_n N_A_452_288#_c_348_n
+ N_A_452_288#_c_349_n N_A_452_288#_c_350_n N_A_452_288#_c_351_n
+ N_A_452_288#_c_352_n N_A_452_288#_c_353_n
+ PM_SKY130_FD_SC_MS__XOR3_1%A_452_288#
x_PM_SKY130_FD_SC_MS__XOR3_1%B N_B_M1012_g N_B_M1015_g N_B_c_461_n N_B_c_462_n
+ N_B_c_448_n N_B_c_449_n N_B_M1009_g N_B_c_464_n N_B_M1014_g N_B_c_451_n
+ N_B_c_452_n N_B_c_453_n N_B_M1021_g N_B_M1011_g N_B_c_467_n N_B_c_455_n
+ N_B_c_456_n B N_B_c_457_n N_B_c_458_n N_B_c_459_n PM_SKY130_FD_SC_MS__XOR3_1%B
x_PM_SKY130_FD_SC_MS__XOR3_1%A_1157_298# N_A_1157_298#_M1017_s
+ N_A_1157_298#_M1013_s N_A_1157_298#_M1001_g N_A_1157_298#_M1016_g
+ N_A_1157_298#_c_589_n N_A_1157_298#_c_590_n N_A_1157_298#_c_591_n
+ N_A_1157_298#_c_592_n N_A_1157_298#_c_584_n N_A_1157_298#_c_585_n
+ N_A_1157_298#_c_604_p N_A_1157_298#_c_594_n N_A_1157_298#_c_586_n
+ N_A_1157_298#_c_587_n PM_SKY130_FD_SC_MS__XOR3_1%A_1157_298#
x_PM_SKY130_FD_SC_MS__XOR3_1%C N_C_M1003_g N_C_c_674_n N_C_M1007_g N_C_c_675_n
+ N_C_c_676_n N_C_c_677_n N_C_M1013_g N_C_c_679_n N_C_M1017_g N_C_c_680_n
+ N_C_c_681_n C PM_SKY130_FD_SC_MS__XOR3_1%C
x_PM_SKY130_FD_SC_MS__XOR3_1%A_1218_396# N_A_1218_396#_M1016_d
+ N_A_1218_396#_M1001_d N_A_1218_396#_M1004_g N_A_1218_396#_M1018_g
+ N_A_1218_396#_c_770_n N_A_1218_396#_c_762_n N_A_1218_396#_c_763_n
+ N_A_1218_396#_c_764_n N_A_1218_396#_c_765_n N_A_1218_396#_c_766_n
+ N_A_1218_396#_c_767_n N_A_1218_396#_c_768_n
+ PM_SKY130_FD_SC_MS__XOR3_1%A_1218_396#
x_PM_SKY130_FD_SC_MS__XOR3_1%A_27_134# N_A_27_134#_M1019_s N_A_27_134#_M1006_d
+ N_A_27_134#_M1005_s N_A_27_134#_M1008_d N_A_27_134#_c_847_n
+ N_A_27_134#_c_848_n N_A_27_134#_c_849_n N_A_27_134#_c_850_n
+ N_A_27_134#_c_851_n N_A_27_134#_c_852_n N_A_27_134#_c_853_n
+ N_A_27_134#_c_854_n N_A_27_134#_c_855_n N_A_27_134#_c_856_n
+ N_A_27_134#_c_861_n N_A_27_134#_c_857_n N_A_27_134#_c_858_n
+ N_A_27_134#_c_859_n PM_SKY130_FD_SC_MS__XOR3_1%A_27_134#
x_PM_SKY130_FD_SC_MS__XOR3_1%VPWR N_VPWR_M1005_d N_VPWR_M1021_d N_VPWR_M1013_d
+ N_VPWR_c_933_n N_VPWR_c_934_n N_VPWR_c_935_n N_VPWR_c_936_n N_VPWR_c_937_n
+ VPWR N_VPWR_c_938_n N_VPWR_c_939_n N_VPWR_c_940_n N_VPWR_c_932_n
+ N_VPWR_c_942_n N_VPWR_c_943_n PM_SKY130_FD_SC_MS__XOR3_1%VPWR
x_PM_SKY130_FD_SC_MS__XOR3_1%A_387_392# N_A_387_392#_M1014_d
+ N_A_387_392#_M1016_s N_A_387_392#_M1012_d N_A_387_392#_M1003_d
+ N_A_387_392#_c_1016_n N_A_387_392#_c_1017_n N_A_387_392#_c_1018_n
+ N_A_387_392#_c_1008_n N_A_387_392#_c_1009_n N_A_387_392#_c_1010_n
+ N_A_387_392#_c_1057_n N_A_387_392#_c_1011_n N_A_387_392#_c_1061_n
+ N_A_387_392#_c_1012_n N_A_387_392#_c_1013_n N_A_387_392#_c_1014_n
+ N_A_387_392#_c_1020_n N_A_387_392#_c_1021_n N_A_387_392#_c_1022_n
+ N_A_387_392#_c_1015_n PM_SKY130_FD_SC_MS__XOR3_1%A_387_392#
x_PM_SKY130_FD_SC_MS__XOR3_1%A_416_86# N_A_416_86#_M1015_d N_A_416_86#_M1007_d
+ N_A_416_86#_M1009_d N_A_416_86#_M1001_s N_A_416_86#_c_1135_n
+ N_A_416_86#_c_1136_n N_A_416_86#_c_1137_n N_A_416_86#_c_1148_n
+ N_A_416_86#_c_1246_n N_A_416_86#_c_1138_n N_A_416_86#_c_1139_n
+ N_A_416_86#_c_1200_n N_A_416_86#_c_1140_n N_A_416_86#_c_1149_n
+ N_A_416_86#_c_1141_n N_A_416_86#_c_1142_n N_A_416_86#_c_1143_n
+ N_A_416_86#_c_1144_n N_A_416_86#_c_1145_n N_A_416_86#_c_1146_n
+ N_A_416_86#_c_1147_n PM_SKY130_FD_SC_MS__XOR3_1%A_416_86#
x_PM_SKY130_FD_SC_MS__XOR3_1%X N_X_M1018_d N_X_M1004_d X X X X X X X
+ PM_SKY130_FD_SC_MS__XOR3_1%X
x_PM_SKY130_FD_SC_MS__XOR3_1%VGND N_VGND_M1019_d N_VGND_M1011_d N_VGND_M1017_d
+ N_VGND_c_1276_n N_VGND_c_1277_n VGND N_VGND_c_1278_n N_VGND_c_1279_n
+ N_VGND_c_1280_n N_VGND_c_1281_n N_VGND_c_1282_n N_VGND_c_1283_n
+ N_VGND_c_1284_n N_VGND_c_1285_n PM_SKY130_FD_SC_MS__XOR3_1%VGND
cc_1 VNB N_A_84_108#_M1019_g 0.0280523f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.99
cc_2 VNB N_A_84_108#_c_189_n 0.00302548f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.635
cc_3 VNB N_A_84_108#_c_190_n 0.0194956f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.635
cc_4 VNB N_A_84_108#_c_191_n 0.00870462f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.165
cc_5 VNB N_A_84_108#_c_192_n 0.00280308f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=1.905
cc_6 VNB N_A_84_108#_c_193_n 8.32769e-19 $X=-0.19 $Y=-0.245 $X2=4.31 $Y2=1.1
cc_7 VNB N_A_c_302_n 0.0208818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB A 0.00138047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_c_304_n 0.0295388f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.99
cc_10 VNB N_A_452_288#_M1008_g 0.0054618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_452_288#_M1006_g 0.0364361f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.47
cc_12 VNB N_A_452_288#_c_340_n 0.0448275f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.99
cc_13 VNB N_A_452_288#_c_341_n 0.0161727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_452_288#_M1010_g 0.00432669f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.46
cc_15 VNB N_A_452_288#_M1020_g 0.0192074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_452_288#_c_344_n 0.0112372f $X=-0.19 $Y=-0.245 $X2=1.535 $Y2=2.105
cc_17 VNB N_A_452_288#_c_345_n 0.00121722f $X=-0.19 $Y=-0.245 $X2=1.535
+ $Y2=2.815
cc_18 VNB N_A_452_288#_c_346_n 0.00662046f $X=-0.19 $Y=-0.245 $X2=1.535
+ $Y2=2.815
cc_19 VNB N_A_452_288#_c_347_n 3.26207e-19 $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.92
cc_20 VNB N_A_452_288#_c_348_n 0.00209964f $X=-0.19 $Y=-0.245 $X2=3.725 $Y2=2.99
cc_21 VNB N_A_452_288#_c_349_n 0.00521677f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=2.905
cc_22 VNB N_A_452_288#_c_350_n 0.00121966f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=2.755
cc_23 VNB N_A_452_288#_c_351_n 0.0215802f $X=-0.19 $Y=-0.245 $X2=4.15 $Y2=1.1
cc_24 VNB N_A_452_288#_c_352_n 0.00171652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_452_288#_c_353_n 0.0171849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B_M1015_g 0.0269244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B_c_448_n 0.0680104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B_c_449_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B_M1014_g 0.021965f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.92
cc_30 VNB N_B_c_451_n 0.089017f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.635
cc_31 VNB N_B_c_452_n 0.00731819f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=2.005
cc_32 VNB N_B_c_453_n 0.0651912f $X=-0.19 $Y=-0.245 $X2=1.535 $Y2=2.09
cc_33 VNB N_B_M1011_g 0.0294207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_B_c_455_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=2.755
cc_35 VNB N_B_c_456_n 0.00741352f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=2.905
cc_36 VNB N_B_c_457_n 0.0148671f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=2.07
cc_37 VNB N_B_c_458_n 0.0325472f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=2.755
cc_38 VNB N_B_c_459_n 0.00289172f $X=-0.19 $Y=-0.245 $X2=4.15 $Y2=1.1
cc_39 VNB N_A_1157_298#_M1016_g 0.0284968f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.47
cc_40 VNB N_A_1157_298#_c_584_n 0.00230372f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=1.635
cc_41 VNB N_A_1157_298#_c_585_n 0.00579654f $X=-0.19 $Y=-0.245 $X2=1.37
+ $Y2=2.005
cc_42 VNB N_A_1157_298#_c_586_n 7.49477e-19 $X=-0.19 $Y=-0.245 $X2=1.7 $Y2=2.99
cc_43 VNB N_A_1157_298#_c_587_n 0.024308f $X=-0.19 $Y=-0.245 $X2=4.31 $Y2=1.905
cc_44 VNB N_C_c_674_n 0.020737f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_C_c_675_n 0.0482695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_C_c_676_n 0.0369866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_C_c_677_n 0.0207623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_C_M1013_g 0.00345753f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.99
cc_49 VNB N_C_c_679_n 0.0167509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_C_c_680_n 0.0265346f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.92
cc_51 VNB N_C_c_681_n 0.0113569f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.635
cc_52 VNB C 9.91118e-19 $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.635
cc_53 VNB N_A_1218_396#_M1018_g 0.0259845f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.47
cc_54 VNB N_A_1218_396#_c_762_n 0.00504306f $X=-0.19 $Y=-0.245 $X2=0.587
+ $Y2=1.92
cc_55 VNB N_A_1218_396#_c_763_n 0.0111402f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=1.635
cc_56 VNB N_A_1218_396#_c_764_n 0.00732547f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=1.635
cc_57 VNB N_A_1218_396#_c_765_n 0.00301031f $X=-0.19 $Y=-0.245 $X2=0.75
+ $Y2=2.005
cc_58 VNB N_A_1218_396#_c_766_n 3.72864e-19 $X=-0.19 $Y=-0.245 $X2=1.535
+ $Y2=2.105
cc_59 VNB N_A_1218_396#_c_767_n 0.00273385f $X=-0.19 $Y=-0.245 $X2=1.54
+ $Y2=1.165
cc_60 VNB N_A_1218_396#_c_768_n 0.0358854f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.165
cc_61 VNB N_A_27_134#_c_847_n 0.0122281f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.47
cc_62 VNB N_A_27_134#_c_848_n 0.0113703f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.99
cc_63 VNB N_A_27_134#_c_849_n 0.00553396f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.8
cc_64 VNB N_A_27_134#_c_850_n 0.00189123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_27_134#_c_851_n 0.0135701f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.92
cc_66 VNB N_A_27_134#_c_852_n 0.00382875f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.635
cc_67 VNB N_A_27_134#_c_853_n 5.75772e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_27_134#_c_854_n 5.55082e-19 $X=-0.19 $Y=-0.245 $X2=1.535 $Y2=2.905
cc_69 VNB N_A_27_134#_c_855_n 0.0028476f $X=-0.19 $Y=-0.245 $X2=1.535 $Y2=2.815
cc_70 VNB N_A_27_134#_c_856_n 0.00710642f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.165
cc_71 VNB N_A_27_134#_c_857_n 0.0169882f $X=-0.19 $Y=-0.245 $X2=3.725 $Y2=2.99
cc_72 VNB N_A_27_134#_c_858_n 0.00227978f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=2.755
cc_73 VNB N_A_27_134#_c_859_n 0.0014917f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=2.905
cc_74 VNB N_VPWR_c_932_n 0.382608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_387_392#_c_1008_n 0.00288672f $X=-0.19 $Y=-0.245 $X2=0.587
+ $Y2=1.635
cc_76 VNB N_A_387_392#_c_1009_n 0.0231598f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=1.635
cc_77 VNB N_A_387_392#_c_1010_n 0.00220727f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=1.635
cc_78 VNB N_A_387_392#_c_1011_n 0.00792656f $X=-0.19 $Y=-0.245 $X2=0.75
+ $Y2=2.005
cc_79 VNB N_A_387_392#_c_1012_n 0.00980532f $X=-0.19 $Y=-0.245 $X2=1.535
+ $Y2=2.815
cc_80 VNB N_A_387_392#_c_1013_n 0.0415815f $X=-0.19 $Y=-0.245 $X2=1.535
+ $Y2=2.815
cc_81 VNB N_A_387_392#_c_1014_n 0.0051092f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.92
cc_82 VNB N_A_387_392#_c_1015_n 0.0231253f $X=-0.19 $Y=-0.245 $X2=4.31 $Y2=1.265
cc_83 VNB N_A_416_86#_c_1135_n 0.00446365f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.99
cc_84 VNB N_A_416_86#_c_1136_n 0.0105037f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=2.46
cc_85 VNB N_A_416_86#_c_1137_n 0.00413213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_416_86#_c_1138_n 0.0125189f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=2.005
cc_87 VNB N_A_416_86#_c_1139_n 0.00510991f $X=-0.19 $Y=-0.245 $X2=1.535 $Y2=2.09
cc_88 VNB N_A_416_86#_c_1140_n 0.00111875f $X=-0.19 $Y=-0.245 $X2=1.535
+ $Y2=2.815
cc_89 VNB N_A_416_86#_c_1141_n 0.00685889f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=2.905
cc_90 VNB N_A_416_86#_c_1142_n 0.00325158f $X=-0.19 $Y=-0.245 $X2=4.31 $Y2=1.265
cc_91 VNB N_A_416_86#_c_1143_n 0.00927332f $X=-0.19 $Y=-0.245 $X2=1.37 $Y2=1.92
cc_92 VNB N_A_416_86#_c_1144_n 5.75165e-19 $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=2.07
cc_93 VNB N_A_416_86#_c_1145_n 0.00519916f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=2.755
cc_94 VNB N_A_416_86#_c_1146_n 0.00193968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_416_86#_c_1147_n 0.00620674f $X=-0.19 $Y=-0.245 $X2=4.31 $Y2=1.1
cc_96 VNB X 0.0563853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1276_n 0.0122953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1277_n 0.0139149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1278_n 0.101468f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=2.005
cc_100 VNB N_VGND_c_1279_n 0.0658973f $X=-0.19 $Y=-0.245 $X2=1.54 $Y2=1.165
cc_101 VNB N_VGND_c_1280_n 0.01773f $X=-0.19 $Y=-0.245 $X2=4.31 $Y2=1.265
cc_102 VNB N_VGND_c_1281_n 0.487308f $X=-0.19 $Y=-0.245 $X2=4.31 $Y2=1.905
cc_103 VNB N_VGND_c_1282_n 0.0197198f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=2.755
cc_104 VNB N_VGND_c_1283_n 0.037346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1284_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1285_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.8
cc_107 VPB N_A_84_108#_M1005_g 0.0288846f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=2.46
cc_108 VPB N_A_84_108#_c_189_n 0.0011055f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.635
cc_109 VPB N_A_84_108#_c_190_n 0.015385f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.635
cc_110 VPB N_A_84_108#_c_197_n 0.00888963f $X=-0.19 $Y=1.66 $X2=1.37 $Y2=2.005
cc_111 VPB N_A_84_108#_c_198_n 3.7562e-19 $X=-0.19 $Y=1.66 $X2=0.75 $Y2=2.005
cc_112 VPB N_A_84_108#_c_199_n 0.0010148f $X=-0.19 $Y=1.66 $X2=1.535 $Y2=2.105
cc_113 VPB N_A_84_108#_c_191_n 0.00610311f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.165
cc_114 VPB N_A_84_108#_c_201_n 0.0378013f $X=-0.19 $Y=1.66 $X2=3.725 $Y2=2.99
cc_115 VPB N_A_84_108#_c_202_n 0.0021839f $X=-0.19 $Y=1.66 $X2=1.7 $Y2=2.99
cc_116 VPB N_A_84_108#_c_203_n 0.00513258f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=2.905
cc_117 VPB N_A_84_108#_c_204_n 0.00576231f $X=-0.19 $Y=1.66 $X2=1.37 $Y2=1.92
cc_118 VPB N_A_84_108#_c_205_n 0.00854388f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=2.07
cc_119 VPB N_A_84_108#_c_192_n 0.00308986f $X=-0.19 $Y=1.66 $X2=4.06 $Y2=1.905
cc_120 VPB N_A_M1002_g 0.0272603f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.96
cc_121 VPB A 0.00242481f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_c_304_n 0.0152507f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.99
cc_123 VPB N_A_452_288#_M1008_g 0.0294109f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_452_288#_M1010_g 0.0279362f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=2.46
cc_125 VPB N_A_452_288#_c_349_n 0.00480236f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=2.905
cc_126 VPB N_A_452_288#_c_350_n 2.52059e-19 $X=-0.19 $Y=1.66 $X2=4.06 $Y2=2.755
cc_127 VPB N_A_452_288#_c_351_n 0.0170489f $X=-0.19 $Y=1.66 $X2=4.15 $Y2=1.1
cc_128 VPB N_B_M1012_g 0.0344702f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.96
cc_129 VPB N_B_c_461_n 0.0524398f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_B_c_462_n 0.0138933f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_B_M1009_g 0.0458417f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.99
cc_132 VPB N_B_c_464_n 0.108109f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.8
cc_133 VPB N_B_c_452_n 0.088932f $X=-0.19 $Y=1.66 $X2=1.37 $Y2=2.005
cc_134 VPB N_B_M1021_g 0.0252231f $X=-0.19 $Y=1.66 $X2=1.535 $Y2=2.815
cc_135 VPB N_B_c_467_n 0.00898883f $X=-0.19 $Y=1.66 $X2=1.7 $Y2=2.99
cc_136 VPB N_B_c_458_n 0.00940712f $X=-0.19 $Y=1.66 $X2=4.06 $Y2=2.755
cc_137 VPB N_B_c_459_n 0.00441473f $X=-0.19 $Y=1.66 $X2=4.15 $Y2=1.1
cc_138 VPB N_A_1157_298#_M1001_g 0.0264749f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_1157_298#_c_589_n 0.00217808f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_1157_298#_c_590_n 0.038367f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.8
cc_141 VPB N_A_1157_298#_c_591_n 0.00632848f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=2.46
cc_142 VPB N_A_1157_298#_c_592_n 0.0123461f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_1157_298#_c_585_n 0.00144102f $X=-0.19 $Y=1.66 $X2=1.37 $Y2=2.005
cc_144 VPB N_A_1157_298#_c_594_n 0.00793251f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_1157_298#_c_587_n 0.0249626f $X=-0.19 $Y=1.66 $X2=4.31 $Y2=1.905
cc_146 VPB N_C_M1003_g 0.0344864f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=1.96
cc_147 VPB N_C_c_676_n 0.0129179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_C_M1013_g 0.0298561f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.99
cc_149 VPB C 0.00111319f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.635
cc_150 VPB N_A_1218_396#_M1004_g 0.027851f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_1218_396#_c_770_n 0.00251474f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.8
cc_152 VPB N_A_1218_396#_c_763_n 0.0146357f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.635
cc_153 VPB N_A_1218_396#_c_764_n 0.00204527f $X=-0.19 $Y=1.66 $X2=0.585
+ $Y2=1.635
cc_154 VPB N_A_1218_396#_c_765_n 4.48504e-19 $X=-0.19 $Y=1.66 $X2=0.75 $Y2=2.005
cc_155 VPB N_A_1218_396#_c_766_n 0.00230679f $X=-0.19 $Y=1.66 $X2=1.535
+ $Y2=2.105
cc_156 VPB N_A_1218_396#_c_767_n 0.00142224f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.165
cc_157 VPB N_A_1218_396#_c_768_n 0.00936406f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.165
cc_158 VPB N_A_27_134#_c_853_n 0.0012385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_A_27_134#_c_861_n 0.039423f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_A_27_134#_c_857_n 0.0285325f $X=-0.19 $Y=1.66 $X2=3.725 $Y2=2.99
cc_161 VPB N_VPWR_c_933_n 0.009508f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_934_n 0.00893245f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_935_n 0.014412f $X=-0.19 $Y=1.66 $X2=0.587 $Y2=1.635
cc_164 VPB N_VPWR_c_936_n 0.0226387f $X=-0.19 $Y=1.66 $X2=0.75 $Y2=2.005
cc_165 VPB N_VPWR_c_937_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.535 $Y2=2.09
cc_166 VPB N_VPWR_c_938_n 0.0943098f $X=-0.19 $Y=1.66 $X2=1.54 $Y2=1.165
cc_167 VPB N_VPWR_c_939_n 0.0786989f $X=-0.19 $Y=1.66 $X2=4.31 $Y2=1.265
cc_168 VPB N_VPWR_c_940_n 0.0180274f $X=-0.19 $Y=1.66 $X2=4.31 $Y2=1.1
cc_169 VPB N_VPWR_c_932_n 0.115289f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_942_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.8
cc_171 VPB N_VPWR_c_943_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_387_392#_c_1016_n 0.00509183f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.99
cc_173 VPB N_A_387_392#_c_1017_n 0.0040615f $X=-0.19 $Y=1.66 $X2=0.66 $Y2=1.8
cc_174 VPB N_A_387_392#_c_1018_n 4.44827e-19 $X=-0.19 $Y=1.66 $X2=0.66 $Y2=2.46
cc_175 VPB N_A_387_392#_c_1008_n 0.0029387f $X=-0.19 $Y=1.66 $X2=0.587 $Y2=1.635
cc_176 VPB N_A_387_392#_c_1020_n 0.00754215f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_387_392#_c_1021_n 0.0105785f $X=-0.19 $Y=1.66 $X2=1.7 $Y2=2.99
cc_178 VPB N_A_387_392#_c_1022_n 0.00372676f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=2.755
cc_179 VPB N_A_387_392#_c_1015_n 0.00448988f $X=-0.19 $Y=1.66 $X2=4.31 $Y2=1.265
cc_180 VPB N_A_416_86#_c_1148_n 0.00112438f $X=-0.19 $Y=1.66 $X2=0.587 $Y2=1.92
cc_181 VPB N_A_416_86#_c_1149_n 0.0168997f $X=-0.19 $Y=1.66 $X2=3.725 $Y2=2.99
cc_182 VPB N_A_416_86#_c_1143_n 0.0205858f $X=-0.19 $Y=1.66 $X2=1.37 $Y2=1.92
cc_183 VPB N_A_416_86#_c_1144_n 0.00316813f $X=-0.19 $Y=1.66 $X2=4.06 $Y2=2.07
cc_184 VPB N_A_416_86#_c_1145_n 0.00298281f $X=-0.19 $Y=1.66 $X2=4.06 $Y2=2.755
cc_185 VPB N_A_416_86#_c_1146_n 0.00273373f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_416_86#_c_1147_n 0.00628502f $X=-0.19 $Y=1.66 $X2=4.31 $Y2=1.1
cc_187 VPB X 0.0534992f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 N_A_84_108#_c_189_n N_A_M1002_g 9.43893e-19 $X=0.585 $Y=1.635 $X2=0 $Y2=0
cc_189 N_A_84_108#_c_190_n N_A_M1002_g 0.0206452f $X=0.585 $Y=1.635 $X2=0 $Y2=0
cc_190 N_A_84_108#_c_197_n N_A_M1002_g 0.0164362f $X=1.37 $Y=2.005 $X2=0 $Y2=0
cc_191 N_A_84_108#_c_199_n N_A_M1002_g 0.0126826f $X=1.535 $Y=2.105 $X2=0 $Y2=0
cc_192 N_A_84_108#_c_202_n N_A_M1002_g 0.00413657f $X=1.7 $Y=2.99 $X2=0 $Y2=0
cc_193 N_A_84_108#_c_204_n N_A_M1002_g 0.00246831f $X=1.37 $Y=1.92 $X2=0 $Y2=0
cc_194 N_A_84_108#_M1019_g N_A_c_302_n 0.0147715f $X=0.495 $Y=0.99 $X2=0 $Y2=0
cc_195 N_A_84_108#_c_191_n N_A_c_302_n 0.0167722f $X=1.54 $Y=1.165 $X2=0 $Y2=0
cc_196 N_A_84_108#_M1019_g A 0.00388715f $X=0.495 $Y=0.99 $X2=0 $Y2=0
cc_197 N_A_84_108#_c_189_n A 0.0177031f $X=0.585 $Y=1.635 $X2=0 $Y2=0
cc_198 N_A_84_108#_c_190_n A 9.75282e-19 $X=0.585 $Y=1.635 $X2=0 $Y2=0
cc_199 N_A_84_108#_c_197_n A 0.0252129f $X=1.37 $Y=2.005 $X2=0 $Y2=0
cc_200 N_A_84_108#_c_191_n A 0.0378174f $X=1.54 $Y=1.165 $X2=0 $Y2=0
cc_201 N_A_84_108#_M1019_g N_A_c_304_n 0.00172878f $X=0.495 $Y=0.99 $X2=0 $Y2=0
cc_202 N_A_84_108#_c_189_n N_A_c_304_n 0.00102935f $X=0.585 $Y=1.635 $X2=0 $Y2=0
cc_203 N_A_84_108#_c_190_n N_A_c_304_n 0.0174427f $X=0.585 $Y=1.635 $X2=0 $Y2=0
cc_204 N_A_84_108#_c_197_n N_A_c_304_n 0.00182581f $X=1.37 $Y=2.005 $X2=0 $Y2=0
cc_205 N_A_84_108#_c_201_n N_A_452_288#_M1008_g 5.95459e-19 $X=3.725 $Y=2.99
+ $X2=0 $Y2=0
cc_206 N_A_84_108#_c_191_n N_A_452_288#_c_341_n 0.00918212f $X=1.54 $Y=1.165
+ $X2=0 $Y2=0
cc_207 N_A_84_108#_c_201_n N_A_452_288#_M1010_g 0.00137965f $X=3.725 $Y=2.99
+ $X2=0 $Y2=0
cc_208 N_A_84_108#_c_205_n N_A_452_288#_M1010_g 0.00916167f $X=3.81 $Y=2.07
+ $X2=0 $Y2=0
cc_209 N_A_84_108#_c_192_n N_A_452_288#_M1020_g 4.85181e-19 $X=4.06 $Y=1.905
+ $X2=0 $Y2=0
cc_210 N_A_84_108#_c_193_n N_A_452_288#_M1020_g 0.00119421f $X=4.31 $Y=1.1 $X2=0
+ $Y2=0
cc_211 N_A_84_108#_c_192_n N_A_452_288#_c_345_n 0.00794442f $X=4.06 $Y=1.905
+ $X2=0 $Y2=0
cc_212 N_A_84_108#_M1020_d N_A_452_288#_c_346_n 0.0066978f $X=3.84 $Y=0.625
+ $X2=0 $Y2=0
cc_213 N_A_84_108#_c_193_n N_A_452_288#_c_346_n 0.0252586f $X=4.31 $Y=1.1 $X2=0
+ $Y2=0
cc_214 N_A_84_108#_c_193_n N_A_452_288#_c_348_n 0.0234597f $X=4.31 $Y=1.1 $X2=0
+ $Y2=0
cc_215 N_A_84_108#_c_192_n N_A_452_288#_c_349_n 0.103684f $X=4.06 $Y=1.905 $X2=0
+ $Y2=0
cc_216 N_A_84_108#_c_205_n N_A_452_288#_c_350_n 0.0228172f $X=3.81 $Y=2.07 $X2=0
+ $Y2=0
cc_217 N_A_84_108#_c_192_n N_A_452_288#_c_350_n 0.0215059f $X=4.06 $Y=1.905
+ $X2=0 $Y2=0
cc_218 N_A_84_108#_c_205_n N_A_452_288#_c_351_n 0.00605898f $X=3.81 $Y=2.07
+ $X2=0 $Y2=0
cc_219 N_A_84_108#_c_192_n N_A_452_288#_c_351_n 0.00106938f $X=4.06 $Y=1.905
+ $X2=0 $Y2=0
cc_220 N_A_84_108#_c_199_n N_B_M1012_g 0.00675063f $X=1.535 $Y=2.105 $X2=0 $Y2=0
cc_221 N_A_84_108#_c_191_n N_B_M1012_g 0.00202908f $X=1.54 $Y=1.165 $X2=0 $Y2=0
cc_222 N_A_84_108#_c_201_n N_B_M1012_g 0.0186438f $X=3.725 $Y=2.99 $X2=0 $Y2=0
cc_223 N_A_84_108#_c_204_n N_B_M1012_g 0.00150482f $X=1.37 $Y=1.92 $X2=0 $Y2=0
cc_224 N_A_84_108#_c_191_n N_B_M1015_g 5.48946e-19 $X=1.54 $Y=1.165 $X2=0 $Y2=0
cc_225 N_A_84_108#_c_201_n N_B_c_461_n 0.011796f $X=3.725 $Y=2.99 $X2=0 $Y2=0
cc_226 N_A_84_108#_c_201_n N_B_M1009_g 0.0149959f $X=3.725 $Y=2.99 $X2=0 $Y2=0
cc_227 N_A_84_108#_c_201_n N_B_c_464_n 0.0182198f $X=3.725 $Y=2.99 $X2=0 $Y2=0
cc_228 N_A_84_108#_c_205_n N_B_c_464_n 0.00629714f $X=3.81 $Y=2.07 $X2=0 $Y2=0
cc_229 N_A_84_108#_c_201_n N_B_c_452_n 0.00546456f $X=3.725 $Y=2.99 $X2=0 $Y2=0
cc_230 N_A_84_108#_c_203_n N_B_c_452_n 0.00399845f $X=3.81 $Y=2.905 $X2=0 $Y2=0
cc_231 N_A_84_108#_c_205_n N_B_c_452_n 0.0349822f $X=3.81 $Y=2.07 $X2=0 $Y2=0
cc_232 N_A_84_108#_c_192_n N_B_c_452_n 0.00936063f $X=4.06 $Y=1.905 $X2=0 $Y2=0
cc_233 N_A_84_108#_c_192_n N_B_c_453_n 0.00202234f $X=4.06 $Y=1.905 $X2=0 $Y2=0
cc_234 N_A_84_108#_c_193_n N_B_c_453_n 0.00916826f $X=4.31 $Y=1.1 $X2=0 $Y2=0
cc_235 N_A_84_108#_c_192_n N_B_c_456_n 0.00544619f $X=4.06 $Y=1.905 $X2=0 $Y2=0
cc_236 N_A_84_108#_c_193_n N_B_c_456_n 4.52447e-19 $X=4.31 $Y=1.1 $X2=0 $Y2=0
cc_237 N_A_84_108#_c_198_n N_A_27_134#_M1005_s 0.00240221f $X=0.75 $Y=2.005
+ $X2=0 $Y2=0
cc_238 N_A_84_108#_M1019_g N_A_27_134#_c_847_n 0.00162247f $X=0.495 $Y=0.99
+ $X2=0 $Y2=0
cc_239 N_A_84_108#_M1019_g N_A_27_134#_c_848_n 0.0126033f $X=0.495 $Y=0.99 $X2=0
+ $Y2=0
cc_240 N_A_84_108#_M1000_d N_A_27_134#_c_849_n 0.0132999f $X=1.4 $Y=0.67 $X2=0
+ $Y2=0
cc_241 N_A_84_108#_M1019_g N_A_27_134#_c_849_n 0.0110445f $X=0.495 $Y=0.99 $X2=0
+ $Y2=0
cc_242 N_A_84_108#_c_189_n N_A_27_134#_c_849_n 0.00721272f $X=0.585 $Y=1.635
+ $X2=0 $Y2=0
cc_243 N_A_84_108#_c_190_n N_A_27_134#_c_849_n 6.97809e-19 $X=0.585 $Y=1.635
+ $X2=0 $Y2=0
cc_244 N_A_84_108#_c_191_n N_A_27_134#_c_849_n 0.0135869f $X=1.54 $Y=1.165 $X2=0
+ $Y2=0
cc_245 N_A_84_108#_M1000_d N_A_27_134#_c_850_n 0.00300777f $X=1.4 $Y=0.67 $X2=0
+ $Y2=0
cc_246 N_A_84_108#_c_191_n N_A_27_134#_c_850_n 0.0191f $X=1.54 $Y=1.165 $X2=0
+ $Y2=0
cc_247 N_A_84_108#_c_191_n N_A_27_134#_c_852_n 0.0142913f $X=1.54 $Y=1.165 $X2=0
+ $Y2=0
cc_248 N_A_84_108#_M1019_g N_A_27_134#_c_856_n 0.00542664f $X=0.495 $Y=0.99
+ $X2=0 $Y2=0
cc_249 N_A_84_108#_c_189_n N_A_27_134#_c_856_n 0.00150787f $X=0.585 $Y=1.635
+ $X2=0 $Y2=0
cc_250 N_A_84_108#_M1005_g N_A_27_134#_c_861_n 0.00937548f $X=0.66 $Y=2.46 $X2=0
+ $Y2=0
cc_251 N_A_84_108#_c_190_n N_A_27_134#_c_861_n 6.97701e-19 $X=0.585 $Y=1.635
+ $X2=0 $Y2=0
cc_252 N_A_84_108#_c_198_n N_A_27_134#_c_861_n 0.0103204f $X=0.75 $Y=2.005 $X2=0
+ $Y2=0
cc_253 N_A_84_108#_M1019_g N_A_27_134#_c_857_n 0.0115559f $X=0.495 $Y=0.99 $X2=0
+ $Y2=0
cc_254 N_A_84_108#_M1005_g N_A_27_134#_c_857_n 0.0050467f $X=0.66 $Y=2.46 $X2=0
+ $Y2=0
cc_255 N_A_84_108#_c_189_n N_A_27_134#_c_857_n 0.0342332f $X=0.585 $Y=1.635
+ $X2=0 $Y2=0
cc_256 N_A_84_108#_c_198_n N_A_27_134#_c_857_n 0.0141272f $X=0.75 $Y=2.005 $X2=0
+ $Y2=0
cc_257 N_A_84_108#_c_197_n N_VPWR_M1005_d 0.00633139f $X=1.37 $Y=2.005 $X2=-0.19
+ $Y2=-0.245
cc_258 N_A_84_108#_M1005_g N_VPWR_c_933_n 0.00360519f $X=0.66 $Y=2.46 $X2=0
+ $Y2=0
cc_259 N_A_84_108#_c_197_n N_VPWR_c_933_n 0.0237567f $X=1.37 $Y=2.005 $X2=0
+ $Y2=0
cc_260 N_A_84_108#_c_199_n N_VPWR_c_933_n 0.0350928f $X=1.535 $Y=2.105 $X2=0
+ $Y2=0
cc_261 N_A_84_108#_c_202_n N_VPWR_c_933_n 0.00998657f $X=1.7 $Y=2.99 $X2=0 $Y2=0
cc_262 N_A_84_108#_M1005_g N_VPWR_c_936_n 0.005209f $X=0.66 $Y=2.46 $X2=0 $Y2=0
cc_263 N_A_84_108#_c_201_n N_VPWR_c_938_n 0.140901f $X=3.725 $Y=2.99 $X2=0 $Y2=0
cc_264 N_A_84_108#_c_202_n N_VPWR_c_938_n 0.0235512f $X=1.7 $Y=2.99 $X2=0 $Y2=0
cc_265 N_A_84_108#_c_205_n N_VPWR_c_938_n 0.0112583f $X=3.81 $Y=2.07 $X2=0 $Y2=0
cc_266 N_A_84_108#_M1005_g N_VPWR_c_932_n 0.00987476f $X=0.66 $Y=2.46 $X2=0
+ $Y2=0
cc_267 N_A_84_108#_c_201_n N_VPWR_c_932_n 0.0738164f $X=3.725 $Y=2.99 $X2=0
+ $Y2=0
cc_268 N_A_84_108#_c_202_n N_VPWR_c_932_n 0.0126924f $X=1.7 $Y=2.99 $X2=0 $Y2=0
cc_269 N_A_84_108#_c_205_n N_VPWR_c_932_n 0.01371f $X=3.81 $Y=2.07 $X2=0 $Y2=0
cc_270 N_A_84_108#_c_204_n N_A_387_392#_c_1016_n 0.00515165f $X=1.37 $Y=1.92
+ $X2=0 $Y2=0
cc_271 N_A_84_108#_M1010_d N_A_387_392#_c_1017_n 0.00235582f $X=3.445 $Y=1.895
+ $X2=0 $Y2=0
cc_272 N_A_84_108#_c_201_n N_A_387_392#_c_1017_n 0.0865756f $X=3.725 $Y=2.99
+ $X2=0 $Y2=0
cc_273 N_A_84_108#_c_205_n N_A_387_392#_c_1017_n 0.0152396f $X=3.81 $Y=2.07
+ $X2=0 $Y2=0
cc_274 N_A_84_108#_c_201_n N_A_387_392#_c_1018_n 0.0233833f $X=3.725 $Y=2.99
+ $X2=0 $Y2=0
cc_275 N_A_84_108#_M1010_d N_A_387_392#_c_1008_n 0.00723342f $X=3.445 $Y=1.895
+ $X2=0 $Y2=0
cc_276 N_A_84_108#_c_205_n N_A_387_392#_c_1008_n 0.0533467f $X=3.81 $Y=2.07
+ $X2=0 $Y2=0
cc_277 N_A_84_108#_c_192_n N_A_387_392#_c_1008_n 0.00492429f $X=4.06 $Y=1.905
+ $X2=0 $Y2=0
cc_278 N_A_84_108#_c_205_n N_A_416_86#_c_1143_n 0.0134146f $X=3.81 $Y=2.07 $X2=0
+ $Y2=0
cc_279 N_A_84_108#_c_192_n N_A_416_86#_c_1143_n 0.0168015f $X=4.06 $Y=1.905
+ $X2=0 $Y2=0
cc_280 N_A_84_108#_c_193_n N_A_416_86#_c_1143_n 0.0048888f $X=4.31 $Y=1.1 $X2=0
+ $Y2=0
cc_281 N_A_84_108#_M1019_g N_VGND_c_1281_n 0.00457172f $X=0.495 $Y=0.99 $X2=0
+ $Y2=0
cc_282 N_A_84_108#_M1019_g N_VGND_c_1282_n 0.00305419f $X=0.495 $Y=0.99 $X2=0
+ $Y2=0
cc_283 N_A_M1002_g N_B_M1012_g 0.0207378f $X=1.31 $Y=2.46 $X2=0 $Y2=0
cc_284 N_A_c_302_n N_B_M1015_g 0.0106761f $X=1.325 $Y=1.42 $X2=0 $Y2=0
cc_285 N_A_c_302_n N_A_27_134#_c_849_n 0.0172797f $X=1.325 $Y=1.42 $X2=0 $Y2=0
cc_286 A N_A_27_134#_c_849_n 0.0123447f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_287 N_A_c_304_n N_A_27_134#_c_849_n 0.00102726f $X=1.325 $Y=1.585 $X2=0 $Y2=0
cc_288 N_A_c_302_n N_A_27_134#_c_850_n 0.00321996f $X=1.325 $Y=1.42 $X2=0 $Y2=0
cc_289 A N_A_27_134#_c_856_n 0.0039539f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_290 N_A_M1002_g N_VPWR_c_933_n 0.00875689f $X=1.31 $Y=2.46 $X2=0 $Y2=0
cc_291 N_A_M1002_g N_VPWR_c_938_n 0.00517089f $X=1.31 $Y=2.46 $X2=0 $Y2=0
cc_292 N_A_M1002_g N_VPWR_c_932_n 0.00981147f $X=1.31 $Y=2.46 $X2=0 $Y2=0
cc_293 A N_VGND_M1019_d 0.00592605f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_294 N_A_c_302_n N_VGND_c_1278_n 0.00305517f $X=1.325 $Y=1.42 $X2=0 $Y2=0
cc_295 N_A_c_302_n N_VGND_c_1281_n 0.00457172f $X=1.325 $Y=1.42 $X2=0 $Y2=0
cc_296 N_A_452_288#_M1008_g N_B_M1012_g 0.00859419f $X=2.35 $Y=2.28 $X2=0 $Y2=0
cc_297 N_A_452_288#_M1006_g N_B_M1015_g 0.0108525f $X=2.505 $Y=0.86 $X2=0 $Y2=0
cc_298 N_A_452_288#_M1008_g N_B_c_461_n 0.00543199f $X=2.35 $Y=2.28 $X2=0 $Y2=0
cc_299 N_A_452_288#_M1006_g N_B_c_448_n 0.00642456f $X=2.505 $Y=0.86 $X2=0 $Y2=0
cc_300 N_A_452_288#_M1008_g N_B_M1009_g 0.0224379f $X=2.35 $Y=2.28 $X2=0 $Y2=0
cc_301 N_A_452_288#_c_340_n N_B_M1009_g 0.0115956f $X=3.265 $Y=1.515 $X2=0 $Y2=0
cc_302 N_A_452_288#_M1010_g N_B_M1009_g 0.0267162f $X=3.355 $Y=2.315 $X2=0 $Y2=0
cc_303 N_A_452_288#_M1010_g N_B_c_464_n 0.0105864f $X=3.355 $Y=2.315 $X2=0 $Y2=0
cc_304 N_A_452_288#_M1006_g N_B_M1014_g 0.00822803f $X=2.505 $Y=0.86 $X2=0 $Y2=0
cc_305 N_A_452_288#_c_340_n N_B_M1014_g 0.00888281f $X=3.265 $Y=1.515 $X2=0
+ $Y2=0
cc_306 N_A_452_288#_M1020_g N_B_M1014_g 0.0127716f $X=3.765 $Y=0.945 $X2=0 $Y2=0
cc_307 N_A_452_288#_M1020_g N_B_c_451_n 0.00737859f $X=3.765 $Y=0.945 $X2=0
+ $Y2=0
cc_308 N_A_452_288#_c_349_n N_B_c_452_n 0.0135784f $X=4.665 $Y=1.985 $X2=0 $Y2=0
cc_309 N_A_452_288#_M1020_g N_B_c_453_n 0.0163701f $X=3.765 $Y=0.945 $X2=0 $Y2=0
cc_310 N_A_452_288#_c_345_n N_B_c_453_n 2.52437e-19 $X=3.81 $Y=1.435 $X2=0 $Y2=0
cc_311 N_A_452_288#_c_346_n N_B_c_453_n 0.0149558f $X=4.58 $Y=0.68 $X2=0 $Y2=0
cc_312 N_A_452_288#_c_348_n N_B_c_453_n 0.0076468f $X=4.72 $Y=0.86 $X2=0 $Y2=0
cc_313 N_A_452_288#_c_349_n N_B_M1011_g 0.00336399f $X=4.665 $Y=1.985 $X2=0
+ $Y2=0
cc_314 N_A_452_288#_c_352_n N_B_M1011_g 7.81465e-19 $X=4.692 $Y=1.13 $X2=0 $Y2=0
cc_315 N_A_452_288#_M1020_g N_B_c_456_n 0.00124076f $X=3.765 $Y=0.945 $X2=0
+ $Y2=0
cc_316 N_A_452_288#_c_345_n N_B_c_456_n 2.08589e-19 $X=3.81 $Y=1.435 $X2=0 $Y2=0
cc_317 N_A_452_288#_c_350_n N_B_c_456_n 4.0729e-19 $X=3.89 $Y=1.57 $X2=0 $Y2=0
cc_318 N_A_452_288#_c_351_n N_B_c_456_n 0.0180764f $X=3.89 $Y=1.57 $X2=0 $Y2=0
cc_319 N_A_452_288#_c_349_n N_B_c_457_n 0.0132684f $X=4.665 $Y=1.985 $X2=0 $Y2=0
cc_320 N_A_452_288#_c_352_n N_B_c_457_n 8.86982e-19 $X=4.692 $Y=1.13 $X2=0 $Y2=0
cc_321 N_A_452_288#_c_349_n N_B_c_458_n 0.00359336f $X=4.665 $Y=1.985 $X2=0
+ $Y2=0
cc_322 N_A_452_288#_c_349_n N_B_c_459_n 0.0307414f $X=4.665 $Y=1.985 $X2=0 $Y2=0
cc_323 N_A_452_288#_M1006_g N_A_27_134#_c_850_n 0.001394f $X=2.505 $Y=0.86 $X2=0
+ $Y2=0
cc_324 N_A_452_288#_c_341_n N_A_27_134#_c_851_n 0.00838583f $X=2.58 $Y=1.515
+ $X2=0 $Y2=0
cc_325 N_A_452_288#_M1008_g N_A_27_134#_c_853_n 0.0238758f $X=2.35 $Y=2.28 $X2=0
+ $Y2=0
cc_326 N_A_452_288#_M1006_g N_A_27_134#_c_853_n 5.71278e-19 $X=2.505 $Y=0.86
+ $X2=0 $Y2=0
cc_327 N_A_452_288#_c_340_n N_A_27_134#_c_853_n 0.0112599f $X=3.265 $Y=1.515
+ $X2=0 $Y2=0
cc_328 N_A_452_288#_c_341_n N_A_27_134#_c_853_n 0.00962286f $X=2.58 $Y=1.515
+ $X2=0 $Y2=0
cc_329 N_A_452_288#_M1006_g N_A_27_134#_c_854_n 0.00428797f $X=2.505 $Y=0.86
+ $X2=0 $Y2=0
cc_330 N_A_452_288#_M1006_g N_A_27_134#_c_858_n 0.0171903f $X=2.505 $Y=0.86
+ $X2=0 $Y2=0
cc_331 N_A_452_288#_c_340_n N_A_27_134#_c_859_n 0.00284831f $X=3.265 $Y=1.515
+ $X2=0 $Y2=0
cc_332 N_A_452_288#_c_349_n N_VPWR_c_934_n 0.0331578f $X=4.665 $Y=1.985 $X2=0
+ $Y2=0
cc_333 N_A_452_288#_c_349_n N_VPWR_c_938_n 0.00749631f $X=4.665 $Y=1.985 $X2=0
+ $Y2=0
cc_334 N_A_452_288#_c_349_n N_VPWR_c_932_n 0.0062048f $X=4.665 $Y=1.985 $X2=0
+ $Y2=0
cc_335 N_A_452_288#_M1008_g N_A_387_392#_c_1017_n 0.0131657f $X=2.35 $Y=2.28
+ $X2=0 $Y2=0
cc_336 N_A_452_288#_M1010_g N_A_387_392#_c_1017_n 0.014666f $X=3.355 $Y=2.315
+ $X2=0 $Y2=0
cc_337 N_A_452_288#_M1008_g N_A_387_392#_c_1018_n 0.00170314f $X=2.35 $Y=2.28
+ $X2=0 $Y2=0
cc_338 N_A_452_288#_M1010_g N_A_387_392#_c_1008_n 0.0284023f $X=3.355 $Y=2.315
+ $X2=0 $Y2=0
cc_339 N_A_452_288#_M1020_g N_A_387_392#_c_1008_n 0.0118517f $X=3.765 $Y=0.945
+ $X2=0 $Y2=0
cc_340 N_A_452_288#_c_344_n N_A_387_392#_c_1008_n 0.00434477f $X=3.355 $Y=1.515
+ $X2=0 $Y2=0
cc_341 N_A_452_288#_c_345_n N_A_387_392#_c_1008_n 0.0471932f $X=3.81 $Y=1.435
+ $X2=0 $Y2=0
cc_342 N_A_452_288#_c_347_n N_A_387_392#_c_1008_n 0.0133618f $X=3.895 $Y=0.68
+ $X2=0 $Y2=0
cc_343 N_A_452_288#_c_350_n N_A_387_392#_c_1008_n 0.0208077f $X=3.89 $Y=1.57
+ $X2=0 $Y2=0
cc_344 N_A_452_288#_c_351_n N_A_387_392#_c_1008_n 7.0374e-19 $X=3.89 $Y=1.57
+ $X2=0 $Y2=0
cc_345 N_A_452_288#_c_353_n N_A_387_392#_c_1008_n 0.00877596f $X=3.69 $Y=1.57
+ $X2=0 $Y2=0
cc_346 N_A_452_288#_M1011_s N_A_387_392#_c_1009_n 0.00231738f $X=4.585 $Y=0.37
+ $X2=0 $Y2=0
cc_347 N_A_452_288#_M1020_g N_A_387_392#_c_1009_n 0.00174767f $X=3.765 $Y=0.945
+ $X2=0 $Y2=0
cc_348 N_A_452_288#_c_346_n N_A_387_392#_c_1009_n 0.0643236f $X=4.58 $Y=0.68
+ $X2=0 $Y2=0
cc_349 N_A_452_288#_c_347_n N_A_387_392#_c_1009_n 0.0129683f $X=3.895 $Y=0.68
+ $X2=0 $Y2=0
cc_350 N_A_452_288#_M1006_g N_A_416_86#_c_1135_n 0.00415017f $X=2.505 $Y=0.86
+ $X2=0 $Y2=0
cc_351 N_A_452_288#_M1006_g N_A_416_86#_c_1136_n 0.00378345f $X=2.505 $Y=0.86
+ $X2=0 $Y2=0
cc_352 N_A_452_288#_c_340_n N_A_416_86#_c_1148_n 0.00170244f $X=3.265 $Y=1.515
+ $X2=0 $Y2=0
cc_353 N_A_452_288#_c_349_n N_A_416_86#_c_1139_n 0.00510874f $X=4.665 $Y=1.985
+ $X2=0 $Y2=0
cc_354 N_A_452_288#_M1010_g N_A_416_86#_c_1143_n 0.00924211f $X=3.355 $Y=2.315
+ $X2=0 $Y2=0
cc_355 N_A_452_288#_c_345_n N_A_416_86#_c_1143_n 8.6696e-19 $X=3.81 $Y=1.435
+ $X2=0 $Y2=0
cc_356 N_A_452_288#_c_349_n N_A_416_86#_c_1143_n 0.0199562f $X=4.665 $Y=1.985
+ $X2=0 $Y2=0
cc_357 N_A_452_288#_c_350_n N_A_416_86#_c_1143_n 0.017006f $X=3.89 $Y=1.57 $X2=0
+ $Y2=0
cc_358 N_A_452_288#_c_351_n N_A_416_86#_c_1143_n 0.0039441f $X=3.89 $Y=1.57
+ $X2=0 $Y2=0
cc_359 N_A_452_288#_c_352_n N_A_416_86#_c_1143_n 0.00207179f $X=4.692 $Y=1.13
+ $X2=0 $Y2=0
cc_360 N_A_452_288#_c_353_n N_A_416_86#_c_1143_n 0.00382019f $X=3.69 $Y=1.57
+ $X2=0 $Y2=0
cc_361 N_A_452_288#_c_340_n N_A_416_86#_c_1144_n 0.00374115f $X=3.265 $Y=1.515
+ $X2=0 $Y2=0
cc_362 N_A_452_288#_M1010_g N_A_416_86#_c_1144_n 0.00305294f $X=3.355 $Y=2.315
+ $X2=0 $Y2=0
cc_363 N_A_452_288#_c_344_n N_A_416_86#_c_1144_n 3.65068e-19 $X=3.355 $Y=1.515
+ $X2=0 $Y2=0
cc_364 N_A_452_288#_M1008_g N_A_416_86#_c_1145_n 7.51956e-19 $X=2.35 $Y=2.28
+ $X2=0 $Y2=0
cc_365 N_A_452_288#_M1006_g N_A_416_86#_c_1145_n 0.00268112f $X=2.505 $Y=0.86
+ $X2=0 $Y2=0
cc_366 N_A_452_288#_c_340_n N_A_416_86#_c_1145_n 0.0136802f $X=3.265 $Y=1.515
+ $X2=0 $Y2=0
cc_367 N_A_452_288#_M1010_g N_A_416_86#_c_1145_n 0.00596353f $X=3.355 $Y=2.315
+ $X2=0 $Y2=0
cc_368 N_A_452_288#_c_349_n N_A_416_86#_c_1147_n 0.00333463f $X=4.665 $Y=1.985
+ $X2=0 $Y2=0
cc_369 N_B_c_458_n N_A_1157_298#_c_587_n 0.00334116f $X=5.085 $Y=1.515 $X2=0
+ $Y2=0
cc_370 N_B_M1015_g N_A_27_134#_c_849_n 0.00578498f $X=2.005 $Y=0.75 $X2=0 $Y2=0
cc_371 N_B_M1015_g N_A_27_134#_c_850_n 0.00996021f $X=2.005 $Y=0.75 $X2=0 $Y2=0
cc_372 N_B_M1015_g N_A_27_134#_c_851_n 0.00536183f $X=2.005 $Y=0.75 $X2=0 $Y2=0
cc_373 N_B_M1012_g N_A_27_134#_c_852_n 0.00519185f $X=1.845 $Y=2.38 $X2=0 $Y2=0
cc_374 N_B_M1012_g N_A_27_134#_c_853_n 6.06199e-19 $X=1.845 $Y=2.38 $X2=0 $Y2=0
cc_375 N_B_M1009_g N_A_27_134#_c_853_n 0.00981834f $X=2.82 $Y=2.28 $X2=0 $Y2=0
cc_376 N_B_M1014_g N_A_27_134#_c_854_n 0.00151817f $X=3.175 $Y=0.75 $X2=0 $Y2=0
cc_377 N_B_M1014_g N_A_27_134#_c_855_n 3.58404e-19 $X=3.175 $Y=0.75 $X2=0 $Y2=0
cc_378 N_B_c_462_n N_VPWR_c_933_n 0.00181942f $X=1.935 $Y=3.15 $X2=0 $Y2=0
cc_379 N_B_c_464_n N_VPWR_c_934_n 0.00229165f $X=4.295 $Y=3.15 $X2=0 $Y2=0
cc_380 N_B_c_452_n N_VPWR_c_934_n 7.81718e-19 $X=4.37 $Y=3.075 $X2=0 $Y2=0
cc_381 N_B_M1021_g N_VPWR_c_934_n 0.0180017f $X=4.89 $Y=2.4 $X2=0 $Y2=0
cc_382 N_B_c_458_n N_VPWR_c_934_n 0.00120263f $X=5.085 $Y=1.515 $X2=0 $Y2=0
cc_383 N_B_c_459_n N_VPWR_c_934_n 0.0177783f $X=5.085 $Y=1.515 $X2=0 $Y2=0
cc_384 N_B_c_462_n N_VPWR_c_938_n 0.0600103f $X=1.935 $Y=3.15 $X2=0 $Y2=0
cc_385 N_B_M1021_g N_VPWR_c_938_n 0.00460063f $X=4.89 $Y=2.4 $X2=0 $Y2=0
cc_386 N_B_c_461_n N_VPWR_c_932_n 0.0187316f $X=2.73 $Y=3.15 $X2=0 $Y2=0
cc_387 N_B_c_462_n N_VPWR_c_932_n 0.0067422f $X=1.935 $Y=3.15 $X2=0 $Y2=0
cc_388 N_B_c_464_n N_VPWR_c_932_n 0.0417446f $X=4.295 $Y=3.15 $X2=0 $Y2=0
cc_389 N_B_M1021_g N_VPWR_c_932_n 0.00909358f $X=4.89 $Y=2.4 $X2=0 $Y2=0
cc_390 N_B_c_467_n N_VPWR_c_932_n 0.00445015f $X=2.82 $Y=3.15 $X2=0 $Y2=0
cc_391 N_B_M1012_g N_A_387_392#_c_1016_n 0.00707946f $X=1.845 $Y=2.38 $X2=0
+ $Y2=0
cc_392 N_B_M1009_g N_A_387_392#_c_1017_n 0.016695f $X=2.82 $Y=2.28 $X2=0 $Y2=0
cc_393 N_B_M1012_g N_A_387_392#_c_1018_n 0.00313279f $X=1.845 $Y=2.38 $X2=0
+ $Y2=0
cc_394 N_B_M1009_g N_A_387_392#_c_1008_n 9.65487e-19 $X=2.82 $Y=2.28 $X2=0 $Y2=0
cc_395 N_B_M1014_g N_A_387_392#_c_1008_n 0.00677596f $X=3.175 $Y=0.75 $X2=0
+ $Y2=0
cc_396 N_B_c_451_n N_A_387_392#_c_1009_n 0.0143527f $X=4.36 $Y=0.18 $X2=0 $Y2=0
cc_397 N_B_c_453_n N_A_387_392#_c_1009_n 0.0121042f $X=4.435 $Y=1.35 $X2=0 $Y2=0
cc_398 N_B_M1011_g N_A_387_392#_c_1009_n 0.0134432f $X=4.935 $Y=0.74 $X2=0 $Y2=0
cc_399 N_B_M1014_g N_A_387_392#_c_1010_n 0.00428767f $X=3.175 $Y=0.75 $X2=0
+ $Y2=0
cc_400 N_B_c_451_n N_A_387_392#_c_1010_n 0.00420304f $X=4.36 $Y=0.18 $X2=0 $Y2=0
cc_401 N_B_c_453_n N_A_387_392#_c_1057_n 9.69016e-19 $X=4.435 $Y=1.35 $X2=0
+ $Y2=0
cc_402 N_B_M1011_g N_A_387_392#_c_1057_n 0.0131592f $X=4.935 $Y=0.74 $X2=0 $Y2=0
cc_403 N_B_c_458_n N_A_387_392#_c_1011_n 6.33323e-19 $X=5.085 $Y=1.515 $X2=0
+ $Y2=0
cc_404 N_B_c_459_n N_A_387_392#_c_1011_n 0.00419509f $X=5.085 $Y=1.515 $X2=0
+ $Y2=0
cc_405 N_B_M1011_g N_A_387_392#_c_1061_n 0.00669508f $X=4.935 $Y=0.74 $X2=0
+ $Y2=0
cc_406 N_B_c_458_n N_A_387_392#_c_1061_n 7.49096e-19 $X=5.085 $Y=1.515 $X2=0
+ $Y2=0
cc_407 N_B_c_459_n N_A_387_392#_c_1061_n 0.00628567f $X=5.085 $Y=1.515 $X2=0
+ $Y2=0
cc_408 N_B_c_448_n N_A_416_86#_c_1136_n 0.0120727f $X=3.1 $Y=0.18 $X2=0 $Y2=0
cc_409 N_B_M1014_g N_A_416_86#_c_1136_n 0.00809565f $X=3.175 $Y=0.75 $X2=0 $Y2=0
cc_410 N_B_M1015_g N_A_416_86#_c_1137_n 0.0064969f $X=2.005 $Y=0.75 $X2=0 $Y2=0
cc_411 N_B_c_448_n N_A_416_86#_c_1137_n 0.00524214f $X=3.1 $Y=0.18 $X2=0 $Y2=0
cc_412 N_B_M1009_g N_A_416_86#_c_1148_n 0.00310476f $X=2.82 $Y=2.28 $X2=0 $Y2=0
cc_413 N_B_M1011_g N_A_416_86#_c_1139_n 0.00313168f $X=4.935 $Y=0.74 $X2=0 $Y2=0
cc_414 N_B_c_458_n N_A_416_86#_c_1139_n 2.72398e-19 $X=5.085 $Y=1.515 $X2=0
+ $Y2=0
cc_415 N_B_c_459_n N_A_416_86#_c_1139_n 8.43333e-19 $X=5.085 $Y=1.515 $X2=0
+ $Y2=0
cc_416 N_B_c_452_n N_A_416_86#_c_1143_n 0.00524423f $X=4.37 $Y=3.075 $X2=0 $Y2=0
cc_417 N_B_M1021_g N_A_416_86#_c_1143_n 0.00537789f $X=4.89 $Y=2.4 $X2=0 $Y2=0
cc_418 N_B_c_457_n N_A_416_86#_c_1143_n 0.00133956f $X=4.8 $Y=1.515 $X2=0 $Y2=0
cc_419 N_B_c_458_n N_A_416_86#_c_1143_n 0.00605591f $X=5.085 $Y=1.515 $X2=0
+ $Y2=0
cc_420 N_B_c_459_n N_A_416_86#_c_1143_n 0.0215037f $X=5.085 $Y=1.515 $X2=0 $Y2=0
cc_421 N_B_M1009_g N_A_416_86#_c_1145_n 3.82365e-19 $X=2.82 $Y=2.28 $X2=0 $Y2=0
cc_422 N_B_M1014_g N_A_416_86#_c_1145_n 0.020973f $X=3.175 $Y=0.75 $X2=0 $Y2=0
cc_423 N_B_c_458_n N_A_416_86#_c_1146_n 8.53932e-19 $X=5.085 $Y=1.515 $X2=0
+ $Y2=0
cc_424 N_B_c_459_n N_A_416_86#_c_1146_n 0.00272458f $X=5.085 $Y=1.515 $X2=0
+ $Y2=0
cc_425 N_B_M1021_g N_A_416_86#_c_1147_n 0.00298486f $X=4.89 $Y=2.4 $X2=0 $Y2=0
cc_426 N_B_c_458_n N_A_416_86#_c_1147_n 0.00504527f $X=5.085 $Y=1.515 $X2=0
+ $Y2=0
cc_427 N_B_c_459_n N_A_416_86#_c_1147_n 0.0301947f $X=5.085 $Y=1.515 $X2=0 $Y2=0
cc_428 N_B_M1011_g N_VGND_c_1276_n 0.00266853f $X=4.935 $Y=0.74 $X2=0 $Y2=0
cc_429 N_B_c_449_n N_VGND_c_1278_n 0.0607067f $X=2.08 $Y=0.18 $X2=0 $Y2=0
cc_430 N_B_M1011_g N_VGND_c_1278_n 0.00278237f $X=4.935 $Y=0.74 $X2=0 $Y2=0
cc_431 N_B_c_448_n N_VGND_c_1281_n 0.0260329f $X=3.1 $Y=0.18 $X2=0 $Y2=0
cc_432 N_B_c_449_n N_VGND_c_1281_n 0.0104612f $X=2.08 $Y=0.18 $X2=0 $Y2=0
cc_433 N_B_c_451_n N_VGND_c_1281_n 0.0367758f $X=4.36 $Y=0.18 $X2=0 $Y2=0
cc_434 N_B_M1011_g N_VGND_c_1281_n 0.00359083f $X=4.935 $Y=0.74 $X2=0 $Y2=0
cc_435 N_B_c_455_n N_VGND_c_1281_n 0.00501319f $X=3.175 $Y=0.18 $X2=0 $Y2=0
cc_436 N_A_1157_298#_M1001_g N_C_M1003_g 0.0113625f $X=6 $Y=2.4 $X2=0 $Y2=0
cc_437 N_A_1157_298#_c_589_n N_C_M1003_g 0.00397264f $X=6.11 $Y=2.905 $X2=0
+ $Y2=0
cc_438 N_A_1157_298#_c_590_n N_C_M1003_g 0.0124373f $X=7.435 $Y=2.99 $X2=0 $Y2=0
cc_439 N_A_1157_298#_c_592_n N_C_M1003_g 0.00377356f $X=7.52 $Y=2.905 $X2=0
+ $Y2=0
cc_440 N_A_1157_298#_M1016_g N_C_c_674_n 0.00807795f $X=6.155 $Y=0.925 $X2=0
+ $Y2=0
cc_441 N_A_1157_298#_c_585_n N_C_c_675_n 0.00273498f $X=7.9 $Y=2.195 $X2=0 $Y2=0
cc_442 N_A_1157_298#_c_594_n N_C_c_675_n 0.0040882f $X=7.9 $Y=2.36 $X2=0 $Y2=0
cc_443 N_A_1157_298#_c_604_p N_C_c_676_n 2.34839e-19 $X=6.11 $Y=1.675 $X2=0
+ $Y2=0
cc_444 N_A_1157_298#_c_587_n N_C_c_676_n 0.0146706f $X=6.155 $Y=1.655 $X2=0
+ $Y2=0
cc_445 N_A_1157_298#_c_585_n N_C_c_677_n 0.0116958f $X=7.9 $Y=2.195 $X2=0 $Y2=0
cc_446 N_A_1157_298#_c_592_n N_C_M1013_g 0.00247829f $X=7.52 $Y=2.905 $X2=0
+ $Y2=0
cc_447 N_A_1157_298#_c_585_n N_C_M1013_g 0.0223158f $X=7.9 $Y=2.195 $X2=0 $Y2=0
cc_448 N_A_1157_298#_c_594_n N_C_M1013_g 0.0110328f $X=7.9 $Y=2.36 $X2=0 $Y2=0
cc_449 N_A_1157_298#_c_584_n N_C_c_679_n 0.00442451f $X=7.9 $Y=0.63 $X2=0 $Y2=0
cc_450 N_A_1157_298#_c_585_n N_C_c_679_n 0.00125427f $X=7.9 $Y=2.195 $X2=0 $Y2=0
cc_451 N_A_1157_298#_c_586_n N_C_c_679_n 0.00302306f $X=7.94 $Y=0.86 $X2=0 $Y2=0
cc_452 N_A_1157_298#_c_585_n N_C_c_680_n 0.00942884f $X=7.9 $Y=2.195 $X2=0 $Y2=0
cc_453 N_A_1157_298#_c_586_n N_C_c_680_n 0.00241658f $X=7.94 $Y=0.86 $X2=0 $Y2=0
cc_454 N_A_1157_298#_c_585_n N_C_c_681_n 0.005861f $X=7.9 $Y=2.195 $X2=0 $Y2=0
cc_455 N_A_1157_298#_c_589_n N_A_1218_396#_M1001_d 0.00835578f $X=6.11 $Y=2.905
+ $X2=0 $Y2=0
cc_456 N_A_1157_298#_c_585_n N_A_1218_396#_M1004_g 9.01237e-19 $X=7.9 $Y=2.195
+ $X2=0 $Y2=0
cc_457 N_A_1157_298#_c_585_n N_A_1218_396#_M1018_g 9.59011e-19 $X=7.9 $Y=2.195
+ $X2=0 $Y2=0
cc_458 N_A_1157_298#_M1001_g N_A_1218_396#_c_770_n 0.00304464f $X=6 $Y=2.4 $X2=0
+ $Y2=0
cc_459 N_A_1157_298#_c_589_n N_A_1218_396#_c_770_n 0.0705476f $X=6.11 $Y=2.905
+ $X2=0 $Y2=0
cc_460 N_A_1157_298#_c_590_n N_A_1218_396#_c_770_n 0.0236382f $X=7.435 $Y=2.99
+ $X2=0 $Y2=0
cc_461 N_A_1157_298#_M1016_g N_A_1218_396#_c_762_n 0.00470692f $X=6.155 $Y=0.925
+ $X2=0 $Y2=0
cc_462 N_A_1157_298#_c_604_p N_A_1218_396#_c_762_n 8.40914e-19 $X=6.11 $Y=1.675
+ $X2=0 $Y2=0
cc_463 N_A_1157_298#_c_585_n N_A_1218_396#_c_763_n 0.0173001f $X=7.9 $Y=2.195
+ $X2=0 $Y2=0
cc_464 N_A_1157_298#_c_594_n N_A_1218_396#_c_763_n 0.00751637f $X=7.9 $Y=2.36
+ $X2=0 $Y2=0
cc_465 N_A_1157_298#_c_604_p N_A_1218_396#_c_764_n 0.00748663f $X=6.11 $Y=1.675
+ $X2=0 $Y2=0
cc_466 N_A_1157_298#_c_587_n N_A_1218_396#_c_764_n 0.004852f $X=6.155 $Y=1.655
+ $X2=0 $Y2=0
cc_467 N_A_1157_298#_c_604_p N_A_1218_396#_c_765_n 0.0185876f $X=6.11 $Y=1.675
+ $X2=0 $Y2=0
cc_468 N_A_1157_298#_c_587_n N_A_1218_396#_c_765_n 0.00241039f $X=6.155 $Y=1.655
+ $X2=0 $Y2=0
cc_469 N_A_1157_298#_c_585_n N_A_1218_396#_c_766_n 0.00219668f $X=7.9 $Y=2.195
+ $X2=0 $Y2=0
cc_470 N_A_1157_298#_c_585_n N_A_1218_396#_c_767_n 0.0188137f $X=7.9 $Y=2.195
+ $X2=0 $Y2=0
cc_471 N_A_1157_298#_c_585_n N_A_1218_396#_c_768_n 0.00120897f $X=7.9 $Y=2.195
+ $X2=0 $Y2=0
cc_472 N_A_1157_298#_c_590_n N_VPWR_c_935_n 0.00609169f $X=7.435 $Y=2.99 $X2=0
+ $Y2=0
cc_473 N_A_1157_298#_c_592_n N_VPWR_c_935_n 0.0121857f $X=7.52 $Y=2.905 $X2=0
+ $Y2=0
cc_474 N_A_1157_298#_c_585_n N_VPWR_c_935_n 0.0139215f $X=7.9 $Y=2.195 $X2=0
+ $Y2=0
cc_475 N_A_1157_298#_c_594_n N_VPWR_c_935_n 0.0204024f $X=7.9 $Y=2.36 $X2=0
+ $Y2=0
cc_476 N_A_1157_298#_M1001_g N_VPWR_c_939_n 0.00398971f $X=6 $Y=2.4 $X2=0 $Y2=0
cc_477 N_A_1157_298#_c_590_n N_VPWR_c_939_n 0.0918162f $X=7.435 $Y=2.99 $X2=0
+ $Y2=0
cc_478 N_A_1157_298#_c_591_n N_VPWR_c_939_n 0.0121867f $X=6.195 $Y=2.99 $X2=0
+ $Y2=0
cc_479 N_A_1157_298#_M1001_g N_VPWR_c_932_n 0.00385171f $X=6 $Y=2.4 $X2=0 $Y2=0
cc_480 N_A_1157_298#_c_590_n N_VPWR_c_932_n 0.0531866f $X=7.435 $Y=2.99 $X2=0
+ $Y2=0
cc_481 N_A_1157_298#_c_591_n N_VPWR_c_932_n 0.00660921f $X=6.195 $Y=2.99 $X2=0
+ $Y2=0
cc_482 N_A_1157_298#_c_594_n N_VPWR_c_932_n 0.0138596f $X=7.9 $Y=2.36 $X2=0
+ $Y2=0
cc_483 N_A_1157_298#_M1016_g N_A_387_392#_c_1012_n 0.0050953f $X=6.155 $Y=0.925
+ $X2=0 $Y2=0
cc_484 N_A_1157_298#_M1016_g N_A_387_392#_c_1013_n 0.00650284f $X=6.155 $Y=0.925
+ $X2=0 $Y2=0
cc_485 N_A_1157_298#_c_584_n N_A_387_392#_c_1013_n 0.00216124f $X=7.9 $Y=0.63
+ $X2=0 $Y2=0
cc_486 N_A_1157_298#_c_590_n N_A_387_392#_c_1020_n 0.0244008f $X=7.435 $Y=2.99
+ $X2=0 $Y2=0
cc_487 N_A_1157_298#_c_592_n N_A_387_392#_c_1020_n 0.0134807f $X=7.52 $Y=2.905
+ $X2=0 $Y2=0
cc_488 N_A_1157_298#_c_594_n N_A_387_392#_c_1020_n 0.0230767f $X=7.9 $Y=2.36
+ $X2=0 $Y2=0
cc_489 N_A_1157_298#_M1013_s N_A_387_392#_c_1021_n 0.00516465f $X=7.455 $Y=1.865
+ $X2=0 $Y2=0
cc_490 N_A_1157_298#_c_585_n N_A_387_392#_c_1021_n 0.00798748f $X=7.9 $Y=2.195
+ $X2=0 $Y2=0
cc_491 N_A_1157_298#_c_594_n N_A_387_392#_c_1021_n 0.0168712f $X=7.9 $Y=2.36
+ $X2=0 $Y2=0
cc_492 N_A_1157_298#_c_584_n N_A_387_392#_c_1015_n 0.105953f $X=7.9 $Y=0.63
+ $X2=0 $Y2=0
cc_493 N_A_1157_298#_M1016_g N_A_416_86#_c_1138_n 0.016605f $X=6.155 $Y=0.925
+ $X2=0 $Y2=0
cc_494 N_A_1157_298#_c_604_p N_A_416_86#_c_1138_n 0.0285588f $X=6.11 $Y=1.675
+ $X2=0 $Y2=0
cc_495 N_A_1157_298#_c_587_n N_A_416_86#_c_1138_n 0.00773078f $X=6.155 $Y=1.655
+ $X2=0 $Y2=0
cc_496 N_A_1157_298#_M1016_g N_A_416_86#_c_1200_n 0.0147634f $X=6.155 $Y=0.925
+ $X2=0 $Y2=0
cc_497 N_A_1157_298#_M1016_g N_A_416_86#_c_1140_n 0.00532072f $X=6.155 $Y=0.925
+ $X2=0 $Y2=0
cc_498 N_A_1157_298#_M1001_g N_A_416_86#_c_1149_n 0.0133313f $X=6 $Y=2.4 $X2=0
+ $Y2=0
cc_499 N_A_1157_298#_c_589_n N_A_416_86#_c_1149_n 0.0235442f $X=6.11 $Y=2.905
+ $X2=0 $Y2=0
cc_500 N_A_1157_298#_c_604_p N_A_416_86#_c_1149_n 0.00400233f $X=6.11 $Y=1.675
+ $X2=0 $Y2=0
cc_501 N_A_1157_298#_c_587_n N_A_416_86#_c_1149_n 0.00175309f $X=6.155 $Y=1.655
+ $X2=0 $Y2=0
cc_502 N_A_1157_298#_c_604_p N_A_416_86#_c_1146_n 0.00752565f $X=6.11 $Y=1.675
+ $X2=0 $Y2=0
cc_503 N_A_1157_298#_c_587_n N_A_416_86#_c_1146_n 0.00598257f $X=6.155 $Y=1.655
+ $X2=0 $Y2=0
cc_504 N_A_1157_298#_M1001_g N_A_416_86#_c_1147_n 0.00252015f $X=6 $Y=2.4 $X2=0
+ $Y2=0
cc_505 N_A_1157_298#_M1016_g N_A_416_86#_c_1147_n 0.00334445f $X=6.155 $Y=0.925
+ $X2=0 $Y2=0
cc_506 N_A_1157_298#_c_589_n N_A_416_86#_c_1147_n 0.00495515f $X=6.11 $Y=2.905
+ $X2=0 $Y2=0
cc_507 N_A_1157_298#_c_604_p N_A_416_86#_c_1147_n 0.0187176f $X=6.11 $Y=1.675
+ $X2=0 $Y2=0
cc_508 N_A_1157_298#_c_587_n N_A_416_86#_c_1147_n 0.00585289f $X=6.155 $Y=1.655
+ $X2=0 $Y2=0
cc_509 N_A_1157_298#_c_584_n N_VGND_c_1277_n 0.0172844f $X=7.9 $Y=0.63 $X2=0
+ $Y2=0
cc_510 N_A_1157_298#_c_585_n N_VGND_c_1277_n 0.0177801f $X=7.9 $Y=2.195 $X2=0
+ $Y2=0
cc_511 N_A_1157_298#_c_584_n N_VGND_c_1279_n 0.00906588f $X=7.9 $Y=0.63 $X2=0
+ $Y2=0
cc_512 N_A_1157_298#_c_584_n N_VGND_c_1281_n 0.00881689f $X=7.9 $Y=0.63 $X2=0
+ $Y2=0
cc_513 N_C_M1013_g N_A_1218_396#_M1004_g 0.0111129f $X=7.925 $Y=2.185 $X2=0
+ $Y2=0
cc_514 N_C_c_677_n N_A_1218_396#_M1018_g 0.00454574f $X=7.91 $Y=1.355 $X2=0
+ $Y2=0
cc_515 N_C_c_679_n N_A_1218_396#_M1018_g 0.012648f $X=8.115 $Y=0.915 $X2=0 $Y2=0
cc_516 N_C_M1003_g N_A_1218_396#_c_770_n 0.0218948f $X=6.755 $Y=2.4 $X2=0 $Y2=0
cc_517 N_C_c_674_n N_A_1218_396#_c_762_n 0.00340146f $X=6.835 $Y=1.355 $X2=0
+ $Y2=0
cc_518 N_C_c_676_n N_A_1218_396#_c_762_n 0.00129045f $X=7.205 $Y=1.43 $X2=0
+ $Y2=0
cc_519 C N_A_1218_396#_c_762_n 0.0341858f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_520 N_C_M1003_g N_A_1218_396#_c_763_n 0.00658635f $X=6.755 $Y=2.4 $X2=0 $Y2=0
cc_521 N_C_c_675_n N_A_1218_396#_c_763_n 0.0103253f $X=7.835 $Y=1.43 $X2=0 $Y2=0
cc_522 N_C_c_676_n N_A_1218_396#_c_763_n 0.010922f $X=7.205 $Y=1.43 $X2=0 $Y2=0
cc_523 N_C_M1013_g N_A_1218_396#_c_763_n 0.00228157f $X=7.925 $Y=2.185 $X2=0
+ $Y2=0
cc_524 N_C_c_680_n N_A_1218_396#_c_763_n 0.00394827f $X=8.115 $Y=0.99 $X2=0
+ $Y2=0
cc_525 N_C_c_681_n N_A_1218_396#_c_763_n 5.15044e-19 $X=7.835 $Y=1.355 $X2=0
+ $Y2=0
cc_526 C N_A_1218_396#_c_763_n 0.0222255f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_527 C N_A_1218_396#_c_764_n 2.70695e-19 $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_528 N_C_M1003_g N_A_1218_396#_c_765_n 0.00124812f $X=6.755 $Y=2.4 $X2=0 $Y2=0
cc_529 N_C_c_676_n N_A_1218_396#_c_765_n 0.00363065f $X=7.205 $Y=1.43 $X2=0
+ $Y2=0
cc_530 N_C_M1013_g N_A_1218_396#_c_766_n 7.19809e-19 $X=7.925 $Y=2.185 $X2=0
+ $Y2=0
cc_531 N_C_c_681_n N_A_1218_396#_c_766_n 2.41308e-19 $X=7.835 $Y=1.355 $X2=0
+ $Y2=0
cc_532 N_C_c_677_n N_A_1218_396#_c_767_n 6.83592e-19 $X=7.91 $Y=1.355 $X2=0
+ $Y2=0
cc_533 N_C_M1013_g N_A_1218_396#_c_767_n 6.77156e-19 $X=7.925 $Y=2.185 $X2=0
+ $Y2=0
cc_534 N_C_c_681_n N_A_1218_396#_c_767_n 6.3673e-19 $X=7.835 $Y=1.355 $X2=0
+ $Y2=0
cc_535 N_C_c_677_n N_A_1218_396#_c_768_n 0.0074916f $X=7.91 $Y=1.355 $X2=0 $Y2=0
cc_536 N_C_c_681_n N_A_1218_396#_c_768_n 0.00988772f $X=7.835 $Y=1.355 $X2=0
+ $Y2=0
cc_537 N_C_M1013_g N_VPWR_c_935_n 0.00639038f $X=7.925 $Y=2.185 $X2=0 $Y2=0
cc_538 N_C_M1003_g N_VPWR_c_939_n 8.29751e-19 $X=6.755 $Y=2.4 $X2=0 $Y2=0
cc_539 N_C_M1013_g N_VPWR_c_939_n 0.00388757f $X=7.925 $Y=2.185 $X2=0 $Y2=0
cc_540 N_C_M1013_g N_VPWR_c_932_n 0.00501024f $X=7.925 $Y=2.185 $X2=0 $Y2=0
cc_541 N_C_c_674_n N_A_387_392#_c_1013_n 0.00455332f $X=6.835 $Y=1.355 $X2=0
+ $Y2=0
cc_542 N_C_c_679_n N_A_387_392#_c_1013_n 0.00226061f $X=8.115 $Y=0.915 $X2=0
+ $Y2=0
cc_543 N_C_M1013_g N_A_387_392#_c_1020_n 0.00156757f $X=7.925 $Y=2.185 $X2=0
+ $Y2=0
cc_544 N_C_c_675_n N_A_387_392#_c_1021_n 0.00759068f $X=7.835 $Y=1.43 $X2=0
+ $Y2=0
cc_545 N_C_M1013_g N_A_387_392#_c_1021_n 0.00128696f $X=7.925 $Y=2.185 $X2=0
+ $Y2=0
cc_546 N_C_M1003_g N_A_387_392#_c_1022_n 0.00307356f $X=6.755 $Y=2.4 $X2=0 $Y2=0
cc_547 N_C_c_676_n N_A_387_392#_c_1022_n 0.00258432f $X=7.205 $Y=1.43 $X2=0
+ $Y2=0
cc_548 C N_A_387_392#_c_1022_n 0.0231272f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_549 N_C_M1003_g N_A_387_392#_c_1015_n 0.00319825f $X=6.755 $Y=2.4 $X2=0 $Y2=0
cc_550 N_C_c_674_n N_A_387_392#_c_1015_n 0.00922302f $X=6.835 $Y=1.355 $X2=0
+ $Y2=0
cc_551 N_C_c_675_n N_A_387_392#_c_1015_n 0.0148537f $X=7.835 $Y=1.43 $X2=0 $Y2=0
cc_552 N_C_c_676_n N_A_387_392#_c_1015_n 0.00151744f $X=7.205 $Y=1.43 $X2=0
+ $Y2=0
cc_553 N_C_c_679_n N_A_387_392#_c_1015_n 7.49501e-19 $X=8.115 $Y=0.915 $X2=0
+ $Y2=0
cc_554 N_C_c_680_n N_A_387_392#_c_1015_n 0.00294884f $X=8.115 $Y=0.99 $X2=0
+ $Y2=0
cc_555 N_C_c_681_n N_A_387_392#_c_1015_n 0.00177524f $X=7.835 $Y=1.355 $X2=0
+ $Y2=0
cc_556 C N_A_387_392#_c_1015_n 0.0258981f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_557 C N_A_416_86#_M1007_d 0.00392197f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_558 N_C_c_674_n N_A_416_86#_c_1200_n 0.00166996f $X=6.835 $Y=1.355 $X2=0
+ $Y2=0
cc_559 N_C_c_674_n N_A_416_86#_c_1141_n 0.0040941f $X=6.835 $Y=1.355 $X2=0 $Y2=0
cc_560 N_C_c_676_n N_A_416_86#_c_1141_n 0.00382945f $X=7.205 $Y=1.43 $X2=0 $Y2=0
cc_561 C N_A_416_86#_c_1141_n 0.0159889f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_562 N_C_c_674_n N_A_416_86#_c_1142_n 0.0113393f $X=6.835 $Y=1.355 $X2=0 $Y2=0
cc_563 C N_A_416_86#_c_1142_n 3.08063e-19 $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_564 N_C_c_677_n N_VGND_c_1277_n 9.50408e-19 $X=7.91 $Y=1.355 $X2=0 $Y2=0
cc_565 N_C_c_679_n N_VGND_c_1277_n 0.00636152f $X=8.115 $Y=0.915 $X2=0 $Y2=0
cc_566 N_C_c_679_n N_VGND_c_1279_n 0.00517302f $X=8.115 $Y=0.915 $X2=0 $Y2=0
cc_567 N_C_c_679_n N_VGND_c_1281_n 0.00529924f $X=8.115 $Y=0.915 $X2=0 $Y2=0
cc_568 N_A_1218_396#_M1004_g N_VPWR_c_935_n 0.021239f $X=8.615 $Y=2.4 $X2=0
+ $Y2=0
cc_569 N_A_1218_396#_c_763_n N_VPWR_c_935_n 0.00143929f $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_570 N_A_1218_396#_c_766_n N_VPWR_c_935_n 0.00246002f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_571 N_A_1218_396#_c_767_n N_VPWR_c_935_n 0.0197205f $X=8.42 $Y=1.515 $X2=0
+ $Y2=0
cc_572 N_A_1218_396#_c_768_n N_VPWR_c_935_n 0.00151227f $X=8.615 $Y=1.515 $X2=0
+ $Y2=0
cc_573 N_A_1218_396#_M1004_g N_VPWR_c_940_n 0.00460063f $X=8.615 $Y=2.4 $X2=0
+ $Y2=0
cc_574 N_A_1218_396#_M1004_g N_VPWR_c_932_n 0.00912296f $X=8.615 $Y=2.4 $X2=0
+ $Y2=0
cc_575 N_A_1218_396#_c_763_n N_A_387_392#_c_1021_n 0.012851f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_576 N_A_1218_396#_c_770_n N_A_387_392#_c_1022_n 0.0122192f $X=6.53 $Y=2.125
+ $X2=0 $Y2=0
cc_577 N_A_1218_396#_c_763_n N_A_387_392#_c_1022_n 0.0091904f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_578 N_A_1218_396#_c_763_n N_A_387_392#_c_1015_n 0.0141719f $X=8.255 $Y=1.665
+ $X2=0 $Y2=0
cc_579 N_A_1218_396#_M1016_d N_A_416_86#_c_1138_n 5.22721e-19 $X=6.23 $Y=0.605
+ $X2=0 $Y2=0
cc_580 N_A_1218_396#_c_762_n N_A_416_86#_c_1138_n 0.0141867f $X=6.62 $Y=1.1
+ $X2=0 $Y2=0
cc_581 N_A_1218_396#_c_764_n N_A_416_86#_c_1138_n 0.00161571f $X=6.625 $Y=1.665
+ $X2=0 $Y2=0
cc_582 N_A_1218_396#_M1016_d N_A_416_86#_c_1200_n 0.00463943f $X=6.23 $Y=0.605
+ $X2=0 $Y2=0
cc_583 N_A_1218_396#_c_762_n N_A_416_86#_c_1200_n 0.0184851f $X=6.62 $Y=1.1
+ $X2=0 $Y2=0
cc_584 N_A_1218_396#_M1016_d N_A_416_86#_c_1142_n 0.0097578f $X=6.23 $Y=0.605
+ $X2=0 $Y2=0
cc_585 N_A_1218_396#_c_762_n N_A_416_86#_c_1142_n 0.0135869f $X=6.62 $Y=1.1
+ $X2=0 $Y2=0
cc_586 N_A_1218_396#_M1018_g X 0.0138917f $X=8.625 $Y=0.79 $X2=0 $Y2=0
cc_587 N_A_1218_396#_c_766_n X 0.00157351f $X=8.4 $Y=1.665 $X2=0 $Y2=0
cc_588 N_A_1218_396#_c_767_n X 0.0316568f $X=8.42 $Y=1.515 $X2=0 $Y2=0
cc_589 N_A_1218_396#_c_768_n X 0.0104194f $X=8.615 $Y=1.515 $X2=0 $Y2=0
cc_590 N_A_1218_396#_M1018_g N_VGND_c_1277_n 0.0167539f $X=8.625 $Y=0.79 $X2=0
+ $Y2=0
cc_591 N_A_1218_396#_c_763_n N_VGND_c_1277_n 3.56247e-19 $X=8.255 $Y=1.665 $X2=0
+ $Y2=0
cc_592 N_A_1218_396#_c_766_n N_VGND_c_1277_n 0.00156605f $X=8.4 $Y=1.665 $X2=0
+ $Y2=0
cc_593 N_A_1218_396#_c_767_n N_VGND_c_1277_n 0.0258718f $X=8.42 $Y=1.515 $X2=0
+ $Y2=0
cc_594 N_A_1218_396#_c_768_n N_VGND_c_1277_n 0.00232457f $X=8.615 $Y=1.515 $X2=0
+ $Y2=0
cc_595 N_A_1218_396#_M1018_g N_VGND_c_1280_n 0.00449979f $X=8.625 $Y=0.79 $X2=0
+ $Y2=0
cc_596 N_A_1218_396#_M1018_g N_VGND_c_1281_n 0.00445136f $X=8.625 $Y=0.79 $X2=0
+ $Y2=0
cc_597 N_A_27_134#_c_861_n N_VPWR_c_933_n 0.0297094f $X=0.435 $Y=2.425 $X2=0
+ $Y2=0
cc_598 N_A_27_134#_c_861_n N_VPWR_c_936_n 0.0228676f $X=0.435 $Y=2.425 $X2=0
+ $Y2=0
cc_599 N_A_27_134#_c_861_n N_VPWR_c_932_n 0.0188319f $X=0.435 $Y=2.425 $X2=0
+ $Y2=0
cc_600 N_A_27_134#_c_851_n N_A_387_392#_c_1016_n 0.0115589f $X=2.43 $Y=1.345
+ $X2=0 $Y2=0
cc_601 N_A_27_134#_c_852_n N_A_387_392#_c_1016_n 0.00146236f $X=1.965 $Y=1.345
+ $X2=0 $Y2=0
cc_602 N_A_27_134#_c_853_n N_A_387_392#_c_1016_n 0.0359609f $X=2.595 $Y=2.205
+ $X2=0 $Y2=0
cc_603 N_A_27_134#_M1008_d N_A_387_392#_c_1017_n 0.00187091f $X=2.44 $Y=1.96
+ $X2=0 $Y2=0
cc_604 N_A_27_134#_c_853_n N_A_387_392#_c_1017_n 0.0171295f $X=2.595 $Y=2.205
+ $X2=0 $Y2=0
cc_605 N_A_27_134#_c_850_n N_A_416_86#_c_1135_n 0.00953553f $X=1.88 $Y=1.26
+ $X2=0 $Y2=0
cc_606 N_A_27_134#_c_851_n N_A_416_86#_c_1135_n 0.0209457f $X=2.43 $Y=1.345
+ $X2=0 $Y2=0
cc_607 N_A_27_134#_c_854_n N_A_416_86#_c_1135_n 0.00266566f $X=2.765 $Y=0.86
+ $X2=0 $Y2=0
cc_608 N_A_27_134#_M1006_d N_A_416_86#_c_1136_n 0.00897407f $X=2.58 $Y=0.65
+ $X2=0 $Y2=0
cc_609 N_A_27_134#_c_854_n N_A_416_86#_c_1136_n 0.0197667f $X=2.765 $Y=0.86
+ $X2=0 $Y2=0
cc_610 N_A_27_134#_c_853_n N_A_416_86#_c_1148_n 0.0197348f $X=2.595 $Y=2.205
+ $X2=0 $Y2=0
cc_611 N_A_27_134#_c_853_n N_A_416_86#_c_1144_n 0.00712425f $X=2.595 $Y=2.205
+ $X2=0 $Y2=0
cc_612 N_A_27_134#_M1006_d N_A_416_86#_c_1145_n 0.00695839f $X=2.58 $Y=0.65
+ $X2=0 $Y2=0
cc_613 N_A_27_134#_c_853_n N_A_416_86#_c_1145_n 0.0216652f $X=2.595 $Y=2.205
+ $X2=0 $Y2=0
cc_614 N_A_27_134#_c_854_n N_A_416_86#_c_1145_n 0.0348734f $X=2.765 $Y=0.86
+ $X2=0 $Y2=0
cc_615 N_A_27_134#_c_855_n N_A_416_86#_c_1145_n 0.00956728f $X=2.675 $Y=1.26
+ $X2=0 $Y2=0
cc_616 N_A_27_134#_c_858_n N_A_416_86#_c_1145_n 0.010767f $X=2.595 $Y=1.345
+ $X2=0 $Y2=0
cc_617 N_A_27_134#_c_849_n N_VGND_M1019_d 0.0217869f $X=1.795 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_618 N_A_27_134#_c_849_n N_VGND_c_1278_n 0.0125374f $X=1.795 $Y=0.745 $X2=0
+ $Y2=0
cc_619 N_A_27_134#_c_847_n N_VGND_c_1281_n 0.0107619f $X=0.265 $Y=0.83 $X2=0
+ $Y2=0
cc_620 N_A_27_134#_c_849_n N_VGND_c_1281_n 0.0288798f $X=1.795 $Y=0.745 $X2=0
+ $Y2=0
cc_621 N_A_27_134#_c_847_n N_VGND_c_1282_n 0.00699929f $X=0.265 $Y=0.83 $X2=0
+ $Y2=0
cc_622 N_A_27_134#_c_849_n N_VGND_c_1282_n 0.00286374f $X=1.795 $Y=0.745 $X2=0
+ $Y2=0
cc_623 N_A_27_134#_c_849_n N_VGND_c_1283_n 0.0436747f $X=1.795 $Y=0.745 $X2=0
+ $Y2=0
cc_624 N_VPWR_c_934_n N_A_416_86#_c_1149_n 0.0637424f $X=5.115 $Y=2.115 $X2=0
+ $Y2=0
cc_625 N_VPWR_c_939_n N_A_416_86#_c_1149_n 0.0127204f $X=8.225 $Y=3.33 $X2=0
+ $Y2=0
cc_626 N_VPWR_c_932_n N_A_416_86#_c_1149_n 0.0150935f $X=8.88 $Y=3.33 $X2=0
+ $Y2=0
cc_627 N_VPWR_c_934_n N_A_416_86#_c_1143_n 0.00189255f $X=5.115 $Y=2.115 $X2=0
+ $Y2=0
cc_628 N_VPWR_c_935_n X 0.0346097f $X=8.39 $Y=2.115 $X2=0 $Y2=0
cc_629 N_VPWR_c_940_n X 0.011066f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_630 N_VPWR_c_932_n X 0.00915947f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_631 N_A_387_392#_c_1017_n N_A_416_86#_M1009_d 0.00420616f $X=3.385 $Y=2.65
+ $X2=0 $Y2=0
cc_632 N_A_387_392#_c_1008_n N_A_416_86#_c_1136_n 0.00271974f $X=3.47 $Y=0.575
+ $X2=0 $Y2=0
cc_633 N_A_387_392#_c_1010_n N_A_416_86#_c_1136_n 0.0120353f $X=3.555 $Y=0.34
+ $X2=0 $Y2=0
cc_634 N_A_387_392#_c_1017_n N_A_416_86#_c_1246_n 0.0195146f $X=3.385 $Y=2.65
+ $X2=0 $Y2=0
cc_635 N_A_387_392#_M1016_s N_A_416_86#_c_1138_n 0.00260133f $X=5.805 $Y=0.605
+ $X2=0 $Y2=0
cc_636 N_A_387_392#_c_1011_n N_A_416_86#_c_1138_n 0.0313943f $X=5.775 $Y=0.935
+ $X2=0 $Y2=0
cc_637 N_A_387_392#_c_1011_n N_A_416_86#_c_1139_n 0.0166871f $X=5.775 $Y=0.935
+ $X2=0 $Y2=0
cc_638 N_A_387_392#_c_1012_n N_A_416_86#_c_1140_n 0.00752165f $X=5.94 $Y=0.8
+ $X2=0 $Y2=0
cc_639 N_A_387_392#_c_1013_n N_A_416_86#_c_1140_n 0.0132904f $X=7.475 $Y=0.34
+ $X2=0 $Y2=0
cc_640 N_A_387_392#_c_1015_n N_A_416_86#_c_1141_n 0.0271845f $X=7.56 $Y=1.855
+ $X2=0 $Y2=0
cc_641 N_A_387_392#_c_1013_n N_A_416_86#_c_1142_n 0.0675114f $X=7.475 $Y=0.34
+ $X2=0 $Y2=0
cc_642 N_A_387_392#_c_1008_n N_A_416_86#_c_1143_n 0.0202635f $X=3.47 $Y=0.575
+ $X2=0 $Y2=0
cc_643 N_A_387_392#_c_1011_n N_A_416_86#_c_1143_n 0.00435893f $X=5.775 $Y=0.935
+ $X2=0 $Y2=0
cc_644 N_A_387_392#_c_1061_n N_A_416_86#_c_1143_n 9.19195e-19 $X=5.145 $Y=0.935
+ $X2=0 $Y2=0
cc_645 N_A_387_392#_c_1008_n N_A_416_86#_c_1144_n 0.00230122f $X=3.47 $Y=0.575
+ $X2=0 $Y2=0
cc_646 N_A_387_392#_c_1008_n N_A_416_86#_c_1145_n 0.118341f $X=3.47 $Y=0.575
+ $X2=0 $Y2=0
cc_647 N_A_387_392#_c_1011_n N_A_416_86#_c_1146_n 0.00236341f $X=5.775 $Y=0.935
+ $X2=0 $Y2=0
cc_648 N_A_387_392#_c_1009_n N_VGND_M1011_d 6.10141e-19 $X=4.975 $Y=0.34 $X2=0
+ $Y2=0
cc_649 N_A_387_392#_c_1057_n N_VGND_M1011_d 0.00596645f $X=5.06 $Y=0.85 $X2=0
+ $Y2=0
cc_650 N_A_387_392#_c_1011_n N_VGND_M1011_d 0.0146644f $X=5.775 $Y=0.935 $X2=0
+ $Y2=0
cc_651 N_A_387_392#_c_1061_n N_VGND_M1011_d 9.32214e-19 $X=5.145 $Y=0.935 $X2=0
+ $Y2=0
cc_652 N_A_387_392#_c_1009_n N_VGND_c_1276_n 0.0145685f $X=4.975 $Y=0.34 $X2=0
+ $Y2=0
cc_653 N_A_387_392#_c_1057_n N_VGND_c_1276_n 0.0190358f $X=5.06 $Y=0.85 $X2=0
+ $Y2=0
cc_654 N_A_387_392#_c_1011_n N_VGND_c_1276_n 0.0198396f $X=5.775 $Y=0.935 $X2=0
+ $Y2=0
cc_655 N_A_387_392#_c_1012_n N_VGND_c_1276_n 0.0175231f $X=5.94 $Y=0.8 $X2=0
+ $Y2=0
cc_656 N_A_387_392#_c_1014_n N_VGND_c_1276_n 0.0127057f $X=6.025 $Y=0.34 $X2=0
+ $Y2=0
cc_657 N_A_387_392#_c_1013_n N_VGND_c_1277_n 0.00528234f $X=7.475 $Y=0.34 $X2=0
+ $Y2=0
cc_658 N_A_387_392#_c_1009_n N_VGND_c_1278_n 0.102695f $X=4.975 $Y=0.34 $X2=0
+ $Y2=0
cc_659 N_A_387_392#_c_1010_n N_VGND_c_1278_n 0.0115893f $X=3.555 $Y=0.34 $X2=0
+ $Y2=0
cc_660 N_A_387_392#_c_1013_n N_VGND_c_1279_n 0.105535f $X=7.475 $Y=0.34 $X2=0
+ $Y2=0
cc_661 N_A_387_392#_c_1014_n N_VGND_c_1279_n 0.0179217f $X=6.025 $Y=0.34 $X2=0
+ $Y2=0
cc_662 N_A_387_392#_c_1009_n N_VGND_c_1281_n 0.0553872f $X=4.975 $Y=0.34 $X2=0
+ $Y2=0
cc_663 N_A_387_392#_c_1010_n N_VGND_c_1281_n 0.00583135f $X=3.555 $Y=0.34 $X2=0
+ $Y2=0
cc_664 N_A_387_392#_c_1011_n N_VGND_c_1281_n 0.0138386f $X=5.775 $Y=0.935 $X2=0
+ $Y2=0
cc_665 N_A_387_392#_c_1013_n N_VGND_c_1281_n 0.061118f $X=7.475 $Y=0.34 $X2=0
+ $Y2=0
cc_666 N_A_387_392#_c_1014_n N_VGND_c_1281_n 0.00971942f $X=6.025 $Y=0.34 $X2=0
+ $Y2=0
cc_667 N_A_416_86#_c_1136_n N_VGND_c_1278_n 0.0445568f $X=3.02 $Y=0.375 $X2=0
+ $Y2=0
cc_668 N_A_416_86#_c_1137_n N_VGND_c_1278_n 0.0146589f $X=2.385 $Y=0.375 $X2=0
+ $Y2=0
cc_669 N_A_416_86#_c_1136_n N_VGND_c_1281_n 0.0273833f $X=3.02 $Y=0.375 $X2=0
+ $Y2=0
cc_670 N_A_416_86#_c_1137_n N_VGND_c_1281_n 0.00855245f $X=2.385 $Y=0.375 $X2=0
+ $Y2=0
cc_671 X N_VGND_c_1277_n 0.0294122f $X=8.795 $Y=0.47 $X2=0 $Y2=0
cc_672 X N_VGND_c_1280_n 0.00920966f $X=8.795 $Y=0.47 $X2=0 $Y2=0
cc_673 X N_VGND_c_1281_n 0.00887807f $X=8.795 $Y=0.47 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__o32a_4.pex.spice
* Created: Fri Aug 28 18:03:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O32A_4%A_83_256# 1 2 3 4 15 19 21 25 29 33 37 41 45
+ 47 48 55 56 58 59 62 64 68 72 74
c170 74 0 1.29542e-19 $X=2.27 $Y=1.195
c171 64 0 6.51508e-20 $X=4.23 $Y=1.015
c172 59 0 7.30872e-20 $X=3.395 $Y=1.92
c173 55 0 2.93174e-19 $X=2.1 $Y=1.445
c174 29 0 8.40338e-20 $X=1.065 $Y=0.74
c175 25 0 1.0009e-19 $X=0.955 $Y=2.4
c176 15 0 3.54028e-20 $X=0.505 $Y=2.4
r177 86 87 67.3763 $w=2.79e-07 $l=3.9e-07 $layer=POLY_cond $X=1.635 $Y=1.445
+ $X2=2.025 $Y2=1.445
r178 85 86 31.0968 $w=2.79e-07 $l=1.8e-07 $layer=POLY_cond $X=1.455 $Y=1.445
+ $X2=1.635 $Y2=1.445
r179 78 79 7.46939 $w=2.94e-07 $l=1.8e-07 $layer=LI1_cond $X=3.395 $Y=1.015
+ $X2=3.395 $Y2=1.195
r180 70 72 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=4.395 $Y=0.93
+ $X2=4.395 $Y2=0.81
r181 66 81 4.74481 $w=1.7e-07 $l=1.96415e-07 $layer=LI1_cond $X=3.575 $Y=2.105
+ $X2=3.402 $Y2=2.055
r182 66 68 119.064 $w=1.68e-07 $l=1.825e-06 $layer=LI1_cond $X=3.575 $Y=2.105
+ $X2=5.4 $Y2=2.105
r183 65 78 3.94234 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.56 $Y=1.015
+ $X2=3.395 $Y2=1.015
r184 64 70 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.23 $Y=1.015
+ $X2=4.395 $Y2=0.93
r185 64 65 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.23 $Y=1.015
+ $X2=3.56 $Y2=1.015
r186 60 78 3.72042 $w=2.94e-07 $l=1.00995e-07 $layer=LI1_cond $X=3.43 $Y=0.93
+ $X2=3.395 $Y2=1.015
r187 60 62 5.31897 $w=2.58e-07 $l=1.2e-07 $layer=LI1_cond $X=3.43 $Y=0.93
+ $X2=3.43 $Y2=0.81
r188 59 81 3.02136 $w=3.3e-07 $l=1.38456e-07 $layer=LI1_cond $X=3.395 $Y=1.92
+ $X2=3.402 $Y2=2.055
r189 58 79 3.3163 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.395 $Y=1.28
+ $X2=3.395 $Y2=1.195
r190 58 59 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=3.395 $Y=1.28
+ $X2=3.395 $Y2=1.92
r191 57 74 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.355 $Y=1.195
+ $X2=2.27 $Y2=1.195
r192 56 79 3.94234 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.23 $Y=1.195
+ $X2=3.395 $Y2=1.195
r193 56 57 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=3.23 $Y=1.195
+ $X2=2.355 $Y2=1.195
r194 55 89 15.5484 $w=2.79e-07 $l=9e-08 $layer=POLY_cond $X=2.1 $Y=1.445
+ $X2=2.19 $Y2=1.445
r195 55 87 12.957 $w=2.79e-07 $l=7.5e-08 $layer=POLY_cond $X=2.1 $Y=1.445
+ $X2=2.025 $Y2=1.445
r196 54 55 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.1
+ $Y=1.445 $X2=2.1 $Y2=1.445
r197 51 85 6.0466 $w=2.79e-07 $l=3.5e-08 $layer=POLY_cond $X=1.42 $Y=1.445
+ $X2=1.455 $Y2=1.445
r198 50 54 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.42 $Y=1.445
+ $X2=2.1 $Y2=1.445
r199 50 51 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.42
+ $Y=1.445 $X2=1.42 $Y2=1.445
r200 48 74 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.27 $Y=1.445
+ $X2=2.27 $Y2=1.195
r201 48 54 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.185 $Y=1.445
+ $X2=2.1 $Y2=1.445
r202 43 89 17.2686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.19 $Y=1.28
+ $X2=2.19 $Y2=1.445
r203 43 45 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.19 $Y=1.28
+ $X2=2.19 $Y2=0.74
r204 39 87 13.0446 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.025 $Y=1.61
+ $X2=2.025 $Y2=1.445
r205 39 41 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=2.025 $Y=1.61
+ $X2=2.025 $Y2=2.4
r206 35 86 17.2686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.635 $Y=1.28
+ $X2=1.635 $Y2=1.445
r207 35 37 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.635 $Y=1.28
+ $X2=1.635 $Y2=0.74
r208 31 85 13.0446 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.455 $Y=1.61
+ $X2=1.455 $Y2=1.445
r209 31 33 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=1.455 $Y=1.61
+ $X2=1.455 $Y2=2.4
r210 27 51 61.3298 $w=2.79e-07 $l=4.29651e-07 $layer=POLY_cond $X=1.065 $Y=1.28
+ $X2=1.42 $Y2=1.445
r211 27 29 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.065 $Y=1.28
+ $X2=1.065 $Y2=0.74
r212 23 27 19.0036 $w=2.79e-07 $l=1.97484e-07 $layer=POLY_cond $X=0.955 $Y=1.43
+ $X2=1.065 $Y2=1.28
r213 23 25 377.048 $w=1.8e-07 $l=9.7e-07 $layer=POLY_cond $X=0.955 $Y=1.43
+ $X2=0.955 $Y2=2.4
r214 22 47 6.66866 $w=1.5e-07 $l=1.48e-07 $layer=POLY_cond $X=0.71 $Y=1.355
+ $X2=0.562 $Y2=1.355
r215 21 23 25.7874 $w=2.79e-07 $l=1.21861e-07 $layer=POLY_cond $X=0.865 $Y=1.355
+ $X2=0.955 $Y2=1.43
r216 21 22 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=0.865 $Y=1.355
+ $X2=0.71 $Y2=1.355
r217 17 47 18.8402 $w=1.65e-07 $l=1.05357e-07 $layer=POLY_cond $X=0.635 $Y=1.28
+ $X2=0.562 $Y2=1.355
r218 17 19 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=0.635 $Y=1.28
+ $X2=0.635 $Y2=0.74
r219 13 47 18.8402 $w=1.65e-07 $l=9.94987e-08 $layer=POLY_cond $X=0.505 $Y=1.43
+ $X2=0.562 $Y2=1.355
r220 13 15 377.048 $w=1.8e-07 $l=9.7e-07 $layer=POLY_cond $X=0.505 $Y=1.43
+ $X2=0.505 $Y2=2.4
r221 4 68 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.265
+ $Y=1.96 $X2=5.4 $Y2=2.105
r222 3 81 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=3.275
+ $Y=1.94 $X2=3.41 $Y2=2.095
r223 2 72 182 $w=1.7e-07 $l=5.3479e-07 $layer=licon1_NDIFF $count=1 $X=4.185
+ $Y=0.37 $X2=4.395 $Y2=0.81
r224 1 62 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=3.255
+ $Y=0.37 $X2=3.395 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_4%B1 3 6 7 8 9 11 12 14 16 17 19 20 21 23 24 26
+ 27 28 29 32 34 35 39 46 54
c144 54 0 1.62575e-19 $X=2.77 $Y=1.615
c145 35 0 6.51508e-20 $X=4.66 $Y=1.615
c146 34 0 7.47943e-20 $X=4.66 $Y=1.615
c147 12 0 7.30872e-20 $X=3.535 $Y=1.165
c148 8 0 1.29542e-19 $X=2.855 $Y=1.165
r149 44 46 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.69 $Y=1.615
+ $X2=2.78 $Y2=1.615
r150 41 44 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=2.595 $Y=1.615
+ $X2=2.69 $Y2=1.615
r151 39 54 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=2.64 $Y=1.615
+ $X2=2.77 $Y2=1.615
r152 39 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.615 $X2=2.69 $Y2=1.615
r153 35 50 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.66 $Y=1.615
+ $X2=4.66 $Y2=1.78
r154 34 37 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.66 $Y=1.615
+ $X2=4.66 $Y2=1.765
r155 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.66
+ $Y=1.615 $X2=4.66 $Y2=1.615
r156 31 32 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.82 $Y=1.85
+ $X2=5.82 $Y2=2.36
r157 30 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.825 $Y=1.765
+ $X2=4.66 $Y2=1.765
r158 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.735 $Y=1.765
+ $X2=5.82 $Y2=1.85
r159 29 30 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=5.735 $Y=1.765
+ $X2=4.825 $Y2=1.765
r160 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.735 $Y=2.445
+ $X2=5.82 $Y2=2.36
r161 27 28 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=5.735 $Y=2.445
+ $X2=2.855 $Y2=2.445
r162 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.77 $Y=2.36
+ $X2=2.855 $Y2=2.445
r163 25 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.77 $Y=1.78
+ $X2=2.77 $Y2=1.615
r164 25 26 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=2.77 $Y=1.78
+ $X2=2.77 $Y2=2.36
r165 23 50 633.266 $w=1.5e-07 $l=1.235e-06 $layer=POLY_cond $X=4.655 $Y=3.015
+ $X2=4.655 $Y2=1.78
r166 20 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.58 $Y=3.09
+ $X2=4.655 $Y2=3.015
r167 20 21 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=4.58 $Y=3.09
+ $X2=4.175 $Y2=3.09
r168 17 21 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.085 $Y=3.015
+ $X2=4.175 $Y2=3.09
r169 17 19 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.085 $Y=3.015
+ $X2=4.085 $Y2=2.44
r170 14 16 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.61 $Y=1.09 $X2=3.61
+ $Y2=0.69
r171 13 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.255 $Y=1.165
+ $X2=3.18 $Y2=1.165
r172 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.535 $Y=1.165
+ $X2=3.61 $Y2=1.09
r173 12 13 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.535 $Y=1.165
+ $X2=3.255 $Y2=1.165
r174 9 24 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.18 $Y=1.09
+ $X2=3.18 $Y2=1.165
r175 9 11 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.18 $Y=1.09 $X2=3.18
+ $Y2=0.69
r176 7 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.105 $Y=1.165
+ $X2=3.18 $Y2=1.165
r177 7 8 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=3.105 $Y=1.165
+ $X2=2.855 $Y2=1.165
r178 6 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.78 $Y=1.45
+ $X2=2.78 $Y2=1.615
r179 5 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.78 $Y=1.24
+ $X2=2.855 $Y2=1.165
r180 5 6 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.78 $Y=1.24 $X2=2.78
+ $Y2=1.45
r181 1 41 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.595 $Y=1.78
+ $X2=2.595 $Y2=1.615
r182 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.595 $Y=1.78
+ $X2=2.595 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_4%B2 1 3 4 5 6 8 9 11 13 14 16 18 22 24 27 28
r77 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.09
+ $Y=1.435 $X2=4.09 $Y2=1.435
r78 24 28 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=4.09 $Y=1.665
+ $X2=4.09 $Y2=1.435
r79 23 27 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.09 $Y=1.45
+ $X2=4.09 $Y2=1.435
r80 21 27 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=4.09 $Y=1.24
+ $X2=4.09 $Y2=1.435
r81 21 22 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=4.09 $Y=1.24
+ $X2=4.09 $Y2=1.165
r82 19 20 79.8313 $w=1.6e-07 $l=2.65e-07 $layer=POLY_cond $X=3.635 $Y=1.525
+ $X2=3.635 $Y2=1.79
r83 16 18 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.61 $Y=1.09 $X2=4.61
+ $Y2=0.69
r84 15 22 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.255 $Y=1.165
+ $X2=4.09 $Y2=1.165
r85 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.535 $Y=1.165
+ $X2=4.61 $Y2=1.09
r86 14 15 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.535 $Y=1.165
+ $X2=4.255 $Y2=1.165
r87 11 22 13.5877 $w=2.4e-07 $l=8.44097e-08 $layer=POLY_cond $X=4.11 $Y=1.09
+ $X2=4.09 $Y2=1.165
r88 11 13 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.11 $Y=1.09 $X2=4.11
+ $Y2=0.69
r89 10 19 4.37345 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.725 $Y=1.525
+ $X2=3.635 $Y2=1.525
r90 9 23 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.925 $Y=1.525
+ $X2=4.09 $Y2=1.45
r91 9 10 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=3.925 $Y=1.525
+ $X2=3.725 $Y2=1.525
r92 6 20 20.7934 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.635 $Y=1.865
+ $X2=3.635 $Y2=1.79
r93 6 8 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.635 $Y=1.865
+ $X2=3.635 $Y2=2.44
r94 4 20 4.37345 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.545 $Y=1.79 $X2=3.635
+ $Y2=1.79
r95 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.545 $Y=1.79
+ $X2=3.275 $Y2=1.79
r96 1 5 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.185 $Y=1.865
+ $X2=3.275 $Y2=1.79
r97 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.185 $Y=1.865
+ $X2=3.185 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_4%A3 3 7 9 11 14 18 19 27
c63 27 0 7.47943e-20 $X=5.66 $Y=1.345
c64 3 0 3.01827e-20 $X=5.14 $Y=0.69
r65 25 27 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.57 $Y=1.345 $X2=5.66
+ $Y2=1.345
r66 23 25 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=5.175 $Y=1.345
+ $X2=5.57 $Y2=1.345
r67 21 23 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=5.14 $Y=1.345
+ $X2=5.175 $Y2=1.345
r68 19 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.57
+ $Y=1.345 $X2=5.57 $Y2=1.345
r69 16 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.66 $Y=1.51
+ $X2=5.66 $Y2=1.345
r70 16 18 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=5.66 $Y=1.51
+ $X2=5.66 $Y2=1.75
r71 12 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.66 $Y=1.18
+ $X2=5.66 $Y2=1.345
r72 12 14 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=5.66 $Y=1.18
+ $X2=5.66 $Y2=0.69
r73 9 18 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.645 $Y=1.84 $X2=5.645
+ $Y2=1.75
r74 9 11 166.022 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=5.645 $Y=1.84
+ $X2=5.645 $Y2=2.46
r75 5 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.175 $Y=1.51
+ $X2=5.175 $Y2=1.345
r76 5 7 369.274 $w=1.8e-07 $l=9.5e-07 $layer=POLY_cond $X=5.175 $Y=1.51
+ $X2=5.175 $Y2=2.46
r77 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.14 $Y=1.18
+ $X2=5.14 $Y2=1.345
r78 1 3 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=5.14 $Y=1.18 $X2=5.14
+ $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_4%A2 3 5 7 8 10 13 17 20 21 22 23 24 32 33 35
+ 42 54
c92 21 0 1.50094e-19 $X=6.395 $Y=1.58
c93 8 0 1.91837e-19 $X=6.61 $Y=1.085
r94 40 42 4.15909 $w=1.98e-07 $l=7.5e-08 $layer=LI1_cond $X=6.405 $Y=1.68
+ $X2=6.48 $Y2=1.68
r95 36 54 7.53752 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.73 $Y=1.615
+ $X2=7.565 $Y2=1.615
r96 35 38 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.73 $Y=1.615
+ $X2=7.73 $Y2=1.78
r97 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.73
+ $Y=1.615 $X2=7.73 $Y2=1.615
r98 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.24
+ $Y=1.295 $X2=6.24 $Y2=1.295
r99 24 36 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=7.92 $Y=1.615
+ $X2=7.73 $Y2=1.615
r100 23 54 6.93182 $w=1.98e-07 $l=1.25e-07 $layer=LI1_cond $X=7.44 $Y=1.68
+ $X2=7.565 $Y2=1.68
r101 22 23 26.6182 $w=1.98e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.68
+ $X2=7.44 $Y2=1.68
r102 21 40 4.52169 $w=2e-07 $l=1.69926e-07 $layer=LI1_cond $X=6.24 $Y=1.69
+ $X2=6.405 $Y2=1.68
r103 21 33 9.66018 $w=3.38e-07 $l=2.85e-07 $layer=LI1_cond $X=6.24 $Y=1.58
+ $X2=6.24 $Y2=1.295
r104 21 22 26.3409 $w=1.98e-07 $l=4.75e-07 $layer=LI1_cond $X=6.485 $Y=1.68
+ $X2=6.96 $Y2=1.68
r105 21 42 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=6.485 $Y=1.68
+ $X2=6.48 $Y2=1.68
r106 19 32 42.4067 $w=4e-07 $l=3.05e-07 $layer=POLY_cond $X=6.205 $Y=1.6
+ $X2=6.205 $Y2=1.295
r107 19 20 44.8438 $w=4e-07 $l=2e-07 $layer=POLY_cond $X=6.205 $Y=1.6 $X2=6.205
+ $Y2=1.8
r108 17 32 8.34231 $w=4e-07 $l=6e-08 $layer=POLY_cond $X=6.205 $Y=1.235
+ $X2=6.205 $Y2=1.295
r109 17 18 131.899 $w=1.48e-07 $l=4.05e-07 $layer=POLY_cond $X=6.205 $Y=1.16
+ $X2=6.61 $Y2=1.16
r110 15 17 30.9392 $w=1.48e-07 $l=9.5e-08 $layer=POLY_cond $X=6.11 $Y=1.16
+ $X2=6.205 $Y2=1.16
r111 13 38 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=7.655 $Y=2.46
+ $X2=7.655 $Y2=1.78
r112 8 18 2.50663 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.61 $Y=1.085
+ $X2=6.61 $Y2=1.16
r113 8 10 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.61 $Y=1.085
+ $X2=6.61 $Y2=0.69
r114 5 15 2.50663 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.11 $Y=1.085
+ $X2=6.11 $Y2=1.16
r115 5 7 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.11 $Y=1.085
+ $X2=6.11 $Y2=0.69
r116 3 20 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=6.095 $Y=2.46
+ $X2=6.095 $Y2=1.8
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_4%A1 1 3 4 6 7 9 10 12 14 22 23 26 27
c62 7 0 2.39531e-19 $X=7.205 $Y=1.885
c63 1 0 8.99845e-20 $X=6.735 $Y=1.885
r64 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.13
+ $Y=1.285 $X2=7.13 $Y2=1.285
r65 23 27 6.7557 $w=2.88e-07 $l=1.7e-07 $layer=LI1_cond $X=6.96 $Y=1.265
+ $X2=7.13 $Y2=1.265
r66 21 26 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=7.13 $Y=1.24
+ $X2=7.13 $Y2=1.285
r67 21 22 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=7.13 $Y=1.24
+ $X2=7.13 $Y2=1.165
r68 18 26 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=7.13 $Y=1.735
+ $X2=7.13 $Y2=1.285
r69 12 14 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=7.665 $Y=1.09
+ $X2=7.665 $Y2=0.69
r70 11 22 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.295 $Y=1.165
+ $X2=7.13 $Y2=1.165
r71 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.59 $Y=1.165
+ $X2=7.665 $Y2=1.09
r72 10 11 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=7.59 $Y=1.165
+ $X2=7.295 $Y2=1.165
r73 7 18 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.205 $Y=1.81
+ $X2=7.13 $Y2=1.81
r74 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.205 $Y=1.885
+ $X2=7.205 $Y2=2.46
r75 4 22 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=7.04 $Y=1.09
+ $X2=7.13 $Y2=1.165
r76 4 6 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=7.04 $Y=1.09 $X2=7.04
+ $Y2=0.69
r77 1 18 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.735 $Y=1.81
+ $X2=7.13 $Y2=1.81
r78 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.735 $Y=1.885
+ $X2=6.735 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_4%VPWR 1 2 3 4 5 16 18 24 26 30 36 40 43 44 45
+ 47 59 68 69 75 78 81
r99 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r100 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r101 76 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r102 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r103 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r104 69 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=6.96 $Y2=3.33
r105 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r106 66 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.135 $Y=3.33
+ $X2=6.97 $Y2=3.33
r107 66 68 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=7.135 $Y=3.33
+ $X2=7.92 $Y2=3.33
r108 65 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r109 64 65 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r110 62 65 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r111 61 64 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r112 61 62 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r113 59 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.805 $Y=3.33
+ $X2=6.97 $Y2=3.33
r114 59 64 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.805 $Y=3.33
+ $X2=6.48 $Y2=3.33
r115 55 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r116 54 57 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r117 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r118 52 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=3.33
+ $X2=2.25 $Y2=3.33
r119 52 54 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.415 $Y=3.33
+ $X2=2.64 $Y2=3.33
r120 51 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r121 51 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r122 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r123 48 72 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r124 48 50 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r125 47 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.23 $Y2=3.33
r126 47 50 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.72 $Y2=3.33
r127 45 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r128 45 55 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r129 45 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r130 43 57 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.195 $Y=3.33
+ $X2=4.08 $Y2=3.33
r131 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.195 $Y=3.33
+ $X2=4.36 $Y2=3.33
r132 42 61 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.525 $Y=3.33
+ $X2=4.56 $Y2=3.33
r133 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.525 $Y=3.33
+ $X2=4.36 $Y2=3.33
r134 38 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.97 $Y=3.245
+ $X2=6.97 $Y2=3.33
r135 38 40 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.97 $Y=3.245
+ $X2=6.97 $Y2=2.815
r136 34 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.36 $Y=3.245
+ $X2=4.36 $Y2=3.33
r137 34 36 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=4.36 $Y=3.245
+ $X2=4.36 $Y2=2.79
r138 30 33 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=2.25 $Y=2.115
+ $X2=2.25 $Y2=2.815
r139 28 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.25 $Y=3.245
+ $X2=2.25 $Y2=3.33
r140 28 33 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.25 $Y=3.245
+ $X2=2.25 $Y2=2.815
r141 27 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.23 $Y2=3.33
r142 26 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=2.25 $Y2=3.33
r143 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=1.395 $Y2=3.33
r144 22 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=3.33
r145 22 24 33.5256 $w=3.28e-07 $l=9.6e-07 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=2.285
r146 18 21 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.24 $Y=1.985
+ $X2=0.24 $Y2=2.815
r147 16 72 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r148 16 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r149 5 40 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.825
+ $Y=1.96 $X2=6.97 $Y2=2.815
r150 4 36 600 $w=1.7e-07 $l=9.3795e-07 $layer=licon1_PDIFF $count=1 $X=4.175
+ $Y=1.94 $X2=4.36 $Y2=2.79
r151 3 33 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.115
+ $Y=1.84 $X2=2.25 $Y2=2.815
r152 3 30 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.115
+ $Y=1.84 $X2=2.25 $Y2=2.115
r153 2 24 300 $w=1.7e-07 $l=5.29481e-07 $layer=licon1_PDIFF $count=2 $X=1.045
+ $Y=1.84 $X2=1.23 $Y2=2.285
r154 1 21 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r155 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_4%X 1 2 3 4 13 15 16 19 25 27 29 33 39 42 45 48
+ 51
c73 42 0 1.30599e-19 $X=0.73 $Y=1.565
c74 27 0 3.54028e-20 $X=1.565 $Y=1.865
c75 15 0 1.0009e-19 $X=0.565 $Y=1.565
c76 13 0 8.40338e-20 $X=0.685 $Y=1.225
r77 48 51 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=1.225 $X2=0.24
+ $Y2=1.31
r78 48 51 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.24 $Y=1.345
+ $X2=0.24 $Y2=1.31
r79 45 46 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.85 $Y=1.025 $X2=0.85
+ $Y2=1.225
r80 42 44 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=0.73 $Y=1.565 $X2=0.73
+ $Y2=1.865
r81 41 48 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.24 $Y=1.48
+ $X2=0.24 $Y2=1.345
r82 37 39 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.85 $Y=0.94
+ $X2=1.85 $Y2=0.515
r83 33 35 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.73 $Y=1.985
+ $X2=1.73 $Y2=2.815
r84 31 33 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=1.73 $Y=1.95
+ $X2=1.73 $Y2=1.985
r85 30 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=1.025
+ $X2=0.85 $Y2=1.025
r86 29 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.685 $Y=1.025
+ $X2=1.85 $Y2=0.94
r87 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.685 $Y=1.025
+ $X2=1.015 $Y2=1.025
r88 28 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=1.865
+ $X2=0.73 $Y2=1.865
r89 27 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.565 $Y=1.865
+ $X2=1.73 $Y2=1.95
r90 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.565 $Y=1.865
+ $X2=0.895 $Y2=1.865
r91 23 45 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=0.94
+ $X2=0.85 $Y2=1.025
r92 23 25 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=0.85 $Y=0.94
+ $X2=0.85 $Y2=0.515
r93 19 21 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.73 $Y=1.985
+ $X2=0.73 $Y2=2.815
r94 17 44 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.95
+ $X2=0.73 $Y2=1.865
r95 17 19 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.73 $Y=1.95
+ $X2=0.73 $Y2=1.985
r96 16 41 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.565
+ $X2=0.24 $Y2=1.48
r97 15 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=1.565
+ $X2=0.73 $Y2=1.565
r98 15 16 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.565 $Y=1.565
+ $X2=0.355 $Y2=1.565
r99 14 48 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.355 $Y=1.225
+ $X2=0.24 $Y2=1.225
r100 13 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.685 $Y=1.225
+ $X2=0.85 $Y2=1.225
r101 13 14 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.685 $Y=1.225
+ $X2=0.355 $Y2=1.225
r102 4 35 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.84 $X2=1.73 $Y2=2.815
r103 4 33 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.84 $X2=1.73 $Y2=1.985
r104 3 21 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=2.815
r105 3 19 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.73 $Y2=1.985
r106 2 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.71
+ $Y=0.37 $X2=1.85 $Y2=0.515
r107 1 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.71
+ $Y=0.37 $X2=0.85 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_4%A_537_388# 1 2 11
r17 8 11 42.995 $w=2.58e-07 $l=9.7e-07 $layer=LI1_cond $X=2.89 $Y=2.83 $X2=3.86
+ $Y2=2.83
r18 2 11 600 $w=1.7e-07 $l=9.15014e-07 $layer=licon1_PDIFF $count=1 $X=3.725
+ $Y=1.94 $X2=3.86 $Y2=2.79
r19 1 8 600 $w=1.7e-07 $l=9.4194e-07 $layer=licon1_PDIFF $count=1 $X=2.685
+ $Y=1.94 $X2=2.89 $Y2=2.785
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_4%A_961_392# 1 2 3 10 17 18 19 22 26 28
r51 24 28 3.10218 $w=3.05e-07 $l=9.66954e-08 $layer=LI1_cond $X=7.905 $Y=2.39
+ $X2=7.88 $Y2=2.475
r52 24 26 11.3186 $w=2.78e-07 $l=2.75e-07 $layer=LI1_cond $X=7.905 $Y=2.39
+ $X2=7.905 $Y2=2.115
r53 20 28 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.88 $Y=2.56
+ $X2=7.88 $Y2=2.475
r54 20 22 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=7.88 $Y=2.56
+ $X2=7.88 $Y2=2.815
r55 18 28 3.51065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.715 $Y=2.475
+ $X2=7.88 $Y2=2.475
r56 18 19 95.9037 $w=1.68e-07 $l=1.47e-06 $layer=LI1_cond $X=7.715 $Y=2.475
+ $X2=6.245 $Y2=2.475
r57 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.16 $Y=2.56
+ $X2=6.245 $Y2=2.475
r58 16 17 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.16 $Y=2.56
+ $X2=6.16 $Y2=2.7
r59 12 15 37.866 $w=2.78e-07 $l=9.2e-07 $layer=LI1_cond $X=4.95 $Y=2.84 $X2=5.87
+ $Y2=2.84
r60 10 17 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=6.075 $Y=2.84
+ $X2=6.16 $Y2=2.7
r61 10 15 8.43753 $w=2.78e-07 $l=2.05e-07 $layer=LI1_cond $X=6.075 $Y=2.84
+ $X2=5.87 $Y2=2.84
r62 3 26 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=7.745
+ $Y=1.96 $X2=7.88 $Y2=2.115
r63 3 22 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.745
+ $Y=1.96 $X2=7.88 $Y2=2.815
r64 2 15 600 $w=1.7e-07 $l=9.04986e-07 $layer=licon1_PDIFF $count=1 $X=5.735
+ $Y=1.96 $X2=5.87 $Y2=2.8
r65 1 12 600 $w=1.7e-07 $l=9.09615e-07 $layer=licon1_PDIFF $count=1 $X=4.805
+ $Y=1.96 $X2=4.95 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_4%A_1237_392# 1 2 7 13 15 16
c21 15 0 8.99845e-20 $X=7.43 $Y=2.115
c22 13 0 8.94372e-20 $X=6.675 $Y=2.095
r23 15 16 7.69997 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=7.43 $Y=2.075
+ $X2=7.265 $Y2=2.075
r24 13 16 29.5627 $w=2.28e-07 $l=5.9e-07 $layer=LI1_cond $X=6.675 $Y=2.085
+ $X2=7.265 $Y2=2.085
r25 7 13 5.85606 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.55 $Y=2.095
+ $X2=6.675 $Y2=2.095
r26 7 9 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=6.55 $Y=2.095
+ $X2=6.415 $Y2=2.095
r27 2 15 600 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=7.295
+ $Y=1.96 $X2=7.43 $Y2=2.115
r28 1 9 600 $w=1.7e-07 $l=3.05205e-07 $layer=licon1_PDIFF $count=1 $X=6.185
+ $Y=1.96 $X2=6.415 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_4%VGND 1 2 3 4 5 6 19 21 23 27 31 35 39 43 46
+ 47 49 50 52 53 54 69 75 76 82 85
r107 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r108 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r109 80 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r110 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r111 76 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r112 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r113 73 85 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=7.545 $Y=0
+ $X2=7.352 $Y2=0
r114 73 75 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.545 $Y=0
+ $X2=7.92 $Y2=0
r115 72 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r116 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r117 69 85 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=7.16 $Y=0 $X2=7.352
+ $Y2=0
r118 69 71 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=7.16 $Y=0 $X2=6.96
+ $Y2=0
r119 68 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r120 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r121 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r122 64 65 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r123 61 64 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=5.04
+ $Y2=0
r124 61 62 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r125 59 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r126 59 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r127 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r128 56 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=0 $X2=1.35
+ $Y2=0
r129 56 58 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.515 $Y=0
+ $X2=2.16 $Y2=0
r130 54 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r131 54 62 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=2.64 $Y2=0
r132 52 67 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.23 $Y=0 $X2=6
+ $Y2=0
r133 52 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.23 $Y=0 $X2=6.395
+ $Y2=0
r134 51 71 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=6.56 $Y=0 $X2=6.96
+ $Y2=0
r135 51 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.56 $Y=0 $X2=6.395
+ $Y2=0
r136 49 64 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.23 $Y=0 $X2=5.04
+ $Y2=0
r137 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.23 $Y=0 $X2=5.395
+ $Y2=0
r138 48 67 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.56 $Y=0 $X2=6
+ $Y2=0
r139 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.56 $Y=0 $X2=5.395
+ $Y2=0
r140 46 58 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.24 $Y=0 $X2=2.16
+ $Y2=0
r141 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=0 $X2=2.405
+ $Y2=0
r142 45 61 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.57 $Y=0 $X2=2.64
+ $Y2=0
r143 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.57 $Y=0 $X2=2.405
+ $Y2=0
r144 41 85 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=7.352 $Y=0.085
+ $X2=7.352 $Y2=0
r145 41 43 12.8714 $w=3.83e-07 $l=4.3e-07 $layer=LI1_cond $X=7.352 $Y=0.085
+ $X2=7.352 $Y2=0.515
r146 37 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.395 $Y=0.085
+ $X2=6.395 $Y2=0
r147 37 39 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=6.395 $Y=0.085
+ $X2=6.395 $Y2=0.52
r148 33 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=0.085
+ $X2=5.395 $Y2=0
r149 33 35 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=5.395 $Y=0.085
+ $X2=5.395 $Y2=0.525
r150 29 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.405 $Y=0.085
+ $X2=2.405 $Y2=0
r151 29 31 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.405 $Y=0.085
+ $X2=2.405 $Y2=0.515
r152 25 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.35 $Y=0.085
+ $X2=1.35 $Y2=0
r153 25 27 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=1.35 $Y=0.085
+ $X2=1.35 $Y2=0.56
r154 24 79 4.59558 $w=1.7e-07 $l=2.58e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.257 $Y2=0
r155 23 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.185 $Y=0 $X2=1.35
+ $Y2=0
r156 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.185 $Y=0
+ $X2=0.515 $Y2=0
r157 19 79 3.17059 $w=3.3e-07 $l=1.28662e-07 $layer=LI1_cond $X=0.35 $Y=0.085
+ $X2=0.257 $Y2=0
r158 19 21 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.35 $Y=0.085
+ $X2=0.35 $Y2=0.515
r159 6 43 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=7.115
+ $Y=0.37 $X2=7.35 $Y2=0.515
r160 5 39 182 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_NDIFF $count=1 $X=6.185
+ $Y=0.37 $X2=6.395 $Y2=0.52
r161 4 35 182 $w=1.7e-07 $l=2.45561e-07 $layer=licon1_NDIFF $count=1 $X=5.215
+ $Y=0.37 $X2=5.395 $Y2=0.525
r162 3 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.265
+ $Y=0.37 $X2=2.405 $Y2=0.515
r163 2 27 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=1.14
+ $Y=0.37 $X2=1.35 $Y2=0.56
r164 1 21 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.205
+ $Y=0.37 $X2=0.35 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O32A_4%A_564_74# 1 2 3 4 5 6 21 23 24 27 29 32 35 39
+ 41 45 47 51 53 56 58
c99 56 0 7.70569e-20 $X=5.895 $Y=0.87
c100 45 0 1.44963e-19 $X=6.825 $Y=0.515
r101 49 51 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=7.88 $Y=0.78
+ $X2=7.88 $Y2=0.515
r102 48 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.99 $Y=0.865
+ $X2=6.865 $Y2=0.865
r103 47 49 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.715 $Y=0.865
+ $X2=7.88 $Y2=0.78
r104 47 48 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=7.715 $Y=0.865
+ $X2=6.99 $Y2=0.865
r105 43 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.865 $Y=0.78
+ $X2=6.865 $Y2=0.865
r106 43 45 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=6.865 $Y=0.78
+ $X2=6.865 $Y2=0.515
r107 42 56 8.61065 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=6.06 $Y=0.865
+ $X2=5.895 $Y2=0.87
r108 41 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.74 $Y=0.865
+ $X2=6.865 $Y2=0.865
r109 41 42 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.74 $Y=0.865
+ $X2=6.06 $Y2=0.865
r110 37 56 0.89609 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=5.895 $Y=0.78
+ $X2=5.895 $Y2=0.87
r111 37 39 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=5.895 $Y=0.78
+ $X2=5.895 $Y2=0.515
r112 36 55 4.91858 $w=1.7e-07 $l=1.77059e-07 $layer=LI1_cond $X=5.06 $Y=0.875
+ $X2=4.895 $Y2=0.9
r113 35 56 8.61065 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=5.73 $Y=0.875
+ $X2=5.895 $Y2=0.87
r114 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.73 $Y=0.875
+ $X2=5.06 $Y2=0.875
r115 32 55 2.8476 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.895 $Y=0.79
+ $X2=4.895 $Y2=0.9
r116 32 34 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.895 $Y=0.79
+ $X2=4.895 $Y2=0.515
r117 31 34 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.895 $Y=0.425
+ $X2=4.895 $Y2=0.515
r118 30 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.06 $Y=0.34
+ $X2=3.895 $Y2=0.34
r119 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.73 $Y=0.34
+ $X2=4.895 $Y2=0.425
r120 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.73 $Y=0.34
+ $X2=4.06 $Y2=0.34
r121 25 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.895 $Y=0.425
+ $X2=3.895 $Y2=0.34
r122 25 27 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.895 $Y=0.425
+ $X2=3.895 $Y2=0.595
r123 23 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.73 $Y=0.34
+ $X2=3.895 $Y2=0.34
r124 23 24 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.73 $Y=0.34 $X2=3.13
+ $Y2=0.34
r125 19 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.965 $Y=0.425
+ $X2=3.13 $Y2=0.34
r126 19 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.965 $Y=0.425
+ $X2=2.965 $Y2=0.515
r127 6 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.74
+ $Y=0.37 $X2=7.88 $Y2=0.515
r128 5 58 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=6.685
+ $Y=0.37 $X2=6.825 $Y2=0.865
r129 5 45 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.685
+ $Y=0.37 $X2=6.825 $Y2=0.515
r130 4 39 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=5.735
+ $Y=0.37 $X2=5.895 $Y2=0.515
r131 3 55 182 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_NDIFF $count=1 $X=4.685
+ $Y=0.37 $X2=4.895 $Y2=0.885
r132 3 34 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=4.685
+ $Y=0.37 $X2=4.895 $Y2=0.515
r133 2 27 182 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_NDIFF $count=1 $X=3.685
+ $Y=0.37 $X2=3.895 $Y2=0.595
r134 1 21 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=2.82
+ $Y=0.37 $X2=2.965 $Y2=0.515
.ends


* File: sky130_fd_sc_ms__dfsbp_1.pex.spice
* Created: Fri Aug 28 17:23:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DFSBP_1%D 2 5 9 11 12 16 17 20
c32 17 0 1.1887e-19 $X=0.64 $Y=1.175
r33 20 22 39.7991 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.855
+ $X2=0.61 $Y2=2.02
r34 20 21 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.855 $X2=0.64 $Y2=1.855
r35 16 18 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.175
+ $X2=0.61 $Y2=1.01
r36 16 17 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.175 $X2=0.64 $Y2=1.175
r37 12 21 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=0.64 $Y=1.665
+ $X2=0.64 $Y2=1.855
r38 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.665
r39 11 17 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.175
r40 9 18 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.495 $Y=0.61 $X2=0.495
+ $Y2=1.01
r41 5 22 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=0.505 $Y=2.75
+ $X2=0.505 $Y2=2.02
r42 2 20 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=0.61 $Y=1.825 $X2=0.61
+ $Y2=1.855
r43 1 16 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=0.61 $Y=1.205 $X2=0.61
+ $Y2=1.175
r44 1 2 88.4142 $w=3.9e-07 $l=6.2e-07 $layer=POLY_cond $X=0.61 $Y=1.205 $X2=0.61
+ $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_1%CLK 3 6 8 11 13
c38 11 0 3.27893e-19 $X=1.465 $Y=1.385
c39 6 0 1.1887e-19 $X=1.515 $Y=2.35
r40 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.385
+ $X2=1.465 $Y2=1.55
r41 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.385
+ $X2=1.465 $Y2=1.22
r42 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.465
+ $Y=1.385 $X2=1.465 $Y2=1.385
r43 8 12 6.69663 $w=3.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=1.465 $Y2=1.365
r44 6 14 310.968 $w=1.8e-07 $l=8e-07 $layer=POLY_cond $X=1.515 $Y=2.35 $X2=1.515
+ $Y2=1.55
r45 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.485 $Y=0.74
+ $X2=1.485 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_1%A_398_74# 1 2 7 8 11 17 21 24 26 29 33 35 36
+ 37 38 41 48 49 52 53 56 57 58 60 61 62 64 65 66 68 70 71 72 75 76 80 81 84 85
+ 86 90 94
c291 84 0 1.22752e-19 $X=7.395 $Y=2.185
c292 66 0 2.3488e-20 $X=6.035 $Y=1.705
c293 65 0 1.57368e-19 $X=6.435 $Y=1.705
c294 62 0 1.42192e-19 $X=5.54 $Y=2.21
c295 35 0 8.72473e-20 $X=3.025 $Y=0.34
c296 26 0 1.32821e-19 $X=3.03 $Y=2.105
r297 89 90 16.2455 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.665 $Y=1.525
+ $X2=3.59 $Y2=1.525
r298 85 97 17.8806 $w=3.1e-07 $l=1.15e-07 $layer=POLY_cond $X=7.395 $Y=2.185
+ $X2=7.51 $Y2=2.185
r299 84 86 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.395 $Y=2.185
+ $X2=7.395 $Y2=2.02
r300 84 85 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.395
+ $Y=2.185 $X2=7.395 $Y2=2.185
r301 81 94 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.715 $Y=1.285
+ $X2=6.715 $Y2=1.12
r302 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.715
+ $Y=1.285 $X2=6.715 $Y2=1.285
r303 77 80 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=6.52 $Y=1.285
+ $X2=6.715 $Y2=1.285
r304 73 86 104.059 $w=1.68e-07 $l=1.595e-06 $layer=LI1_cond $X=7.475 $Y=0.425
+ $X2=7.475 $Y2=2.02
r305 71 73 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.39 $Y=0.34
+ $X2=7.475 $Y2=0.425
r306 71 72 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=7.39 $Y=0.34
+ $X2=6.605 $Y2=0.34
r307 69 77 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.52 $Y=1.45
+ $X2=6.52 $Y2=1.285
r308 69 70 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.52 $Y=1.45
+ $X2=6.52 $Y2=1.62
r309 68 77 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.52 $Y=1.12
+ $X2=6.52 $Y2=1.285
r310 67 72 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.52 $Y=0.425
+ $X2=6.605 $Y2=0.34
r311 67 68 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.52 $Y=0.425
+ $X2=6.52 $Y2=1.12
r312 65 70 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.435 $Y=1.705
+ $X2=6.52 $Y2=1.62
r313 65 66 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=6.435 $Y=1.705
+ $X2=6.035 $Y2=1.705
r314 63 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.95 $Y=1.79
+ $X2=6.035 $Y2=1.705
r315 63 64 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.95 $Y=1.79
+ $X2=5.95 $Y2=2.125
r316 61 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.865 $Y=2.21
+ $X2=5.95 $Y2=2.125
r317 61 62 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.865 $Y=2.21
+ $X2=5.54 $Y2=2.21
r318 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.455 $Y=2.295
+ $X2=5.54 $Y2=2.21
r319 59 60 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.455 $Y=2.295
+ $X2=5.455 $Y2=2.905
r320 57 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.37 $Y=2.99
+ $X2=5.455 $Y2=2.905
r321 57 58 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.37 $Y=2.99
+ $X2=4.78 $Y2=2.99
r322 56 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.695 $Y=2.905
+ $X2=4.78 $Y2=2.99
r323 55 56 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.695 $Y=2.335
+ $X2=4.695 $Y2=2.905
r324 54 76 2.0246 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.945 $Y=2.25
+ $X2=3.825 $Y2=2.25
r325 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.61 $Y=2.25
+ $X2=4.695 $Y2=2.335
r326 53 54 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.61 $Y=2.25
+ $X2=3.945 $Y2=2.25
r327 51 76 4.40882 $w=2.05e-07 $l=1.00995e-07 $layer=LI1_cond $X=3.79 $Y=2.335
+ $X2=3.825 $Y2=2.25
r328 51 52 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.79 $Y=2.335
+ $X2=3.79 $Y2=2.905
r329 49 89 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=3.825 $Y=1.525
+ $X2=3.665 $Y2=1.525
r330 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.825
+ $Y=1.525 $X2=3.825 $Y2=1.525
r331 46 76 4.40882 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.825 $Y=2.165
+ $X2=3.825 $Y2=2.25
r332 46 48 30.7318 $w=2.38e-07 $l=6.4e-07 $layer=LI1_cond $X=3.825 $Y=2.165
+ $X2=3.825 $Y2=1.525
r333 44 75 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.11 $Y=0.425
+ $X2=3.11 $Y2=1.435
r334 41 75 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.03 $Y=1.6
+ $X2=3.03 $Y2=1.435
r335 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.03
+ $Y=1.6 $X2=3.03 $Y2=1.6
r336 37 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.705 $Y=2.99
+ $X2=3.79 $Y2=2.905
r337 37 38 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=3.705 $Y=2.99
+ $X2=2.355 $Y2=2.99
r338 35 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.025 $Y=0.34
+ $X2=3.11 $Y2=0.425
r339 35 36 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.025 $Y=0.34
+ $X2=2.295 $Y2=0.34
r340 31 38 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.23 $Y=2.905
+ $X2=2.355 $Y2=2.99
r341 31 33 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=2.23 $Y=2.905
+ $X2=2.23 $Y2=2.565
r342 27 36 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.17 $Y=0.425
+ $X2=2.295 $Y2=0.34
r343 27 29 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=2.17 $Y=0.425
+ $X2=2.17 $Y2=0.515
r344 22 97 15.4789 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.51 $Y=2.35
+ $X2=7.51 $Y2=2.185
r345 22 24 155.484 $w=1.8e-07 $l=4e-07 $layer=POLY_cond $X=7.51 $Y=2.35 $X2=7.51
+ $Y2=2.75
r346 21 94 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.725 $Y=0.69
+ $X2=6.725 $Y2=1.12
r347 15 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.665 $Y=1.36
+ $X2=3.665 $Y2=1.525
r348 15 17 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=3.665 $Y=1.36
+ $X2=3.665 $Y2=0.615
r349 14 42 15.4923 $w=2.55e-07 $l=1.65e-07 $layer=POLY_cond $X=3.195 $Y=1.562
+ $X2=3.03 $Y2=1.562
r350 14 90 96.2149 $w=2.55e-07 $l=3.95e-07 $layer=POLY_cond $X=3.195 $Y=1.562
+ $X2=3.59 $Y2=1.562
r351 11 26 163.258 $w=1.8e-07 $l=4.2e-07 $layer=POLY_cond $X=3.065 $Y=2.525
+ $X2=3.065 $Y2=2.105
r352 8 26 36.5727 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.03 $Y=1.94
+ $X2=3.03 $Y2=2.105
r353 7 42 12.0182 $w=3.3e-07 $l=1.28e-07 $layer=POLY_cond $X=3.03 $Y=1.69
+ $X2=3.03 $Y2=1.562
r354 7 8 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.03 $Y=1.69 $X2=3.03
+ $Y2=1.94
r355 2 33 600 $w=1.7e-07 $l=8.39792e-07 $layer=licon1_PDIFF $count=1 $X=2.055
+ $Y=1.79 $X2=2.19 $Y2=2.565
r356 1 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.99
+ $Y=0.37 $X2=2.13 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_1%A_779_380# 1 2 9 11 13 14 15 16 17 20 23 27
+ 30 35 38
c87 35 0 9.58642e-20 $X=4.395 $Y=1.72
c88 20 0 1.31064e-19 $X=4.95 $Y=1.885
c89 9 0 1.14714e-19 $X=3.985 $Y=2.525
r90 35 41 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.485 $Y=1.72
+ $X2=4.485 $Y2=1.265
r91 33 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.575 $Y=1.1
+ $X2=4.575 $Y2=1.265
r92 33 38 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.575 $Y=1.1 $X2=4.575
+ $Y2=1.01
r93 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.575
+ $Y=1.1 $X2=4.575 $Y2=1.1
r94 30 32 13.3188 $w=4.58e-07 $l=6.09098e-07 $layer=LI1_cond $X=4.817 $Y=0.6
+ $X2=4.575 $Y2=1.1
r95 25 27 23.9708 $w=2.48e-07 $l=5.2e-07 $layer=LI1_cond $X=5.075 $Y=1.995
+ $X2=5.075 $Y2=2.515
r96 23 36 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.395 $Y=1.885
+ $X2=4.395 $Y2=1.975
r97 23 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.395 $Y=1.885
+ $X2=4.395 $Y2=1.72
r98 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.395
+ $Y=1.885 $X2=4.395 $Y2=1.885
r99 20 25 6.85268 $w=2.2e-07 $l=1.71391e-07 $layer=LI1_cond $X=4.95 $Y=1.885
+ $X2=5.075 $Y2=1.995
r100 20 22 29.073 $w=2.18e-07 $l=5.55e-07 $layer=LI1_cond $X=4.95 $Y=1.885
+ $X2=4.395 $Y2=1.885
r101 16 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.41 $Y=1.01
+ $X2=4.575 $Y2=1.01
r102 16 17 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.41 $Y=1.01
+ $X2=4.13 $Y2=1.01
r103 14 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.23 $Y=1.975
+ $X2=4.395 $Y2=1.975
r104 14 15 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=4.23 $Y=1.975
+ $X2=4.075 $Y2=1.975
r105 11 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.055 $Y=0.935
+ $X2=4.13 $Y2=1.01
r106 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.055 $Y=0.935
+ $X2=4.055 $Y2=0.615
r107 7 15 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.985 $Y=2.05
+ $X2=4.075 $Y2=1.975
r108 7 9 184.637 $w=1.8e-07 $l=4.75e-07 $layer=POLY_cond $X=3.985 $Y=2.05
+ $X2=3.985 $Y2=2.525
r109 2 27 600 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_PDIFF $count=1 $X=4.98
+ $Y=2.315 $X2=5.115 $Y2=2.515
r110 1 30 182 $w=1.7e-07 $l=2.85745e-07 $layer=licon1_NDIFF $count=1 $X=4.89
+ $Y=0.37 $X2=5.015 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_1%A_596_81# 1 2 9 12 15 19 23 26 30 34 37 38
+ 39 40 41 42 45 46 48 52 56 61 64
c158 46 0 1.14714e-19 $X=3.355 $Y=2.295
c159 45 0 1.32821e-19 $X=3.34 $Y=2.515
c160 40 0 9.58642e-20 $X=5.092 $Y=1.29
c161 12 0 1.19393e-19 $X=5.025 $Y=1.57
c162 9 0 1.42192e-19 $X=4.89 $Y=2.525
r163 56 65 39.5669 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=6.122 $Y=1.285
+ $X2=6.122 $Y2=1.45
r164 56 64 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=6.122 $Y=1.285
+ $X2=6.122 $Y2=1.12
r165 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.1
+ $Y=1.285 $X2=6.1 $Y2=1.285
r166 52 55 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=6.1 $Y=1.205 $X2=6.1
+ $Y2=1.285
r167 51 61 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=5.115 $Y=1.22
+ $X2=5.23 $Y2=1.22
r168 51 58 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.115 $Y=1.22
+ $X2=5.025 $Y2=1.22
r169 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.115
+ $Y=1.22 $X2=5.115 $Y2=1.22
r170 45 46 10.2717 $w=3.58e-07 $l=2.2e-07 $layer=LI1_cond $X=3.355 $Y=2.515
+ $X2=3.355 $Y2=2.295
r171 43 50 4.42914 $w=1.7e-07 $l=1.58644e-07 $layer=LI1_cond $X=5.235 $Y=1.205
+ $X2=5.092 $Y2=1.172
r172 42 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.935 $Y=1.205
+ $X2=6.1 $Y2=1.205
r173 42 43 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=5.935 $Y=1.205
+ $X2=5.235 $Y2=1.205
r174 40 50 2.96953 $w=2.85e-07 $l=1.18e-07 $layer=LI1_cond $X=5.092 $Y=1.29
+ $X2=5.092 $Y2=1.172
r175 40 41 5.86331 $w=2.83e-07 $l=1.45e-07 $layer=LI1_cond $X=5.092 $Y=1.29
+ $X2=5.092 $Y2=1.435
r176 38 41 7.39867 $w=1.7e-07 $l=1.79538e-07 $layer=LI1_cond $X=4.95 $Y=1.52
+ $X2=5.092 $Y2=1.435
r177 38 39 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.95 $Y=1.52
+ $X2=4.285 $Y2=1.52
r178 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.2 $Y=1.435
+ $X2=4.285 $Y2=1.52
r179 36 37 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.2 $Y=1.055
+ $X2=4.2 $Y2=1.435
r180 35 48 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.615 $Y=0.97
+ $X2=3.49 $Y2=0.97
r181 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.115 $Y=0.97
+ $X2=4.2 $Y2=1.055
r182 34 35 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=4.115 $Y=0.97
+ $X2=3.615 $Y2=0.97
r183 32 48 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=3.45 $Y=1.055
+ $X2=3.49 $Y2=0.97
r184 32 46 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=3.45 $Y=1.055
+ $X2=3.45 $Y2=2.295
r185 28 48 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.49 $Y=0.885
+ $X2=3.49 $Y2=0.97
r186 28 30 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=3.49 $Y=0.885
+ $X2=3.49 $Y2=0.615
r187 23 64 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.235 $Y=0.69
+ $X2=6.235 $Y2=1.12
r188 19 65 293.476 $w=1.8e-07 $l=7.55e-07 $layer=POLY_cond $X=6.195 $Y=2.205
+ $X2=6.195 $Y2=1.45
r189 13 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.23 $Y=1.055
+ $X2=5.23 $Y2=1.22
r190 13 15 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=5.23 $Y=1.055
+ $X2=5.23 $Y2=0.58
r191 12 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.025 $Y=1.57
+ $X2=5.025 $Y2=1.645
r192 11 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.025 $Y=1.385
+ $X2=5.025 $Y2=1.22
r193 11 12 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=5.025 $Y=1.385
+ $X2=5.025 $Y2=1.57
r194 7 26 69.2234 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.89 $Y=1.645
+ $X2=5.025 $Y2=1.645
r195 7 9 312.911 $w=1.8e-07 $l=8.05e-07 $layer=POLY_cond $X=4.89 $Y=1.72
+ $X2=4.89 $Y2=2.525
r196 2 45 600 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_PDIFF $count=1 $X=3.155
+ $Y=2.315 $X2=3.34 $Y2=2.515
r197 1 30 182 $w=1.7e-07 $l=5.65332e-07 $layer=licon1_NDIFF $count=1 $X=2.98
+ $Y=0.405 $X2=3.45 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_1%SET_B 3 7 11 13 14 17 21 22 23 24 27 29 36
+ 38 42
c146 27 0 1.19393e-19 $X=5.52 $Y=1.665
c147 24 0 1.31064e-19 $X=5.665 $Y=1.665
c148 23 0 1.03271e-19 $X=8.255 $Y=1.665
c149 14 0 2.58188e-20 $X=8.09 $Y=1.3
r150 42 50 8.23174 $w=3.83e-07 $l=2.75e-07 $layer=LI1_cond $X=8.477 $Y=1.39
+ $X2=8.477 $Y2=1.665
r151 41 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.505 $Y=1.39
+ $X2=8.505 $Y2=1.555
r152 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.505
+ $Y=1.39 $X2=8.505 $Y2=1.39
r153 38 41 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.505 $Y=1.3
+ $X2=8.505 $Y2=1.39
r154 34 36 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.53 $Y=1.79 $X2=5.62
+ $Y2=1.79
r155 31 34 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=5.4 $Y=1.79 $X2=5.53
+ $Y2=1.79
r156 29 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=1.665
+ $X2=8.4 $Y2=1.665
r157 27 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.53
+ $Y=1.79 $X2=5.53 $Y2=1.79
r158 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.665
+ $X2=5.52 $Y2=1.665
r159 24 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=1.665
+ $X2=5.52 $Y2=1.665
r160 23 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=8.4 $Y2=1.665
r161 23 24 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=5.665 $Y2=1.665
r162 21 22 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=8.39 $Y=2.155
+ $X2=8.39 $Y2=2.305
r163 21 43 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=8.415 $Y=2.155
+ $X2=8.415 $Y2=1.555
r164 17 22 172.976 $w=1.8e-07 $l=4.45e-07 $layer=POLY_cond $X=8.38 $Y=2.75
+ $X2=8.38 $Y2=2.305
r165 13 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.34 $Y=1.3
+ $X2=8.505 $Y2=1.3
r166 13 14 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=8.34 $Y=1.3
+ $X2=8.09 $Y2=1.3
r167 9 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.015 $Y=1.225
+ $X2=8.09 $Y2=1.3
r168 9 11 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=8.015 $Y=1.225
+ $X2=8.015 $Y2=0.58
r169 5 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.62 $Y=1.625
+ $X2=5.62 $Y2=1.79
r170 5 7 535.84 $w=1.5e-07 $l=1.045e-06 $layer=POLY_cond $X=5.62 $Y=1.625
+ $X2=5.62 $Y2=0.58
r171 1 31 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.4 $Y=1.955
+ $X2=5.4 $Y2=1.79
r172 1 3 221.565 $w=1.8e-07 $l=5.7e-07 $layer=POLY_cond $X=5.4 $Y=1.955 $X2=5.4
+ $Y2=2.525
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_1%A_225_74# 1 2 9 13 16 17 19 20 23 27 29 34
+ 35 36 39 42 43 46 47 49 50 51 54 58 62 65
c171 58 0 1.8808e-19 $X=2.19 $Y=1.465
c172 54 0 2.99812e-20 $X=2.025 $Y=1.805
c173 39 0 1.57368e-19 $X=7.235 $Y=0.58
c174 34 0 1.22752e-19 $X=6.7 $Y=2.385
c175 27 0 1.25383e-19 $X=3.565 $Y=2.525
c176 17 0 8.72473e-20 $X=2.83 $Y=1.12
r177 62 64 17.8607 $w=4.58e-07 $l=4.95e-07 $layer=LI1_cond $X=1.205 $Y=0.515
+ $X2=1.205 $Y2=1.01
r178 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.19
+ $Y=1.465 $X2=2.19 $Y2=1.465
r179 56 58 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.19 $Y=1.72
+ $X2=2.19 $Y2=1.465
r180 54 56 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.025 $Y=1.805
+ $X2=2.19 $Y2=1.72
r181 54 65 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.025 $Y=1.805
+ $X2=1.455 $Y2=1.805
r182 51 53 5.57014 $w=2.98e-07 $l=1.45e-07 $layer=LI1_cond $X=1.145 $Y=1.87
+ $X2=1.29 $Y2=1.87
r183 50 65 7.90841 $w=2.98e-07 $l=1.5e-07 $layer=LI1_cond $X=1.305 $Y=1.87
+ $X2=1.455 $Y2=1.87
r184 50 53 0.576222 $w=2.98e-07 $l=1.5e-08 $layer=LI1_cond $X=1.305 $Y=1.87
+ $X2=1.29 $Y2=1.87
r185 49 51 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=1.06 $Y=1.72
+ $X2=1.145 $Y2=1.87
r186 49 64 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.06 $Y=1.72
+ $X2=1.06 $Y2=1.01
r187 46 59 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=2.41 $Y=1.465
+ $X2=2.19 $Y2=1.465
r188 43 46 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=2.485 $Y=1.12
+ $X2=2.485 $Y2=1.465
r189 41 59 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.055 $Y=1.465
+ $X2=2.19 $Y2=1.465
r190 41 42 3.90195 $w=3.3e-07 $l=2.85832e-07 $layer=POLY_cond $X=2.055 $Y=1.465
+ $X2=1.84 $Y2=1.3
r191 37 39 553.787 $w=1.5e-07 $l=1.08e-06 $layer=POLY_cond $X=7.235 $Y=1.66
+ $X2=7.235 $Y2=0.58
r192 35 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.16 $Y=1.735
+ $X2=7.235 $Y2=1.66
r193 35 36 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.16 $Y=1.735
+ $X2=6.79 $Y2=1.735
r194 32 34 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=6.7 $Y=3.075 $X2=6.7
+ $Y2=2.385
r195 31 36 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.7 $Y=1.81
+ $X2=6.79 $Y2=1.735
r196 31 34 223.508 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.7 $Y=1.81
+ $X2=6.7 $Y2=2.385
r197 30 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.655 $Y=3.15
+ $X2=3.565 $Y2=3.15
r198 29 32 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.61 $Y=3.15
+ $X2=6.7 $Y2=3.075
r199 29 30 1515.22 $w=1.5e-07 $l=2.955e-06 $layer=POLY_cond $X=6.61 $Y=3.15
+ $X2=3.655 $Y2=3.15
r200 25 47 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.565 $Y=3.075
+ $X2=3.565 $Y2=3.15
r201 25 27 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=3.565 $Y=3.075
+ $X2=3.565 $Y2=2.525
r202 21 23 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.905 $Y=1.045
+ $X2=2.905 $Y2=0.615
r203 19 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.475 $Y=3.15
+ $X2=3.565 $Y2=3.15
r204 19 20 469.181 $w=1.5e-07 $l=9.15e-07 $layer=POLY_cond $X=3.475 $Y=3.15
+ $X2=2.56 $Y2=3.15
r205 18 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.56 $Y=1.12
+ $X2=2.485 $Y2=1.12
r206 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.83 $Y=1.12
+ $X2=2.905 $Y2=1.045
r207 17 18 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.83 $Y=1.12
+ $X2=2.56 $Y2=1.12
r208 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.485 $Y=3.075
+ $X2=2.56 $Y2=3.15
r209 15 46 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.485 $Y=1.63
+ $X2=2.485 $Y2=1.465
r210 15 16 740.947 $w=1.5e-07 $l=1.445e-06 $layer=POLY_cond $X=2.485 $Y=1.63
+ $X2=2.485 $Y2=3.075
r211 11 42 34.7346 $w=1.65e-07 $l=3.87492e-07 $layer=POLY_cond $X=1.965 $Y=1.63
+ $X2=1.84 $Y2=1.3
r212 11 13 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.965 $Y=1.63
+ $X2=1.965 $Y2=2.35
r213 7 42 34.7346 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=1.915 $Y=1.3
+ $X2=1.84 $Y2=1.3
r214 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.915 $Y=1.3
+ $X2=1.915 $Y2=0.74
r215 2 53 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.79 $X2=1.29 $Y2=1.935
r216 1 62 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.125
+ $Y=0.37 $X2=1.27 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_1%A_1510_48# 1 2 9 13 17 20 21 24 28 30 32 33
+ 35 36 38
c116 38 0 7.00183e-20 $X=7.93 $Y=1.75
r117 34 35 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=9.65 $Y=1.01
+ $X2=9.65 $Y2=2.39
r118 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.565 $Y=2.475
+ $X2=9.65 $Y2=2.39
r119 32 33 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.565 $Y=2.475
+ $X2=9.33 $Y2=2.475
r120 31 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.255 $Y=0.925
+ $X2=9.09 $Y2=0.925
r121 30 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.565 $Y=0.925
+ $X2=9.65 $Y2=1.01
r122 30 31 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=9.565 $Y=0.925
+ $X2=9.255 $Y2=0.925
r123 26 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.165 $Y=2.56
+ $X2=9.33 $Y2=2.475
r124 26 28 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=9.165 $Y=2.56
+ $X2=9.165 $Y2=2.75
r125 22 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.09 $Y=0.84
+ $X2=9.09 $Y2=0.925
r126 22 24 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=9.09 $Y=0.84
+ $X2=9.09 $Y2=0.58
r127 20 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.925 $Y=0.925
+ $X2=9.09 $Y2=0.925
r128 20 21 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=8.925 $Y=0.925
+ $X2=8.1 $Y2=0.925
r129 18 38 0.934109 $w=2.58e-07 $l=5e-09 $layer=POLY_cond $X=7.935 $Y=1.75
+ $X2=7.93 $Y2=1.75
r130 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.935
+ $Y=1.75 $X2=7.935 $Y2=1.75
r131 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.935 $Y=1.01
+ $X2=8.1 $Y2=0.925
r132 15 17 25.8427 $w=3.28e-07 $l=7.4e-07 $layer=LI1_cond $X=7.935 $Y=1.01
+ $X2=7.935 $Y2=1.75
r133 11 38 11.2427 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.93 $Y=1.915
+ $X2=7.93 $Y2=1.75
r134 11 13 324.573 $w=1.8e-07 $l=8.35e-07 $layer=POLY_cond $X=7.93 $Y=1.915
+ $X2=7.93 $Y2=2.75
r135 7 38 56.9806 $w=2.58e-07 $l=3.78616e-07 $layer=POLY_cond $X=7.625 $Y=1.585
+ $X2=7.93 $Y2=1.75
r136 7 9 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=7.625 $Y=1.585
+ $X2=7.625 $Y2=0.58
r137 2 28 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=9.02
+ $Y=2.54 $X2=9.165 $Y2=2.75
r138 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.95
+ $Y=0.37 $X2=9.09 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_1%A_1358_377# 1 2 3 10 12 14 16 17 19 21 23 26
+ 28 29 32 38 41 43 44 45 49 50 51 53 56 60 62 64 66 69 74 78 79 80 81
c197 69 0 7.00183e-20 $X=6.885 $Y=1.882
c198 56 0 2.58188e-20 $X=8.44 $Y=2.265
c199 43 0 1.55237e-19 $X=10.925 $Y=1.41
r200 89 90 6.25673 $w=4e-07 $l=4.5e-08 $layer=POLY_cond $X=9.935 $Y=1.41
+ $X2=9.98 $Y2=1.41
r201 83 84 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=9.23
+ $Y=2.055 $X2=9.23 $Y2=2.055
r202 79 80 8.9189 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.73 $Y=2.35 $X2=7.9
+ $Y2=2.35
r203 78 79 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.45 $Y=2.565
+ $X2=7.73 $Y2=2.565
r204 77 78 8.76046 $w=4.23e-07 $l=1.65e-07 $layer=LI1_cond $X=7.285 $Y=2.692
+ $X2=7.45 $Y2=2.692
r205 72 74 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=6.94 $Y=0.76
+ $X2=7.135 $Y2=0.76
r206 67 85 12.5135 $w=4e-07 $l=9e-08 $layer=POLY_cond $X=9.23 $Y=1.41 $X2=9.14
+ $Y2=1.41
r207 66 67 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=9.23
+ $Y=1.375 $X2=9.23 $Y2=1.375
r208 64 83 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.23 $Y=2.05 $X2=9.23
+ $Y2=2.135
r209 64 66 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=9.23 $Y=2.05
+ $X2=9.23 $Y2=1.375
r210 63 81 5.58832 $w=3e-07 $l=2.20624e-07 $layer=LI1_cond $X=8.77 $Y=2.135
+ $X2=8.605 $Y2=2.265
r211 62 83 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.065 $Y=2.135
+ $X2=9.23 $Y2=2.135
r212 62 63 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.065 $Y=2.135
+ $X2=8.77 $Y2=2.135
r213 58 81 1.0017 $w=3.3e-07 $l=2.15e-07 $layer=LI1_cond $X=8.605 $Y=2.48
+ $X2=8.605 $Y2=2.265
r214 58 60 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=8.605 $Y=2.48
+ $X2=8.605 $Y2=2.75
r215 56 81 5.58832 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=8.44 $Y=2.265
+ $X2=8.605 $Y2=2.265
r216 56 80 14.4725 $w=4.28e-07 $l=5.4e-07 $layer=LI1_cond $X=8.44 $Y=2.265
+ $X2=7.9 $Y2=2.265
r217 53 69 12.249 $w=2.49e-07 $l=3.36155e-07 $layer=LI1_cond $X=7.135 $Y=1.68
+ $X2=6.885 $Y2=1.882
r218 52 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.135 $Y=0.925
+ $X2=7.135 $Y2=0.76
r219 52 53 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=7.135 $Y=0.925
+ $X2=7.135 $Y2=1.68
r220 50 77 1.27447 $w=4.23e-07 $l=4.7e-08 $layer=LI1_cond $X=7.238 $Y=2.692
+ $X2=7.285 $Y2=2.692
r221 50 51 6.18252 $w=4.23e-07 $l=2.28e-07 $layer=LI1_cond $X=7.238 $Y=2.692
+ $X2=7.01 $Y2=2.692
r222 47 51 7.42997 $w=4.25e-07 $l=2.6729e-07 $layer=LI1_cond $X=6.885 $Y=2.48
+ $X2=7.01 $Y2=2.692
r223 47 49 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=6.885 $Y=2.48
+ $X2=6.885 $Y2=2.26
r224 46 69 0.692029 $w=2.5e-07 $l=2.03e-07 $layer=LI1_cond $X=6.885 $Y=2.085
+ $X2=6.885 $Y2=1.882
r225 46 49 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=6.885 $Y=2.085
+ $X2=6.885 $Y2=2.26
r226 44 45 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=10.965 $Y=1.79
+ $X2=10.965 $Y2=1.94
r227 39 41 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=8.875 $Y=0.94
+ $X2=9.14 $Y2=0.94
r228 38 45 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=10.99 $Y=2.435
+ $X2=10.99 $Y2=1.94
r229 34 43 42.0026 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=10.925 $Y=1.61
+ $X2=10.925 $Y2=1.41
r230 34 44 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=10.925 $Y=1.61
+ $X2=10.925 $Y2=1.79
r231 30 43 42.0026 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=10.925 $Y=1.21
+ $X2=10.925 $Y2=1.41
r232 30 32 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=10.925 $Y=1.21
+ $X2=10.925 $Y2=0.645
r233 29 90 12.5135 $w=4e-07 $l=9e-08 $layer=POLY_cond $X=10.07 $Y=1.41 $X2=9.98
+ $Y2=1.41
r234 28 43 7.17539 $w=4e-07 $l=7.5e-08 $layer=POLY_cond $X=10.85 $Y=1.41
+ $X2=10.925 $Y2=1.41
r235 28 29 108.45 $w=4e-07 $l=7.8e-07 $layer=POLY_cond $X=10.85 $Y=1.41
+ $X2=10.07 $Y2=1.41
r236 24 90 21.4623 $w=1.8e-07 $l=2e-07 $layer=POLY_cond $X=9.98 $Y=1.61 $X2=9.98
+ $Y2=1.41
r237 24 26 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=9.98 $Y=1.61
+ $X2=9.98 $Y2=2.4
r238 21 89 25.8619 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=9.935 $Y=1.21
+ $X2=9.935 $Y2=1.41
r239 21 23 151.027 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=9.935 $Y=1.21
+ $X2=9.935 $Y2=0.74
r240 17 84 45.6296 $w=3.89e-07 $l=3.25308e-07 $layer=POLY_cond $X=9.475 $Y=2.31
+ $X2=9.315 $Y2=2.055
r241 17 19 171.032 $w=1.8e-07 $l=4.4e-07 $layer=POLY_cond $X=9.475 $Y=2.31
+ $X2=9.475 $Y2=2.75
r242 16 84 8.75288 $w=4.7e-07 $l=7.71362e-08 $layer=POLY_cond $X=9.3 $Y=1.985
+ $X2=9.315 $Y2=2.055
r243 15 89 88.2894 $w=4e-07 $l=6.35e-07 $layer=POLY_cond $X=9.3 $Y=1.41
+ $X2=9.935 $Y2=1.41
r244 15 67 9.73269 $w=4e-07 $l=7e-08 $layer=POLY_cond $X=9.3 $Y=1.41 $X2=9.23
+ $Y2=1.41
r245 15 16 44.374 $w=4.7e-07 $l=3.75e-07 $layer=POLY_cond $X=9.3 $Y=1.61 $X2=9.3
+ $Y2=1.985
r246 14 85 25.8619 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=9.14 $Y=1.21 $X2=9.14
+ $Y2=1.41
r247 13 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.14 $Y=1.015
+ $X2=9.14 $Y2=0.94
r248 13 14 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=9.14 $Y=1.015
+ $X2=9.14 $Y2=1.21
r249 10 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.875 $Y=0.865
+ $X2=8.875 $Y2=0.94
r250 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.875 $Y=0.865
+ $X2=8.875 $Y2=0.58
r251 3 60 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=8.47
+ $Y=2.54 $X2=8.605 $Y2=2.75
r252 2 77 300 $w=1.7e-07 $l=1.07436e-06 $layer=licon1_PDIFF $count=2 $X=6.79
+ $Y=1.885 $X2=7.285 $Y2=2.74
r253 2 49 600 $w=1.7e-07 $l=4.37321e-07 $layer=licon1_PDIFF $count=1 $X=6.79
+ $Y=1.885 $X2=6.925 $Y2=2.26
r254 1 72 182 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_NDIFF $count=1 $X=6.8
+ $Y=0.37 $X2=6.94 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_1%A_2113_74# 1 2 9 13 16 19 22 26 27 29 30 32
c56 19 0 1.55237e-19 $X=10.777 $Y=1.22
r57 27 33 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.42 $Y=1.385
+ $X2=11.42 $Y2=1.55
r58 27 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.42 $Y=1.385
+ $X2=11.42 $Y2=1.22
r59 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.42
+ $Y=1.385 $X2=11.42 $Y2=1.385
r60 24 30 0.674692 $w=3.3e-07 $l=9.8e-08 $layer=LI1_cond $X=10.875 $Y=1.385
+ $X2=10.777 $Y2=1.385
r61 24 26 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=10.875 $Y=1.385
+ $X2=11.42 $Y2=1.385
r62 20 30 8.18839 $w=1.82e-07 $l=1.70895e-07 $layer=LI1_cond $X=10.765 $Y=1.55
+ $X2=10.777 $Y2=1.385
r63 20 22 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=10.765 $Y=1.55
+ $X2=10.765 $Y2=2.16
r64 19 30 8.18839 $w=1.82e-07 $l=1.65e-07 $layer=LI1_cond $X=10.777 $Y=1.22
+ $X2=10.777 $Y2=1.385
r65 19 29 15.9254 $w=1.93e-07 $l=2.8e-07 $layer=LI1_cond $X=10.777 $Y=1.22
+ $X2=10.777 $Y2=0.94
r66 14 29 7.67512 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=10.71 $Y=0.775
+ $X2=10.71 $Y2=0.94
r67 14 16 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=10.71 $Y=0.775
+ $X2=10.71 $Y2=0.645
r68 13 32 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=11.505 $Y=0.74
+ $X2=11.505 $Y2=1.22
r69 9 33 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=11.495 $Y=2.4
+ $X2=11.495 $Y2=1.55
r70 2 22 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=10.62
+ $Y=2.015 $X2=10.765 $Y2=2.16
r71 1 16 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=10.565
+ $Y=0.37 $X2=10.71 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_1%A_27_80# 1 2 3 4 15 18 21 23 25 28 29 30 31
+ 36
c67 25 0 1.25383e-19 $X=2.525 $Y=2.145
r68 36 38 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=0.68
+ $X2=2.69 $Y2=0.845
r69 31 33 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.71 $Y=2.145
+ $X2=1.71 $Y2=2.275
r70 28 38 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=2.61 $Y=2.06
+ $X2=2.61 $Y2=0.845
r71 26 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=2.145
+ $X2=1.71 $Y2=2.145
r72 25 41 12.1344 $w=3.72e-07 $l=4.75079e-07 $layer=LI1_cond $X=2.525 $Y=2.145
+ $X2=2.765 $Y2=2.515
r73 25 28 6.42219 $w=3.72e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.525 $Y=2.145
+ $X2=2.61 $Y2=2.06
r74 25 26 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.525 $Y=2.145
+ $X2=1.795 $Y2=2.145
r75 24 30 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=2.275
+ $X2=0.24 $Y2=2.275
r76 23 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=2.275
+ $X2=1.71 $Y2=2.275
r77 23 24 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=1.625 $Y=2.275
+ $X2=0.365 $Y2=2.275
r78 19 30 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.36 $X2=0.24
+ $Y2=2.275
r79 19 21 17.9781 $w=2.48e-07 $l=3.9e-07 $layer=LI1_cond $X=0.24 $Y=2.36
+ $X2=0.24 $Y2=2.75
r80 18 30 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.2 $Y=2.19
+ $X2=0.24 $Y2=2.275
r81 18 29 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=0.2 $Y=2.19 $X2=0.2
+ $Y2=0.84
r82 13 29 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=0.715
+ $X2=0.24 $Y2=0.84
r83 13 15 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=0.24 $Y=0.715
+ $X2=0.24 $Y2=0.61
r84 4 41 600 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=2.695
+ $Y=2.315 $X2=2.84 $Y2=2.515
r85 3 21 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.28 $Y2=2.75
r86 2 36 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=2.545
+ $Y=0.405 $X2=2.69 $Y2=0.68
r87 1 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.4 $X2=0.28 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_1%VPWR 1 2 3 4 5 6 7 24 28 32 36 40 44 48 51
+ 52 53 55 60 65 70 82 89 96 97 100 103 106 109 112 115
c136 28 0 2.99812e-20 $X=1.74 $Y=2.695
c137 4 0 1.03271e-19 $X=5.49 $Y=2.315
r138 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r139 112 113 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r140 106 107 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r141 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r142 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r143 97 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=11.28 $Y2=3.33
r144 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r145 94 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.38 $Y=3.33
+ $X2=11.215 $Y2=3.33
r146 94 96 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=11.38 $Y=3.33
+ $X2=11.76 $Y2=3.33
r147 93 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r148 93 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=9.84 $Y2=3.33
r149 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r150 90 112 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=9.91 $Y=3.33
+ $X2=9.735 $Y2=3.33
r151 90 92 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=9.91 $Y=3.33
+ $X2=10.8 $Y2=3.33
r152 89 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.05 $Y=3.33
+ $X2=11.215 $Y2=3.33
r153 89 92 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=11.05 $Y=3.33
+ $X2=10.8 $Y2=3.33
r154 88 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r155 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r156 85 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r157 84 87 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.4 $Y=3.33 $X2=9.36
+ $Y2=3.33
r158 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r159 82 112 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=9.56 $Y=3.33
+ $X2=9.735 $Y2=3.33
r160 82 87 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=9.56 $Y=3.33 $X2=9.36
+ $Y2=3.33
r161 81 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r162 80 81 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r163 78 109 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.05 $Y=3.33
+ $X2=5.88 $Y2=3.33
r164 78 80 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=6.05 $Y=3.33 $X2=7.92
+ $Y2=3.33
r165 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r166 74 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r167 74 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r168 73 76 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r169 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r170 71 106 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=4.44 $Y=3.33
+ $X2=4.242 $Y2=3.33
r171 71 73 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.44 $Y=3.33
+ $X2=4.56 $Y2=3.33
r172 70 109 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.71 $Y=3.33
+ $X2=5.88 $Y2=3.33
r173 70 76 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.71 $Y=3.33
+ $X2=5.52 $Y2=3.33
r174 69 107 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r175 69 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r176 68 69 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r177 66 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=1.74 $Y2=3.33
r178 66 68 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=2.16 $Y2=3.33
r179 65 106 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=4.242 $Y2=3.33
r180 65 68 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=2.16 $Y2=3.33
r181 64 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r182 64 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r183 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r184 61 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r185 61 63 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r186 60 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.74 $Y2=3.33
r187 60 63 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.2 $Y2=3.33
r188 58 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r189 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r190 55 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r191 55 57 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r192 53 81 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=7.92 $Y2=3.33
r193 53 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r194 53 109 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r195 51 80 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=8.07 $Y=3.33
+ $X2=7.92 $Y2=3.33
r196 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.07 $Y=3.33
+ $X2=8.155 $Y2=3.33
r197 50 84 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=8.24 $Y=3.33
+ $X2=8.4 $Y2=3.33
r198 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.24 $Y=3.33
+ $X2=8.155 $Y2=3.33
r199 46 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.215 $Y=3.245
+ $X2=11.215 $Y2=3.33
r200 46 48 37.8909 $w=3.28e-07 $l=1.085e-06 $layer=LI1_cond $X=11.215 $Y=3.245
+ $X2=11.215 $Y2=2.16
r201 42 112 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.735 $Y=3.245
+ $X2=9.735 $Y2=3.33
r202 42 44 14.1586 $w=3.48e-07 $l=4.3e-07 $layer=LI1_cond $X=9.735 $Y=3.245
+ $X2=9.735 $Y2=2.815
r203 38 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.155 $Y=3.245
+ $X2=8.155 $Y2=3.33
r204 38 40 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.155 $Y=3.245
+ $X2=8.155 $Y2=2.815
r205 34 109 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=5.88 $Y=3.245
+ $X2=5.88 $Y2=3.33
r206 34 36 20.8457 $w=3.38e-07 $l=6.15e-07 $layer=LI1_cond $X=5.88 $Y=3.245
+ $X2=5.88 $Y2=2.63
r207 30 106 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=4.242 $Y=3.245
+ $X2=4.242 $Y2=3.33
r208 30 32 19.1101 $w=3.93e-07 $l=6.55e-07 $layer=LI1_cond $X=4.242 $Y=3.245
+ $X2=4.242 $Y2=2.59
r209 26 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=3.245
+ $X2=1.74 $Y2=3.33
r210 26 28 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=1.74 $Y=3.245
+ $X2=1.74 $Y2=2.695
r211 22 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r212 22 24 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.755
r213 7 48 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=11.08
+ $Y=2.015 $X2=11.215 $Y2=2.16
r214 6 44 600 $w=1.7e-07 $l=3.49821e-07 $layer=licon1_PDIFF $count=1 $X=9.565
+ $Y=2.54 $X2=9.735 $Y2=2.815
r215 5 40 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=8.02
+ $Y=2.54 $X2=8.155 $Y2=2.815
r216 4 36 600 $w=1.7e-07 $l=4.82442e-07 $layer=licon1_PDIFF $count=1 $X=5.49
+ $Y=2.315 $X2=5.84 $Y2=2.63
r217 3 32 600 $w=1.7e-07 $l=3.47851e-07 $layer=licon1_PDIFF $count=1 $X=4.075
+ $Y=2.315 $X2=4.24 $Y2=2.59
r218 2 28 600 $w=1.7e-07 $l=9.70155e-07 $layer=licon1_PDIFF $count=1 $X=1.605
+ $Y=1.79 $X2=1.74 $Y2=2.695
r219 1 24 600 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=2.54 $X2=0.73 $Y2=2.755
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_1%Q_N 1 2 9 11 12 13 14 15 22 39
r29 22 39 1.62667 $w=3.15e-07 $l=8.54576e-08 $layer=LI1_cond $X=10.277 $Y=1.337
+ $X2=10.21 $Y2=1.295
r30 15 35 1.46342 $w=3.13e-07 $l=4e-08 $layer=LI1_cond $X=10.277 $Y=2.775
+ $X2=10.277 $Y2=2.815
r31 14 15 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=10.277 $Y=2.405
+ $X2=10.277 $Y2=2.775
r32 13 14 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=10.277 $Y=2.035
+ $X2=10.277 $Y2=2.405
r33 13 27 1.82927 $w=3.13e-07 $l=5e-08 $layer=LI1_cond $X=10.277 $Y=2.035
+ $X2=10.277 $Y2=1.985
r34 12 27 11.7074 $w=3.13e-07 $l=3.2e-07 $layer=LI1_cond $X=10.277 $Y=1.665
+ $X2=10.277 $Y2=1.985
r35 11 39 0.88 $w=3.05e-07 $l=2.2e-08 $layer=LI1_cond $X=10.21 $Y=1.273
+ $X2=10.21 $Y2=1.295
r36 11 12 11.2317 $w=3.13e-07 $l=3.07e-07 $layer=LI1_cond $X=10.277 $Y=1.358
+ $X2=10.277 $Y2=1.665
r37 11 22 0.768295 $w=3.13e-07 $l=2.1e-08 $layer=LI1_cond $X=10.277 $Y=1.358
+ $X2=10.277 $Y2=1.337
r38 7 11 11.4767 $w=3.3e-07 $l=3.36666e-07 $layer=LI1_cond $X=10.15 $Y=0.965
+ $X2=10.21 $Y2=1.273
r39 7 9 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=10.15 $Y=0.965
+ $X2=10.15 $Y2=0.515
r40 2 35 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.07
+ $Y=1.84 $X2=10.205 $Y2=2.815
r41 2 27 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.07
+ $Y=1.84 $X2=10.205 $Y2=1.985
r42 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.01
+ $Y=0.37 $X2=10.15 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_1%Q 1 2 9 13 14 15 16 24 33
r19 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=11.72 $Y=2.405
+ $X2=11.72 $Y2=2.775
r20 14 24 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=11.72 $Y=1.967
+ $X2=11.72 $Y2=1.985
r21 14 33 7.83357 $w=3.28e-07 $l=1.47e-07 $layer=LI1_cond $X=11.72 $Y=1.967
+ $X2=11.72 $Y2=1.82
r22 14 15 12.3276 $w=3.28e-07 $l=3.53e-07 $layer=LI1_cond $X=11.72 $Y=2.052
+ $X2=11.72 $Y2=2.405
r23 14 24 2.33981 $w=3.28e-07 $l=6.7e-08 $layer=LI1_cond $X=11.72 $Y=2.052
+ $X2=11.72 $Y2=1.985
r24 13 33 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=11.8 $Y=1.05
+ $X2=11.8 $Y2=1.82
r25 7 13 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=11.72 $Y=0.885
+ $X2=11.72 $Y2=1.05
r26 7 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=11.72 $Y=0.885
+ $X2=11.72 $Y2=0.515
r27 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=11.585
+ $Y=1.84 $X2=11.72 $Y2=2.815
r28 2 24 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=11.585
+ $Y=1.84 $X2=11.72 $Y2=1.985
r29 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.58
+ $Y=0.37 $X2=11.72 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFSBP_1%VGND 1 2 3 4 5 6 7 24 26 30 34 38 42 46 49
+ 50 52 53 54 56 68 75 87 96 97 100 103 106 110 116
c130 38 0 2.3488e-20 $X=6.02 $Y=0.495
c131 30 0 1.39813e-19 $X=1.7 $Y=0.505
r132 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r133 110 113 9.62063 $w=6.88e-07 $l=5.55e-07 $layer=LI1_cond $X=8.41 $Y=0
+ $X2=8.41 $Y2=0.555
r134 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r135 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r136 101 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=1.68 $Y2=0
r137 100 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r138 97 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r139 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r140 94 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.385 $Y=0
+ $X2=11.22 $Y2=0
r141 94 96 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.385 $Y=0
+ $X2=11.76 $Y2=0
r142 93 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r143 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r144 90 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=10.8
+ $Y2=0
r145 89 92 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=9.84 $Y=0 $X2=10.8
+ $Y2=0
r146 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r147 87 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.055 $Y=0
+ $X2=11.22 $Y2=0
r148 87 92 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.055 $Y=0
+ $X2=10.8 $Y2=0
r149 86 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=9.84
+ $Y2=0
r150 86 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=8.4
+ $Y2=0
r151 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r152 83 110 9.22683 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=8.755 $Y=0
+ $X2=8.41 $Y2=0
r153 83 85 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=8.755 $Y=0
+ $X2=9.36 $Y2=0
r154 82 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r155 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r156 79 82 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=7.92 $Y2=0
r157 78 81 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.48 $Y=0 $X2=7.92
+ $Y2=0
r158 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r159 76 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.185 $Y=0
+ $X2=6.02 $Y2=0
r160 76 78 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.185 $Y=0 $X2=6.48
+ $Y2=0
r161 75 110 9.22683 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=8.065 $Y=0
+ $X2=8.41 $Y2=0
r162 75 81 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=8.065 $Y=0
+ $X2=7.92 $Y2=0
r163 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r164 71 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r165 70 73 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r166 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r167 68 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.855 $Y=0
+ $X2=6.02 $Y2=0
r168 68 73 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.855 $Y=0
+ $X2=5.52 $Y2=0
r169 67 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r170 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r171 64 67 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=4.08 $Y2=0
r172 64 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r173 63 66 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r174 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r175 61 103 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.865 $Y=0
+ $X2=1.735 $Y2=0
r176 61 63 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.16
+ $Y2=0
r177 59 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r178 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r179 56 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.67 $Y2=0
r180 56 58 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r181 54 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r182 54 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r183 54 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r184 52 85 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=9.485 $Y=0
+ $X2=9.36 $Y2=0
r185 52 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.485 $Y=0 $X2=9.65
+ $Y2=0
r186 51 89 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=9.815 $Y=0 $X2=9.84
+ $Y2=0
r187 51 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.815 $Y=0 $X2=9.65
+ $Y2=0
r188 49 66 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.105 $Y=0 $X2=4.08
+ $Y2=0
r189 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.105 $Y=0 $X2=4.27
+ $Y2=0
r190 48 70 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.435 $Y=0
+ $X2=4.56 $Y2=0
r191 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.435 $Y=0 $X2=4.27
+ $Y2=0
r192 44 116 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.22 $Y=0.085
+ $X2=11.22 $Y2=0
r193 44 46 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=11.22 $Y=0.085
+ $X2=11.22 $Y2=0.495
r194 40 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.65 $Y=0.085
+ $X2=9.65 $Y2=0
r195 40 42 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=9.65 $Y=0.085
+ $X2=9.65 $Y2=0.55
r196 36 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.02 $Y=0.085
+ $X2=6.02 $Y2=0
r197 36 38 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.02 $Y=0.085
+ $X2=6.02 $Y2=0.495
r198 32 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.27 $Y=0.085
+ $X2=4.27 $Y2=0
r199 32 34 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.27 $Y=0.085
+ $X2=4.27 $Y2=0.55
r200 28 103 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.735 $Y=0.085
+ $X2=1.735 $Y2=0
r201 28 30 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=1.735 $Y=0.085
+ $X2=1.735 $Y2=0.505
r202 27 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=0
+ $X2=0.67 $Y2=0
r203 26 103 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.605 $Y=0
+ $X2=1.735 $Y2=0
r204 26 27 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=1.605 $Y=0
+ $X2=0.795 $Y2=0
r205 22 100 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0
r206 22 24 24.2013 $w=2.48e-07 $l=5.25e-07 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0.61
r207 7 46 91 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=2 $X=11 $Y=0.37
+ $X2=11.22 $Y2=0.495
r208 6 42 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=9.505
+ $Y=0.37 $X2=9.65 $Y2=0.55
r209 5 113 91 $w=1.7e-07 $l=5.85235e-07 $layer=licon1_NDIFF $count=2 $X=8.09
+ $Y=0.37 $X2=8.59 $Y2=0.555
r210 4 38 91 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=2 $X=5.695
+ $Y=0.37 $X2=6.02 $Y2=0.495
r211 3 34 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.13
+ $Y=0.405 $X2=4.27 $Y2=0.55
r212 2 30 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=1.56
+ $Y=0.37 $X2=1.7 $Y2=0.505
r213 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.4 $X2=0.71 $Y2=0.61
.ends


* File: sky130_fd_sc_ms__o21a_4.spice
* Created: Fri Aug 28 17:54:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o21a_4.pex.spice"
.subckt sky130_fd_sc_ms__o21a_4  VNB VPB A2 A1 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_A1_M1015_g N_A_27_125#_M1015_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1136 AS=0.1824 PD=0.995 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.7 A=0.096 P=1.58 MULT=1
MM1003 N_A_27_125#_M1003_d N_A2_M1003_g N_VGND_M1015_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1136 PD=0.92 PS=0.995 NRD=0 NRS=0.936 M=1 R=4.26667 SA=75000.7
+ SB=75002.2 A=0.096 P=1.58 MULT=1
MM1004 N_A_27_125#_M1003_d N_A2_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1376 PD=0.92 PS=1.07 NRD=0 NRS=14.988 M=1 R=4.26667 SA=75001.1
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1018 N_VGND_M1004_s N_A1_M1018_g N_A_27_125#_M1018_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1376 AS=0.0896 PD=1.07 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75001.7
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1010 N_A_27_125#_M1018_s N_B1_M1010_g N_A_219_387#_M1010_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1019 N_A_27_125#_M1019_d N_B1_M1019_g N_A_219_387#_M1010_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.2336 AS=0.0896 PD=2.01 PS=0.92 NRD=14.988 NRS=0 M=1 R=4.26667
+ SA=75002.6 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1001 N_VGND_M1001_d N_A_219_387#_M1001_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_A_219_387#_M1002_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.11655 AS=0.1036 PD=1.055 PS=1.02 NRD=2.424 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1002_d N_A_219_387#_M1005_g N_X_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.11655 AS=0.1036 PD=1.055 PS=1.02 NRD=3.24 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_A_219_387#_M1006_g N_X_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1014 N_VPWR_M1014_d N_A1_M1014_g N_A_119_387#_M1014_s VPB PSHORT L=0.18 W=1
+ AD=0.28 AS=0.16 PD=2.56 PS=1.32 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90000.2
+ SB=90004.4 A=0.18 P=2.36 MULT=1
MM1011 N_A_219_387#_M1011_d N_A2_M1011_g N_A_119_387#_M1014_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.16 PD=1.27 PS=1.32 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.7
+ SB=90003.9 A=0.18 P=2.36 MULT=1
MM1013 N_A_219_387#_M1011_d N_A2_M1013_g N_A_119_387#_M1013_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.16 PD=1.27 PS=1.32 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90001.1
+ SB=90003.5 A=0.18 P=2.36 MULT=1
MM1016 N_VPWR_M1016_d N_A1_M1016_g N_A_119_387#_M1013_s VPB PSHORT L=0.18 W=1
+ AD=0.186087 AS=0.16 PD=1.47826 PS=1.32 NRD=8.8453 NRS=0 M=1 R=5.55556
+ SA=90001.6 SB=90003 A=0.18 P=2.36 MULT=1
MM1000 N_A_219_387#_M1000_d N_B1_M1000_g N_VPWR_M1016_d VPB PSHORT L=0.18 W=0.84
+ AD=0.147 AS=0.156313 PD=1.19 PS=1.24174 NRD=1.1623 NRS=8.1952 M=1 R=4.66667
+ SA=90002.2 SB=90002.9 A=0.1512 P=2.04 MULT=1
MM1008 N_A_219_387#_M1000_d N_B1_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=0.84
+ AD=0.147 AS=0.228 PD=1.19 PS=1.43143 NRD=15.2281 NRS=24.625 M=1 R=4.66667
+ SA=90002.7 SB=90002.4 A=0.1512 P=2.04 MULT=1
MM1007 N_X_M1007_d N_A_219_387#_M1007_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.304 PD=1.39 PS=1.90857 NRD=0 NRS=29.0181 M=1 R=6.22222
+ SA=90002.6 SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1009 N_X_M1007_d N_A_219_387#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003.1
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1012 N_X_M1012_d N_A_219_387#_M1012_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003.6
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1017 N_X_M1012_d N_A_219_387#_M1017_g N_VPWR_M1017_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90004.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4204 P=16
*
.include "sky130_fd_sc_ms__o21a_4.pxi.spice"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfxtp_1 CLK D VGND VNB VPB VPWR Q
X0 a_457_503# a_209_368# a_564_463# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X1 VPWR a_564_463# a_713_458# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X2 VGND a_1210_314# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VPWR a_27_74# a_209_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X4 a_1210_314# a_1014_424# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X5 a_564_463# a_209_368# a_731_101# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X6 VGND D a_457_503# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X7 a_1014_424# a_27_74# a_1168_124# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X8 VPWR D a_457_503# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X9 a_1168_124# a_1210_314# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X10 a_27_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X11 a_1121_508# a_1210_314# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X12 VGND a_27_74# a_209_368# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_1210_314# a_1014_424# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X14 VPWR a_1210_314# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 a_564_463# a_27_74# a_671_503# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X16 VGND a_564_463# a_713_458# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X17 a_713_458# a_27_74# a_1014_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X18 a_731_101# a_713_458# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X19 a_713_458# a_209_368# a_1014_424# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X20 a_457_503# a_27_74# a_564_463# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X21 a_1014_424# a_209_368# a_1121_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X22 a_27_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 a_671_503# a_713_458# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
.ends

* File: sky130_fd_sc_ms__dfbbp_1.pxi.spice
* Created: Fri Aug 28 17:21:49 2020
* 
x_PM_SKY130_FD_SC_MS__DFBBP_1%CLK N_CLK_M1029_g N_CLK_M1018_g CLK N_CLK_c_266_n
+ N_CLK_c_267_n PM_SKY130_FD_SC_MS__DFBBP_1%CLK
x_PM_SKY130_FD_SC_MS__DFBBP_1%D N_D_M1032_g N_D_M1013_g D N_D_c_305_n
+ PM_SKY130_FD_SC_MS__DFBBP_1%D
x_PM_SKY130_FD_SC_MS__DFBBP_1%A_671_93# N_A_671_93#_M1022_d N_A_671_93#_M1020_d
+ N_A_671_93#_c_336_n N_A_671_93#_M1036_g N_A_671_93#_M1009_g
+ N_A_671_93#_M1003_g N_A_671_93#_c_339_n N_A_671_93#_c_340_n
+ N_A_671_93#_M1006_g N_A_671_93#_c_341_n N_A_671_93#_c_342_n
+ N_A_671_93#_c_356_p N_A_671_93#_c_379_p N_A_671_93#_c_350_n
+ N_A_671_93#_c_351_n N_A_671_93#_c_352_n N_A_671_93#_c_343_n
+ N_A_671_93#_c_344_n N_A_671_93#_c_406_p N_A_671_93#_c_345_n
+ N_A_671_93#_c_346_n N_A_671_93#_c_347_n PM_SKY130_FD_SC_MS__DFBBP_1%A_671_93#
x_PM_SKY130_FD_SC_MS__DFBBP_1%SET_B N_SET_B_M1033_g N_SET_B_M1020_g
+ N_SET_B_M1034_g N_SET_B_M1023_g N_SET_B_c_500_n N_SET_B_c_501_n
+ N_SET_B_c_502_n N_SET_B_c_503_n N_SET_B_c_526_n N_SET_B_c_530_n
+ N_SET_B_c_504_n N_SET_B_c_505_n N_SET_B_c_506_n N_SET_B_c_507_n
+ N_SET_B_c_508_n N_SET_B_c_509_n N_SET_B_c_494_n SET_B N_SET_B_c_496_n
+ N_SET_B_c_497_n PM_SKY130_FD_SC_MS__DFBBP_1%SET_B
x_PM_SKY130_FD_SC_MS__DFBBP_1%A_520_87# N_A_520_87#_M1004_d N_A_520_87#_M1016_d
+ N_A_520_87#_M1022_g N_A_520_87#_M1035_g N_A_520_87#_c_656_n
+ N_A_520_87#_c_657_n N_A_520_87#_c_666_n N_A_520_87#_c_658_n
+ N_A_520_87#_c_659_n N_A_520_87#_c_660_n N_A_520_87#_c_661_n
+ N_A_520_87#_c_662_n N_A_520_87#_c_663_n N_A_520_87#_c_664_n
+ PM_SKY130_FD_SC_MS__DFBBP_1%A_520_87#
x_PM_SKY130_FD_SC_MS__DFBBP_1%A_1062_93# N_A_1062_93#_M1007_s
+ N_A_1062_93#_M1000_s N_A_1062_93#_M1030_g N_A_1062_93#_M1011_g
+ N_A_1062_93#_M1024_g N_A_1062_93#_c_759_n N_A_1062_93#_M1031_g
+ N_A_1062_93#_c_760_n N_A_1062_93#_c_761_n N_A_1062_93#_c_762_n
+ N_A_1062_93#_c_776_n N_A_1062_93#_c_777_n N_A_1062_93#_c_763_n
+ N_A_1062_93#_c_764_n N_A_1062_93#_c_765_n N_A_1062_93#_c_766_n
+ N_A_1062_93#_c_767_n N_A_1062_93#_c_768_n N_A_1062_93#_c_769_n
+ N_A_1062_93#_c_770_n N_A_1062_93#_c_771_n N_A_1062_93#_c_772_n
+ PM_SKY130_FD_SC_MS__DFBBP_1%A_1062_93#
x_PM_SKY130_FD_SC_MS__DFBBP_1%A_27_74# N_A_27_74#_M1029_s N_A_27_74#_M1018_s
+ N_A_27_74#_M1017_g N_A_27_74#_M1028_g N_A_27_74#_c_904_n N_A_27_74#_c_905_n
+ N_A_27_74#_c_906_n N_A_27_74#_c_907_n N_A_27_74#_c_908_n N_A_27_74#_c_926_n
+ N_A_27_74#_c_927_n N_A_27_74#_M1004_g N_A_27_74#_M1039_g N_A_27_74#_c_929_n
+ N_A_27_74#_M1005_g N_A_27_74#_M1014_g N_A_27_74#_c_910_n N_A_27_74#_c_931_n
+ N_A_27_74#_c_911_n N_A_27_74#_c_912_n N_A_27_74#_c_933_n N_A_27_74#_c_934_n
+ N_A_27_74#_c_913_n N_A_27_74#_c_914_n N_A_27_74#_c_915_n N_A_27_74#_c_916_n
+ N_A_27_74#_c_917_n N_A_27_74#_c_918_n N_A_27_74#_c_936_n N_A_27_74#_c_919_n
+ N_A_27_74#_c_920_n N_A_27_74#_c_921_n N_A_27_74#_c_922_n N_A_27_74#_c_923_n
+ PM_SKY130_FD_SC_MS__DFBBP_1%A_27_74#
x_PM_SKY130_FD_SC_MS__DFBBP_1%A_214_74# N_A_214_74#_M1017_d N_A_214_74#_M1028_d
+ N_A_214_74#_c_1121_n N_A_214_74#_M1025_g N_A_214_74#_M1016_g
+ N_A_214_74#_c_1124_n N_A_214_74#_c_1125_n N_A_214_74#_M1012_g
+ N_A_214_74#_M1001_g N_A_214_74#_c_1127_n N_A_214_74#_c_1128_n
+ N_A_214_74#_c_1129_n N_A_214_74#_c_1138_n N_A_214_74#_c_1130_n
+ N_A_214_74#_c_1131_n N_A_214_74#_c_1132_n N_A_214_74#_c_1133_n
+ N_A_214_74#_c_1134_n PM_SKY130_FD_SC_MS__DFBBP_1%A_214_74#
x_PM_SKY130_FD_SC_MS__DFBBP_1%A_1474_446# N_A_1474_446#_M1027_d
+ N_A_1474_446#_M1023_d N_A_1474_446#_M1015_g N_A_1474_446#_c_1271_n
+ N_A_1474_446#_M1021_g N_A_1474_446#_M1008_g N_A_1474_446#_M1002_g
+ N_A_1474_446#_c_1261_n N_A_1474_446#_c_1262_n N_A_1474_446#_c_1263_n
+ N_A_1474_446#_c_1275_n N_A_1474_446#_M1026_g N_A_1474_446#_c_1264_n
+ N_A_1474_446#_M1019_g N_A_1474_446#_c_1276_n N_A_1474_446#_c_1265_n
+ N_A_1474_446#_c_1266_n N_A_1474_446#_c_1277_n N_A_1474_446#_c_1278_n
+ N_A_1474_446#_c_1267_n N_A_1474_446#_c_1280_n N_A_1474_446#_c_1281_n
+ N_A_1474_446#_c_1282_n N_A_1474_446#_c_1302_n N_A_1474_446#_c_1324_n
+ N_A_1474_446#_c_1268_n N_A_1474_446#_c_1269_n
+ PM_SKY130_FD_SC_MS__DFBBP_1%A_1474_446#
x_PM_SKY130_FD_SC_MS__DFBBP_1%A_1314_424# N_A_1314_424#_M1012_d
+ N_A_1314_424#_M1005_d N_A_1314_424#_M1027_g N_A_1314_424#_M1010_g
+ N_A_1314_424#_c_1448_n N_A_1314_424#_c_1439_n N_A_1314_424#_c_1440_n
+ N_A_1314_424#_c_1441_n N_A_1314_424#_c_1442_n N_A_1314_424#_c_1450_n
+ N_A_1314_424#_c_1443_n N_A_1314_424#_c_1444_n N_A_1314_424#_c_1445_n
+ N_A_1314_424#_c_1446_n PM_SKY130_FD_SC_MS__DFBBP_1%A_1314_424#
x_PM_SKY130_FD_SC_MS__DFBBP_1%RESET_B N_RESET_B_M1007_g N_RESET_B_M1000_g
+ N_RESET_B_c_1544_n N_RESET_B_c_1545_n RESET_B N_RESET_B_c_1546_n
+ N_RESET_B_c_1547_n PM_SKY130_FD_SC_MS__DFBBP_1%RESET_B
x_PM_SKY130_FD_SC_MS__DFBBP_1%A_2320_410# N_A_2320_410#_M1019_s
+ N_A_2320_410#_M1026_s N_A_2320_410#_M1037_g N_A_2320_410#_M1038_g
+ N_A_2320_410#_c_1590_n N_A_2320_410#_c_1591_n N_A_2320_410#_c_1592_n
+ N_A_2320_410#_c_1597_n N_A_2320_410#_c_1598_n N_A_2320_410#_c_1593_n
+ N_A_2320_410#_c_1594_n N_A_2320_410#_c_1595_n
+ PM_SKY130_FD_SC_MS__DFBBP_1%A_2320_410#
x_PM_SKY130_FD_SC_MS__DFBBP_1%VPWR N_VPWR_M1018_d N_VPWR_M1013_s N_VPWR_M1009_d
+ N_VPWR_M1011_d N_VPWR_M1015_d N_VPWR_M1024_d N_VPWR_M1000_d N_VPWR_M1026_d
+ N_VPWR_c_1650_n N_VPWR_c_1651_n N_VPWR_c_1652_n N_VPWR_c_1653_n
+ N_VPWR_c_1654_n N_VPWR_c_1655_n N_VPWR_c_1656_n N_VPWR_c_1657_n
+ N_VPWR_c_1658_n VPWR N_VPWR_c_1659_n N_VPWR_c_1660_n N_VPWR_c_1661_n
+ N_VPWR_c_1662_n N_VPWR_c_1663_n N_VPWR_c_1664_n N_VPWR_c_1649_n
+ N_VPWR_c_1666_n N_VPWR_c_1667_n N_VPWR_c_1668_n N_VPWR_c_1669_n
+ N_VPWR_c_1670_n N_VPWR_c_1671_n N_VPWR_c_1672_n N_VPWR_c_1673_n
+ PM_SKY130_FD_SC_MS__DFBBP_1%VPWR
x_PM_SKY130_FD_SC_MS__DFBBP_1%A_422_125# N_A_422_125#_M1032_d
+ N_A_422_125#_M1013_d N_A_422_125#_c_1795_n N_A_422_125#_c_1796_n
+ N_A_422_125#_c_1797_n N_A_422_125#_c_1799_n N_A_422_125#_c_1798_n
+ PM_SKY130_FD_SC_MS__DFBBP_1%A_422_125#
x_PM_SKY130_FD_SC_MS__DFBBP_1%Q_N N_Q_N_M1002_d N_Q_N_M1008_d N_Q_N_c_1851_n
+ N_Q_N_c_1852_n Q_N Q_N Q_N Q_N N_Q_N_c_1853_n PM_SKY130_FD_SC_MS__DFBBP_1%Q_N
x_PM_SKY130_FD_SC_MS__DFBBP_1%Q N_Q_M1038_d N_Q_M1037_d Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_MS__DFBBP_1%Q
x_PM_SKY130_FD_SC_MS__DFBBP_1%VGND N_VGND_M1029_d N_VGND_M1032_s N_VGND_M1036_d
+ N_VGND_M1006_s N_VGND_M1021_d N_VGND_M1007_d N_VGND_M1019_d N_VGND_c_1902_n
+ N_VGND_c_1903_n N_VGND_c_1904_n N_VGND_c_1905_n N_VGND_c_1935_n
+ N_VGND_c_1906_n N_VGND_c_1907_n N_VGND_c_1908_n N_VGND_c_1909_n
+ N_VGND_c_1910_n N_VGND_c_1911_n N_VGND_c_1912_n N_VGND_c_1913_n VGND
+ N_VGND_c_1914_n N_VGND_c_1915_n N_VGND_c_1916_n N_VGND_c_1917_n
+ N_VGND_c_1918_n N_VGND_c_1919_n N_VGND_c_1920_n N_VGND_c_1921_n
+ N_VGND_c_1922_n N_VGND_c_1923_n PM_SKY130_FD_SC_MS__DFBBP_1%VGND
x_PM_SKY130_FD_SC_MS__DFBBP_1%A_872_119# N_A_872_119#_M1033_d
+ N_A_872_119#_M1030_d N_A_872_119#_c_2063_n N_A_872_119#_c_2064_n
+ N_A_872_119#_c_2065_n PM_SKY130_FD_SC_MS__DFBBP_1%A_872_119#
x_PM_SKY130_FD_SC_MS__DFBBP_1%A_1708_74# N_A_1708_74#_M1034_d
+ N_A_1708_74#_M1031_d N_A_1708_74#_c_2096_n N_A_1708_74#_c_2093_n
+ N_A_1708_74#_c_2094_n N_A_1708_74#_c_2100_n
+ PM_SKY130_FD_SC_MS__DFBBP_1%A_1708_74#
cc_1 VNB N_CLK_M1018_g 0.00667765f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.4
cc_2 VNB CLK 0.00713458f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_CLK_c_266_n 0.0313968f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.385
cc_4 VNB N_CLK_c_267_n 0.021865f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.22
cc_5 VNB N_D_M1032_g 0.0416847f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_6 VNB N_A_671_93#_c_336_n 0.0177094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_671_93#_M1009_g 0.0120618f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.385
cc_8 VNB N_A_671_93#_M1003_g 0.00480377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_671_93#_c_339_n 0.0275397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_671_93#_c_340_n 0.0138218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_671_93#_c_341_n 0.00318059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_671_93#_c_342_n 0.0535566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_671_93#_c_343_n 0.00450078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_671_93#_c_344_n 9.76271e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_671_93#_c_345_n 0.00235757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_671_93#_c_346_n 0.00434991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_671_93#_c_347_n 0.0395513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_SET_B_M1033_g 0.0246772f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_19 VNB N_SET_B_M1034_g 0.0295617f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.385
cc_20 VNB N_SET_B_c_494_n 0.00194515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB SET_B 0.00463034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_SET_B_c_496_n 0.025082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_SET_B_c_497_n 0.0162335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_520_87#_M1035_g 0.00432871f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.385
cc_25 VNB N_A_520_87#_c_656_n 0.00623074f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.55
cc_26 VNB N_A_520_87#_c_657_n 0.0111246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_520_87#_c_658_n 0.00274783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_520_87#_c_659_n 0.0032561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_520_87#_c_660_n 0.0198117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_520_87#_c_661_n 0.00185643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_520_87#_c_662_n 0.00362121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_520_87#_c_663_n 0.0285461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_520_87#_c_664_n 0.0165111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_1062_93#_M1011_g 0.00427276f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.385
cc_35 VNB N_A_1062_93#_M1024_g 0.013722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_1062_93#_c_759_n 0.0188807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_1062_93#_c_760_n 0.0191354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_1062_93#_c_761_n 0.00591265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_1062_93#_c_762_n 0.00268812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_1062_93#_c_763_n 0.0181401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_1062_93#_c_764_n 0.0339695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1062_93#_c_765_n 0.00239212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1062_93#_c_766_n 0.00248349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1062_93#_c_767_n 0.00786335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1062_93#_c_768_n 0.00351751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_1062_93#_c_769_n 0.0309621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1062_93#_c_770_n 0.0162912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1062_93#_c_771_n 0.0360877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1062_93#_c_772_n 0.00811013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_27_74#_M1017_g 0.0224989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_27_74#_M1028_g 0.0016208f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.22
cc_52 VNB N_A_27_74#_c_904_n 0.00816286f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.365
cc_53 VNB N_A_27_74#_c_905_n 0.0569175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_27_74#_c_906_n 0.0683039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_27_74#_c_907_n 0.0123817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_27_74#_c_908_n 0.00940304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_27_74#_M1004_g 0.0197931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_27_74#_c_910_n 0.0122917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_27_74#_c_911_n 0.021853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_27_74#_c_912_n 0.0299666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_27_74#_c_913_n 3.17047e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_27_74#_c_914_n 0.00769092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_27_74#_c_915_n 0.00166555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_27_74#_c_916_n 0.00203856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_27_74#_c_917_n 0.0390929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_27_74#_c_918_n 0.00710642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_27_74#_c_919_n 6.96084e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_27_74#_c_920_n 0.0117531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_27_74#_c_921_n 0.0107725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_27_74#_c_922_n 0.0304326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_27_74#_c_923_n 0.0177878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_214_74#_c_1121_n 0.0183009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_214_74#_M1025_g 0.0355213f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.385
cc_74 VNB N_A_214_74#_M1016_g 0.0143717f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.365
cc_75 VNB N_A_214_74#_c_1124_n 0.286458f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.365
cc_76 VNB N_A_214_74#_c_1125_n 0.00962308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_214_74#_M1012_g 0.0235622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_214_74#_c_1127_n 0.00690488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_214_74#_c_1128_n 0.0250872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_214_74#_c_1129_n 0.0218065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_214_74#_c_1130_n 0.00299917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_214_74#_c_1131_n 0.00526652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_214_74#_c_1132_n 0.00123797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_214_74#_c_1133_n 0.0192504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_214_74#_c_1134_n 0.0339982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1474_446#_M1021_g 0.065314f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.365
cc_87 VNB N_A_1474_446#_M1008_g 5.47829e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1474_446#_M1002_g 0.0290725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1474_446#_c_1261_n 0.0432697f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1474_446#_c_1262_n 0.0167158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1474_446#_c_1263_n 5.77437e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1474_446#_c_1264_n 0.0186482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1474_446#_c_1265_n 0.0305356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1474_446#_c_1266_n 0.00972803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1474_446#_c_1267_n 0.00337358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1474_446#_c_1268_n 0.00229347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1474_446#_c_1269_n 0.0223175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1314_424#_M1010_g 0.00626735f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=1.385
cc_99 VNB N_A_1314_424#_c_1439_n 0.0044036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1314_424#_c_1440_n 6.58668e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1314_424#_c_1441_n 0.0156357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1314_424#_c_1442_n 0.0146937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1314_424#_c_1443_n 0.00342912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1314_424#_c_1444_n 0.00465144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1314_424#_c_1445_n 0.0314409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1314_424#_c_1446_n 0.0162593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_RESET_B_M1007_g 0.0265205f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_108 VNB N_RESET_B_M1000_g 5.85784e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_RESET_B_c_1544_n 0.0211328f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.385
cc_110 VNB N_RESET_B_c_1545_n 0.0150632f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.385
cc_111 VNB N_RESET_B_c_1546_n 0.0194514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_RESET_B_c_1547_n 0.0111244f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.365
cc_113 VNB N_A_2320_410#_M1037_g 0.00566674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_2320_410#_M1038_g 0.0260646f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.22
cc_115 VNB N_A_2320_410#_c_1590_n 0.0380679f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=1.365
cc_116 VNB N_A_2320_410#_c_1591_n 0.0173865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_2320_410#_c_1592_n 0.0097541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_2320_410#_c_1593_n 0.00322651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_2320_410#_c_1594_n 4.84981e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_2320_410#_c_1595_n 0.00100541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VPWR_c_1649_n 0.541827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_422_125#_c_1795_n 7.66685e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_A_422_125#_c_1796_n 0.00845715f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=1.385
cc_124 VNB N_A_422_125#_c_1797_n 0.00204574f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=1.385
cc_125 VNB N_A_422_125#_c_1798_n 0.00468724f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=1.365
cc_126 VNB N_Q_N_c_1851_n 0.00922224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_Q_N_c_1852_n 0.00591911f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.22
cc_128 VNB N_Q_N_c_1853_n 0.00272629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB Q 0.0550644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1902_n 0.00641543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1903_n 0.0185285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1904_n 0.0142221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1905_n 0.00445932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1906_n 0.00796047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1907_n 0.0144974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1908_n 0.00638918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1909_n 0.0441488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1910_n 0.00492725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_1911_n 0.00285168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_1912_n 0.0318016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_1913_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_1914_n 0.0189171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_1915_n 0.0594655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_1916_n 0.0411788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_1917_n 0.0533685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_1918_n 0.0203853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_1919_n 0.655422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_1920_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_1921_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_1922_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_1923_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_A_872_119#_c_2063_n 0.0140742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_A_872_119#_c_2064_n 0.00771386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_A_872_119#_c_2065_n 0.00899945f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=1.55
cc_155 VNB N_A_1708_74#_c_2093_n 0.00591279f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=1.385
cc_156 VNB N_A_1708_74#_c_2094_n 0.00338117f $X=-0.19 $Y=-0.245 $X2=0.52
+ $Y2=1.385
cc_157 VPB N_CLK_M1018_g 0.0302268f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=2.4
cc_158 VPB N_D_M1032_g 0.0104669f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_159 VPB N_D_M1013_g 0.0225044f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB D 0.00549977f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_D_c_305_n 0.056611f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.22
cc_162 VPB N_A_671_93#_M1009_g 0.026313f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.385
cc_163 VPB N_A_671_93#_M1003_g 0.0243756f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_A_671_93#_c_350_n 9.60827e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_A_671_93#_c_351_n 0.0113529f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_A_671_93#_c_352_n 0.00255343f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_SET_B_M1020_g 0.0227667f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_SET_B_M1023_g 0.0243689f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.365
cc_169 VPB N_SET_B_c_500_n 0.00408097f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_SET_B_c_501_n 0.0189453f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_SET_B_c_502_n 0.00177503f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_SET_B_c_503_n 0.00375549f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_SET_B_c_504_n 0.00166884f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_SET_B_c_505_n 0.00545982f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_SET_B_c_506_n 0.00246631f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_SET_B_c_507_n 0.00782661f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_SET_B_c_508_n 0.0113159f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_SET_B_c_509_n 0.00326001f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB SET_B 0.00379486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_SET_B_c_496_n 0.0115495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_SET_B_c_497_n 0.0127766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_520_87#_M1035_g 0.023585f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.385
cc_183 VPB N_A_520_87#_c_666_n 0.00705551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_520_87#_c_658_n 0.00912385f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_520_87#_c_662_n 0.00122969f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_1062_93#_M1011_g 0.02233f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.385
cc_187 VPB N_A_1062_93#_M1024_g 0.0304583f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_1062_93#_c_762_n 0.00426589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_1062_93#_c_776_n 0.0067531f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_1062_93#_c_777_n 0.0079042f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_27_74#_M1028_g 0.0240917f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.22
cc_192 VPB N_A_27_74#_c_908_n 0.083363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_27_74#_c_926_n 0.120382f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_27_74#_c_927_n 0.0123574f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_27_74#_M1039_g 0.0636487f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_27_74#_c_929_n 0.217425f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_27_74#_M1005_g 0.0187322f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_27_74#_c_931_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_27_74#_c_912_n 0.00278822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_27_74#_c_933_n 0.0514224f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_27_74#_c_934_n 0.00496437f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_27_74#_c_913_n 6.23525e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_27_74#_c_936_n 0.0135811f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_27_74#_c_919_n 0.00186525f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_27_74#_c_920_n 0.0279406f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_214_74#_M1016_g 0.0496632f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.365
cc_207 VPB N_A_214_74#_M1001_g 0.0247823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_208 VPB N_A_214_74#_c_1129_n 0.0313477f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_A_214_74#_c_1138_n 0.0114116f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_A_214_74#_c_1132_n 0.0164251f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_A_1474_446#_M1015_g 0.0258561f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_A_1474_446#_c_1271_n 0.01118f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.385
cc_213 VPB N_A_1474_446#_M1021_g 0.00586386f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.365
cc_214 VPB N_A_1474_446#_M1008_g 0.028708f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_A_1474_446#_c_1263_n 0.00855823f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_A_1474_446#_c_1275_n 0.0454609f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_1474_446#_c_1276_n 0.0136284f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_A_1474_446#_c_1277_n 0.0507018f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_1474_446#_c_1278_n 0.00203805f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_A_1474_446#_c_1267_n 0.00283937f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_1474_446#_c_1280_n 0.0158064f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_1474_446#_c_1281_n 0.00176398f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_A_1474_446#_c_1282_n 0.00479737f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_A_1314_424#_M1010_g 0.0307087f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.385
cc_225 VPB N_A_1314_424#_c_1448_n 0.00217643f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_1314_424#_c_1440_n 0.00368906f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_A_1314_424#_c_1450_n 0.00817579f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_RESET_B_M1000_g 0.0291849f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_2320_410#_M1037_g 0.0308782f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_A_2320_410#_c_1597_n 4.97507e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_A_2320_410#_c_1598_n 0.0022931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_2320_410#_c_1595_n 0.00298449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1650_n 0.00978155f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1651_n 0.0193804f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1652_n 0.0129015f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1653_n 0.00396484f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1654_n 0.0238731f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1655_n 0.0241773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1656_n 0.0152785f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1657_n 0.0310952f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1658_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1659_n 0.0214552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1660_n 0.0446599f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1661_n 0.0304123f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1662_n 0.0250757f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1663_n 0.0322037f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1664_n 0.0197489f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1649_n 0.131021f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1666_n 0.0273996f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1667_n 0.00803083f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1668_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1669_n 0.00490136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1670_n 0.0409001f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1671_n 0.0261359f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1672_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1673_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_A_422_125#_c_1799_n 0.00897263f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_A_422_125#_c_1798_n 0.00703237f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.365
cc_259 VPB Q_N 0.00508159f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.55
cc_260 VPB Q_N 0.0151096f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_Q_N_c_1853_n 0.00183998f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB Q 0.0542187f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 CLK N_A_27_74#_M1017_g 0.00134224f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_264 N_CLK_c_266_n N_A_27_74#_M1017_g 0.00404399f $X=0.52 $Y=1.385 $X2=0 $Y2=0
cc_265 N_CLK_c_267_n N_A_27_74#_M1017_g 0.0175656f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_266 N_CLK_M1018_g N_A_27_74#_M1028_g 0.0224977f $X=0.595 $Y=2.4 $X2=0 $Y2=0
cc_267 N_CLK_c_267_n N_A_27_74#_c_911_n 0.00593943f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_268 N_CLK_M1018_g N_A_27_74#_c_912_n 0.00383326f $X=0.595 $Y=2.4 $X2=0 $Y2=0
cc_269 CLK N_A_27_74#_c_912_n 0.0280545f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_270 N_CLK_c_266_n N_A_27_74#_c_912_n 0.00804857f $X=0.52 $Y=1.385 $X2=0 $Y2=0
cc_271 N_CLK_c_267_n N_A_27_74#_c_912_n 0.00404717f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_272 N_CLK_M1018_g N_A_27_74#_c_933_n 0.0159368f $X=0.595 $Y=2.4 $X2=0 $Y2=0
cc_273 N_CLK_M1018_g N_A_27_74#_c_934_n 0.0135649f $X=0.595 $Y=2.4 $X2=0 $Y2=0
cc_274 CLK N_A_27_74#_c_934_n 0.0203789f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_275 N_CLK_M1018_g N_A_27_74#_c_913_n 0.00169956f $X=0.595 $Y=2.4 $X2=0 $Y2=0
cc_276 CLK N_A_27_74#_c_913_n 0.0191154f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_277 N_CLK_c_266_n N_A_27_74#_c_913_n 6.75433e-19 $X=0.52 $Y=1.385 $X2=0 $Y2=0
cc_278 CLK N_A_27_74#_c_918_n 0.0015257f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_279 N_CLK_c_266_n N_A_27_74#_c_918_n 0.00144239f $X=0.52 $Y=1.385 $X2=0 $Y2=0
cc_280 N_CLK_c_267_n N_A_27_74#_c_918_n 0.00211436f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_281 N_CLK_M1018_g N_A_27_74#_c_936_n 0.00349541f $X=0.595 $Y=2.4 $X2=0 $Y2=0
cc_282 CLK N_A_27_74#_c_936_n 0.00921466f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_283 N_CLK_c_266_n N_A_27_74#_c_936_n 0.0053098f $X=0.52 $Y=1.385 $X2=0 $Y2=0
cc_284 CLK N_A_27_74#_c_922_n 0.00179043f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_285 N_CLK_c_266_n N_A_27_74#_c_922_n 0.0211768f $X=0.52 $Y=1.385 $X2=0 $Y2=0
cc_286 CLK N_A_214_74#_c_1131_n 0.00462759f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_287 N_CLK_M1018_g N_VPWR_c_1650_n 0.00348921f $X=0.595 $Y=2.4 $X2=0 $Y2=0
cc_288 N_CLK_M1018_g N_VPWR_c_1649_n 0.00986825f $X=0.595 $Y=2.4 $X2=0 $Y2=0
cc_289 N_CLK_M1018_g N_VPWR_c_1666_n 0.005209f $X=0.595 $Y=2.4 $X2=0 $Y2=0
cc_290 CLK N_VGND_c_1902_n 0.0160287f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_291 N_CLK_c_266_n N_VGND_c_1902_n 4.54296e-19 $X=0.52 $Y=1.385 $X2=0 $Y2=0
cc_292 N_CLK_c_267_n N_VGND_c_1902_n 0.00659657f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_293 N_CLK_c_267_n N_VGND_c_1914_n 0.00434272f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_294 N_CLK_c_267_n N_VGND_c_1919_n 0.00824429f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_295 N_D_M1032_g N_A_520_87#_c_656_n 4.05638e-19 $X=2.035 $Y=0.835 $X2=0 $Y2=0
cc_296 N_D_M1032_g N_A_27_74#_c_905_n 0.0170648f $X=2.035 $Y=0.835 $X2=0 $Y2=0
cc_297 N_D_M1032_g N_A_27_74#_c_906_n 0.00895007f $X=2.035 $Y=0.835 $X2=0 $Y2=0
cc_298 N_D_M1013_g N_A_27_74#_c_908_n 0.00819217f $X=2.52 $Y=2.525 $X2=0 $Y2=0
cc_299 D N_A_27_74#_c_908_n 0.00115219f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_300 N_D_c_305_n N_A_27_74#_c_908_n 0.0267093f $X=2.125 $Y=1.99 $X2=0 $Y2=0
cc_301 N_D_M1013_g N_A_27_74#_c_926_n 0.0123594f $X=2.52 $Y=2.525 $X2=0 $Y2=0
cc_302 N_D_M1032_g N_A_27_74#_M1004_g 0.00957963f $X=2.035 $Y=0.835 $X2=0 $Y2=0
cc_303 N_D_M1032_g N_A_27_74#_c_910_n 0.0267093f $X=2.035 $Y=0.835 $X2=0 $Y2=0
cc_304 D N_A_214_74#_M1016_g 2.98598e-19 $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_305 N_D_c_305_n N_A_214_74#_M1016_g 0.0246178f $X=2.125 $Y=1.99 $X2=0 $Y2=0
cc_306 N_D_M1032_g N_A_214_74#_c_1131_n 9.0931e-19 $X=2.035 $Y=0.835 $X2=0 $Y2=0
cc_307 D N_A_214_74#_c_1132_n 0.0135932f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_308 N_D_M1032_g N_A_214_74#_c_1133_n 0.0195775f $X=2.035 $Y=0.835 $X2=0 $Y2=0
cc_309 D N_A_214_74#_c_1133_n 0.0195142f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_310 N_D_c_305_n N_A_214_74#_c_1133_n 0.00398163f $X=2.125 $Y=1.99 $X2=0 $Y2=0
cc_311 N_D_M1032_g N_A_214_74#_c_1134_n 0.0213788f $X=2.035 $Y=0.835 $X2=0 $Y2=0
cc_312 N_D_c_305_n N_A_214_74#_c_1134_n 0.00967035f $X=2.125 $Y=1.99 $X2=0 $Y2=0
cc_313 N_D_M1013_g N_VPWR_c_1651_n 0.00434053f $X=2.52 $Y=2.525 $X2=0 $Y2=0
cc_314 D N_VPWR_c_1651_n 0.0190452f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_315 N_D_c_305_n N_VPWR_c_1651_n 0.0060958f $X=2.125 $Y=1.99 $X2=0 $Y2=0
cc_316 N_D_M1013_g N_VPWR_c_1649_n 0.00112709f $X=2.52 $Y=2.525 $X2=0 $Y2=0
cc_317 N_D_M1032_g N_A_422_125#_c_1795_n 0.00393226f $X=2.035 $Y=0.835 $X2=0
+ $Y2=0
cc_318 N_D_M1032_g N_A_422_125#_c_1797_n 0.00363027f $X=2.035 $Y=0.835 $X2=0
+ $Y2=0
cc_319 N_D_M1013_g N_A_422_125#_c_1799_n 0.0121735f $X=2.52 $Y=2.525 $X2=0 $Y2=0
cc_320 N_D_M1032_g N_A_422_125#_c_1798_n 0.00837482f $X=2.035 $Y=0.835 $X2=0
+ $Y2=0
cc_321 D N_A_422_125#_c_1798_n 0.0110926f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_322 N_D_c_305_n N_A_422_125#_c_1798_n 0.00570392f $X=2.125 $Y=1.99 $X2=0
+ $Y2=0
cc_323 N_D_M1032_g N_VGND_c_1904_n 0.00212205f $X=2.035 $Y=0.835 $X2=0 $Y2=0
cc_324 N_D_M1032_g N_VGND_c_1919_n 9.49986e-19 $X=2.035 $Y=0.835 $X2=0 $Y2=0
cc_325 N_A_671_93#_c_336_n N_SET_B_M1033_g 0.00828892f $X=3.43 $Y=1.125 $X2=0
+ $Y2=0
cc_326 N_A_671_93#_c_341_n N_SET_B_M1033_g 0.00327032f $X=3.59 $Y=1.29 $X2=0
+ $Y2=0
cc_327 N_A_671_93#_c_342_n N_SET_B_M1033_g 0.0138119f $X=3.59 $Y=1.29 $X2=0
+ $Y2=0
cc_328 N_A_671_93#_c_356_p N_SET_B_M1033_g 0.013805f $X=5.015 $Y=0.815 $X2=0
+ $Y2=0
cc_329 N_A_671_93#_c_344_n N_SET_B_M1033_g 5.74808e-19 $X=5.335 $Y=0.925 $X2=0
+ $Y2=0
cc_330 N_A_671_93#_M1009_g N_SET_B_M1020_g 0.0150044f $X=3.88 $Y=2.105 $X2=0
+ $Y2=0
cc_331 N_A_671_93#_c_350_n N_SET_B_M1020_g 0.00528862f $X=4.785 $Y=2.04 $X2=0
+ $Y2=0
cc_332 N_A_671_93#_c_352_n N_SET_B_M1020_g 0.00133435f $X=4.95 $Y=1.91 $X2=0
+ $Y2=0
cc_333 N_A_671_93#_M1009_g N_SET_B_c_500_n 0.00222581f $X=3.88 $Y=2.105 $X2=0
+ $Y2=0
cc_334 N_A_671_93#_c_350_n N_SET_B_c_500_n 0.0535111f $X=4.785 $Y=2.04 $X2=0
+ $Y2=0
cc_335 N_A_671_93#_c_352_n N_SET_B_c_500_n 0.0135407f $X=4.95 $Y=1.91 $X2=0
+ $Y2=0
cc_336 N_A_671_93#_c_350_n N_SET_B_c_501_n 0.0168382f $X=4.785 $Y=2.04 $X2=0
+ $Y2=0
cc_337 N_A_671_93#_c_350_n N_SET_B_c_503_n 0.0245375f $X=4.785 $Y=2.04 $X2=0
+ $Y2=0
cc_338 N_A_671_93#_M1003_g N_SET_B_c_526_n 0.0163036f $X=5.94 $Y=2.315 $X2=0
+ $Y2=0
cc_339 N_A_671_93#_c_351_n N_SET_B_c_526_n 0.0407208f $X=5.85 $Y=1.91 $X2=0
+ $Y2=0
cc_340 N_A_671_93#_c_345_n N_SET_B_c_526_n 0.00395021f $X=6.015 $Y=1.42 $X2=0
+ $Y2=0
cc_341 N_A_671_93#_c_347_n N_SET_B_c_526_n 6.8061e-19 $X=6.015 $Y=1.295 $X2=0
+ $Y2=0
cc_342 N_A_671_93#_c_350_n N_SET_B_c_530_n 0.0117007f $X=4.785 $Y=2.04 $X2=0
+ $Y2=0
cc_343 N_A_671_93#_c_351_n N_SET_B_c_530_n 0.0100071f $X=5.85 $Y=1.91 $X2=0
+ $Y2=0
cc_344 N_A_671_93#_M1003_g N_SET_B_c_504_n 0.00356579f $X=5.94 $Y=2.315 $X2=0
+ $Y2=0
cc_345 N_A_671_93#_c_342_n N_SET_B_c_494_n 2.53955e-19 $X=3.59 $Y=1.29 $X2=0
+ $Y2=0
cc_346 N_A_671_93#_M1009_g N_SET_B_c_496_n 0.0101593f $X=3.88 $Y=2.105 $X2=0
+ $Y2=0
cc_347 N_A_671_93#_c_350_n N_A_520_87#_M1035_g 0.0116313f $X=4.785 $Y=2.04 $X2=0
+ $Y2=0
cc_348 N_A_671_93#_c_351_n N_A_520_87#_M1035_g 0.0131068f $X=5.85 $Y=1.91 $X2=0
+ $Y2=0
cc_349 N_A_671_93#_c_352_n N_A_520_87#_M1035_g 0.00173127f $X=4.95 $Y=1.91 $X2=0
+ $Y2=0
cc_350 N_A_671_93#_c_336_n N_A_520_87#_c_656_n 0.00656686f $X=3.43 $Y=1.125
+ $X2=0 $Y2=0
cc_351 N_A_671_93#_c_379_p N_A_520_87#_c_656_n 0.00131642f $X=3.72 $Y=0.815
+ $X2=0 $Y2=0
cc_352 N_A_671_93#_c_336_n N_A_520_87#_c_657_n 0.00569157f $X=3.43 $Y=1.125
+ $X2=0 $Y2=0
cc_353 N_A_671_93#_M1009_g N_A_520_87#_c_657_n 0.00274152f $X=3.88 $Y=2.105
+ $X2=0 $Y2=0
cc_354 N_A_671_93#_c_341_n N_A_520_87#_c_657_n 0.0406769f $X=3.59 $Y=1.29 $X2=0
+ $Y2=0
cc_355 N_A_671_93#_c_379_p N_A_520_87#_c_657_n 0.0121462f $X=3.72 $Y=0.815 $X2=0
+ $Y2=0
cc_356 N_A_671_93#_M1009_g N_A_520_87#_c_666_n 0.00183175f $X=3.88 $Y=2.105
+ $X2=0 $Y2=0
cc_357 N_A_671_93#_M1009_g N_A_520_87#_c_658_n 0.0187049f $X=3.88 $Y=2.105 $X2=0
+ $Y2=0
cc_358 N_A_671_93#_c_341_n N_A_520_87#_c_658_n 0.0202187f $X=3.59 $Y=1.29 $X2=0
+ $Y2=0
cc_359 N_A_671_93#_c_342_n N_A_520_87#_c_658_n 0.00469367f $X=3.59 $Y=1.29 $X2=0
+ $Y2=0
cc_360 N_A_671_93#_M1009_g N_A_520_87#_c_659_n 0.00509465f $X=3.88 $Y=2.105
+ $X2=0 $Y2=0
cc_361 N_A_671_93#_c_341_n N_A_520_87#_c_659_n 0.0152467f $X=3.59 $Y=1.29 $X2=0
+ $Y2=0
cc_362 N_A_671_93#_c_342_n N_A_520_87#_c_659_n 0.00598734f $X=3.59 $Y=1.29 $X2=0
+ $Y2=0
cc_363 N_A_671_93#_c_356_p N_A_520_87#_c_660_n 0.0534303f $X=5.015 $Y=0.815
+ $X2=0 $Y2=0
cc_364 N_A_671_93#_c_351_n N_A_520_87#_c_660_n 0.00813741f $X=5.85 $Y=1.91 $X2=0
+ $Y2=0
cc_365 N_A_671_93#_c_352_n N_A_520_87#_c_660_n 0.0153161f $X=4.95 $Y=1.91 $X2=0
+ $Y2=0
cc_366 N_A_671_93#_c_344_n N_A_520_87#_c_660_n 0.00259022f $X=5.335 $Y=0.925
+ $X2=0 $Y2=0
cc_367 N_A_671_93#_c_341_n N_A_520_87#_c_661_n 0.014307f $X=3.59 $Y=1.29 $X2=0
+ $Y2=0
cc_368 N_A_671_93#_c_342_n N_A_520_87#_c_661_n 0.0011591f $X=3.59 $Y=1.29 $X2=0
+ $Y2=0
cc_369 N_A_671_93#_c_356_p N_A_520_87#_c_661_n 0.0139549f $X=5.015 $Y=0.815
+ $X2=0 $Y2=0
cc_370 N_A_671_93#_c_342_n N_A_520_87#_c_662_n 0.00305459f $X=3.59 $Y=1.29 $X2=0
+ $Y2=0
cc_371 N_A_671_93#_c_356_p N_A_520_87#_c_663_n 4.11778e-19 $X=5.015 $Y=0.815
+ $X2=0 $Y2=0
cc_372 N_A_671_93#_c_352_n N_A_520_87#_c_663_n 0.00113523f $X=4.95 $Y=1.91 $X2=0
+ $Y2=0
cc_373 N_A_671_93#_c_356_p N_A_520_87#_c_664_n 0.00948817f $X=5.015 $Y=0.815
+ $X2=0 $Y2=0
cc_374 N_A_671_93#_c_344_n N_A_520_87#_c_664_n 0.00360733f $X=5.335 $Y=0.925
+ $X2=0 $Y2=0
cc_375 N_A_671_93#_M1003_g N_A_1062_93#_M1011_g 0.036113f $X=5.94 $Y=2.315 $X2=0
+ $Y2=0
cc_376 N_A_671_93#_c_350_n N_A_1062_93#_M1011_g 0.00109562f $X=4.785 $Y=2.04
+ $X2=0 $Y2=0
cc_377 N_A_671_93#_c_351_n N_A_1062_93#_M1011_g 0.0121906f $X=5.85 $Y=1.91 $X2=0
+ $Y2=0
cc_378 N_A_671_93#_c_406_p N_A_1062_93#_M1011_g 0.00148114f $X=5.935 $Y=1.825
+ $X2=0 $Y2=0
cc_379 N_A_671_93#_c_339_n N_A_1062_93#_c_764_n 0.0198682f $X=6.44 $Y=1.295
+ $X2=0 $Y2=0
cc_380 N_A_671_93#_c_351_n N_A_1062_93#_c_764_n 0.00631979f $X=5.85 $Y=1.91
+ $X2=0 $Y2=0
cc_381 N_A_671_93#_c_343_n N_A_1062_93#_c_764_n 0.00798804f $X=5.85 $Y=0.925
+ $X2=0 $Y2=0
cc_382 N_A_671_93#_c_345_n N_A_1062_93#_c_764_n 0.025397f $X=6.015 $Y=1.42 $X2=0
+ $Y2=0
cc_383 N_A_671_93#_c_346_n N_A_1062_93#_c_764_n 0.00954547f $X=6.015 $Y=1.255
+ $X2=0 $Y2=0
cc_384 N_A_671_93#_c_347_n N_A_1062_93#_c_764_n 0.00372139f $X=6.015 $Y=1.295
+ $X2=0 $Y2=0
cc_385 N_A_671_93#_c_351_n N_A_1062_93#_c_765_n 0.00223748f $X=5.85 $Y=1.91
+ $X2=0 $Y2=0
cc_386 N_A_671_93#_c_343_n N_A_1062_93#_c_765_n 0.00322139f $X=5.85 $Y=0.925
+ $X2=0 $Y2=0
cc_387 N_A_671_93#_c_345_n N_A_1062_93#_c_765_n 0.00128921f $X=6.015 $Y=1.42
+ $X2=0 $Y2=0
cc_388 N_A_671_93#_c_346_n N_A_1062_93#_c_765_n 0.00129148f $X=6.015 $Y=1.255
+ $X2=0 $Y2=0
cc_389 N_A_671_93#_c_347_n N_A_1062_93#_c_765_n 7.67181e-19 $X=6.015 $Y=1.295
+ $X2=0 $Y2=0
cc_390 N_A_671_93#_c_351_n N_A_1062_93#_c_766_n 0.017358f $X=5.85 $Y=1.91 $X2=0
+ $Y2=0
cc_391 N_A_671_93#_c_343_n N_A_1062_93#_c_766_n 0.0181773f $X=5.85 $Y=0.925
+ $X2=0 $Y2=0
cc_392 N_A_671_93#_c_344_n N_A_1062_93#_c_766_n 0.00188106f $X=5.335 $Y=0.925
+ $X2=0 $Y2=0
cc_393 N_A_671_93#_c_346_n N_A_1062_93#_c_766_n 0.0230094f $X=6.015 $Y=1.255
+ $X2=0 $Y2=0
cc_394 N_A_671_93#_c_347_n N_A_1062_93#_c_766_n 0.00141195f $X=6.015 $Y=1.295
+ $X2=0 $Y2=0
cc_395 N_A_671_93#_c_351_n N_A_1062_93#_c_769_n 9.67991e-19 $X=5.85 $Y=1.91
+ $X2=0 $Y2=0
cc_396 N_A_671_93#_c_343_n N_A_1062_93#_c_769_n 9.21407e-19 $X=5.85 $Y=0.925
+ $X2=0 $Y2=0
cc_397 N_A_671_93#_c_345_n N_A_1062_93#_c_769_n 0.00110037f $X=6.015 $Y=1.42
+ $X2=0 $Y2=0
cc_398 N_A_671_93#_c_347_n N_A_1062_93#_c_769_n 0.0215457f $X=6.015 $Y=1.295
+ $X2=0 $Y2=0
cc_399 N_A_671_93#_c_343_n N_A_1062_93#_c_770_n 0.00971016f $X=5.85 $Y=0.925
+ $X2=0 $Y2=0
cc_400 N_A_671_93#_c_344_n N_A_1062_93#_c_770_n 0.00976139f $X=5.335 $Y=0.925
+ $X2=0 $Y2=0
cc_401 N_A_671_93#_c_346_n N_A_1062_93#_c_770_n 0.00482672f $X=6.015 $Y=1.255
+ $X2=0 $Y2=0
cc_402 N_A_671_93#_c_347_n N_A_1062_93#_c_770_n 0.00110364f $X=6.015 $Y=1.295
+ $X2=0 $Y2=0
cc_403 N_A_671_93#_M1009_g N_A_27_74#_M1039_g 0.0413784f $X=3.88 $Y=2.105 $X2=0
+ $Y2=0
cc_404 N_A_671_93#_c_342_n N_A_27_74#_M1039_g 0.00720464f $X=3.59 $Y=1.29 $X2=0
+ $Y2=0
cc_405 N_A_671_93#_M1009_g N_A_27_74#_c_929_n 0.00384162f $X=3.88 $Y=2.105 $X2=0
+ $Y2=0
cc_406 N_A_671_93#_M1003_g N_A_27_74#_c_929_n 0.0124167f $X=5.94 $Y=2.315 $X2=0
+ $Y2=0
cc_407 N_A_671_93#_M1003_g N_A_27_74#_c_919_n 0.00113329f $X=5.94 $Y=2.315 $X2=0
+ $Y2=0
cc_408 N_A_671_93#_c_339_n N_A_27_74#_c_919_n 0.00113069f $X=6.44 $Y=1.295 $X2=0
+ $Y2=0
cc_409 N_A_671_93#_c_351_n N_A_27_74#_c_919_n 0.00441009f $X=5.85 $Y=1.91 $X2=0
+ $Y2=0
cc_410 N_A_671_93#_c_406_p N_A_27_74#_c_919_n 0.00737995f $X=5.935 $Y=1.825
+ $X2=0 $Y2=0
cc_411 N_A_671_93#_M1003_g N_A_27_74#_c_920_n 0.0372909f $X=5.94 $Y=2.315 $X2=0
+ $Y2=0
cc_412 N_A_671_93#_c_339_n N_A_27_74#_c_920_n 0.011622f $X=6.44 $Y=1.295 $X2=0
+ $Y2=0
cc_413 N_A_671_93#_c_351_n N_A_27_74#_c_920_n 8.09982e-19 $X=5.85 $Y=1.91 $X2=0
+ $Y2=0
cc_414 N_A_671_93#_c_406_p N_A_27_74#_c_920_n 9.19564e-19 $X=5.935 $Y=1.825
+ $X2=0 $Y2=0
cc_415 N_A_671_93#_M1003_g N_A_27_74#_c_921_n 3.5569e-19 $X=5.94 $Y=2.315 $X2=0
+ $Y2=0
cc_416 N_A_671_93#_c_340_n N_A_27_74#_c_921_n 0.00527455f $X=6.515 $Y=1.22 $X2=0
+ $Y2=0
cc_417 N_A_671_93#_c_406_p N_A_27_74#_c_921_n 6.80646e-19 $X=5.935 $Y=1.825
+ $X2=0 $Y2=0
cc_418 N_A_671_93#_c_345_n N_A_27_74#_c_921_n 0.0110962f $X=6.015 $Y=1.42 $X2=0
+ $Y2=0
cc_419 N_A_671_93#_c_346_n N_A_27_74#_c_921_n 0.00391001f $X=6.015 $Y=1.255
+ $X2=0 $Y2=0
cc_420 N_A_671_93#_c_347_n N_A_27_74#_c_921_n 0.00400932f $X=6.015 $Y=1.295
+ $X2=0 $Y2=0
cc_421 N_A_671_93#_c_336_n N_A_214_74#_M1025_g 0.0238128f $X=3.43 $Y=1.125 $X2=0
+ $Y2=0
cc_422 N_A_671_93#_c_336_n N_A_214_74#_c_1124_n 0.0102834f $X=3.43 $Y=1.125
+ $X2=0 $Y2=0
cc_423 N_A_671_93#_c_340_n N_A_214_74#_c_1124_n 0.0104164f $X=6.515 $Y=1.22
+ $X2=0 $Y2=0
cc_424 N_A_671_93#_c_356_p N_A_214_74#_c_1124_n 0.00342121f $X=5.015 $Y=0.815
+ $X2=0 $Y2=0
cc_425 N_A_671_93#_c_379_p N_A_214_74#_c_1124_n 7.47729e-19 $X=3.72 $Y=0.815
+ $X2=0 $Y2=0
cc_426 N_A_671_93#_c_343_n N_A_214_74#_c_1124_n 0.0057641f $X=5.85 $Y=0.925
+ $X2=0 $Y2=0
cc_427 N_A_671_93#_c_340_n N_A_214_74#_M1012_g 0.0248811f $X=6.515 $Y=1.22 $X2=0
+ $Y2=0
cc_428 N_A_671_93#_c_342_n N_A_214_74#_c_1127_n 0.00785896f $X=3.59 $Y=1.29
+ $X2=0 $Y2=0
cc_429 N_A_671_93#_c_339_n N_A_214_74#_c_1128_n 0.0248811f $X=6.44 $Y=1.295
+ $X2=0 $Y2=0
cc_430 N_A_671_93#_M1003_g N_A_1314_424#_c_1448_n 2.07201e-19 $X=5.94 $Y=2.315
+ $X2=0 $Y2=0
cc_431 N_A_671_93#_M1003_g N_A_1314_424#_c_1450_n 3.4362e-19 $X=5.94 $Y=2.315
+ $X2=0 $Y2=0
cc_432 N_A_671_93#_c_351_n N_VPWR_M1011_d 0.00230172f $X=5.85 $Y=1.91 $X2=0
+ $Y2=0
cc_433 N_A_671_93#_M1009_g N_VPWR_c_1652_n 0.0110678f $X=3.88 $Y=2.105 $X2=0
+ $Y2=0
cc_434 N_A_671_93#_M1003_g N_VPWR_c_1653_n 0.0059978f $X=5.94 $Y=2.315 $X2=0
+ $Y2=0
cc_435 N_A_671_93#_M1009_g N_VPWR_c_1649_n 9.48371e-19 $X=3.88 $Y=2.105 $X2=0
+ $Y2=0
cc_436 N_A_671_93#_M1003_g N_VPWR_c_1649_n 0.00100812f $X=5.94 $Y=2.315 $X2=0
+ $Y2=0
cc_437 N_A_671_93#_c_351_n A_1020_379# 0.00130751f $X=5.85 $Y=1.91 $X2=-0.19
+ $Y2=-0.245
cc_438 N_A_671_93#_c_341_n N_VGND_M1036_d 0.001911f $X=3.59 $Y=1.29 $X2=0 $Y2=0
cc_439 N_A_671_93#_c_356_p N_VGND_M1036_d 0.0118141f $X=5.015 $Y=0.815 $X2=0
+ $Y2=0
cc_440 N_A_671_93#_c_379_p N_VGND_M1036_d 0.00183319f $X=3.72 $Y=0.815 $X2=0
+ $Y2=0
cc_441 N_A_671_93#_c_340_n N_VGND_c_1905_n 0.00570252f $X=6.515 $Y=1.22 $X2=0
+ $Y2=0
cc_442 N_A_671_93#_c_339_n N_VGND_c_1935_n 0.00900609f $X=6.44 $Y=1.295 $X2=0
+ $Y2=0
cc_443 N_A_671_93#_c_343_n N_VGND_c_1935_n 0.0144604f $X=5.85 $Y=0.925 $X2=0
+ $Y2=0
cc_444 N_A_671_93#_c_346_n N_VGND_c_1935_n 0.00565417f $X=6.015 $Y=1.255 $X2=0
+ $Y2=0
cc_445 N_A_671_93#_c_356_p N_VGND_c_1909_n 0.00283998f $X=5.015 $Y=0.815 $X2=0
+ $Y2=0
cc_446 N_A_671_93#_c_345_n N_VGND_c_1911_n 0.00189302f $X=6.015 $Y=1.42 $X2=0
+ $Y2=0
cc_447 N_A_671_93#_c_347_n N_VGND_c_1911_n 0.00248751f $X=6.015 $Y=1.295 $X2=0
+ $Y2=0
cc_448 N_A_671_93#_c_336_n N_VGND_c_1915_n 0.00136819f $X=3.43 $Y=1.125 $X2=0
+ $Y2=0
cc_449 N_A_671_93#_c_342_n N_VGND_c_1915_n 6.15763e-19 $X=3.59 $Y=1.29 $X2=0
+ $Y2=0
cc_450 N_A_671_93#_c_356_p N_VGND_c_1915_n 0.0339583f $X=5.015 $Y=0.815 $X2=0
+ $Y2=0
cc_451 N_A_671_93#_c_379_p N_VGND_c_1915_n 0.0147547f $X=3.72 $Y=0.815 $X2=0
+ $Y2=0
cc_452 N_A_671_93#_c_336_n N_VGND_c_1919_n 9.39239e-19 $X=3.43 $Y=1.125 $X2=0
+ $Y2=0
cc_453 N_A_671_93#_c_340_n N_VGND_c_1919_n 9.39239e-19 $X=6.515 $Y=1.22 $X2=0
+ $Y2=0
cc_454 N_A_671_93#_c_356_p N_VGND_c_1919_n 0.00860021f $X=5.015 $Y=0.815 $X2=0
+ $Y2=0
cc_455 N_A_671_93#_c_379_p N_VGND_c_1919_n 0.00299379f $X=3.72 $Y=0.815 $X2=0
+ $Y2=0
cc_456 N_A_671_93#_c_343_n N_VGND_c_1919_n 0.00734385f $X=5.85 $Y=0.925 $X2=0
+ $Y2=0
cc_457 N_A_671_93#_c_356_p N_A_872_119#_M1033_d 0.00925221f $X=5.015 $Y=0.815
+ $X2=-0.19 $Y2=-0.245
cc_458 N_A_671_93#_c_343_n N_A_872_119#_M1030_d 0.00779711f $X=5.85 $Y=0.925
+ $X2=0 $Y2=0
cc_459 N_A_671_93#_c_356_p N_A_872_119#_c_2063_n 0.00694096f $X=5.015 $Y=0.815
+ $X2=0 $Y2=0
cc_460 N_A_671_93#_c_343_n N_A_872_119#_c_2063_n 0.00499238f $X=5.85 $Y=0.925
+ $X2=0 $Y2=0
cc_461 N_A_671_93#_c_344_n N_A_872_119#_c_2063_n 0.019569f $X=5.335 $Y=0.925
+ $X2=0 $Y2=0
cc_462 N_A_671_93#_c_356_p N_A_872_119#_c_2064_n 0.0300357f $X=5.015 $Y=0.815
+ $X2=0 $Y2=0
cc_463 N_A_671_93#_c_343_n N_A_872_119#_c_2065_n 0.0238389f $X=5.85 $Y=0.925
+ $X2=0 $Y2=0
cc_464 N_SET_B_c_500_n N_A_520_87#_M1035_g 0.00186845f $X=4.445 $Y=2.905 $X2=0
+ $Y2=0
cc_465 N_SET_B_c_501_n N_A_520_87#_M1035_g 0.00396457f $X=5.16 $Y=2.99 $X2=0
+ $Y2=0
cc_466 N_SET_B_c_503_n N_A_520_87#_M1035_g 0.00442072f $X=5.245 $Y=2.905 $X2=0
+ $Y2=0
cc_467 N_SET_B_c_530_n N_A_520_87#_M1035_g 0.00143241f $X=5.33 $Y=2.25 $X2=0
+ $Y2=0
cc_468 N_SET_B_c_494_n N_A_520_87#_M1035_g 4.1388e-19 $X=4.445 $Y=1.532 $X2=0
+ $Y2=0
cc_469 N_SET_B_c_496_n N_A_520_87#_M1035_g 0.0272139f $X=4.47 $Y=1.53 $X2=0
+ $Y2=0
cc_470 N_SET_B_M1020_g N_A_520_87#_c_658_n 4.64982e-19 $X=4.47 $Y=2.315 $X2=0
+ $Y2=0
cc_471 N_SET_B_c_500_n N_A_520_87#_c_658_n 0.00779985f $X=4.445 $Y=2.905 $X2=0
+ $Y2=0
cc_472 N_SET_B_c_494_n N_A_520_87#_c_658_n 0.00245753f $X=4.445 $Y=1.532 $X2=0
+ $Y2=0
cc_473 N_SET_B_c_496_n N_A_520_87#_c_658_n 5.85823e-19 $X=4.47 $Y=1.53 $X2=0
+ $Y2=0
cc_474 N_SET_B_M1033_g N_A_520_87#_c_659_n 0.00497141f $X=4.285 $Y=0.87 $X2=0
+ $Y2=0
cc_475 N_SET_B_c_494_n N_A_520_87#_c_659_n 0.0161246f $X=4.445 $Y=1.532 $X2=0
+ $Y2=0
cc_476 N_SET_B_M1033_g N_A_520_87#_c_660_n 0.015008f $X=4.285 $Y=0.87 $X2=0
+ $Y2=0
cc_477 N_SET_B_c_494_n N_A_520_87#_c_660_n 0.0368787f $X=4.445 $Y=1.532 $X2=0
+ $Y2=0
cc_478 N_SET_B_c_496_n N_A_520_87#_c_660_n 0.00713696f $X=4.47 $Y=1.53 $X2=0
+ $Y2=0
cc_479 N_SET_B_M1033_g N_A_520_87#_c_663_n 0.00275729f $X=4.285 $Y=0.87 $X2=0
+ $Y2=0
cc_480 N_SET_B_c_494_n N_A_520_87#_c_663_n 2.07915e-19 $X=4.445 $Y=1.532 $X2=0
+ $Y2=0
cc_481 N_SET_B_c_496_n N_A_520_87#_c_663_n 0.0141879f $X=4.47 $Y=1.53 $X2=0
+ $Y2=0
cc_482 N_SET_B_M1033_g N_A_520_87#_c_664_n 0.0168362f $X=4.285 $Y=0.87 $X2=0
+ $Y2=0
cc_483 N_SET_B_c_503_n N_A_1062_93#_M1011_g 0.00262459f $X=5.245 $Y=2.905 $X2=0
+ $Y2=0
cc_484 N_SET_B_c_526_n N_A_1062_93#_M1011_g 0.0157762f $X=6.04 $Y=2.25 $X2=0
+ $Y2=0
cc_485 N_SET_B_M1034_g N_A_1062_93#_c_764_n 0.00213786f $X=8.465 $Y=0.74 $X2=0
+ $Y2=0
cc_486 N_SET_B_c_508_n N_A_1062_93#_c_764_n 0.00560703f $X=8.24 $Y=1.825 $X2=0
+ $Y2=0
cc_487 SET_B N_A_1062_93#_c_764_n 0.00844095f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_488 N_SET_B_M1020_g N_A_27_74#_c_929_n 0.011501f $X=4.47 $Y=2.315 $X2=0 $Y2=0
cc_489 N_SET_B_c_501_n N_A_27_74#_c_929_n 0.0154848f $X=5.16 $Y=2.99 $X2=0 $Y2=0
cc_490 N_SET_B_c_502_n N_A_27_74#_c_929_n 0.00169616f $X=4.53 $Y=2.99 $X2=0
+ $Y2=0
cc_491 N_SET_B_c_505_n N_A_27_74#_c_929_n 0.00211038f $X=7.28 $Y=2.99 $X2=0
+ $Y2=0
cc_492 N_SET_B_c_506_n N_A_27_74#_c_929_n 0.00420304f $X=6.21 $Y=2.99 $X2=0
+ $Y2=0
cc_493 N_SET_B_c_526_n N_A_27_74#_M1005_g 0.00166795f $X=6.04 $Y=2.25 $X2=0
+ $Y2=0
cc_494 N_SET_B_c_504_n N_A_27_74#_M1005_g 0.00741364f $X=6.125 $Y=2.905 $X2=0
+ $Y2=0
cc_495 N_SET_B_c_505_n N_A_27_74#_M1005_g 0.0173018f $X=7.28 $Y=2.99 $X2=0 $Y2=0
cc_496 N_SET_B_M1033_g N_A_214_74#_c_1124_n 0.00991925f $X=4.285 $Y=0.87 $X2=0
+ $Y2=0
cc_497 N_SET_B_c_505_n N_A_214_74#_M1001_g 0.0130081f $X=7.28 $Y=2.99 $X2=0
+ $Y2=0
cc_498 N_SET_B_c_507_n N_A_214_74#_M1001_g 0.00672345f $X=7.365 $Y=2.905 $X2=0
+ $Y2=0
cc_499 N_SET_B_c_507_n N_A_214_74#_c_1129_n 0.00347575f $X=7.365 $Y=2.905 $X2=0
+ $Y2=0
cc_500 N_SET_B_c_509_n N_A_214_74#_c_1129_n 0.00176185f $X=7.45 $Y=1.825 $X2=0
+ $Y2=0
cc_501 N_SET_B_c_505_n N_A_1474_446#_M1015_g 0.00488481f $X=7.28 $Y=2.99 $X2=0
+ $Y2=0
cc_502 N_SET_B_c_507_n N_A_1474_446#_M1015_g 0.0189067f $X=7.365 $Y=2.905 $X2=0
+ $Y2=0
cc_503 N_SET_B_M1023_g N_A_1474_446#_c_1271_n 0.0136746f $X=8.48 $Y=2.46 $X2=0
+ $Y2=0
cc_504 N_SET_B_c_507_n N_A_1474_446#_c_1271_n 0.00269073f $X=7.365 $Y=2.905
+ $X2=0 $Y2=0
cc_505 N_SET_B_c_508_n N_A_1474_446#_c_1271_n 0.00319331f $X=8.24 $Y=1.825 $X2=0
+ $Y2=0
cc_506 N_SET_B_M1034_g N_A_1474_446#_M1021_g 0.0263478f $X=8.465 $Y=0.74 $X2=0
+ $Y2=0
cc_507 SET_B N_A_1474_446#_M1021_g 0.00125179f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_508 N_SET_B_c_497_n N_A_1474_446#_M1021_g 0.0204448f $X=8.405 $Y=1.635 $X2=0
+ $Y2=0
cc_509 N_SET_B_M1023_g N_A_1474_446#_c_1276_n 0.00273304f $X=8.48 $Y=2.46 $X2=0
+ $Y2=0
cc_510 N_SET_B_c_508_n N_A_1474_446#_c_1276_n 0.0111733f $X=8.24 $Y=1.825 $X2=0
+ $Y2=0
cc_511 N_SET_B_c_507_n N_A_1474_446#_c_1277_n 0.00696429f $X=7.365 $Y=2.905
+ $X2=0 $Y2=0
cc_512 N_SET_B_c_508_n N_A_1474_446#_c_1277_n 0.00974498f $X=8.24 $Y=1.825 $X2=0
+ $Y2=0
cc_513 N_SET_B_M1023_g N_A_1474_446#_c_1278_n 0.00875105f $X=8.48 $Y=2.46 $X2=0
+ $Y2=0
cc_514 SET_B N_A_1474_446#_c_1267_n 0.00683367f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_515 N_SET_B_M1023_g N_A_1474_446#_c_1282_n 0.0243251f $X=8.48 $Y=2.46 $X2=0
+ $Y2=0
cc_516 N_SET_B_c_507_n N_A_1474_446#_c_1282_n 0.0232576f $X=7.365 $Y=2.905 $X2=0
+ $Y2=0
cc_517 N_SET_B_c_508_n N_A_1474_446#_c_1282_n 0.0466911f $X=8.24 $Y=1.825 $X2=0
+ $Y2=0
cc_518 SET_B N_A_1474_446#_c_1282_n 0.0225793f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_519 N_SET_B_c_497_n N_A_1474_446#_c_1282_n 7.20549e-19 $X=8.405 $Y=1.635
+ $X2=0 $Y2=0
cc_520 N_SET_B_M1023_g N_A_1474_446#_c_1302_n 0.00415444f $X=8.48 $Y=2.46 $X2=0
+ $Y2=0
cc_521 N_SET_B_c_505_n N_A_1314_424#_M1005_d 0.00256188f $X=7.28 $Y=2.99 $X2=0
+ $Y2=0
cc_522 SET_B N_A_1314_424#_M1010_g 0.00162477f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_523 N_SET_B_c_497_n N_A_1314_424#_M1010_g 0.0344008f $X=8.405 $Y=1.635 $X2=0
+ $Y2=0
cc_524 N_SET_B_c_526_n N_A_1314_424#_c_1448_n 0.00272807f $X=6.04 $Y=2.25 $X2=0
+ $Y2=0
cc_525 N_SET_B_c_504_n N_A_1314_424#_c_1448_n 0.0177173f $X=6.125 $Y=2.905 $X2=0
+ $Y2=0
cc_526 N_SET_B_c_505_n N_A_1314_424#_c_1448_n 0.0197579f $X=7.28 $Y=2.99 $X2=0
+ $Y2=0
cc_527 N_SET_B_c_507_n N_A_1314_424#_c_1448_n 0.0148375f $X=7.365 $Y=2.905 $X2=0
+ $Y2=0
cc_528 N_SET_B_c_507_n N_A_1314_424#_c_1440_n 0.0142669f $X=7.365 $Y=2.905 $X2=0
+ $Y2=0
cc_529 N_SET_B_c_509_n N_A_1314_424#_c_1440_n 0.0137158f $X=7.45 $Y=1.825 $X2=0
+ $Y2=0
cc_530 N_SET_B_c_508_n N_A_1314_424#_c_1441_n 0.0315946f $X=8.24 $Y=1.825 $X2=0
+ $Y2=0
cc_531 N_SET_B_c_509_n N_A_1314_424#_c_1441_n 0.0135027f $X=7.45 $Y=1.825 $X2=0
+ $Y2=0
cc_532 N_SET_B_M1034_g N_A_1314_424#_c_1442_n 0.0147584f $X=8.465 $Y=0.74 $X2=0
+ $Y2=0
cc_533 N_SET_B_c_508_n N_A_1314_424#_c_1442_n 0.00414643f $X=8.24 $Y=1.825 $X2=0
+ $Y2=0
cc_534 SET_B N_A_1314_424#_c_1442_n 0.0265108f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_535 N_SET_B_c_497_n N_A_1314_424#_c_1442_n 0.00118239f $X=8.405 $Y=1.635
+ $X2=0 $Y2=0
cc_536 N_SET_B_c_526_n N_A_1314_424#_c_1450_n 0.00588951f $X=6.04 $Y=2.25 $X2=0
+ $Y2=0
cc_537 N_SET_B_c_505_n N_A_1314_424#_c_1450_n 0.00507182f $X=7.28 $Y=2.99 $X2=0
+ $Y2=0
cc_538 N_SET_B_c_507_n N_A_1314_424#_c_1450_n 0.013197f $X=7.365 $Y=2.905 $X2=0
+ $Y2=0
cc_539 N_SET_B_M1034_g N_A_1314_424#_c_1444_n 0.00284277f $X=8.465 $Y=0.74 $X2=0
+ $Y2=0
cc_540 N_SET_B_c_508_n N_A_1314_424#_c_1444_n 0.0120262f $X=8.24 $Y=1.825 $X2=0
+ $Y2=0
cc_541 SET_B N_A_1314_424#_c_1444_n 0.00755271f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_542 N_SET_B_c_497_n N_A_1314_424#_c_1444_n 2.92299e-19 $X=8.405 $Y=1.635
+ $X2=0 $Y2=0
cc_543 N_SET_B_M1034_g N_A_1314_424#_c_1445_n 0.0141555f $X=8.465 $Y=0.74 $X2=0
+ $Y2=0
cc_544 SET_B N_A_1314_424#_c_1445_n 2.7904e-19 $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_545 N_SET_B_c_497_n N_A_1314_424#_c_1445_n 0.00503224f $X=8.405 $Y=1.635
+ $X2=0 $Y2=0
cc_546 N_SET_B_M1034_g N_A_1314_424#_c_1446_n 0.0184908f $X=8.465 $Y=0.74 $X2=0
+ $Y2=0
cc_547 N_SET_B_c_526_n N_VPWR_M1011_d 0.00453815f $X=6.04 $Y=2.25 $X2=0 $Y2=0
cc_548 N_SET_B_M1020_g N_VPWR_c_1652_n 0.00461962f $X=4.47 $Y=2.315 $X2=0 $Y2=0
cc_549 N_SET_B_c_500_n N_VPWR_c_1652_n 0.0427355f $X=4.445 $Y=2.905 $X2=0 $Y2=0
cc_550 N_SET_B_c_502_n N_VPWR_c_1652_n 0.0147459f $X=4.53 $Y=2.99 $X2=0 $Y2=0
cc_551 N_SET_B_c_501_n N_VPWR_c_1653_n 0.0151625f $X=5.16 $Y=2.99 $X2=0 $Y2=0
cc_552 N_SET_B_c_503_n N_VPWR_c_1653_n 0.0217628f $X=5.245 $Y=2.905 $X2=0 $Y2=0
cc_553 N_SET_B_c_526_n N_VPWR_c_1653_n 0.0203498f $X=6.04 $Y=2.25 $X2=0 $Y2=0
cc_554 N_SET_B_c_504_n N_VPWR_c_1653_n 0.0217628f $X=6.125 $Y=2.905 $X2=0 $Y2=0
cc_555 N_SET_B_c_506_n N_VPWR_c_1653_n 0.0151624f $X=6.21 $Y=2.99 $X2=0 $Y2=0
cc_556 N_SET_B_M1023_g N_VPWR_c_1657_n 0.00460063f $X=8.48 $Y=2.46 $X2=0 $Y2=0
cc_557 N_SET_B_c_501_n N_VPWR_c_1661_n 0.0521009f $X=5.16 $Y=2.99 $X2=0 $Y2=0
cc_558 N_SET_B_c_502_n N_VPWR_c_1661_n 0.0115893f $X=4.53 $Y=2.99 $X2=0 $Y2=0
cc_559 N_SET_B_M1023_g N_VPWR_c_1649_n 0.00904612f $X=8.48 $Y=2.46 $X2=0 $Y2=0
cc_560 N_SET_B_c_501_n N_VPWR_c_1649_n 0.0269995f $X=5.16 $Y=2.99 $X2=0 $Y2=0
cc_561 N_SET_B_c_502_n N_VPWR_c_1649_n 0.00583135f $X=4.53 $Y=2.99 $X2=0 $Y2=0
cc_562 N_SET_B_c_505_n N_VPWR_c_1649_n 0.044075f $X=7.28 $Y=2.99 $X2=0 $Y2=0
cc_563 N_SET_B_c_506_n N_VPWR_c_1649_n 0.00583135f $X=6.21 $Y=2.99 $X2=0 $Y2=0
cc_564 N_SET_B_c_505_n N_VPWR_c_1670_n 0.0796923f $X=7.28 $Y=2.99 $X2=0 $Y2=0
cc_565 N_SET_B_c_506_n N_VPWR_c_1670_n 0.0115893f $X=6.21 $Y=2.99 $X2=0 $Y2=0
cc_566 N_SET_B_M1023_g N_VPWR_c_1671_n 0.0111395f $X=8.48 $Y=2.46 $X2=0 $Y2=0
cc_567 N_SET_B_c_505_n N_VPWR_c_1671_n 0.0150587f $X=7.28 $Y=2.99 $X2=0 $Y2=0
cc_568 N_SET_B_c_507_n N_VPWR_c_1671_n 0.0200141f $X=7.365 $Y=2.905 $X2=0 $Y2=0
cc_569 N_SET_B_c_503_n A_1020_379# 0.00501624f $X=5.245 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_570 N_SET_B_c_530_n A_1020_379# 0.00292905f $X=5.33 $Y=2.25 $X2=-0.19
+ $Y2=-0.245
cc_571 N_SET_B_c_526_n A_1206_379# 0.00496097f $X=6.04 $Y=2.25 $X2=-0.19
+ $Y2=-0.245
cc_572 N_SET_B_c_504_n A_1206_379# 0.00851041f $X=6.125 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_573 N_SET_B_c_505_n A_1206_379# 0.00465498f $X=7.28 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_574 N_SET_B_c_506_n A_1206_379# 2.13099e-19 $X=6.21 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_575 N_SET_B_c_505_n A_1421_508# 0.0044642f $X=7.28 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_576 N_SET_B_c_507_n A_1421_508# 0.00432504f $X=7.365 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_577 N_SET_B_M1034_g N_VGND_c_1906_n 0.00989595f $X=8.465 $Y=0.74 $X2=0 $Y2=0
cc_578 N_SET_B_M1033_g N_VGND_c_1915_n 0.00136121f $X=4.285 $Y=0.87 $X2=0 $Y2=0
cc_579 N_SET_B_M1034_g N_VGND_c_1917_n 0.00383152f $X=8.465 $Y=0.74 $X2=0 $Y2=0
cc_580 N_SET_B_M1033_g N_VGND_c_1919_n 9.39239e-19 $X=4.285 $Y=0.87 $X2=0 $Y2=0
cc_581 N_SET_B_M1034_g N_VGND_c_1919_n 0.00758251f $X=8.465 $Y=0.74 $X2=0 $Y2=0
cc_582 N_SET_B_M1033_g N_A_872_119#_c_2064_n 0.00114548f $X=4.285 $Y=0.87 $X2=0
+ $Y2=0
cc_583 N_SET_B_M1034_g N_A_1708_74#_c_2094_n 0.00133752f $X=8.465 $Y=0.74 $X2=0
+ $Y2=0
cc_584 N_A_520_87#_M1035_g N_A_1062_93#_M1011_g 0.0650816f $X=5.01 $Y=2.315
+ $X2=0 $Y2=0
cc_585 N_A_520_87#_c_660_n N_A_1062_93#_c_765_n 0.00139777f $X=4.745 $Y=1.155
+ $X2=0 $Y2=0
cc_586 N_A_520_87#_c_660_n N_A_1062_93#_c_766_n 0.0224887f $X=4.745 $Y=1.155
+ $X2=0 $Y2=0
cc_587 N_A_520_87#_c_663_n N_A_1062_93#_c_766_n 4.1682e-19 $X=4.935 $Y=1.42
+ $X2=0 $Y2=0
cc_588 N_A_520_87#_c_664_n N_A_1062_93#_c_766_n 2.64981e-19 $X=4.935 $Y=1.255
+ $X2=0 $Y2=0
cc_589 N_A_520_87#_c_660_n N_A_1062_93#_c_769_n 0.00115066f $X=4.745 $Y=1.155
+ $X2=0 $Y2=0
cc_590 N_A_520_87#_c_663_n N_A_1062_93#_c_769_n 0.020758f $X=4.935 $Y=1.42 $X2=0
+ $Y2=0
cc_591 N_A_520_87#_c_660_n N_A_1062_93#_c_770_n 7.50369e-19 $X=4.745 $Y=1.155
+ $X2=0 $Y2=0
cc_592 N_A_520_87#_c_664_n N_A_1062_93#_c_770_n 0.0175976f $X=4.935 $Y=1.255
+ $X2=0 $Y2=0
cc_593 N_A_520_87#_c_656_n N_A_27_74#_M1004_g 0.00653675f $X=3.125 $Y=0.58 $X2=0
+ $Y2=0
cc_594 N_A_520_87#_c_666_n N_A_27_74#_M1039_g 0.0134394f $X=3.265 $Y=2.17 $X2=0
+ $Y2=0
cc_595 N_A_520_87#_c_658_n N_A_27_74#_M1039_g 0.0084238f $X=3.89 $Y=1.71 $X2=0
+ $Y2=0
cc_596 N_A_520_87#_c_662_n N_A_27_74#_M1039_g 6.59953e-19 $X=3.277 $Y=1.71 $X2=0
+ $Y2=0
cc_597 N_A_520_87#_M1035_g N_A_27_74#_c_929_n 0.0105864f $X=5.01 $Y=2.315 $X2=0
+ $Y2=0
cc_598 N_A_520_87#_c_656_n N_A_214_74#_c_1121_n 4.50715e-19 $X=3.125 $Y=0.58
+ $X2=0 $Y2=0
cc_599 N_A_520_87#_c_656_n N_A_214_74#_M1025_g 0.0157186f $X=3.125 $Y=0.58 $X2=0
+ $Y2=0
cc_600 N_A_520_87#_c_657_n N_A_214_74#_M1025_g 0.00629505f $X=3.21 $Y=1.625
+ $X2=0 $Y2=0
cc_601 N_A_520_87#_c_666_n N_A_214_74#_M1016_g 0.0044257f $X=3.265 $Y=2.17 $X2=0
+ $Y2=0
cc_602 N_A_520_87#_c_662_n N_A_214_74#_M1016_g 0.0035635f $X=3.277 $Y=1.71 $X2=0
+ $Y2=0
cc_603 N_A_520_87#_c_656_n N_A_214_74#_c_1124_n 0.00397316f $X=3.125 $Y=0.58
+ $X2=0 $Y2=0
cc_604 N_A_520_87#_c_664_n N_A_214_74#_c_1124_n 0.00882199f $X=4.935 $Y=1.255
+ $X2=0 $Y2=0
cc_605 N_A_520_87#_c_657_n N_A_214_74#_c_1127_n 0.00550783f $X=3.21 $Y=1.625
+ $X2=0 $Y2=0
cc_606 N_A_520_87#_c_666_n N_VPWR_c_1652_n 0.0110142f $X=3.265 $Y=2.17 $X2=0
+ $Y2=0
cc_607 N_A_520_87#_c_658_n N_VPWR_c_1652_n 0.00811661f $X=3.89 $Y=1.71 $X2=0
+ $Y2=0
cc_608 N_A_520_87#_c_656_n N_A_422_125#_c_1795_n 0.00863643f $X=3.125 $Y=0.58
+ $X2=0 $Y2=0
cc_609 N_A_520_87#_c_656_n N_A_422_125#_c_1796_n 0.0257208f $X=3.125 $Y=0.58
+ $X2=0 $Y2=0
cc_610 N_A_520_87#_c_657_n N_A_422_125#_c_1796_n 0.0134534f $X=3.21 $Y=1.625
+ $X2=0 $Y2=0
cc_611 N_A_520_87#_c_657_n N_A_422_125#_c_1798_n 0.0384791f $X=3.21 $Y=1.625
+ $X2=0 $Y2=0
cc_612 N_A_520_87#_c_666_n N_A_422_125#_c_1798_n 0.0405723f $X=3.265 $Y=2.17
+ $X2=0 $Y2=0
cc_613 N_A_520_87#_c_662_n N_A_422_125#_c_1798_n 0.0137143f $X=3.277 $Y=1.71
+ $X2=0 $Y2=0
cc_614 N_A_520_87#_c_660_n N_VGND_M1036_d 9.80362e-19 $X=4.745 $Y=1.155 $X2=0
+ $Y2=0
cc_615 N_A_520_87#_c_661_n N_VGND_M1036_d 0.00132245f $X=4.06 $Y=1.155 $X2=0
+ $Y2=0
cc_616 N_A_520_87#_c_656_n N_VGND_c_1904_n 0.00540135f $X=3.125 $Y=0.58 $X2=0
+ $Y2=0
cc_617 N_A_520_87#_c_656_n N_VGND_c_1915_n 0.0338125f $X=3.125 $Y=0.58 $X2=0
+ $Y2=0
cc_618 N_A_520_87#_c_656_n N_VGND_c_1919_n 0.0230527f $X=3.125 $Y=0.58 $X2=0
+ $Y2=0
cc_619 N_A_520_87#_c_656_n A_606_87# 0.00465801f $X=3.125 $Y=0.58 $X2=-0.19
+ $Y2=-0.245
cc_620 N_A_520_87#_c_657_n A_606_87# 0.00637288f $X=3.21 $Y=1.625 $X2=-0.19
+ $Y2=-0.245
cc_621 N_A_520_87#_c_660_n N_A_872_119#_M1033_d 0.00457168f $X=4.745 $Y=1.155
+ $X2=-0.19 $Y2=-0.245
cc_622 N_A_520_87#_c_664_n N_A_872_119#_c_2063_n 0.00141486f $X=4.935 $Y=1.255
+ $X2=0 $Y2=0
cc_623 N_A_520_87#_c_664_n N_A_872_119#_c_2064_n 0.00295816f $X=4.935 $Y=1.255
+ $X2=0 $Y2=0
cc_624 N_A_1062_93#_M1011_g N_A_27_74#_c_929_n 0.0124167f $X=5.43 $Y=2.315 $X2=0
+ $Y2=0
cc_625 N_A_1062_93#_c_764_n N_A_27_74#_c_916_n 0.0195501f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_626 N_A_1062_93#_c_764_n N_A_27_74#_c_917_n 0.00369898f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_627 N_A_1062_93#_c_764_n N_A_27_74#_c_919_n 0.0060273f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_628 N_A_1062_93#_c_764_n N_A_27_74#_c_920_n 3.41598e-19 $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_629 N_A_1062_93#_c_764_n N_A_27_74#_c_921_n 0.0203746f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_630 N_A_1062_93#_c_770_n N_A_214_74#_c_1124_n 0.00882199f $X=5.475 $Y=1.255
+ $X2=0 $Y2=0
cc_631 N_A_1062_93#_c_764_n N_A_214_74#_c_1128_n 0.0114635f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_632 N_A_1062_93#_c_764_n N_A_1474_446#_M1021_g 0.00322586f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_633 N_A_1062_93#_c_777_n N_A_1474_446#_M1008_g 2.23317e-19 $X=10.24 $Y=1.985
+ $X2=0 $Y2=0
cc_634 N_A_1062_93#_M1024_g N_A_1474_446#_c_1278_n 0.00195126f $X=9.41 $Y=2.46
+ $X2=0 $Y2=0
cc_635 N_A_1062_93#_M1024_g N_A_1474_446#_c_1267_n 0.0138367f $X=9.41 $Y=2.46
+ $X2=0 $Y2=0
cc_636 N_A_1062_93#_c_759_n N_A_1474_446#_c_1267_n 0.00671177f $X=9.4 $Y=1.22
+ $X2=0 $Y2=0
cc_637 N_A_1062_93#_c_761_n N_A_1474_446#_c_1267_n 0.00374461f $X=9.41 $Y=1.295
+ $X2=0 $Y2=0
cc_638 N_A_1062_93#_c_776_n N_A_1474_446#_c_1267_n 0.00747985f $X=10.065
+ $Y=1.945 $X2=0 $Y2=0
cc_639 N_A_1062_93#_c_764_n N_A_1474_446#_c_1267_n 0.0121037f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_640 N_A_1062_93#_c_767_n N_A_1474_446#_c_1267_n 0.00228603f $X=9.84 $Y=1.295
+ $X2=0 $Y2=0
cc_641 N_A_1062_93#_c_768_n N_A_1474_446#_c_1267_n 0.0252649f $X=9.84 $Y=1.295
+ $X2=0 $Y2=0
cc_642 N_A_1062_93#_c_771_n N_A_1474_446#_c_1267_n 4.9787e-19 $X=9.875 $Y=1.295
+ $X2=0 $Y2=0
cc_643 N_A_1062_93#_c_772_n N_A_1474_446#_c_1267_n 0.00518815f $X=9.887 $Y=1.19
+ $X2=0 $Y2=0
cc_644 N_A_1062_93#_M1000_s N_A_1474_446#_c_1280_n 0.0105889f $X=10.115 $Y=1.84
+ $X2=0 $Y2=0
cc_645 N_A_1062_93#_M1024_g N_A_1474_446#_c_1280_n 0.0150681f $X=9.41 $Y=2.46
+ $X2=0 $Y2=0
cc_646 N_A_1062_93#_c_776_n N_A_1474_446#_c_1280_n 0.0297197f $X=10.065 $Y=1.945
+ $X2=0 $Y2=0
cc_647 N_A_1062_93#_c_777_n N_A_1474_446#_c_1280_n 0.0210811f $X=10.24 $Y=1.985
+ $X2=0 $Y2=0
cc_648 N_A_1062_93#_c_771_n N_A_1474_446#_c_1280_n 8.3656e-19 $X=9.875 $Y=1.295
+ $X2=0 $Y2=0
cc_649 N_A_1062_93#_c_777_n N_A_1474_446#_c_1281_n 0.0106031f $X=10.24 $Y=1.985
+ $X2=0 $Y2=0
cc_650 N_A_1062_93#_M1024_g N_A_1474_446#_c_1302_n 0.0192274f $X=9.41 $Y=2.46
+ $X2=0 $Y2=0
cc_651 N_A_1062_93#_c_776_n N_A_1474_446#_c_1302_n 0.00526144f $X=10.065
+ $Y=1.945 $X2=0 $Y2=0
cc_652 N_A_1062_93#_c_764_n N_A_1474_446#_c_1302_n 0.00906167f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_653 N_A_1062_93#_c_759_n N_A_1474_446#_c_1324_n 0.00573501f $X=9.4 $Y=1.22
+ $X2=0 $Y2=0
cc_654 N_A_1062_93#_c_764_n N_A_1474_446#_c_1324_n 0.00638392f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_655 N_A_1062_93#_M1024_g N_A_1314_424#_M1010_g 0.0826966f $X=9.41 $Y=2.46
+ $X2=0 $Y2=0
cc_656 N_A_1062_93#_c_764_n N_A_1314_424#_c_1439_n 0.0340295f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_657 N_A_1062_93#_c_764_n N_A_1314_424#_c_1441_n 0.0302998f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_658 N_A_1062_93#_c_759_n N_A_1314_424#_c_1442_n 2.35854e-19 $X=9.4 $Y=1.22
+ $X2=0 $Y2=0
cc_659 N_A_1062_93#_c_761_n N_A_1314_424#_c_1442_n 3.7036e-19 $X=9.41 $Y=1.295
+ $X2=0 $Y2=0
cc_660 N_A_1062_93#_c_764_n N_A_1314_424#_c_1442_n 0.046608f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_661 N_A_1062_93#_c_764_n N_A_1314_424#_c_1444_n 0.0183069f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_662 N_A_1062_93#_c_761_n N_A_1314_424#_c_1445_n 0.021255f $X=9.41 $Y=1.295
+ $X2=0 $Y2=0
cc_663 N_A_1062_93#_c_764_n N_A_1314_424#_c_1445_n 0.00365831f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_664 N_A_1062_93#_c_759_n N_A_1314_424#_c_1446_n 0.0247919f $X=9.4 $Y=1.22
+ $X2=0 $Y2=0
cc_665 N_A_1062_93#_c_763_n N_RESET_B_M1007_g 0.00698007f $X=10.22 $Y=0.58 $X2=0
+ $Y2=0
cc_666 N_A_1062_93#_c_772_n N_RESET_B_M1007_g 0.00507751f $X=9.887 $Y=1.19 $X2=0
+ $Y2=0
cc_667 N_A_1062_93#_c_762_n N_RESET_B_M1000_g 0.00555304f $X=9.875 $Y=1.385
+ $X2=0 $Y2=0
cc_668 N_A_1062_93#_c_777_n N_RESET_B_M1000_g 0.00520656f $X=10.24 $Y=1.985
+ $X2=0 $Y2=0
cc_669 N_A_1062_93#_c_768_n N_RESET_B_c_1544_n 0.00112633f $X=9.84 $Y=1.295
+ $X2=0 $Y2=0
cc_670 N_A_1062_93#_c_771_n N_RESET_B_c_1544_n 0.0214207f $X=9.875 $Y=1.295
+ $X2=0 $Y2=0
cc_671 N_A_1062_93#_c_762_n N_RESET_B_c_1545_n 0.00112633f $X=9.875 $Y=1.385
+ $X2=0 $Y2=0
cc_672 N_A_1062_93#_c_777_n N_RESET_B_c_1545_n 0.00327725f $X=10.24 $Y=1.985
+ $X2=0 $Y2=0
cc_673 N_A_1062_93#_c_763_n N_RESET_B_c_1546_n 0.0029184f $X=10.22 $Y=0.58 $X2=0
+ $Y2=0
cc_674 N_A_1062_93#_c_772_n N_RESET_B_c_1546_n 0.00112633f $X=9.887 $Y=1.19
+ $X2=0 $Y2=0
cc_675 N_A_1062_93#_c_777_n N_RESET_B_c_1547_n 0.0138414f $X=10.24 $Y=1.985
+ $X2=0 $Y2=0
cc_676 N_A_1062_93#_c_763_n N_RESET_B_c_1547_n 0.0127967f $X=10.22 $Y=0.58 $X2=0
+ $Y2=0
cc_677 N_A_1062_93#_c_767_n N_RESET_B_c_1547_n 0.00145843f $X=9.84 $Y=1.295
+ $X2=0 $Y2=0
cc_678 N_A_1062_93#_c_771_n N_RESET_B_c_1547_n 0.00103133f $X=9.875 $Y=1.295
+ $X2=0 $Y2=0
cc_679 N_A_1062_93#_c_772_n N_RESET_B_c_1547_n 0.0538379f $X=9.887 $Y=1.19 $X2=0
+ $Y2=0
cc_680 N_A_1062_93#_c_776_n N_VPWR_M1024_d 0.00245171f $X=10.065 $Y=1.945 $X2=0
+ $Y2=0
cc_681 N_A_1062_93#_M1011_g N_VPWR_c_1653_n 0.00592421f $X=5.43 $Y=2.315 $X2=0
+ $Y2=0
cc_682 N_A_1062_93#_M1024_g N_VPWR_c_1654_n 0.0131496f $X=9.41 $Y=2.46 $X2=0
+ $Y2=0
cc_683 N_A_1062_93#_M1024_g N_VPWR_c_1657_n 0.00460063f $X=9.41 $Y=2.46 $X2=0
+ $Y2=0
cc_684 N_A_1062_93#_M1011_g N_VPWR_c_1649_n 0.00100812f $X=5.43 $Y=2.315 $X2=0
+ $Y2=0
cc_685 N_A_1062_93#_M1024_g N_VPWR_c_1649_n 0.0090832f $X=9.41 $Y=2.46 $X2=0
+ $Y2=0
cc_686 N_A_1062_93#_c_764_n N_VGND_c_1935_n 0.0120438f $X=9.695 $Y=1.295 $X2=0
+ $Y2=0
cc_687 N_A_1062_93#_c_764_n N_VGND_c_1906_n 0.00223229f $X=9.695 $Y=1.295 $X2=0
+ $Y2=0
cc_688 N_A_1062_93#_c_763_n N_VGND_c_1907_n 0.0189715f $X=10.22 $Y=0.58 $X2=0
+ $Y2=0
cc_689 N_A_1062_93#_c_764_n N_VGND_c_1911_n 0.00249368f $X=9.695 $Y=1.295 $X2=0
+ $Y2=0
cc_690 N_A_1062_93#_c_759_n N_VGND_c_1917_n 0.00278271f $X=9.4 $Y=1.22 $X2=0
+ $Y2=0
cc_691 N_A_1062_93#_c_763_n N_VGND_c_1917_n 0.0210954f $X=10.22 $Y=0.58 $X2=0
+ $Y2=0
cc_692 N_A_1062_93#_c_759_n N_VGND_c_1919_n 0.00358571f $X=9.4 $Y=1.22 $X2=0
+ $Y2=0
cc_693 N_A_1062_93#_c_763_n N_VGND_c_1919_n 0.0177302f $X=10.22 $Y=0.58 $X2=0
+ $Y2=0
cc_694 N_A_1062_93#_c_770_n N_A_872_119#_c_2063_n 0.00157384f $X=5.475 $Y=1.255
+ $X2=0 $Y2=0
cc_695 N_A_1062_93#_c_770_n N_A_872_119#_c_2065_n 0.00691858f $X=5.475 $Y=1.255
+ $X2=0 $Y2=0
cc_696 N_A_1062_93#_c_759_n N_A_1708_74#_c_2096_n 4.90836e-19 $X=9.4 $Y=1.22
+ $X2=0 $Y2=0
cc_697 N_A_1062_93#_c_764_n N_A_1708_74#_c_2096_n 0.00223048f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_698 N_A_1062_93#_c_759_n N_A_1708_74#_c_2093_n 0.0120308f $X=9.4 $Y=1.22
+ $X2=0 $Y2=0
cc_699 N_A_1062_93#_c_763_n N_A_1708_74#_c_2093_n 0.00666958f $X=10.22 $Y=0.58
+ $X2=0 $Y2=0
cc_700 N_A_1062_93#_c_760_n N_A_1708_74#_c_2100_n 0.00610556f $X=9.71 $Y=1.295
+ $X2=0 $Y2=0
cc_701 N_A_1062_93#_c_763_n N_A_1708_74#_c_2100_n 0.0310232f $X=10.22 $Y=0.58
+ $X2=0 $Y2=0
cc_702 N_A_1062_93#_c_764_n N_A_1708_74#_c_2100_n 0.0065442f $X=9.695 $Y=1.295
+ $X2=0 $Y2=0
cc_703 N_A_1062_93#_c_767_n N_A_1708_74#_c_2100_n 0.00126143f $X=9.84 $Y=1.295
+ $X2=0 $Y2=0
cc_704 N_A_1062_93#_c_768_n N_A_1708_74#_c_2100_n 9.59633e-19 $X=9.84 $Y=1.295
+ $X2=0 $Y2=0
cc_705 N_A_1062_93#_c_772_n N_A_1708_74#_c_2100_n 0.0155328f $X=9.887 $Y=1.19
+ $X2=0 $Y2=0
cc_706 N_A_27_74#_M1004_g N_A_214_74#_M1025_g 0.01308f $X=2.525 $Y=0.645 $X2=0
+ $Y2=0
cc_707 N_A_27_74#_c_926_n N_A_214_74#_M1016_g 0.0121418f $X=3.4 $Y=3.15 $X2=0
+ $Y2=0
cc_708 N_A_27_74#_M1039_g N_A_214_74#_M1016_g 0.0326246f $X=3.49 $Y=2.105 $X2=0
+ $Y2=0
cc_709 N_A_27_74#_c_915_n N_A_214_74#_c_1124_n 0.00410612f $X=6.77 $Y=0.34 $X2=0
+ $Y2=0
cc_710 N_A_27_74#_c_923_n N_A_214_74#_c_1124_n 0.0105927f $X=7.505 $Y=0.9 $X2=0
+ $Y2=0
cc_711 N_A_27_74#_c_906_n N_A_214_74#_c_1125_n 0.01308f $X=2.45 $Y=0.18 $X2=0
+ $Y2=0
cc_712 N_A_27_74#_c_914_n N_A_214_74#_M1012_g 0.0156389f $X=7.345 $Y=0.34 $X2=0
+ $Y2=0
cc_713 N_A_27_74#_c_916_n N_A_214_74#_M1012_g 9.92945e-19 $X=7.505 $Y=1.065
+ $X2=0 $Y2=0
cc_714 N_A_27_74#_c_917_n N_A_214_74#_M1012_g 0.0105927f $X=7.505 $Y=1.065 $X2=0
+ $Y2=0
cc_715 N_A_27_74#_c_921_n N_A_214_74#_M1012_g 0.00586547f $X=6.605 $Y=1.61 $X2=0
+ $Y2=0
cc_716 N_A_27_74#_c_929_n N_A_214_74#_M1001_g 0.00926378f $X=6.39 $Y=3.15 $X2=0
+ $Y2=0
cc_717 N_A_27_74#_c_917_n N_A_214_74#_c_1128_n 6.51839e-19 $X=7.505 $Y=1.065
+ $X2=0 $Y2=0
cc_718 N_A_27_74#_M1005_g N_A_214_74#_c_1129_n 0.00534854f $X=6.48 $Y=2.54 $X2=0
+ $Y2=0
cc_719 N_A_27_74#_c_919_n N_A_214_74#_c_1129_n 3.84827e-19 $X=6.605 $Y=1.775
+ $X2=0 $Y2=0
cc_720 N_A_27_74#_c_920_n N_A_214_74#_c_1129_n 0.0207569f $X=6.605 $Y=1.775
+ $X2=0 $Y2=0
cc_721 N_A_27_74#_c_921_n N_A_214_74#_c_1129_n 0.00155147f $X=6.605 $Y=1.61
+ $X2=0 $Y2=0
cc_722 N_A_27_74#_M1005_g N_A_214_74#_c_1138_n 0.00926378f $X=6.48 $Y=2.54 $X2=0
+ $Y2=0
cc_723 N_A_27_74#_M1017_g N_A_214_74#_c_1130_n 5.04179e-19 $X=0.995 $Y=0.74
+ $X2=0 $Y2=0
cc_724 N_A_27_74#_c_905_n N_A_214_74#_c_1130_n 0.0148152f $X=1.525 $Y=1.3 $X2=0
+ $Y2=0
cc_725 N_A_27_74#_M1017_g N_A_214_74#_c_1131_n 0.00269942f $X=0.995 $Y=0.74
+ $X2=0 $Y2=0
cc_726 N_A_27_74#_c_904_n N_A_214_74#_c_1131_n 0.00748749f $X=1.45 $Y=1.375
+ $X2=0 $Y2=0
cc_727 N_A_27_74#_c_905_n N_A_214_74#_c_1131_n 0.0134812f $X=1.525 $Y=1.3 $X2=0
+ $Y2=0
cc_728 N_A_27_74#_c_910_n N_A_214_74#_c_1131_n 0.00313259f $X=1.675 $Y=1.375
+ $X2=0 $Y2=0
cc_729 N_A_27_74#_c_913_n N_A_214_74#_c_1131_n 0.023994f $X=1.06 $Y=1.465 $X2=0
+ $Y2=0
cc_730 N_A_27_74#_c_922_n N_A_214_74#_c_1131_n 0.00882834f $X=1.265 $Y=1.465
+ $X2=0 $Y2=0
cc_731 N_A_27_74#_c_908_n N_A_214_74#_c_1132_n 0.0229188f $X=1.675 $Y=3.075
+ $X2=0 $Y2=0
cc_732 N_A_27_74#_c_934_n N_A_214_74#_c_1132_n 0.0119282f $X=0.975 $Y=1.805
+ $X2=0 $Y2=0
cc_733 N_A_27_74#_c_913_n N_A_214_74#_c_1132_n 0.00985303f $X=1.06 $Y=1.465
+ $X2=0 $Y2=0
cc_734 N_A_27_74#_c_922_n N_A_214_74#_c_1132_n 0.00258611f $X=1.265 $Y=1.465
+ $X2=0 $Y2=0
cc_735 N_A_27_74#_c_905_n N_A_214_74#_c_1133_n 0.00237249f $X=1.525 $Y=1.3 $X2=0
+ $Y2=0
cc_736 N_A_27_74#_c_908_n N_A_214_74#_c_1133_n 0.0117473f $X=1.675 $Y=3.075
+ $X2=0 $Y2=0
cc_737 N_A_27_74#_c_910_n N_A_214_74#_c_1133_n 0.00620701f $X=1.675 $Y=1.375
+ $X2=0 $Y2=0
cc_738 N_A_27_74#_M1004_g N_A_214_74#_c_1134_n 0.00680601f $X=2.525 $Y=0.645
+ $X2=0 $Y2=0
cc_739 N_A_27_74#_c_914_n N_A_1474_446#_M1021_g 0.00176953f $X=7.345 $Y=0.34
+ $X2=0 $Y2=0
cc_740 N_A_27_74#_c_916_n N_A_1474_446#_M1021_g 0.00609261f $X=7.505 $Y=1.065
+ $X2=0 $Y2=0
cc_741 N_A_27_74#_c_917_n N_A_1474_446#_M1021_g 0.0203391f $X=7.505 $Y=1.065
+ $X2=0 $Y2=0
cc_742 N_A_27_74#_c_923_n N_A_1474_446#_M1021_g 0.0170701f $X=7.505 $Y=0.9 $X2=0
+ $Y2=0
cc_743 N_A_27_74#_c_914_n N_A_1314_424#_M1012_d 0.00514156f $X=7.345 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_744 N_A_27_74#_M1005_g N_A_1314_424#_c_1448_n 0.00730563f $X=6.48 $Y=2.54
+ $X2=0 $Y2=0
cc_745 N_A_27_74#_c_914_n N_A_1314_424#_c_1439_n 0.0155805f $X=7.345 $Y=0.34
+ $X2=0 $Y2=0
cc_746 N_A_27_74#_c_916_n N_A_1314_424#_c_1439_n 0.0480163f $X=7.505 $Y=1.065
+ $X2=0 $Y2=0
cc_747 N_A_27_74#_c_921_n N_A_1314_424#_c_1439_n 0.037512f $X=6.605 $Y=1.61
+ $X2=0 $Y2=0
cc_748 N_A_27_74#_c_923_n N_A_1314_424#_c_1439_n 0.00463634f $X=7.505 $Y=0.9
+ $X2=0 $Y2=0
cc_749 N_A_27_74#_M1005_g N_A_1314_424#_c_1440_n 0.00295298f $X=6.48 $Y=2.54
+ $X2=0 $Y2=0
cc_750 N_A_27_74#_c_920_n N_A_1314_424#_c_1440_n 0.0017734f $X=6.605 $Y=1.775
+ $X2=0 $Y2=0
cc_751 N_A_27_74#_c_921_n N_A_1314_424#_c_1440_n 0.0277379f $X=6.605 $Y=1.61
+ $X2=0 $Y2=0
cc_752 N_A_27_74#_c_916_n N_A_1314_424#_c_1441_n 0.0201659f $X=7.505 $Y=1.065
+ $X2=0 $Y2=0
cc_753 N_A_27_74#_c_917_n N_A_1314_424#_c_1441_n 0.00246536f $X=7.505 $Y=1.065
+ $X2=0 $Y2=0
cc_754 N_A_27_74#_M1005_g N_A_1314_424#_c_1450_n 0.00349838f $X=6.48 $Y=2.54
+ $X2=0 $Y2=0
cc_755 N_A_27_74#_c_919_n N_A_1314_424#_c_1450_n 0.0179252f $X=6.605 $Y=1.775
+ $X2=0 $Y2=0
cc_756 N_A_27_74#_c_920_n N_A_1314_424#_c_1450_n 0.00140285f $X=6.605 $Y=1.775
+ $X2=0 $Y2=0
cc_757 N_A_27_74#_c_921_n N_A_1314_424#_c_1443_n 0.0143562f $X=6.605 $Y=1.61
+ $X2=0 $Y2=0
cc_758 N_A_27_74#_c_916_n N_A_1314_424#_c_1444_n 0.00555387f $X=7.505 $Y=1.065
+ $X2=0 $Y2=0
cc_759 N_A_27_74#_c_917_n N_A_1314_424#_c_1444_n 3.38303e-19 $X=7.505 $Y=1.065
+ $X2=0 $Y2=0
cc_760 N_A_27_74#_c_934_n N_VPWR_M1018_d 0.00314765f $X=0.975 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_761 N_A_27_74#_M1028_g N_VPWR_c_1650_n 0.00880174f $X=1.175 $Y=2.4 $X2=0
+ $Y2=0
cc_762 N_A_27_74#_c_908_n N_VPWR_c_1650_n 0.00231241f $X=1.675 $Y=3.075 $X2=0
+ $Y2=0
cc_763 N_A_27_74#_c_933_n N_VPWR_c_1650_n 0.0369884f $X=0.37 $Y=1.985 $X2=0
+ $Y2=0
cc_764 N_A_27_74#_c_934_n N_VPWR_c_1650_n 0.0236498f $X=0.975 $Y=1.805 $X2=0
+ $Y2=0
cc_765 N_A_27_74#_c_922_n N_VPWR_c_1650_n 4.14145e-19 $X=1.265 $Y=1.465 $X2=0
+ $Y2=0
cc_766 N_A_27_74#_c_908_n N_VPWR_c_1651_n 0.0131353f $X=1.675 $Y=3.075 $X2=0
+ $Y2=0
cc_767 N_A_27_74#_c_926_n N_VPWR_c_1651_n 0.03981f $X=3.4 $Y=3.15 $X2=0 $Y2=0
cc_768 N_A_27_74#_M1039_g N_VPWR_c_1652_n 0.0203571f $X=3.49 $Y=2.105 $X2=0
+ $Y2=0
cc_769 N_A_27_74#_c_929_n N_VPWR_c_1652_n 0.0215035f $X=6.39 $Y=3.15 $X2=0 $Y2=0
cc_770 N_A_27_74#_c_929_n N_VPWR_c_1653_n 0.0275116f $X=6.39 $Y=3.15 $X2=0 $Y2=0
cc_771 N_A_27_74#_M1005_g N_VPWR_c_1653_n 6.745e-19 $X=6.48 $Y=2.54 $X2=0 $Y2=0
cc_772 N_A_27_74#_M1028_g N_VPWR_c_1659_n 0.00553757f $X=1.175 $Y=2.4 $X2=0
+ $Y2=0
cc_773 N_A_27_74#_c_927_n N_VPWR_c_1659_n 0.00796123f $X=1.75 $Y=3.15 $X2=0
+ $Y2=0
cc_774 N_A_27_74#_c_926_n N_VPWR_c_1660_n 0.0510543f $X=3.4 $Y=3.15 $X2=0 $Y2=0
cc_775 N_A_27_74#_c_929_n N_VPWR_c_1661_n 0.0314889f $X=6.39 $Y=3.15 $X2=0 $Y2=0
cc_776 N_A_27_74#_M1028_g N_VPWR_c_1649_n 0.010905f $X=1.175 $Y=2.4 $X2=0 $Y2=0
cc_777 N_A_27_74#_c_926_n N_VPWR_c_1649_n 0.0413038f $X=3.4 $Y=3.15 $X2=0 $Y2=0
cc_778 N_A_27_74#_c_927_n N_VPWR_c_1649_n 0.0114361f $X=1.75 $Y=3.15 $X2=0 $Y2=0
cc_779 N_A_27_74#_c_929_n N_VPWR_c_1649_n 0.07478f $X=6.39 $Y=3.15 $X2=0 $Y2=0
cc_780 N_A_27_74#_c_931_n N_VPWR_c_1649_n 0.0111208f $X=3.49 $Y=3.15 $X2=0 $Y2=0
cc_781 N_A_27_74#_c_933_n N_VPWR_c_1649_n 0.0164063f $X=0.37 $Y=1.985 $X2=0
+ $Y2=0
cc_782 N_A_27_74#_c_933_n N_VPWR_c_1666_n 0.0199035f $X=0.37 $Y=1.985 $X2=0
+ $Y2=0
cc_783 N_A_27_74#_c_929_n N_VPWR_c_1670_n 0.0176354f $X=6.39 $Y=3.15 $X2=0 $Y2=0
cc_784 N_A_27_74#_c_906_n N_A_422_125#_c_1795_n 0.00440091f $X=2.45 $Y=0.18
+ $X2=0 $Y2=0
cc_785 N_A_27_74#_M1004_g N_A_422_125#_c_1795_n 0.00529615f $X=2.525 $Y=0.645
+ $X2=0 $Y2=0
cc_786 N_A_27_74#_c_906_n N_A_422_125#_c_1796_n 5.05855e-19 $X=2.45 $Y=0.18
+ $X2=0 $Y2=0
cc_787 N_A_27_74#_M1004_g N_A_422_125#_c_1796_n 0.00946624f $X=2.525 $Y=0.645
+ $X2=0 $Y2=0
cc_788 N_A_27_74#_c_926_n N_A_422_125#_c_1799_n 0.00567784f $X=3.4 $Y=3.15 $X2=0
+ $Y2=0
cc_789 N_A_27_74#_M1039_g N_A_422_125#_c_1799_n 0.00210566f $X=3.49 $Y=2.105
+ $X2=0 $Y2=0
cc_790 N_A_27_74#_M1039_g N_A_422_125#_c_1798_n 2.60695e-19 $X=3.49 $Y=2.105
+ $X2=0 $Y2=0
cc_791 N_A_27_74#_M1017_g N_VGND_c_1902_n 0.0125459f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_792 N_A_27_74#_c_905_n N_VGND_c_1902_n 4.60892e-19 $X=1.525 $Y=1.3 $X2=0
+ $Y2=0
cc_793 N_A_27_74#_c_907_n N_VGND_c_1902_n 0.00286132f $X=1.6 $Y=0.18 $X2=0 $Y2=0
cc_794 N_A_27_74#_c_911_n N_VGND_c_1902_n 0.0258493f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_795 N_A_27_74#_M1017_g N_VGND_c_1903_n 0.00383152f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_796 N_A_27_74#_c_907_n N_VGND_c_1903_n 0.00748834f $X=1.6 $Y=0.18 $X2=0 $Y2=0
cc_797 N_A_27_74#_c_905_n N_VGND_c_1904_n 0.0117703f $X=1.525 $Y=1.3 $X2=0 $Y2=0
cc_798 N_A_27_74#_c_906_n N_VGND_c_1904_n 0.0200453f $X=2.45 $Y=0.18 $X2=0 $Y2=0
cc_799 N_A_27_74#_M1004_g N_VGND_c_1904_n 0.00534265f $X=2.525 $Y=0.645 $X2=0
+ $Y2=0
cc_800 N_A_27_74#_c_910_n N_VGND_c_1904_n 6.48816e-19 $X=1.675 $Y=1.375 $X2=0
+ $Y2=0
cc_801 N_A_27_74#_c_915_n N_VGND_c_1905_n 0.015162f $X=6.77 $Y=0.34 $X2=0 $Y2=0
cc_802 N_A_27_74#_c_921_n N_VGND_c_1905_n 0.0134343f $X=6.605 $Y=1.61 $X2=0
+ $Y2=0
cc_803 N_A_27_74#_c_914_n N_VGND_c_1906_n 0.00670281f $X=7.345 $Y=0.34 $X2=0
+ $Y2=0
cc_804 N_A_27_74#_c_916_n N_VGND_c_1906_n 0.0148625f $X=7.505 $Y=1.065 $X2=0
+ $Y2=0
cc_805 N_A_27_74#_c_911_n N_VGND_c_1914_n 0.0158845f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_806 N_A_27_74#_c_906_n N_VGND_c_1915_n 0.0223339f $X=2.45 $Y=0.18 $X2=0 $Y2=0
cc_807 N_A_27_74#_c_914_n N_VGND_c_1916_n 0.0593225f $X=7.345 $Y=0.34 $X2=0
+ $Y2=0
cc_808 N_A_27_74#_c_915_n N_VGND_c_1916_n 0.0115893f $X=6.77 $Y=0.34 $X2=0 $Y2=0
cc_809 N_A_27_74#_c_923_n N_VGND_c_1916_n 0.0027813f $X=7.505 $Y=0.9 $X2=0 $Y2=0
cc_810 N_A_27_74#_M1017_g N_VGND_c_1919_n 0.00758454f $X=0.995 $Y=0.74 $X2=0
+ $Y2=0
cc_811 N_A_27_74#_c_906_n N_VGND_c_1919_n 0.0328412f $X=2.45 $Y=0.18 $X2=0 $Y2=0
cc_812 N_A_27_74#_c_907_n N_VGND_c_1919_n 0.0101927f $X=1.6 $Y=0.18 $X2=0 $Y2=0
cc_813 N_A_27_74#_c_911_n N_VGND_c_1919_n 0.0130993f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_814 N_A_27_74#_c_914_n N_VGND_c_1919_n 0.0327286f $X=7.345 $Y=0.34 $X2=0
+ $Y2=0
cc_815 N_A_27_74#_c_915_n N_VGND_c_1919_n 0.00583135f $X=6.77 $Y=0.34 $X2=0
+ $Y2=0
cc_816 N_A_27_74#_c_923_n N_VGND_c_1919_n 0.00355475f $X=7.505 $Y=0.9 $X2=0
+ $Y2=0
cc_817 N_A_27_74#_c_921_n A_1318_119# 0.00287467f $X=6.605 $Y=1.61 $X2=-0.19
+ $Y2=-0.245
cc_818 N_A_27_74#_c_914_n A_1498_74# 7.09228e-19 $X=7.345 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_819 N_A_27_74#_c_916_n A_1498_74# 0.00458644f $X=7.505 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_820 N_A_214_74#_c_1129_n N_A_1474_446#_c_1276_n 0.00313657f $X=7.027 $Y=2.18
+ $X2=0 $Y2=0
cc_821 N_A_214_74#_M1001_g N_A_1474_446#_c_1277_n 0.0344219f $X=7.015 $Y=2.75
+ $X2=0 $Y2=0
cc_822 N_A_214_74#_c_1129_n N_A_1474_446#_c_1277_n 0.00315962f $X=7.027 $Y=2.18
+ $X2=0 $Y2=0
cc_823 N_A_214_74#_c_1138_n N_A_1474_446#_c_1277_n 0.00509396f $X=7.027 $Y=2.33
+ $X2=0 $Y2=0
cc_824 N_A_214_74#_c_1138_n N_A_1314_424#_c_1448_n 0.00426858f $X=7.027 $Y=2.33
+ $X2=0 $Y2=0
cc_825 N_A_214_74#_M1012_g N_A_1314_424#_c_1439_n 0.00871573f $X=6.875 $Y=0.87
+ $X2=0 $Y2=0
cc_826 N_A_214_74#_c_1128_n N_A_1314_424#_c_1439_n 0.0107525f $X=7.055 $Y=1.295
+ $X2=0 $Y2=0
cc_827 N_A_214_74#_c_1129_n N_A_1314_424#_c_1439_n 0.00122492f $X=7.027 $Y=2.18
+ $X2=0 $Y2=0
cc_828 N_A_214_74#_c_1129_n N_A_1314_424#_c_1440_n 0.0175654f $X=7.027 $Y=2.18
+ $X2=0 $Y2=0
cc_829 N_A_214_74#_c_1138_n N_A_1314_424#_c_1440_n 3.01272e-19 $X=7.027 $Y=2.33
+ $X2=0 $Y2=0
cc_830 N_A_214_74#_c_1129_n N_A_1314_424#_c_1450_n 0.0026461f $X=7.027 $Y=2.18
+ $X2=0 $Y2=0
cc_831 N_A_214_74#_c_1138_n N_A_1314_424#_c_1450_n 0.00957612f $X=7.027 $Y=2.33
+ $X2=0 $Y2=0
cc_832 N_A_214_74#_c_1129_n N_A_1314_424#_c_1443_n 0.0100462f $X=7.027 $Y=2.18
+ $X2=0 $Y2=0
cc_833 N_A_214_74#_c_1132_n N_VPWR_c_1650_n 0.00109322f $X=1.4 $Y=1.985 $X2=0
+ $Y2=0
cc_834 N_A_214_74#_c_1132_n N_VPWR_c_1651_n 0.037269f $X=1.4 $Y=1.985 $X2=0
+ $Y2=0
cc_835 N_A_214_74#_c_1132_n N_VPWR_c_1659_n 0.011066f $X=1.4 $Y=1.985 $X2=0
+ $Y2=0
cc_836 N_A_214_74#_M1016_g N_VPWR_c_1649_n 0.00112709f $X=2.97 $Y=2.525 $X2=0
+ $Y2=0
cc_837 N_A_214_74#_M1001_g N_VPWR_c_1649_n 0.00423612f $X=7.015 $Y=2.75 $X2=0
+ $Y2=0
cc_838 N_A_214_74#_c_1132_n N_VPWR_c_1649_n 0.00915947f $X=1.4 $Y=1.985 $X2=0
+ $Y2=0
cc_839 N_A_214_74#_M1001_g N_VPWR_c_1670_n 0.00333926f $X=7.015 $Y=2.75 $X2=0
+ $Y2=0
cc_840 N_A_214_74#_M1025_g N_A_422_125#_c_1796_n 0.00663728f $X=2.955 $Y=0.645
+ $X2=0 $Y2=0
cc_841 N_A_214_74#_c_1133_n N_A_422_125#_c_1796_n 0.0210062f $X=2.485 $Y=1.42
+ $X2=0 $Y2=0
cc_842 N_A_214_74#_c_1134_n N_A_422_125#_c_1796_n 0.00972455f $X=2.485 $Y=1.33
+ $X2=0 $Y2=0
cc_843 N_A_214_74#_c_1131_n N_A_422_125#_c_1797_n 5.65197e-19 $X=1.44 $Y=1.585
+ $X2=0 $Y2=0
cc_844 N_A_214_74#_c_1133_n N_A_422_125#_c_1797_n 0.0212522f $X=2.485 $Y=1.42
+ $X2=0 $Y2=0
cc_845 N_A_214_74#_c_1134_n N_A_422_125#_c_1797_n 3.45666e-19 $X=2.485 $Y=1.33
+ $X2=0 $Y2=0
cc_846 N_A_214_74#_M1016_g N_A_422_125#_c_1799_n 0.0123044f $X=2.97 $Y=2.525
+ $X2=0 $Y2=0
cc_847 N_A_214_74#_c_1121_n N_A_422_125#_c_1798_n 0.00746444f $X=2.88 $Y=1.33
+ $X2=0 $Y2=0
cc_848 N_A_214_74#_M1025_g N_A_422_125#_c_1798_n 0.00499504f $X=2.955 $Y=0.645
+ $X2=0 $Y2=0
cc_849 N_A_214_74#_M1016_g N_A_422_125#_c_1798_n 0.021377f $X=2.97 $Y=2.525
+ $X2=0 $Y2=0
cc_850 N_A_214_74#_c_1127_n N_A_422_125#_c_1798_n 0.00216139f $X=2.97 $Y=1.33
+ $X2=0 $Y2=0
cc_851 N_A_214_74#_c_1133_n N_A_422_125#_c_1798_n 0.0256544f $X=2.485 $Y=1.42
+ $X2=0 $Y2=0
cc_852 N_A_214_74#_c_1134_n N_A_422_125#_c_1798_n 0.00108296f $X=2.485 $Y=1.33
+ $X2=0 $Y2=0
cc_853 N_A_214_74#_c_1130_n N_VGND_c_1902_n 0.0222741f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_854 N_A_214_74#_c_1130_n N_VGND_c_1903_n 0.0158727f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_855 N_A_214_74#_c_1130_n N_VGND_c_1904_n 0.0467131f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_856 N_A_214_74#_c_1131_n N_VGND_c_1904_n 0.00900433f $X=1.44 $Y=1.585 $X2=0
+ $Y2=0
cc_857 N_A_214_74#_c_1133_n N_VGND_c_1904_n 0.0202767f $X=2.485 $Y=1.42 $X2=0
+ $Y2=0
cc_858 N_A_214_74#_c_1124_n N_VGND_c_1905_n 0.0279578f $X=6.8 $Y=0.18 $X2=0
+ $Y2=0
cc_859 N_A_214_74#_M1012_g N_VGND_c_1905_n 8.86009e-19 $X=6.875 $Y=0.87 $X2=0
+ $Y2=0
cc_860 N_A_214_74#_c_1124_n N_VGND_c_1909_n 0.0430985f $X=6.8 $Y=0.18 $X2=0
+ $Y2=0
cc_861 N_A_214_74#_M1025_g N_VGND_c_1915_n 0.00465262f $X=2.955 $Y=0.645 $X2=0
+ $Y2=0
cc_862 N_A_214_74#_c_1124_n N_VGND_c_1915_n 0.038842f $X=6.8 $Y=0.18 $X2=0 $Y2=0
cc_863 N_A_214_74#_c_1125_n N_VGND_c_1915_n 0.0185119f $X=3.03 $Y=0.18 $X2=0
+ $Y2=0
cc_864 N_A_214_74#_c_1124_n N_VGND_c_1916_n 0.0138999f $X=6.8 $Y=0.18 $X2=0
+ $Y2=0
cc_865 N_A_214_74#_c_1124_n N_VGND_c_1919_n 0.0798093f $X=6.8 $Y=0.18 $X2=0
+ $Y2=0
cc_866 N_A_214_74#_c_1125_n N_VGND_c_1919_n 0.00475067f $X=3.03 $Y=0.18 $X2=0
+ $Y2=0
cc_867 N_A_214_74#_c_1130_n N_VGND_c_1919_n 0.0130581f $X=1.21 $Y=0.515 $X2=0
+ $Y2=0
cc_868 N_A_214_74#_c_1124_n N_A_872_119#_c_2063_n 0.0110768f $X=6.8 $Y=0.18
+ $X2=0 $Y2=0
cc_869 N_A_214_74#_c_1124_n N_A_872_119#_c_2064_n 0.0097718f $X=6.8 $Y=0.18
+ $X2=0 $Y2=0
cc_870 N_A_214_74#_c_1124_n N_A_872_119#_c_2065_n 0.00794104f $X=6.8 $Y=0.18
+ $X2=0 $Y2=0
cc_871 N_A_1474_446#_c_1278_n N_A_1314_424#_M1010_g 0.0110058f $X=8.77 $Y=2.475
+ $X2=0 $Y2=0
cc_872 N_A_1474_446#_c_1267_n N_A_1314_424#_M1010_g 0.00628602f $X=9.3 $Y=1.97
+ $X2=0 $Y2=0
cc_873 N_A_1474_446#_c_1302_n N_A_1314_424#_M1010_g 0.0236248f $X=9.385 $Y=2.19
+ $X2=0 $Y2=0
cc_874 N_A_1474_446#_M1021_g N_A_1314_424#_c_1441_n 0.00542998f $X=7.955 $Y=0.58
+ $X2=0 $Y2=0
cc_875 N_A_1474_446#_c_1276_n N_A_1314_424#_c_1441_n 0.00207291f $X=7.955
+ $Y=1.81 $X2=0 $Y2=0
cc_876 N_A_1474_446#_c_1277_n N_A_1314_424#_c_1441_n 3.7868e-19 $X=7.785
+ $Y=2.215 $X2=0 $Y2=0
cc_877 N_A_1474_446#_M1021_g N_A_1314_424#_c_1442_n 4.92684e-19 $X=7.955 $Y=0.58
+ $X2=0 $Y2=0
cc_878 N_A_1474_446#_c_1267_n N_A_1314_424#_c_1442_n 0.0305515f $X=9.3 $Y=1.97
+ $X2=0 $Y2=0
cc_879 N_A_1474_446#_c_1302_n N_A_1314_424#_c_1442_n 0.00927806f $X=9.385
+ $Y=2.19 $X2=0 $Y2=0
cc_880 N_A_1474_446#_M1021_g N_A_1314_424#_c_1444_n 0.020561f $X=7.955 $Y=0.58
+ $X2=0 $Y2=0
cc_881 N_A_1474_446#_c_1267_n N_A_1314_424#_c_1445_n 0.00180678f $X=9.3 $Y=1.97
+ $X2=0 $Y2=0
cc_882 N_A_1474_446#_c_1302_n N_A_1314_424#_c_1445_n 5.85637e-19 $X=9.385
+ $Y=2.19 $X2=0 $Y2=0
cc_883 N_A_1474_446#_c_1324_n N_A_1314_424#_c_1445_n 7.03158e-19 $X=9.3 $Y=0.777
+ $X2=0 $Y2=0
cc_884 N_A_1474_446#_c_1267_n N_A_1314_424#_c_1446_n 0.00375181f $X=9.3 $Y=1.97
+ $X2=0 $Y2=0
cc_885 N_A_1474_446#_M1002_g N_RESET_B_M1007_g 0.0154694f $X=11.015 $Y=0.74
+ $X2=0 $Y2=0
cc_886 N_A_1474_446#_M1008_g N_RESET_B_M1000_g 0.0317942f $X=10.98 $Y=2.4 $X2=0
+ $Y2=0
cc_887 N_A_1474_446#_c_1280_n N_RESET_B_M1000_g 0.0206719f $X=10.78 $Y=2.325
+ $X2=0 $Y2=0
cc_888 N_A_1474_446#_c_1281_n N_RESET_B_M1000_g 0.00872838f $X=10.865 $Y=2.24
+ $X2=0 $Y2=0
cc_889 N_A_1474_446#_c_1268_n N_RESET_B_c_1544_n 0.00113328f $X=10.955 $Y=1.485
+ $X2=0 $Y2=0
cc_890 N_A_1474_446#_c_1269_n N_RESET_B_c_1544_n 0.0214892f $X=10.955 $Y=1.485
+ $X2=0 $Y2=0
cc_891 N_A_1474_446#_M1002_g N_RESET_B_c_1546_n 0.0102574f $X=11.015 $Y=0.74
+ $X2=0 $Y2=0
cc_892 N_A_1474_446#_M1002_g N_RESET_B_c_1547_n 0.00167795f $X=11.015 $Y=0.74
+ $X2=0 $Y2=0
cc_893 N_A_1474_446#_c_1280_n N_RESET_B_c_1547_n 0.00443777f $X=10.78 $Y=2.325
+ $X2=0 $Y2=0
cc_894 N_A_1474_446#_c_1268_n N_RESET_B_c_1547_n 0.0232735f $X=10.955 $Y=1.485
+ $X2=0 $Y2=0
cc_895 N_A_1474_446#_c_1269_n N_RESET_B_c_1547_n 4.00949e-19 $X=10.955 $Y=1.485
+ $X2=0 $Y2=0
cc_896 N_A_1474_446#_c_1275_n N_A_2320_410#_M1037_g 0.0184448f $X=11.95 $Y=1.975
+ $X2=0 $Y2=0
cc_897 N_A_1474_446#_c_1266_n N_A_2320_410#_M1037_g 0.00223102f $X=11.71
+ $Y=1.485 $X2=0 $Y2=0
cc_898 N_A_1474_446#_c_1262_n N_A_2320_410#_M1038_g 0.00198036f $X=11.71 $Y=1.32
+ $X2=0 $Y2=0
cc_899 N_A_1474_446#_c_1264_n N_A_2320_410#_M1038_g 0.0134505f $X=12.005
+ $Y=0.865 $X2=0 $Y2=0
cc_900 N_A_1474_446#_c_1262_n N_A_2320_410#_c_1590_n 0.018228f $X=11.71 $Y=1.32
+ $X2=0 $Y2=0
cc_901 N_A_1474_446#_c_1275_n N_A_2320_410#_c_1590_n 9.3041e-19 $X=11.95
+ $Y=1.975 $X2=0 $Y2=0
cc_902 N_A_1474_446#_c_1265_n N_A_2320_410#_c_1590_n 0.00329796f $X=12.005
+ $Y=0.94 $X2=0 $Y2=0
cc_903 N_A_1474_446#_M1002_g N_A_2320_410#_c_1592_n 0.00105741f $X=11.015
+ $Y=0.74 $X2=0 $Y2=0
cc_904 N_A_1474_446#_c_1262_n N_A_2320_410#_c_1592_n 0.00613665f $X=11.71
+ $Y=1.32 $X2=0 $Y2=0
cc_905 N_A_1474_446#_c_1264_n N_A_2320_410#_c_1592_n 0.00300625f $X=12.005
+ $Y=0.865 $X2=0 $Y2=0
cc_906 N_A_1474_446#_c_1265_n N_A_2320_410#_c_1592_n 0.0142998f $X=12.005
+ $Y=0.94 $X2=0 $Y2=0
cc_907 N_A_1474_446#_c_1275_n N_A_2320_410#_c_1597_n 0.00371718f $X=11.95
+ $Y=1.975 $X2=0 $Y2=0
cc_908 N_A_1474_446#_c_1275_n N_A_2320_410#_c_1598_n 0.0124878f $X=11.95
+ $Y=1.975 $X2=0 $Y2=0
cc_909 N_A_1474_446#_c_1275_n N_A_2320_410#_c_1593_n 0.00609223f $X=11.95
+ $Y=1.975 $X2=0 $Y2=0
cc_910 N_A_1474_446#_c_1265_n N_A_2320_410#_c_1593_n 0.0061315f $X=12.005
+ $Y=0.94 $X2=0 $Y2=0
cc_911 N_A_1474_446#_c_1262_n N_A_2320_410#_c_1594_n 0.00183591f $X=11.71
+ $Y=1.32 $X2=0 $Y2=0
cc_912 N_A_1474_446#_c_1275_n N_A_2320_410#_c_1594_n 0.00152885f $X=11.95
+ $Y=1.975 $X2=0 $Y2=0
cc_913 N_A_1474_446#_c_1266_n N_A_2320_410#_c_1594_n 0.0103185f $X=11.71
+ $Y=1.485 $X2=0 $Y2=0
cc_914 N_A_1474_446#_M1008_g N_A_2320_410#_c_1595_n 2.23836e-19 $X=10.98 $Y=2.4
+ $X2=0 $Y2=0
cc_915 N_A_1474_446#_c_1263_n N_A_2320_410#_c_1595_n 0.00397831f $X=11.71
+ $Y=1.825 $X2=0 $Y2=0
cc_916 N_A_1474_446#_c_1275_n N_A_2320_410#_c_1595_n 0.0111151f $X=11.95
+ $Y=1.975 $X2=0 $Y2=0
cc_917 N_A_1474_446#_c_1266_n N_A_2320_410#_c_1595_n 0.00234039f $X=11.71
+ $Y=1.485 $X2=0 $Y2=0
cc_918 N_A_1474_446#_c_1282_n N_VPWR_M1015_d 0.00564423f $X=8.685 $Y=2.19 $X2=0
+ $Y2=0
cc_919 N_A_1474_446#_c_1280_n N_VPWR_M1024_d 0.00982282f $X=10.78 $Y=2.325 $X2=0
+ $Y2=0
cc_920 N_A_1474_446#_c_1280_n N_VPWR_M1000_d 0.00872266f $X=10.78 $Y=2.325 $X2=0
+ $Y2=0
cc_921 N_A_1474_446#_c_1281_n N_VPWR_M1000_d 0.0047678f $X=10.865 $Y=2.24 $X2=0
+ $Y2=0
cc_922 N_A_1474_446#_c_1278_n N_VPWR_c_1654_n 0.011484f $X=8.77 $Y=2.475 $X2=0
+ $Y2=0
cc_923 N_A_1474_446#_c_1280_n N_VPWR_c_1654_n 0.0219568f $X=10.78 $Y=2.325 $X2=0
+ $Y2=0
cc_924 N_A_1474_446#_M1008_g N_VPWR_c_1655_n 0.0137845f $X=10.98 $Y=2.4 $X2=0
+ $Y2=0
cc_925 N_A_1474_446#_c_1280_n N_VPWR_c_1655_n 0.0217894f $X=10.78 $Y=2.325 $X2=0
+ $Y2=0
cc_926 N_A_1474_446#_c_1275_n N_VPWR_c_1656_n 0.00917765f $X=11.95 $Y=1.975
+ $X2=0 $Y2=0
cc_927 N_A_1474_446#_c_1278_n N_VPWR_c_1657_n 0.0108405f $X=8.77 $Y=2.475 $X2=0
+ $Y2=0
cc_928 N_A_1474_446#_M1008_g N_VPWR_c_1663_n 0.00460063f $X=10.98 $Y=2.4 $X2=0
+ $Y2=0
cc_929 N_A_1474_446#_c_1275_n N_VPWR_c_1663_n 0.00604985f $X=11.95 $Y=1.975
+ $X2=0 $Y2=0
cc_930 N_A_1474_446#_M1015_g N_VPWR_c_1649_n 0.00797798f $X=7.46 $Y=2.75 $X2=0
+ $Y2=0
cc_931 N_A_1474_446#_M1008_g N_VPWR_c_1649_n 0.00913687f $X=10.98 $Y=2.4 $X2=0
+ $Y2=0
cc_932 N_A_1474_446#_c_1275_n N_VPWR_c_1649_n 0.00628405f $X=11.95 $Y=1.975
+ $X2=0 $Y2=0
cc_933 N_A_1474_446#_c_1278_n N_VPWR_c_1649_n 0.00896536f $X=8.77 $Y=2.475 $X2=0
+ $Y2=0
cc_934 N_A_1474_446#_M1015_g N_VPWR_c_1670_n 0.00455976f $X=7.46 $Y=2.75 $X2=0
+ $Y2=0
cc_935 N_A_1474_446#_M1015_g N_VPWR_c_1671_n 0.00448951f $X=7.46 $Y=2.75 $X2=0
+ $Y2=0
cc_936 N_A_1474_446#_c_1277_n N_VPWR_c_1671_n 0.00775326f $X=7.785 $Y=2.215
+ $X2=0 $Y2=0
cc_937 N_A_1474_446#_c_1278_n N_VPWR_c_1671_n 0.0188859f $X=8.77 $Y=2.475 $X2=0
+ $Y2=0
cc_938 N_A_1474_446#_c_1282_n N_VPWR_c_1671_n 0.0437847f $X=8.685 $Y=2.19 $X2=0
+ $Y2=0
cc_939 N_A_1474_446#_c_1267_n A_1817_392# 2.52189e-19 $X=9.3 $Y=1.97 $X2=-0.19
+ $Y2=-0.245
cc_940 N_A_1474_446#_c_1302_n A_1817_392# 0.0069992f $X=9.385 $Y=2.19 $X2=-0.19
+ $Y2=-0.245
cc_941 N_A_1474_446#_M1002_g N_Q_N_c_1851_n 0.00921093f $X=11.015 $Y=0.74 $X2=0
+ $Y2=0
cc_942 N_A_1474_446#_c_1265_n N_Q_N_c_1851_n 0.00216172f $X=12.005 $Y=0.94 $X2=0
+ $Y2=0
cc_943 N_A_1474_446#_M1002_g N_Q_N_c_1852_n 0.00419661f $X=11.015 $Y=0.74 $X2=0
+ $Y2=0
cc_944 N_A_1474_446#_c_1261_n N_Q_N_c_1852_n 0.00478419f $X=11.635 $Y=1.485
+ $X2=0 $Y2=0
cc_945 N_A_1474_446#_c_1262_n N_Q_N_c_1852_n 0.00216172f $X=11.71 $Y=1.32 $X2=0
+ $Y2=0
cc_946 N_A_1474_446#_c_1268_n N_Q_N_c_1852_n 0.00404482f $X=10.955 $Y=1.485
+ $X2=0 $Y2=0
cc_947 N_A_1474_446#_M1008_g Q_N 0.00169947f $X=10.98 $Y=2.4 $X2=0 $Y2=0
cc_948 N_A_1474_446#_c_1261_n Q_N 0.00585625f $X=11.635 $Y=1.485 $X2=0 $Y2=0
cc_949 N_A_1474_446#_c_1275_n Q_N 0.00162322f $X=11.95 $Y=1.975 $X2=0 $Y2=0
cc_950 N_A_1474_446#_c_1281_n Q_N 0.0149941f $X=10.865 $Y=2.24 $X2=0 $Y2=0
cc_951 N_A_1474_446#_c_1275_n Q_N 0.00343581f $X=11.95 $Y=1.975 $X2=0 $Y2=0
cc_952 N_A_1474_446#_M1008_g N_Q_N_c_1853_n 0.00113201f $X=10.98 $Y=2.4 $X2=0
+ $Y2=0
cc_953 N_A_1474_446#_M1002_g N_Q_N_c_1853_n 0.00312482f $X=11.015 $Y=0.74 $X2=0
+ $Y2=0
cc_954 N_A_1474_446#_c_1261_n N_Q_N_c_1853_n 0.0224523f $X=11.635 $Y=1.485 $X2=0
+ $Y2=0
cc_955 N_A_1474_446#_c_1263_n N_Q_N_c_1853_n 0.00162322f $X=11.71 $Y=1.825 $X2=0
+ $Y2=0
cc_956 N_A_1474_446#_c_1281_n N_Q_N_c_1853_n 0.00510544f $X=10.865 $Y=2.24 $X2=0
+ $Y2=0
cc_957 N_A_1474_446#_c_1268_n N_Q_N_c_1853_n 0.0236023f $X=10.955 $Y=1.485 $X2=0
+ $Y2=0
cc_958 N_A_1474_446#_c_1264_n Q 9.2113e-19 $X=12.005 $Y=0.865 $X2=0 $Y2=0
cc_959 N_A_1474_446#_M1021_g N_VGND_c_1906_n 0.00608281f $X=7.955 $Y=0.58 $X2=0
+ $Y2=0
cc_960 N_A_1474_446#_M1002_g N_VGND_c_1907_n 0.00611132f $X=11.015 $Y=0.74 $X2=0
+ $Y2=0
cc_961 N_A_1474_446#_c_1268_n N_VGND_c_1907_n 0.0038303f $X=10.955 $Y=1.485
+ $X2=0 $Y2=0
cc_962 N_A_1474_446#_c_1269_n N_VGND_c_1907_n 0.00189639f $X=10.955 $Y=1.485
+ $X2=0 $Y2=0
cc_963 N_A_1474_446#_c_1264_n N_VGND_c_1908_n 0.0122327f $X=12.005 $Y=0.865
+ $X2=0 $Y2=0
cc_964 N_A_1474_446#_M1002_g N_VGND_c_1912_n 0.00434272f $X=11.015 $Y=0.74 $X2=0
+ $Y2=0
cc_965 N_A_1474_446#_c_1264_n N_VGND_c_1912_n 0.00383152f $X=12.005 $Y=0.865
+ $X2=0 $Y2=0
cc_966 N_A_1474_446#_M1021_g N_VGND_c_1916_n 0.00461464f $X=7.955 $Y=0.58 $X2=0
+ $Y2=0
cc_967 N_A_1474_446#_M1021_g N_VGND_c_1919_n 0.00910155f $X=7.955 $Y=0.58 $X2=0
+ $Y2=0
cc_968 N_A_1474_446#_M1002_g N_VGND_c_1919_n 0.00826383f $X=11.015 $Y=0.74 $X2=0
+ $Y2=0
cc_969 N_A_1474_446#_c_1264_n N_VGND_c_1919_n 0.00762539f $X=12.005 $Y=0.865
+ $X2=0 $Y2=0
cc_970 N_A_1474_446#_c_1265_n N_VGND_c_1919_n 0.00127635f $X=12.005 $Y=0.94
+ $X2=0 $Y2=0
cc_971 N_A_1474_446#_M1027_d N_A_1708_74#_c_2093_n 0.00182219f $X=9.04 $Y=0.37
+ $X2=0 $Y2=0
cc_972 N_A_1474_446#_c_1324_n N_A_1708_74#_c_2093_n 0.0163672f $X=9.3 $Y=0.777
+ $X2=0 $Y2=0
cc_973 N_A_1474_446#_c_1267_n N_A_1708_74#_c_2100_n 0.00421225f $X=9.3 $Y=1.97
+ $X2=0 $Y2=0
cc_974 N_A_1474_446#_c_1324_n N_A_1708_74#_c_2100_n 0.0267408f $X=9.3 $Y=0.777
+ $X2=0 $Y2=0
cc_975 N_A_1314_424#_M1010_g N_VPWR_c_1654_n 0.00167187f $X=8.995 $Y=2.46 $X2=0
+ $Y2=0
cc_976 N_A_1314_424#_M1010_g N_VPWR_c_1657_n 0.005209f $X=8.995 $Y=2.46 $X2=0
+ $Y2=0
cc_977 N_A_1314_424#_M1010_g N_VPWR_c_1649_n 0.00983825f $X=8.995 $Y=2.46 $X2=0
+ $Y2=0
cc_978 N_A_1314_424#_M1010_g N_VPWR_c_1671_n 6.41206e-19 $X=8.995 $Y=2.46 $X2=0
+ $Y2=0
cc_979 N_A_1314_424#_c_1442_n N_VGND_c_1906_n 0.0225846f $X=8.78 $Y=1.215 $X2=0
+ $Y2=0
cc_980 N_A_1314_424#_c_1446_n N_VGND_c_1906_n 3.01761e-19 $X=8.945 $Y=1.22 $X2=0
+ $Y2=0
cc_981 N_A_1314_424#_c_1446_n N_VGND_c_1917_n 0.00278247f $X=8.945 $Y=1.22 $X2=0
+ $Y2=0
cc_982 N_A_1314_424#_c_1446_n N_VGND_c_1919_n 0.00354282f $X=8.945 $Y=1.22 $X2=0
+ $Y2=0
cc_983 N_A_1314_424#_c_1442_n N_A_1708_74#_c_2096_n 0.0228868f $X=8.78 $Y=1.215
+ $X2=0 $Y2=0
cc_984 N_A_1314_424#_c_1445_n N_A_1708_74#_c_2096_n 5.40259e-19 $X=8.945
+ $Y=1.385 $X2=0 $Y2=0
cc_985 N_A_1314_424#_c_1446_n N_A_1708_74#_c_2096_n 0.0072469f $X=8.945 $Y=1.22
+ $X2=0 $Y2=0
cc_986 N_A_1314_424#_c_1446_n N_A_1708_74#_c_2093_n 0.010054f $X=8.945 $Y=1.22
+ $X2=0 $Y2=0
cc_987 N_A_1314_424#_c_1446_n N_A_1708_74#_c_2094_n 0.00188363f $X=8.945 $Y=1.22
+ $X2=0 $Y2=0
cc_988 N_RESET_B_M1000_g N_VPWR_c_1654_n 7.4425e-19 $X=10.465 $Y=2.16 $X2=0
+ $Y2=0
cc_989 N_RESET_B_M1000_g N_VPWR_c_1655_n 8.6256e-19 $X=10.465 $Y=2.16 $X2=0
+ $Y2=0
cc_990 N_RESET_B_M1000_g N_VPWR_c_1662_n 0.00377165f $X=10.465 $Y=2.16 $X2=0
+ $Y2=0
cc_991 N_RESET_B_M1000_g N_VPWR_c_1649_n 0.00493777f $X=10.465 $Y=2.16 $X2=0
+ $Y2=0
cc_992 N_RESET_B_M1007_g N_Q_N_c_1851_n 8.54515e-19 $X=10.435 $Y=0.58 $X2=0
+ $Y2=0
cc_993 N_RESET_B_c_1547_n N_Q_N_c_1852_n 0.00485681f $X=10.415 $Y=1.145 $X2=0
+ $Y2=0
cc_994 N_RESET_B_M1007_g N_VGND_c_1907_n 0.00611788f $X=10.435 $Y=0.58 $X2=0
+ $Y2=0
cc_995 N_RESET_B_c_1546_n N_VGND_c_1907_n 3.75842e-19 $X=10.415 $Y=1.145 $X2=0
+ $Y2=0
cc_996 N_RESET_B_c_1547_n N_VGND_c_1907_n 0.001241f $X=10.415 $Y=1.145 $X2=0
+ $Y2=0
cc_997 N_RESET_B_M1007_g N_VGND_c_1917_n 0.00433162f $X=10.435 $Y=0.58 $X2=0
+ $Y2=0
cc_998 N_RESET_B_M1007_g N_VGND_c_1919_n 0.00822956f $X=10.435 $Y=0.58 $X2=0
+ $Y2=0
cc_999 N_RESET_B_M1007_g N_A_1708_74#_c_2093_n 0.00260004f $X=10.435 $Y=0.58
+ $X2=0 $Y2=0
cc_1000 N_RESET_B_M1007_g N_A_1708_74#_c_2100_n 6.08874e-19 $X=10.435 $Y=0.58
+ $X2=0 $Y2=0
cc_1001 N_A_2320_410#_M1037_g N_VPWR_c_1656_n 0.00462997f $X=12.465 $Y=2.4 $X2=0
+ $Y2=0
cc_1002 N_A_2320_410#_c_1590_n N_VPWR_c_1656_n 0.00557956f $X=12.375 $Y=1.42
+ $X2=0 $Y2=0
cc_1003 N_A_2320_410#_c_1597_n N_VPWR_c_1656_n 0.0309652f $X=11.765 $Y=2.155
+ $X2=0 $Y2=0
cc_1004 N_A_2320_410#_c_1593_n N_VPWR_c_1656_n 0.016421f $X=12.19 $Y=1.42 $X2=0
+ $Y2=0
cc_1005 N_A_2320_410#_c_1595_n N_VPWR_c_1656_n 0.011338f $X=11.765 $Y=2.03 $X2=0
+ $Y2=0
cc_1006 N_A_2320_410#_c_1598_n N_VPWR_c_1663_n 0.00854762f $X=11.725 $Y=2.195
+ $X2=0 $Y2=0
cc_1007 N_A_2320_410#_M1037_g N_VPWR_c_1664_n 0.005209f $X=12.465 $Y=2.4 $X2=0
+ $Y2=0
cc_1008 N_A_2320_410#_M1037_g N_VPWR_c_1649_n 0.00991105f $X=12.465 $Y=2.4 $X2=0
+ $Y2=0
cc_1009 N_A_2320_410#_c_1598_n N_VPWR_c_1649_n 0.00873555f $X=11.725 $Y=2.195
+ $X2=0 $Y2=0
cc_1010 N_A_2320_410#_c_1592_n N_Q_N_c_1851_n 0.0696665f $X=11.79 $Y=0.58 $X2=0
+ $Y2=0
cc_1011 N_A_2320_410#_c_1597_n Q_N 0.0331074f $X=11.765 $Y=2.155 $X2=0 $Y2=0
cc_1012 N_A_2320_410#_c_1598_n Q_N 0.0331074f $X=11.725 $Y=2.195 $X2=0 $Y2=0
cc_1013 N_A_2320_410#_c_1594_n N_Q_N_c_1853_n 0.0243109f $X=11.757 $Y=1.42 $X2=0
+ $Y2=0
cc_1014 N_A_2320_410#_c_1595_n N_Q_N_c_1853_n 0.0331074f $X=11.765 $Y=2.03 $X2=0
+ $Y2=0
cc_1015 N_A_2320_410#_M1037_g Q 0.0310822f $X=12.465 $Y=2.4 $X2=0 $Y2=0
cc_1016 N_A_2320_410#_M1038_g Q 0.0195724f $X=12.48 $Y=0.74 $X2=0 $Y2=0
cc_1017 N_A_2320_410#_c_1591_n Q 0.0121736f $X=12.465 $Y=1.42 $X2=0 $Y2=0
cc_1018 N_A_2320_410#_c_1592_n Q 0.0117429f $X=11.79 $Y=0.58 $X2=0 $Y2=0
cc_1019 N_A_2320_410#_c_1593_n Q 0.0263169f $X=12.19 $Y=1.42 $X2=0 $Y2=0
cc_1020 N_A_2320_410#_M1038_g N_VGND_c_1908_n 0.00461951f $X=12.48 $Y=0.74 $X2=0
+ $Y2=0
cc_1021 N_A_2320_410#_c_1590_n N_VGND_c_1908_n 0.00443885f $X=12.375 $Y=1.42
+ $X2=0 $Y2=0
cc_1022 N_A_2320_410#_c_1592_n N_VGND_c_1908_n 0.0172426f $X=11.79 $Y=0.58 $X2=0
+ $Y2=0
cc_1023 N_A_2320_410#_c_1593_n N_VGND_c_1908_n 0.00981145f $X=12.19 $Y=1.42
+ $X2=0 $Y2=0
cc_1024 N_A_2320_410#_c_1592_n N_VGND_c_1912_n 0.0103967f $X=11.79 $Y=0.58 $X2=0
+ $Y2=0
cc_1025 N_A_2320_410#_M1038_g N_VGND_c_1918_n 0.00428607f $X=12.48 $Y=0.74 $X2=0
+ $Y2=0
cc_1026 N_A_2320_410#_M1038_g N_VGND_c_1919_n 0.00807033f $X=12.48 $Y=0.74 $X2=0
+ $Y2=0
cc_1027 N_A_2320_410#_c_1592_n N_VGND_c_1919_n 0.00860547f $X=11.79 $Y=0.58
+ $X2=0 $Y2=0
cc_1028 N_VPWR_c_1651_n N_A_422_125#_c_1799_n 0.0134933f $X=2.29 $Y=2.59 $X2=0
+ $Y2=0
cc_1029 N_VPWR_c_1660_n N_A_422_125#_c_1799_n 0.00821391f $X=3.94 $Y=3.33 $X2=0
+ $Y2=0
cc_1030 N_VPWR_c_1649_n N_A_422_125#_c_1799_n 0.0101208f $X=12.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1031 N_VPWR_c_1655_n Q_N 0.0138864f $X=10.755 $Y=2.745 $X2=0 $Y2=0
cc_1032 N_VPWR_c_1656_n Q_N 0.00231337f $X=12.24 $Y=1.985 $X2=0 $Y2=0
cc_1033 N_VPWR_c_1663_n Q_N 0.0150819f $X=12.075 $Y=3.33 $X2=0 $Y2=0
cc_1034 N_VPWR_c_1649_n Q_N 0.0124835f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_1035 N_VPWR_c_1656_n Q 0.0396567f $X=12.24 $Y=1.985 $X2=0 $Y2=0
cc_1036 N_VPWR_c_1664_n Q 0.0147721f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_1037 N_VPWR_c_1649_n Q 0.0121589f $X=12.72 $Y=3.33 $X2=0 $Y2=0
cc_1038 N_A_422_125#_c_1795_n N_VGND_c_1904_n 0.0113416f $X=2.25 $Y=0.835 $X2=0
+ $Y2=0
cc_1039 N_A_422_125#_c_1797_n N_VGND_c_1904_n 0.00676472f $X=2.335 $Y=1 $X2=0
+ $Y2=0
cc_1040 N_A_422_125#_c_1795_n N_VGND_c_1915_n 0.00503013f $X=2.25 $Y=0.835 $X2=0
+ $Y2=0
cc_1041 N_A_422_125#_c_1795_n N_VGND_c_1919_n 0.00656676f $X=2.25 $Y=0.835 $X2=0
+ $Y2=0
cc_1042 N_Q_N_c_1851_n N_VGND_c_1907_n 0.0185323f $X=11.23 $Y=0.515 $X2=0 $Y2=0
cc_1043 N_Q_N_c_1851_n N_VGND_c_1912_n 0.0174643f $X=11.23 $Y=0.515 $X2=0 $Y2=0
cc_1044 N_Q_N_c_1851_n N_VGND_c_1919_n 0.014399f $X=11.23 $Y=0.515 $X2=0 $Y2=0
cc_1045 Q N_VGND_c_1908_n 0.028733f $X=12.635 $Y=0.47 $X2=0 $Y2=0
cc_1046 Q N_VGND_c_1918_n 0.0147721f $X=12.635 $Y=0.47 $X2=0 $Y2=0
cc_1047 Q N_VGND_c_1919_n 0.0121589f $X=12.635 $Y=0.47 $X2=0 $Y2=0
cc_1048 N_VGND_c_1909_n N_A_872_119#_c_2063_n 0.0441117f $X=6.06 $Y=0 $X2=0
+ $Y2=0
cc_1049 N_VGND_c_1919_n N_A_872_119#_c_2063_n 0.0230249f $X=12.72 $Y=0 $X2=0
+ $Y2=0
cc_1050 N_VGND_c_1909_n N_A_872_119#_c_2064_n 0.0262823f $X=6.06 $Y=0 $X2=0
+ $Y2=0
cc_1051 N_VGND_c_1915_n N_A_872_119#_c_2064_n 0.02008f $X=3.56 $Y=0 $X2=0 $Y2=0
cc_1052 N_VGND_c_1919_n N_A_872_119#_c_2064_n 0.013689f $X=12.72 $Y=0 $X2=0
+ $Y2=0
cc_1053 N_VGND_c_1905_n N_A_872_119#_c_2065_n 0.0290702f $X=6.245 $Y=0.485 $X2=0
+ $Y2=0
cc_1054 N_VGND_c_1909_n N_A_872_119#_c_2065_n 0.0215843f $X=6.06 $Y=0 $X2=0
+ $Y2=0
cc_1055 N_VGND_c_1919_n N_A_872_119#_c_2065_n 0.0110944f $X=12.72 $Y=0 $X2=0
+ $Y2=0
cc_1056 N_VGND_c_1917_n N_A_1708_74#_c_2093_n 0.0525586f $X=10.565 $Y=0 $X2=0
+ $Y2=0
cc_1057 N_VGND_c_1919_n N_A_1708_74#_c_2093_n 0.0294129f $X=12.72 $Y=0 $X2=0
+ $Y2=0
cc_1058 N_VGND_c_1906_n N_A_1708_74#_c_2094_n 0.0117237f $X=8.25 $Y=0.495 $X2=0
+ $Y2=0
cc_1059 N_VGND_c_1917_n N_A_1708_74#_c_2094_n 0.023633f $X=10.565 $Y=0 $X2=0
+ $Y2=0
cc_1060 N_VGND_c_1919_n N_A_1708_74#_c_2094_n 0.0127274f $X=12.72 $Y=0 $X2=0
+ $Y2=0

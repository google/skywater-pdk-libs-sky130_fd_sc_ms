* File: sky130_fd_sc_ms__o32ai_4.pxi.spice
* Created: Fri Aug 28 18:04:25 2020
* 
x_PM_SKY130_FD_SC_MS__O32AI_4%B2 N_B2_M1015_g N_B2_M1022_g N_B2_M1030_g
+ N_B2_M1016_g N_B2_M1019_g N_B2_M1031_g N_B2_M1020_g N_B2_M1032_g B2 B2 B2 B2
+ N_B2_c_158_n PM_SKY130_FD_SC_MS__O32AI_4%B2
x_PM_SKY130_FD_SC_MS__O32AI_4%B1 N_B1_M1012_g N_B1_M1000_g N_B1_M1023_g
+ N_B1_M1004_g N_B1_M1025_g N_B1_M1011_g N_B1_M1028_g N_B1_M1014_g B1 B1 B1 B1
+ B1 N_B1_c_242_n PM_SKY130_FD_SC_MS__O32AI_4%B1
x_PM_SKY130_FD_SC_MS__O32AI_4%A3 N_A3_M1001_g N_A3_c_335_n N_A3_c_336_n
+ N_A3_M1006_g N_A3_M1033_g N_A3_M1013_g N_A3_M1036_g N_A3_M1029_g N_A3_M1038_g
+ N_A3_M1037_g A3 A3 A3 N_A3_c_341_n PM_SKY130_FD_SC_MS__O32AI_4%A3
x_PM_SKY130_FD_SC_MS__O32AI_4%A2 N_A2_c_436_n N_A2_M1003_g N_A2_M1005_g
+ N_A2_M1007_g N_A2_M1008_g N_A2_M1009_g N_A2_M1017_g N_A2_M1010_g N_A2_M1034_g
+ A2 A2 A2 A2 A2 N_A2_c_435_n PM_SKY130_FD_SC_MS__O32AI_4%A2
x_PM_SKY130_FD_SC_MS__O32AI_4%A1 N_A1_M1002_g N_A1_M1021_g N_A1_M1018_g
+ N_A1_M1024_g N_A1_M1027_g N_A1_M1026_g N_A1_M1039_g N_A1_M1035_g A1 A1 A1 A1
+ A1 N_A1_c_532_n PM_SKY130_FD_SC_MS__O32AI_4%A1
x_PM_SKY130_FD_SC_MS__O32AI_4%A_27_368# N_A_27_368#_M1015_s N_A_27_368#_M1016_s
+ N_A_27_368#_M1020_s N_A_27_368#_M1023_d N_A_27_368#_M1028_d
+ N_A_27_368#_c_610_n N_A_27_368#_c_611_n N_A_27_368#_c_612_n
+ N_A_27_368#_c_623_n N_A_27_368#_c_613_n N_A_27_368#_c_629_n
+ N_A_27_368#_c_630_n N_A_27_368#_c_632_n N_A_27_368#_c_634_n
+ N_A_27_368#_c_614_n N_A_27_368#_c_615_n N_A_27_368#_c_616_n
+ PM_SKY130_FD_SC_MS__O32AI_4%A_27_368#
x_PM_SKY130_FD_SC_MS__O32AI_4%Y N_Y_M1022_s N_Y_M1031_s N_Y_M1000_s N_Y_M1011_s
+ N_Y_M1015_d N_Y_M1019_d N_Y_M1006_d N_Y_M1029_d N_Y_c_689_n N_Y_c_692_n
+ N_Y_c_678_n N_Y_c_679_n N_Y_c_704_n N_Y_c_687_n N_Y_c_680_n N_Y_c_729_n
+ N_Y_c_681_n N_Y_c_735_n N_Y_c_682_n N_Y_c_757_n N_Y_c_683_n N_Y_c_707_n
+ N_Y_c_709_n N_Y_c_684_n N_Y_c_685_n N_Y_c_686_n N_Y_c_767_n N_Y_c_772_n Y
+ PM_SKY130_FD_SC_MS__O32AI_4%Y
x_PM_SKY130_FD_SC_MS__O32AI_4%VPWR N_VPWR_M1012_s N_VPWR_M1025_s N_VPWR_M1021_s
+ N_VPWR_M1024_s N_VPWR_M1035_s N_VPWR_c_837_n N_VPWR_c_838_n N_VPWR_c_839_n
+ N_VPWR_c_840_n N_VPWR_c_841_n N_VPWR_c_842_n N_VPWR_c_843_n N_VPWR_c_844_n
+ N_VPWR_c_845_n N_VPWR_c_846_n N_VPWR_c_847_n N_VPWR_c_848_n VPWR
+ N_VPWR_c_849_n N_VPWR_c_850_n N_VPWR_c_851_n N_VPWR_c_836_n
+ PM_SKY130_FD_SC_MS__O32AI_4%VPWR
x_PM_SKY130_FD_SC_MS__O32AI_4%A_861_368# N_A_861_368#_M1006_s
+ N_A_861_368#_M1013_s N_A_861_368#_M1037_s N_A_861_368#_M1007_s
+ N_A_861_368#_M1010_s N_A_861_368#_c_955_n N_A_861_368#_c_956_n
+ N_A_861_368#_c_957_n N_A_861_368#_c_985_n N_A_861_368#_c_958_n
+ N_A_861_368#_c_970_n N_A_861_368#_c_959_n N_A_861_368#_c_973_n
+ N_A_861_368#_c_960_n N_A_861_368#_c_961_n N_A_861_368#_c_962_n
+ N_A_861_368#_c_963_n N_A_861_368#_c_964_n
+ PM_SKY130_FD_SC_MS__O32AI_4%A_861_368#
x_PM_SKY130_FD_SC_MS__O32AI_4%A_1333_368# N_A_1333_368#_M1003_d
+ N_A_1333_368#_M1009_d N_A_1333_368#_M1021_d N_A_1333_368#_M1026_d
+ N_A_1333_368#_c_1017_n N_A_1333_368#_c_1014_n N_A_1333_368#_c_1015_n
+ N_A_1333_368#_c_1038_n N_A_1333_368#_c_1042_n N_A_1333_368#_c_1016_n
+ N_A_1333_368#_c_1024_n N_A_1333_368#_c_1029_n N_A_1333_368#_c_1049_n
+ PM_SKY130_FD_SC_MS__O32AI_4%A_1333_368#
x_PM_SKY130_FD_SC_MS__O32AI_4%A_27_74# N_A_27_74#_M1022_d N_A_27_74#_M1030_d
+ N_A_27_74#_M1032_d N_A_27_74#_M1004_d N_A_27_74#_M1014_d N_A_27_74#_M1033_d
+ N_A_27_74#_M1038_d N_A_27_74#_M1008_s N_A_27_74#_M1034_s N_A_27_74#_M1018_s
+ N_A_27_74#_M1039_s N_A_27_74#_c_1073_n N_A_27_74#_c_1074_n N_A_27_74#_c_1075_n
+ N_A_27_74#_c_1099_n N_A_27_74#_c_1076_n N_A_27_74#_c_1104_n
+ N_A_27_74#_c_1077_n N_A_27_74#_c_1108_n N_A_27_74#_c_1078_n
+ N_A_27_74#_c_1115_n N_A_27_74#_c_1117_n N_A_27_74#_c_1119_n
+ N_A_27_74#_c_1079_n N_A_27_74#_c_1123_n N_A_27_74#_c_1080_n
+ N_A_27_74#_c_1081_n N_A_27_74#_c_1082_n N_A_27_74#_c_1083_n
+ N_A_27_74#_c_1084_n N_A_27_74#_c_1085_n N_A_27_74#_c_1086_n
+ N_A_27_74#_c_1087_n N_A_27_74#_c_1088_n N_A_27_74#_c_1089_n
+ N_A_27_74#_c_1090_n N_A_27_74#_c_1125_n N_A_27_74#_c_1091_n
+ N_A_27_74#_c_1092_n N_A_27_74#_c_1093_n N_A_27_74#_c_1094_n
+ PM_SKY130_FD_SC_MS__O32AI_4%A_27_74#
x_PM_SKY130_FD_SC_MS__O32AI_4%VGND N_VGND_M1001_s N_VGND_M1036_s N_VGND_M1005_d
+ N_VGND_M1017_d N_VGND_M1002_d N_VGND_M1027_d N_VGND_c_1257_n N_VGND_c_1258_n
+ N_VGND_c_1259_n N_VGND_c_1260_n N_VGND_c_1261_n N_VGND_c_1262_n
+ N_VGND_c_1263_n N_VGND_c_1264_n N_VGND_c_1265_n N_VGND_c_1266_n VGND
+ N_VGND_c_1267_n N_VGND_c_1268_n N_VGND_c_1269_n N_VGND_c_1270_n
+ N_VGND_c_1271_n N_VGND_c_1272_n N_VGND_c_1273_n N_VGND_c_1274_n
+ N_VGND_c_1275_n N_VGND_c_1276_n PM_SKY130_FD_SC_MS__O32AI_4%VGND
cc_1 VNB N_B2_M1022_g 0.0309142f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_B2_M1030_g 0.0225305f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_3 VNB N_B2_M1031_g 0.0227565f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_4 VNB N_B2_M1032_g 0.0227237f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_5 VNB B2 0.0149358f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_6 VNB N_B2_c_158_n 0.0768688f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.515
cc_7 VNB N_B1_M1000_g 0.0234867f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_8 VNB N_B1_M1004_g 0.023521f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_9 VNB N_B1_M1011_g 0.023521f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_10 VNB N_B1_M1014_g 0.0236802f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_11 VNB B1 0.00801322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B1_c_242_n 0.081983f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.605
cc_13 VNB N_A3_M1001_g 0.0252062f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_14 VNB N_A3_c_335_n 0.00823166f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_15 VNB N_A3_c_336_n 0.0105593f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_16 VNB N_A3_M1033_g 0.0252948f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.68
cc_17 VNB N_A3_M1036_g 0.0228207f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.35
cc_18 VNB N_A3_M1038_g 0.0257126f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.35
cc_19 VNB A3 0.00134275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A3_c_341_n 0.0753012f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.515
cc_21 VNB N_A2_M1005_g 0.029538f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_22 VNB N_A2_M1008_g 0.024924f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_23 VNB N_A2_M1017_g 0.024924f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_24 VNB N_A2_M1034_g 0.0263392f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_25 VNB A2 0.00778854f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_26 VNB N_A2_c_435_n 0.0904757f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.515
cc_27 VNB N_A1_M1002_g 0.0249391f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_28 VNB N_A1_M1018_g 0.0240482f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_29 VNB N_A1_M1027_g 0.0240482f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_30 VNB N_A1_M1039_g 0.0328666f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_31 VNB A1 0.0267679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A1_c_532_n 0.0930779f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=1.515
cc_33 VNB N_Y_c_678_n 0.00314141f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_34 VNB N_Y_c_679_n 0.00228572f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_35 VNB N_Y_c_680_n 0.00578048f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_36 VNB N_Y_c_681_n 0.00304954f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.515
cc_37 VNB N_Y_c_682_n 0.0188349f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.515
cc_38 VNB N_Y_c_683_n 0.00308421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_Y_c_684_n 0.00184947f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.605
cc_40 VNB N_Y_c_685_n 0.00227118f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=1.605
cc_41 VNB N_Y_c_686_n 0.00227118f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.605
cc_42 VNB N_VPWR_c_836_n 0.462217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_27_74#_c_1073_n 0.0293003f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_44 VNB N_A_27_74#_c_1074_n 0.0026914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_27_74#_c_1075_n 0.00931596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_27_74#_c_1076_n 0.00230691f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.515
cc_47 VNB N_A_27_74#_c_1077_n 0.00280532f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.515
cc_48 VNB N_A_27_74#_c_1078_n 0.00502477f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=1.515
cc_49 VNB N_A_27_74#_c_1079_n 0.00291301f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.605
cc_50 VNB N_A_27_74#_c_1080_n 0.00323083f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.605
cc_51 VNB N_A_27_74#_c_1081_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_27_74#_c_1082_n 0.00323083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_27_74#_c_1083_n 0.00280455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_27_74#_c_1084_n 0.00418647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_27_74#_c_1085_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_27_74#_c_1086_n 0.0128173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_27_74#_c_1087_n 0.0281704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_27_74#_c_1088_n 0.00221218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_27_74#_c_1089_n 0.00221218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_27_74#_c_1090_n 0.00221218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_27_74#_c_1091_n 0.0104699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_27_74#_c_1092_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_27_74#_c_1093_n 0.00772133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_27_74#_c_1094_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1257_n 0.00830625f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.35
cc_66 VNB N_VGND_c_1258_n 0.0174979f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.74
cc_67 VNB N_VGND_c_1259_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_68 VNB N_VGND_c_1260_n 0.00891319f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.74
cc_69 VNB N_VGND_c_1261_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_70 VNB N_VGND_c_1262_n 0.00830803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1263_n 0.0185368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1264_n 0.00516528f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.515
cc_73 VNB N_VGND_c_1265_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.515
cc_74 VNB N_VGND_c_1266_n 0.00571618f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.515
cc_75 VNB N_VGND_c_1267_n 0.10355f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=1.515
cc_76 VNB N_VGND_c_1268_n 0.025997f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.515
cc_77 VNB N_VGND_c_1269_n 0.0271081f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=1.605
cc_78 VNB N_VGND_c_1270_n 0.573724f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.605
cc_79 VNB N_VGND_c_1271_n 0.00632082f $X=-0.19 $Y=-0.245 $X2=1.6 $Y2=1.605
cc_80 VNB N_VGND_c_1272_n 0.00601569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1273_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1274_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1275_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1276_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VPB N_B2_M1015_g 0.0252759f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_86 VPB N_B2_M1016_g 0.0196343f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_87 VPB N_B2_M1019_g 0.0196385f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_88 VPB N_B2_M1020_g 0.0203407f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_89 VPB B2 0.0169612f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_90 VPB N_B2_c_158_n 0.0119229f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.515
cc_91 VPB N_B1_M1012_g 0.0202515f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_92 VPB N_B1_M1023_g 0.020498f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_93 VPB N_B1_M1025_g 0.0206164f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_94 VPB N_B1_M1028_g 0.0259328f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_95 VPB B1 0.0154157f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_B1_c_242_n 0.0173478f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.605
cc_97 VPB N_A3_M1006_g 0.0252952f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.35
cc_98 VPB N_A3_M1013_g 0.0196374f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.68
cc_99 VPB N_A3_M1029_g 0.02001f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.68
cc_100 VPB N_A3_M1037_g 0.0211225f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_101 VPB A3 0.00738419f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_A3_c_341_n 0.0118378f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.515
cc_103 VPB N_A2_c_436_n 0.0164723f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.68
cc_104 VPB N_A2_M1007_g 0.0202197f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_105 VPB N_A2_M1009_g 0.0207967f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_106 VPB N_A2_M1010_g 0.0256828f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_107 VPB A2 0.0159288f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_108 VPB N_A2_c_435_n 0.0275216f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.515
cc_109 VPB N_A1_M1021_g 0.0246442f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_110 VPB N_A1_M1024_g 0.0215821f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_111 VPB N_A1_M1026_g 0.0215821f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.74
cc_112 VPB N_A1_M1035_g 0.0246442f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=0.74
cc_113 VPB A1 0.0210348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A1_c_532_n 0.0236019f $X=-0.19 $Y=1.66 $X2=1.6 $Y2=1.515
cc_115 VPB N_A_27_368#_c_610_n 0.0366851f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_116 VPB N_A_27_368#_c_611_n 0.00192243f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.74
cc_117 VPB N_A_27_368#_c_612_n 0.00965867f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.74
cc_118 VPB N_A_27_368#_c_613_n 0.00422173f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_27_368#_c_614_n 0.00160153f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_27_368#_c_615_n 0.00231675f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.515
cc_121 VPB N_A_27_368#_c_616_n 0.00891286f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.515
cc_122 VPB N_Y_c_687_n 0.0146673f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_Y_c_683_n 0.00116077f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_837_n 0.00768031f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_125 VPB N_VPWR_c_838_n 0.00798265f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=0.74
cc_126 VPB N_VPWR_c_839_n 0.0150737f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_127 VPB N_VPWR_c_840_n 0.00969617f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=0.74
cc_128 VPB N_VPWR_c_841_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_842_n 0.0498587f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_130 VPB N_VPWR_c_843_n 0.0592423f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_844_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_845_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_846_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.515
cc_134 VPB N_VPWR_c_847_n 0.121777f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.515
cc_135 VPB N_VPWR_c_848_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.515
cc_136 VPB N_VPWR_c_849_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.605
cc_137 VPB N_VPWR_c_850_n 0.0196495f $X=-0.19 $Y=1.66 $X2=1.6 $Y2=1.605
cc_138 VPB N_VPWR_c_851_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_836_n 0.117572f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_861_368#_c_955_n 0.00557161f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_141 VPB N_A_861_368#_c_956_n 0.0026202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_861_368#_c_957_n 0.00446997f $X=-0.19 $Y=1.66 $X2=1.425 $Y2=1.35
cc_143 VPB N_A_861_368#_c_958_n 0.0024778f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_144 VPB N_A_861_368#_c_959_n 0.00219299f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_145 VPB N_A_861_368#_c_960_n 0.00697634f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_A_861_368#_c_961_n 0.00559862f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.515
cc_147 VPB N_A_861_368#_c_962_n 0.00123754f $X=-0.19 $Y=1.66 $X2=0.92 $Y2=1.515
cc_148 VPB N_A_861_368#_c_963_n 0.00237203f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=1.515
cc_149 VPB N_A_861_368#_c_964_n 0.0021839f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.515
cc_150 VPB N_A_1333_368#_c_1014_n 0.0175099f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_151 VPB N_A_1333_368#_c_1015_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.425
+ $Y2=0.74
cc_152 VPB N_A_1333_368#_c_1016_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.87 $Y2=1.35
cc_153 N_B2_M1020_g N_B1_M1012_g 0.0258548f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_154 N_B2_M1032_g N_B1_M1000_g 0.0255777f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_155 B2 B1 0.0231673f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_156 N_B2_c_158_n B1 0.00343679f $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_157 B2 N_B1_c_242_n 2.74134e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_158 N_B2_c_158_n N_B1_c_242_n 0.0258548f $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_159 N_B2_M1015_g N_A_27_368#_c_610_n 0.0128843f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_160 N_B2_M1016_g N_A_27_368#_c_610_n 6.27116e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_161 B2 N_A_27_368#_c_610_n 0.0249908f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_162 N_B2_M1015_g N_A_27_368#_c_611_n 0.0116345f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_163 N_B2_M1016_g N_A_27_368#_c_611_n 0.0116345f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_164 N_B2_M1015_g N_A_27_368#_c_612_n 0.00291744f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_165 N_B2_M1015_g N_A_27_368#_c_623_n 5.74986e-19 $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_166 N_B2_M1016_g N_A_27_368#_c_623_n 0.00892729f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_167 N_B2_M1019_g N_A_27_368#_c_613_n 0.0140221f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_168 N_B2_M1020_g N_A_27_368#_c_613_n 0.0139518f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_169 N_B2_M1016_g N_A_27_368#_c_614_n 0.00194226f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_170 N_B2_M1022_g N_Y_c_689_n 0.00698434f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_171 N_B2_M1030_g N_Y_c_689_n 0.00817703f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_172 N_B2_M1031_g N_Y_c_689_n 9.19396e-19 $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_173 N_B2_M1016_g N_Y_c_692_n 0.0142562f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_174 N_B2_M1019_g N_Y_c_692_n 0.0128923f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_175 B2 N_Y_c_692_n 0.042718f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_176 N_B2_c_158_n N_Y_c_692_n 4.90767e-19 $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_177 N_B2_M1030_g N_Y_c_678_n 0.00962629f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_178 N_B2_M1031_g N_Y_c_678_n 0.012847f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_179 B2 N_Y_c_678_n 0.0502387f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_180 N_B2_c_158_n N_Y_c_678_n 0.00453387f $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_181 N_B2_M1022_g N_Y_c_679_n 0.00895201f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_182 N_B2_M1030_g N_Y_c_679_n 0.00277825f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_183 B2 N_Y_c_679_n 0.0276692f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_184 N_B2_c_158_n N_Y_c_679_n 0.00266872f $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_185 N_B2_M1032_g N_Y_c_704_n 0.00731251f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_186 N_B2_M1020_g N_Y_c_687_n 0.0174429f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_187 N_B2_M1032_g N_Y_c_680_n 0.0146095f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_188 B2 N_Y_c_707_n 0.0141726f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_189 N_B2_c_158_n N_Y_c_707_n 5.53716e-19 $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_190 N_B2_M1019_g N_Y_c_709_n 8.84614e-19 $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_191 N_B2_M1020_g N_Y_c_709_n 8.84614e-19 $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_192 B2 N_Y_c_709_n 0.0231165f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_193 N_B2_c_158_n N_Y_c_709_n 5.54423e-19 $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_194 N_B2_M1032_g N_Y_c_684_n 0.00274828f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_195 B2 N_Y_c_684_n 0.0202859f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_196 N_B2_c_158_n N_Y_c_684_n 0.0030744f $X=1.87 $Y=1.515 $X2=0 $Y2=0
cc_197 N_B2_M1016_g Y 4.47651e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_198 N_B2_M1019_g Y 0.00987781f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_199 N_B2_M1020_g Y 0.00966359f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_200 N_B2_M1015_g N_VPWR_c_843_n 0.00333896f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_201 N_B2_M1016_g N_VPWR_c_843_n 0.00333896f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_202 N_B2_M1019_g N_VPWR_c_843_n 0.00333926f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_203 N_B2_M1020_g N_VPWR_c_843_n 0.00333926f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_204 N_B2_M1015_g N_VPWR_c_836_n 0.00426427f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_205 N_B2_M1016_g N_VPWR_c_836_n 0.00422685f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_206 N_B2_M1019_g N_VPWR_c_836_n 0.00422687f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_207 N_B2_M1020_g N_VPWR_c_836_n 0.00422798f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_208 N_B2_M1022_g N_A_27_74#_c_1073_n 0.00159289f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_209 B2 N_A_27_74#_c_1073_n 0.0142937f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_210 N_B2_M1022_g N_A_27_74#_c_1074_n 0.0132617f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_211 N_B2_M1030_g N_A_27_74#_c_1074_n 0.0114512f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_212 N_B2_M1031_g N_A_27_74#_c_1099_n 0.00812239f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_213 N_B2_M1032_g N_A_27_74#_c_1099_n 6.41487e-19 $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_214 N_B2_M1031_g N_A_27_74#_c_1076_n 0.00824471f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_215 N_B2_M1032_g N_A_27_74#_c_1076_n 0.0116325f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_216 N_B2_M1031_g N_A_27_74#_c_1088_n 0.00294698f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_217 N_B2_M1022_g N_VGND_c_1267_n 0.00278271f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_218 N_B2_M1030_g N_VGND_c_1267_n 0.00278271f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_219 N_B2_M1031_g N_VGND_c_1267_n 0.00278247f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_220 N_B2_M1032_g N_VGND_c_1267_n 0.00278271f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_221 N_B2_M1022_g N_VGND_c_1270_n 0.00357086f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_222 N_B2_M1030_g N_VGND_c_1270_n 0.00354087f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_223 N_B2_M1031_g N_VGND_c_1270_n 0.00354233f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_224 N_B2_M1032_g N_VGND_c_1270_n 0.00354163f $X=1.87 $Y=0.74 $X2=0 $Y2=0
cc_225 N_B1_M1014_g N_A3_M1001_g 0.0181896f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_226 B1 N_A3_c_336_n 8.29026e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_227 N_B1_c_242_n N_A3_c_336_n 0.0181896f $X=3.855 $Y=1.515 $X2=0 $Y2=0
cc_228 N_B1_M1028_g A3 3.38614e-19 $X=3.665 $Y=2.4 $X2=0 $Y2=0
cc_229 B1 A3 0.0245233f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_230 N_B1_c_242_n A3 5.89412e-19 $X=3.855 $Y=1.515 $X2=0 $Y2=0
cc_231 B1 N_A3_c_341_n 0.00124924f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_232 N_B1_c_242_n N_A3_c_341_n 0.00205346f $X=3.855 $Y=1.515 $X2=0 $Y2=0
cc_233 N_B1_M1012_g N_A_27_368#_c_613_n 0.00347836f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_234 N_B1_M1012_g N_A_27_368#_c_629_n 8.84614e-19 $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_235 N_B1_M1012_g N_A_27_368#_c_630_n 0.00649085f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_236 N_B1_M1023_g N_A_27_368#_c_630_n 5.41755e-19 $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_237 N_B1_M1012_g N_A_27_368#_c_632_n 0.012696f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_238 N_B1_M1023_g N_A_27_368#_c_632_n 0.0126573f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_239 N_B1_M1025_g N_A_27_368#_c_634_n 0.0127584f $X=3.205 $Y=2.4 $X2=0 $Y2=0
cc_240 N_B1_M1028_g N_A_27_368#_c_634_n 0.0127584f $X=3.665 $Y=2.4 $X2=0 $Y2=0
cc_241 N_B1_M1012_g N_A_27_368#_c_615_n 5.64228e-19 $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_242 N_B1_M1023_g N_A_27_368#_c_615_n 0.00877121f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_243 N_B1_M1025_g N_A_27_368#_c_615_n 0.00881385f $X=3.205 $Y=2.4 $X2=0 $Y2=0
cc_244 N_B1_M1028_g N_A_27_368#_c_615_n 5.64931e-19 $X=3.665 $Y=2.4 $X2=0 $Y2=0
cc_245 N_B1_M1025_g N_A_27_368#_c_616_n 5.69921e-19 $X=3.205 $Y=2.4 $X2=0 $Y2=0
cc_246 N_B1_M1028_g N_A_27_368#_c_616_n 0.00905697f $X=3.665 $Y=2.4 $X2=0 $Y2=0
cc_247 N_B1_M1000_g N_Y_c_704_n 6.35897e-19 $X=2.355 $Y=0.74 $X2=0 $Y2=0
cc_248 N_B1_M1012_g N_Y_c_687_n 0.0116236f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_249 N_B1_M1023_g N_Y_c_687_n 0.0116623f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_250 N_B1_M1025_g N_Y_c_687_n 0.0117247f $X=3.205 $Y=2.4 $X2=0 $Y2=0
cc_251 N_B1_M1028_g N_Y_c_687_n 0.0138478f $X=3.665 $Y=2.4 $X2=0 $Y2=0
cc_252 B1 N_Y_c_687_n 0.147317f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_253 N_B1_c_242_n N_Y_c_687_n 0.00235029f $X=3.855 $Y=1.515 $X2=0 $Y2=0
cc_254 N_B1_M1000_g N_Y_c_680_n 0.0130134f $X=2.355 $Y=0.74 $X2=0 $Y2=0
cc_255 B1 N_Y_c_680_n 0.0325718f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_256 N_B1_c_242_n N_Y_c_680_n 0.00188144f $X=3.855 $Y=1.515 $X2=0 $Y2=0
cc_257 N_B1_M1004_g N_Y_c_729_n 0.00829713f $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_258 N_B1_M1011_g N_Y_c_729_n 6.51423e-19 $X=3.355 $Y=0.74 $X2=0 $Y2=0
cc_259 N_B1_M1004_g N_Y_c_681_n 0.00962629f $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_260 N_B1_M1011_g N_Y_c_681_n 0.0131496f $X=3.355 $Y=0.74 $X2=0 $Y2=0
cc_261 B1 N_Y_c_681_n 0.0494836f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_262 N_B1_c_242_n N_Y_c_681_n 0.00489921f $X=3.855 $Y=1.515 $X2=0 $Y2=0
cc_263 N_B1_M1014_g N_Y_c_735_n 0.00817927f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_264 N_B1_M1014_g N_Y_c_682_n 0.00956562f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_265 B1 N_Y_c_682_n 0.0300444f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_266 N_B1_M1004_g N_Y_c_685_n 0.00317618f $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_267 B1 N_Y_c_685_n 0.02778f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_268 N_B1_c_242_n N_Y_c_685_n 0.00484877f $X=3.855 $Y=1.515 $X2=0 $Y2=0
cc_269 N_B1_M1014_g N_Y_c_686_n 0.00317618f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_270 B1 N_Y_c_686_n 0.02778f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_271 N_B1_c_242_n N_Y_c_686_n 0.00508543f $X=3.855 $Y=1.515 $X2=0 $Y2=0
cc_272 N_B1_M1012_g Y 7.42905e-19 $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_273 N_B1_M1012_g N_VPWR_c_837_n 0.00120619f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_274 N_B1_M1023_g N_VPWR_c_837_n 0.0027763f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_275 N_B1_M1025_g N_VPWR_c_838_n 0.00279439f $X=3.205 $Y=2.4 $X2=0 $Y2=0
cc_276 N_B1_M1028_g N_VPWR_c_838_n 0.0038624f $X=3.665 $Y=2.4 $X2=0 $Y2=0
cc_277 N_B1_M1012_g N_VPWR_c_843_n 0.00517089f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_278 N_B1_M1023_g N_VPWR_c_845_n 0.005209f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_279 N_B1_M1025_g N_VPWR_c_845_n 0.005209f $X=3.205 $Y=2.4 $X2=0 $Y2=0
cc_280 N_B1_M1028_g N_VPWR_c_847_n 0.005209f $X=3.665 $Y=2.4 $X2=0 $Y2=0
cc_281 N_B1_M1012_g N_VPWR_c_836_n 0.00977588f $X=2.305 $Y=2.4 $X2=0 $Y2=0
cc_282 N_B1_M1023_g N_VPWR_c_836_n 0.00982266f $X=2.755 $Y=2.4 $X2=0 $Y2=0
cc_283 N_B1_M1025_g N_VPWR_c_836_n 0.00982367f $X=3.205 $Y=2.4 $X2=0 $Y2=0
cc_284 N_B1_M1028_g N_VPWR_c_836_n 0.00987724f $X=3.665 $Y=2.4 $X2=0 $Y2=0
cc_285 N_B1_M1028_g N_A_861_368#_c_957_n 0.00292778f $X=3.665 $Y=2.4 $X2=0 $Y2=0
cc_286 N_B1_M1000_g N_A_27_74#_c_1104_n 0.00827017f $X=2.355 $Y=0.74 $X2=0 $Y2=0
cc_287 N_B1_M1004_g N_A_27_74#_c_1104_n 6.42138e-19 $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_288 N_B1_M1000_g N_A_27_74#_c_1077_n 0.00854735f $X=2.355 $Y=0.74 $X2=0 $Y2=0
cc_289 N_B1_M1004_g N_A_27_74#_c_1077_n 0.0118445f $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_290 N_B1_M1011_g N_A_27_74#_c_1108_n 0.00830243f $X=3.355 $Y=0.74 $X2=0 $Y2=0
cc_291 N_B1_M1014_g N_A_27_74#_c_1108_n 6.42138e-19 $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_292 N_B1_M1011_g N_A_27_74#_c_1078_n 0.00854735f $X=3.355 $Y=0.74 $X2=0 $Y2=0
cc_293 N_B1_M1014_g N_A_27_74#_c_1078_n 0.0117838f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_294 N_B1_M1000_g N_A_27_74#_c_1089_n 0.00280918f $X=2.355 $Y=0.74 $X2=0 $Y2=0
cc_295 N_B1_M1011_g N_A_27_74#_c_1090_n 0.00294698f $X=3.355 $Y=0.74 $X2=0 $Y2=0
cc_296 N_B1_M1000_g N_VGND_c_1267_n 0.00278247f $X=2.355 $Y=0.74 $X2=0 $Y2=0
cc_297 N_B1_M1004_g N_VGND_c_1267_n 0.00278271f $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_298 N_B1_M1011_g N_VGND_c_1267_n 0.00278247f $X=3.355 $Y=0.74 $X2=0 $Y2=0
cc_299 N_B1_M1014_g N_VGND_c_1267_n 0.00278271f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_300 N_B1_M1000_g N_VGND_c_1270_n 0.00354671f $X=2.355 $Y=0.74 $X2=0 $Y2=0
cc_301 N_B1_M1004_g N_VGND_c_1270_n 0.00354745f $X=2.855 $Y=0.74 $X2=0 $Y2=0
cc_302 N_B1_M1011_g N_VGND_c_1270_n 0.00354743f $X=3.355 $Y=0.74 $X2=0 $Y2=0
cc_303 N_B1_M1014_g N_VGND_c_1270_n 0.00354798f $X=3.855 $Y=0.74 $X2=0 $Y2=0
cc_304 N_A3_M1038_g N_A2_M1005_g 0.00994657f $X=5.875 $Y=0.74 $X2=0 $Y2=0
cc_305 N_A3_c_341_n A2 0.00346788f $X=5.875 $Y=1.515 $X2=0 $Y2=0
cc_306 N_A3_M1037_g N_A2_c_435_n 0.0119473f $X=6.025 $Y=2.4 $X2=0 $Y2=0
cc_307 N_A3_c_341_n N_A2_c_435_n 0.00704011f $X=5.875 $Y=1.515 $X2=0 $Y2=0
cc_308 N_A3_c_335_n N_Y_c_687_n 4.54065e-19 $X=4.585 $Y=1.425 $X2=0 $Y2=0
cc_309 N_A3_c_336_n N_Y_c_687_n 0.00508082f $X=4.43 $Y=1.425 $X2=0 $Y2=0
cc_310 N_A3_M1006_g N_Y_c_687_n 0.0150541f $X=4.675 $Y=2.4 $X2=0 $Y2=0
cc_311 A3 N_Y_c_687_n 0.0196242f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_312 N_A3_M1001_g N_Y_c_735_n 9.19175e-19 $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_313 N_A3_M1001_g N_Y_c_682_n 0.0154867f $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_314 N_A3_c_335_n N_Y_c_682_n 0.00699187f $X=4.585 $Y=1.425 $X2=0 $Y2=0
cc_315 N_A3_M1033_g N_Y_c_682_n 0.0116606f $X=4.945 $Y=0.74 $X2=0 $Y2=0
cc_316 N_A3_M1036_g N_Y_c_682_n 0.010843f $X=5.44 $Y=0.74 $X2=0 $Y2=0
cc_317 N_A3_M1038_g N_Y_c_682_n 0.00829246f $X=5.875 $Y=0.74 $X2=0 $Y2=0
cc_318 A3 N_Y_c_682_n 0.0886829f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_319 N_A3_c_341_n N_Y_c_682_n 0.00904029f $X=5.875 $Y=1.515 $X2=0 $Y2=0
cc_320 N_A3_M1013_g N_Y_c_757_n 0.012931f $X=5.125 $Y=2.4 $X2=0 $Y2=0
cc_321 N_A3_M1029_g N_Y_c_757_n 0.012931f $X=5.575 $Y=2.4 $X2=0 $Y2=0
cc_322 A3 N_Y_c_757_n 0.0384651f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_323 N_A3_c_341_n N_Y_c_757_n 4.84419e-19 $X=5.875 $Y=1.515 $X2=0 $Y2=0
cc_324 N_A3_M1036_g N_Y_c_683_n 5.51338e-19 $X=5.44 $Y=0.74 $X2=0 $Y2=0
cc_325 N_A3_M1029_g N_Y_c_683_n 0.00412904f $X=5.575 $Y=2.4 $X2=0 $Y2=0
cc_326 N_A3_M1038_g N_Y_c_683_n 0.00324012f $X=5.875 $Y=0.74 $X2=0 $Y2=0
cc_327 N_A3_M1037_g N_Y_c_683_n 0.00667908f $X=6.025 $Y=2.4 $X2=0 $Y2=0
cc_328 A3 N_Y_c_683_n 0.0268369f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_329 N_A3_c_341_n N_Y_c_683_n 0.0169033f $X=5.875 $Y=1.515 $X2=0 $Y2=0
cc_330 N_A3_M1006_g N_Y_c_767_n 0.0150733f $X=4.675 $Y=2.4 $X2=0 $Y2=0
cc_331 N_A3_M1013_g N_Y_c_767_n 0.010564f $X=5.125 $Y=2.4 $X2=0 $Y2=0
cc_332 N_A3_M1029_g N_Y_c_767_n 5.73047e-19 $X=5.575 $Y=2.4 $X2=0 $Y2=0
cc_333 A3 N_Y_c_767_n 0.0231165f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_334 N_A3_c_341_n N_Y_c_767_n 5.48413e-19 $X=5.875 $Y=1.515 $X2=0 $Y2=0
cc_335 N_A3_M1013_g N_Y_c_772_n 5.73047e-19 $X=5.125 $Y=2.4 $X2=0 $Y2=0
cc_336 N_A3_M1029_g N_Y_c_772_n 0.0115803f $X=5.575 $Y=2.4 $X2=0 $Y2=0
cc_337 N_A3_M1037_g N_Y_c_772_n 0.0107914f $X=6.025 $Y=2.4 $X2=0 $Y2=0
cc_338 N_A3_c_341_n N_Y_c_772_n 0.00217346f $X=5.875 $Y=1.515 $X2=0 $Y2=0
cc_339 N_A3_M1006_g N_VPWR_c_847_n 0.00333926f $X=4.675 $Y=2.4 $X2=0 $Y2=0
cc_340 N_A3_M1013_g N_VPWR_c_847_n 0.00333926f $X=5.125 $Y=2.4 $X2=0 $Y2=0
cc_341 N_A3_M1029_g N_VPWR_c_847_n 0.00333926f $X=5.575 $Y=2.4 $X2=0 $Y2=0
cc_342 N_A3_M1037_g N_VPWR_c_847_n 0.00333926f $X=6.025 $Y=2.4 $X2=0 $Y2=0
cc_343 N_A3_M1006_g N_VPWR_c_836_n 0.0042782f $X=4.675 $Y=2.4 $X2=0 $Y2=0
cc_344 N_A3_M1013_g N_VPWR_c_836_n 0.00422687f $X=5.125 $Y=2.4 $X2=0 $Y2=0
cc_345 N_A3_M1029_g N_VPWR_c_836_n 0.00422687f $X=5.575 $Y=2.4 $X2=0 $Y2=0
cc_346 N_A3_M1037_g N_VPWR_c_836_n 0.0042367f $X=6.025 $Y=2.4 $X2=0 $Y2=0
cc_347 N_A3_M1006_g N_A_861_368#_c_956_n 0.0149887f $X=4.675 $Y=2.4 $X2=0 $Y2=0
cc_348 N_A3_M1013_g N_A_861_368#_c_956_n 0.0140221f $X=5.125 $Y=2.4 $X2=0 $Y2=0
cc_349 N_A3_M1029_g N_A_861_368#_c_958_n 0.0139779f $X=5.575 $Y=2.4 $X2=0 $Y2=0
cc_350 N_A3_M1037_g N_A_861_368#_c_958_n 0.0143573f $X=6.025 $Y=2.4 $X2=0 $Y2=0
cc_351 N_A3_M1001_g N_A_27_74#_c_1078_n 0.00431215f $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_352 N_A3_M1001_g N_A_27_74#_c_1115_n 0.00528993f $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_353 N_A3_M1033_g N_A_27_74#_c_1115_n 7.96365e-19 $X=4.945 $Y=0.74 $X2=0 $Y2=0
cc_354 N_A3_M1001_g N_A_27_74#_c_1117_n 0.0095689f $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_355 N_A3_M1033_g N_A_27_74#_c_1117_n 0.0095689f $X=4.945 $Y=0.74 $X2=0 $Y2=0
cc_356 N_A3_M1001_g N_A_27_74#_c_1119_n 0.00183649f $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_357 N_A3_M1001_g N_A_27_74#_c_1079_n 8.15591e-19 $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_358 N_A3_M1033_g N_A_27_74#_c_1079_n 0.00681679f $X=4.945 $Y=0.74 $X2=0 $Y2=0
cc_359 N_A3_M1036_g N_A_27_74#_c_1079_n 0.00231544f $X=5.44 $Y=0.74 $X2=0 $Y2=0
cc_360 N_A3_M1036_g N_A_27_74#_c_1123_n 0.0123473f $X=5.44 $Y=0.74 $X2=0 $Y2=0
cc_361 N_A3_M1038_g N_A_27_74#_c_1123_n 0.0133708f $X=5.875 $Y=0.74 $X2=0 $Y2=0
cc_362 N_A3_M1033_g N_A_27_74#_c_1125_n 7.15561e-19 $X=4.945 $Y=0.74 $X2=0 $Y2=0
cc_363 N_A3_M1038_g N_A_27_74#_c_1091_n 0.00824209f $X=5.875 $Y=0.74 $X2=0 $Y2=0
cc_364 N_A3_c_341_n N_A_27_74#_c_1091_n 0.00342133f $X=5.875 $Y=1.515 $X2=0
+ $Y2=0
cc_365 N_A3_M1001_g N_VGND_c_1257_n 0.00280479f $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_366 N_A3_M1033_g N_VGND_c_1257_n 0.00426833f $X=4.945 $Y=0.74 $X2=0 $Y2=0
cc_367 N_A3_M1033_g N_VGND_c_1258_n 0.00331f $X=4.945 $Y=0.74 $X2=0 $Y2=0
cc_368 N_A3_M1036_g N_VGND_c_1258_n 0.00292409f $X=5.44 $Y=0.74 $X2=0 $Y2=0
cc_369 N_A3_M1033_g N_VGND_c_1259_n 5.11412e-19 $X=4.945 $Y=0.74 $X2=0 $Y2=0
cc_370 N_A3_M1036_g N_VGND_c_1259_n 0.0064019f $X=5.44 $Y=0.74 $X2=0 $Y2=0
cc_371 N_A3_M1038_g N_VGND_c_1259_n 0.00879163f $X=5.875 $Y=0.74 $X2=0 $Y2=0
cc_372 N_A3_M1001_g N_VGND_c_1267_n 0.00328073f $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_373 N_A3_M1038_g N_VGND_c_1268_n 0.00281141f $X=5.875 $Y=0.74 $X2=0 $Y2=0
cc_374 N_A3_M1001_g N_VGND_c_1270_n 0.00428419f $X=4.355 $Y=0.74 $X2=0 $Y2=0
cc_375 N_A3_M1033_g N_VGND_c_1270_n 0.00428003f $X=4.945 $Y=0.74 $X2=0 $Y2=0
cc_376 N_A3_M1036_g N_VGND_c_1270_n 0.00380101f $X=5.44 $Y=0.74 $X2=0 $Y2=0
cc_377 N_A3_M1038_g N_VGND_c_1270_n 0.00367885f $X=5.875 $Y=0.74 $X2=0 $Y2=0
cc_378 N_A2_M1034_g N_A1_M1002_g 0.0176969f $X=8.29 $Y=0.74 $X2=0 $Y2=0
cc_379 A2 N_A1_M1021_g 4.77705e-19 $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_380 N_A2_M1010_g A1 3.60426e-19 $X=8.025 $Y=2.4 $X2=0 $Y2=0
cc_381 A2 A1 0.0290088f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_382 N_A2_c_435_n A1 3.10114e-19 $X=8.04 $Y=1.515 $X2=0 $Y2=0
cc_383 A2 N_A1_c_532_n 0.00315089f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_384 N_A2_c_435_n N_A1_c_532_n 0.0176969f $X=8.04 $Y=1.515 $X2=0 $Y2=0
cc_385 N_A2_M1005_g N_Y_c_682_n 0.00162132f $X=6.72 $Y=0.74 $X2=0 $Y2=0
cc_386 N_A2_c_436_n N_Y_c_683_n 7.28528e-19 $X=6.575 $Y=1.77 $X2=0 $Y2=0
cc_387 N_A2_M1005_g N_Y_c_683_n 0.00119795f $X=6.72 $Y=0.74 $X2=0 $Y2=0
cc_388 A2 N_Y_c_683_n 0.0193245f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_389 N_A2_c_435_n N_Y_c_683_n 7.50276e-19 $X=8.04 $Y=1.515 $X2=0 $Y2=0
cc_390 N_A2_M1010_g N_VPWR_c_839_n 8.0317e-19 $X=8.025 $Y=2.4 $X2=0 $Y2=0
cc_391 N_A2_c_436_n N_VPWR_c_847_n 0.00333926f $X=6.575 $Y=1.77 $X2=0 $Y2=0
cc_392 N_A2_M1007_g N_VPWR_c_847_n 0.00333926f $X=7.025 $Y=2.4 $X2=0 $Y2=0
cc_393 N_A2_M1009_g N_VPWR_c_847_n 0.00333896f $X=7.525 $Y=2.4 $X2=0 $Y2=0
cc_394 N_A2_M1010_g N_VPWR_c_847_n 0.00333926f $X=8.025 $Y=2.4 $X2=0 $Y2=0
cc_395 N_A2_c_436_n N_VPWR_c_836_n 0.0042367f $X=6.575 $Y=1.77 $X2=0 $Y2=0
cc_396 N_A2_M1007_g N_VPWR_c_836_n 0.00423176f $X=7.025 $Y=2.4 $X2=0 $Y2=0
cc_397 N_A2_M1009_g N_VPWR_c_836_n 0.00423662f $X=7.525 $Y=2.4 $X2=0 $Y2=0
cc_398 N_A2_M1010_g N_VPWR_c_836_n 0.00428309f $X=8.025 $Y=2.4 $X2=0 $Y2=0
cc_399 A2 N_A_861_368#_c_970_n 0.00713561f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_400 N_A2_c_436_n N_A_861_368#_c_959_n 0.0143573f $X=6.575 $Y=1.77 $X2=0 $Y2=0
cc_401 N_A2_M1007_g N_A_861_368#_c_959_n 0.0142213f $X=7.025 $Y=2.4 $X2=0 $Y2=0
cc_402 N_A2_M1009_g N_A_861_368#_c_973_n 0.00895541f $X=7.525 $Y=2.4 $X2=0 $Y2=0
cc_403 N_A2_M1010_g N_A_861_368#_c_973_n 5.88728e-19 $X=8.025 $Y=2.4 $X2=0 $Y2=0
cc_404 N_A2_M1009_g N_A_861_368#_c_960_n 0.0119307f $X=7.525 $Y=2.4 $X2=0 $Y2=0
cc_405 N_A2_M1010_g N_A_861_368#_c_960_n 0.0153671f $X=8.025 $Y=2.4 $X2=0 $Y2=0
cc_406 N_A2_M1009_g N_A_861_368#_c_964_n 0.00214324f $X=7.525 $Y=2.4 $X2=0 $Y2=0
cc_407 N_A2_M1007_g N_A_1333_368#_c_1017_n 0.0132272f $X=7.025 $Y=2.4 $X2=0
+ $Y2=0
cc_408 N_A2_M1009_g N_A_1333_368#_c_1017_n 0.0145524f $X=7.525 $Y=2.4 $X2=0
+ $Y2=0
cc_409 A2 N_A_1333_368#_c_1017_n 0.046225f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_410 N_A2_c_435_n N_A_1333_368#_c_1017_n 7.5354e-19 $X=8.04 $Y=1.515 $X2=0
+ $Y2=0
cc_411 N_A2_M1010_g N_A_1333_368#_c_1014_n 0.0150541f $X=8.025 $Y=2.4 $X2=0
+ $Y2=0
cc_412 A2 N_A_1333_368#_c_1014_n 0.0407943f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_413 N_A2_c_435_n N_A_1333_368#_c_1014_n 0.00124336f $X=8.04 $Y=1.515 $X2=0
+ $Y2=0
cc_414 N_A2_c_436_n N_A_1333_368#_c_1024_n 0.0104807f $X=6.575 $Y=1.77 $X2=0
+ $Y2=0
cc_415 N_A2_M1007_g N_A_1333_368#_c_1024_n 0.0105922f $X=7.025 $Y=2.4 $X2=0
+ $Y2=0
cc_416 N_A2_M1009_g N_A_1333_368#_c_1024_n 4.54422e-19 $X=7.525 $Y=2.4 $X2=0
+ $Y2=0
cc_417 A2 N_A_1333_368#_c_1024_n 0.0235495f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_418 N_A2_c_435_n N_A_1333_368#_c_1024_n 5.48413e-19 $X=8.04 $Y=1.515 $X2=0
+ $Y2=0
cc_419 N_A2_M1010_g N_A_1333_368#_c_1029_n 0.0147083f $X=8.025 $Y=2.4 $X2=0
+ $Y2=0
cc_420 A2 N_A_1333_368#_c_1029_n 0.0246996f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_421 N_A2_c_435_n N_A_1333_368#_c_1029_n 8.53086e-19 $X=8.04 $Y=1.515 $X2=0
+ $Y2=0
cc_422 N_A2_M1005_g N_A_27_74#_c_1080_n 0.0118691f $X=6.72 $Y=0.74 $X2=0 $Y2=0
cc_423 N_A2_M1008_g N_A_27_74#_c_1080_n 0.0118691f $X=7.29 $Y=0.74 $X2=0 $Y2=0
cc_424 A2 N_A_27_74#_c_1080_n 0.050393f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_425 N_A2_c_435_n N_A_27_74#_c_1080_n 0.00632651f $X=8.04 $Y=1.515 $X2=0 $Y2=0
cc_426 N_A2_M1005_g N_A_27_74#_c_1081_n 6.2873e-19 $X=6.72 $Y=0.74 $X2=0 $Y2=0
cc_427 N_A2_M1008_g N_A_27_74#_c_1081_n 0.00968013f $X=7.29 $Y=0.74 $X2=0 $Y2=0
cc_428 N_A2_M1017_g N_A_27_74#_c_1081_n 0.00968263f $X=7.72 $Y=0.74 $X2=0 $Y2=0
cc_429 N_A2_M1034_g N_A_27_74#_c_1081_n 6.28869e-19 $X=8.29 $Y=0.74 $X2=0 $Y2=0
cc_430 N_A2_M1017_g N_A_27_74#_c_1082_n 0.0118691f $X=7.72 $Y=0.74 $X2=0 $Y2=0
cc_431 N_A2_M1034_g N_A_27_74#_c_1082_n 0.0118691f $X=8.29 $Y=0.74 $X2=0 $Y2=0
cc_432 A2 N_A_27_74#_c_1082_n 0.050393f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_433 N_A2_c_435_n N_A_27_74#_c_1082_n 0.00628711f $X=8.04 $Y=1.515 $X2=0 $Y2=0
cc_434 N_A2_M1017_g N_A_27_74#_c_1083_n 6.28869e-19 $X=7.72 $Y=0.74 $X2=0 $Y2=0
cc_435 N_A2_M1034_g N_A_27_74#_c_1083_n 0.00968736f $X=8.29 $Y=0.74 $X2=0 $Y2=0
cc_436 N_A2_M1005_g N_A_27_74#_c_1091_n 0.0188409f $X=6.72 $Y=0.74 $X2=0 $Y2=0
cc_437 N_A2_M1008_g N_A_27_74#_c_1091_n 6.31055e-19 $X=7.29 $Y=0.74 $X2=0 $Y2=0
cc_438 A2 N_A_27_74#_c_1091_n 0.0267257f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_439 N_A2_c_435_n N_A_27_74#_c_1091_n 0.00365802f $X=8.04 $Y=1.515 $X2=0 $Y2=0
cc_440 N_A2_M1008_g N_A_27_74#_c_1092_n 0.00157732f $X=7.29 $Y=0.74 $X2=0 $Y2=0
cc_441 N_A2_M1017_g N_A_27_74#_c_1092_n 0.00157732f $X=7.72 $Y=0.74 $X2=0 $Y2=0
cc_442 A2 N_A_27_74#_c_1092_n 0.0281223f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_443 N_A2_c_435_n N_A_27_74#_c_1092_n 0.00272398f $X=8.04 $Y=1.515 $X2=0 $Y2=0
cc_444 N_A2_M1034_g N_A_27_74#_c_1093_n 0.00171391f $X=8.29 $Y=0.74 $X2=0 $Y2=0
cc_445 A2 N_A_27_74#_c_1093_n 0.0155598f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_446 N_A2_M1005_g N_VGND_c_1260_n 0.00582842f $X=6.72 $Y=0.74 $X2=0 $Y2=0
cc_447 N_A2_M1008_g N_VGND_c_1260_n 0.00484409f $X=7.29 $Y=0.74 $X2=0 $Y2=0
cc_448 N_A2_M1008_g N_VGND_c_1261_n 0.00434272f $X=7.29 $Y=0.74 $X2=0 $Y2=0
cc_449 N_A2_M1017_g N_VGND_c_1261_n 0.00434272f $X=7.72 $Y=0.74 $X2=0 $Y2=0
cc_450 N_A2_M1017_g N_VGND_c_1262_n 0.00484409f $X=7.72 $Y=0.74 $X2=0 $Y2=0
cc_451 N_A2_M1034_g N_VGND_c_1262_n 0.00484409f $X=8.29 $Y=0.74 $X2=0 $Y2=0
cc_452 N_A2_M1034_g N_VGND_c_1263_n 0.00434272f $X=8.29 $Y=0.74 $X2=0 $Y2=0
cc_453 N_A2_M1034_g N_VGND_c_1264_n 4.99121e-19 $X=8.29 $Y=0.74 $X2=0 $Y2=0
cc_454 N_A2_M1005_g N_VGND_c_1268_n 0.00432683f $X=6.72 $Y=0.74 $X2=0 $Y2=0
cc_455 N_A2_M1005_g N_VGND_c_1270_n 0.00820125f $X=6.72 $Y=0.74 $X2=0 $Y2=0
cc_456 N_A2_M1008_g N_VGND_c_1270_n 0.00821294f $X=7.29 $Y=0.74 $X2=0 $Y2=0
cc_457 N_A2_M1017_g N_VGND_c_1270_n 0.00821294f $X=7.72 $Y=0.74 $X2=0 $Y2=0
cc_458 N_A2_M1034_g N_VGND_c_1270_n 0.00822005f $X=8.29 $Y=0.74 $X2=0 $Y2=0
cc_459 N_A1_M1021_g N_VPWR_c_839_n 0.00501904f $X=9.085 $Y=2.4 $X2=0 $Y2=0
cc_460 N_A1_M1024_g N_VPWR_c_840_n 0.00343717f $X=9.535 $Y=2.4 $X2=0 $Y2=0
cc_461 N_A1_M1026_g N_VPWR_c_840_n 0.00343717f $X=10.085 $Y=2.4 $X2=0 $Y2=0
cc_462 N_A1_M1035_g N_VPWR_c_842_n 0.00501904f $X=10.535 $Y=2.4 $X2=0 $Y2=0
cc_463 A1 N_VPWR_c_842_n 0.0208754f $X=10.715 $Y=1.58 $X2=0 $Y2=0
cc_464 N_A1_M1021_g N_VPWR_c_849_n 0.005209f $X=9.085 $Y=2.4 $X2=0 $Y2=0
cc_465 N_A1_M1024_g N_VPWR_c_849_n 0.005209f $X=9.535 $Y=2.4 $X2=0 $Y2=0
cc_466 N_A1_M1026_g N_VPWR_c_850_n 0.005209f $X=10.085 $Y=2.4 $X2=0 $Y2=0
cc_467 N_A1_M1035_g N_VPWR_c_850_n 0.005209f $X=10.535 $Y=2.4 $X2=0 $Y2=0
cc_468 N_A1_M1021_g N_VPWR_c_836_n 0.00987399f $X=9.085 $Y=2.4 $X2=0 $Y2=0
cc_469 N_A1_M1024_g N_VPWR_c_836_n 0.00982526f $X=9.535 $Y=2.4 $X2=0 $Y2=0
cc_470 N_A1_M1026_g N_VPWR_c_836_n 0.00982526f $X=10.085 $Y=2.4 $X2=0 $Y2=0
cc_471 N_A1_M1035_g N_VPWR_c_836_n 0.00986008f $X=10.535 $Y=2.4 $X2=0 $Y2=0
cc_472 N_A1_M1021_g N_A_1333_368#_c_1014_n 0.0150541f $X=9.085 $Y=2.4 $X2=0
+ $Y2=0
cc_473 A1 N_A_1333_368#_c_1014_n 0.0271602f $X=10.715 $Y=1.58 $X2=0 $Y2=0
cc_474 N_A1_c_532_n N_A_1333_368#_c_1014_n 0.00300231f $X=10.22 $Y=1.515 $X2=0
+ $Y2=0
cc_475 N_A1_M1021_g N_A_1333_368#_c_1015_n 0.0166062f $X=9.085 $Y=2.4 $X2=0
+ $Y2=0
cc_476 N_A1_M1024_g N_A_1333_368#_c_1015_n 0.0119199f $X=9.535 $Y=2.4 $X2=0
+ $Y2=0
cc_477 N_A1_M1026_g N_A_1333_368#_c_1015_n 6.00071e-19 $X=10.085 $Y=2.4 $X2=0
+ $Y2=0
cc_478 N_A1_M1024_g N_A_1333_368#_c_1038_n 0.0134861f $X=9.535 $Y=2.4 $X2=0
+ $Y2=0
cc_479 N_A1_M1026_g N_A_1333_368#_c_1038_n 0.0134861f $X=10.085 $Y=2.4 $X2=0
+ $Y2=0
cc_480 A1 N_A_1333_368#_c_1038_n 0.0471519f $X=10.715 $Y=1.58 $X2=0 $Y2=0
cc_481 N_A1_c_532_n N_A_1333_368#_c_1038_n 0.00102407f $X=10.22 $Y=1.515 $X2=0
+ $Y2=0
cc_482 N_A1_M1026_g N_A_1333_368#_c_1042_n 8.84614e-19 $X=10.085 $Y=2.4 $X2=0
+ $Y2=0
cc_483 N_A1_M1035_g N_A_1333_368#_c_1042_n 0.0025567f $X=10.535 $Y=2.4 $X2=0
+ $Y2=0
cc_484 A1 N_A_1333_368#_c_1042_n 0.0235495f $X=10.715 $Y=1.58 $X2=0 $Y2=0
cc_485 N_A1_c_532_n N_A_1333_368#_c_1042_n 5.57028e-19 $X=10.22 $Y=1.515 $X2=0
+ $Y2=0
cc_486 N_A1_M1024_g N_A_1333_368#_c_1016_n 6.00071e-19 $X=9.535 $Y=2.4 $X2=0
+ $Y2=0
cc_487 N_A1_M1026_g N_A_1333_368#_c_1016_n 0.0119199f $X=10.085 $Y=2.4 $X2=0
+ $Y2=0
cc_488 N_A1_M1035_g N_A_1333_368#_c_1016_n 0.0112644f $X=10.535 $Y=2.4 $X2=0
+ $Y2=0
cc_489 N_A1_M1021_g N_A_1333_368#_c_1049_n 8.84614e-19 $X=9.085 $Y=2.4 $X2=0
+ $Y2=0
cc_490 N_A1_M1024_g N_A_1333_368#_c_1049_n 8.84614e-19 $X=9.535 $Y=2.4 $X2=0
+ $Y2=0
cc_491 A1 N_A_1333_368#_c_1049_n 0.0235495f $X=10.715 $Y=1.58 $X2=0 $Y2=0
cc_492 N_A1_c_532_n N_A_1333_368#_c_1049_n 5.48413e-19 $X=10.22 $Y=1.515 $X2=0
+ $Y2=0
cc_493 N_A1_M1002_g N_A_27_74#_c_1083_n 0.00350341f $X=8.79 $Y=0.74 $X2=0 $Y2=0
cc_494 N_A1_M1002_g N_A_27_74#_c_1084_n 0.0164698f $X=8.79 $Y=0.74 $X2=0 $Y2=0
cc_495 N_A1_M1018_g N_A_27_74#_c_1084_n 0.0115433f $X=9.29 $Y=0.74 $X2=0 $Y2=0
cc_496 A1 N_A_27_74#_c_1084_n 0.0432333f $X=10.715 $Y=1.58 $X2=0 $Y2=0
cc_497 N_A1_c_532_n N_A_27_74#_c_1084_n 0.00432368f $X=10.22 $Y=1.515 $X2=0
+ $Y2=0
cc_498 N_A1_M1002_g N_A_27_74#_c_1085_n 6.94971e-19 $X=8.79 $Y=0.74 $X2=0 $Y2=0
cc_499 N_A1_M1018_g N_A_27_74#_c_1085_n 0.00957028f $X=9.29 $Y=0.74 $X2=0 $Y2=0
cc_500 N_A1_M1027_g N_A_27_74#_c_1085_n 0.00957028f $X=9.72 $Y=0.74 $X2=0 $Y2=0
cc_501 N_A1_M1039_g N_A_27_74#_c_1085_n 6.94971e-19 $X=10.22 $Y=0.74 $X2=0 $Y2=0
cc_502 N_A1_M1027_g N_A_27_74#_c_1086_n 0.0115433f $X=9.72 $Y=0.74 $X2=0 $Y2=0
cc_503 N_A1_M1039_g N_A_27_74#_c_1086_n 0.0162853f $X=10.22 $Y=0.74 $X2=0 $Y2=0
cc_504 A1 N_A_27_74#_c_1086_n 0.0802423f $X=10.715 $Y=1.58 $X2=0 $Y2=0
cc_505 N_A1_c_532_n N_A_27_74#_c_1086_n 0.00607837f $X=10.22 $Y=1.515 $X2=0
+ $Y2=0
cc_506 N_A1_M1039_g N_A_27_74#_c_1087_n 0.0128452f $X=10.22 $Y=0.74 $X2=0 $Y2=0
cc_507 N_A1_M1018_g N_A_27_74#_c_1094_n 0.00157732f $X=9.29 $Y=0.74 $X2=0 $Y2=0
cc_508 N_A1_M1027_g N_A_27_74#_c_1094_n 0.00157732f $X=9.72 $Y=0.74 $X2=0 $Y2=0
cc_509 A1 N_A_27_74#_c_1094_n 0.0281223f $X=10.715 $Y=1.58 $X2=0 $Y2=0
cc_510 N_A1_c_532_n N_A_27_74#_c_1094_n 0.00272398f $X=10.22 $Y=1.515 $X2=0
+ $Y2=0
cc_511 N_A1_M1002_g N_VGND_c_1263_n 0.00383152f $X=8.79 $Y=0.74 $X2=0 $Y2=0
cc_512 N_A1_M1002_g N_VGND_c_1264_n 0.0105599f $X=8.79 $Y=0.74 $X2=0 $Y2=0
cc_513 N_A1_M1018_g N_VGND_c_1264_n 0.00432843f $X=9.29 $Y=0.74 $X2=0 $Y2=0
cc_514 N_A1_M1018_g N_VGND_c_1265_n 0.00434272f $X=9.29 $Y=0.74 $X2=0 $Y2=0
cc_515 N_A1_M1027_g N_VGND_c_1265_n 0.00434272f $X=9.72 $Y=0.74 $X2=0 $Y2=0
cc_516 N_A1_M1027_g N_VGND_c_1266_n 0.00432843f $X=9.72 $Y=0.74 $X2=0 $Y2=0
cc_517 N_A1_M1039_g N_VGND_c_1266_n 0.0132583f $X=10.22 $Y=0.74 $X2=0 $Y2=0
cc_518 N_A1_M1039_g N_VGND_c_1269_n 0.00383152f $X=10.22 $Y=0.74 $X2=0 $Y2=0
cc_519 N_A1_M1002_g N_VGND_c_1270_n 0.00758251f $X=8.79 $Y=0.74 $X2=0 $Y2=0
cc_520 N_A1_M1018_g N_VGND_c_1270_n 0.00820718f $X=9.29 $Y=0.74 $X2=0 $Y2=0
cc_521 N_A1_M1027_g N_VGND_c_1270_n 0.00820718f $X=9.72 $Y=0.74 $X2=0 $Y2=0
cc_522 N_A1_M1039_g N_VGND_c_1270_n 0.00762539f $X=10.22 $Y=0.74 $X2=0 $Y2=0
cc_523 N_A_27_368#_c_611_n N_Y_M1015_d 0.00165831f $X=1.015 $Y=2.99 $X2=0 $Y2=0
cc_524 N_A_27_368#_c_613_n N_Y_M1019_d 0.00165831f $X=1.995 $Y=2.99 $X2=0 $Y2=0
cc_525 N_A_27_368#_M1016_s N_Y_c_692_n 0.00314376f $X=1.045 $Y=1.84 $X2=0 $Y2=0
cc_526 N_A_27_368#_c_623_n N_Y_c_692_n 0.0148589f $X=1.18 $Y=2.455 $X2=0 $Y2=0
cc_527 N_A_27_368#_M1020_s N_Y_c_687_n 0.00450314f $X=1.945 $Y=1.84 $X2=0 $Y2=0
cc_528 N_A_27_368#_M1023_d N_Y_c_687_n 0.00314376f $X=2.845 $Y=1.84 $X2=0 $Y2=0
cc_529 N_A_27_368#_M1028_d N_Y_c_687_n 0.00544479f $X=3.755 $Y=1.84 $X2=0 $Y2=0
cc_530 N_A_27_368#_c_629_n N_Y_c_687_n 0.0149351f $X=2.12 $Y=2.46 $X2=0 $Y2=0
cc_531 N_A_27_368#_c_632_n N_Y_c_687_n 0.0315971f $X=2.815 $Y=2.375 $X2=0 $Y2=0
cc_532 N_A_27_368#_c_634_n N_Y_c_687_n 0.0323235f $X=3.725 $Y=2.375 $X2=0 $Y2=0
cc_533 N_A_27_368#_c_615_n N_Y_c_687_n 0.0171986f $X=2.98 $Y=2.455 $X2=0 $Y2=0
cc_534 N_A_27_368#_c_616_n N_Y_c_687_n 0.0221016f $X=3.89 $Y=2.455 $X2=0 $Y2=0
cc_535 N_A_27_368#_c_611_n N_Y_c_707_n 0.0118736f $X=1.015 $Y=2.99 $X2=0 $Y2=0
cc_536 N_A_27_368#_c_613_n Y 0.0159318f $X=1.995 $Y=2.99 $X2=0 $Y2=0
cc_537 N_A_27_368#_c_632_n N_VPWR_M1012_s 0.00324075f $X=2.815 $Y=2.375
+ $X2=-0.19 $Y2=1.66
cc_538 N_A_27_368#_c_634_n N_VPWR_M1025_s 0.00340221f $X=3.725 $Y=2.375 $X2=0
+ $Y2=0
cc_539 N_A_27_368#_c_613_n N_VPWR_c_837_n 0.0101219f $X=1.995 $Y=2.99 $X2=0
+ $Y2=0
cc_540 N_A_27_368#_c_632_n N_VPWR_c_837_n 0.0126919f $X=2.815 $Y=2.375 $X2=0
+ $Y2=0
cc_541 N_A_27_368#_c_615_n N_VPWR_c_837_n 0.0121684f $X=2.98 $Y=2.455 $X2=0
+ $Y2=0
cc_542 N_A_27_368#_c_634_n N_VPWR_c_838_n 0.0131801f $X=3.725 $Y=2.375 $X2=0
+ $Y2=0
cc_543 N_A_27_368#_c_615_n N_VPWR_c_838_n 0.0121684f $X=2.98 $Y=2.455 $X2=0
+ $Y2=0
cc_544 N_A_27_368#_c_616_n N_VPWR_c_838_n 0.021987f $X=3.89 $Y=2.455 $X2=0 $Y2=0
cc_545 N_A_27_368#_c_611_n N_VPWR_c_843_n 0.0357927f $X=1.015 $Y=2.99 $X2=0
+ $Y2=0
cc_546 N_A_27_368#_c_612_n N_VPWR_c_843_n 0.0235512f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_547 N_A_27_368#_c_613_n N_VPWR_c_843_n 0.0637354f $X=1.995 $Y=2.99 $X2=0
+ $Y2=0
cc_548 N_A_27_368#_c_614_n N_VPWR_c_843_n 0.0178163f $X=1.14 $Y=2.99 $X2=0 $Y2=0
cc_549 N_A_27_368#_c_615_n N_VPWR_c_845_n 0.0144776f $X=2.98 $Y=2.455 $X2=0
+ $Y2=0
cc_550 N_A_27_368#_c_616_n N_VPWR_c_847_n 0.0145644f $X=3.89 $Y=2.455 $X2=0
+ $Y2=0
cc_551 N_A_27_368#_c_611_n N_VPWR_c_836_n 0.0200586f $X=1.015 $Y=2.99 $X2=0
+ $Y2=0
cc_552 N_A_27_368#_c_612_n N_VPWR_c_836_n 0.0126924f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_553 N_A_27_368#_c_613_n N_VPWR_c_836_n 0.0353823f $X=1.995 $Y=2.99 $X2=0
+ $Y2=0
cc_554 N_A_27_368#_c_614_n N_VPWR_c_836_n 0.00958215f $X=1.14 $Y=2.99 $X2=0
+ $Y2=0
cc_555 N_A_27_368#_c_615_n N_VPWR_c_836_n 0.0118404f $X=2.98 $Y=2.455 $X2=0
+ $Y2=0
cc_556 N_A_27_368#_c_616_n N_VPWR_c_836_n 0.0119803f $X=3.89 $Y=2.455 $X2=0
+ $Y2=0
cc_557 N_A_27_368#_c_616_n N_A_861_368#_c_955_n 0.0412426f $X=3.89 $Y=2.455
+ $X2=0 $Y2=0
cc_558 N_A_27_368#_c_616_n N_A_861_368#_c_957_n 0.00536542f $X=3.89 $Y=2.455
+ $X2=0 $Y2=0
cc_559 N_Y_c_687_n N_VPWR_M1012_s 0.0031478f $X=4.735 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_560 N_Y_c_687_n N_VPWR_M1025_s 0.00329864f $X=4.735 $Y=2.035 $X2=0 $Y2=0
cc_561 N_Y_c_687_n N_A_861_368#_M1006_s 0.00613628f $X=4.735 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_562 N_Y_c_757_n N_A_861_368#_M1013_s 0.00314376f $X=5.635 $Y=2.035 $X2=0
+ $Y2=0
cc_563 N_Y_c_687_n N_A_861_368#_c_955_n 0.0197477f $X=4.735 $Y=2.035 $X2=0 $Y2=0
cc_564 N_Y_M1006_d N_A_861_368#_c_956_n 0.00165831f $X=4.765 $Y=1.84 $X2=0 $Y2=0
cc_565 N_Y_c_767_n N_A_861_368#_c_956_n 0.0159318f $X=4.9 $Y=2.115 $X2=0 $Y2=0
cc_566 N_Y_c_757_n N_A_861_368#_c_985_n 0.0126919f $X=5.635 $Y=2.035 $X2=0 $Y2=0
cc_567 N_Y_M1029_d N_A_861_368#_c_958_n 0.00165831f $X=5.665 $Y=1.84 $X2=0 $Y2=0
cc_568 N_Y_c_772_n N_A_861_368#_c_958_n 0.0159318f $X=5.8 $Y=2.115 $X2=0 $Y2=0
cc_569 N_Y_c_678_n N_A_27_74#_M1030_d 0.00250873f $X=1.555 $Y=1.175 $X2=0 $Y2=0
cc_570 N_Y_c_680_n N_A_27_74#_M1032_d 0.00234927f $X=2.475 $Y=1.175 $X2=0 $Y2=0
cc_571 N_Y_c_681_n N_A_27_74#_M1004_d 0.00250873f $X=3.475 $Y=1.175 $X2=0 $Y2=0
cc_572 N_Y_c_682_n N_A_27_74#_M1014_d 0.00250873f $X=5.805 $Y=1.175 $X2=0 $Y2=0
cc_573 N_Y_c_682_n N_A_27_74#_M1033_d 0.00245557f $X=5.805 $Y=1.175 $X2=0 $Y2=0
cc_574 N_Y_c_679_n N_A_27_74#_c_1073_n 0.00233987f $X=0.875 $Y=1.175 $X2=0 $Y2=0
cc_575 N_Y_M1022_s N_A_27_74#_c_1074_n 0.00176461f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_576 N_Y_c_689_n N_A_27_74#_c_1074_n 0.0160271f $X=0.71 $Y=0.86 $X2=0 $Y2=0
cc_577 N_Y_c_678_n N_A_27_74#_c_1074_n 0.00270072f $X=1.555 $Y=1.175 $X2=0 $Y2=0
cc_578 N_Y_c_678_n N_A_27_74#_c_1099_n 0.0209904f $X=1.555 $Y=1.175 $X2=0 $Y2=0
cc_579 N_Y_M1031_s N_A_27_74#_c_1076_n 0.00192406f $X=1.5 $Y=0.37 $X2=0 $Y2=0
cc_580 N_Y_c_678_n N_A_27_74#_c_1076_n 0.00270072f $X=1.555 $Y=1.175 $X2=0 $Y2=0
cc_581 N_Y_c_704_n N_A_27_74#_c_1076_n 0.0143929f $X=1.64 $Y=0.86 $X2=0 $Y2=0
cc_582 N_Y_c_680_n N_A_27_74#_c_1076_n 0.0030261f $X=2.475 $Y=1.175 $X2=0 $Y2=0
cc_583 N_Y_c_680_n N_A_27_74#_c_1104_n 0.0197723f $X=2.475 $Y=1.175 $X2=0 $Y2=0
cc_584 N_Y_M1000_s N_A_27_74#_c_1077_n 0.00250873f $X=2.43 $Y=0.37 $X2=0 $Y2=0
cc_585 N_Y_c_680_n N_A_27_74#_c_1077_n 0.00270072f $X=2.475 $Y=1.175 $X2=0 $Y2=0
cc_586 N_Y_c_729_n N_A_27_74#_c_1077_n 0.0196388f $X=2.64 $Y=0.86 $X2=0 $Y2=0
cc_587 N_Y_c_681_n N_A_27_74#_c_1077_n 0.00270072f $X=3.475 $Y=1.175 $X2=0 $Y2=0
cc_588 N_Y_c_681_n N_A_27_74#_c_1108_n 0.0209904f $X=3.475 $Y=1.175 $X2=0 $Y2=0
cc_589 N_Y_M1011_s N_A_27_74#_c_1078_n 0.00250873f $X=3.43 $Y=0.37 $X2=0 $Y2=0
cc_590 N_Y_c_681_n N_A_27_74#_c_1078_n 0.00270072f $X=3.475 $Y=1.175 $X2=0 $Y2=0
cc_591 N_Y_c_735_n N_A_27_74#_c_1078_n 0.0196388f $X=3.64 $Y=0.86 $X2=0 $Y2=0
cc_592 N_Y_c_682_n N_A_27_74#_c_1078_n 0.00270072f $X=5.805 $Y=1.175 $X2=0 $Y2=0
cc_593 N_Y_c_682_n N_A_27_74#_c_1117_n 0.0405558f $X=5.805 $Y=1.175 $X2=0 $Y2=0
cc_594 N_Y_c_682_n N_A_27_74#_c_1119_n 0.0210664f $X=5.805 $Y=1.175 $X2=0 $Y2=0
cc_595 N_Y_c_682_n N_A_27_74#_c_1123_n 0.0339378f $X=5.805 $Y=1.175 $X2=0 $Y2=0
cc_596 N_Y_c_682_n N_A_27_74#_c_1125_n 0.0204193f $X=5.805 $Y=1.175 $X2=0 $Y2=0
cc_597 N_Y_c_682_n N_A_27_74#_c_1091_n 0.0044173f $X=5.805 $Y=1.175 $X2=0 $Y2=0
cc_598 N_Y_c_682_n N_VGND_M1001_s 0.00355802f $X=5.805 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_599 N_Y_c_682_n N_VGND_M1036_s 0.00182219f $X=5.805 $Y=1.175 $X2=0 $Y2=0
cc_600 N_VPWR_c_847_n N_A_861_368#_c_956_n 0.0459191f $X=8.695 $Y=3.33 $X2=0
+ $Y2=0
cc_601 N_VPWR_c_836_n N_A_861_368#_c_956_n 0.0258001f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_602 N_VPWR_c_847_n N_A_861_368#_c_957_n 0.0179217f $X=8.695 $Y=3.33 $X2=0
+ $Y2=0
cc_603 N_VPWR_c_836_n N_A_861_368#_c_957_n 0.00971942f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_604 N_VPWR_c_847_n N_A_861_368#_c_958_n 0.0446307f $X=8.695 $Y=3.33 $X2=0
+ $Y2=0
cc_605 N_VPWR_c_836_n N_A_861_368#_c_958_n 0.0250482f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_606 N_VPWR_c_847_n N_A_861_368#_c_959_n 0.042054f $X=8.695 $Y=3.33 $X2=0
+ $Y2=0
cc_607 N_VPWR_c_836_n N_A_861_368#_c_959_n 0.0235443f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_608 N_VPWR_c_839_n N_A_861_368#_c_960_n 0.0119251f $X=8.86 $Y=2.455 $X2=0
+ $Y2=0
cc_609 N_VPWR_c_847_n N_A_861_368#_c_960_n 0.0658009f $X=8.695 $Y=3.33 $X2=0
+ $Y2=0
cc_610 N_VPWR_c_836_n N_A_861_368#_c_960_n 0.036511f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_611 N_VPWR_c_839_n N_A_861_368#_c_961_n 0.0405754f $X=8.86 $Y=2.455 $X2=0
+ $Y2=0
cc_612 N_VPWR_c_847_n N_A_861_368#_c_962_n 0.0121867f $X=8.695 $Y=3.33 $X2=0
+ $Y2=0
cc_613 N_VPWR_c_836_n N_A_861_368#_c_962_n 0.00660921f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_614 N_VPWR_c_847_n N_A_861_368#_c_963_n 0.0229398f $X=8.695 $Y=3.33 $X2=0
+ $Y2=0
cc_615 N_VPWR_c_836_n N_A_861_368#_c_963_n 0.0124409f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_616 N_VPWR_c_847_n N_A_861_368#_c_964_n 0.0235512f $X=8.695 $Y=3.33 $X2=0
+ $Y2=0
cc_617 N_VPWR_c_836_n N_A_861_368#_c_964_n 0.0126924f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_618 N_VPWR_M1021_s N_A_1333_368#_c_1014_n 0.00543031f $X=8.715 $Y=1.84 $X2=0
+ $Y2=0
cc_619 N_VPWR_c_839_n N_A_1333_368#_c_1014_n 0.0197477f $X=8.86 $Y=2.455 $X2=0
+ $Y2=0
cc_620 N_VPWR_c_839_n N_A_1333_368#_c_1015_n 0.0234083f $X=8.86 $Y=2.455 $X2=0
+ $Y2=0
cc_621 N_VPWR_c_840_n N_A_1333_368#_c_1015_n 0.0266809f $X=9.81 $Y=2.455 $X2=0
+ $Y2=0
cc_622 N_VPWR_c_849_n N_A_1333_368#_c_1015_n 0.0144623f $X=9.645 $Y=3.33 $X2=0
+ $Y2=0
cc_623 N_VPWR_c_836_n N_A_1333_368#_c_1015_n 0.0118344f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_624 N_VPWR_M1024_s N_A_1333_368#_c_1038_n 0.00516882f $X=9.625 $Y=1.84 $X2=0
+ $Y2=0
cc_625 N_VPWR_c_840_n N_A_1333_368#_c_1038_n 0.0208278f $X=9.81 $Y=2.455 $X2=0
+ $Y2=0
cc_626 N_VPWR_c_840_n N_A_1333_368#_c_1016_n 0.0266809f $X=9.81 $Y=2.455 $X2=0
+ $Y2=0
cc_627 N_VPWR_c_842_n N_A_1333_368#_c_1016_n 0.0289761f $X=10.76 $Y=2.115 $X2=0
+ $Y2=0
cc_628 N_VPWR_c_850_n N_A_1333_368#_c_1016_n 0.0144623f $X=10.675 $Y=3.33 $X2=0
+ $Y2=0
cc_629 N_VPWR_c_836_n N_A_1333_368#_c_1016_n 0.0118344f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_630 N_A_861_368#_c_959_n N_A_1333_368#_M1003_d 0.00165831f $X=7.135 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_631 N_A_861_368#_c_960_n N_A_1333_368#_M1009_d 0.00218982f $X=8.135 $Y=2.99
+ $X2=0 $Y2=0
cc_632 N_A_861_368#_M1007_s N_A_1333_368#_c_1017_n 0.00410979f $X=7.115 $Y=1.84
+ $X2=0 $Y2=0
cc_633 N_A_861_368#_c_973_n N_A_1333_368#_c_1017_n 0.0189268f $X=7.3 $Y=2.455
+ $X2=0 $Y2=0
cc_634 N_A_861_368#_M1010_s N_A_1333_368#_c_1014_n 0.00682663f $X=8.115 $Y=1.84
+ $X2=0 $Y2=0
cc_635 N_A_861_368#_c_961_n N_A_1333_368#_c_1014_n 0.0238156f $X=8.3 $Y=2.455
+ $X2=0 $Y2=0
cc_636 N_A_861_368#_c_959_n N_A_1333_368#_c_1024_n 0.0159318f $X=7.135 $Y=2.99
+ $X2=0 $Y2=0
cc_637 N_A_861_368#_c_960_n N_A_1333_368#_c_1029_n 0.0177084f $X=8.135 $Y=2.99
+ $X2=0 $Y2=0
cc_638 N_A_27_74#_c_1117_n N_VGND_M1001_s 0.00724158f $X=4.995 $Y=0.835
+ $X2=-0.19 $Y2=-0.245
cc_639 N_A_27_74#_c_1123_n N_VGND_M1036_s 0.00345243f $X=5.995 $Y=0.835 $X2=0
+ $Y2=0
cc_640 N_A_27_74#_c_1080_n N_VGND_M1005_d 0.00358162f $X=7.34 $Y=1.095 $X2=0
+ $Y2=0
cc_641 N_A_27_74#_c_1082_n N_VGND_M1017_d 0.00358162f $X=8.34 $Y=1.095 $X2=0
+ $Y2=0
cc_642 N_A_27_74#_c_1084_n N_VGND_M1002_d 0.00250873f $X=9.34 $Y=1.095 $X2=0
+ $Y2=0
cc_643 N_A_27_74#_c_1086_n N_VGND_M1027_d 0.00250873f $X=10.34 $Y=1.095 $X2=0
+ $Y2=0
cc_644 N_A_27_74#_c_1078_n N_VGND_c_1257_n 0.0114117f $X=3.975 $Y=0.34 $X2=0
+ $Y2=0
cc_645 N_A_27_74#_c_1117_n N_VGND_c_1257_n 0.0256608f $X=4.995 $Y=0.835 $X2=0
+ $Y2=0
cc_646 N_A_27_74#_c_1079_n N_VGND_c_1257_n 0.0105187f $X=5.16 $Y=0.495 $X2=0
+ $Y2=0
cc_647 N_A_27_74#_c_1117_n N_VGND_c_1258_n 0.00197156f $X=4.995 $Y=0.835 $X2=0
+ $Y2=0
cc_648 N_A_27_74#_c_1079_n N_VGND_c_1258_n 0.0156726f $X=5.16 $Y=0.495 $X2=0
+ $Y2=0
cc_649 N_A_27_74#_c_1123_n N_VGND_c_1258_n 0.00193113f $X=5.995 $Y=0.835 $X2=0
+ $Y2=0
cc_650 N_A_27_74#_c_1079_n N_VGND_c_1259_n 0.0110032f $X=5.16 $Y=0.495 $X2=0
+ $Y2=0
cc_651 N_A_27_74#_c_1123_n N_VGND_c_1259_n 0.0165453f $X=5.995 $Y=0.835 $X2=0
+ $Y2=0
cc_652 N_A_27_74#_c_1091_n N_VGND_c_1259_n 0.0112413f $X=6.505 $Y=0.9 $X2=0
+ $Y2=0
cc_653 N_A_27_74#_c_1080_n N_VGND_c_1260_n 0.0248957f $X=7.34 $Y=1.095 $X2=0
+ $Y2=0
cc_654 N_A_27_74#_c_1081_n N_VGND_c_1260_n 0.0191765f $X=7.505 $Y=0.515 $X2=0
+ $Y2=0
cc_655 N_A_27_74#_c_1091_n N_VGND_c_1260_n 0.0230929f $X=6.505 $Y=0.9 $X2=0
+ $Y2=0
cc_656 N_A_27_74#_c_1081_n N_VGND_c_1261_n 0.0144922f $X=7.505 $Y=0.515 $X2=0
+ $Y2=0
cc_657 N_A_27_74#_c_1081_n N_VGND_c_1262_n 0.0191765f $X=7.505 $Y=0.515 $X2=0
+ $Y2=0
cc_658 N_A_27_74#_c_1082_n N_VGND_c_1262_n 0.0248957f $X=8.34 $Y=1.095 $X2=0
+ $Y2=0
cc_659 N_A_27_74#_c_1083_n N_VGND_c_1262_n 0.0191765f $X=8.505 $Y=0.515 $X2=0
+ $Y2=0
cc_660 N_A_27_74#_c_1083_n N_VGND_c_1263_n 0.0145639f $X=8.505 $Y=0.515 $X2=0
+ $Y2=0
cc_661 N_A_27_74#_c_1083_n N_VGND_c_1264_n 0.0191765f $X=8.505 $Y=0.515 $X2=0
+ $Y2=0
cc_662 N_A_27_74#_c_1084_n N_VGND_c_1264_n 0.0210288f $X=9.34 $Y=1.095 $X2=0
+ $Y2=0
cc_663 N_A_27_74#_c_1085_n N_VGND_c_1264_n 0.0191765f $X=9.505 $Y=0.515 $X2=0
+ $Y2=0
cc_664 N_A_27_74#_c_1085_n N_VGND_c_1265_n 0.0144922f $X=9.505 $Y=0.515 $X2=0
+ $Y2=0
cc_665 N_A_27_74#_c_1085_n N_VGND_c_1266_n 0.0191765f $X=9.505 $Y=0.515 $X2=0
+ $Y2=0
cc_666 N_A_27_74#_c_1086_n N_VGND_c_1266_n 0.0210288f $X=10.34 $Y=1.095 $X2=0
+ $Y2=0
cc_667 N_A_27_74#_c_1087_n N_VGND_c_1266_n 0.0191765f $X=10.505 $Y=0.515 $X2=0
+ $Y2=0
cc_668 N_A_27_74#_c_1074_n N_VGND_c_1267_n 0.0428729f $X=1.045 $Y=0.34 $X2=0
+ $Y2=0
cc_669 N_A_27_74#_c_1075_n N_VGND_c_1267_n 0.0179217f $X=0.365 $Y=0.34 $X2=0
+ $Y2=0
cc_670 N_A_27_74#_c_1076_n N_VGND_c_1267_n 0.0377951f $X=1.975 $Y=0.34 $X2=0
+ $Y2=0
cc_671 N_A_27_74#_c_1077_n N_VGND_c_1267_n 0.0423044f $X=2.975 $Y=0.34 $X2=0
+ $Y2=0
cc_672 N_A_27_74#_c_1078_n N_VGND_c_1267_n 0.0658334f $X=3.975 $Y=0.34 $X2=0
+ $Y2=0
cc_673 N_A_27_74#_c_1117_n N_VGND_c_1267_n 0.00197156f $X=4.995 $Y=0.835 $X2=0
+ $Y2=0
cc_674 N_A_27_74#_c_1088_n N_VGND_c_1267_n 0.0235293f $X=1.21 $Y=0.34 $X2=0
+ $Y2=0
cc_675 N_A_27_74#_c_1089_n N_VGND_c_1267_n 0.0235293f $X=2.14 $Y=0.34 $X2=0
+ $Y2=0
cc_676 N_A_27_74#_c_1090_n N_VGND_c_1267_n 0.0235293f $X=3.14 $Y=0.34 $X2=0
+ $Y2=0
cc_677 N_A_27_74#_c_1123_n N_VGND_c_1268_n 0.00190416f $X=5.995 $Y=0.835 $X2=0
+ $Y2=0
cc_678 N_A_27_74#_c_1091_n N_VGND_c_1268_n 0.032496f $X=6.505 $Y=0.9 $X2=0 $Y2=0
cc_679 N_A_27_74#_c_1087_n N_VGND_c_1269_n 0.0146357f $X=10.505 $Y=0.515 $X2=0
+ $Y2=0
cc_680 N_A_27_74#_c_1074_n N_VGND_c_1270_n 0.0241933f $X=1.045 $Y=0.34 $X2=0
+ $Y2=0
cc_681 N_A_27_74#_c_1075_n N_VGND_c_1270_n 0.00971942f $X=0.365 $Y=0.34 $X2=0
+ $Y2=0
cc_682 N_A_27_74#_c_1076_n N_VGND_c_1270_n 0.0212998f $X=1.975 $Y=0.34 $X2=0
+ $Y2=0
cc_683 N_A_27_74#_c_1077_n N_VGND_c_1270_n 0.0239316f $X=2.975 $Y=0.34 $X2=0
+ $Y2=0
cc_684 N_A_27_74#_c_1078_n N_VGND_c_1270_n 0.0366393f $X=3.975 $Y=0.34 $X2=0
+ $Y2=0
cc_685 N_A_27_74#_c_1117_n N_VGND_c_1270_n 0.00943478f $X=4.995 $Y=0.835 $X2=0
+ $Y2=0
cc_686 N_A_27_74#_c_1079_n N_VGND_c_1270_n 0.0120869f $X=5.16 $Y=0.495 $X2=0
+ $Y2=0
cc_687 N_A_27_74#_c_1123_n N_VGND_c_1270_n 0.00885587f $X=5.995 $Y=0.835 $X2=0
+ $Y2=0
cc_688 N_A_27_74#_c_1081_n N_VGND_c_1270_n 0.0118826f $X=7.505 $Y=0.515 $X2=0
+ $Y2=0
cc_689 N_A_27_74#_c_1083_n N_VGND_c_1270_n 0.0119984f $X=8.505 $Y=0.515 $X2=0
+ $Y2=0
cc_690 N_A_27_74#_c_1085_n N_VGND_c_1270_n 0.0118826f $X=9.505 $Y=0.515 $X2=0
+ $Y2=0
cc_691 N_A_27_74#_c_1087_n N_VGND_c_1270_n 0.0121141f $X=10.505 $Y=0.515 $X2=0
+ $Y2=0
cc_692 N_A_27_74#_c_1088_n N_VGND_c_1270_n 0.0127078f $X=1.21 $Y=0.34 $X2=0
+ $Y2=0
cc_693 N_A_27_74#_c_1089_n N_VGND_c_1270_n 0.0127078f $X=2.14 $Y=0.34 $X2=0
+ $Y2=0
cc_694 N_A_27_74#_c_1090_n N_VGND_c_1270_n 0.0127078f $X=3.14 $Y=0.34 $X2=0
+ $Y2=0
cc_695 N_A_27_74#_c_1091_n N_VGND_c_1270_n 0.0250488f $X=6.505 $Y=0.9 $X2=0
+ $Y2=0

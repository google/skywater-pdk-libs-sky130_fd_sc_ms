* NGSPICE file created from sky130_fd_sc_ms__a222oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__a222oi_1 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR Y
M1000 VGND C2 a_119_74# VNB nlowvt w=640000u l=150000u
+  ad=9.312e+11p pd=5.47e+06u as=1.536e+11p ps=1.76e+06u
M1001 a_119_392# C1 Y VPB pshort w=1e+06u l=180000u
+  ad=6.4e+11p pd=5.28e+06u as=6.1e+11p ps=5.22e+06u
M1002 a_461_74# B2 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1003 a_119_74# C1 Y VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=5.92e+11p ps=4.41e+06u
M1004 Y B1 a_461_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A2 a_697_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.536e+11p ps=1.76e+06u
M1006 a_697_74# A1 Y VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_369_392# A2 VPWR VPB pshort w=1e+06u l=180000u
+  ad=8.8e+11p pd=7.76e+06u as=4.2e+11p ps=2.84e+06u
M1008 VPWR A1 a_369_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_119_392# B2 a_369_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_369_392# B1 a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y C2 a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


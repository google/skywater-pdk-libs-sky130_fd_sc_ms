* File: sky130_fd_sc_ms__a31o_1.pxi.spice
* Created: Wed Sep  2 11:55:01 2020
* 
x_PM_SKY130_FD_SC_MS__A31O_1%A_81_270# N_A_81_270#_M1009_d N_A_81_270#_M1002_d
+ N_A_81_270#_M1007_g N_A_81_270#_M1006_g N_A_81_270#_c_60_n N_A_81_270#_c_97_p
+ N_A_81_270#_c_61_n N_A_81_270#_c_62_n N_A_81_270#_c_63_n N_A_81_270#_c_64_n
+ N_A_81_270#_c_65_n N_A_81_270#_c_66_n PM_SKY130_FD_SC_MS__A31O_1%A_81_270#
x_PM_SKY130_FD_SC_MS__A31O_1%A3 N_A3_M1003_g N_A3_M1008_g A3 N_A3_c_138_n
+ PM_SKY130_FD_SC_MS__A31O_1%A3
x_PM_SKY130_FD_SC_MS__A31O_1%A2 N_A2_M1005_g N_A2_M1004_g A2 N_A2_c_176_n
+ PM_SKY130_FD_SC_MS__A31O_1%A2
x_PM_SKY130_FD_SC_MS__A31O_1%A1 N_A1_M1009_g N_A1_M1001_g A1 N_A1_c_211_n
+ PM_SKY130_FD_SC_MS__A31O_1%A1
x_PM_SKY130_FD_SC_MS__A31O_1%B1 N_B1_M1002_g N_B1_M1000_g N_B1_c_248_n B1 B1 B1
+ N_B1_c_249_n N_B1_c_250_n PM_SKY130_FD_SC_MS__A31O_1%B1
x_PM_SKY130_FD_SC_MS__A31O_1%X N_X_M1006_s N_X_M1007_s N_X_c_285_n N_X_c_286_n X
+ X X X N_X_c_287_n PM_SKY130_FD_SC_MS__A31O_1%X
x_PM_SKY130_FD_SC_MS__A31O_1%VPWR N_VPWR_M1007_d N_VPWR_M1004_d N_VPWR_c_308_n
+ N_VPWR_c_309_n N_VPWR_c_310_n N_VPWR_c_311_n VPWR N_VPWR_c_312_n
+ N_VPWR_c_313_n N_VPWR_c_307_n N_VPWR_c_315_n PM_SKY130_FD_SC_MS__A31O_1%VPWR
x_PM_SKY130_FD_SC_MS__A31O_1%A_253_392# N_A_253_392#_M1003_d
+ N_A_253_392#_M1001_d N_A_253_392#_c_351_n N_A_253_392#_c_349_n
+ N_A_253_392#_c_352_n N_A_253_392#_c_353_n N_A_253_392#_c_350_n
+ PM_SKY130_FD_SC_MS__A31O_1%A_253_392#
x_PM_SKY130_FD_SC_MS__A31O_1%VGND N_VGND_M1006_d N_VGND_M1000_d N_VGND_c_386_n
+ N_VGND_c_387_n N_VGND_c_388_n N_VGND_c_389_n VGND N_VGND_c_390_n
+ N_VGND_c_391_n N_VGND_c_392_n N_VGND_c_393_n PM_SKY130_FD_SC_MS__A31O_1%VGND
cc_1 VNB N_A_81_270#_c_60_n 0.0121926f $X=-0.19 $Y=-0.245 $X2=2.28 $Y2=1.235
cc_2 VNB N_A_81_270#_c_61_n 0.0088318f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=1.235
cc_3 VNB N_A_81_270#_c_62_n 0.0173236f $X=-0.19 $Y=-0.245 $X2=2.93 $Y2=2.105
cc_4 VNB N_A_81_270#_c_63_n 0.00531266f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.235
cc_5 VNB N_A_81_270#_c_64_n 0.0289898f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.515
cc_6 VNB N_A_81_270#_c_65_n 0.00437417f $X=-0.19 $Y=-0.245 $X2=2.445 $Y2=1.235
cc_7 VNB N_A_81_270#_c_66_n 0.0221308f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.35
cc_8 VNB N_A3_M1008_g 0.0237957f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.68
cc_9 VNB A3 0.0021755f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_10 VNB N_A3_c_138_n 0.0155404f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.87
cc_11 VNB N_A2_M1005_g 0.0226062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_c_176_n 0.0173271f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.87
cc_13 VNB N_A1_M1009_g 0.0235943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB A1 0.00279888f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_15 VNB N_A1_c_211_n 0.0153346f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.87
cc_16 VNB N_B1_M1002_g 0.0042235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B1_M1000_g 0.0179075f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_18 VNB N_B1_c_248_n 0.0115349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_c_249_n 0.0473693f $X=-0.19 $Y=-0.245 $X2=2.445 $Y2=0.955
cc_20 VNB N_B1_c_250_n 0.0142364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_X_c_285_n 0.0248845f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_22 VNB N_X_c_286_n 0.00743257f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.87
cc_23 VNB N_X_c_287_n 0.0221277f $X=-0.19 $Y=-0.245 $X2=2.445 $Y2=1.235
cc_24 VNB N_VPWR_c_307_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_386_n 0.0209501f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.4
cc_26 VNB N_VGND_c_387_n 0.0120067f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.35
cc_27 VNB N_VGND_c_388_n 0.0295961f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.87
cc_28 VNB N_VGND_c_389_n 0.00921063f $X=-0.19 $Y=-0.245 $X2=2.445 $Y2=1.15
cc_29 VNB N_VGND_c_390_n 0.0196766f $X=-0.19 $Y=-0.245 $X2=2.845 $Y2=1.235
cc_30 VNB N_VGND_c_391_n 0.0448011f $X=-0.19 $Y=-0.245 $X2=2.97 $Y2=2.815
cc_31 VNB N_VGND_c_392_n 0.0111562f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.35
cc_32 VNB N_VGND_c_393_n 0.219881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VPB N_A_81_270#_M1007_g 0.029133f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_34 VPB N_A_81_270#_c_62_n 0.0568125f $X=-0.19 $Y=1.66 $X2=2.93 $Y2=2.105
cc_35 VPB N_A_81_270#_c_63_n 0.00341417f $X=-0.19 $Y=1.66 $X2=0.625 $Y2=1.235
cc_36 VPB N_A_81_270#_c_64_n 0.0063159f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.515
cc_37 VPB N_A3_M1003_g 0.02445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB A3 0.00256767f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_39 VPB N_A3_c_138_n 0.0129815f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.87
cc_40 VPB N_A2_M1004_g 0.0240563f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.68
cc_41 VPB A2 0.00138051f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_42 VPB N_A2_c_176_n 0.0137752f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.87
cc_43 VPB N_A1_M1001_g 0.0240551f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.68
cc_44 VPB A1 0.00235147f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_45 VPB N_A1_c_211_n 0.0115364f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=0.87
cc_46 VPB N_B1_M1002_g 0.0340492f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB X 0.00695105f $X=-0.19 $Y=1.66 $X2=2.28 $Y2=1.235
cc_48 VPB X 0.0406888f $X=-0.19 $Y=1.66 $X2=2.97 $Y2=2.105
cc_49 VPB N_X_c_287_n 0.00901974f $X=-0.19 $Y=1.66 $X2=2.445 $Y2=1.235
cc_50 VPB N_VPWR_c_308_n 0.0104132f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_51 VPB N_VPWR_c_309_n 0.00987068f $X=-0.19 $Y=1.66 $X2=0.825 $Y2=1.235
cc_52 VPB N_VPWR_c_310_n 0.0186948f $X=-0.19 $Y=1.66 $X2=2.445 $Y2=0.955
cc_53 VPB N_VPWR_c_311_n 0.00786036f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_312_n 0.018677f $X=-0.19 $Y=1.66 $X2=2.97 $Y2=1.32
cc_55 VPB N_VPWR_c_313_n 0.0363074f $X=-0.19 $Y=1.66 $X2=0.58 $Y2=1.68
cc_56 VPB N_VPWR_c_307_n 0.0643112f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_315_n 0.0088221f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_A_253_392#_c_349_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.4
cc_59 VPB N_A_253_392#_c_350_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.825 $Y2=1.235
cc_60 N_A_81_270#_M1007_g N_A3_M1003_g 0.021138f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_61 N_A_81_270#_c_60_n N_A3_M1008_g 0.0149586f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_62 N_A_81_270#_c_63_n N_A3_M1008_g 0.00309045f $X=0.625 $Y=1.235 $X2=0 $Y2=0
cc_63 N_A_81_270#_c_64_n N_A3_M1008_g 0.00287123f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_64 N_A_81_270#_c_66_n N_A3_M1008_g 0.00806675f $X=0.58 $Y=1.35 $X2=0 $Y2=0
cc_65 N_A_81_270#_M1007_g A3 6.91928e-19 $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_66 N_A_81_270#_c_60_n A3 0.0241217f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_67 N_A_81_270#_c_63_n A3 0.0153381f $X=0.625 $Y=1.235 $X2=0 $Y2=0
cc_68 N_A_81_270#_c_64_n A3 2.0879e-19 $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_69 N_A_81_270#_M1007_g N_A3_c_138_n 0.00308451f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_70 N_A_81_270#_c_60_n N_A3_c_138_n 0.00449386f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_71 N_A_81_270#_c_63_n N_A3_c_138_n 0.00117732f $X=0.625 $Y=1.235 $X2=0 $Y2=0
cc_72 N_A_81_270#_c_64_n N_A3_c_138_n 0.0115055f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_73 N_A_81_270#_c_60_n N_A2_M1005_g 0.0127685f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_74 N_A_81_270#_c_60_n A2 0.024098f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_75 N_A_81_270#_c_60_n N_A2_c_176_n 0.00425501f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_76 N_A_81_270#_c_60_n N_A1_M1009_g 0.0134426f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_77 N_A_81_270#_c_60_n A1 0.0171013f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_78 N_A_81_270#_c_62_n A1 0.0117728f $X=2.93 $Y=2.105 $X2=0 $Y2=0
cc_79 N_A_81_270#_c_65_n A1 0.0102517f $X=2.445 $Y=1.235 $X2=0 $Y2=0
cc_80 N_A_81_270#_c_60_n N_A1_c_211_n 0.00148156f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_81 N_A_81_270#_c_65_n N_A1_c_211_n 0.00321516f $X=2.445 $Y=1.235 $X2=0 $Y2=0
cc_82 N_A_81_270#_c_62_n N_B1_M1002_g 0.0129369f $X=2.93 $Y=2.105 $X2=0 $Y2=0
cc_83 N_A_81_270#_c_61_n N_B1_M1000_g 0.0184507f $X=2.845 $Y=1.235 $X2=0 $Y2=0
cc_84 N_A_81_270#_c_62_n N_B1_M1000_g 0.00983966f $X=2.93 $Y=2.105 $X2=0 $Y2=0
cc_85 N_A_81_270#_c_61_n N_B1_c_248_n 0.00188154f $X=2.845 $Y=1.235 $X2=0 $Y2=0
cc_86 N_A_81_270#_c_97_p N_B1_c_249_n 6.83819e-19 $X=2.445 $Y=0.955 $X2=0 $Y2=0
cc_87 N_A_81_270#_M1009_d N_B1_c_250_n 0.00355368f $X=2.225 $Y=0.615 $X2=0 $Y2=0
cc_88 N_A_81_270#_c_60_n N_B1_c_250_n 0.0174185f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_89 N_A_81_270#_c_97_p N_B1_c_250_n 0.0266869f $X=2.445 $Y=0.955 $X2=0 $Y2=0
cc_90 N_A_81_270#_c_61_n N_B1_c_250_n 0.00368593f $X=2.845 $Y=1.235 $X2=0 $Y2=0
cc_91 N_A_81_270#_c_66_n N_X_c_285_n 0.00629257f $X=0.58 $Y=1.35 $X2=0 $Y2=0
cc_92 N_A_81_270#_c_63_n N_X_c_286_n 0.00146264f $X=0.625 $Y=1.235 $X2=0 $Y2=0
cc_93 N_A_81_270#_c_66_n N_X_c_286_n 0.00702486f $X=0.58 $Y=1.35 $X2=0 $Y2=0
cc_94 N_A_81_270#_M1007_g X 0.00397838f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_95 N_A_81_270#_c_63_n X 7.22171e-19 $X=0.625 $Y=1.235 $X2=0 $Y2=0
cc_96 N_A_81_270#_M1007_g X 0.0120548f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_97 N_A_81_270#_c_63_n N_X_c_287_n 0.0307829f $X=0.625 $Y=1.235 $X2=0 $Y2=0
cc_98 N_A_81_270#_c_64_n N_X_c_287_n 0.0119308f $X=0.59 $Y=1.515 $X2=0 $Y2=0
cc_99 N_A_81_270#_c_66_n N_X_c_287_n 0.00249972f $X=0.58 $Y=1.35 $X2=0 $Y2=0
cc_100 N_A_81_270#_M1007_g N_VPWR_c_308_n 0.0114459f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_101 N_A_81_270#_c_60_n N_VPWR_c_308_n 0.00527561f $X=2.28 $Y=1.235 $X2=0
+ $Y2=0
cc_102 N_A_81_270#_c_63_n N_VPWR_c_308_n 0.011642f $X=0.625 $Y=1.235 $X2=0 $Y2=0
cc_103 N_A_81_270#_c_64_n N_VPWR_c_308_n 9.63158e-19 $X=0.59 $Y=1.515 $X2=0
+ $Y2=0
cc_104 N_A_81_270#_M1007_g N_VPWR_c_312_n 0.005209f $X=0.495 $Y=2.4 $X2=0 $Y2=0
cc_105 N_A_81_270#_c_62_n N_VPWR_c_313_n 0.011066f $X=2.93 $Y=2.105 $X2=0 $Y2=0
cc_106 N_A_81_270#_M1007_g N_VPWR_c_307_n 0.00987203f $X=0.495 $Y=2.4 $X2=0
+ $Y2=0
cc_107 N_A_81_270#_c_62_n N_VPWR_c_307_n 0.00915947f $X=2.93 $Y=2.105 $X2=0
+ $Y2=0
cc_108 N_A_81_270#_c_60_n N_A_253_392#_c_351_n 0.00561552f $X=2.28 $Y=1.235
+ $X2=0 $Y2=0
cc_109 N_A_81_270#_c_60_n N_A_253_392#_c_352_n 0.00507286f $X=2.28 $Y=1.235
+ $X2=0 $Y2=0
cc_110 N_A_81_270#_c_61_n N_A_253_392#_c_353_n 8.93138e-19 $X=2.845 $Y=1.235
+ $X2=0 $Y2=0
cc_111 N_A_81_270#_c_65_n N_A_253_392#_c_353_n 0.00608946f $X=2.445 $Y=1.235
+ $X2=0 $Y2=0
cc_112 N_A_81_270#_c_62_n N_A_253_392#_c_350_n 0.0283172f $X=2.93 $Y=2.105 $X2=0
+ $Y2=0
cc_113 N_A_81_270#_c_60_n N_VGND_M1006_d 0.00351422f $X=2.28 $Y=1.235 $X2=-0.19
+ $Y2=-0.245
cc_114 N_A_81_270#_c_63_n N_VGND_M1006_d 0.00221237f $X=0.625 $Y=1.235 $X2=-0.19
+ $Y2=-0.245
cc_115 N_A_81_270#_c_61_n N_VGND_M1000_d 0.00280144f $X=2.845 $Y=1.235 $X2=0
+ $Y2=0
cc_116 N_A_81_270#_c_60_n N_VGND_c_386_n 0.0255877f $X=2.28 $Y=1.235 $X2=0 $Y2=0
cc_117 N_A_81_270#_c_63_n N_VGND_c_386_n 0.0162002f $X=0.625 $Y=1.235 $X2=0
+ $Y2=0
cc_118 N_A_81_270#_c_64_n N_VGND_c_386_n 6.25171e-19 $X=0.59 $Y=1.515 $X2=0
+ $Y2=0
cc_119 N_A_81_270#_c_66_n N_VGND_c_386_n 0.00650193f $X=0.58 $Y=1.35 $X2=0 $Y2=0
cc_120 N_A_81_270#_c_61_n N_VGND_c_389_n 0.0198501f $X=2.845 $Y=1.235 $X2=0
+ $Y2=0
cc_121 N_A_81_270#_c_66_n N_VGND_c_390_n 0.00475875f $X=0.58 $Y=1.35 $X2=0 $Y2=0
cc_122 N_A_81_270#_c_66_n N_VGND_c_393_n 0.00505379f $X=0.58 $Y=1.35 $X2=0 $Y2=0
cc_123 N_A_81_270#_c_60_n A_265_120# 0.00366293f $X=2.28 $Y=1.235 $X2=-0.19
+ $Y2=-0.245
cc_124 N_A_81_270#_c_60_n A_337_120# 0.00521091f $X=2.28 $Y=1.235 $X2=-0.19
+ $Y2=-0.245
cc_125 N_A3_M1008_g N_A2_M1005_g 0.0416465f $X=1.25 $Y=0.92 $X2=0 $Y2=0
cc_126 N_A3_M1003_g N_A2_M1004_g 0.0144965f $X=1.175 $Y=2.46 $X2=0 $Y2=0
cc_127 A3 A2 0.0196026f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_128 N_A3_c_138_n A2 3.89032e-19 $X=1.16 $Y=1.635 $X2=0 $Y2=0
cc_129 A3 N_A2_c_176_n 0.0010743f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_130 N_A3_c_138_n N_A2_c_176_n 0.0416465f $X=1.16 $Y=1.635 $X2=0 $Y2=0
cc_131 N_A3_M1008_g N_B1_c_250_n 5.34903e-19 $X=1.25 $Y=0.92 $X2=0 $Y2=0
cc_132 N_A3_M1003_g X 6.73872e-19 $X=1.175 $Y=2.46 $X2=0 $Y2=0
cc_133 N_A3_M1003_g N_VPWR_c_308_n 0.00994014f $X=1.175 $Y=2.46 $X2=0 $Y2=0
cc_134 A3 N_VPWR_c_308_n 0.00405759f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_135 N_A3_c_138_n N_VPWR_c_308_n 0.0014977f $X=1.16 $Y=1.635 $X2=0 $Y2=0
cc_136 N_A3_M1003_g N_VPWR_c_310_n 0.005209f $X=1.175 $Y=2.46 $X2=0 $Y2=0
cc_137 N_A3_M1003_g N_VPWR_c_307_n 0.00983608f $X=1.175 $Y=2.46 $X2=0 $Y2=0
cc_138 N_A3_M1003_g N_A_253_392#_c_351_n 0.00238276f $X=1.175 $Y=2.46 $X2=0
+ $Y2=0
cc_139 A3 N_A_253_392#_c_351_n 0.00471696f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_140 N_A3_c_138_n N_A_253_392#_c_351_n 0.00146071f $X=1.16 $Y=1.635 $X2=0
+ $Y2=0
cc_141 N_A3_M1003_g N_A_253_392#_c_349_n 0.01015f $X=1.175 $Y=2.46 $X2=0 $Y2=0
cc_142 N_A3_M1008_g N_VGND_c_386_n 0.013823f $X=1.25 $Y=0.92 $X2=0 $Y2=0
cc_143 N_A3_M1008_g N_VGND_c_391_n 0.00356352f $X=1.25 $Y=0.92 $X2=0 $Y2=0
cc_144 N_A3_M1008_g N_VGND_c_393_n 0.00400172f $X=1.25 $Y=0.92 $X2=0 $Y2=0
cc_145 N_A2_M1005_g N_A1_M1009_g 0.0326149f $X=1.61 $Y=0.92 $X2=0 $Y2=0
cc_146 N_A2_M1004_g N_A1_M1001_g 0.0274079f $X=1.625 $Y=2.46 $X2=0 $Y2=0
cc_147 A2 A1 0.0236226f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_148 N_A2_c_176_n A1 0.00175997f $X=1.7 $Y=1.635 $X2=0 $Y2=0
cc_149 A2 N_A1_c_211_n 3.63175e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_150 N_A2_c_176_n N_A1_c_211_n 0.0209153f $X=1.7 $Y=1.635 $X2=0 $Y2=0
cc_151 N_A2_M1005_g N_B1_c_250_n 0.0115129f $X=1.61 $Y=0.92 $X2=0 $Y2=0
cc_152 N_A2_M1004_g N_VPWR_c_309_n 0.00681871f $X=1.625 $Y=2.46 $X2=0 $Y2=0
cc_153 N_A2_M1004_g N_VPWR_c_310_n 0.005209f $X=1.625 $Y=2.46 $X2=0 $Y2=0
cc_154 N_A2_M1004_g N_VPWR_c_307_n 0.00983279f $X=1.625 $Y=2.46 $X2=0 $Y2=0
cc_155 N_A2_M1004_g N_A_253_392#_c_351_n 8.8334e-19 $X=1.625 $Y=2.46 $X2=0 $Y2=0
cc_156 A2 N_A_253_392#_c_351_n 0.00231658f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_157 N_A2_M1004_g N_A_253_392#_c_349_n 0.0118578f $X=1.625 $Y=2.46 $X2=0 $Y2=0
cc_158 N_A2_M1004_g N_A_253_392#_c_352_n 0.0137624f $X=1.625 $Y=2.46 $X2=0 $Y2=0
cc_159 A2 N_A_253_392#_c_352_n 0.0196054f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_160 N_A2_c_176_n N_A_253_392#_c_352_n 9.26001e-19 $X=1.7 $Y=1.635 $X2=0 $Y2=0
cc_161 N_A2_M1004_g N_A_253_392#_c_350_n 8.65935e-19 $X=1.625 $Y=2.46 $X2=0
+ $Y2=0
cc_162 N_A2_M1005_g N_VGND_c_386_n 0.00212757f $X=1.61 $Y=0.92 $X2=0 $Y2=0
cc_163 N_A2_M1005_g N_VGND_c_391_n 0.0013085f $X=1.61 $Y=0.92 $X2=0 $Y2=0
cc_164 N_A2_M1005_g N_VGND_c_393_n 9.5279e-19 $X=1.61 $Y=0.92 $X2=0 $Y2=0
cc_165 N_A1_M1001_g N_B1_M1002_g 0.014321f $X=2.255 $Y=2.46 $X2=0 $Y2=0
cc_166 N_A1_M1009_g N_B1_M1000_g 0.0223483f $X=2.15 $Y=0.935 $X2=0 $Y2=0
cc_167 N_A1_M1009_g N_B1_c_248_n 0.00117875f $X=2.15 $Y=0.935 $X2=0 $Y2=0
cc_168 A1 N_B1_c_248_n 0.00114373f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_169 N_A1_c_211_n N_B1_c_248_n 0.0200553f $X=2.24 $Y=1.635 $X2=0 $Y2=0
cc_170 N_A1_M1009_g N_B1_c_249_n 9.92136e-19 $X=2.15 $Y=0.935 $X2=0 $Y2=0
cc_171 N_A1_M1009_g N_B1_c_250_n 0.013629f $X=2.15 $Y=0.935 $X2=0 $Y2=0
cc_172 N_A1_M1001_g N_VPWR_c_309_n 0.00828598f $X=2.255 $Y=2.46 $X2=0 $Y2=0
cc_173 N_A1_M1001_g N_VPWR_c_313_n 0.005209f $X=2.255 $Y=2.46 $X2=0 $Y2=0
cc_174 N_A1_M1001_g N_VPWR_c_307_n 0.00983279f $X=2.255 $Y=2.46 $X2=0 $Y2=0
cc_175 N_A1_M1001_g N_A_253_392#_c_349_n 8.65935e-19 $X=2.255 $Y=2.46 $X2=0
+ $Y2=0
cc_176 N_A1_M1001_g N_A_253_392#_c_352_n 0.0137686f $X=2.255 $Y=2.46 $X2=0 $Y2=0
cc_177 A1 N_A_253_392#_c_352_n 0.0174944f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_178 N_A1_c_211_n N_A_253_392#_c_352_n 0.00224739f $X=2.24 $Y=1.635 $X2=0
+ $Y2=0
cc_179 N_A1_M1001_g N_A_253_392#_c_353_n 8.84614e-19 $X=2.255 $Y=2.46 $X2=0
+ $Y2=0
cc_180 A1 N_A_253_392#_c_353_n 0.00471696f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_181 N_A1_c_211_n N_A_253_392#_c_353_n 0.00122405f $X=2.24 $Y=1.635 $X2=0
+ $Y2=0
cc_182 N_A1_M1001_g N_A_253_392#_c_350_n 0.0118578f $X=2.255 $Y=2.46 $X2=0 $Y2=0
cc_183 N_A1_M1009_g N_VGND_c_391_n 5.46057e-19 $X=2.15 $Y=0.935 $X2=0 $Y2=0
cc_184 N_B1_M1002_g N_VPWR_c_313_n 0.005209f $X=2.705 $Y=2.46 $X2=0 $Y2=0
cc_185 N_B1_M1002_g N_VPWR_c_307_n 0.00987636f $X=2.705 $Y=2.46 $X2=0 $Y2=0
cc_186 N_B1_M1002_g N_A_253_392#_c_353_n 0.00288529f $X=2.705 $Y=2.46 $X2=0
+ $Y2=0
cc_187 N_B1_M1002_g N_A_253_392#_c_350_n 0.0110096f $X=2.705 $Y=2.46 $X2=0 $Y2=0
cc_188 N_B1_c_250_n N_VGND_c_386_n 0.0192005f $X=2.65 $Y=0.34 $X2=0 $Y2=0
cc_189 N_B1_M1000_g N_VGND_c_388_n 0.00399579f $X=2.74 $Y=0.935 $X2=0 $Y2=0
cc_190 N_B1_c_249_n N_VGND_c_388_n 0.00511411f $X=2.65 $Y=0.34 $X2=0 $Y2=0
cc_191 N_B1_c_250_n N_VGND_c_388_n 0.0305341f $X=2.65 $Y=0.34 $X2=0 $Y2=0
cc_192 N_B1_M1000_g N_VGND_c_389_n 0.00244045f $X=2.74 $Y=0.935 $X2=0 $Y2=0
cc_193 N_B1_c_250_n N_VGND_c_389_n 0.00172851f $X=2.65 $Y=0.34 $X2=0 $Y2=0
cc_194 N_B1_c_249_n N_VGND_c_391_n 0.00659816f $X=2.65 $Y=0.34 $X2=0 $Y2=0
cc_195 N_B1_c_250_n N_VGND_c_391_n 0.084256f $X=2.65 $Y=0.34 $X2=0 $Y2=0
cc_196 N_B1_c_249_n N_VGND_c_393_n 0.0102618f $X=2.65 $Y=0.34 $X2=0 $Y2=0
cc_197 N_B1_c_250_n N_VGND_c_393_n 0.0463662f $X=2.65 $Y=0.34 $X2=0 $Y2=0
cc_198 N_B1_c_250_n A_337_120# 0.00524643f $X=2.65 $Y=0.34 $X2=-0.19 $Y2=-0.245
cc_199 X N_VPWR_c_308_n 0.0390338f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_200 X N_VPWR_c_312_n 0.0154414f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_201 X N_VPWR_c_307_n 0.0127129f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_202 N_X_c_285_n N_VGND_c_386_n 0.0199137f $X=0.295 $Y=0.645 $X2=0 $Y2=0
cc_203 N_X_c_285_n N_VGND_c_390_n 0.0105642f $X=0.295 $Y=0.645 $X2=0 $Y2=0
cc_204 N_X_c_285_n N_VGND_c_393_n 0.0123086f $X=0.295 $Y=0.645 $X2=0 $Y2=0
cc_205 N_VPWR_c_308_n N_A_253_392#_c_349_n 0.0323124f $X=0.835 $Y=2.135 $X2=0
+ $Y2=0
cc_206 N_VPWR_c_309_n N_A_253_392#_c_349_n 0.0259568f $X=1.94 $Y=2.42 $X2=0
+ $Y2=0
cc_207 N_VPWR_c_310_n N_A_253_392#_c_349_n 0.0144623f $X=1.735 $Y=3.33 $X2=0
+ $Y2=0
cc_208 N_VPWR_c_307_n N_A_253_392#_c_349_n 0.0118344f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_209 N_VPWR_M1004_d N_A_253_392#_c_352_n 0.00948736f $X=1.715 $Y=1.96 $X2=0
+ $Y2=0
cc_210 N_VPWR_c_309_n N_A_253_392#_c_352_n 0.0273365f $X=1.94 $Y=2.42 $X2=0
+ $Y2=0
cc_211 N_VPWR_c_309_n N_A_253_392#_c_350_n 0.0259568f $X=1.94 $Y=2.42 $X2=0
+ $Y2=0
cc_212 N_VPWR_c_313_n N_A_253_392#_c_350_n 0.0144623f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_213 N_VPWR_c_307_n N_A_253_392#_c_350_n 0.0118344f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__sdfrtp_2.pxi.spice
* Created: Wed Sep  2 12:30:39 2020
* 
x_PM_SKY130_FD_SC_MS__SDFRTP_2%A_27_74# N_A_27_74#_M1036_s N_A_27_74#_M1011_s
+ N_A_27_74#_c_291_n N_A_27_74#_c_292_n N_A_27_74#_M1014_g N_A_27_74#_M1038_g
+ N_A_27_74#_c_293_n N_A_27_74#_c_294_n N_A_27_74#_c_300_n N_A_27_74#_c_295_n
+ N_A_27_74#_c_301_n N_A_27_74#_c_296_n N_A_27_74#_c_302_n N_A_27_74#_c_303_n
+ N_A_27_74#_c_304_n N_A_27_74#_c_297_n PM_SKY130_FD_SC_MS__SDFRTP_2%A_27_74#
x_PM_SKY130_FD_SC_MS__SDFRTP_2%SCE N_SCE_M1011_g N_SCE_M1036_g N_SCE_M1012_g
+ N_SCE_M1008_g N_SCE_c_375_n N_SCE_c_376_n N_SCE_c_377_n N_SCE_c_378_n
+ N_SCE_c_379_n N_SCE_c_380_n N_SCE_c_381_n SCE SCE SCE N_SCE_c_382_n
+ N_SCE_c_383_n SCE N_SCE_c_384_n PM_SKY130_FD_SC_MS__SDFRTP_2%SCE
x_PM_SKY130_FD_SC_MS__SDFRTP_2%D N_D_M1015_g N_D_M1000_g D N_D_c_460_n
+ N_D_c_461_n N_D_c_462_n PM_SKY130_FD_SC_MS__SDFRTP_2%D
x_PM_SKY130_FD_SC_MS__SDFRTP_2%SCD N_SCD_M1039_g N_SCD_M1035_g N_SCD_c_504_n
+ N_SCD_c_509_n SCD SCD N_SCD_c_506_n PM_SKY130_FD_SC_MS__SDFRTP_2%SCD
x_PM_SKY130_FD_SC_MS__SDFRTP_2%CLK N_CLK_c_551_n N_CLK_M1016_g N_CLK_M1027_g CLK
+ N_CLK_c_553_n N_CLK_c_554_n N_CLK_c_555_n PM_SKY130_FD_SC_MS__SDFRTP_2%CLK
x_PM_SKY130_FD_SC_MS__SDFRTP_2%A_1037_119# N_A_1037_119#_M1017_d
+ N_A_1037_119#_M1034_d N_A_1037_119#_M1002_g N_A_1037_119#_c_611_n
+ N_A_1037_119#_c_612_n N_A_1037_119#_M1032_g N_A_1037_119#_c_614_n
+ N_A_1037_119#_M1028_g N_A_1037_119#_c_615_n N_A_1037_119#_c_616_n
+ N_A_1037_119#_M1021_g N_A_1037_119#_c_617_n N_A_1037_119#_c_618_n
+ N_A_1037_119#_c_619_n N_A_1037_119#_c_620_n N_A_1037_119#_c_621_n
+ N_A_1037_119#_c_622_n N_A_1037_119#_c_803_p N_A_1037_119#_c_623_n
+ N_A_1037_119#_c_624_n N_A_1037_119#_c_684_p N_A_1037_119#_c_625_n
+ N_A_1037_119#_c_626_n N_A_1037_119#_c_627_n N_A_1037_119#_c_628_n
+ N_A_1037_119#_c_629_n N_A_1037_119#_c_630_n N_A_1037_119#_c_631_n
+ N_A_1037_119#_c_632_n N_A_1037_119#_c_641_n
+ PM_SKY130_FD_SC_MS__SDFRTP_2%A_1037_119#
x_PM_SKY130_FD_SC_MS__SDFRTP_2%A_1383_349# N_A_1383_349#_M1040_d
+ N_A_1383_349#_M1006_d N_A_1383_349#_M1033_g N_A_1383_349#_M1022_g
+ N_A_1383_349#_c_826_n N_A_1383_349#_c_833_n N_A_1383_349#_c_827_n
+ N_A_1383_349#_c_848_n N_A_1383_349#_c_834_n N_A_1383_349#_c_828_n
+ N_A_1383_349#_c_835_n N_A_1383_349#_c_829_n
+ PM_SKY130_FD_SC_MS__SDFRTP_2%A_1383_349#
x_PM_SKY130_FD_SC_MS__SDFRTP_2%RESET_B N_RESET_B_c_917_n N_RESET_B_M1023_g
+ N_RESET_B_M1004_g N_RESET_B_c_919_n N_RESET_B_c_920_n N_RESET_B_M1007_g
+ N_RESET_B_M1013_g N_RESET_B_c_922_n N_RESET_B_M1026_g N_RESET_B_M1019_g
+ N_RESET_B_c_924_n N_RESET_B_c_932_n N_RESET_B_c_925_n N_RESET_B_c_933_n
+ N_RESET_B_c_934_n N_RESET_B_c_935_n N_RESET_B_c_936_n N_RESET_B_c_937_n
+ RESET_B N_RESET_B_c_938_n N_RESET_B_c_939_n N_RESET_B_c_940_n
+ N_RESET_B_c_941_n N_RESET_B_c_1052_p PM_SKY130_FD_SC_MS__SDFRTP_2%RESET_B
x_PM_SKY130_FD_SC_MS__SDFRTP_2%A_1235_119# N_A_1235_119#_M1031_d
+ N_A_1235_119#_M1002_d N_A_1235_119#_M1013_d N_A_1235_119#_M1040_g
+ N_A_1235_119#_M1006_g N_A_1235_119#_c_1138_n N_A_1235_119#_c_1139_n
+ N_A_1235_119#_c_1148_n N_A_1235_119#_c_1140_n N_A_1235_119#_c_1177_n
+ N_A_1235_119#_c_1141_n N_A_1235_119#_c_1142_n N_A_1235_119#_c_1143_n
+ N_A_1235_119#_c_1144_n N_A_1235_119#_c_1151_n
+ PM_SKY130_FD_SC_MS__SDFRTP_2%A_1235_119#
x_PM_SKY130_FD_SC_MS__SDFRTP_2%A_837_119# N_A_837_119#_M1016_s
+ N_A_837_119#_M1027_s N_A_837_119#_M1034_g N_A_837_119#_M1017_g
+ N_A_837_119#_c_1256_n N_A_837_119#_c_1257_n N_A_837_119#_c_1272_n
+ N_A_837_119#_c_1273_n N_A_837_119#_c_1258_n N_A_837_119#_c_1259_n
+ N_A_837_119#_c_1274_n N_A_837_119#_c_1275_n N_A_837_119#_c_1260_n
+ N_A_837_119#_M1031_g N_A_837_119#_M1025_g N_A_837_119#_c_1277_n
+ N_A_837_119#_M1020_g N_A_837_119#_c_1261_n N_A_837_119#_c_1280_n
+ N_A_837_119#_c_1262_n N_A_837_119#_M1009_g N_A_837_119#_c_1264_n
+ N_A_837_119#_c_1265_n N_A_837_119#_c_1282_n N_A_837_119#_c_1266_n
+ N_A_837_119#_c_1288_n N_A_837_119#_c_1291_n N_A_837_119#_c_1267_n
+ N_A_837_119#_c_1283_n N_A_837_119#_c_1268_n N_A_837_119#_c_1300_n
+ N_A_837_119#_c_1269_n N_A_837_119#_c_1270_n N_A_837_119#_c_1271_n
+ N_A_837_119#_c_1286_n PM_SKY130_FD_SC_MS__SDFRTP_2%A_837_119#
x_PM_SKY130_FD_SC_MS__SDFRTP_2%A_2082_446# N_A_2082_446#_M1018_d
+ N_A_2082_446#_M1019_d N_A_2082_446#_M1005_g N_A_2082_446#_M1010_g
+ N_A_2082_446#_c_1469_n N_A_2082_446#_c_1481_n N_A_2082_446#_c_1460_n
+ N_A_2082_446#_c_1461_n N_A_2082_446#_c_1472_n N_A_2082_446#_c_1528_p
+ N_A_2082_446#_c_1473_n N_A_2082_446#_c_1462_n N_A_2082_446#_c_1463_n
+ N_A_2082_446#_c_1464_n N_A_2082_446#_c_1465_n N_A_2082_446#_c_1466_n
+ N_A_2082_446#_c_1467_n PM_SKY130_FD_SC_MS__SDFRTP_2%A_2082_446#
x_PM_SKY130_FD_SC_MS__SDFRTP_2%A_1824_74# N_A_1824_74#_M1028_d
+ N_A_1824_74#_M1020_d N_A_1824_74#_M1018_g N_A_1824_74#_c_1592_n
+ N_A_1824_74#_M1024_g N_A_1824_74#_c_1579_n N_A_1824_74#_c_1580_n
+ N_A_1824_74#_M1037_g N_A_1824_74#_c_1582_n N_A_1824_74#_M1029_g
+ N_A_1824_74#_c_1583_n N_A_1824_74#_c_1584_n N_A_1824_74#_c_1601_n
+ N_A_1824_74#_c_1585_n N_A_1824_74#_c_1595_n N_A_1824_74#_c_1596_n
+ N_A_1824_74#_c_1586_n N_A_1824_74#_c_1587_n N_A_1824_74#_c_1588_n
+ N_A_1824_74#_c_1589_n N_A_1824_74#_c_1590_n N_A_1824_74#_c_1591_n
+ PM_SKY130_FD_SC_MS__SDFRTP_2%A_1824_74#
x_PM_SKY130_FD_SC_MS__SDFRTP_2%A_2495_392# N_A_2495_392#_M1029_d
+ N_A_2495_392#_M1037_d N_A_2495_392#_M1001_g N_A_2495_392#_M1003_g
+ N_A_2495_392#_M1041_g N_A_2495_392#_M1030_g N_A_2495_392#_c_1726_n
+ N_A_2495_392#_c_1727_n N_A_2495_392#_c_1719_n N_A_2495_392#_c_1720_n
+ N_A_2495_392#_c_1721_n N_A_2495_392#_c_1722_n N_A_2495_392#_c_1723_n
+ PM_SKY130_FD_SC_MS__SDFRTP_2%A_2495_392#
x_PM_SKY130_FD_SC_MS__SDFRTP_2%VPWR N_VPWR_M1011_d N_VPWR_M1039_d N_VPWR_M1027_d
+ N_VPWR_M1033_d N_VPWR_M1006_s N_VPWR_M1005_d N_VPWR_M1024_d N_VPWR_M1001_d
+ N_VPWR_M1041_d N_VPWR_c_1778_n N_VPWR_c_1779_n N_VPWR_c_1780_n N_VPWR_c_1781_n
+ N_VPWR_c_1782_n N_VPWR_c_1783_n N_VPWR_c_1784_n N_VPWR_c_1785_n
+ N_VPWR_c_1786_n N_VPWR_c_1787_n N_VPWR_c_1788_n N_VPWR_c_1789_n
+ N_VPWR_c_1790_n N_VPWR_c_1791_n VPWR N_VPWR_c_1792_n N_VPWR_c_1793_n
+ N_VPWR_c_1794_n N_VPWR_c_1795_n N_VPWR_c_1796_n N_VPWR_c_1797_n
+ N_VPWR_c_1798_n N_VPWR_c_1799_n N_VPWR_c_1800_n N_VPWR_c_1801_n
+ N_VPWR_c_1802_n N_VPWR_c_1777_n PM_SKY130_FD_SC_MS__SDFRTP_2%VPWR
x_PM_SKY130_FD_SC_MS__SDFRTP_2%A_390_81# N_A_390_81#_M1015_d N_A_390_81#_M1031_s
+ N_A_390_81#_M1000_d N_A_390_81#_M1023_d N_A_390_81#_M1002_s
+ N_A_390_81#_c_1956_n N_A_390_81#_c_1947_n N_A_390_81#_c_1957_n
+ N_A_390_81#_c_1958_n N_A_390_81#_c_1948_n N_A_390_81#_c_1949_n
+ N_A_390_81#_c_1950_n N_A_390_81#_c_1951_n N_A_390_81#_c_1960_n
+ N_A_390_81#_c_1961_n N_A_390_81#_c_1952_n N_A_390_81#_c_1962_n
+ N_A_390_81#_c_1963_n N_A_390_81#_c_1953_n N_A_390_81#_c_1954_n
+ N_A_390_81#_c_1955_n N_A_390_81#_c_1965_n
+ PM_SKY130_FD_SC_MS__SDFRTP_2%A_390_81#
x_PM_SKY130_FD_SC_MS__SDFRTP_2%Q N_Q_M1003_d N_Q_M1001_s N_Q_c_2116_n Q Q Q Q
+ PM_SKY130_FD_SC_MS__SDFRTP_2%Q
x_PM_SKY130_FD_SC_MS__SDFRTP_2%VGND N_VGND_M1036_d N_VGND_M1004_d N_VGND_M1016_d
+ N_VGND_M1007_d N_VGND_M1010_d N_VGND_M1029_s N_VGND_M1003_s N_VGND_M1030_s
+ N_VGND_c_2137_n N_VGND_c_2138_n N_VGND_c_2139_n N_VGND_c_2140_n
+ N_VGND_c_2141_n N_VGND_c_2142_n N_VGND_c_2143_n N_VGND_c_2144_n
+ N_VGND_c_2145_n N_VGND_c_2146_n N_VGND_c_2147_n N_VGND_c_2148_n VGND
+ N_VGND_c_2149_n N_VGND_c_2150_n N_VGND_c_2151_n N_VGND_c_2152_n
+ N_VGND_c_2153_n N_VGND_c_2154_n N_VGND_c_2155_n N_VGND_c_2156_n
+ N_VGND_c_2157_n N_VGND_c_2158_n N_VGND_c_2159_n
+ PM_SKY130_FD_SC_MS__SDFRTP_2%VGND
x_PM_SKY130_FD_SC_MS__SDFRTP_2%noxref_24 N_noxref_24_M1014_s N_noxref_24_M1035_d
+ N_noxref_24_c_2273_n N_noxref_24_c_2289_n N_noxref_24_c_2274_n
+ PM_SKY130_FD_SC_MS__SDFRTP_2%noxref_24
cc_1 VNB N_A_27_74#_c_291_n 0.0258189f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_2 VNB N_A_27_74#_c_292_n 0.0202565f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.935
cc_3 VNB N_A_27_74#_c_293_n 0.0257773f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_4 VNB N_A_27_74#_c_294_n 0.0190417f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.005
cc_5 VNB N_A_27_74#_c_295_n 0.00987534f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_6 VNB N_A_27_74#_c_296_n 0.018224f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_7 VNB N_A_27_74#_c_297_n 0.0395906f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.01
cc_8 VNB N_SCE_M1036_g 0.0668709f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_9 VNB N_SCE_c_375_n 0.00775502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_SCE_c_376_n 0.0420243f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.265
cc_11 VNB N_SCE_c_377_n 0.0151284f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.005
cc_12 VNB N_SCE_c_378_n 0.0142876f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.175
cc_13 VNB N_SCE_c_379_n 0.0118824f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.465
cc_14 VNB N_SCE_c_380_n 0.0057985f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.1
cc_15 VNB N_SCE_c_381_n 0.0297083f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_16 VNB N_SCE_c_382_n 0.01224f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_17 VNB N_SCE_c_383_n 0.0106235f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=2.16
cc_18 VNB N_SCE_c_384_n 0.00168276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_D_M1000_g 0.0271007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_D_c_460_n 0.0364471f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_21 VNB N_D_c_461_n 0.00754927f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.16
cc_22 VNB N_D_c_462_n 0.016179f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.735
cc_23 VNB N_SCD_M1035_g 0.0417173f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_24 VNB N_SCD_c_504_n 9.06233e-19 $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_25 VNB SCD 0.00275067f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.735
cc_26 VNB N_SCD_c_506_n 0.0155389f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_27 VNB N_CLK_c_551_n 0.0223227f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=0.37
cc_28 VNB CLK 0.0200716f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_29 VNB N_CLK_c_553_n 0.0322566f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.735
cc_30 VNB N_CLK_c_554_n 0.0215445f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_31 VNB N_CLK_c_555_n 0.0149759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_1037_119#_c_611_n 0.00800051f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.615
cc_33 VNB N_A_1037_119#_c_612_n 0.0267885f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.735
cc_34 VNB N_A_1037_119#_M1032_g 0.027122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_1037_119#_c_614_n 0.0171555f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_36 VNB N_A_1037_119#_c_615_n 0.0222225f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.265
cc_37 VNB N_A_1037_119#_c_616_n 0.0102361f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.005
cc_38 VNB N_A_1037_119#_c_617_n 0.00215883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_1037_119#_c_618_n 0.00105427f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=2.09
cc_40 VNB N_A_1037_119#_c_619_n 0.0412395f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_41 VNB N_A_1037_119#_c_620_n 0.00358858f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.09
cc_42 VNB N_A_1037_119#_c_621_n 0.00213605f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_43 VNB N_A_1037_119#_c_622_n 0.00235278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_1037_119#_c_623_n 0.00854373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_1037_119#_c_624_n 0.00229566f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_46 VNB N_A_1037_119#_c_625_n 0.00595338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1037_119#_c_626_n 0.00363165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1037_119#_c_627_n 0.0322711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1037_119#_c_628_n 0.0101868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1037_119#_c_629_n 0.00285652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1037_119#_c_630_n 2.38103e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1037_119#_c_631_n 0.0046617f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1037_119#_c_632_n 0.0117715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1383_349#_M1022_g 0.0389668f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.735
cc_55 VNB N_A_1383_349#_c_826_n 0.00413621f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_56 VNB N_A_1383_349#_c_827_n 0.00304711f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.265
cc_57 VNB N_A_1383_349#_c_828_n 0.00239154f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_58 VNB N_A_1383_349#_c_829_n 0.0143226f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=1.995
cc_59 VNB N_RESET_B_c_917_n 0.0293798f $X=-0.19 $Y=-0.245 $X2=0.135 $Y2=2.32
cc_60 VNB N_RESET_B_M1004_g 0.0143778f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_61 VNB N_RESET_B_c_919_n 0.284303f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.615
cc_62 VNB N_RESET_B_c_920_n 0.012806f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.16
cc_63 VNB N_RESET_B_M1007_g 0.03552f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.935
cc_64 VNB N_RESET_B_c_922_n 0.0189013f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=2.175
cc_65 VNB N_RESET_B_M1026_g 0.0531601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_RESET_B_c_924_n 0.0155543f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=2.09
cc_67 VNB N_RESET_B_c_925_n 0.0224087f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_68 VNB N_A_1235_119#_M1040_g 0.0241865f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.16
cc_69 VNB N_A_1235_119#_c_1138_n 0.0274099f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_70 VNB N_A_1235_119#_c_1139_n 0.0172233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1235_119#_c_1140_n 0.00406303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1235_119#_c_1141_n 5.47821e-19 $X=-0.19 $Y=-0.245 $X2=0.975
+ $Y2=1.1
cc_73 VNB N_A_1235_119#_c_1142_n 0.00159936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1235_119#_c_1143_n 0.00560512f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=2.09
cc_75 VNB N_A_1235_119#_c_1144_n 0.00436197f $X=-0.19 $Y=-0.245 $X2=2.5
+ $Y2=1.995
cc_76 VNB N_A_837_119#_c_1256_n 0.00915784f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.735
cc_77 VNB N_A_837_119#_c_1257_n 0.00896212f $X=-0.19 $Y=-0.245 $X2=0.24
+ $Y2=0.935
cc_78 VNB N_A_837_119#_c_1258_n 0.0323794f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.005
cc_79 VNB N_A_837_119#_c_1259_n 0.00946783f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.175
cc_80 VNB N_A_837_119#_c_1260_n 0.0168105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_837_119#_c_1261_n 0.012531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_837_119#_c_1262_n 0.0236403f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.01
cc_83 VNB N_A_837_119#_M1009_g 0.027022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_837_119#_c_1264_n 0.00731326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_837_119#_c_1265_n 0.00504746f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=2.16
cc_86 VNB N_A_837_119#_c_1266_n 0.0209137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_837_119#_c_1267_n 0.00164026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_837_119#_c_1268_n 0.00522229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_837_119#_c_1269_n 0.00177279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_837_119#_c_1270_n 0.0175279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_837_119#_c_1271_n 0.0155629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_2082_446#_M1010_g 0.0407896f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.735
cc_93 VNB N_A_2082_446#_c_1460_n 0.00604102f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.175
cc_94 VNB N_A_2082_446#_c_1461_n 0.00978233f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.465
cc_95 VNB N_A_2082_446#_c_1462_n 0.00743589f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.1
cc_96 VNB N_A_2082_446#_c_1463_n 0.00688415f $X=-0.19 $Y=-0.245 $X2=2.54
+ $Y2=1.995
cc_97 VNB N_A_2082_446#_c_1464_n 0.00281201f $X=-0.19 $Y=-0.245 $X2=2.5
+ $Y2=1.995
cc_98 VNB N_A_2082_446#_c_1465_n 0.00528256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_2082_446#_c_1466_n 0.00129589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_2082_446#_c_1467_n 0.0231274f $X=-0.19 $Y=-0.245 $X2=0.975
+ $Y2=1.01
cc_101 VNB N_A_1824_74#_M1018_g 0.0313995f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.935
cc_102 VNB N_A_1824_74#_c_1579_n 0.0313227f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=0.58
cc_103 VNB N_A_1824_74#_c_1580_n 0.0323107f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=0.58
cc_104 VNB N_A_1824_74#_M1037_g 0.0156535f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.005
cc_105 VNB N_A_1824_74#_c_1582_n 0.0193338f $X=-0.19 $Y=-0.245 $X2=0.28
+ $Y2=2.465
cc_106 VNB N_A_1824_74#_c_1583_n 0.0143534f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.1
cc_107 VNB N_A_1824_74#_c_1584_n 0.0203145f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_108 VNB N_A_1824_74#_c_1585_n 0.00728448f $X=-0.19 $Y=-0.245 $X2=0.445
+ $Y2=2.09
cc_109 VNB N_A_1824_74#_c_1586_n 0.00580575f $X=-0.19 $Y=-0.245 $X2=0.975
+ $Y2=1.01
cc_110 VNB N_A_1824_74#_c_1587_n 0.00783827f $X=-0.19 $Y=-0.245 $X2=0.975
+ $Y2=1.1
cc_111 VNB N_A_1824_74#_c_1588_n 0.0103967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_1824_74#_c_1589_n 4.11765e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_1824_74#_c_1590_n 0.0164314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_1824_74#_c_1591_n 0.00253069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_2495_392#_M1001_g 0.00189158f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=0.935
cc_116 VNB N_A_2495_392#_M1003_g 0.0229518f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.735
cc_117 VNB N_A_2495_392#_M1041_g 0.00231818f $X=-0.19 $Y=-0.245 $X2=0.24
+ $Y2=0.58
cc_118 VNB N_A_2495_392#_M1030_g 0.0260209f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=2.005
cc_119 VNB N_A_2495_392#_c_1719_n 0.0162202f $X=-0.19 $Y=-0.245 $X2=2.375
+ $Y2=2.09
cc_120 VNB N_A_2495_392#_c_1720_n 0.0113264f $X=-0.19 $Y=-0.245 $X2=2.5
+ $Y2=1.995
cc_121 VNB N_A_2495_392#_c_1721_n 7.87382e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_2495_392#_c_1722_n 0.00922601f $X=-0.19 $Y=-0.245 $X2=0.975
+ $Y2=1.01
cc_123 VNB N_A_2495_392#_c_1723_n 0.0847287f $X=-0.19 $Y=-0.245 $X2=2.5
+ $Y2=1.995
cc_124 VNB N_VPWR_c_1777_n 0.601534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_390_81#_c_1947_n 0.00863948f $X=-0.19 $Y=-0.245 $X2=0.2 $Y2=1.265
cc_126 VNB N_A_390_81#_c_1948_n 0.00280061f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_127 VNB N_A_390_81#_c_1949_n 0.014315f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_128 VNB N_A_390_81#_c_1950_n 0.00270766f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_129 VNB N_A_390_81#_c_1951_n 0.00249563f $X=-0.19 $Y=-0.245 $X2=2.375
+ $Y2=2.09
cc_130 VNB N_A_390_81#_c_1952_n 0.00151767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_A_390_81#_c_1953_n 0.00953662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_A_390_81#_c_1954_n 0.00360151f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=1.995
cc_133 VNB N_A_390_81#_c_1955_n 0.00170226f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=2.16
cc_134 VNB N_Q_c_2116_n 2.86109e-19 $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.935
cc_135 VNB Q 0.00240191f $X=-0.19 $Y=-0.245 $X2=2.495 $Y2=2.735
cc_136 VNB N_VGND_c_2137_n 0.0110567f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_137 VNB N_VGND_c_2138_n 0.0133929f $X=-0.19 $Y=-0.245 $X2=2.375 $Y2=2.09
cc_138 VNB N_VGND_c_2139_n 0.00960261f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=1.995
cc_139 VNB N_VGND_c_2140_n 0.0067048f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=2.09
cc_140 VNB N_VGND_c_2141_n 0.00861345f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.1
cc_141 VNB N_VGND_c_2142_n 0.0169646f $X=-0.19 $Y=-0.245 $X2=2.5 $Y2=2.16
cc_142 VNB N_VGND_c_2143_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2144_n 0.0505973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2145_n 0.0659799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2146_n 0.00399507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2147_n 0.0204564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2148_n 0.0034624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2149_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2150_n 0.0784397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2151_n 0.0684884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2152_n 0.0296745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2153_n 0.0187654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2154_n 0.0193312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2155_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2156_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2157_n 0.00613227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_2158_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2159_n 0.748115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_noxref_24_c_2273_n 0.0172763f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.01
cc_160 VNB N_noxref_24_c_2274_n 0.00655627f $X=-0.19 $Y=-0.245 $X2=2.495
+ $Y2=2.735
cc_161 VPB N_A_27_74#_M1038_g 0.0271114f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.735
cc_162 VPB N_A_27_74#_c_294_n 0.016494f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.005
cc_163 VPB N_A_27_74#_c_300_n 0.0337004f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_164 VPB N_A_27_74#_c_301_n 0.0343789f $X=-0.19 $Y=1.66 $X2=2.375 $Y2=2.09
cc_165 VPB N_A_27_74#_c_302_n 0.0129728f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_166 VPB N_A_27_74#_c_303_n 0.0060227f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_167 VPB N_A_27_74#_c_304_n 0.0277775f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_168 VPB N_SCE_M1011_g 0.0591491f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_SCE_M1012_g 0.0569663f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_170 VPB N_SCE_c_375_n 0.00782879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_SCE_c_376_n 0.0410198f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.265
cc_172 VPB N_SCE_c_380_n 0.00211749f $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_173 VPB N_SCE_c_384_n 0.0026972f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_D_M1000_g 0.0555291f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_SCD_M1039_g 0.0276542f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_SCD_c_504_n 0.0258731f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_177 VPB N_SCD_c_509_n 0.0143222f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.16
cc_178 VPB SCD 0.00440777f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.735
cc_179 VPB N_CLK_M1027_g 0.0255463f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=1.01
cc_180 VPB CLK 0.00482818f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.615
cc_181 VPB N_CLK_c_554_n 0.0127548f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_182 VPB N_A_1037_119#_M1002_g 0.0291921f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.935
cc_183 VPB N_A_1037_119#_c_611_n 0.00961448f $X=-0.19 $Y=1.66 $X2=1.485
+ $Y2=0.615
cc_184 VPB N_A_1037_119#_c_612_n 0.00971273f $X=-0.19 $Y=1.66 $X2=2.495
+ $Y2=2.735
cc_185 VPB N_A_1037_119#_M1021_g 0.0280945f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_186 VPB N_A_1037_119#_c_621_n 0.00174889f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_187 VPB N_A_1037_119#_c_628_n 0.0064161f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_1037_119#_c_630_n 0.00270697f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_189 VPB N_A_1037_119#_c_632_n 0.0240192f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_190 VPB N_A_1037_119#_c_641_n 0.0394518f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_191 VPB N_A_1383_349#_M1033_g 0.0244689f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.935
cc_192 VPB N_A_1383_349#_M1022_g 0.00462646f $X=-0.19 $Y=1.66 $X2=2.495
+ $Y2=2.735
cc_193 VPB N_A_1383_349#_c_826_n 0.00156886f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.58
cc_194 VPB N_A_1383_349#_c_833_n 0.0453043f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_195 VPB N_A_1383_349#_c_834_n 5.83247e-19 $X=-0.19 $Y=1.66 $X2=0.365 $Y2=1.1
cc_196 VPB N_A_1383_349#_c_835_n 0.00551405f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_197 VPB N_A_1383_349#_c_829_n 0.00449421f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=1.995
cc_198 VPB N_RESET_B_c_917_n 0.0102676f $X=-0.19 $Y=1.66 $X2=0.135 $Y2=2.32
cc_199 VPB N_RESET_B_M1023_g 0.0312081f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_RESET_B_M1013_g 0.0256766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_RESET_B_c_922_n 0.0105327f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.175
cc_202 VPB N_RESET_B_M1026_g 0.0132171f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_RESET_B_M1019_g 0.0324286f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_204 VPB N_RESET_B_c_932_n 0.0127772f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_205 VPB N_RESET_B_c_933_n 0.0193703f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=2.09
cc_206 VPB N_RESET_B_c_934_n 0.00173686f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_RESET_B_c_935_n 0.0135889f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.01
cc_208 VPB N_RESET_B_c_936_n 3.23518e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_209 VPB N_RESET_B_c_937_n 0.0118766f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_210 VPB N_RESET_B_c_938_n 0.0516141f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_211 VPB N_RESET_B_c_939_n 0.00288093f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_212 VPB N_RESET_B_c_940_n 0.0528936f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_213 VPB N_RESET_B_c_941_n 0.0351975f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_1235_119#_M1006_g 0.0267004f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.935
cc_215 VPB N_A_1235_119#_c_1138_n 0.00914718f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_216 VPB N_A_1235_119#_c_1139_n 0.00381103f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_A_1235_119#_c_1148_n 0.00280501f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.265
cc_218 VPB N_A_1235_119#_c_1140_n 0.0101341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_A_1235_119#_c_1141_n 0.0105848f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_220 VPB N_A_1235_119#_c_1151_n 0.00191608f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_A_837_119#_c_1272_n 0.00460432f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_A_837_119#_c_1273_n 0.0511184f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=1.265
cc_223 VPB N_A_837_119#_c_1274_n 0.0569553f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_224 VPB N_A_837_119#_c_1275_n 0.0111463f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_225 VPB N_A_837_119#_M1025_g 0.0404743f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_A_837_119#_c_1277_n 0.19503f $X=-0.19 $Y=1.66 $X2=0.445 $Y2=2.09
cc_227 VPB N_A_837_119#_M1020_g 0.026642f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_228 VPB N_A_837_119#_c_1261_n 0.03645f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_A_837_119#_c_1280_n 0.00994735f $X=-0.19 $Y=1.66 $X2=2.54 $Y2=2.09
cc_230 VPB N_A_837_119#_c_1265_n 0.0230177f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=2.16
cc_231 VPB N_A_837_119#_c_1282_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_A_837_119#_c_1283_n 0.00248018f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_A_837_119#_c_1269_n 9.43952e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_A_837_119#_c_1270_n 0.0153562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_A_837_119#_c_1286_n 0.0165206f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_A_2082_446#_M1005_g 0.0228197f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.935
cc_237 VPB N_A_2082_446#_c_1469_n 0.0217114f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.58
cc_238 VPB N_A_2082_446#_c_1460_n 0.0447354f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.175
cc_239 VPB N_A_2082_446#_c_1461_n 0.0137444f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_240 VPB N_A_2082_446#_c_1472_n 0.00779622f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_241 VPB N_A_2082_446#_c_1473_n 0.0023101f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_242 VPB N_A_1824_74#_c_1592_n 0.00554553f $X=-0.19 $Y=1.66 $X2=1.485
+ $Y2=0.615
cc_243 VPB N_A_1824_74#_M1024_g 0.0606802f $X=-0.19 $Y=1.66 $X2=2.495 $Y2=2.735
cc_244 VPB N_A_1824_74#_M1037_g 0.0342788f $X=-0.19 $Y=1.66 $X2=0.2 $Y2=2.005
cc_245 VPB N_A_1824_74#_c_1595_n 0.00597636f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_246 VPB N_A_1824_74#_c_1596_n 0.00270733f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_247 VPB N_A_1824_74#_c_1587_n 0.0143637f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_248 VPB N_A_2495_392#_M1001_g 0.0259836f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.935
cc_249 VPB N_A_2495_392#_M1041_g 0.0274054f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=0.58
cc_250 VPB N_A_2495_392#_c_1726_n 0.00488438f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_251 VPB N_A_2495_392#_c_1727_n 0.0103543f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_252 VPB N_A_2495_392#_c_1721_n 0.00694126f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1778_n 0.00151893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1779_n 0.00151893f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_255 VPB N_VPWR_c_1780_n 0.0153422f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1781_n 0.0188146f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1782_n 0.019438f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1783_n 0.0184521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1784_n 0.0121909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1785_n 0.0688078f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1786_n 0.0327672f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1787_n 0.00485379f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1788_n 0.0582875f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1789_n 0.00443527f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1790_n 0.0198404f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1791_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1792_n 0.0191816f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1793_n 0.0437698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1794_n 0.0206273f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1795_n 0.0534696f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1796_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1797_n 0.0174925f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1798_n 0.0292631f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1799_n 0.00485691f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1800_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1801_n 0.0230715f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1802_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1777_n 0.109393f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_279 VPB N_A_390_81#_c_1956_n 0.00203831f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=0.58
cc_280 VPB N_A_390_81#_c_1957_n 0.0134125f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.465
cc_281 VPB N_A_390_81#_c_1958_n 0.00239826f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_282 VPB N_A_390_81#_c_1951_n 0.0116459f $X=-0.19 $Y=1.66 $X2=2.375 $Y2=2.09
cc_283 VPB N_A_390_81#_c_1960_n 0.0116707f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=2.09
cc_284 VPB N_A_390_81#_c_1961_n 0.00475312f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=1.995
cc_285 VPB N_A_390_81#_c_1962_n 0.00128301f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_286 VPB N_A_390_81#_c_1963_n 0.00322424f $X=-0.19 $Y=1.66 $X2=0.975 $Y2=1.1
cc_287 VPB N_A_390_81#_c_1955_n 0.00509989f $X=-0.19 $Y=1.66 $X2=2.5 $Y2=2.16
cc_288 VPB N_A_390_81#_c_1965_n 0.0159146f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_289 VPB N_Q_c_2116_n 0.00380841f $X=-0.19 $Y=1.66 $X2=1.485 $Y2=0.935
cc_290 N_A_27_74#_c_300_n N_SCE_M1011_g 0.0184741f $X=0.28 $Y=2.465 $X2=0 $Y2=0
cc_291 N_A_27_74#_c_301_n N_SCE_M1011_g 0.0195433f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_292 N_A_27_74#_c_302_n N_SCE_M1011_g 0.00544367f $X=0.28 $Y=2.09 $X2=0 $Y2=0
cc_293 N_A_27_74#_c_293_n N_SCE_M1036_g 0.00686809f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_294 N_A_27_74#_c_294_n N_SCE_M1036_g 0.00830473f $X=0.2 $Y=2.005 $X2=0 $Y2=0
cc_295 N_A_27_74#_c_295_n N_SCE_M1036_g 0.0281157f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_296 N_A_27_74#_c_297_n N_SCE_M1036_g 0.0181297f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_297 N_A_27_74#_c_301_n N_SCE_M1012_g 0.0181012f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_298 N_A_27_74#_c_294_n N_SCE_c_375_n 0.0158921f $X=0.2 $Y=2.005 $X2=0 $Y2=0
cc_299 N_A_27_74#_c_295_n N_SCE_c_375_n 0.00162366f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_300 N_A_27_74#_c_291_n N_SCE_c_376_n 0.0106974f $X=1.41 $Y=1.01 $X2=0 $Y2=0
cc_301 N_A_27_74#_c_295_n N_SCE_c_376_n 0.00180358f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_302 N_A_27_74#_c_301_n N_SCE_c_376_n 0.0170396f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_303 N_A_27_74#_c_297_n N_SCE_c_376_n 0.0175645f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_304 N_A_27_74#_c_301_n N_SCE_c_379_n 0.0251991f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_305 N_A_27_74#_c_304_n N_SCE_c_379_n 3.04821e-19 $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_306 N_A_27_74#_c_303_n N_SCE_c_380_n 0.0268647f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_307 N_A_27_74#_c_304_n N_SCE_c_380_n 0.00100599f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_308 N_A_27_74#_c_303_n N_SCE_c_381_n 3.17572e-19 $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_309 N_A_27_74#_c_304_n N_SCE_c_381_n 0.0181417f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_310 N_A_27_74#_c_291_n N_SCE_c_383_n 0.00818136f $X=1.41 $Y=1.01 $X2=0 $Y2=0
cc_311 N_A_27_74#_c_294_n N_SCE_c_383_n 0.0170838f $X=0.2 $Y=2.005 $X2=0 $Y2=0
cc_312 N_A_27_74#_c_295_n N_SCE_c_383_n 0.0353374f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_313 N_A_27_74#_c_301_n N_SCE_c_383_n 0.0893268f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_314 N_A_27_74#_c_297_n N_SCE_c_383_n 0.00202099f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_315 N_A_27_74#_M1038_g N_D_M1000_g 0.0191772f $X=2.495 $Y=2.735 $X2=0 $Y2=0
cc_316 N_A_27_74#_c_301_n N_D_M1000_g 0.0169877f $X=2.375 $Y=2.09 $X2=0 $Y2=0
cc_317 N_A_27_74#_c_303_n N_D_M1000_g 0.00117555f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_318 N_A_27_74#_c_304_n N_D_M1000_g 0.0214638f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_319 N_A_27_74#_c_291_n N_D_c_460_n 0.00979672f $X=1.41 $Y=1.01 $X2=0 $Y2=0
cc_320 N_A_27_74#_c_295_n N_D_c_460_n 2.46837e-19 $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_321 N_A_27_74#_c_297_n N_D_c_460_n 0.00223442f $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_322 N_A_27_74#_c_292_n N_D_c_461_n 0.00558783f $X=1.485 $Y=0.935 $X2=0 $Y2=0
cc_323 N_A_27_74#_c_295_n N_D_c_461_n 0.0143876f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_324 N_A_27_74#_c_297_n N_D_c_461_n 8.79717e-19 $X=0.975 $Y=1.01 $X2=0 $Y2=0
cc_325 N_A_27_74#_c_292_n N_D_c_462_n 0.0356736f $X=1.485 $Y=0.935 $X2=0 $Y2=0
cc_326 N_A_27_74#_M1038_g N_SCD_M1039_g 0.0355942f $X=2.495 $Y=2.735 $X2=0 $Y2=0
cc_327 N_A_27_74#_c_303_n N_SCD_M1039_g 5.52836e-19 $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_328 N_A_27_74#_c_304_n N_SCD_M1039_g 3.99404e-19 $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_329 N_A_27_74#_c_303_n N_SCD_c_504_n 0.00210253f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_330 N_A_27_74#_c_304_n N_SCD_c_504_n 0.0199742f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_331 N_A_27_74#_c_303_n SCD 0.019551f $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_332 N_A_27_74#_c_304_n SCD 3.37003e-19 $X=2.5 $Y=1.995 $X2=0 $Y2=0
cc_333 N_A_27_74#_M1038_g N_VPWR_c_1778_n 0.00191337f $X=2.495 $Y=2.735 $X2=0
+ $Y2=0
cc_334 N_A_27_74#_c_300_n N_VPWR_c_1792_n 0.014549f $X=0.28 $Y=2.465 $X2=0 $Y2=0
cc_335 N_A_27_74#_M1038_g N_VPWR_c_1793_n 0.00613344f $X=2.495 $Y=2.735 $X2=0
+ $Y2=0
cc_336 N_A_27_74#_c_300_n N_VPWR_c_1798_n 0.0247088f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_337 N_A_27_74#_c_301_n N_VPWR_c_1798_n 0.0769127f $X=2.375 $Y=2.09 $X2=0
+ $Y2=0
cc_338 N_A_27_74#_M1038_g N_VPWR_c_1777_n 0.00695261f $X=2.495 $Y=2.735 $X2=0
+ $Y2=0
cc_339 N_A_27_74#_c_300_n N_VPWR_c_1777_n 0.0119743f $X=0.28 $Y=2.465 $X2=0
+ $Y2=0
cc_340 N_A_27_74#_M1038_g N_A_390_81#_c_1956_n 0.0120918f $X=2.495 $Y=2.735
+ $X2=0 $Y2=0
cc_341 N_A_27_74#_M1038_g N_A_390_81#_c_1957_n 0.0101887f $X=2.495 $Y=2.735
+ $X2=0 $Y2=0
cc_342 N_A_27_74#_c_303_n N_A_390_81#_c_1957_n 0.0202835f $X=2.5 $Y=1.995 $X2=0
+ $Y2=0
cc_343 N_A_27_74#_c_304_n N_A_390_81#_c_1957_n 5.39896e-19 $X=2.5 $Y=1.995 $X2=0
+ $Y2=0
cc_344 N_A_27_74#_M1038_g N_A_390_81#_c_1958_n 0.00171171f $X=2.495 $Y=2.735
+ $X2=0 $Y2=0
cc_345 N_A_27_74#_c_301_n N_A_390_81#_c_1958_n 0.0226379f $X=2.375 $Y=2.09 $X2=0
+ $Y2=0
cc_346 N_A_27_74#_c_303_n N_A_390_81#_c_1958_n 0.00499989f $X=2.5 $Y=1.995 $X2=0
+ $Y2=0
cc_347 N_A_27_74#_c_304_n N_A_390_81#_c_1958_n 5.24165e-19 $X=2.5 $Y=1.995 $X2=0
+ $Y2=0
cc_348 N_A_27_74#_c_292_n N_VGND_c_2137_n 0.00287309f $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_349 N_A_27_74#_c_293_n N_VGND_c_2137_n 0.0156021f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_350 N_A_27_74#_c_295_n N_VGND_c_2137_n 0.0254818f $X=0.975 $Y=1.1 $X2=0 $Y2=0
cc_351 N_A_27_74#_c_297_n N_VGND_c_2137_n 0.00149092f $X=0.975 $Y=1.01 $X2=0
+ $Y2=0
cc_352 N_A_27_74#_c_292_n N_VGND_c_2145_n 9.09582e-19 $X=1.485 $Y=0.935 $X2=0
+ $Y2=0
cc_353 N_A_27_74#_c_293_n N_VGND_c_2149_n 0.011066f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_354 N_A_27_74#_c_293_n N_VGND_c_2159_n 0.00915947f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_355 N_A_27_74#_c_292_n N_noxref_24_c_2273_n 0.0108727f $X=1.485 $Y=0.935
+ $X2=0 $Y2=0
cc_356 N_A_27_74#_c_292_n N_noxref_24_c_2274_n 0.00859442f $X=1.485 $Y=0.935
+ $X2=0 $Y2=0
cc_357 N_A_27_74#_c_295_n N_noxref_24_c_2274_n 0.00178881f $X=0.975 $Y=1.1 $X2=0
+ $Y2=0
cc_358 N_A_27_74#_c_297_n N_noxref_24_c_2274_n 0.00859402f $X=0.975 $Y=1.01
+ $X2=0 $Y2=0
cc_359 N_SCE_c_376_n N_D_M1000_g 0.0944756f $X=1.535 $Y=1.67 $X2=0 $Y2=0
cc_360 N_SCE_c_379_n N_D_M1000_g 0.0140585f $X=2.375 $Y=1.575 $X2=0 $Y2=0
cc_361 N_SCE_c_380_n N_D_M1000_g 3.24847e-19 $X=2.5 $Y=1.425 $X2=0 $Y2=0
cc_362 N_SCE_c_384_n N_D_M1000_g 0.00483039f $X=1.795 $Y=1.662 $X2=0 $Y2=0
cc_363 N_SCE_c_378_n N_D_c_460_n 0.0112143f $X=2.625 $Y=1.05 $X2=0 $Y2=0
cc_364 N_SCE_c_380_n N_D_c_460_n 0.00141664f $X=2.5 $Y=1.425 $X2=0 $Y2=0
cc_365 N_SCE_c_381_n N_D_c_460_n 0.0214877f $X=2.5 $Y=1.425 $X2=0 $Y2=0
cc_366 N_SCE_c_384_n N_D_c_460_n 0.00432931f $X=1.795 $Y=1.662 $X2=0 $Y2=0
cc_367 N_SCE_c_376_n N_D_c_461_n 0.00106377f $X=1.535 $Y=1.67 $X2=0 $Y2=0
cc_368 N_SCE_c_377_n N_D_c_461_n 0.00118822f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_369 N_SCE_c_378_n N_D_c_461_n 0.00257293f $X=2.625 $Y=1.05 $X2=0 $Y2=0
cc_370 N_SCE_c_383_n N_D_c_461_n 0.0344557f $X=1.623 $Y=1.662 $X2=0 $Y2=0
cc_371 N_SCE_c_377_n N_D_c_462_n 0.00677849f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_372 N_SCE_c_378_n N_D_c_462_n 5.31722e-19 $X=2.625 $Y=1.05 $X2=0 $Y2=0
cc_373 N_SCE_c_377_n N_SCD_M1035_g 0.0414075f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_374 N_SCE_c_380_n N_SCD_M1035_g 0.00373757f $X=2.5 $Y=1.425 $X2=0 $Y2=0
cc_375 N_SCE_c_382_n N_SCD_M1035_g 0.0156026f $X=2.5 $Y=1.26 $X2=0 $Y2=0
cc_376 N_SCE_c_380_n SCD 0.010985f $X=2.5 $Y=1.425 $X2=0 $Y2=0
cc_377 N_SCE_c_380_n N_SCD_c_506_n 0.00236449f $X=2.5 $Y=1.425 $X2=0 $Y2=0
cc_378 N_SCE_c_381_n N_SCD_c_506_n 0.00687648f $X=2.5 $Y=1.425 $X2=0 $Y2=0
cc_379 N_SCE_M1011_g N_VPWR_c_1792_n 0.005209f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_380 N_SCE_M1012_g N_VPWR_c_1793_n 0.00545548f $X=1.625 $Y=2.735 $X2=0 $Y2=0
cc_381 N_SCE_M1011_g N_VPWR_c_1798_n 0.00585939f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_382 N_SCE_M1012_g N_VPWR_c_1798_n 0.0216934f $X=1.625 $Y=2.735 $X2=0 $Y2=0
cc_383 N_SCE_M1011_g N_VPWR_c_1777_n 0.00990469f $X=0.505 $Y=2.64 $X2=0 $Y2=0
cc_384 N_SCE_M1012_g N_VPWR_c_1777_n 0.00962554f $X=1.625 $Y=2.735 $X2=0 $Y2=0
cc_385 N_SCE_M1012_g N_A_390_81#_c_1956_n 0.00154346f $X=1.625 $Y=2.735 $X2=0
+ $Y2=0
cc_386 N_SCE_c_377_n N_A_390_81#_c_1947_n 0.0120699f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_387 N_SCE_c_378_n N_A_390_81#_c_1947_n 0.00236281f $X=2.625 $Y=1.05 $X2=0
+ $Y2=0
cc_388 N_SCE_c_379_n N_A_390_81#_c_1947_n 0.00306381f $X=2.375 $Y=1.575 $X2=0
+ $Y2=0
cc_389 N_SCE_c_380_n N_A_390_81#_c_1947_n 0.0129373f $X=2.5 $Y=1.425 $X2=0 $Y2=0
cc_390 N_SCE_c_381_n N_A_390_81#_c_1947_n 0.00169354f $X=2.5 $Y=1.425 $X2=0
+ $Y2=0
cc_391 N_SCE_M1012_g N_A_390_81#_c_1958_n 4.66801e-19 $X=1.625 $Y=2.735 $X2=0
+ $Y2=0
cc_392 N_SCE_c_377_n N_A_390_81#_c_1948_n 0.00432562f $X=2.625 $Y=0.9 $X2=0
+ $Y2=0
cc_393 N_SCE_c_382_n N_A_390_81#_c_1948_n 0.00177942f $X=2.5 $Y=1.26 $X2=0 $Y2=0
cc_394 N_SCE_c_380_n N_A_390_81#_c_1950_n 0.00442191f $X=2.5 $Y=1.425 $X2=0
+ $Y2=0
cc_395 N_SCE_c_382_n N_A_390_81#_c_1950_n 0.00318428f $X=2.5 $Y=1.26 $X2=0 $Y2=0
cc_396 N_SCE_M1036_g N_VGND_c_2137_n 0.0129468f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_397 N_SCE_c_377_n N_VGND_c_2145_n 9.15902e-19 $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_398 N_SCE_M1036_g N_VGND_c_2149_n 0.00383152f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_399 N_SCE_M1036_g N_VGND_c_2159_n 0.00761198f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_400 N_SCE_c_377_n N_noxref_24_c_2273_n 0.0107628f $X=2.625 $Y=0.9 $X2=0 $Y2=0
cc_401 N_SCE_M1036_g N_noxref_24_c_2274_n 9.19966e-19 $X=0.495 $Y=0.58 $X2=0
+ $Y2=0
cc_402 N_D_M1000_g N_VPWR_c_1793_n 0.0062759f $X=2.035 $Y=2.735 $X2=0 $Y2=0
cc_403 N_D_M1000_g N_VPWR_c_1798_n 0.00292617f $X=2.035 $Y=2.735 $X2=0 $Y2=0
cc_404 N_D_M1000_g N_VPWR_c_1777_n 0.0116416f $X=2.035 $Y=2.735 $X2=0 $Y2=0
cc_405 N_D_c_461_n N_A_390_81#_M1015_d 0.00160203f $X=1.935 $Y=1.1 $X2=-0.19
+ $Y2=-0.245
cc_406 N_D_M1000_g N_A_390_81#_c_1956_n 0.0103048f $X=2.035 $Y=2.735 $X2=0 $Y2=0
cc_407 N_D_c_461_n N_A_390_81#_c_1947_n 0.00298881f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_408 N_D_c_462_n N_A_390_81#_c_1947_n 0.00564096f $X=1.947 $Y=0.935 $X2=0
+ $Y2=0
cc_409 N_D_M1000_g N_A_390_81#_c_1958_n 0.00413459f $X=2.035 $Y=2.735 $X2=0
+ $Y2=0
cc_410 N_D_c_462_n N_VGND_c_2145_n 9.15902e-19 $X=1.947 $Y=0.935 $X2=0 $Y2=0
cc_411 N_D_c_460_n N_noxref_24_c_2273_n 0.00128684f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_412 N_D_c_461_n N_noxref_24_c_2273_n 0.0128576f $X=1.935 $Y=1.1 $X2=0 $Y2=0
cc_413 N_D_c_462_n N_noxref_24_c_2273_n 0.0119231f $X=1.947 $Y=0.935 $X2=0 $Y2=0
cc_414 N_D_c_462_n N_noxref_24_c_2274_n 0.00113655f $X=1.947 $Y=0.935 $X2=0
+ $Y2=0
cc_415 N_D_c_461_n noxref_25 0.00198619f $X=1.935 $Y=1.1 $X2=-0.19 $Y2=-0.245
cc_416 SCD N_RESET_B_c_917_n 0.00401365f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_417 N_SCD_c_506_n N_RESET_B_c_917_n 0.0207959f $X=3.04 $Y=1.645 $X2=0 $Y2=0
cc_418 N_SCD_M1035_g N_RESET_B_M1004_g 0.00851514f $X=3.05 $Y=0.615 $X2=0 $Y2=0
cc_419 N_SCD_M1035_g N_RESET_B_c_924_n 0.0247519f $X=3.05 $Y=0.615 $X2=0 $Y2=0
cc_420 N_SCD_M1039_g N_RESET_B_c_932_n 0.0283007f $X=3.035 $Y=2.735 $X2=0 $Y2=0
cc_421 N_SCD_c_504_n N_RESET_B_c_932_n 0.0207959f $X=3.04 $Y=1.985 $X2=0 $Y2=0
cc_422 N_SCD_M1039_g N_VPWR_c_1778_n 0.0140158f $X=3.035 $Y=2.735 $X2=0 $Y2=0
cc_423 N_SCD_M1039_g N_VPWR_c_1793_n 0.00543892f $X=3.035 $Y=2.735 $X2=0 $Y2=0
cc_424 N_SCD_M1039_g N_VPWR_c_1777_n 0.0053232f $X=3.035 $Y=2.735 $X2=0 $Y2=0
cc_425 N_SCD_M1039_g N_A_390_81#_c_1956_n 0.00198381f $X=3.035 $Y=2.735 $X2=0
+ $Y2=0
cc_426 N_SCD_M1035_g N_A_390_81#_c_1947_n 0.00753213f $X=3.05 $Y=0.615 $X2=0
+ $Y2=0
cc_427 N_SCD_M1039_g N_A_390_81#_c_1957_n 0.0137344f $X=3.035 $Y=2.735 $X2=0
+ $Y2=0
cc_428 N_SCD_c_509_n N_A_390_81#_c_1957_n 0.0033426f $X=3.04 $Y=2.15 $X2=0 $Y2=0
cc_429 SCD N_A_390_81#_c_1957_n 0.0232308f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_430 N_SCD_M1035_g N_A_390_81#_c_1948_n 0.0077301f $X=3.05 $Y=0.615 $X2=0
+ $Y2=0
cc_431 N_SCD_M1035_g N_A_390_81#_c_1949_n 0.00784052f $X=3.05 $Y=0.615 $X2=0
+ $Y2=0
cc_432 SCD N_A_390_81#_c_1949_n 0.0182587f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_433 N_SCD_c_506_n N_A_390_81#_c_1949_n 5.57115e-19 $X=3.04 $Y=1.645 $X2=0
+ $Y2=0
cc_434 N_SCD_M1035_g N_A_390_81#_c_1950_n 0.00328692f $X=3.05 $Y=0.615 $X2=0
+ $Y2=0
cc_435 SCD N_A_390_81#_c_1950_n 0.00853461f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_436 N_SCD_c_506_n N_A_390_81#_c_1950_n 0.00363171f $X=3.04 $Y=1.645 $X2=0
+ $Y2=0
cc_437 N_SCD_M1039_g N_A_390_81#_c_1951_n 0.00107151f $X=3.035 $Y=2.735 $X2=0
+ $Y2=0
cc_438 N_SCD_M1035_g N_A_390_81#_c_1951_n 9.9612e-19 $X=3.05 $Y=0.615 $X2=0
+ $Y2=0
cc_439 SCD N_A_390_81#_c_1951_n 0.0505537f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_440 N_SCD_c_506_n N_A_390_81#_c_1951_n 6.95935e-19 $X=3.04 $Y=1.645 $X2=0
+ $Y2=0
cc_441 N_SCD_M1035_g N_VGND_c_2145_n 9.15902e-19 $X=3.05 $Y=0.615 $X2=0 $Y2=0
cc_442 N_SCD_M1035_g N_noxref_24_c_2273_n 0.0118051f $X=3.05 $Y=0.615 $X2=0
+ $Y2=0
cc_443 N_CLK_c_555_n N_A_1037_119#_c_617_n 5.68491e-19 $X=4.565 $Y=1.41 $X2=0
+ $Y2=0
cc_444 N_CLK_M1027_g N_A_1037_119#_c_630_n 6.37144e-19 $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_445 CLK N_RESET_B_c_917_n 0.00394967f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_446 N_CLK_c_553_n N_RESET_B_c_917_n 0.021258f $X=3.94 $Y=1.445 $X2=0 $Y2=0
cc_447 N_CLK_c_555_n N_RESET_B_c_919_n 0.00984356f $X=4.565 $Y=1.41 $X2=0 $Y2=0
cc_448 CLK N_RESET_B_c_924_n 0.0022828f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_449 CLK N_RESET_B_c_933_n 0.00708182f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_450 N_CLK_M1027_g N_RESET_B_c_934_n 3.38591e-19 $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_451 CLK N_RESET_B_c_934_n 0.00451237f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_452 N_CLK_M1027_g N_RESET_B_c_938_n 0.00516734f $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_453 CLK N_RESET_B_c_938_n 0.00205192f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_454 N_CLK_c_553_n N_RESET_B_c_938_n 0.0201497f $X=3.94 $Y=1.445 $X2=0 $Y2=0
cc_455 N_CLK_c_551_n N_RESET_B_c_939_n 3.32348e-19 $X=4.395 $Y=1.51 $X2=0 $Y2=0
cc_456 N_CLK_M1027_g N_RESET_B_c_939_n 9.55661e-19 $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_457 CLK N_RESET_B_c_939_n 0.0290523f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_458 N_CLK_c_553_n N_RESET_B_c_939_n 3.82941e-19 $X=3.94 $Y=1.445 $X2=0 $Y2=0
cc_459 CLK N_A_837_119#_M1016_s 0.00682239f $X=3.995 $Y=1.21 $X2=-0.19
+ $Y2=-0.245
cc_460 CLK N_A_837_119#_c_1288_n 0.00331534f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_461 N_CLK_c_554_n N_A_837_119#_c_1288_n 0.00278435f $X=4.565 $Y=1.51 $X2=0
+ $Y2=0
cc_462 N_CLK_c_555_n N_A_837_119#_c_1288_n 0.00458006f $X=4.565 $Y=1.41 $X2=0
+ $Y2=0
cc_463 N_CLK_M1027_g N_A_837_119#_c_1291_n 0.0115693f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_464 CLK N_A_837_119#_c_1291_n 0.00402917f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_465 CLK N_A_837_119#_c_1267_n 0.0169963f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_466 N_CLK_c_554_n N_A_837_119#_c_1267_n 2.59598e-19 $X=4.565 $Y=1.51 $X2=0
+ $Y2=0
cc_467 N_CLK_c_555_n N_A_837_119#_c_1267_n 0.00229403f $X=4.565 $Y=1.41 $X2=0
+ $Y2=0
cc_468 N_CLK_M1027_g N_A_837_119#_c_1283_n 0.00263587f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_469 N_CLK_c_551_n N_A_837_119#_c_1268_n 0.00132107f $X=4.395 $Y=1.51 $X2=0
+ $Y2=0
cc_470 CLK N_A_837_119#_c_1268_n 0.0299511f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_471 N_CLK_c_555_n N_A_837_119#_c_1268_n 0.0133462f $X=4.565 $Y=1.41 $X2=0
+ $Y2=0
cc_472 N_CLK_c_551_n N_A_837_119#_c_1300_n 3.66206e-19 $X=4.395 $Y=1.51 $X2=0
+ $Y2=0
cc_473 N_CLK_M1027_g N_A_837_119#_c_1300_n 0.00439741f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_474 CLK N_A_837_119#_c_1300_n 0.0143178f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_475 N_CLK_c_554_n N_A_837_119#_c_1300_n 0.00103337f $X=4.565 $Y=1.51 $X2=0
+ $Y2=0
cc_476 CLK N_A_837_119#_c_1269_n 0.0273204f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_477 N_CLK_c_554_n N_A_837_119#_c_1269_n 0.00249677f $X=4.565 $Y=1.51 $X2=0
+ $Y2=0
cc_478 CLK N_A_837_119#_c_1270_n 2.99534e-19 $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_479 N_CLK_c_554_n N_A_837_119#_c_1270_n 0.0252665f $X=4.565 $Y=1.51 $X2=0
+ $Y2=0
cc_480 N_CLK_c_555_n N_A_837_119#_c_1271_n 0.0200837f $X=4.565 $Y=1.41 $X2=0
+ $Y2=0
cc_481 N_CLK_M1027_g N_A_837_119#_c_1286_n 0.0455485f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_482 N_CLK_M1027_g N_VPWR_c_1779_n 0.017461f $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_483 N_CLK_M1027_g N_VPWR_c_1786_n 0.00401239f $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_484 N_CLK_M1027_g N_VPWR_c_1777_n 0.00589267f $X=4.645 $Y=2.495 $X2=0 $Y2=0
cc_485 CLK N_A_390_81#_c_1949_n 0.0154252f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_486 CLK N_A_390_81#_c_1951_n 0.0273145f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_487 N_CLK_c_553_n N_A_390_81#_c_1951_n 0.00173026f $X=3.94 $Y=1.445 $X2=0
+ $Y2=0
cc_488 N_CLK_M1027_g N_A_390_81#_c_1960_n 0.0166738f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_489 N_CLK_M1027_g N_A_390_81#_c_1965_n 0.0147063f $X=4.645 $Y=2.495 $X2=0
+ $Y2=0
cc_490 CLK N_VGND_c_2138_n 0.0130346f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_491 N_CLK_c_553_n N_VGND_c_2138_n 0.00112289f $X=3.94 $Y=1.445 $X2=0 $Y2=0
cc_492 N_CLK_c_555_n N_VGND_c_2138_n 0.00335971f $X=4.565 $Y=1.41 $X2=0 $Y2=0
cc_493 N_CLK_c_555_n N_VGND_c_2139_n 0.00449587f $X=4.565 $Y=1.41 $X2=0 $Y2=0
cc_494 N_CLK_c_555_n N_VGND_c_2159_n 9.39239e-19 $X=4.565 $Y=1.41 $X2=0 $Y2=0
cc_495 N_A_1037_119#_c_623_n N_A_1383_349#_M1040_d 0.00256188f $X=9.09 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_496 N_A_1037_119#_c_612_n N_A_1383_349#_M1022_g 0.00668757f $X=6.695 $Y=1.355
+ $X2=0 $Y2=0
cc_497 N_A_1037_119#_M1032_g N_A_1383_349#_M1022_g 0.0522788f $X=6.695 $Y=0.805
+ $X2=0 $Y2=0
cc_498 N_A_1037_119#_c_622_n N_A_1383_349#_M1022_g 2.16281e-19 $X=8.25 $Y=0.665
+ $X2=0 $Y2=0
cc_499 N_A_1037_119#_c_631_n N_A_1383_349#_M1022_g 0.0124017f $X=7.135 $Y=0.365
+ $X2=0 $Y2=0
cc_500 N_A_1037_119#_M1032_g N_A_1383_349#_c_826_n 4.19365e-19 $X=6.695 $Y=0.805
+ $X2=0 $Y2=0
cc_501 N_A_1037_119#_M1002_g N_A_1383_349#_c_833_n 0.00260447f $X=6.135 $Y=2.495
+ $X2=0 $Y2=0
cc_502 N_A_1037_119#_c_612_n N_A_1383_349#_c_833_n 0.00193915f $X=6.695 $Y=1.355
+ $X2=0 $Y2=0
cc_503 N_A_1037_119#_c_632_n N_A_1383_349#_c_833_n 0.00175484f $X=6.065 $Y=1.682
+ $X2=0 $Y2=0
cc_504 N_A_1037_119#_c_622_n N_A_1383_349#_c_827_n 0.0713598f $X=8.25 $Y=0.665
+ $X2=0 $Y2=0
cc_505 N_A_1037_119#_c_623_n N_A_1383_349#_c_827_n 0.00354657f $X=9.09 $Y=0.34
+ $X2=0 $Y2=0
cc_506 N_A_1037_119#_M1032_g N_A_1383_349#_c_848_n 2.50187e-19 $X=6.695 $Y=0.805
+ $X2=0 $Y2=0
cc_507 N_A_1037_119#_c_622_n N_A_1383_349#_c_848_n 0.00488151f $X=8.25 $Y=0.665
+ $X2=0 $Y2=0
cc_508 N_A_1037_119#_c_631_n N_A_1383_349#_c_848_n 0.013158f $X=7.135 $Y=0.365
+ $X2=0 $Y2=0
cc_509 N_A_1037_119#_c_614_n N_A_1383_349#_c_828_n 0.00241408f $X=9.045 $Y=1.185
+ $X2=0 $Y2=0
cc_510 N_A_1037_119#_c_623_n N_A_1383_349#_c_828_n 0.0199132f $X=9.09 $Y=0.34
+ $X2=0 $Y2=0
cc_511 N_A_1037_119#_c_626_n N_A_1383_349#_c_828_n 0.0223601f $X=9.26 $Y=1.17
+ $X2=0 $Y2=0
cc_512 N_A_1037_119#_c_616_n N_A_1383_349#_c_835_n 0.00481612f $X=9.12 $Y=1.26
+ $X2=0 $Y2=0
cc_513 N_A_1037_119#_c_626_n N_A_1383_349#_c_835_n 0.0011706f $X=9.26 $Y=1.17
+ $X2=0 $Y2=0
cc_514 N_A_1037_119#_c_628_n N_A_1383_349#_c_835_n 0.0036935f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_515 N_A_1037_119#_c_616_n N_A_1383_349#_c_829_n 0.00241408f $X=9.12 $Y=1.26
+ $X2=0 $Y2=0
cc_516 N_A_1037_119#_M1032_g N_RESET_B_c_919_n 0.00881316f $X=6.695 $Y=0.805
+ $X2=0 $Y2=0
cc_517 N_A_1037_119#_c_619_n N_RESET_B_c_919_n 0.0323956f $X=7.015 $Y=0.365
+ $X2=0 $Y2=0
cc_518 N_A_1037_119#_c_620_n N_RESET_B_c_919_n 0.00590986f $X=5.42 $Y=0.365
+ $X2=0 $Y2=0
cc_519 N_A_1037_119#_c_622_n N_RESET_B_c_919_n 0.0010205f $X=8.25 $Y=0.665 $X2=0
+ $Y2=0
cc_520 N_A_1037_119#_c_631_n N_RESET_B_c_919_n 0.00338531f $X=7.135 $Y=0.365
+ $X2=0 $Y2=0
cc_521 N_A_1037_119#_c_622_n N_RESET_B_M1007_g 0.0127125f $X=8.25 $Y=0.665 $X2=0
+ $Y2=0
cc_522 N_A_1037_119#_c_624_n N_RESET_B_M1007_g 5.42284e-19 $X=8.42 $Y=0.34 $X2=0
+ $Y2=0
cc_523 N_A_1037_119#_c_631_n N_RESET_B_M1007_g 0.00797906f $X=7.135 $Y=0.365
+ $X2=0 $Y2=0
cc_524 N_A_1037_119#_M1002_g N_RESET_B_c_933_n 0.00529886f $X=6.135 $Y=2.495
+ $X2=0 $Y2=0
cc_525 N_A_1037_119#_c_611_n N_RESET_B_c_933_n 0.00476221f $X=6.47 $Y=1.682
+ $X2=0 $Y2=0
cc_526 N_A_1037_119#_c_612_n N_RESET_B_c_933_n 6.19028e-19 $X=6.695 $Y=1.355
+ $X2=0 $Y2=0
cc_527 N_A_1037_119#_c_621_n N_RESET_B_c_933_n 0.0164042f $X=6.065 $Y=1.8 $X2=0
+ $Y2=0
cc_528 N_A_1037_119#_c_630_n N_RESET_B_c_933_n 0.0340128f $X=5.387 $Y=1.8 $X2=0
+ $Y2=0
cc_529 N_A_1037_119#_c_632_n N_RESET_B_c_933_n 0.00570083f $X=6.065 $Y=1.682
+ $X2=0 $Y2=0
cc_530 N_A_1037_119#_c_615_n N_RESET_B_c_935_n 4.12125e-19 $X=9.48 $Y=1.26 $X2=0
+ $Y2=0
cc_531 N_A_1037_119#_c_628_n N_RESET_B_c_935_n 0.0178906f $X=9.95 $Y=2.165 $X2=0
+ $Y2=0
cc_532 N_A_1037_119#_c_641_n N_RESET_B_c_935_n 0.00339488f $X=10.11 $Y=2.165
+ $X2=0 $Y2=0
cc_533 N_A_1037_119#_c_614_n N_A_1235_119#_M1040_g 0.0131362f $X=9.045 $Y=1.185
+ $X2=0 $Y2=0
cc_534 N_A_1037_119#_c_623_n N_A_1235_119#_M1040_g 0.0120273f $X=9.09 $Y=0.34
+ $X2=0 $Y2=0
cc_535 N_A_1037_119#_c_684_p N_A_1235_119#_M1040_g 6.7135e-19 $X=9.175 $Y=1.005
+ $X2=0 $Y2=0
cc_536 N_A_1037_119#_c_616_n N_A_1235_119#_c_1139_n 0.0131362f $X=9.12 $Y=1.26
+ $X2=0 $Y2=0
cc_537 N_A_1037_119#_M1002_g N_A_1235_119#_c_1148_n 0.00402175f $X=6.135
+ $Y=2.495 $X2=0 $Y2=0
cc_538 N_A_1037_119#_c_611_n N_A_1235_119#_c_1148_n 4.35859e-19 $X=6.47 $Y=1.682
+ $X2=0 $Y2=0
cc_539 N_A_1037_119#_c_612_n N_A_1235_119#_c_1148_n 5.25936e-19 $X=6.695
+ $Y=1.355 $X2=0 $Y2=0
cc_540 N_A_1037_119#_M1002_g N_A_1235_119#_c_1140_n 2.50724e-19 $X=6.135
+ $Y=2.495 $X2=0 $Y2=0
cc_541 N_A_1037_119#_c_612_n N_A_1235_119#_c_1140_n 0.00821458f $X=6.695
+ $Y=1.355 $X2=0 $Y2=0
cc_542 N_A_1037_119#_M1032_g N_A_1235_119#_c_1140_n 0.0058207f $X=6.695 $Y=0.805
+ $X2=0 $Y2=0
cc_543 N_A_1037_119#_c_611_n N_A_1235_119#_c_1144_n 5.35933e-19 $X=6.47 $Y=1.682
+ $X2=0 $Y2=0
cc_544 N_A_1037_119#_c_612_n N_A_1235_119#_c_1144_n 0.00406521f $X=6.695
+ $Y=1.355 $X2=0 $Y2=0
cc_545 N_A_1037_119#_M1032_g N_A_1235_119#_c_1144_n 0.0163191f $X=6.695 $Y=0.805
+ $X2=0 $Y2=0
cc_546 N_A_1037_119#_c_619_n N_A_1235_119#_c_1144_n 0.029146f $X=7.015 $Y=0.365
+ $X2=0 $Y2=0
cc_547 N_A_1037_119#_c_631_n N_A_1235_119#_c_1144_n 0.00412857f $X=7.135
+ $Y=0.365 $X2=0 $Y2=0
cc_548 N_A_1037_119#_c_618_n N_A_837_119#_c_1256_n 0.00683949f $X=5.502 $Y=1.635
+ $X2=0 $Y2=0
cc_549 N_A_1037_119#_c_618_n N_A_837_119#_c_1257_n 0.00398951f $X=5.502 $Y=1.635
+ $X2=0 $Y2=0
cc_550 N_A_1037_119#_M1002_g N_A_837_119#_c_1272_n 0.0140717f $X=6.135 $Y=2.495
+ $X2=0 $Y2=0
cc_551 N_A_1037_119#_c_621_n N_A_837_119#_c_1272_n 2.83568e-19 $X=6.065 $Y=1.8
+ $X2=0 $Y2=0
cc_552 N_A_1037_119#_c_630_n N_A_837_119#_c_1272_n 0.00273999f $X=5.387 $Y=1.8
+ $X2=0 $Y2=0
cc_553 N_A_1037_119#_c_619_n N_A_837_119#_c_1258_n 6.93569e-19 $X=7.015 $Y=0.365
+ $X2=0 $Y2=0
cc_554 N_A_1037_119#_c_621_n N_A_837_119#_c_1258_n 0.00390284f $X=6.065 $Y=1.8
+ $X2=0 $Y2=0
cc_555 N_A_1037_119#_c_632_n N_A_837_119#_c_1258_n 0.00919512f $X=6.065 $Y=1.682
+ $X2=0 $Y2=0
cc_556 N_A_1037_119#_c_618_n N_A_837_119#_c_1259_n 5.88192e-19 $X=5.502 $Y=1.635
+ $X2=0 $Y2=0
cc_557 N_A_1037_119#_c_619_n N_A_837_119#_c_1259_n 0.00440089f $X=7.015 $Y=0.365
+ $X2=0 $Y2=0
cc_558 N_A_1037_119#_c_629_n N_A_837_119#_c_1259_n 0.00626502f $X=5.32 $Y=1.11
+ $X2=0 $Y2=0
cc_559 N_A_1037_119#_M1002_g N_A_837_119#_c_1274_n 0.0107342f $X=6.135 $Y=2.495
+ $X2=0 $Y2=0
cc_560 N_A_1037_119#_M1032_g N_A_837_119#_c_1260_n 0.0141831f $X=6.695 $Y=0.805
+ $X2=0 $Y2=0
cc_561 N_A_1037_119#_c_617_n N_A_837_119#_c_1260_n 0.00388823f $X=5.32 $Y=0.74
+ $X2=0 $Y2=0
cc_562 N_A_1037_119#_c_619_n N_A_837_119#_c_1260_n 0.00241808f $X=7.015 $Y=0.365
+ $X2=0 $Y2=0
cc_563 N_A_1037_119#_c_629_n N_A_837_119#_c_1260_n 4.05093e-19 $X=5.32 $Y=1.11
+ $X2=0 $Y2=0
cc_564 N_A_1037_119#_M1002_g N_A_837_119#_M1025_g 0.0153886f $X=6.135 $Y=2.495
+ $X2=0 $Y2=0
cc_565 N_A_1037_119#_c_612_n N_A_837_119#_M1025_g 0.00635016f $X=6.695 $Y=1.355
+ $X2=0 $Y2=0
cc_566 N_A_1037_119#_M1021_g N_A_837_119#_M1020_g 0.00652156f $X=10.11 $Y=2.75
+ $X2=0 $Y2=0
cc_567 N_A_1037_119#_c_628_n N_A_837_119#_M1020_g 0.00195755f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_568 N_A_1037_119#_c_627_n N_A_837_119#_c_1261_n 0.0170653f $X=9.645 $Y=1.17
+ $X2=0 $Y2=0
cc_569 N_A_1037_119#_c_628_n N_A_837_119#_c_1261_n 0.0202931f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_570 N_A_1037_119#_c_641_n N_A_837_119#_c_1261_n 0.0207799f $X=10.11 $Y=2.165
+ $X2=0 $Y2=0
cc_571 N_A_1037_119#_c_615_n N_A_837_119#_c_1280_n 0.0170653f $X=9.48 $Y=1.26
+ $X2=0 $Y2=0
cc_572 N_A_1037_119#_c_625_n N_A_837_119#_c_1280_n 0.00273345f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_573 N_A_1037_119#_c_626_n N_A_837_119#_c_1280_n 6.76091e-19 $X=9.26 $Y=1.17
+ $X2=0 $Y2=0
cc_574 N_A_1037_119#_c_628_n N_A_837_119#_c_1262_n 0.00569302f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_575 N_A_1037_119#_c_618_n N_A_837_119#_c_1264_n 0.00530144f $X=5.502 $Y=1.635
+ $X2=0 $Y2=0
cc_576 N_A_1037_119#_M1002_g N_A_837_119#_c_1265_n 0.00780637f $X=6.135 $Y=2.495
+ $X2=0 $Y2=0
cc_577 N_A_1037_119#_c_618_n N_A_837_119#_c_1265_n 0.0025296f $X=5.502 $Y=1.635
+ $X2=0 $Y2=0
cc_578 N_A_1037_119#_c_621_n N_A_837_119#_c_1265_n 0.00887481f $X=6.065 $Y=1.8
+ $X2=0 $Y2=0
cc_579 N_A_1037_119#_c_630_n N_A_837_119#_c_1265_n 0.0137747f $X=5.387 $Y=1.8
+ $X2=0 $Y2=0
cc_580 N_A_1037_119#_c_632_n N_A_837_119#_c_1265_n 0.0236278f $X=6.065 $Y=1.682
+ $X2=0 $Y2=0
cc_581 N_A_1037_119#_c_625_n N_A_837_119#_c_1266_n 0.00289132f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_582 N_A_1037_119#_c_627_n N_A_837_119#_c_1266_n 0.0181127f $X=9.645 $Y=1.17
+ $X2=0 $Y2=0
cc_583 N_A_1037_119#_c_630_n N_A_837_119#_c_1291_n 0.00844482f $X=5.387 $Y=1.8
+ $X2=0 $Y2=0
cc_584 N_A_1037_119#_c_618_n N_A_837_119#_c_1267_n 0.00670366f $X=5.502 $Y=1.635
+ $X2=0 $Y2=0
cc_585 N_A_1037_119#_c_630_n N_A_837_119#_c_1283_n 0.00732766f $X=5.387 $Y=1.8
+ $X2=0 $Y2=0
cc_586 N_A_1037_119#_c_617_n N_A_837_119#_c_1268_n 0.00435847f $X=5.32 $Y=0.74
+ $X2=0 $Y2=0
cc_587 N_A_1037_119#_c_630_n N_A_837_119#_c_1300_n 0.00445803f $X=5.387 $Y=1.8
+ $X2=0 $Y2=0
cc_588 N_A_1037_119#_c_618_n N_A_837_119#_c_1269_n 0.0143607f $X=5.502 $Y=1.635
+ $X2=0 $Y2=0
cc_589 N_A_1037_119#_c_629_n N_A_837_119#_c_1269_n 0.002722f $X=5.32 $Y=1.11
+ $X2=0 $Y2=0
cc_590 N_A_1037_119#_c_630_n N_A_837_119#_c_1269_n 0.0148843f $X=5.387 $Y=1.8
+ $X2=0 $Y2=0
cc_591 N_A_1037_119#_c_618_n N_A_837_119#_c_1270_n 5.05397e-19 $X=5.502 $Y=1.635
+ $X2=0 $Y2=0
cc_592 N_A_1037_119#_c_629_n N_A_837_119#_c_1270_n 0.00513697f $X=5.32 $Y=1.11
+ $X2=0 $Y2=0
cc_593 N_A_1037_119#_c_630_n N_A_837_119#_c_1270_n 0.00611889f $X=5.387 $Y=1.8
+ $X2=0 $Y2=0
cc_594 N_A_1037_119#_c_617_n N_A_837_119#_c_1271_n 0.00832061f $X=5.32 $Y=0.74
+ $X2=0 $Y2=0
cc_595 N_A_1037_119#_c_618_n N_A_837_119#_c_1271_n 0.00129839f $X=5.502 $Y=1.635
+ $X2=0 $Y2=0
cc_596 N_A_1037_119#_c_629_n N_A_837_119#_c_1271_n 0.00399071f $X=5.32 $Y=1.11
+ $X2=0 $Y2=0
cc_597 N_A_1037_119#_c_630_n N_A_837_119#_c_1286_n 0.0061722f $X=5.387 $Y=1.8
+ $X2=0 $Y2=0
cc_598 N_A_1037_119#_M1021_g N_A_2082_446#_M1005_g 0.0254895f $X=10.11 $Y=2.75
+ $X2=0 $Y2=0
cc_599 N_A_1037_119#_c_641_n N_A_2082_446#_c_1469_n 0.0254895f $X=10.11 $Y=2.165
+ $X2=0 $Y2=0
cc_600 N_A_1037_119#_c_641_n N_A_2082_446#_c_1460_n 0.0127423f $X=10.11 $Y=2.165
+ $X2=0 $Y2=0
cc_601 N_A_1037_119#_c_623_n N_A_1824_74#_M1028_d 0.00248108f $X=9.09 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_602 N_A_1037_119#_c_684_p N_A_1824_74#_M1028_d 0.0130256f $X=9.175 $Y=1.005
+ $X2=-0.19 $Y2=-0.245
cc_603 N_A_1037_119#_c_625_n N_A_1824_74#_M1028_d 0.00450592f $X=9.785 $Y=1.17
+ $X2=-0.19 $Y2=-0.245
cc_604 N_A_1037_119#_M1021_g N_A_1824_74#_c_1601_n 0.0018001f $X=10.11 $Y=2.75
+ $X2=0 $Y2=0
cc_605 N_A_1037_119#_c_625_n N_A_1824_74#_c_1601_n 0.00858049f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_606 N_A_1037_119#_c_628_n N_A_1824_74#_c_1601_n 0.0339542f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_607 N_A_1037_119#_c_641_n N_A_1824_74#_c_1601_n 0.00257809f $X=10.11 $Y=2.165
+ $X2=0 $Y2=0
cc_608 N_A_1037_119#_c_614_n N_A_1824_74#_c_1585_n 0.0018748f $X=9.045 $Y=1.185
+ $X2=0 $Y2=0
cc_609 N_A_1037_119#_c_615_n N_A_1824_74#_c_1585_n 2.42458e-19 $X=9.48 $Y=1.26
+ $X2=0 $Y2=0
cc_610 N_A_1037_119#_c_684_p N_A_1824_74#_c_1585_n 0.026719f $X=9.175 $Y=1.005
+ $X2=0 $Y2=0
cc_611 N_A_1037_119#_c_625_n N_A_1824_74#_c_1585_n 0.0466861f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_612 N_A_1037_119#_c_627_n N_A_1824_74#_c_1585_n 0.0070276f $X=9.645 $Y=1.17
+ $X2=0 $Y2=0
cc_613 N_A_1037_119#_M1021_g N_A_1824_74#_c_1595_n 0.014429f $X=10.11 $Y=2.75
+ $X2=0 $Y2=0
cc_614 N_A_1037_119#_c_628_n N_A_1824_74#_c_1595_n 0.0189574f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_615 N_A_1037_119#_c_641_n N_A_1824_74#_c_1595_n 0.00170014f $X=10.11 $Y=2.165
+ $X2=0 $Y2=0
cc_616 N_A_1037_119#_c_625_n N_A_1824_74#_c_1586_n 0.00187033f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_617 N_A_1037_119#_c_625_n N_A_1824_74#_c_1587_n 0.0107493f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_618 N_A_1037_119#_c_628_n N_A_1824_74#_c_1587_n 0.0746733f $X=9.95 $Y=2.165
+ $X2=0 $Y2=0
cc_619 N_A_1037_119#_c_641_n N_A_1824_74#_c_1587_n 0.00480077f $X=10.11 $Y=2.165
+ $X2=0 $Y2=0
cc_620 N_A_1037_119#_c_625_n N_A_1824_74#_c_1589_n 0.0146626f $X=9.785 $Y=1.17
+ $X2=0 $Y2=0
cc_621 N_A_1037_119#_M1021_g N_VPWR_c_1795_n 0.00370063f $X=10.11 $Y=2.75 $X2=0
+ $Y2=0
cc_622 N_A_1037_119#_M1021_g N_VPWR_c_1801_n 0.00125493f $X=10.11 $Y=2.75 $X2=0
+ $Y2=0
cc_623 N_A_1037_119#_M1002_g N_VPWR_c_1777_n 0.00113998f $X=6.135 $Y=2.495 $X2=0
+ $Y2=0
cc_624 N_A_1037_119#_M1021_g N_VPWR_c_1777_n 0.00455976f $X=10.11 $Y=2.75 $X2=0
+ $Y2=0
cc_625 N_A_1037_119#_M1034_d N_A_390_81#_c_1960_n 0.00583079f $X=5.185 $Y=1.935
+ $X2=0 $Y2=0
cc_626 N_A_1037_119#_c_621_n N_A_390_81#_c_1960_n 0.00200754f $X=6.065 $Y=1.8
+ $X2=0 $Y2=0
cc_627 N_A_1037_119#_c_630_n N_A_390_81#_c_1960_n 0.0278382f $X=5.387 $Y=1.8
+ $X2=0 $Y2=0
cc_628 N_A_1037_119#_M1002_g N_A_390_81#_c_1961_n 2.76323e-19 $X=6.135 $Y=2.495
+ $X2=0 $Y2=0
cc_629 N_A_1037_119#_M1032_g N_A_390_81#_c_1952_n 0.00145669f $X=6.695 $Y=0.805
+ $X2=0 $Y2=0
cc_630 N_A_1037_119#_c_617_n N_A_390_81#_c_1952_n 0.0119409f $X=5.32 $Y=0.74
+ $X2=0 $Y2=0
cc_631 N_A_1037_119#_c_618_n N_A_390_81#_c_1952_n 0.00559071f $X=5.502 $Y=1.635
+ $X2=0 $Y2=0
cc_632 N_A_1037_119#_c_619_n N_A_390_81#_c_1952_n 0.0214205f $X=7.015 $Y=0.365
+ $X2=0 $Y2=0
cc_633 N_A_1037_119#_c_629_n N_A_390_81#_c_1952_n 0.0219181f $X=5.32 $Y=1.11
+ $X2=0 $Y2=0
cc_634 N_A_1037_119#_M1002_g N_A_390_81#_c_1962_n 0.0165116f $X=6.135 $Y=2.495
+ $X2=0 $Y2=0
cc_635 N_A_1037_119#_c_611_n N_A_390_81#_c_1962_n 0.00260156f $X=6.47 $Y=1.682
+ $X2=0 $Y2=0
cc_636 N_A_1037_119#_c_621_n N_A_390_81#_c_1962_n 0.00952002f $X=6.065 $Y=1.8
+ $X2=0 $Y2=0
cc_637 N_A_1037_119#_c_632_n N_A_390_81#_c_1962_n 9.74074e-19 $X=6.065 $Y=1.682
+ $X2=0 $Y2=0
cc_638 N_A_1037_119#_c_621_n N_A_390_81#_c_1963_n 0.0166792f $X=6.065 $Y=1.8
+ $X2=0 $Y2=0
cc_639 N_A_1037_119#_c_630_n N_A_390_81#_c_1963_n 0.0120217f $X=5.387 $Y=1.8
+ $X2=0 $Y2=0
cc_640 N_A_1037_119#_c_632_n N_A_390_81#_c_1963_n 0.00171449f $X=6.065 $Y=1.682
+ $X2=0 $Y2=0
cc_641 N_A_1037_119#_c_612_n N_A_390_81#_c_1953_n 0.00565997f $X=6.695 $Y=1.355
+ $X2=0 $Y2=0
cc_642 N_A_1037_119#_M1032_g N_A_390_81#_c_1953_n 0.00130392f $X=6.695 $Y=0.805
+ $X2=0 $Y2=0
cc_643 N_A_1037_119#_c_621_n N_A_390_81#_c_1953_n 0.00358942f $X=6.065 $Y=1.8
+ $X2=0 $Y2=0
cc_644 N_A_1037_119#_c_632_n N_A_390_81#_c_1953_n 0.00590575f $X=6.065 $Y=1.682
+ $X2=0 $Y2=0
cc_645 N_A_1037_119#_c_618_n N_A_390_81#_c_1954_n 0.0139746f $X=5.502 $Y=1.635
+ $X2=0 $Y2=0
cc_646 N_A_1037_119#_c_621_n N_A_390_81#_c_1954_n 0.0268006f $X=6.065 $Y=1.8
+ $X2=0 $Y2=0
cc_647 N_A_1037_119#_c_632_n N_A_390_81#_c_1954_n 0.00197058f $X=6.065 $Y=1.682
+ $X2=0 $Y2=0
cc_648 N_A_1037_119#_M1002_g N_A_390_81#_c_1955_n 0.00366452f $X=6.135 $Y=2.495
+ $X2=0 $Y2=0
cc_649 N_A_1037_119#_c_611_n N_A_390_81#_c_1955_n 0.00995261f $X=6.47 $Y=1.682
+ $X2=0 $Y2=0
cc_650 N_A_1037_119#_c_612_n N_A_390_81#_c_1955_n 0.00766644f $X=6.695 $Y=1.355
+ $X2=0 $Y2=0
cc_651 N_A_1037_119#_c_621_n N_A_390_81#_c_1955_n 0.0230519f $X=6.065 $Y=1.8
+ $X2=0 $Y2=0
cc_652 N_A_1037_119#_c_632_n N_A_390_81#_c_1955_n 0.00213027f $X=6.065 $Y=1.682
+ $X2=0 $Y2=0
cc_653 N_A_1037_119#_c_622_n N_VGND_M1007_d 0.0214581f $X=8.25 $Y=0.665 $X2=0
+ $Y2=0
cc_654 N_A_1037_119#_c_803_p N_VGND_M1007_d 0.00612573f $X=8.335 $Y=0.58 $X2=0
+ $Y2=0
cc_655 N_A_1037_119#_c_624_n N_VGND_M1007_d 8.42533e-19 $X=8.42 $Y=0.34 $X2=0
+ $Y2=0
cc_656 N_A_1037_119#_c_617_n N_VGND_c_2139_n 0.0153892f $X=5.32 $Y=0.74 $X2=0
+ $Y2=0
cc_657 N_A_1037_119#_c_620_n N_VGND_c_2139_n 0.0173959f $X=5.42 $Y=0.365 $X2=0
+ $Y2=0
cc_658 N_A_1037_119#_c_619_n N_VGND_c_2150_n 0.0977364f $X=7.015 $Y=0.365 $X2=0
+ $Y2=0
cc_659 N_A_1037_119#_c_620_n N_VGND_c_2150_n 0.0168491f $X=5.42 $Y=0.365 $X2=0
+ $Y2=0
cc_660 N_A_1037_119#_c_622_n N_VGND_c_2150_n 0.0423632f $X=8.25 $Y=0.665 $X2=0
+ $Y2=0
cc_661 N_A_1037_119#_c_624_n N_VGND_c_2150_n 0.0139413f $X=8.42 $Y=0.34 $X2=0
+ $Y2=0
cc_662 N_A_1037_119#_c_631_n N_VGND_c_2150_n 0.0229767f $X=7.135 $Y=0.365 $X2=0
+ $Y2=0
cc_663 N_A_1037_119#_c_614_n N_VGND_c_2151_n 0.00278242f $X=9.045 $Y=1.185 $X2=0
+ $Y2=0
cc_664 N_A_1037_119#_c_622_n N_VGND_c_2151_n 0.00335833f $X=8.25 $Y=0.665 $X2=0
+ $Y2=0
cc_665 N_A_1037_119#_c_623_n N_VGND_c_2151_n 0.0544002f $X=9.09 $Y=0.34 $X2=0
+ $Y2=0
cc_666 N_A_1037_119#_c_624_n N_VGND_c_2151_n 0.0118998f $X=8.42 $Y=0.34 $X2=0
+ $Y2=0
cc_667 N_A_1037_119#_c_614_n N_VGND_c_2159_n 0.00359177f $X=9.045 $Y=1.185 $X2=0
+ $Y2=0
cc_668 N_A_1037_119#_c_619_n N_VGND_c_2159_n 0.0534591f $X=7.015 $Y=0.365 $X2=0
+ $Y2=0
cc_669 N_A_1037_119#_c_620_n N_VGND_c_2159_n 0.00867614f $X=5.42 $Y=0.365 $X2=0
+ $Y2=0
cc_670 N_A_1037_119#_c_622_n N_VGND_c_2159_n 0.0165948f $X=8.25 $Y=0.665 $X2=0
+ $Y2=0
cc_671 N_A_1037_119#_c_623_n N_VGND_c_2159_n 0.0304263f $X=9.09 $Y=0.34 $X2=0
+ $Y2=0
cc_672 N_A_1037_119#_c_624_n N_VGND_c_2159_n 0.00655543f $X=8.42 $Y=0.34 $X2=0
+ $Y2=0
cc_673 N_A_1037_119#_c_631_n N_VGND_c_2159_n 0.00817719f $X=7.135 $Y=0.365 $X2=0
+ $Y2=0
cc_674 N_A_1037_119#_c_622_n A_1432_119# 0.00130131f $X=8.25 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_675 N_A_1037_119#_c_631_n A_1432_119# 7.74822e-19 $X=7.135 $Y=0.365 $X2=-0.19
+ $Y2=-0.245
cc_676 N_A_1383_349#_M1022_g N_RESET_B_c_919_n 0.00880383f $X=7.085 $Y=0.805
+ $X2=0 $Y2=0
cc_677 N_A_1383_349#_M1022_g N_RESET_B_M1007_g 0.0465693f $X=7.085 $Y=0.805
+ $X2=0 $Y2=0
cc_678 N_A_1383_349#_c_826_n N_RESET_B_M1007_g 0.00474717f $X=7.165 $Y=1.91
+ $X2=0 $Y2=0
cc_679 N_A_1383_349#_c_827_n N_RESET_B_M1007_g 0.0144265f $X=8.59 $Y=1.005 $X2=0
+ $Y2=0
cc_680 N_A_1383_349#_M1022_g N_RESET_B_c_922_n 0.0108937f $X=7.085 $Y=0.805
+ $X2=0 $Y2=0
cc_681 N_A_1383_349#_c_826_n N_RESET_B_c_922_n 0.00131101f $X=7.165 $Y=1.91
+ $X2=0 $Y2=0
cc_682 N_A_1383_349#_c_833_n N_RESET_B_c_922_n 0.00263372f $X=7.165 $Y=1.91
+ $X2=0 $Y2=0
cc_683 N_A_1383_349#_c_827_n N_RESET_B_c_925_n 0.00473252f $X=8.59 $Y=1.005
+ $X2=0 $Y2=0
cc_684 N_A_1383_349#_M1033_g N_RESET_B_c_933_n 0.00229321f $X=7.005 $Y=2.495
+ $X2=0 $Y2=0
cc_685 N_A_1383_349#_c_826_n N_RESET_B_c_933_n 0.0210957f $X=7.165 $Y=1.91 $X2=0
+ $Y2=0
cc_686 N_A_1383_349#_c_833_n N_RESET_B_c_933_n 0.00910947f $X=7.165 $Y=1.91
+ $X2=0 $Y2=0
cc_687 N_A_1383_349#_M1006_d N_RESET_B_c_935_n 0.00448801f $X=8.73 $Y=1.735
+ $X2=0 $Y2=0
cc_688 N_A_1383_349#_c_834_n N_RESET_B_c_935_n 0.0436783f $X=8.95 $Y=2.235 $X2=0
+ $Y2=0
cc_689 N_A_1383_349#_c_834_n N_RESET_B_c_936_n 0.00263797f $X=8.95 $Y=2.235
+ $X2=0 $Y2=0
cc_690 N_A_1383_349#_c_834_n N_RESET_B_c_937_n 0.00493501f $X=8.95 $Y=2.235
+ $X2=0 $Y2=0
cc_691 N_A_1383_349#_M1033_g N_RESET_B_c_940_n 0.0169494f $X=7.005 $Y=2.495
+ $X2=0 $Y2=0
cc_692 N_A_1383_349#_c_826_n N_RESET_B_c_940_n 3.6329e-19 $X=7.165 $Y=1.91 $X2=0
+ $Y2=0
cc_693 N_A_1383_349#_c_833_n N_RESET_B_c_940_n 0.0183362f $X=7.165 $Y=1.91 $X2=0
+ $Y2=0
cc_694 N_A_1383_349#_c_827_n N_A_1235_119#_M1040_g 0.0149183f $X=8.59 $Y=1.005
+ $X2=0 $Y2=0
cc_695 N_A_1383_349#_c_828_n N_A_1235_119#_M1040_g 0.0150489f $X=8.755 $Y=0.86
+ $X2=0 $Y2=0
cc_696 N_A_1383_349#_c_829_n N_A_1235_119#_M1040_g 0.00617118f $X=8.932 $Y=1.715
+ $X2=0 $Y2=0
cc_697 N_A_1383_349#_c_835_n N_A_1235_119#_M1006_g 0.00832071f $X=8.95 $Y=1.88
+ $X2=0 $Y2=0
cc_698 N_A_1383_349#_c_827_n N_A_1235_119#_c_1138_n 0.00840745f $X=8.59 $Y=1.005
+ $X2=0 $Y2=0
cc_699 N_A_1383_349#_c_828_n N_A_1235_119#_c_1139_n 0.00470883f $X=8.755 $Y=0.86
+ $X2=0 $Y2=0
cc_700 N_A_1383_349#_c_829_n N_A_1235_119#_c_1139_n 0.00832071f $X=8.932
+ $Y=1.715 $X2=0 $Y2=0
cc_701 N_A_1383_349#_M1022_g N_A_1235_119#_c_1140_n 0.0036446f $X=7.085 $Y=0.805
+ $X2=0 $Y2=0
cc_702 N_A_1383_349#_c_826_n N_A_1235_119#_c_1140_n 0.0696484f $X=7.165 $Y=1.91
+ $X2=0 $Y2=0
cc_703 N_A_1383_349#_c_833_n N_A_1235_119#_c_1140_n 0.00708991f $X=7.165 $Y=1.91
+ $X2=0 $Y2=0
cc_704 N_A_1383_349#_M1033_g N_A_1235_119#_c_1177_n 0.0115346f $X=7.005 $Y=2.495
+ $X2=0 $Y2=0
cc_705 N_A_1383_349#_c_826_n N_A_1235_119#_c_1177_n 0.0101422f $X=7.165 $Y=1.91
+ $X2=0 $Y2=0
cc_706 N_A_1383_349#_c_833_n N_A_1235_119#_c_1177_n 0.00173802f $X=7.165 $Y=1.91
+ $X2=0 $Y2=0
cc_707 N_A_1383_349#_M1033_g N_A_1235_119#_c_1141_n 0.00248668f $X=7.005
+ $Y=2.495 $X2=0 $Y2=0
cc_708 N_A_1383_349#_M1022_g N_A_1235_119#_c_1141_n 4.10299e-19 $X=7.085
+ $Y=0.805 $X2=0 $Y2=0
cc_709 N_A_1383_349#_c_826_n N_A_1235_119#_c_1141_n 0.0370159f $X=7.165 $Y=1.91
+ $X2=0 $Y2=0
cc_710 N_A_1383_349#_c_833_n N_A_1235_119#_c_1141_n 0.00171792f $X=7.165 $Y=1.91
+ $X2=0 $Y2=0
cc_711 N_A_1383_349#_M1022_g N_A_1235_119#_c_1142_n 7.98464e-19 $X=7.085
+ $Y=0.805 $X2=0 $Y2=0
cc_712 N_A_1383_349#_c_826_n N_A_1235_119#_c_1142_n 0.0271618f $X=7.165 $Y=1.91
+ $X2=0 $Y2=0
cc_713 N_A_1383_349#_c_827_n N_A_1235_119#_c_1142_n 0.0133025f $X=8.59 $Y=1.005
+ $X2=0 $Y2=0
cc_714 N_A_1383_349#_c_827_n N_A_1235_119#_c_1143_n 0.0573215f $X=8.59 $Y=1.005
+ $X2=0 $Y2=0
cc_715 N_A_1383_349#_c_829_n N_A_1235_119#_c_1143_n 0.0151715f $X=8.932 $Y=1.715
+ $X2=0 $Y2=0
cc_716 N_A_1383_349#_M1022_g N_A_1235_119#_c_1144_n 0.00225945f $X=7.085
+ $Y=0.805 $X2=0 $Y2=0
cc_717 N_A_1383_349#_c_826_n N_A_1235_119#_c_1144_n 0.00282944f $X=7.165 $Y=1.91
+ $X2=0 $Y2=0
cc_718 N_A_1383_349#_c_848_n N_A_1235_119#_c_1144_n 0.0131612f $X=7.315 $Y=1.005
+ $X2=0 $Y2=0
cc_719 N_A_1383_349#_M1033_g N_A_1235_119#_c_1151_n 9.66315e-19 $X=7.005
+ $Y=2.495 $X2=0 $Y2=0
cc_720 N_A_1383_349#_M1033_g N_A_837_119#_M1025_g 0.0375552f $X=7.005 $Y=2.495
+ $X2=0 $Y2=0
cc_721 N_A_1383_349#_M1033_g N_A_837_119#_c_1277_n 0.0103493f $X=7.005 $Y=2.495
+ $X2=0 $Y2=0
cc_722 N_A_1383_349#_c_834_n N_A_837_119#_c_1277_n 0.00668309f $X=8.95 $Y=2.235
+ $X2=0 $Y2=0
cc_723 N_A_1383_349#_c_834_n N_A_837_119#_M1020_g 0.00399773f $X=8.95 $Y=2.235
+ $X2=0 $Y2=0
cc_724 N_A_1383_349#_c_835_n N_A_837_119#_c_1280_n 0.00399773f $X=8.95 $Y=1.88
+ $X2=0 $Y2=0
cc_725 N_A_1383_349#_c_829_n N_A_837_119#_c_1280_n 0.00306438f $X=8.932 $Y=1.715
+ $X2=0 $Y2=0
cc_726 N_A_1383_349#_c_834_n N_A_1824_74#_c_1601_n 0.0227868f $X=8.95 $Y=2.235
+ $X2=0 $Y2=0
cc_727 N_A_1383_349#_M1033_g N_VPWR_c_1780_n 0.00376235f $X=7.005 $Y=2.495 $X2=0
+ $Y2=0
cc_728 N_A_1383_349#_c_834_n N_VPWR_c_1781_n 0.0171249f $X=8.95 $Y=2.235 $X2=0
+ $Y2=0
cc_729 N_A_1383_349#_c_834_n N_VPWR_c_1795_n 0.00804742f $X=8.95 $Y=2.235 $X2=0
+ $Y2=0
cc_730 N_A_1383_349#_M1033_g N_VPWR_c_1777_n 0.00113998f $X=7.005 $Y=2.495 $X2=0
+ $Y2=0
cc_731 N_A_1383_349#_c_834_n N_VPWR_c_1777_n 0.0100639f $X=8.95 $Y=2.235 $X2=0
+ $Y2=0
cc_732 N_A_1383_349#_c_827_n N_VGND_M1007_d 0.0208142f $X=8.59 $Y=1.005 $X2=0
+ $Y2=0
cc_733 N_A_1383_349#_c_827_n A_1432_119# 2.87715e-19 $X=8.59 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_734 N_A_1383_349#_c_848_n A_1432_119# 0.001002f $X=7.315 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_735 N_RESET_B_c_935_n N_A_1235_119#_M1006_g 0.0161199f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_736 N_RESET_B_c_936_n N_A_1235_119#_M1006_g 0.00187394f $X=8.545 $Y=2.035
+ $X2=0 $Y2=0
cc_737 N_RESET_B_c_937_n N_A_1235_119#_M1006_g 0.00290543f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_738 N_RESET_B_c_940_n N_A_1235_119#_M1006_g 0.0086835f $X=7.975 $Y=1.96 $X2=0
+ $Y2=0
cc_739 N_RESET_B_c_925_n N_A_1235_119#_c_1138_n 0.0105479f $X=7.645 $Y=1.26
+ $X2=0 $Y2=0
cc_740 N_RESET_B_c_937_n N_A_1235_119#_c_1138_n 0.00978949f $X=8.4 $Y=2.035
+ $X2=0 $Y2=0
cc_741 N_RESET_B_c_940_n N_A_1235_119#_c_1138_n 0.00287914f $X=7.975 $Y=1.96
+ $X2=0 $Y2=0
cc_742 N_RESET_B_c_936_n N_A_1235_119#_c_1139_n 7.899e-19 $X=8.545 $Y=2.035
+ $X2=0 $Y2=0
cc_743 N_RESET_B_c_933_n N_A_1235_119#_c_1148_n 0.00719547f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_744 N_RESET_B_c_933_n N_A_1235_119#_c_1140_n 0.0221124f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_745 N_RESET_B_c_933_n N_A_1235_119#_c_1177_n 0.0204635f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_746 N_RESET_B_M1013_g N_A_1235_119#_c_1141_n 0.0239921f $X=7.63 $Y=2.495
+ $X2=0 $Y2=0
cc_747 N_RESET_B_c_922_n N_A_1235_119#_c_1141_n 0.0114947f $X=7.645 $Y=1.795
+ $X2=0 $Y2=0
cc_748 N_RESET_B_c_933_n N_A_1235_119#_c_1141_n 0.0293251f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_749 N_RESET_B_c_936_n N_A_1235_119#_c_1141_n 2.61031e-19 $X=8.545 $Y=2.035
+ $X2=0 $Y2=0
cc_750 N_RESET_B_c_937_n N_A_1235_119#_c_1141_n 0.0403674f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_751 N_RESET_B_c_940_n N_A_1235_119#_c_1141_n 0.0133467f $X=7.975 $Y=1.96
+ $X2=0 $Y2=0
cc_752 N_RESET_B_c_922_n N_A_1235_119#_c_1142_n 0.00390473f $X=7.645 $Y=1.795
+ $X2=0 $Y2=0
cc_753 N_RESET_B_c_925_n N_A_1235_119#_c_1142_n 0.00529036f $X=7.645 $Y=1.26
+ $X2=0 $Y2=0
cc_754 N_RESET_B_c_922_n N_A_1235_119#_c_1143_n 0.00624417f $X=7.645 $Y=1.795
+ $X2=0 $Y2=0
cc_755 N_RESET_B_c_925_n N_A_1235_119#_c_1143_n 0.00198801f $X=7.645 $Y=1.26
+ $X2=0 $Y2=0
cc_756 N_RESET_B_c_933_n N_A_1235_119#_c_1143_n 0.0080909f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_757 N_RESET_B_c_936_n N_A_1235_119#_c_1143_n 8.96068e-19 $X=8.545 $Y=2.035
+ $X2=0 $Y2=0
cc_758 N_RESET_B_c_937_n N_A_1235_119#_c_1143_n 0.0351039f $X=8.4 $Y=2.035 $X2=0
+ $Y2=0
cc_759 N_RESET_B_c_940_n N_A_1235_119#_c_1143_n 0.0100276f $X=7.975 $Y=1.96
+ $X2=0 $Y2=0
cc_760 N_RESET_B_c_933_n N_A_837_119#_M1027_s 0.00116422f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_761 N_RESET_B_c_933_n N_A_837_119#_c_1272_n 2.92073e-19 $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_762 N_RESET_B_c_919_n N_A_837_119#_c_1260_n 0.00881316f $X=7.4 $Y=0.18 $X2=0
+ $Y2=0
cc_763 N_RESET_B_c_933_n N_A_837_119#_M1025_g 0.00283681f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_764 N_RESET_B_M1013_g N_A_837_119#_c_1277_n 0.0102838f $X=7.63 $Y=2.495 $X2=0
+ $Y2=0
cc_765 N_RESET_B_c_935_n N_A_837_119#_M1020_g 0.0102815f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_766 N_RESET_B_c_935_n N_A_837_119#_c_1261_n 0.00577012f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_767 N_RESET_B_c_933_n N_A_837_119#_c_1265_n 0.00275836f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_768 N_RESET_B_c_919_n N_A_837_119#_c_1288_n 0.00281183f $X=7.4 $Y=0.18 $X2=0
+ $Y2=0
cc_769 N_RESET_B_c_933_n N_A_837_119#_c_1291_n 0.0225779f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_770 N_RESET_B_c_934_n N_A_837_119#_c_1283_n 5.46046e-19 $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_771 N_RESET_B_c_939_n N_A_837_119#_c_1283_n 0.00314885f $X=3.95 $Y=1.995
+ $X2=0 $Y2=0
cc_772 N_RESET_B_M1004_g N_A_837_119#_c_1268_n 0.00193025f $X=3.515 $Y=0.615
+ $X2=0 $Y2=0
cc_773 N_RESET_B_c_919_n N_A_837_119#_c_1268_n 0.00603673f $X=7.4 $Y=0.18 $X2=0
+ $Y2=0
cc_774 N_RESET_B_c_933_n N_A_837_119#_c_1300_n 0.0114432f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_775 N_RESET_B_c_934_n N_A_837_119#_c_1300_n 0.00200463f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_776 N_RESET_B_c_938_n N_A_837_119#_c_1300_n 6.26563e-19 $X=3.95 $Y=1.995
+ $X2=0 $Y2=0
cc_777 N_RESET_B_c_939_n N_A_837_119#_c_1300_n 0.0150716f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_778 N_RESET_B_c_933_n N_A_837_119#_c_1269_n 0.00588539f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_779 N_RESET_B_c_933_n N_A_837_119#_c_1270_n 5.3491e-19 $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_780 N_RESET_B_c_919_n N_A_837_119#_c_1271_n 0.010225f $X=7.4 $Y=0.18 $X2=0
+ $Y2=0
cc_781 N_RESET_B_c_933_n N_A_837_119#_c_1286_n 0.00385098f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_782 N_RESET_B_M1019_g N_A_2082_446#_M1005_g 0.00463034f $X=11.35 $Y=2.75
+ $X2=0 $Y2=0
cc_783 N_RESET_B_M1026_g N_A_2082_446#_M1010_g 0.0332604f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_784 N_RESET_B_M1019_g N_A_2082_446#_c_1469_n 0.00483575f $X=11.35 $Y=2.75
+ $X2=0 $Y2=0
cc_785 N_RESET_B_c_935_n N_A_2082_446#_c_1469_n 8.58242e-19 $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_786 N_RESET_B_M1019_g N_A_2082_446#_c_1481_n 0.00102797f $X=11.35 $Y=2.75
+ $X2=0 $Y2=0
cc_787 N_RESET_B_c_935_n N_A_2082_446#_c_1481_n 0.0371304f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_788 RESET_B N_A_2082_446#_c_1481_n 5.86564e-19 $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_789 N_RESET_B_c_941_n N_A_2082_446#_c_1481_n 0.00153537f $X=11.275 $Y=2.07
+ $X2=0 $Y2=0
cc_790 N_RESET_B_c_1052_p N_A_2082_446#_c_1481_n 0.0134652f $X=11.28 $Y=2.035
+ $X2=0 $Y2=0
cc_791 N_RESET_B_c_935_n N_A_2082_446#_c_1460_n 0.0118555f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_792 N_RESET_B_c_941_n N_A_2082_446#_c_1460_n 0.031607f $X=11.275 $Y=2.07
+ $X2=0 $Y2=0
cc_793 N_RESET_B_c_1052_p N_A_2082_446#_c_1460_n 0.00107974f $X=11.28 $Y=2.035
+ $X2=0 $Y2=0
cc_794 N_RESET_B_M1026_g N_A_2082_446#_c_1461_n 0.0112646f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_795 N_RESET_B_c_935_n N_A_2082_446#_c_1461_n 0.00766736f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_796 RESET_B N_A_2082_446#_c_1461_n 0.0021857f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_797 N_RESET_B_c_941_n N_A_2082_446#_c_1461_n 0.00568091f $X=11.275 $Y=2.07
+ $X2=0 $Y2=0
cc_798 N_RESET_B_c_1052_p N_A_2082_446#_c_1461_n 0.0208148f $X=11.28 $Y=2.035
+ $X2=0 $Y2=0
cc_799 N_RESET_B_M1019_g N_A_2082_446#_c_1472_n 0.0137018f $X=11.35 $Y=2.75
+ $X2=0 $Y2=0
cc_800 N_RESET_B_c_935_n N_A_2082_446#_c_1472_n 0.00726729f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_801 RESET_B N_A_2082_446#_c_1472_n 0.00176886f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_802 N_RESET_B_c_941_n N_A_2082_446#_c_1472_n 0.00469264f $X=11.275 $Y=2.07
+ $X2=0 $Y2=0
cc_803 N_RESET_B_c_1052_p N_A_2082_446#_c_1472_n 0.0223172f $X=11.28 $Y=2.035
+ $X2=0 $Y2=0
cc_804 N_RESET_B_M1019_g N_A_2082_446#_c_1473_n 0.0110799f $X=11.35 $Y=2.75
+ $X2=0 $Y2=0
cc_805 N_RESET_B_M1026_g N_A_2082_446#_c_1462_n 0.00114233f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_806 N_RESET_B_M1026_g N_A_2082_446#_c_1464_n 7.54334e-19 $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_807 N_RESET_B_M1026_g N_A_2082_446#_c_1466_n 0.00211977f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_808 N_RESET_B_M1026_g N_A_2082_446#_c_1467_n 0.0225188f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_809 N_RESET_B_c_935_n N_A_1824_74#_M1020_d 6.85563e-19 $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_810 N_RESET_B_M1026_g N_A_1824_74#_M1018_g 0.0603983f $X=11.135 $Y=0.58 $X2=0
+ $Y2=0
cc_811 N_RESET_B_M1026_g N_A_1824_74#_c_1592_n 0.00632307f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_812 N_RESET_B_c_941_n N_A_1824_74#_M1024_g 0.0375449f $X=11.275 $Y=2.07 $X2=0
+ $Y2=0
cc_813 N_RESET_B_c_1052_p N_A_1824_74#_M1024_g 0.00121903f $X=11.28 $Y=2.035
+ $X2=0 $Y2=0
cc_814 N_RESET_B_M1026_g N_A_1824_74#_c_1580_n 0.00629822f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_815 N_RESET_B_c_941_n N_A_1824_74#_c_1580_n 2.30537e-19 $X=11.275 $Y=2.07
+ $X2=0 $Y2=0
cc_816 N_RESET_B_M1026_g N_A_1824_74#_c_1583_n 0.00585373f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_817 N_RESET_B_c_935_n N_A_1824_74#_c_1601_n 0.028385f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_818 N_RESET_B_c_935_n N_A_1824_74#_c_1595_n 0.0138331f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_819 N_RESET_B_c_935_n N_A_1824_74#_c_1587_n 0.023417f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_820 N_RESET_B_M1026_g N_A_1824_74#_c_1588_n 0.00517953f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_821 N_RESET_B_M1026_g N_A_1824_74#_c_1591_n 0.0159185f $X=11.135 $Y=0.58
+ $X2=0 $Y2=0
cc_822 N_RESET_B_c_933_n N_VPWR_M1027_d 3.376e-19 $X=8.255 $Y=2.035 $X2=0 $Y2=0
cc_823 N_RESET_B_c_936_n N_VPWR_M1006_s 0.00313047f $X=8.545 $Y=2.035 $X2=0
+ $Y2=0
cc_824 N_RESET_B_c_937_n N_VPWR_M1006_s 0.00634743f $X=8.4 $Y=2.035 $X2=0 $Y2=0
cc_825 N_RESET_B_M1023_g N_VPWR_c_1778_n 0.00944745f $X=3.505 $Y=2.735 $X2=0
+ $Y2=0
cc_826 N_RESET_B_M1013_g N_VPWR_c_1780_n 0.00373896f $X=7.63 $Y=2.495 $X2=0
+ $Y2=0
cc_827 N_RESET_B_M1013_g N_VPWR_c_1781_n 0.00361589f $X=7.63 $Y=2.495 $X2=0
+ $Y2=0
cc_828 N_RESET_B_c_935_n N_VPWR_c_1781_n 0.00146686f $X=11.135 $Y=2.035 $X2=0
+ $Y2=0
cc_829 N_RESET_B_c_936_n N_VPWR_c_1781_n 0.00903602f $X=8.545 $Y=2.035 $X2=0
+ $Y2=0
cc_830 N_RESET_B_c_937_n N_VPWR_c_1781_n 0.017909f $X=8.4 $Y=2.035 $X2=0 $Y2=0
cc_831 RESET_B N_VPWR_c_1782_n 0.00143958f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_832 N_RESET_B_c_1052_p N_VPWR_c_1782_n 0.00812957f $X=11.28 $Y=2.035 $X2=0
+ $Y2=0
cc_833 N_RESET_B_M1023_g N_VPWR_c_1786_n 0.00616631f $X=3.505 $Y=2.735 $X2=0
+ $Y2=0
cc_834 N_RESET_B_M1019_g N_VPWR_c_1790_n 0.005209f $X=11.35 $Y=2.75 $X2=0 $Y2=0
cc_835 N_RESET_B_M1019_g N_VPWR_c_1801_n 0.0043693f $X=11.35 $Y=2.75 $X2=0 $Y2=0
cc_836 N_RESET_B_M1023_g N_VPWR_c_1777_n 0.00680759f $X=3.505 $Y=2.735 $X2=0
+ $Y2=0
cc_837 N_RESET_B_M1013_g N_VPWR_c_1777_n 0.00113998f $X=7.63 $Y=2.495 $X2=0
+ $Y2=0
cc_838 N_RESET_B_M1019_g N_VPWR_c_1777_n 0.00517685f $X=11.35 $Y=2.75 $X2=0
+ $Y2=0
cc_839 N_RESET_B_M1004_g N_A_390_81#_c_1947_n 3.15251e-19 $X=3.515 $Y=0.615
+ $X2=0 $Y2=0
cc_840 N_RESET_B_M1023_g N_A_390_81#_c_1957_n 0.00434499f $X=3.505 $Y=2.735
+ $X2=0 $Y2=0
cc_841 N_RESET_B_M1004_g N_A_390_81#_c_1948_n 2.84226e-19 $X=3.515 $Y=0.615
+ $X2=0 $Y2=0
cc_842 N_RESET_B_c_924_n N_A_390_81#_c_1948_n 0.00129005f $X=3.502 $Y=1.075
+ $X2=0 $Y2=0
cc_843 N_RESET_B_c_917_n N_A_390_81#_c_1949_n 0.015085f $X=3.49 $Y=1.83 $X2=0
+ $Y2=0
cc_844 N_RESET_B_c_924_n N_A_390_81#_c_1949_n 0.00135631f $X=3.502 $Y=1.075
+ $X2=0 $Y2=0
cc_845 N_RESET_B_c_917_n N_A_390_81#_c_1951_n 0.0139879f $X=3.49 $Y=1.83 $X2=0
+ $Y2=0
cc_846 N_RESET_B_M1023_g N_A_390_81#_c_1951_n 0.00699164f $X=3.505 $Y=2.735
+ $X2=0 $Y2=0
cc_847 N_RESET_B_c_932_n N_A_390_81#_c_1951_n 0.00713227f $X=3.505 $Y=1.995
+ $X2=0 $Y2=0
cc_848 N_RESET_B_c_934_n N_A_390_81#_c_1951_n 0.00108729f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_849 N_RESET_B_c_938_n N_A_390_81#_c_1951_n 0.0057826f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_850 N_RESET_B_c_939_n N_A_390_81#_c_1951_n 0.0228135f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_851 N_RESET_B_c_933_n N_A_390_81#_c_1960_n 0.0177348f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_852 N_RESET_B_c_934_n N_A_390_81#_c_1960_n 0.00373288f $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_853 N_RESET_B_c_938_n N_A_390_81#_c_1960_n 0.00248575f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_854 N_RESET_B_c_939_n N_A_390_81#_c_1960_n 0.00754045f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_855 N_RESET_B_c_933_n N_A_390_81#_c_1962_n 0.0115758f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_856 N_RESET_B_c_933_n N_A_390_81#_c_1963_n 0.00767724f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_857 N_RESET_B_c_933_n N_A_390_81#_c_1953_n 0.00410787f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_858 N_RESET_B_c_933_n N_A_390_81#_c_1955_n 0.0156292f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_859 N_RESET_B_M1023_g N_A_390_81#_c_1965_n 0.0203875f $X=3.505 $Y=2.735 $X2=0
+ $Y2=0
cc_860 N_RESET_B_c_934_n N_A_390_81#_c_1965_n 5.00635e-19 $X=4.225 $Y=2.035
+ $X2=0 $Y2=0
cc_861 N_RESET_B_c_938_n N_A_390_81#_c_1965_n 0.0124471f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_862 N_RESET_B_c_939_n N_A_390_81#_c_1965_n 0.017195f $X=3.95 $Y=1.995 $X2=0
+ $Y2=0
cc_863 N_RESET_B_M1004_g N_VGND_c_2138_n 0.0120745f $X=3.515 $Y=0.615 $X2=0
+ $Y2=0
cc_864 N_RESET_B_c_919_n N_VGND_c_2138_n 0.0232366f $X=7.4 $Y=0.18 $X2=0 $Y2=0
cc_865 N_RESET_B_c_919_n N_VGND_c_2139_n 0.0217794f $X=7.4 $Y=0.18 $X2=0 $Y2=0
cc_866 N_RESET_B_M1026_g N_VGND_c_2140_n 0.0122528f $X=11.135 $Y=0.58 $X2=0
+ $Y2=0
cc_867 N_RESET_B_c_920_n N_VGND_c_2145_n 0.00874174f $X=3.59 $Y=0.18 $X2=0 $Y2=0
cc_868 N_RESET_B_c_919_n N_VGND_c_2147_n 0.0226045f $X=7.4 $Y=0.18 $X2=0 $Y2=0
cc_869 N_RESET_B_c_919_n N_VGND_c_2150_n 0.0663838f $X=7.4 $Y=0.18 $X2=0 $Y2=0
cc_870 N_RESET_B_M1026_g N_VGND_c_2152_n 0.00383152f $X=11.135 $Y=0.58 $X2=0
+ $Y2=0
cc_871 N_RESET_B_c_919_n N_VGND_c_2159_n 0.0981736f $X=7.4 $Y=0.18 $X2=0 $Y2=0
cc_872 N_RESET_B_c_920_n N_VGND_c_2159_n 0.0115384f $X=3.59 $Y=0.18 $X2=0 $Y2=0
cc_873 N_RESET_B_M1026_g N_VGND_c_2159_n 0.0075694f $X=11.135 $Y=0.58 $X2=0
+ $Y2=0
cc_874 N_RESET_B_M1004_g N_noxref_24_c_2273_n 0.00196666f $X=3.515 $Y=0.615
+ $X2=0 $Y2=0
cc_875 N_A_1235_119#_c_1140_n N_A_837_119#_c_1258_n 5.0125e-19 $X=6.785 $Y=2.32
+ $X2=0 $Y2=0
cc_876 N_A_1235_119#_c_1148_n N_A_837_119#_c_1274_n 0.00380204f $X=6.7 $Y=2.6
+ $X2=0 $Y2=0
cc_877 N_A_1235_119#_c_1144_n N_A_837_119#_c_1260_n 0.00427553f $X=6.48 $Y=0.81
+ $X2=0 $Y2=0
cc_878 N_A_1235_119#_c_1148_n N_A_837_119#_M1025_g 0.0120094f $X=6.7 $Y=2.6
+ $X2=0 $Y2=0
cc_879 N_A_1235_119#_c_1140_n N_A_837_119#_M1025_g 0.00104602f $X=6.785 $Y=2.32
+ $X2=0 $Y2=0
cc_880 N_A_1235_119#_M1006_g N_A_837_119#_c_1277_n 0.0123711f $X=8.64 $Y=2.235
+ $X2=0 $Y2=0
cc_881 N_A_1235_119#_c_1177_n N_A_837_119#_c_1277_n 0.00162087f $X=7.485
+ $Y=2.405 $X2=0 $Y2=0
cc_882 N_A_1235_119#_c_1141_n N_A_837_119#_c_1277_n 0.00632743f $X=7.57 $Y=2.32
+ $X2=0 $Y2=0
cc_883 N_A_1235_119#_c_1151_n N_A_837_119#_c_1277_n 0.00168131f $X=6.785
+ $Y=2.522 $X2=0 $Y2=0
cc_884 N_A_1235_119#_M1006_g N_A_837_119#_c_1280_n 0.0262478f $X=8.64 $Y=2.235
+ $X2=0 $Y2=0
cc_885 N_A_1235_119#_M1006_g N_A_1824_74#_c_1596_n 4.67625e-19 $X=8.64 $Y=2.235
+ $X2=0 $Y2=0
cc_886 N_A_1235_119#_c_1177_n N_VPWR_M1033_d 0.00755907f $X=7.485 $Y=2.405 $X2=0
+ $Y2=0
cc_887 N_A_1235_119#_c_1177_n N_VPWR_c_1780_n 0.0254917f $X=7.485 $Y=2.405 $X2=0
+ $Y2=0
cc_888 N_A_1235_119#_c_1141_n N_VPWR_c_1780_n 0.00280675f $X=7.57 $Y=2.32 $X2=0
+ $Y2=0
cc_889 N_A_1235_119#_c_1151_n N_VPWR_c_1780_n 0.00118439f $X=6.785 $Y=2.522
+ $X2=0 $Y2=0
cc_890 N_A_1235_119#_M1006_g N_VPWR_c_1781_n 0.0113098f $X=8.64 $Y=2.235 $X2=0
+ $Y2=0
cc_891 N_A_1235_119#_c_1141_n N_VPWR_c_1781_n 0.02806f $X=7.57 $Y=2.32 $X2=0
+ $Y2=0
cc_892 N_A_1235_119#_c_1148_n N_VPWR_c_1788_n 0.00965271f $X=6.7 $Y=2.6 $X2=0
+ $Y2=0
cc_893 N_A_1235_119#_c_1151_n N_VPWR_c_1788_n 0.00364353f $X=6.785 $Y=2.522
+ $X2=0 $Y2=0
cc_894 N_A_1235_119#_c_1141_n N_VPWR_c_1794_n 0.00677432f $X=7.57 $Y=2.32 $X2=0
+ $Y2=0
cc_895 N_A_1235_119#_M1006_g N_VPWR_c_1777_n 9.455e-19 $X=8.64 $Y=2.235 $X2=0
+ $Y2=0
cc_896 N_A_1235_119#_c_1148_n N_VPWR_c_1777_n 0.0127233f $X=6.7 $Y=2.6 $X2=0
+ $Y2=0
cc_897 N_A_1235_119#_c_1177_n N_VPWR_c_1777_n 0.00908852f $X=7.485 $Y=2.405
+ $X2=0 $Y2=0
cc_898 N_A_1235_119#_c_1141_n N_VPWR_c_1777_n 0.015216f $X=7.57 $Y=2.32 $X2=0
+ $Y2=0
cc_899 N_A_1235_119#_c_1151_n N_VPWR_c_1777_n 0.00458771f $X=6.785 $Y=2.522
+ $X2=0 $Y2=0
cc_900 N_A_1235_119#_c_1148_n N_A_390_81#_c_1961_n 0.0098387f $X=6.7 $Y=2.6
+ $X2=0 $Y2=0
cc_901 N_A_1235_119#_c_1140_n N_A_390_81#_c_1952_n 0.00456668f $X=6.785 $Y=2.32
+ $X2=0 $Y2=0
cc_902 N_A_1235_119#_c_1144_n N_A_390_81#_c_1952_n 0.0332844f $X=6.48 $Y=0.81
+ $X2=0 $Y2=0
cc_903 N_A_1235_119#_M1002_d N_A_390_81#_c_1962_n 0.00190768f $X=6.225 $Y=2.285
+ $X2=0 $Y2=0
cc_904 N_A_1235_119#_c_1148_n N_A_390_81#_c_1962_n 0.0162637f $X=6.7 $Y=2.6
+ $X2=0 $Y2=0
cc_905 N_A_1235_119#_c_1140_n N_A_390_81#_c_1962_n 0.0128814f $X=6.785 $Y=2.32
+ $X2=0 $Y2=0
cc_906 N_A_1235_119#_c_1140_n N_A_390_81#_c_1953_n 0.0131857f $X=6.785 $Y=2.32
+ $X2=0 $Y2=0
cc_907 N_A_1235_119#_c_1144_n N_A_390_81#_c_1953_n 0.0191771f $X=6.48 $Y=0.81
+ $X2=0 $Y2=0
cc_908 N_A_1235_119#_c_1140_n N_A_390_81#_c_1955_n 0.048352f $X=6.785 $Y=2.32
+ $X2=0 $Y2=0
cc_909 N_A_1235_119#_M1040_g N_VGND_c_2150_n 0.00115066f $X=8.54 $Y=0.74 $X2=0
+ $Y2=0
cc_910 N_A_1235_119#_M1040_g N_VGND_c_2151_n 0.00278271f $X=8.54 $Y=0.74 $X2=0
+ $Y2=0
cc_911 N_A_1235_119#_M1040_g N_VGND_c_2159_n 0.0035918f $X=8.54 $Y=0.74 $X2=0
+ $Y2=0
cc_912 N_A_1235_119#_c_1144_n A_1354_119# 0.00123907f $X=6.48 $Y=0.81 $X2=-0.19
+ $Y2=-0.245
cc_913 N_A_837_119#_c_1262_n N_A_2082_446#_M1010_g 0.00472321f $X=10.125
+ $Y=1.575 $X2=0 $Y2=0
cc_914 N_A_837_119#_M1009_g N_A_2082_446#_M1010_g 0.0465564f $X=10.315 $Y=0.58
+ $X2=0 $Y2=0
cc_915 N_A_837_119#_c_1261_n N_A_2082_446#_c_1460_n 0.00873113f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_916 N_A_837_119#_c_1262_n N_A_2082_446#_c_1467_n 0.00873113f $X=10.125
+ $Y=1.575 $X2=0 $Y2=0
cc_917 N_A_837_119#_M1020_g N_A_1824_74#_c_1601_n 0.00834084f $X=9.26 $Y=2.33
+ $X2=0 $Y2=0
cc_918 N_A_837_119#_c_1261_n N_A_1824_74#_c_1601_n 0.00614737f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_919 N_A_837_119#_M1009_g N_A_1824_74#_c_1585_n 0.0085841f $X=10.315 $Y=0.58
+ $X2=0 $Y2=0
cc_920 N_A_837_119#_c_1266_n N_A_1824_74#_c_1585_n 0.0073765f $X=10.315 $Y=1.055
+ $X2=0 $Y2=0
cc_921 N_A_837_119#_M1020_g N_A_1824_74#_c_1596_n 0.0060423f $X=9.26 $Y=2.33
+ $X2=0 $Y2=0
cc_922 N_A_837_119#_M1009_g N_A_1824_74#_c_1586_n 0.00682018f $X=10.315 $Y=0.58
+ $X2=0 $Y2=0
cc_923 N_A_837_119#_c_1266_n N_A_1824_74#_c_1586_n 0.00308052f $X=10.315
+ $Y=1.055 $X2=0 $Y2=0
cc_924 N_A_837_119#_c_1262_n N_A_1824_74#_c_1587_n 0.00432791f $X=10.125
+ $Y=1.575 $X2=0 $Y2=0
cc_925 N_A_837_119#_c_1262_n N_A_1824_74#_c_1589_n 7.4004e-19 $X=10.125 $Y=1.575
+ $X2=0 $Y2=0
cc_926 N_A_837_119#_c_1266_n N_A_1824_74#_c_1589_n 0.00823777f $X=10.315
+ $Y=1.055 $X2=0 $Y2=0
cc_927 N_A_837_119#_c_1291_n N_VPWR_M1027_d 0.00325331f $X=4.815 $Y=2.03 $X2=0
+ $Y2=0
cc_928 N_A_837_119#_c_1273_n N_VPWR_c_1779_n 0.00203598f $X=5.61 $Y=3.075 $X2=0
+ $Y2=0
cc_929 N_A_837_119#_c_1275_n N_VPWR_c_1779_n 7.02368e-19 $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_930 N_A_837_119#_c_1286_n N_VPWR_c_1779_n 0.0105232f $X=5.13 $Y=1.86 $X2=0
+ $Y2=0
cc_931 N_A_837_119#_M1025_g N_VPWR_c_1780_n 0.00690475f $X=6.605 $Y=2.495 $X2=0
+ $Y2=0
cc_932 N_A_837_119#_c_1277_n N_VPWR_c_1780_n 0.025635f $X=9.17 $Y=3.15 $X2=0
+ $Y2=0
cc_933 N_A_837_119#_c_1277_n N_VPWR_c_1781_n 0.0257203f $X=9.17 $Y=3.15 $X2=0
+ $Y2=0
cc_934 N_A_837_119#_M1020_g N_VPWR_c_1781_n 0.00568708f $X=9.26 $Y=2.33 $X2=0
+ $Y2=0
cc_935 N_A_837_119#_c_1275_n N_VPWR_c_1788_n 0.047056f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_936 N_A_837_119#_c_1286_n N_VPWR_c_1788_n 0.00401239f $X=5.13 $Y=1.86 $X2=0
+ $Y2=0
cc_937 N_A_837_119#_c_1277_n N_VPWR_c_1794_n 0.0233394f $X=9.17 $Y=3.15 $X2=0
+ $Y2=0
cc_938 N_A_837_119#_c_1277_n N_VPWR_c_1795_n 0.0236738f $X=9.17 $Y=3.15 $X2=0
+ $Y2=0
cc_939 N_A_837_119#_c_1274_n N_VPWR_c_1777_n 0.0244696f $X=6.515 $Y=3.15 $X2=0
+ $Y2=0
cc_940 N_A_837_119#_c_1275_n N_VPWR_c_1777_n 0.00618409f $X=5.69 $Y=3.15 $X2=0
+ $Y2=0
cc_941 N_A_837_119#_c_1277_n N_VPWR_c_1777_n 0.0705251f $X=9.17 $Y=3.15 $X2=0
+ $Y2=0
cc_942 N_A_837_119#_c_1282_n N_VPWR_c_1777_n 0.00508747f $X=6.605 $Y=3.15 $X2=0
+ $Y2=0
cc_943 N_A_837_119#_c_1286_n N_VPWR_c_1777_n 0.00500915f $X=5.13 $Y=1.86 $X2=0
+ $Y2=0
cc_944 N_A_837_119#_M1027_s N_A_390_81#_c_1960_n 0.00770925f $X=4.275 $Y=1.935
+ $X2=0 $Y2=0
cc_945 N_A_837_119#_c_1273_n N_A_390_81#_c_1960_n 0.0145389f $X=5.61 $Y=3.075
+ $X2=0 $Y2=0
cc_946 N_A_837_119#_c_1291_n N_A_390_81#_c_1960_n 0.0110961f $X=4.815 $Y=2.03
+ $X2=0 $Y2=0
cc_947 N_A_837_119#_c_1300_n N_A_390_81#_c_1960_n 0.0137082f $X=4.46 $Y=2.03
+ $X2=0 $Y2=0
cc_948 N_A_837_119#_c_1269_n N_A_390_81#_c_1960_n 0.00140597f $X=5.13 $Y=1.61
+ $X2=0 $Y2=0
cc_949 N_A_837_119#_c_1286_n N_A_390_81#_c_1960_n 0.0160652f $X=5.13 $Y=1.86
+ $X2=0 $Y2=0
cc_950 N_A_837_119#_c_1273_n N_A_390_81#_c_1961_n 0.00637944f $X=5.61 $Y=3.075
+ $X2=0 $Y2=0
cc_951 N_A_837_119#_c_1274_n N_A_390_81#_c_1961_n 0.00421145f $X=6.515 $Y=3.15
+ $X2=0 $Y2=0
cc_952 N_A_837_119#_c_1257_n N_A_390_81#_c_1952_n 0.00112915f $X=5.605 $Y=1.41
+ $X2=0 $Y2=0
cc_953 N_A_837_119#_c_1258_n N_A_390_81#_c_1952_n 0.0179613f $X=6.025 $Y=1.165
+ $X2=0 $Y2=0
cc_954 N_A_837_119#_c_1260_n N_A_390_81#_c_1952_n 0.0090845f $X=6.1 $Y=1.09
+ $X2=0 $Y2=0
cc_955 N_A_837_119#_M1025_g N_A_390_81#_c_1962_n 0.00377426f $X=6.605 $Y=2.495
+ $X2=0 $Y2=0
cc_956 N_A_837_119#_c_1272_n N_A_390_81#_c_1963_n 0.00170292f $X=5.61 $Y=2.275
+ $X2=0 $Y2=0
cc_957 N_A_837_119#_c_1265_n N_A_390_81#_c_1963_n 5.32154e-19 $X=5.61 $Y=2.195
+ $X2=0 $Y2=0
cc_958 N_A_837_119#_c_1258_n N_A_390_81#_c_1953_n 0.00158731f $X=6.025 $Y=1.165
+ $X2=0 $Y2=0
cc_959 N_A_837_119#_c_1257_n N_A_390_81#_c_1954_n 0.00406108f $X=5.605 $Y=1.41
+ $X2=0 $Y2=0
cc_960 N_A_837_119#_c_1264_n N_A_390_81#_c_1955_n 0.00271528f $X=5.605 $Y=1.485
+ $X2=0 $Y2=0
cc_961 N_A_837_119#_c_1265_n N_A_390_81#_c_1955_n 2.11377e-19 $X=5.61 $Y=2.195
+ $X2=0 $Y2=0
cc_962 N_A_837_119#_c_1288_n N_VGND_M1016_d 0.00911076f $X=4.815 $Y=1.005 $X2=0
+ $Y2=0
cc_963 N_A_837_119#_c_1267_n N_VGND_M1016_d 0.0042694f $X=4.9 $Y=1.445 $X2=0
+ $Y2=0
cc_964 N_A_837_119#_c_1268_n N_VGND_c_2138_n 0.0150432f $X=4.31 $Y=0.76 $X2=0
+ $Y2=0
cc_965 N_A_837_119#_c_1288_n N_VGND_c_2139_n 0.0204055f $X=4.815 $Y=1.005 $X2=0
+ $Y2=0
cc_966 N_A_837_119#_c_1268_n N_VGND_c_2139_n 0.0121035f $X=4.31 $Y=0.76 $X2=0
+ $Y2=0
cc_967 N_A_837_119#_c_1271_n N_VGND_c_2139_n 0.00217883f $X=5.13 $Y=1.41 $X2=0
+ $Y2=0
cc_968 N_A_837_119#_M1009_g N_VGND_c_2140_n 0.00155929f $X=10.315 $Y=0.58 $X2=0
+ $Y2=0
cc_969 N_A_837_119#_c_1268_n N_VGND_c_2147_n 0.00785495f $X=4.31 $Y=0.76 $X2=0
+ $Y2=0
cc_970 N_A_837_119#_M1009_g N_VGND_c_2151_n 0.00308264f $X=10.315 $Y=0.58 $X2=0
+ $Y2=0
cc_971 N_A_837_119#_M1009_g N_VGND_c_2159_n 0.00383744f $X=10.315 $Y=0.58 $X2=0
+ $Y2=0
cc_972 N_A_837_119#_c_1268_n N_VGND_c_2159_n 0.0110687f $X=4.31 $Y=0.76 $X2=0
+ $Y2=0
cc_973 N_A_837_119#_c_1271_n N_VGND_c_2159_n 8.45315e-19 $X=5.13 $Y=1.41 $X2=0
+ $Y2=0
cc_974 N_A_2082_446#_c_1462_n N_A_1824_74#_M1018_g 0.00761651f $X=11.71 $Y=0.58
+ $X2=0 $Y2=0
cc_975 N_A_2082_446#_c_1464_n N_A_1824_74#_M1018_g 0.00732912f $X=11.875
+ $Y=0.855 $X2=0 $Y2=0
cc_976 N_A_2082_446#_c_1465_n N_A_1824_74#_M1018_g 0.00376832f $X=12.145 $Y=1.58
+ $X2=0 $Y2=0
cc_977 N_A_2082_446#_c_1461_n N_A_1824_74#_c_1592_n 0.0116511f $X=12.06 $Y=1.665
+ $X2=0 $Y2=0
cc_978 N_A_2082_446#_c_1472_n N_A_1824_74#_M1024_g 0.00477715f $X=11.41 $Y=2.475
+ $X2=0 $Y2=0
cc_979 N_A_2082_446#_c_1473_n N_A_1824_74#_M1024_g 0.00581157f $X=11.575 $Y=2.75
+ $X2=0 $Y2=0
cc_980 N_A_2082_446#_c_1461_n N_A_1824_74#_c_1579_n 0.00220284f $X=12.06
+ $Y=1.665 $X2=0 $Y2=0
cc_981 N_A_2082_446#_c_1465_n N_A_1824_74#_c_1579_n 0.022644f $X=12.145 $Y=1.58
+ $X2=0 $Y2=0
cc_982 N_A_2082_446#_c_1461_n N_A_1824_74#_c_1580_n 0.00461365f $X=12.06
+ $Y=1.665 $X2=0 $Y2=0
cc_983 N_A_2082_446#_c_1463_n N_A_1824_74#_c_1580_n 0.0054249f $X=12.06 $Y=0.855
+ $X2=0 $Y2=0
cc_984 N_A_2082_446#_c_1464_n N_A_1824_74#_c_1580_n 0.00561111f $X=11.875
+ $Y=0.855 $X2=0 $Y2=0
cc_985 N_A_2082_446#_c_1461_n N_A_1824_74#_M1037_g 0.00230014f $X=12.06 $Y=1.665
+ $X2=0 $Y2=0
cc_986 N_A_2082_446#_c_1465_n N_A_1824_74#_M1037_g 0.0017493f $X=12.145 $Y=1.58
+ $X2=0 $Y2=0
cc_987 N_A_2082_446#_c_1462_n N_A_1824_74#_c_1582_n 0.00350124f $X=11.71 $Y=0.58
+ $X2=0 $Y2=0
cc_988 N_A_2082_446#_c_1463_n N_A_1824_74#_c_1582_n 0.00386679f $X=12.06
+ $Y=0.855 $X2=0 $Y2=0
cc_989 N_A_2082_446#_c_1465_n N_A_1824_74#_c_1582_n 0.00324637f $X=12.145
+ $Y=1.58 $X2=0 $Y2=0
cc_990 N_A_2082_446#_c_1461_n N_A_1824_74#_c_1583_n 0.00573299f $X=12.06
+ $Y=1.665 $X2=0 $Y2=0
cc_991 N_A_2082_446#_c_1465_n N_A_1824_74#_c_1583_n 0.00338011f $X=12.145
+ $Y=1.58 $X2=0 $Y2=0
cc_992 N_A_2082_446#_M1010_g N_A_1824_74#_c_1585_n 0.00114145f $X=10.705 $Y=0.58
+ $X2=0 $Y2=0
cc_993 N_A_2082_446#_M1005_g N_A_1824_74#_c_1595_n 0.00128633f $X=10.5 $Y=2.75
+ $X2=0 $Y2=0
cc_994 N_A_2082_446#_c_1528_p N_A_1824_74#_c_1595_n 0.0025825f $X=10.85 $Y=2.475
+ $X2=0 $Y2=0
cc_995 N_A_2082_446#_M1010_g N_A_1824_74#_c_1586_n 0.00142814f $X=10.705 $Y=0.58
+ $X2=0 $Y2=0
cc_996 N_A_2082_446#_M1010_g N_A_1824_74#_c_1587_n 0.00172861f $X=10.705 $Y=0.58
+ $X2=0 $Y2=0
cc_997 N_A_2082_446#_c_1469_n N_A_1824_74#_c_1587_n 0.00204272f $X=10.63 $Y=2.38
+ $X2=0 $Y2=0
cc_998 N_A_2082_446#_c_1528_p N_A_1824_74#_c_1587_n 0.0103498f $X=10.85 $Y=2.475
+ $X2=0 $Y2=0
cc_999 N_A_2082_446#_c_1466_n N_A_1824_74#_c_1587_n 0.0747982f $X=10.685
+ $Y=1.535 $X2=0 $Y2=0
cc_1000 N_A_2082_446#_c_1467_n N_A_1824_74#_c_1587_n 0.0114396f $X=10.685
+ $Y=1.535 $X2=0 $Y2=0
cc_1001 N_A_2082_446#_c_1463_n N_A_1824_74#_c_1588_n 0.00108154f $X=12.06
+ $Y=0.855 $X2=0 $Y2=0
cc_1002 N_A_2082_446#_c_1464_n N_A_1824_74#_c_1588_n 0.0272174f $X=11.875
+ $Y=0.855 $X2=0 $Y2=0
cc_1003 N_A_2082_446#_c_1465_n N_A_1824_74#_c_1588_n 0.0227002f $X=12.145
+ $Y=1.58 $X2=0 $Y2=0
cc_1004 N_A_2082_446#_M1010_g N_A_1824_74#_c_1590_n 0.0143673f $X=10.705 $Y=0.58
+ $X2=0 $Y2=0
cc_1005 N_A_2082_446#_c_1461_n N_A_1824_74#_c_1590_n 0.00732151f $X=12.06
+ $Y=1.665 $X2=0 $Y2=0
cc_1006 N_A_2082_446#_c_1466_n N_A_1824_74#_c_1590_n 0.0224547f $X=10.685
+ $Y=1.535 $X2=0 $Y2=0
cc_1007 N_A_2082_446#_c_1467_n N_A_1824_74#_c_1590_n 0.00598209f $X=10.685
+ $Y=1.535 $X2=0 $Y2=0
cc_1008 N_A_2082_446#_M1010_g N_A_1824_74#_c_1591_n 0.0019127f $X=10.705 $Y=0.58
+ $X2=0 $Y2=0
cc_1009 N_A_2082_446#_c_1461_n N_A_1824_74#_c_1591_n 0.06452f $X=12.06 $Y=1.665
+ $X2=0 $Y2=0
cc_1010 N_A_2082_446#_c_1466_n N_A_1824_74#_c_1591_n 0.00326018f $X=10.685
+ $Y=1.535 $X2=0 $Y2=0
cc_1011 N_A_2082_446#_c_1467_n N_A_1824_74#_c_1591_n 2.45278e-19 $X=10.685
+ $Y=1.535 $X2=0 $Y2=0
cc_1012 N_A_2082_446#_c_1465_n N_A_2495_392#_c_1719_n 0.0135871f $X=12.145
+ $Y=1.58 $X2=0 $Y2=0
cc_1013 N_A_2082_446#_c_1461_n N_A_2495_392#_c_1721_n 0.0058056f $X=12.06
+ $Y=1.665 $X2=0 $Y2=0
cc_1014 N_A_2082_446#_c_1461_n N_A_2495_392#_c_1722_n 0.00268745f $X=12.06
+ $Y=1.665 $X2=0 $Y2=0
cc_1015 N_A_2082_446#_c_1465_n N_A_2495_392#_c_1722_n 0.0131081f $X=12.145
+ $Y=1.58 $X2=0 $Y2=0
cc_1016 N_A_2082_446#_c_1472_n N_VPWR_M1005_d 0.00372166f $X=11.41 $Y=2.475
+ $X2=0 $Y2=0
cc_1017 N_A_2082_446#_c_1528_p N_VPWR_M1005_d 0.00220205f $X=10.85 $Y=2.475
+ $X2=0 $Y2=0
cc_1018 N_A_2082_446#_c_1461_n N_VPWR_c_1782_n 0.0235807f $X=12.06 $Y=1.665
+ $X2=0 $Y2=0
cc_1019 N_A_2082_446#_c_1472_n N_VPWR_c_1782_n 0.0116128f $X=11.41 $Y=2.475
+ $X2=0 $Y2=0
cc_1020 N_A_2082_446#_c_1473_n N_VPWR_c_1782_n 0.0142276f $X=11.575 $Y=2.75
+ $X2=0 $Y2=0
cc_1021 N_A_2082_446#_c_1473_n N_VPWR_c_1790_n 0.0143153f $X=11.575 $Y=2.75
+ $X2=0 $Y2=0
cc_1022 N_A_2082_446#_M1005_g N_VPWR_c_1795_n 0.00461464f $X=10.5 $Y=2.75 $X2=0
+ $Y2=0
cc_1023 N_A_2082_446#_M1005_g N_VPWR_c_1801_n 0.00963833f $X=10.5 $Y=2.75 $X2=0
+ $Y2=0
cc_1024 N_A_2082_446#_c_1469_n N_VPWR_c_1801_n 0.00120202f $X=10.63 $Y=2.38
+ $X2=0 $Y2=0
cc_1025 N_A_2082_446#_c_1472_n N_VPWR_c_1801_n 0.0277252f $X=11.41 $Y=2.475
+ $X2=0 $Y2=0
cc_1026 N_A_2082_446#_c_1528_p N_VPWR_c_1801_n 0.0200749f $X=10.85 $Y=2.475
+ $X2=0 $Y2=0
cc_1027 N_A_2082_446#_c_1473_n N_VPWR_c_1801_n 0.0102623f $X=11.575 $Y=2.75
+ $X2=0 $Y2=0
cc_1028 N_A_2082_446#_M1005_g N_VPWR_c_1777_n 0.00908061f $X=10.5 $Y=2.75 $X2=0
+ $Y2=0
cc_1029 N_A_2082_446#_c_1472_n N_VPWR_c_1777_n 0.00656614f $X=11.41 $Y=2.475
+ $X2=0 $Y2=0
cc_1030 N_A_2082_446#_c_1528_p N_VPWR_c_1777_n 0.00115936f $X=10.85 $Y=2.475
+ $X2=0 $Y2=0
cc_1031 N_A_2082_446#_c_1473_n N_VPWR_c_1777_n 0.0117766f $X=11.575 $Y=2.75
+ $X2=0 $Y2=0
cc_1032 N_A_2082_446#_c_1463_n N_VGND_M1029_s 0.00405314f $X=12.06 $Y=0.855
+ $X2=0 $Y2=0
cc_1033 N_A_2082_446#_c_1465_n N_VGND_M1029_s 8.04296e-19 $X=12.145 $Y=1.58
+ $X2=0 $Y2=0
cc_1034 N_A_2082_446#_M1010_g N_VGND_c_2140_n 0.0119771f $X=10.705 $Y=0.58 $X2=0
+ $Y2=0
cc_1035 N_A_2082_446#_c_1462_n N_VGND_c_2140_n 0.0140354f $X=11.71 $Y=0.58 $X2=0
+ $Y2=0
cc_1036 N_A_2082_446#_c_1464_n N_VGND_c_2140_n 0.00142029f $X=11.875 $Y=0.855
+ $X2=0 $Y2=0
cc_1037 N_A_2082_446#_c_1462_n N_VGND_c_2141_n 0.0168546f $X=11.71 $Y=0.58 $X2=0
+ $Y2=0
cc_1038 N_A_2082_446#_c_1463_n N_VGND_c_2141_n 0.0109002f $X=12.06 $Y=0.855
+ $X2=0 $Y2=0
cc_1039 N_A_2082_446#_M1010_g N_VGND_c_2151_n 0.00383152f $X=10.705 $Y=0.58
+ $X2=0 $Y2=0
cc_1040 N_A_2082_446#_c_1462_n N_VGND_c_2152_n 0.014415f $X=11.71 $Y=0.58 $X2=0
+ $Y2=0
cc_1041 N_A_2082_446#_M1010_g N_VGND_c_2159_n 0.0075725f $X=10.705 $Y=0.58 $X2=0
+ $Y2=0
cc_1042 N_A_2082_446#_c_1462_n N_VGND_c_2159_n 0.0119404f $X=11.71 $Y=0.58 $X2=0
+ $Y2=0
cc_1043 N_A_2082_446#_c_1463_n N_VGND_c_2159_n 0.0092009f $X=12.06 $Y=0.855
+ $X2=0 $Y2=0
cc_1044 N_A_1824_74#_M1037_g N_A_2495_392#_c_1726_n 0.00376928f $X=12.385
+ $Y=2.46 $X2=0 $Y2=0
cc_1045 N_A_1824_74#_c_1584_n N_A_2495_392#_c_1726_n 0.00239754f $X=12.295
+ $Y=1.095 $X2=0 $Y2=0
cc_1046 N_A_1824_74#_M1037_g N_A_2495_392#_c_1727_n 0.0106267f $X=12.385 $Y=2.46
+ $X2=0 $Y2=0
cc_1047 N_A_1824_74#_c_1582_n N_A_2495_392#_c_1719_n 0.00769864f $X=12.485
+ $Y=1.095 $X2=0 $Y2=0
cc_1048 N_A_1824_74#_c_1584_n N_A_2495_392#_c_1719_n 0.00167437f $X=12.295
+ $Y=1.095 $X2=0 $Y2=0
cc_1049 N_A_1824_74#_M1037_g N_A_2495_392#_c_1721_n 0.00969578f $X=12.385
+ $Y=2.46 $X2=0 $Y2=0
cc_1050 N_A_1824_74#_c_1584_n N_A_2495_392#_c_1722_n 0.00471821f $X=12.295
+ $Y=1.095 $X2=0 $Y2=0
cc_1051 N_A_1824_74#_c_1584_n N_A_2495_392#_c_1723_n 0.00503519f $X=12.295
+ $Y=1.095 $X2=0 $Y2=0
cc_1052 N_A_1824_74#_M1024_g N_VPWR_c_1782_n 0.0162693f $X=11.8 $Y=2.75 $X2=0
+ $Y2=0
cc_1053 N_A_1824_74#_c_1579_n N_VPWR_c_1782_n 7.36409e-19 $X=12.295 $Y=1.26
+ $X2=0 $Y2=0
cc_1054 N_A_1824_74#_M1037_g N_VPWR_c_1782_n 0.00369333f $X=12.385 $Y=2.46 $X2=0
+ $Y2=0
cc_1055 N_A_1824_74#_M1037_g N_VPWR_c_1783_n 0.00470925f $X=12.385 $Y=2.46 $X2=0
+ $Y2=0
cc_1056 N_A_1824_74#_M1024_g N_VPWR_c_1790_n 0.005209f $X=11.8 $Y=2.75 $X2=0
+ $Y2=0
cc_1057 N_A_1824_74#_c_1595_n N_VPWR_c_1795_n 0.0193246f $X=10.22 $Y=2.685 $X2=0
+ $Y2=0
cc_1058 N_A_1824_74#_c_1596_n N_VPWR_c_1795_n 0.00809057f $X=9.6 $Y=2.685 $X2=0
+ $Y2=0
cc_1059 N_A_1824_74#_M1037_g N_VPWR_c_1796_n 0.005209f $X=12.385 $Y=2.46 $X2=0
+ $Y2=0
cc_1060 N_A_1824_74#_M1024_g N_VPWR_c_1777_n 0.00983707f $X=11.8 $Y=2.75 $X2=0
+ $Y2=0
cc_1061 N_A_1824_74#_M1037_g N_VPWR_c_1777_n 0.00987945f $X=12.385 $Y=2.46 $X2=0
+ $Y2=0
cc_1062 N_A_1824_74#_c_1595_n N_VPWR_c_1777_n 0.0252724f $X=10.22 $Y=2.685 $X2=0
+ $Y2=0
cc_1063 N_A_1824_74#_c_1596_n N_VPWR_c_1777_n 0.00934828f $X=9.6 $Y=2.685 $X2=0
+ $Y2=0
cc_1064 N_A_1824_74#_c_1595_n A_2040_508# 0.00142071f $X=10.22 $Y=2.685
+ $X2=-0.19 $Y2=-0.245
cc_1065 N_A_1824_74#_M1018_g N_VGND_c_2140_n 0.00182082f $X=11.495 $Y=0.58 $X2=0
+ $Y2=0
cc_1066 N_A_1824_74#_c_1585_n N_VGND_c_2140_n 0.014224f $X=10.22 $Y=0.645 $X2=0
+ $Y2=0
cc_1067 N_A_1824_74#_c_1590_n N_VGND_c_2140_n 0.0229174f $X=11.02 $Y=1.22 $X2=0
+ $Y2=0
cc_1068 N_A_1824_74#_M1018_g N_VGND_c_2141_n 0.00324482f $X=11.495 $Y=0.58 $X2=0
+ $Y2=0
cc_1069 N_A_1824_74#_c_1579_n N_VGND_c_2141_n 0.00356476f $X=12.295 $Y=1.26
+ $X2=0 $Y2=0
cc_1070 N_A_1824_74#_c_1582_n N_VGND_c_2141_n 0.00936719f $X=12.485 $Y=1.095
+ $X2=0 $Y2=0
cc_1071 N_A_1824_74#_c_1582_n N_VGND_c_2142_n 0.00296233f $X=12.485 $Y=1.095
+ $X2=0 $Y2=0
cc_1072 N_A_1824_74#_c_1585_n N_VGND_c_2151_n 0.0249458f $X=10.22 $Y=0.645 $X2=0
+ $Y2=0
cc_1073 N_A_1824_74#_M1018_g N_VGND_c_2152_n 0.00434272f $X=11.495 $Y=0.58 $X2=0
+ $Y2=0
cc_1074 N_A_1824_74#_c_1582_n N_VGND_c_2153_n 0.00383152f $X=12.485 $Y=1.095
+ $X2=0 $Y2=0
cc_1075 N_A_1824_74#_M1018_g N_VGND_c_2159_n 0.00825669f $X=11.495 $Y=0.58 $X2=0
+ $Y2=0
cc_1076 N_A_1824_74#_c_1582_n N_VGND_c_2159_n 0.00762539f $X=12.485 $Y=1.095
+ $X2=0 $Y2=0
cc_1077 N_A_1824_74#_c_1585_n N_VGND_c_2159_n 0.0310203f $X=10.22 $Y=0.645 $X2=0
+ $Y2=0
cc_1078 N_A_2495_392#_c_1726_n N_VPWR_c_1782_n 0.0405667f $X=12.61 $Y=2.105
+ $X2=0 $Y2=0
cc_1079 N_A_2495_392#_M1001_g N_VPWR_c_1783_n 0.0207145f $X=13.395 $Y=2.4 $X2=0
+ $Y2=0
cc_1080 N_A_2495_392#_M1041_g N_VPWR_c_1783_n 7.17218e-19 $X=13.845 $Y=2.4 $X2=0
+ $Y2=0
cc_1081 N_A_2495_392#_c_1720_n N_VPWR_c_1783_n 0.0253895f $X=13.19 $Y=1.465
+ $X2=0 $Y2=0
cc_1082 N_A_2495_392#_c_1721_n N_VPWR_c_1783_n 0.077754f $X=12.61 $Y=1.94 $X2=0
+ $Y2=0
cc_1083 N_A_2495_392#_c_1723_n N_VPWR_c_1783_n 0.00645758f $X=13.845 $Y=1.465
+ $X2=0 $Y2=0
cc_1084 N_A_2495_392#_M1041_g N_VPWR_c_1785_n 0.00540173f $X=13.845 $Y=2.4 $X2=0
+ $Y2=0
cc_1085 N_A_2495_392#_c_1723_n N_VPWR_c_1785_n 9.39066e-19 $X=13.845 $Y=1.465
+ $X2=0 $Y2=0
cc_1086 N_A_2495_392#_c_1727_n N_VPWR_c_1796_n 0.014549f $X=12.61 $Y=2.815 $X2=0
+ $Y2=0
cc_1087 N_A_2495_392#_M1001_g N_VPWR_c_1797_n 0.00460063f $X=13.395 $Y=2.4 $X2=0
+ $Y2=0
cc_1088 N_A_2495_392#_M1041_g N_VPWR_c_1797_n 0.005209f $X=13.845 $Y=2.4 $X2=0
+ $Y2=0
cc_1089 N_A_2495_392#_M1001_g N_VPWR_c_1777_n 0.00908554f $X=13.395 $Y=2.4 $X2=0
+ $Y2=0
cc_1090 N_A_2495_392#_M1041_g N_VPWR_c_1777_n 0.00985497f $X=13.845 $Y=2.4 $X2=0
+ $Y2=0
cc_1091 N_A_2495_392#_c_1727_n N_VPWR_c_1777_n 0.0119743f $X=12.61 $Y=2.815
+ $X2=0 $Y2=0
cc_1092 N_A_2495_392#_M1001_g N_Q_c_2116_n 0.00554343f $X=13.395 $Y=2.4 $X2=0
+ $Y2=0
cc_1093 N_A_2495_392#_M1041_g N_Q_c_2116_n 0.0245288f $X=13.845 $Y=2.4 $X2=0
+ $Y2=0
cc_1094 N_A_2495_392#_c_1723_n N_Q_c_2116_n 0.0194596f $X=13.845 $Y=1.465 $X2=0
+ $Y2=0
cc_1095 N_A_2495_392#_M1003_g Q 0.0138248f $X=13.475 $Y=0.74 $X2=0 $Y2=0
cc_1096 N_A_2495_392#_M1030_g Q 0.0162403f $X=13.905 $Y=0.74 $X2=0 $Y2=0
cc_1097 N_A_2495_392#_c_1719_n Q 0.00465944f $X=12.7 $Y=0.515 $X2=0 $Y2=0
cc_1098 N_A_2495_392#_M1003_g Q 0.0018463f $X=13.475 $Y=0.74 $X2=0 $Y2=0
cc_1099 N_A_2495_392#_M1030_g Q 0.00299044f $X=13.905 $Y=0.74 $X2=0 $Y2=0
cc_1100 N_A_2495_392#_c_1720_n Q 0.02585f $X=13.19 $Y=1.465 $X2=0 $Y2=0
cc_1101 N_A_2495_392#_c_1723_n Q 0.0155405f $X=13.845 $Y=1.465 $X2=0 $Y2=0
cc_1102 N_A_2495_392#_c_1719_n N_VGND_c_2141_n 0.0101431f $X=12.7 $Y=0.515 $X2=0
+ $Y2=0
cc_1103 N_A_2495_392#_M1003_g N_VGND_c_2142_n 0.00647412f $X=13.475 $Y=0.74
+ $X2=0 $Y2=0
cc_1104 N_A_2495_392#_c_1719_n N_VGND_c_2142_n 0.0505719f $X=12.7 $Y=0.515 $X2=0
+ $Y2=0
cc_1105 N_A_2495_392#_c_1720_n N_VGND_c_2142_n 0.0209147f $X=13.19 $Y=1.465
+ $X2=0 $Y2=0
cc_1106 N_A_2495_392#_c_1723_n N_VGND_c_2142_n 0.00593115f $X=13.845 $Y=1.465
+ $X2=0 $Y2=0
cc_1107 N_A_2495_392#_M1030_g N_VGND_c_2144_n 0.00647412f $X=13.905 $Y=0.74
+ $X2=0 $Y2=0
cc_1108 N_A_2495_392#_c_1719_n N_VGND_c_2153_n 0.0115122f $X=12.7 $Y=0.515 $X2=0
+ $Y2=0
cc_1109 N_A_2495_392#_M1003_g N_VGND_c_2154_n 0.00434272f $X=13.475 $Y=0.74
+ $X2=0 $Y2=0
cc_1110 N_A_2495_392#_M1030_g N_VGND_c_2154_n 0.00434272f $X=13.905 $Y=0.74
+ $X2=0 $Y2=0
cc_1111 N_A_2495_392#_M1003_g N_VGND_c_2159_n 0.00825283f $X=13.475 $Y=0.74
+ $X2=0 $Y2=0
cc_1112 N_A_2495_392#_M1030_g N_VGND_c_2159_n 0.00823942f $X=13.905 $Y=0.74
+ $X2=0 $Y2=0
cc_1113 N_A_2495_392#_c_1719_n N_VGND_c_2159_n 0.0095288f $X=12.7 $Y=0.515 $X2=0
+ $Y2=0
cc_1114 N_VPWR_c_1778_n N_A_390_81#_c_1956_n 0.00942884f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1115 N_VPWR_c_1793_n N_A_390_81#_c_1956_n 0.0233446f $X=3.095 $Y=3.33 $X2=0
+ $Y2=0
cc_1116 N_VPWR_c_1798_n N_A_390_81#_c_1956_n 0.0172244f $X=0.78 $Y=2.465 $X2=0
+ $Y2=0
cc_1117 N_VPWR_c_1777_n N_A_390_81#_c_1956_n 0.0125323f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1118 N_VPWR_M1039_d N_A_390_81#_c_1957_n 0.00184188f $X=3.125 $Y=2.415 $X2=0
+ $Y2=0
cc_1119 N_VPWR_c_1778_n N_A_390_81#_c_1957_n 0.016715f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1120 N_VPWR_c_1777_n N_A_390_81#_c_1957_n 0.0228237f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1121 N_VPWR_c_1798_n N_A_390_81#_c_1958_n 0.00553242f $X=0.78 $Y=2.465 $X2=0
+ $Y2=0
cc_1122 N_VPWR_M1027_d N_A_390_81#_c_1960_n 0.00371121f $X=4.735 $Y=1.935 $X2=0
+ $Y2=0
cc_1123 N_VPWR_c_1779_n N_A_390_81#_c_1960_n 0.016342f $X=4.87 $Y=2.88 $X2=0
+ $Y2=0
cc_1124 N_VPWR_c_1786_n N_A_390_81#_c_1960_n 0.0103633f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1125 N_VPWR_c_1788_n N_A_390_81#_c_1960_n 0.0100794f $X=7.15 $Y=3.33 $X2=0
+ $Y2=0
cc_1126 N_VPWR_c_1777_n N_A_390_81#_c_1960_n 0.0373206f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1127 N_VPWR_c_1788_n N_A_390_81#_c_1961_n 0.0053294f $X=7.15 $Y=3.33 $X2=0
+ $Y2=0
cc_1128 N_VPWR_c_1777_n N_A_390_81#_c_1961_n 0.00671812f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1129 N_VPWR_c_1778_n N_A_390_81#_c_1965_n 0.0141328f $X=3.26 $Y=2.79 $X2=0
+ $Y2=0
cc_1130 N_VPWR_c_1786_n N_A_390_81#_c_1965_n 0.0270976f $X=4.705 $Y=3.33 $X2=0
+ $Y2=0
cc_1131 N_VPWR_c_1777_n N_A_390_81#_c_1965_n 0.0203696f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1132 N_VPWR_c_1783_n N_Q_c_2116_n 0.0412253f $X=13.17 $Y=1.985 $X2=0 $Y2=0
cc_1133 N_VPWR_c_1785_n N_Q_c_2116_n 0.0435456f $X=14.12 $Y=1.985 $X2=0 $Y2=0
cc_1134 N_VPWR_c_1797_n N_Q_c_2116_n 0.0114255f $X=13.955 $Y=3.33 $X2=0 $Y2=0
cc_1135 N_VPWR_c_1777_n N_Q_c_2116_n 0.00938892f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1136 N_A_390_81#_c_1957_n A_517_483# 0.00483994f $X=3.445 $Y=2.43 $X2=-0.19
+ $Y2=-0.245
cc_1137 N_A_390_81#_M1015_d N_noxref_24_c_2273_n 0.0102044f $X=1.95 $Y=0.405
+ $X2=0 $Y2=0
cc_1138 N_A_390_81#_c_1947_n N_noxref_24_c_2273_n 0.0420252f $X=2.875 $Y=0.72
+ $X2=0 $Y2=0
cc_1139 N_A_390_81#_c_1947_n N_noxref_24_c_2289_n 0.0147071f $X=2.875 $Y=0.72
+ $X2=0 $Y2=0
cc_1140 N_A_390_81#_c_1949_n N_noxref_24_c_2289_n 0.00859185f $X=3.445 $Y=1.225
+ $X2=0 $Y2=0
cc_1141 N_A_390_81#_c_1947_n noxref_26 0.00129814f $X=2.875 $Y=0.72 $X2=-0.19
+ $Y2=-0.245
cc_1142 Q N_VGND_c_2142_n 0.0294122f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1143 Q N_VGND_c_2144_n 0.0294122f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1144 Q N_VGND_c_2154_n 0.0144922f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1145 Q N_VGND_c_2159_n 0.0118826f $X=13.595 $Y=0.47 $X2=0 $Y2=0
cc_1146 N_VGND_c_2138_n N_noxref_24_c_2273_n 0.010604f $X=3.79 $Y=0.615 $X2=0
+ $Y2=0
cc_1147 N_VGND_c_2145_n N_noxref_24_c_2273_n 0.128699f $X=3.665 $Y=0 $X2=0 $Y2=0
cc_1148 N_VGND_c_2159_n N_noxref_24_c_2273_n 0.0746443f $X=14.16 $Y=0 $X2=0
+ $Y2=0
cc_1149 N_VGND_c_2137_n N_noxref_24_c_2274_n 0.0259561f $X=0.71 $Y=0.555 $X2=0
+ $Y2=0
cc_1150 N_VGND_c_2145_n N_noxref_24_c_2274_n 0.0225398f $X=3.665 $Y=0 $X2=0
+ $Y2=0
cc_1151 N_VGND_c_2159_n N_noxref_24_c_2274_n 0.0125704f $X=14.16 $Y=0 $X2=0
+ $Y2=0
cc_1152 N_noxref_24_c_2273_n noxref_25 0.00198134f $X=3.215 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1153 N_noxref_24_c_2273_n noxref_26 0.00134156f $X=3.215 $Y=0.34 $X2=-0.19
+ $Y2=-0.245

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 a_34_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.3e+11p pd=5.06e+06u as=6.766e+11p ps=5.55e+06u
M1001 X a_194_136# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1002 a_122_136# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=5.6545e+11p ps=5.75e+06u
M1003 X a_194_136# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1004 VGND a_272_110# a_194_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.496e+11p ps=2.06e+06u
M1005 a_194_136# a_272_110# a_34_392# VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
M1006 VPWR A2 a_34_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR B1_N a_272_110# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.184e+11p ps=2.2e+06u
M1008 VGND B1_N a_272_110# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1009 a_194_136# A1 a_122_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

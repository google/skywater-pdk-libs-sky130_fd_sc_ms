# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__dfrtp_1
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.000000 0.515000 2.170000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.591700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  9.725000 1.885000 10.425000 2.980000 ;
        RECT 10.165000 0.350000 10.495000 1.130000 ;
        RECT 10.165000 1.130000 10.425000 1.885000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.055000 1.920000 1.345000 1.965000 ;
        RECT 1.055000 1.965000 8.065000 2.105000 ;
        RECT 1.055000 2.105000 1.345000 2.150000 ;
        RECT 4.895000 1.920000 5.185000 1.965000 ;
        RECT 4.895000 2.105000 5.185000 2.150000 ;
        RECT 7.775000 1.920000 8.065000 1.965000 ;
        RECT 7.775000 2.105000 8.065000 2.150000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.261000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.795000 1.310000 2.275000 1.775000 ;
        RECT 2.045000 1.775000 2.275000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.040000 0.085000 ;
      RECT  0.000000  3.245000 11.040000 3.415000 ;
      RECT  0.105000  2.520000  0.355000 3.245000 ;
      RECT  0.130000  0.370000  0.460000 0.660000 ;
      RECT  0.130000  0.660000  0.855000 0.830000 ;
      RECT  0.555000  2.520000  3.290000 2.560000 ;
      RECT  0.555000  2.560000  0.860000 2.605000 ;
      RECT  0.555000  2.605000  0.835000 2.640000 ;
      RECT  0.555000  2.640000  0.810000 2.980000 ;
      RECT  0.685000  0.830000  0.855000 2.310000 ;
      RECT  0.685000  2.310000  1.435000 2.335000 ;
      RECT  0.685000  2.335000  1.465000 2.360000 ;
      RECT  0.685000  2.360000  1.490000 2.375000 ;
      RECT  0.685000  2.375000  1.510000 2.390000 ;
      RECT  0.685000  2.390000  1.530000 2.410000 ;
      RECT  0.685000  2.410000  3.290000 2.520000 ;
      RECT  0.980000  2.730000  1.310000 3.245000 ;
      RECT  1.025000  1.130000  1.285000 2.140000 ;
      RECT  1.030000  0.085000  1.280000 0.830000 ;
      RECT  1.405000  2.560000  3.290000 2.570000 ;
      RECT  1.405000  2.570000  1.925000 2.575000 ;
      RECT  1.405000  2.575000  1.910000 2.580000 ;
      RECT  1.405000  2.580000  1.890000 2.585000 ;
      RECT  1.435000  2.585000  1.890000 2.590000 ;
      RECT  1.435000  2.590000  1.860000 2.610000 ;
      RECT  1.455000  0.350000  1.840000 0.970000 ;
      RECT  1.455000  0.970000  2.505000 0.975000 ;
      RECT  1.455000  0.975000  2.695000 1.140000 ;
      RECT  1.455000  1.140000  1.625000 1.945000 ;
      RECT  1.455000  1.945000  1.865000 2.140000 ;
      RECT  1.615000  2.140000  1.865000 2.205000 ;
      RECT  1.615000  2.205000  1.785000 2.240000 ;
      RECT  1.835000  2.405000  3.290000 2.410000 ;
      RECT  1.850000  2.400000  3.290000 2.405000 ;
      RECT  1.870000  2.390000  3.290000 2.400000 ;
      RECT  1.895000  2.375000  3.290000 2.390000 ;
      RECT  1.985000  2.740000  2.315000 3.245000 ;
      RECT  2.060000  0.085000  2.390000 0.800000 ;
      RECT  2.445000  1.140000  2.695000 1.490000 ;
      RECT  2.445000  1.490000  2.775000 1.695000 ;
      RECT  2.445000  1.865000  3.420000 1.985000 ;
      RECT  2.445000  1.985000  3.060000 2.035000 ;
      RECT  2.445000  2.035000  2.775000 2.205000 ;
      RECT  2.560000  0.330000  4.440000 0.500000 ;
      RECT  2.560000  0.500000  3.035000 0.805000 ;
      RECT  2.865000  0.805000  3.035000 1.195000 ;
      RECT  2.865000  1.195000  3.115000 1.345000 ;
      RECT  2.900000  1.820000  3.420000 1.865000 ;
      RECT  2.945000  1.345000  3.115000 1.560000 ;
      RECT  2.945000  1.560000  3.420000 1.820000 ;
      RECT  3.010000  2.205000  3.760000 2.325000 ;
      RECT  3.010000  2.325000  3.335000 2.370000 ;
      RECT  3.010000  2.370000  3.290000 2.375000 ;
      RECT  3.010000  2.570000  3.290000 2.725000 ;
      RECT  3.185000  2.155000  3.760000 2.205000 ;
      RECT  3.205000  0.670000  3.455000 1.045000 ;
      RECT  3.285000  1.045000  3.455000 1.220000 ;
      RECT  3.285000  1.220000  3.760000 1.390000 ;
      RECT  3.460000  2.495000  5.250000 2.570000 ;
      RECT  3.460000  2.570000  4.215000 2.725000 ;
      RECT  3.590000  1.390000  3.760000 2.155000 ;
      RECT  3.625000  0.670000  4.100000 1.050000 ;
      RECT  3.930000  1.050000  4.100000 2.400000 ;
      RECT  3.930000  2.400000  5.250000 2.495000 ;
      RECT  4.270000  0.500000  4.440000 0.565000 ;
      RECT  4.270000  0.565000  5.650000 0.735000 ;
      RECT  4.270000  0.905000  6.150000 1.075000 ;
      RECT  4.270000  1.075000  4.445000 2.125000 ;
      RECT  4.385000  2.740000  4.715000 3.245000 ;
      RECT  4.615000  1.245000  5.650000 1.575000 ;
      RECT  4.615000  1.575000  4.785000 2.320000 ;
      RECT  4.615000  2.320000  5.250000 2.400000 ;
      RECT  4.915000  0.085000  5.310000 0.395000 ;
      RECT  4.955000  1.795000  5.285000 2.150000 ;
      RECT  5.480000  0.255000  7.420000 0.425000 ;
      RECT  5.480000  0.425000  5.650000 0.565000 ;
      RECT  5.480000  1.745000  5.810000 3.245000 ;
      RECT  5.820000  0.665000  6.150000 0.905000 ;
      RECT  5.820000  1.075000  6.150000 1.130000 ;
      RECT  5.980000  1.130000  6.150000 1.865000 ;
      RECT  5.980000  1.865000  6.310000 2.755000 ;
      RECT  6.320000  0.595000  7.080000 0.845000 ;
      RECT  6.320000  0.845000  6.490000 1.515000 ;
      RECT  6.320000  1.515000  6.650000 1.685000 ;
      RECT  6.480000  1.685000  6.650000 2.475000 ;
      RECT  6.480000  2.475000  7.635000 2.805000 ;
      RECT  6.690000  1.015000  7.420000 1.345000 ;
      RECT  6.965000  1.345000  7.295000 2.305000 ;
      RECT  7.250000  0.425000  7.420000 1.015000 ;
      RECT  7.465000  1.515000  8.850000 1.685000 ;
      RECT  7.465000  1.685000  7.635000 2.475000 ;
      RECT  7.590000  1.015000  9.190000 1.185000 ;
      RECT  7.590000  1.185000  7.920000 1.345000 ;
      RECT  7.745000  0.085000  8.075000 0.845000 ;
      RECT  7.805000  1.920000  8.345000 2.255000 ;
      RECT  7.805000  2.445000  8.135000 3.245000 ;
      RECT  8.320000  2.445000  8.685000 2.905000 ;
      RECT  8.515000  1.855000  9.190000 2.025000 ;
      RECT  8.515000  2.025000  8.685000 2.445000 ;
      RECT  8.520000  1.355000  8.850000 1.515000 ;
      RECT  8.615000  0.385000  8.945000 1.015000 ;
      RECT  8.855000  2.195000  9.185000 3.245000 ;
      RECT  9.020000  1.185000  9.190000 1.855000 ;
      RECT  9.175000  0.085000  9.425000 0.845000 ;
      RECT  9.385000  1.385000  9.935000 1.715000 ;
      RECT  9.385000  1.715000  9.555000 2.905000 ;
      RECT  9.605000  0.350000  9.935000 1.385000 ;
      RECT 10.595000  1.820000 10.925000 3.245000 ;
      RECT 10.675000  0.085000 10.925000 1.130000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  1.950000  1.285000 2.120000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  1.950000  5.125000 2.120000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.950000  8.005000 2.120000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
  END
END sky130_fd_sc_ms__dfrtp_1

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfstp_4 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
M1000 Q a_2580_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=2.9103e+12p ps=2.649e+07u
M1001 Q a_2580_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=5.291e+11p pd=4.39e+06u as=2.27325e+12p ps=1.996e+07u
M1002 a_1017_81# a_616_74# a_291_464# VNB nlowvt w=420000u l=150000u
+  ad=2.226e+11p pd=1.9e+06u as=3.592e+11p ps=3.44e+06u
M1003 VGND SET_B a_1445_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1004 a_2227_74# a_2191_180# a_2149_74# VNB nlowvt w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=1.008e+11p ps=1.32e+06u
M1005 VGND a_1823_524# a_2580_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1006 a_1823_524# a_803_74# a_1677_74# VNB nlowvt w=640000u l=150000u
+  ad=3.963e+11p pd=3.85e+06u as=3.584e+11p ps=3.68e+06u
M1007 VPWR a_2191_180# a_2106_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.869e+11p ps=1.73e+06u
M1008 a_1017_81# a_803_74# a_291_464# VPB pshort w=420000u l=180000u
+  ad=1.8235e+11p pd=1.93e+06u as=4.056e+11p ps=3.58e+06u
M1009 a_2580_74# a_1823_524# VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1010 VPWR a_1201_55# a_1143_495# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.6975e+11p ps=1.87e+06u
M1011 a_1823_524# SET_B VPWR VPB pshort w=420000u l=180000u
+  ad=5.793e+11p pd=5.97e+06u as=0p ps=0u
M1012 VGND a_1017_81# a_1677_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1143_495# a_616_74# a_1017_81# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_1823_524# a_2580_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Q a_2580_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_417_74# SCE a_291_464# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1017 VGND SCD a_417_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_1201_55# a_1153_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1019 a_1153_81# a_803_74# a_1017_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_803_74# a_616_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1021 VGND a_2580_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1445_74# a_1017_81# a_1201_55# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1023 VPWR SET_B a_1201_55# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1024 a_1623_373# a_1017_81# VPWR VPB pshort w=840000u l=180000u
+  ad=4.536e+11p pd=4.44e+06u as=0p ps=0u
M1025 VGND CLK a_616_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1026 a_2149_74# a_616_74# a_1823_524# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_417_464# a_27_74# a_291_464# VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1028 a_1201_55# a_1017_81# VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_1017_81# a_1623_373# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR a_2580_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND a_2580_74# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_2106_508# a_803_74# a_1823_524# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR SCE a_27_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1034 a_207_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1035 VPWR SCD a_417_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1677_74# a_803_74# a_1823_524# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR a_1823_524# a_2191_180# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1038 VGND SET_B a_2227_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_2191_180# a_1823_524# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1040 a_222_74# a_27_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1041 a_291_464# D a_222_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VPWR CLK a_616_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1043 a_1623_373# a_616_74# a_1823_524# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_291_464# D a_207_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VGND SCE a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1046 Q a_2580_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1047 a_1823_524# a_616_74# a_1623_373# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_803_74# a_616_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.088e+11p pd=2.9e+06u as=0p ps=0u
M1049 a_1677_74# a_1017_81# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1050 VPWR a_2580_74# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

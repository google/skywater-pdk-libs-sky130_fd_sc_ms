* NGSPICE file created from sky130_fd_sc_ms__o22a_4.ext - technology: sky130A

.subckt sky130_fd_sc_ms__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 VPWR A1 a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=2.0354e+12p pd=1.451e+07u as=5.9e+11p ps=5.18e+06u
M1001 a_119_392# A2 a_209_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=6.4e+11p ps=5.28e+06u
M1002 a_119_392# A1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_209_392# A2 a_119_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_209_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.44e+11p pd=5.63e+06u as=0p ps=0u
M1005 a_27_136# B1 a_209_392# VNB nlowvt w=640000u l=150000u
+  ad=1.0112e+12p pd=9.56e+06u as=3.616e+11p ps=3.69e+06u
M1006 VGND a_209_392# X VNB nlowvt w=740000u l=150000u
+  ad=1.1945e+12p pd=1.055e+07u as=4.144e+11p ps=4.08e+06u
M1007 X a_209_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_209_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_209_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_209_392# B2 a_27_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_209_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_136# B2 a_209_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_136# A2 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A2 a_27_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_209_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_136# A1 VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A1 a_27_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_209_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_519_392# B1 VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=0p ps=0u
M1020 a_209_392# B1 a_27_136# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR B1 a_519_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_519_392# B2 a_209_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_209_392# B2 a_519_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


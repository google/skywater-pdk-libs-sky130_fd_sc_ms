* File: sky130_fd_sc_ms__sdfrtn_1.pex.spice
* Created: Wed Sep  2 12:30:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SDFRTN_1%SCE 3 7 10 13 17 24 25 27 28 29 35 37
c70 24 0 8.65763e-20 $X=0.7 $Y=1.575
r71 34 37 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=2.385 $Y=1.12
+ $X2=2.615 $Y2=1.12
r72 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.385
+ $Y=1.12 $X2=2.385 $Y2=1.12
r73 29 35 5.91467 $w=4.53e-07 $l=2.25e-07 $layer=LI1_cond $X=2.16 $Y=1.182
+ $X2=2.385 $Y2=1.182
r74 28 29 3.02306 $w=4.53e-07 $l=1.15e-07 $layer=LI1_cond $X=2.045 $Y=1.182
+ $X2=2.16 $Y2=1.182
r75 27 28 9.38335 $w=4.53e-07 $l=1.7e-07 $layer=LI1_cond $X=1.875 $Y=1.267
+ $X2=2.045 $Y2=1.267
r76 25 32 46.8028 $w=4.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.642 $Y=1.575
+ $X2=0.642 $Y2=1.41
r77 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.7
+ $Y=1.575 $X2=0.7 $Y2=1.575
r78 22 24 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=1.495
+ $X2=0.7 $Y2=1.495
r79 22 27 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=0.865 $Y=1.495
+ $X2=1.875 $Y2=1.495
r80 15 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.615 $Y=0.955
+ $X2=2.615 $Y2=1.12
r81 15 17 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.615 $Y=0.955
+ $X2=2.615 $Y2=0.615
r82 9 25 7.12377 $w=4.45e-07 $l=5.7e-08 $layer=POLY_cond $X=0.642 $Y=1.632
+ $X2=0.642 $Y2=1.575
r83 9 10 37.2436 $w=4.45e-07 $l=2.98e-07 $layer=POLY_cond $X=0.642 $Y=1.632
+ $X2=0.642 $Y2=1.93
r84 7 32 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.495 $Y=0.65
+ $X2=0.495 $Y2=1.41
r85 1 10 15.786 $w=4.58e-07 $l=3.80682e-07 $layer=POLY_cond $X=0.955 $Y=2.08
+ $X2=0.642 $Y2=1.93
r86 1 13 217.677 $w=1.8e-07 $l=5.6e-07 $layer=POLY_cond $X=0.955 $Y=2.08
+ $X2=0.955 $Y2=2.64
r87 1 3 182.694 $w=1.8e-07 $l=4.7e-07 $layer=POLY_cond $X=0.505 $Y=2.17
+ $X2=0.505 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTN_1%A_27_88# 1 2 9 12 16 19 22 24 30 31 33 34
+ 36 37 38 41
c88 12 0 1.86156e-19 $X=2.28 $Y=2.64
r89 37 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.455 $Y=1.1
+ $X2=1.455 $Y2=0.935
r90 36 38 7.86356 $w=3.03e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=1.087
+ $X2=1.29 $Y2=1.087
r91 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.455
+ $Y=1.1 $X2=1.455 $Y2=1.1
r92 31 43 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=2.38 $Y=1.72 $X2=2.28
+ $Y2=1.72
r93 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.38
+ $Y=1.72 $X2=2.38 $Y2=1.72
r94 28 30 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=2.38 $Y=2.29
+ $X2=2.38 $Y2=1.72
r95 27 33 2.90107 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=1.145
+ $X2=0.28 $Y2=1.145
r96 27 38 49.3254 $w=1.88e-07 $l=8.45e-07 $layer=LI1_cond $X=0.445 $Y=1.145
+ $X2=1.29 $Y2=1.145
r97 25 34 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=2.375
+ $X2=0.24 $Y2=2.375
r98 24 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.215 $Y=2.375
+ $X2=2.38 $Y2=2.29
r99 24 25 120.695 $w=1.68e-07 $l=1.85e-06 $layer=LI1_cond $X=2.215 $Y=2.375
+ $X2=0.365 $Y2=2.375
r100 20 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.46
+ $X2=0.24 $Y2=2.375
r101 20 22 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.24 $Y=2.46
+ $X2=0.24 $Y2=2.465
r102 19 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.29
+ $X2=0.24 $Y2=2.375
r103 18 33 3.58697 $w=2.9e-07 $l=1.13248e-07 $layer=LI1_cond $X=0.24 $Y=1.24
+ $X2=0.28 $Y2=1.145
r104 18 19 48.4026 $w=2.48e-07 $l=1.05e-06 $layer=LI1_cond $X=0.24 $Y=1.24
+ $X2=0.24 $Y2=2.29
r105 14 33 3.58697 $w=2.9e-07 $l=9.5e-08 $layer=LI1_cond $X=0.28 $Y=1.05
+ $X2=0.28 $Y2=1.145
r106 14 16 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=0.28 $Y=1.05 $X2=0.28
+ $Y2=0.65
r107 10 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.28 $Y=1.885
+ $X2=2.28 $Y2=1.72
r108 10 12 293.476 $w=1.8e-07 $l=7.55e-07 $layer=POLY_cond $X=2.28 $Y=1.885
+ $X2=2.28 $Y2=2.64
r109 9 41 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.545 $Y=0.615
+ $X2=1.545 $Y2=0.935
r110 2 22 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.465
r111 1 16 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.44 $X2=0.28 $Y2=0.65
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTN_1%D 3 5 6 9 11 12 16 17
c39 17 0 1.86156e-19 $X=1.815 $Y=1.945
c40 6 0 8.65763e-20 $X=1.435 $Y=2.035
r41 16 19 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.815 $Y=1.945
+ $X2=1.815 $Y2=2.035
r42 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.945
+ $X2=1.815 $Y2=1.78
r43 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.815
+ $Y=1.945 $X2=1.815 $Y2=1.945
r44 12 17 4.57588 $w=3.38e-07 $l=1.35e-07 $layer=LI1_cond $X=1.68 $Y=1.95
+ $X2=1.815 $Y2=1.95
r45 11 12 16.2698 $w=3.38e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.95 $X2=1.68
+ $Y2=1.95
r46 9 18 597.372 $w=1.5e-07 $l=1.165e-06 $layer=POLY_cond $X=1.905 $Y=0.615
+ $X2=1.905 $Y2=1.78
r47 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.65 $Y=2.035
+ $X2=1.815 $Y2=2.035
r48 5 6 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.65 $Y=2.035
+ $X2=1.435 $Y2=2.035
r49 1 6 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.345 $Y=2.11
+ $X2=1.435 $Y2=2.035
r50 1 3 206.016 $w=1.8e-07 $l=5.3e-07 $layer=POLY_cond $X=1.345 $Y=2.11
+ $X2=1.345 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTN_1%SCD 1 3 5 8 12 14 15 19
c48 5 0 1.38402e-19 $X=2.875 $Y=2.095
r49 19 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.965 $Y=1.69
+ $X2=2.965 $Y2=1.855
r50 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.965 $Y=1.69
+ $X2=2.965 $Y2=1.525
r51 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.965
+ $Y=1.69 $X2=2.965 $Y2=1.69
r52 15 20 9.14007 $w=4.33e-07 $l=3.45e-07 $layer=LI1_cond $X=3.017 $Y=2.035
+ $X2=3.017 $Y2=1.69
r53 14 20 0.662324 $w=4.33e-07 $l=2.5e-08 $layer=LI1_cond $X=3.017 $Y=1.665
+ $X2=3.017 $Y2=1.69
r54 8 21 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=3.005 $Y=0.615
+ $X2=3.005 $Y2=1.525
r55 5 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.875 $Y=2.095
+ $X2=2.875 $Y2=2.17
r56 5 22 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.875 $Y=2.095
+ $X2=2.875 $Y2=1.855
r57 1 12 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.67 $Y=2.17
+ $X2=2.875 $Y2=2.17
r58 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.67 $Y=2.245
+ $X2=2.67 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTN_1%CLK_N 1 3 4 6 7 8 9
c45 1 0 1.33645e-19 $X=4.71 $Y=1.66
r46 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.44
+ $Y=1.385 $X2=4.44 $Y2=1.385
r47 9 13 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=4.56 $Y=1.38 $X2=4.44
+ $Y2=1.38
r48 7 12 22.2462 $w=4.5e-07 $l=1.8e-07 $layer=POLY_cond $X=4.62 $Y=1.435
+ $X2=4.44 $Y2=1.435
r49 7 8 7.41388 $w=4.5e-07 $l=9e-08 $layer=POLY_cond $X=4.62 $Y=1.435 $X2=4.71
+ $Y2=1.435
r50 4 8 42.5959 $w=1.65e-07 $l=2.32379e-07 $layer=POLY_cond $X=4.725 $Y=1.21
+ $X2=4.71 $Y2=1.435
r51 4 6 151.027 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=4.725 $Y=1.21
+ $X2=4.725 $Y2=0.74
r52 1 8 42.5959 $w=1.65e-07 $l=2.25e-07 $layer=POLY_cond $X=4.71 $Y=1.66
+ $X2=4.71 $Y2=1.435
r53 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.71 $Y=1.66 $X2=4.71
+ $Y2=2.235
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTN_1%A_1069_74# 1 2 9 13 15 19 21 25 27 31 34 35
+ 38 39 41 44 45 46 48 49 50 52 53 55 59 60 62 63 67
c184 63 0 1.94919e-19 $X=6.415 $Y=0.36
c185 59 0 1.33645e-19 $X=5.525 $Y=1.915
c186 53 0 6.18583e-20 $X=9.24 $Y=1.115
c187 52 0 1.42542e-19 $X=9.155 $Y=1.03
c188 35 0 8.56593e-20 $X=5.735 $Y=0.36
c189 25 0 1.98659e-19 $X=10.29 $Y=0.58
c190 15 0 1.33753e-19 $X=6.815 $Y=2.495
c191 13 0 4.67055e-20 $X=6.815 $Y=2.055
r192 60 62 28.4849 $w=2.63e-07 $l=6.55e-07 $layer=LI1_cond $X=5.602 $Y=1.745
+ $X2=5.602 $Y2=1.09
r193 59 60 6.23097 $w=3.73e-07 $l=1.7e-07 $layer=LI1_cond $X=5.547 $Y=1.915
+ $X2=5.547 $Y2=1.745
r194 56 70 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.66 $Y=1.115
+ $X2=9.66 $Y2=1.28
r195 56 67 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=9.66 $Y=1.115
+ $X2=9.66 $Y2=1.005
r196 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.66
+ $Y=1.115 $X2=9.66 $Y2=1.115
r197 53 55 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=9.24 $Y=1.115
+ $X2=9.66 $Y2=1.115
r198 52 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.155 $Y=1.03
+ $X2=9.24 $Y2=1.115
r199 51 52 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=9.155 $Y=0.53
+ $X2=9.155 $Y2=1.03
r200 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.07 $Y=0.445
+ $X2=9.155 $Y2=0.53
r201 49 50 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=9.07 $Y=0.445
+ $X2=8.56 $Y2=0.445
r202 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.475 $Y=0.53
+ $X2=8.56 $Y2=0.445
r203 47 48 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=8.475 $Y=0.53
+ $X2=8.475 $Y2=0.79
r204 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.39 $Y=0.875
+ $X2=8.475 $Y2=0.79
r205 45 46 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=8.39 $Y=0.875
+ $X2=7.26 $Y2=0.875
r206 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.175 $Y=0.79
+ $X2=7.26 $Y2=0.875
r207 43 44 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.175 $Y=0.465
+ $X2=7.175 $Y2=0.79
r208 42 63 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.5 $Y=0.36 $X2=6.415
+ $Y2=0.36
r209 41 43 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=7.09 $Y=0.36
+ $X2=7.175 $Y2=0.465
r210 41 42 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=7.09 $Y=0.36
+ $X2=6.5 $Y2=0.36
r211 39 66 70.8282 $w=2.62e-07 $l=3.85e-07 $layer=POLY_cond $X=6.415 $Y=1.43
+ $X2=6.8 $Y2=1.43
r212 39 64 22.9962 $w=2.62e-07 $l=1.25e-07 $layer=POLY_cond $X=6.415 $Y=1.43
+ $X2=6.29 $Y2=1.43
r213 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.415
+ $Y=1.43 $X2=6.415 $Y2=1.43
r214 36 63 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.415 $Y=0.465
+ $X2=6.415 $Y2=0.36
r215 36 38 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=6.415 $Y=0.465
+ $X2=6.415 $Y2=1.43
r216 34 63 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.33 $Y=0.36
+ $X2=6.415 $Y2=0.36
r217 34 35 31.4242 $w=2.08e-07 $l=5.95e-07 $layer=LI1_cond $X=6.33 $Y=0.36
+ $X2=5.735 $Y2=0.36
r218 29 62 5.88737 $w=2.93e-07 $l=1.47e-07 $layer=LI1_cond $X=5.587 $Y=0.943
+ $X2=5.587 $Y2=1.09
r219 29 31 14.9622 $w=2.93e-07 $l=3.83e-07 $layer=LI1_cond $X=5.587 $Y=0.943
+ $X2=5.587 $Y2=0.56
r220 28 35 7.07071 $w=2.1e-07 $l=1.93505e-07 $layer=LI1_cond $X=5.587 $Y=0.465
+ $X2=5.735 $Y2=0.36
r221 28 31 3.71126 $w=2.93e-07 $l=9.5e-08 $layer=LI1_cond $X=5.587 $Y=0.465
+ $X2=5.587 $Y2=0.56
r222 23 25 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=10.29 $Y=0.93
+ $X2=10.29 $Y2=0.58
r223 22 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.825 $Y=1.005
+ $X2=9.66 $Y2=1.005
r224 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.215 $Y=1.005
+ $X2=10.29 $Y2=0.93
r225 21 22 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=10.215 $Y=1.005
+ $X2=9.825 $Y2=1.005
r226 19 70 458.677 $w=1.8e-07 $l=1.18e-06 $layer=POLY_cond $X=9.62 $Y=2.46
+ $X2=9.62 $Y2=1.28
r227 13 27 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.815 $Y=2.055
+ $X2=6.815 $Y2=1.965
r228 13 15 171.032 $w=1.8e-07 $l=4.4e-07 $layer=POLY_cond $X=6.815 $Y=2.055
+ $X2=6.815 $Y2=2.495
r229 11 66 15.8058 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.8 $Y=1.595
+ $X2=6.8 $Y2=1.43
r230 11 27 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.8 $Y=1.595
+ $X2=6.8 $Y2=1.965
r231 7 64 15.8058 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.29 $Y=1.265
+ $X2=6.29 $Y2=1.43
r232 7 9 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=6.29 $Y=1.265 $X2=6.29
+ $Y2=0.865
r233 2 59 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=5.385
+ $Y=1.735 $X2=5.525 $Y2=1.915
r234 1 31 91 $w=1.7e-07 $l=2.65141e-07 $layer=licon1_NDIFF $count=2 $X=5.345
+ $Y=0.37 $X2=5.525 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTN_1%A_1417_294# 1 2 9 13 17 18 21 27 30 31 32
+ 35 37 38
c97 13 0 1.82775e-19 $X=7.34 $Y=0.865
r98 37 39 0.577631 $w=7.63e-07 $l=3e-08 $layer=LI1_cond $X=9.112 $Y=2.135
+ $X2=9.112 $Y2=2.165
r99 37 38 11.2171 $w=7.63e-07 $l=1.65e-07 $layer=LI1_cond $X=9.112 $Y=2.135
+ $X2=9.112 $Y2=1.97
r100 31 42 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.25 $Y=1.635
+ $X2=7.25 $Y2=1.8
r101 31 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.25 $Y=1.635
+ $X2=7.25 $Y2=1.47
r102 30 32 8.13106 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=7.245 $Y=1.635
+ $X2=7.245 $Y2=1.47
r103 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.25
+ $Y=1.635 $X2=7.25 $Y2=1.635
r104 27 39 11.1064 $w=6.98e-07 $l=6.5e-07 $layer=LI1_cond $X=9.145 $Y=2.815
+ $X2=9.145 $Y2=2.165
r105 23 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.815 $Y=1.3
+ $X2=8.815 $Y2=1.215
r106 23 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.815 $Y=1.3
+ $X2=8.815 $Y2=1.97
r107 19 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.815 $Y=1.13
+ $X2=8.815 $Y2=1.215
r108 19 21 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.815 $Y=1.13
+ $X2=8.815 $Y2=0.865
r109 17 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.73 $Y=1.215
+ $X2=8.815 $Y2=1.215
r110 17 18 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=8.73 $Y=1.215
+ $X2=7.415 $Y2=1.215
r111 15 18 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=7.325 $Y=1.3
+ $X2=7.415 $Y2=1.215
r112 15 32 10.4747 $w=1.78e-07 $l=1.7e-07 $layer=LI1_cond $X=7.325 $Y=1.3
+ $X2=7.325 $Y2=1.47
r113 13 41 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=7.34 $Y=0.865
+ $X2=7.34 $Y2=1.47
r114 9 42 270.153 $w=1.8e-07 $l=6.95e-07 $layer=POLY_cond $X=7.235 $Y=2.495
+ $X2=7.235 $Y2=1.8
r115 2 37 200 $w=1.7e-07 $l=2.5807e-07 $layer=licon1_PDIFF $count=3 $X=8.775
+ $Y=1.96 $X2=8.96 $Y2=2.135
r116 2 27 200 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=3 $X=8.775
+ $Y=1.96 $X2=8.96 $Y2=2.815
r117 1 35 182 $w=1.7e-07 $l=6.61872e-07 $layer=licon1_NDIFF $count=1 $X=8.425
+ $Y=0.72 $X2=8.815 $Y2=1.215
r118 1 21 182 $w=1.7e-07 $l=4.56782e-07 $layer=licon1_NDIFF $count=1 $X=8.425
+ $Y=0.72 $X2=8.815 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTN_1%RESET_B 4 7 10 11 12 15 20 23 29 30 31 32
+ 33 34 35 40 43 46 47 50 51 55 56
c221 55 0 1.97052e-19 $X=11.16 $Y=1.375
c222 47 0 1.38402e-19 $X=3.57 $Y=1.52
c223 35 0 6.65468e-20 $X=8.065 $Y=1.665
c224 31 0 9.59361e-20 $X=11.292 $Y=2.435
r225 55 58 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.16 $Y=1.375
+ $X2=11.16 $Y2=1.54
r226 55 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.16 $Y=1.375
+ $X2=11.16 $Y2=1.21
r227 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.16
+ $Y=1.375 $X2=11.16 $Y2=1.375
r228 50 53 39.7991 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=7.82 $Y=1.635
+ $X2=7.82 $Y2=1.8
r229 50 52 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=7.82 $Y=1.635
+ $X2=7.82 $Y2=1.47
r230 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.82
+ $Y=1.635 $X2=7.82 $Y2=1.635
r231 46 48 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=3.552 $Y=1.52
+ $X2=3.552 $Y2=1.355
r232 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.57
+ $Y=1.52 $X2=3.57 $Y2=1.52
r233 43 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=1.665
+ $X2=3.6 $Y2=1.665
r234 41 56 11.2317 $w=3.15e-07 $l=2.9e-07 $layer=LI1_cond $X=11.195 $Y=1.665
+ $X2=11.195 $Y2=1.375
r235 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=1.665
+ $X2=11.28 $Y2=1.665
r236 37 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=1.665
+ $X2=7.92 $Y2=1.665
r237 35 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.065 $Y=1.665
+ $X2=7.92 $Y2=1.665
r238 34 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.135 $Y=1.665
+ $X2=11.28 $Y2=1.665
r239 34 35 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=11.135 $Y=1.665
+ $X2=8.065 $Y2=1.665
r240 33 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.745 $Y=1.665
+ $X2=3.6 $Y2=1.665
r241 32 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=1.665
+ $X2=7.92 $Y2=1.665
r242 32 33 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=7.775 $Y=1.665
+ $X2=3.745 $Y2=1.665
r243 30 31 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=11.292 $Y=2.285
+ $X2=11.292 $Y2=2.435
r244 30 58 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=11.25 $Y=2.285
+ $X2=11.25 $Y2=1.54
r245 29 31 84.35 $w=1.8e-07 $l=3.15e-07 $layer=POLY_cond $X=11.32 $Y=2.75
+ $X2=11.32 $Y2=2.435
r246 23 57 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=11.25 $Y=0.58
+ $X2=11.25 $Y2=1.21
r247 20 53 270.153 $w=1.8e-07 $l=6.95e-07 $layer=POLY_cond $X=7.715 $Y=2.495
+ $X2=7.715 $Y2=1.8
r248 18 20 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=7.715 $Y=3.075
+ $X2=7.715 $Y2=2.495
r249 15 52 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=7.7 $Y=0.865
+ $X2=7.7 $Y2=1.47
r250 11 18 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=7.625 $Y=3.15
+ $X2=7.715 $Y2=3.075
r251 11 12 2176.69 $w=1.5e-07 $l=4.245e-06 $layer=POLY_cond $X=7.625 $Y=3.15
+ $X2=3.38 $Y2=3.15
r252 9 46 2.68759 $w=3.65e-07 $l=1.7e-08 $layer=POLY_cond $X=3.552 $Y=1.537
+ $X2=3.552 $Y2=1.52
r253 9 10 48.3767 $w=3.65e-07 $l=3.06e-07 $layer=POLY_cond $X=3.552 $Y=1.537
+ $X2=3.552 $Y2=1.843
r254 7 48 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.445 $Y=0.615
+ $X2=3.445 $Y2=1.355
r255 2 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.29 $Y=3.075
+ $X2=3.38 $Y2=3.15
r256 2 4 169.089 $w=1.8e-07 $l=4.35e-07 $layer=POLY_cond $X=3.29 $Y=3.075
+ $X2=3.29 $Y2=2.64
r257 1 10 62.5045 $w=3.1e-07 $l=5.16651e-07 $layer=POLY_cond $X=3.29 $Y=2.245
+ $X2=3.552 $Y2=1.843
r258 1 4 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.29 $Y=2.245
+ $X2=3.29 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTN_1%A_1273_131# 1 2 3 10 12 15 17 21 22 23 24
+ 26 30 36 42
c105 30 0 8.58467e-20 $X=8.39 $Y=1.635
c106 22 0 6.65468e-20 $X=7.785 $Y=2.08
c107 21 0 4.67055e-20 $X=6.76 $Y=1.97
c108 17 0 1.82775e-19 $X=6.795 $Y=0.95
c109 10 0 2.044e-19 $X=8.35 $Y=1.47
r110 31 42 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=8.39 $Y=1.635
+ $X2=8.685 $Y2=1.635
r111 31 39 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=8.39 $Y=1.635
+ $X2=8.35 $Y2=1.635
r112 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.39
+ $Y=1.635 $X2=8.39 $Y2=1.635
r113 28 30 14.5686 $w=2.63e-07 $l=3.35e-07 $layer=LI1_cond $X=8.357 $Y=1.97
+ $X2=8.357 $Y2=1.635
r114 24 28 25.2804 $w=1.94e-07 $l=4.02e-07 $layer=LI1_cond $X=7.955 $Y=2.08
+ $X2=8.357 $Y2=2.08
r115 24 26 11.355 $w=3.38e-07 $l=3.35e-07 $layer=LI1_cond $X=7.955 $Y=2.19
+ $X2=7.955 $Y2=2.525
r116 23 35 16.5015 $w=3.29e-07 $l=5.43171e-07 $layer=LI1_cond $X=6.85 $Y=2.08
+ $X2=6.632 $Y2=2.525
r117 22 24 9.62821 $w=2.2e-07 $l=1.7e-07 $layer=LI1_cond $X=7.785 $Y=2.08
+ $X2=7.955 $Y2=2.08
r118 22 23 48.9788 $w=2.18e-07 $l=9.35e-07 $layer=LI1_cond $X=7.785 $Y=2.08
+ $X2=6.85 $Y2=2.08
r119 21 23 6.56333 $w=3.29e-07 $l=1.48324e-07 $layer=LI1_cond $X=6.76 $Y=1.97
+ $X2=6.85 $Y2=2.08
r120 21 36 55.1465 $w=1.78e-07 $l=8.95e-07 $layer=LI1_cond $X=6.76 $Y=1.97
+ $X2=6.76 $Y2=1.075
r121 17 36 6.68437 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.795 $Y=0.95
+ $X2=6.795 $Y2=1.075
r122 17 19 0.976 $w=2.5e-07 $l=2e-08 $layer=LI1_cond $X=6.795 $Y=0.95 $X2=6.795
+ $Y2=0.93
r123 13 42 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.685 $Y=1.8
+ $X2=8.685 $Y2=1.635
r124 13 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=8.685 $Y=1.8
+ $X2=8.685 $Y2=2.46
r125 10 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.35 $Y=1.47
+ $X2=8.35 $Y2=1.635
r126 10 12 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.35 $Y=1.47
+ $X2=8.35 $Y2=1.04
r127 3 26 600 $w=1.7e-07 $l=3e-07 $layer=licon1_PDIFF $count=1 $X=7.805 $Y=2.285
+ $X2=7.94 $Y2=2.525
r128 2 35 600 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_PDIFF $count=1 $X=6.445
+ $Y=2.285 $X2=6.585 $Y2=2.525
r129 1 19 182 $w=1.7e-07 $l=5.09264e-07 $layer=licon1_NDIFF $count=1 $X=6.365
+ $Y=0.655 $X2=6.755 $Y2=0.93
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTN_1%A_859_347# 1 2 7 9 10 12 14 16 17 18 19 20
+ 21 23 26 28 33 36 38 39 45 47 48 52 56 58 60 64 67 68 69 75
c202 18 0 8.56593e-20 $X=5.875 $Y=0.18
r203 74 75 62.4128 $w=4.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.295 $Y=1.435
+ $X2=5.8 $Y2=1.435
r204 73 74 3.08974 $w=4.5e-07 $l=2.5e-08 $layer=POLY_cond $X=5.27 $Y=1.435
+ $X2=5.295 $Y2=1.435
r205 68 81 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=10.23 $Y=1.455
+ $X2=10.135 $Y2=1.455
r206 67 69 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=10.23 $Y=1.415
+ $X2=10.065 $Y2=1.415
r207 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.23
+ $Y=1.455 $X2=10.23 $Y2=1.455
r208 64 77 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=9.155 $Y=1.635
+ $X2=9.06 $Y2=1.635
r209 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.155
+ $Y=1.635 $X2=9.155 $Y2=1.635
r210 60 63 7.40856 $w=2.78e-07 $l=1.8e-07 $layer=LI1_cond $X=9.21 $Y=1.455
+ $X2=9.21 $Y2=1.635
r211 57 73 6.79744 $w=4.5e-07 $l=5.5e-08 $layer=POLY_cond $X=5.215 $Y=1.435
+ $X2=5.27 $Y2=1.435
r212 56 59 6.36939 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.12 $Y=1.41
+ $X2=5.12 $Y2=1.575
r213 56 58 6.18336 $w=3.58e-07 $l=1.9e-07 $layer=LI1_cond $X=5.12 $Y=1.41
+ $X2=5.12 $Y2=1.22
r214 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.215
+ $Y=1.41 $X2=5.215 $Y2=1.41
r215 54 60 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=9.35 $Y=1.455
+ $X2=9.21 $Y2=1.455
r216 54 69 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=9.35 $Y=1.455
+ $X2=10.065 $Y2=1.455
r217 52 59 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=5.065 $Y=1.82
+ $X2=5.065 $Y2=1.575
r218 49 58 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=5.105 $Y=1.01
+ $X2=5.105 $Y2=1.22
r219 47 49 7.36389 $w=2e-07 $l=2.09105e-07 $layer=LI1_cond $X=4.94 $Y=0.91
+ $X2=5.105 $Y2=1.01
r220 47 48 15.5273 $w=1.98e-07 $l=2.8e-07 $layer=LI1_cond $X=4.94 $Y=0.91
+ $X2=4.66 $Y2=0.91
r221 43 48 7.39673 $w=2e-07 $l=2.12189e-07 $layer=LI1_cond $X=4.492 $Y=0.81
+ $X2=4.66 $Y2=0.91
r222 43 45 8.60032 $w=3.33e-07 $l=2.5e-07 $layer=LI1_cond $X=4.492 $Y=0.81
+ $X2=4.492 $Y2=0.56
r223 39 52 6.98266 $w=1.9e-07 $l=1.65831e-07 $layer=LI1_cond $X=4.94 $Y=1.915
+ $X2=5.065 $Y2=1.82
r224 39 41 27.1435 $w=1.88e-07 $l=4.65e-07 $layer=LI1_cond $X=4.94 $Y=1.915
+ $X2=4.475 $Y2=1.915
r225 34 81 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.135 $Y=1.62
+ $X2=10.135 $Y2=1.455
r226 34 36 439.242 $w=1.8e-07 $l=1.13e-06 $layer=POLY_cond $X=10.135 $Y=1.62
+ $X2=10.135 $Y2=2.75
r227 31 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.06 $Y=1.47
+ $X2=9.06 $Y2=1.635
r228 31 33 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.06 $Y=1.47
+ $X2=9.06 $Y2=1.04
r229 30 33 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=9.06 $Y=0.255
+ $X2=9.06 $Y2=1.04
r230 29 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.045 $Y=0.18
+ $X2=6.97 $Y2=0.18
r231 28 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.985 $Y=0.18
+ $X2=9.06 $Y2=0.255
r232 28 29 994.766 $w=1.5e-07 $l=1.94e-06 $layer=POLY_cond $X=8.985 $Y=0.18
+ $X2=7.045 $Y2=0.18
r233 24 38 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.97 $Y=0.255
+ $X2=6.97 $Y2=0.18
r234 24 26 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.97 $Y=0.255
+ $X2=6.97 $Y2=0.865
r235 21 23 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.355 $Y=2.21
+ $X2=6.355 $Y2=2.495
r236 19 21 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.265 $Y=2.135
+ $X2=6.355 $Y2=2.21
r237 19 20 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=6.265 $Y=2.135
+ $X2=5.875 $Y2=2.135
r238 17 38 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.895 $Y=0.18
+ $X2=6.97 $Y2=0.18
r239 17 18 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=6.895 $Y=0.18
+ $X2=5.875 $Y2=0.18
r240 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.8 $Y=2.06
+ $X2=5.875 $Y2=2.135
r241 15 75 28.7666 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=5.8 $Y=1.66
+ $X2=5.8 $Y2=1.435
r242 15 16 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=5.8 $Y=1.66 $X2=5.8
+ $Y2=2.06
r243 14 75 28.7666 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=5.8 $Y=1.21
+ $X2=5.8 $Y2=1.435
r244 13 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.8 $Y=0.255
+ $X2=5.875 $Y2=0.18
r245 13 14 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=5.8 $Y=0.255
+ $X2=5.8 $Y2=1.21
r246 10 74 24.2915 $w=1.8e-07 $l=2.25e-07 $layer=POLY_cond $X=5.295 $Y=1.66
+ $X2=5.295 $Y2=1.435
r247 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.295 $Y=1.66
+ $X2=5.295 $Y2=2.235
r248 7 73 28.7666 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=5.27 $Y=1.21
+ $X2=5.27 $Y2=1.435
r249 7 9 151.027 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=5.27 $Y=1.21 $X2=5.27
+ $Y2=0.74
r250 2 41 600 $w=1.7e-07 $l=2.54558e-07 $layer=licon1_PDIFF $count=1 $X=4.295
+ $Y=1.735 $X2=4.475 $Y2=1.915
r251 1 45 91 $w=1.7e-07 $l=2.61534e-07 $layer=licon1_NDIFF $count=2 $X=4.32
+ $Y=0.37 $X2=4.49 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTN_1%A_2087_410# 1 2 9 13 15 19 21 25 28 30 31
+ 35
c91 30 0 9.59361e-20 $X=10.6 $Y=2.215
r92 31 38 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.6 $Y=2.215
+ $X2=10.6 $Y2=2.38
r93 31 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.6 $Y=2.215
+ $X2=10.6 $Y2=2.05
r94 30 33 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=10.56 $Y=2.215
+ $X2=10.56 $Y2=2.375
r95 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.6
+ $Y=2.215 $X2=10.6 $Y2=2.215
r96 27 28 103.733 $w=1.68e-07 $l=1.59e-06 $layer=LI1_cond $X=12.15 $Y=0.7
+ $X2=12.15 $Y2=2.29
r97 26 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.71 $Y=2.375
+ $X2=11.545 $Y2=2.375
r98 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.065 $Y=2.375
+ $X2=12.15 $Y2=2.29
r99 25 26 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=12.065 $Y=2.375
+ $X2=11.71 $Y2=2.375
r100 21 27 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=12.065 $Y=0.575
+ $X2=12.15 $Y2=0.7
r101 21 23 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=12.065 $Y=0.575
+ $X2=11.96 $Y2=0.575
r102 17 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.545 $Y=2.46
+ $X2=11.545 $Y2=2.375
r103 17 19 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=11.545 $Y=2.46
+ $X2=11.545 $Y2=2.75
r104 16 33 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.685 $Y=2.375
+ $X2=10.56 $Y2=2.375
r105 15 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.38 $Y=2.375
+ $X2=11.545 $Y2=2.375
r106 15 16 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=11.38 $Y=2.375
+ $X2=10.685 $Y2=2.375
r107 13 37 753.766 $w=1.5e-07 $l=1.47e-06 $layer=POLY_cond $X=10.69 $Y=0.58
+ $X2=10.69 $Y2=2.05
r108 9 38 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=10.545 $Y=2.75
+ $X2=10.545 $Y2=2.38
r109 2 19 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=11.41
+ $Y=2.54 $X2=11.545 $Y2=2.75
r110 1 23 182 $w=1.7e-07 $l=3.46482e-07 $layer=licon1_NDIFF $count=1 $X=11.715
+ $Y=0.37 $X2=11.96 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTN_1%A_1827_144# 1 2 7 9 11 13 16 18 20 22 24 25
+ 27 28 29 30 38 42 43 44 46 51 52 57
c145 57 0 1.97052e-19 $X=10.94 $Y=1.795
c146 44 0 1.98659e-19 $X=11.565 $Y=0.955
c147 20 0 1.07922e-19 $X=12.77 $Y=1.07
c148 18 0 1.07922e-19 $X=12.74 $Y=1.97
r149 57 59 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=10.94 $Y=1.795
+ $X2=10.94 $Y2=2.035
r150 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.73
+ $Y=1.065 $X2=11.73 $Y2=1.065
r151 49 51 30.9064 $w=3.28e-07 $l=8.85e-07 $layer=LI1_cond $X=11.73 $Y=1.95
+ $X2=11.73 $Y2=1.065
r152 48 51 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=11.73 $Y=1.04
+ $X2=11.73 $Y2=1.065
r153 47 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.025 $Y=2.035
+ $X2=10.94 $Y2=2.035
r154 46 49 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.565 $Y=2.035
+ $X2=11.73 $Y2=1.95
r155 46 47 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=11.565 $Y=2.035
+ $X2=11.025 $Y2=2.035
r156 45 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.475 $Y=0.955
+ $X2=10.39 $Y2=0.955
r157 44 48 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.565 $Y=0.955
+ $X2=11.73 $Y2=1.04
r158 44 45 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=11.565 $Y=0.955
+ $X2=10.475 $Y2=0.955
r159 42 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.855 $Y=1.795
+ $X2=10.94 $Y2=1.795
r160 42 43 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=10.855 $Y=1.795
+ $X2=10.065 $Y2=1.795
r161 38 40 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=9.9 $Y=2.135
+ $X2=9.9 $Y2=2.815
r162 36 43 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.9 $Y=1.88
+ $X2=10.065 $Y2=1.795
r163 36 38 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=9.9 $Y=1.88
+ $X2=9.9 $Y2=2.135
r164 32 35 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=9.495 $Y=0.695
+ $X2=10.075 $Y2=0.695
r165 30 55 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=10.39 $Y=0.695
+ $X2=10.39 $Y2=0.955
r166 30 35 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=10.305 $Y=0.695
+ $X2=10.075 $Y2=0.695
r167 25 27 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=12.845 $Y=0.995
+ $X2=12.845 $Y2=0.645
r168 22 24 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=12.83 $Y=2.045
+ $X2=12.83 $Y2=2.54
r169 21 52 12.1617 $w=1.5e-07 $l=1.8747e-07 $layer=POLY_cond $X=11.895 $Y=1.07
+ $X2=11.73 $Y2=1.022
r170 20 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.77 $Y=1.07
+ $X2=12.845 $Y2=0.995
r171 20 21 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=12.77 $Y=1.07
+ $X2=11.895 $Y2=1.07
r172 19 29 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=11.86 $Y=1.97
+ $X2=11.77 $Y2=1.97
r173 18 22 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=12.74 $Y=1.97
+ $X2=12.83 $Y2=2.045
r174 18 19 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=12.74 $Y=1.97
+ $X2=11.86 $Y2=1.97
r175 14 29 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=11.77 $Y=2.045
+ $X2=11.77 $Y2=1.97
r176 14 16 274.04 $w=1.8e-07 $l=7.05e-07 $layer=POLY_cond $X=11.77 $Y=2.045
+ $X2=11.77 $Y2=2.75
r177 13 29 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=11.755
+ $Y=1.895 $X2=11.77 $Y2=1.97
r178 13 28 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=11.755 $Y=1.895
+ $X2=11.755 $Y2=1.57
r179 11 28 38.9318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.73 $Y=1.405
+ $X2=11.73 $Y2=1.57
r180 10 52 13.5877 $w=2.4e-07 $l=1.23e-07 $layer=POLY_cond $X=11.73 $Y=1.145
+ $X2=11.73 $Y2=1.022
r181 10 11 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=11.73 $Y=1.145
+ $X2=11.73 $Y2=1.405
r182 7 52 13.5877 $w=2.4e-07 $l=1.60823e-07 $layer=POLY_cond $X=11.64 $Y=0.9
+ $X2=11.73 $Y2=1.022
r183 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.64 $Y=0.9
+ $X2=11.64 $Y2=0.58
r184 2 40 600 $w=1.7e-07 $l=9.45238e-07 $layer=licon1_PDIFF $count=1 $X=9.71
+ $Y=1.96 $X2=9.9 $Y2=2.815
r185 2 38 300 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=2 $X=9.71
+ $Y=1.96 $X2=9.845 $Y2=2.135
r186 1 35 182 $w=1.7e-07 $l=9.9111e-07 $layer=licon1_NDIFF $count=1 $X=9.135
+ $Y=0.72 $X2=10.075 $Y2=0.615
r187 1 32 182 $w=1.7e-07 $l=3.7229e-07 $layer=licon1_NDIFF $count=1 $X=9.135
+ $Y=0.72 $X2=9.495 $Y2=0.695
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTN_1%A_2492_424# 1 2 9 13 15 16 19 23 26
c44 26 0 2.15844e-19 $X=12.645 $Y=1.52
r45 26 29 5.13927 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=12.625 $Y=1.52
+ $X2=12.625 $Y2=1.685
r46 26 28 5.13927 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=12.625 $Y=1.52
+ $X2=12.625 $Y2=1.355
r47 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.645
+ $Y=1.52 $X2=12.645 $Y2=1.52
r48 23 29 18.8286 $w=3.53e-07 $l=5.8e-07 $layer=LI1_cond $X=12.617 $Y=2.265
+ $X2=12.617 $Y2=1.685
r49 19 28 23.0489 $w=3.53e-07 $l=7.1e-07 $layer=LI1_cond $X=12.617 $Y=0.645
+ $X2=12.617 $Y2=1.355
r50 15 27 118.031 $w=3.3e-07 $l=6.75e-07 $layer=POLY_cond $X=13.32 $Y=1.52
+ $X2=12.645 $Y2=1.52
r51 15 16 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=13.32 $Y=1.52
+ $X2=13.41 $Y2=1.52
r52 11 16 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=13.425 $Y=1.355
+ $X2=13.41 $Y2=1.52
r53 11 13 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=13.425 $Y=1.355
+ $X2=13.425 $Y2=0.74
r54 7 16 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=13.41 $Y=1.685
+ $X2=13.41 $Y2=1.52
r55 7 9 277.927 $w=1.8e-07 $l=7.15e-07 $layer=POLY_cond $X=13.41 $Y=1.685
+ $X2=13.41 $Y2=2.4
r56 2 23 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=12.46
+ $Y=2.12 $X2=12.605 $Y2=2.265
r57 1 19 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=12.485
+ $Y=0.37 $X2=12.63 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTN_1%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 47 52
+ 53 54 56 61 69 74 82 87 99 105 106 109 112 119 122 125 128 135
c139 5 0 8.58467e-20 $X=8.335 $Y=1.96
r140 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r141 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r142 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r143 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r144 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r145 112 115 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.98 $Y=3.055
+ $X2=2.98 $Y2=3.33
r146 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r147 106 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=13.2 $Y2=3.33
r148 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r149 103 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.305 $Y=3.33
+ $X2=13.14 $Y2=3.33
r150 103 105 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.305 $Y=3.33
+ $X2=13.68 $Y2=3.33
r151 102 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r152 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r153 99 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.975 $Y=3.33
+ $X2=13.14 $Y2=3.33
r154 99 101 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=12.975 $Y=3.33
+ $X2=12.72 $Y2=3.33
r155 98 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.72 $Y2=3.33
r156 98 132 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=10.8 $Y2=3.33
r157 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r158 95 97 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=11.21 $Y=3.33
+ $X2=11.76 $Y2=3.33
r159 94 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r160 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r161 91 94 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r162 91 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r163 90 93 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=10.32 $Y2=3.33
r164 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r165 88 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.625 $Y=3.33
+ $X2=8.46 $Y2=3.33
r166 88 90 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.625 $Y=3.33
+ $X2=8.88 $Y2=3.33
r167 87 95 8.37032 $w=1.7e-07 $l=3.03e-07 $layer=LI1_cond $X=10.907 $Y=3.33
+ $X2=11.21 $Y2=3.33
r168 87 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r169 87 128 10.1815 $w=6.03e-07 $l=5.15e-07 $layer=LI1_cond $X=10.907 $Y=3.33
+ $X2=10.907 $Y2=2.815
r170 87 93 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=10.605 $Y=3.33
+ $X2=10.32 $Y2=3.33
r171 86 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r172 86 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r173 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r174 83 122 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.545 $Y=3.33
+ $X2=7.42 $Y2=3.33
r175 83 85 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.545 $Y=3.33
+ $X2=7.92 $Y2=3.33
r176 82 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.295 $Y=3.33
+ $X2=8.46 $Y2=3.33
r177 82 85 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.295 $Y=3.33
+ $X2=7.92 $Y2=3.33
r178 78 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r179 77 80 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=6.96 $Y2=3.33
r180 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r181 75 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.17 $Y=3.33
+ $X2=5.005 $Y2=3.33
r182 75 77 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=5.17 $Y=3.33
+ $X2=5.52 $Y2=3.33
r183 74 122 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.295 $Y=3.33
+ $X2=7.42 $Y2=3.33
r184 74 80 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.295 $Y=3.33
+ $X2=6.96 $Y2=3.33
r185 73 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r186 73 116 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=3.12 $Y2=3.33
r187 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r188 70 115 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.145 $Y=3.33
+ $X2=2.98 $Y2=3.33
r189 70 72 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=3.145 $Y=3.33
+ $X2=4.56 $Y2=3.33
r190 69 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.84 $Y=3.33
+ $X2=5.005 $Y2=3.33
r191 69 72 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.84 $Y=3.33
+ $X2=4.56 $Y2=3.33
r192 68 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r193 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r194 65 68 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r195 65 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r196 64 67 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r197 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r198 62 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r199 62 64 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r200 61 115 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=3.33
+ $X2=2.98 $Y2=3.33
r201 61 67 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.815 $Y=3.33
+ $X2=2.64 $Y2=3.33
r202 59 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r203 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r204 56 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r205 56 58 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r206 54 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r207 54 78 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=5.52 $Y2=3.33
r208 54 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r209 52 97 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=11.88 $Y=3.33
+ $X2=11.76 $Y2=3.33
r210 52 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.88 $Y=3.33
+ $X2=12.045 $Y2=3.33
r211 51 101 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=12.21 $Y=3.33
+ $X2=12.72 $Y2=3.33
r212 51 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.21 $Y=3.33
+ $X2=12.045 $Y2=3.33
r213 47 50 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=13.14 $Y=1.985
+ $X2=13.14 $Y2=2.4
r214 45 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.14 $Y=3.245
+ $X2=13.14 $Y2=3.33
r215 45 50 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=13.14 $Y=3.245
+ $X2=13.14 $Y2=2.4
r216 41 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.045 $Y=3.245
+ $X2=12.045 $Y2=3.33
r217 41 43 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=12.045 $Y=3.245
+ $X2=12.045 $Y2=2.805
r218 37 125 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.46 $Y=3.245
+ $X2=8.46 $Y2=3.33
r219 37 39 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=8.46 $Y=3.245
+ $X2=8.46 $Y2=2.395
r220 33 122 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.42 $Y=3.245
+ $X2=7.42 $Y2=3.33
r221 33 35 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=7.42 $Y=3.245
+ $X2=7.42 $Y2=2.525
r222 29 119 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.005 $Y=3.245
+ $X2=5.005 $Y2=3.33
r223 29 31 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=5.005 $Y=3.245
+ $X2=5.005 $Y2=2.635
r224 25 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r225 25 27 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.805
r226 8 50 300 $w=1.7e-07 $l=3.74166e-07 $layer=licon1_PDIFF $count=2 $X=12.92
+ $Y=2.12 $X2=13.14 $Y2=2.4
r227 8 47 600 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_PDIFF $count=1 $X=12.92
+ $Y=2.12 $X2=13.14 $Y2=1.985
r228 7 43 600 $w=1.7e-07 $l=3.45326e-07 $layer=licon1_PDIFF $count=1 $X=11.86
+ $Y=2.54 $X2=12.045 $Y2=2.805
r229 6 128 600 $w=1.7e-07 $l=3.87137e-07 $layer=licon1_PDIFF $count=1 $X=10.635
+ $Y=2.54 $X2=10.905 $Y2=2.815
r230 5 39 300 $w=1.7e-07 $l=4.93559e-07 $layer=licon1_PDIFF $count=2 $X=8.335
+ $Y=1.96 $X2=8.46 $Y2=2.395
r231 4 35 600 $w=1.7e-07 $l=3e-07 $layer=licon1_PDIFF $count=1 $X=7.325 $Y=2.285
+ $X2=7.46 $Y2=2.525
r232 3 31 600 $w=1.7e-07 $l=9.97246e-07 $layer=licon1_PDIFF $count=1 $X=4.8
+ $Y=1.735 $X2=5.005 $Y2=2.635
r233 2 112 600 $w=1.7e-07 $l=8.3781e-07 $layer=licon1_PDIFF $count=1 $X=2.76
+ $Y=2.32 $X2=2.98 $Y2=3.055
r234 1 27 600 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=2.32 $X2=0.73 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTN_1%A_287_464# 1 2 3 4 5 18 22 25 26 27 29 30
+ 32 36 38 39 42 45 46 53 55
c131 55 0 2.66294e-20 $X=6.072 $Y=2.28
c132 39 0 1.07123e-19 $X=6.072 $Y=2.18
r133 47 49 2.37047 $w=3.86e-07 $l=7.5e-08 $layer=LI1_cond $X=3.752 $Y=2.39
+ $X2=3.752 $Y2=2.465
r134 45 46 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.055 $Y=2.795
+ $X2=2.22 $Y2=2.795
r135 40 55 3.66998 $w=2.97e-07 $l=1.13137e-07 $layer=LI1_cond $X=6.1 $Y=2.38
+ $X2=6.072 $Y2=2.28
r136 40 42 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.1 $Y=2.38
+ $X2=6.1 $Y2=2.525
r137 39 55 3.66998 $w=2.97e-07 $l=1e-07 $layer=LI1_cond $X=6.072 $Y=2.18
+ $X2=6.072 $Y2=2.28
r138 38 54 6.38767 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=6.072 $Y=2.002
+ $X2=6.072 $Y2=1.84
r139 38 39 6.31184 $w=3.23e-07 $l=1.78e-07 $layer=LI1_cond $X=6.072 $Y=2.002
+ $X2=6.072 $Y2=2.18
r140 36 54 44.9453 $w=2.48e-07 $l=9.75e-07 $layer=LI1_cond $X=6.035 $Y=0.865
+ $X2=6.035 $Y2=1.84
r141 32 55 2.80448 $w=2e-07 $l=1.62e-07 $layer=LI1_cond $X=5.91 $Y=2.28
+ $X2=6.072 $Y2=2.28
r142 32 53 77.3591 $w=1.98e-07 $l=1.395e-06 $layer=LI1_cond $X=5.91 $Y=2.28
+ $X2=4.515 $Y2=2.28
r143 31 47 0.194975 $w=4.2e-07 $l=3.23e-07 $layer=LI1_cond $X=4.075 $Y=2.39
+ $X2=3.752 $Y2=2.39
r144 30 53 8.93948 $w=4.18e-07 $l=2.1e-07 $layer=LI1_cond $X=4.305 $Y=2.39
+ $X2=4.515 $Y2=2.39
r145 30 31 6.311 $w=4.18e-07 $l=2.3e-07 $layer=LI1_cond $X=4.305 $Y=2.39
+ $X2=4.075 $Y2=2.39
r146 29 47 10.5186 $w=3.86e-07 $l=3.26533e-07 $layer=LI1_cond $X=3.99 $Y=2.18
+ $X2=3.752 $Y2=2.39
r147 28 29 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=3.99 $Y=1.185
+ $X2=3.99 $Y2=2.18
r148 26 28 6.9898 $w=2.25e-07 $l=1.49579e-07 $layer=LI1_cond $X=3.905 $Y=1.072
+ $X2=3.99 $Y2=1.185
r149 26 27 51.988 $w=2.23e-07 $l=1.015e-06 $layer=LI1_cond $X=3.905 $Y=1.072
+ $X2=2.89 $Y2=1.072
r150 25 27 6.9898 $w=2.25e-07 $l=1.4854e-07 $layer=LI1_cond $X=2.805 $Y=0.96
+ $X2=2.89 $Y2=1.072
r151 24 25 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.805 $Y=0.765
+ $X2=2.805 $Y2=0.96
r152 22 52 3.16062 $w=3.86e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.43 $Y=2.715
+ $X2=3.515 $Y2=2.815
r153 22 49 7.90155 $w=3.86e-07 $l=4.29167e-07 $layer=LI1_cond $X=3.43 $Y=2.715
+ $X2=3.752 $Y2=2.465
r154 22 46 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=3.43 $Y=2.715
+ $X2=2.22 $Y2=2.715
r155 18 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.72 $Y=0.68
+ $X2=2.805 $Y2=0.765
r156 18 20 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.72 $Y=0.68
+ $X2=2.26 $Y2=0.68
r157 5 42 600 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_PDIFF $count=1 $X=5.985
+ $Y=2.285 $X2=6.125 $Y2=2.525
r158 4 52 600 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_PDIFF $count=1 $X=3.38
+ $Y=2.32 $X2=3.515 $Y2=2.815
r159 4 49 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.38
+ $Y=2.32 $X2=3.515 $Y2=2.465
r160 3 45 300 $w=1.7e-07 $l=8.23954e-07 $layer=licon1_PDIFF $count=2 $X=1.435
+ $Y=2.32 $X2=2.055 $Y2=2.795
r161 2 36 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=5.95
+ $Y=0.655 $X2=6.075 $Y2=0.865
r162 1 20 182 $w=1.7e-07 $l=3.94208e-07 $layer=licon1_NDIFF $count=1 $X=1.98
+ $Y=0.405 $X2=2.26 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTN_1%Q 1 2 7 8 9 10 11 12 13
r13 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=13.64 $Y=2.405
+ $X2=13.64 $Y2=2.775
r14 11 12 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=13.64 $Y=1.985
+ $X2=13.64 $Y2=2.405
r15 10 11 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=13.64 $Y=1.665
+ $X2=13.64 $Y2=1.985
r16 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=13.64 $Y=1.295
+ $X2=13.64 $Y2=1.665
r17 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=13.64 $Y=0.925
+ $X2=13.64 $Y2=1.295
r18 7 8 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=13.64 $Y=0.515
+ $X2=13.64 $Y2=0.925
r19 2 13 400 $w=1.7e-07 $l=1.04265e-06 $layer=licon1_PDIFF $count=1 $X=13.5
+ $Y=1.84 $X2=13.64 $Y2=2.815
r20 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.5
+ $Y=1.84 $X2=13.64 $Y2=1.985
r21 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.5
+ $Y=0.37 $X2=13.64 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTN_1%VGND 1 2 3 4 5 6 21 25 29 33 37 41 46 47 48
+ 50 62 66 71 76 86 87 90 93 96 99 102
r125 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r126 99 100 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r127 96 97 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r128 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r129 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r130 87 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r131 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r132 84 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.305 $Y=0
+ $X2=13.14 $Y2=0
r133 84 86 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.305 $Y=0
+ $X2=13.68 $Y2=0
r134 83 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r135 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r136 80 83 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=12.72 $Y2=0
r137 80 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r138 79 82 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=11.28 $Y=0
+ $X2=12.72 $Y2=0
r139 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r140 77 99 10.873 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=11.2 $Y=0 $X2=10.965
+ $Y2=0
r141 77 79 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=11.2 $Y=0 $X2=11.28
+ $Y2=0
r142 76 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.975 $Y=0
+ $X2=13.14 $Y2=0
r143 76 82 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=12.975 $Y=0
+ $X2=12.72 $Y2=0
r144 75 100 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.4 $Y=0 $X2=10.8
+ $Y2=0
r145 75 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r146 74 75 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r147 72 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.22 $Y=0 $X2=8.055
+ $Y2=0
r148 72 74 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.22 $Y=0 $X2=8.4
+ $Y2=0
r149 71 99 10.873 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=10.73 $Y=0
+ $X2=10.965 $Y2=0
r150 71 74 152.011 $w=1.68e-07 $l=2.33e-06 $layer=LI1_cond $X=10.73 $Y=0 $X2=8.4
+ $Y2=0
r151 70 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r152 69 70 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r153 67 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.165 $Y=0 $X2=5
+ $Y2=0
r154 67 69 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.165 $Y=0
+ $X2=5.52 $Y2=0
r155 66 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.89 $Y=0 $X2=8.055
+ $Y2=0
r156 66 69 154.62 $w=1.68e-07 $l=2.37e-06 $layer=LI1_cond $X=7.89 $Y=0 $X2=5.52
+ $Y2=0
r157 65 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r158 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r159 62 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=0 $X2=5
+ $Y2=0
r160 62 64 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.835 $Y=0
+ $X2=4.56 $Y2=0
r161 61 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r162 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r163 58 61 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r164 58 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r165 57 60 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r166 57 58 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r167 55 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r168 55 57 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r169 53 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r170 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r171 50 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r172 50 52 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r173 48 97 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r174 48 70 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=5.52 $Y2=0
r175 46 60 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.655 $Y=0 $X2=3.6
+ $Y2=0
r176 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.655 $Y=0 $X2=3.82
+ $Y2=0
r177 45 64 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=3.985 $Y=0
+ $X2=4.56 $Y2=0
r178 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.985 $Y=0 $X2=3.82
+ $Y2=0
r179 41 43 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=13.14 $Y=0.555
+ $X2=13.14 $Y2=0.965
r180 39 102 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.14 $Y=0.085
+ $X2=13.14 $Y2=0
r181 39 41 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=13.14 $Y=0.085
+ $X2=13.14 $Y2=0.555
r182 35 99 1.91284 $w=4.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.965 $Y=0.085
+ $X2=10.965 $Y2=0
r183 35 37 10.9428 $w=4.68e-07 $l=4.3e-07 $layer=LI1_cond $X=10.965 $Y=0.085
+ $X2=10.965 $Y2=0.515
r184 31 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.055 $Y=0.085
+ $X2=8.055 $Y2=0
r185 31 33 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=8.055 $Y=0.085
+ $X2=8.055 $Y2=0.535
r186 27 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0
r187 27 29 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=5 $Y=0.085 $X2=5
+ $Y2=0.535
r188 23 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.82 $Y=0.085
+ $X2=3.82 $Y2=0
r189 23 25 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=3.82 $Y=0.085
+ $X2=3.82 $Y2=0.615
r190 19 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r191 19 21 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.65
r192 6 43 182 $w=1.7e-07 $l=7.25655e-07 $layer=licon1_NDIFF $count=1 $X=12.92
+ $Y=0.37 $X2=13.21 $Y2=0.965
r193 6 41 182 $w=1.7e-07 $l=2.98496e-07 $layer=licon1_NDIFF $count=1 $X=12.92
+ $Y=0.37 $X2=13.14 $Y2=0.555
r194 5 37 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=10.765
+ $Y=0.37 $X2=10.965 $Y2=0.515
r195 4 33 182 $w=1.7e-07 $l=3.34664e-07 $layer=licon1_NDIFF $count=1 $X=7.775
+ $Y=0.655 $X2=8.055 $Y2=0.535
r196 3 29 182 $w=1.7e-07 $l=2.70185e-07 $layer=licon1_NDIFF $count=1 $X=4.8
+ $Y=0.37 $X2=5 $Y2=0.535
r197 2 25 182 $w=1.7e-07 $l=3.91152e-07 $layer=licon1_NDIFF $count=1 $X=3.52
+ $Y=0.405 $X2=3.82 $Y2=0.615
r198 1 21 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.44 $X2=0.78 $Y2=0.65
.ends

.subckt PM_SKY130_FD_SC_MS__SDFRTN_1%noxref_24 1 2 9 11 12 15
r34 13 15 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.225 $Y=0.425
+ $X2=3.225 $Y2=0.615
r35 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.06 $Y=0.34
+ $X2=3.225 $Y2=0.425
r36 11 12 102.102 $w=1.68e-07 $l=1.565e-06 $layer=LI1_cond $X=3.06 $Y=0.34
+ $X2=1.495 $Y2=0.34
r37 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.33 $Y=0.425
+ $X2=1.495 $Y2=0.34
r38 7 9 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.33 $Y=0.425 $X2=1.33
+ $Y2=0.575
r39 2 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.08
+ $Y=0.405 $X2=3.225 $Y2=0.615
r40 1 9 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1 $X=1.195
+ $Y=0.405 $X2=1.33 $Y2=0.575
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_ms__sdfrtn_1 CLK_N D RESET_B SCD SCE VGND VNB VPB VPWR Q
*.PININFO CLK_N:I D:I RESET_B:I SCD:I SCE:I VGND:I VNB:I VPB:I VPWR:I
*.PININFO Q:O
MI642 clkpos CLK_N VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI636 clkneg clkpos VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI42 db clkneg M0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI656 net87 s0 net121 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI657 net121 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI33 net114 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI634 sceb SCE VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI4 M0 clkpos net102 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI34 net102 M1 net114 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI655 s0 clkneg net97 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI652 net182 s0 VGND VNB nfet_01v8_lvt m=1 w=0.55 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI653 Q net182 VGND VNB nfet_01v8_lvt m=1 w=0.74 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI654 net97 net87 VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI647 M1 M0 VGND VNB nfet_01v8_lvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI649 M1 clkpos s0 VNB nfet_01v8_lvt m=1 w=0.64 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI666 net137 RESET_B VGND VNB nfet_01v8_lvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI98 db D n0 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI103 n1 SCD net137 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI120 db SCE n1 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI104 n0 sceb net137 VNB nfet_01v8_lvt m=1 w=0.42 l=0.15 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.525 perim=3.1
MI643 clkpos CLK_N VPWR VPB pfet_01v8 m=1 w=1 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI635 clkneg clkpos VPWR VPB pfet_01v8 m=1 w=1 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI43 db clkpos M0 VPB pfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI662 net210 net87 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.18 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI659 net87 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.18 mult=1
+ sa=0.265 sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI664 s0 clkpos net210 VPB pfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI658 net87 s0 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI30 net189 M1 VPWR VPB pfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI31 M0 clkneg net189 VPB pfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI32 M0 RESET_B VPWR VPB pfet_01v8 m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI663 net182 s0 VPWR VPB pfet_01v8 m=1 w=0.84 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI660 Q net182 VPWR VPB pfet_01v8 m=1 w=1.12 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI648 M1 M0 VPWR VPB pfet_01v8 m=1 w=1.0 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI650 M1 clkneg s0 VPB pfet_01v8 m=1 w=1.0 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI633 sceb SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI101 db sceb p1 VPB pfet_01v8 m=1 w=0.64 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI107 p0 SCE VPWR VPB pfet_01v8 m=1 w=0.64 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI94 db D p0 VPB pfet_01v8 m=1 w=0.64 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MI108 p1 SCD VPWR VPB pfet_01v8 m=1 w=0.64 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MI665 db RESET_B VPWR VPB pfet_01v8 m=1 w=0.64 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_ms__sdfrtn_1

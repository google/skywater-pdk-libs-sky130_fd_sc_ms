* File: sky130_fd_sc_ms__dlrbn_2.pex.spice
* Created: Fri Aug 28 17:26:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLRBN_2%D 2 5 9 11 12 15
r36 15 17 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.425
+ $X2=0.585 $Y2=1.26
r37 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.425 $X2=0.59 $Y2=1.425
r38 12 16 2.32075 $w=6.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.72 $Y=1.595
+ $X2=0.59 $Y2=1.595
r39 9 17 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=0.495 $Y=0.835
+ $X2=0.495 $Y2=1.26
r40 5 11 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=0.505 $Y=2.54
+ $X2=0.505 $Y2=1.93
r41 2 11 41.5618 $w=3.4e-07 $l=1.7e-07 $layer=POLY_cond $X=0.585 $Y=1.76
+ $X2=0.585 $Y2=1.93
r42 1 15 0.848592 $w=3.4e-07 $l=5e-09 $layer=POLY_cond $X=0.585 $Y=1.43
+ $X2=0.585 $Y2=1.425
r43 1 2 56.007 $w=3.4e-07 $l=3.3e-07 $layer=POLY_cond $X=0.585 $Y=1.43 $X2=0.585
+ $Y2=1.76
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_2%GATE_N 3 7 11 12 13 16 17
r39 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.13
+ $Y=1.425 $X2=1.13 $Y2=1.425
r40 13 17 8.92214 $w=3.08e-07 $l=2.4e-07 $layer=LI1_cond $X=1.13 $Y=1.665
+ $X2=1.13 $Y2=1.425
r41 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.13 $Y=1.765
+ $X2=1.13 $Y2=1.425
r42 11 12 38.198 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.765
+ $X2=1.13 $Y2=1.93
r43 10 16 41.3509 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.26
+ $X2=1.13 $Y2=1.425
r44 7 12 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=1.185 $Y=2.54
+ $X2=1.185 $Y2=1.93
r45 3 10 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.075 $Y=0.74
+ $X2=1.075 $Y2=1.26
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_2%A_230_74# 1 2 9 12 16 19 22 23 26 27 30 32
+ 33 34 37 38 41 48 49 53 57 63 66 69
c148 63 0 4.17599e-20 $X=3.365 $Y=1.285
c149 53 0 9.56297e-20 $X=2.285 $Y=1.385
c150 37 0 1.2913e-19 $X=4 $Y=2.215
c151 27 0 1.15905e-19 $X=3.155 $Y=1.215
r152 63 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.365 $Y=1.285
+ $X2=3.365 $Y2=1.12
r153 62 64 8.55446 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=3.342 $Y=1.285
+ $X2=3.342 $Y2=1.45
r154 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.365
+ $Y=1.285 $X2=3.365 $Y2=1.285
r155 55 57 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.095 $Y=2.055
+ $X2=3.24 $Y2=2.055
r156 53 67 40.7727 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=1.385
+ $X2=2.275 $Y2=1.55
r157 53 66 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=1.385
+ $X2=2.275 $Y2=1.22
r158 52 54 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=1.385
+ $X2=2.305 $Y2=1.55
r159 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.285
+ $Y=1.385 $X2=2.285 $Y2=1.385
r160 49 52 5.76222 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=2.305 $Y=1.215
+ $X2=2.305 $Y2=1.385
r161 47 48 6.145 $w=3.78e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=2.29
+ $X2=1.625 $Y2=2.29
r162 45 47 3.94257 $w=3.78e-07 $l=1.3e-07 $layer=LI1_cond $X=1.41 $Y=2.29
+ $X2=1.54 $Y2=2.29
r163 41 43 19.325 $w=4.98e-07 $l=5.75e-07 $layer=LI1_cond $X=1.375 $Y=0.515
+ $X2=1.375 $Y2=1.09
r164 38 71 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=4 $Y=2.215 $X2=3.84
+ $Y2=2.215
r165 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4
+ $Y=2.215 $X2=4 $Y2=2.215
r166 35 37 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=4 $Y=2.905 $X2=4
+ $Y2=2.215
r167 33 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.835 $Y=2.99
+ $X2=4 $Y2=2.905
r168 33 34 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.835 $Y=2.99
+ $X2=3.18 $Y2=2.99
r169 32 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.24 $Y=1.97
+ $X2=3.24 $Y2=2.055
r170 32 64 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.24 $Y=1.97
+ $X2=3.24 $Y2=1.45
r171 30 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.095 $Y=2.905
+ $X2=3.18 $Y2=2.99
r172 29 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=2.14
+ $X2=3.095 $Y2=2.055
r173 29 30 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=3.095 $Y=2.14
+ $X2=3.095 $Y2=2.905
r174 28 49 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.475 $Y=1.215
+ $X2=2.305 $Y2=1.215
r175 27 62 2.15123 $w=3.73e-07 $l=7e-08 $layer=LI1_cond $X=3.342 $Y=1.215
+ $X2=3.342 $Y2=1.285
r176 27 28 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.155 $Y=1.215
+ $X2=2.475 $Y2=1.215
r177 26 54 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.39 $Y=2.14
+ $X2=2.39 $Y2=1.55
r178 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.305 $Y=2.225
+ $X2=2.39 $Y2=2.14
r179 23 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.305 $Y=2.225
+ $X2=1.625 $Y2=2.225
r180 22 47 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.54 $Y=2.1 $X2=1.54
+ $Y2=2.29
r181 22 43 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=1.54 $Y=2.1
+ $X2=1.54 $Y2=1.09
r182 17 71 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.84 $Y=2.38
+ $X2=3.84 $Y2=2.215
r183 17 19 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=3.84 $Y=2.38
+ $X2=3.84 $Y2=2.75
r184 16 69 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.275 $Y=0.69
+ $X2=3.275 $Y2=1.12
r185 12 67 322.629 $w=1.8e-07 $l=8.3e-07 $layer=POLY_cond $X=2.28 $Y=2.38
+ $X2=2.28 $Y2=1.55
r186 9 66 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.175 $Y=0.74
+ $X2=2.175 $Y2=1.22
r187 2 45 600 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_PDIFF $count=1 $X=1.275
+ $Y=2.12 $X2=1.41 $Y2=2.29
r188 1 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.15
+ $Y=0.37 $X2=1.29 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_2%A_27_112# 1 2 9 13 15 19 22 25 26 27 28 31
+ 32 34 35 40 41
c102 40 0 2.18845e-19 $X=2.825 $Y=1.635
c103 31 0 2.08259e-19 $X=2.745 $Y=2.48
c104 9 0 4.2215e-20 $X=2.885 $Y=0.69
r105 41 46 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.825 $Y=1.635
+ $X2=2.825 $Y2=1.8
r106 41 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.825 $Y=1.635
+ $X2=2.825 $Y2=1.47
r107 40 43 8.46017 $w=3.23e-07 $l=1.65e-07 $layer=LI1_cond $X=2.822 $Y=1.635
+ $X2=2.822 $Y2=1.8
r108 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.825
+ $Y=1.635 $X2=2.825 $Y2=1.635
r109 35 37 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.88 $Y=2.565
+ $X2=1.88 $Y2=2.735
r110 31 43 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.745 $Y=2.48
+ $X2=2.745 $Y2=1.8
r111 29 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.965 $Y=2.565
+ $X2=1.88 $Y2=2.565
r112 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.66 $Y=2.565
+ $X2=2.745 $Y2=2.48
r113 28 29 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.66 $Y=2.565
+ $X2=1.965 $Y2=2.565
r114 26 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=2.735
+ $X2=1.88 $Y2=2.735
r115 26 27 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.795 $Y=2.735
+ $X2=1.155 $Y2=2.735
r116 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.07 $Y=2.65
+ $X2=1.155 $Y2=2.735
r117 24 25 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.07 $Y=2.27
+ $X2=1.07 $Y2=2.65
r118 23 34 2.98021 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.445 $Y=2.185
+ $X2=0.265 $Y2=2.185
r119 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.985 $Y=2.185
+ $X2=1.07 $Y2=2.27
r120 22 23 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=0.985 $Y=2.185
+ $X2=0.445 $Y2=2.185
r121 19 34 3.52026 $w=2.65e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.17 $Y=2.1
+ $X2=0.265 $Y2=2.185
r122 19 32 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=0.17 $Y=2.1
+ $X2=0.17 $Y2=1.09
r123 15 32 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.265 $Y=0.91
+ $X2=0.265 $Y2=1.09
r124 15 17 3.21944 $w=3.6e-07 $l=9.5e-08 $layer=LI1_cond $X=0.265 $Y=0.91
+ $X2=0.265 $Y2=0.815
r125 13 46 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.9 $Y=2.46 $X2=2.9
+ $Y2=1.8
r126 9 45 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.885 $Y=0.69
+ $X2=2.885 $Y2=1.47
r127 2 34 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.265
r128 1 17 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.28 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_2%A_363_74# 1 2 7 9 10 11 14 18 21 22 25 26 30
+ 35 36
c103 36 0 1.2913e-19 $X=3.965 $Y=1.39
c104 26 0 4.2215e-20 $X=1.96 $Y=0.87
c105 25 0 5.79271e-20 $X=3.8 $Y=1.225
c106 22 0 1.49993e-19 $X=3.715 $Y=0.865
c107 14 0 1.15905e-19 $X=3.875 $Y=0.58
c108 11 0 2.84074e-19 $X=3.38 $Y=1.765
r109 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.965
+ $Y=1.39 $X2=3.965 $Y2=1.39
r110 27 30 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.88 $Y=1.845
+ $X2=1.97 $Y2=1.845
r111 25 35 6.03661 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=3.8 $Y=1.382
+ $X2=3.965 $Y2=1.382
r112 24 25 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.8 $Y=0.95
+ $X2=3.8 $Y2=1.225
r113 23 26 2.76166 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=2.125 $Y=0.865
+ $X2=1.96 $Y2=0.87
r114 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.715 $Y=0.865
+ $X2=3.8 $Y2=0.95
r115 22 23 103.733 $w=1.68e-07 $l=1.59e-06 $layer=LI1_cond $X=3.715 $Y=0.865
+ $X2=2.125 $Y2=0.865
r116 21 27 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.88 $Y=1.72
+ $X2=1.88 $Y2=1.845
r117 20 26 3.70735 $w=2.5e-07 $l=1.23693e-07 $layer=LI1_cond $X=1.88 $Y=0.96
+ $X2=1.96 $Y2=0.87
r118 20 21 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=1.88 $Y=0.96
+ $X2=1.88 $Y2=1.72
r119 16 26 3.70735 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=1.96 $Y=0.78 $X2=1.96
+ $Y2=0.87
r120 16 18 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=1.96 $Y=0.78
+ $X2=1.96 $Y2=0.515
r121 12 36 39.6178 $w=2.46e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.875 $Y=1.225
+ $X2=3.965 $Y2=1.39
r122 12 14 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=3.875 $Y=1.225
+ $X2=3.875 $Y2=0.58
r123 10 36 73.4756 $w=2.46e-07 $l=4.5e-07 $layer=POLY_cond $X=3.8 $Y=1.765
+ $X2=3.965 $Y2=1.39
r124 10 11 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.8 $Y=1.765
+ $X2=3.38 $Y2=1.765
r125 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.29 $Y=1.84
+ $X2=3.38 $Y2=1.765
r126 7 9 166.022 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=3.29 $Y=1.84 $X2=3.29
+ $Y2=2.46
r127 2 30 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.74 $X2=1.97 $Y2=1.885
r128 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.815
+ $Y=0.37 $X2=1.96 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_2%A_838_48# 1 2 7 9 14 18 22 28 32 36 40 44 46
+ 47 50 53 54 56 58 61 63 71 76 79 83
c171 71 0 1.27392e-19 $X=6.79 $Y=1.485
c172 61 0 1.25688e-19 $X=6.87 $Y=2.24
c173 44 0 1.1451e-19 $X=4.45 $Y=0.94
c174 7 0 9.34102e-20 $X=4.265 $Y=0.865
r175 82 83 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=7.155 $Y=1.485
+ $X2=7.165 $Y2=1.485
r176 78 80 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.65 $Y=1.485
+ $X2=6.665 $Y2=1.485
r177 78 79 33.0969 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.65 $Y=1.485
+ $X2=6.56 $Y2=1.485
r178 72 82 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=6.79 $Y=1.485
+ $X2=7.155 $Y2=1.485
r179 72 80 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=6.79 $Y=1.485
+ $X2=6.665 $Y2=1.485
r180 71 74 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.79 $Y=1.485
+ $X2=6.79 $Y2=1.65
r181 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.79
+ $Y=1.485 $X2=6.79 $Y2=1.485
r182 68 69 3.80299 $w=4.01e-07 $l=1.25e-07 $layer=LI1_cond $X=5.435 $Y=2.2
+ $X2=5.435 $Y2=2.325
r183 67 68 6.54115 $w=4.01e-07 $l=2.15e-07 $layer=LI1_cond $X=5.435 $Y=1.985
+ $X2=5.435 $Y2=2.2
r184 63 65 19.9249 $w=5.23e-07 $l=6.15e-07 $layer=LI1_cond $X=5.137 $Y=0.515
+ $X2=5.137 $Y2=1.13
r185 61 74 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=6.87 $Y=2.24
+ $X2=6.87 $Y2=1.65
r186 59 69 5.79359 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=5.64 $Y=2.325
+ $X2=5.435 $Y2=2.325
r187 58 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.785 $Y=2.325
+ $X2=6.87 $Y2=2.24
r188 58 59 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=6.785 $Y=2.325
+ $X2=5.64 $Y2=2.325
r189 54 69 3.0046 $w=4.01e-07 $l=1.03078e-07 $layer=LI1_cond $X=5.475 $Y=2.41
+ $X2=5.435 $Y2=2.325
r190 54 56 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=5.475 $Y=2.41
+ $X2=5.475 $Y2=2.815
r191 53 67 9.15896 $w=4.01e-07 $l=2.16852e-07 $layer=LI1_cond $X=5.315 $Y=1.82
+ $X2=5.435 $Y2=1.985
r192 53 65 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.315 $Y=1.82
+ $X2=5.315 $Y2=1.13
r193 50 77 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.54 $Y=2.2
+ $X2=4.54 $Y2=2.365
r194 50 76 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.54 $Y=2.2
+ $X2=4.54 $Y2=2.035
r195 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.54
+ $Y=2.2 $X2=4.54 $Y2=2.2
r196 47 68 2.43857 $w=3e-07 $l=2.05e-07 $layer=LI1_cond $X=5.23 $Y=2.2 $X2=5.435
+ $Y2=2.2
r197 47 49 26.5062 $w=2.98e-07 $l=6.9e-07 $layer=LI1_cond $X=5.23 $Y=2.2
+ $X2=4.54 $Y2=2.2
r198 42 44 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=4.265 $Y=0.94
+ $X2=4.45 $Y2=0.94
r199 38 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.165 $Y=1.32
+ $X2=7.165 $Y2=1.485
r200 38 40 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=7.165 $Y=1.32
+ $X2=7.165 $Y2=0.69
r201 34 82 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.155 $Y=1.65
+ $X2=7.155 $Y2=1.485
r202 34 36 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=7.155 $Y=1.65
+ $X2=7.155 $Y2=2.34
r203 30 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.665 $Y=1.32
+ $X2=6.665 $Y2=1.485
r204 30 32 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.665 $Y=1.32
+ $X2=6.665 $Y2=0.74
r205 26 78 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.65 $Y=1.65
+ $X2=6.65 $Y2=1.485
r206 26 28 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=6.65 $Y=1.65
+ $X2=6.65 $Y2=2.4
r207 25 46 6.66866 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=6.31 $Y=1.395
+ $X2=6.21 $Y2=1.395
r208 25 79 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=6.31 $Y=1.395
+ $X2=6.56 $Y2=1.395
r209 20 46 18.8402 $w=1.65e-07 $l=8.66025e-08 $layer=POLY_cond $X=6.235 $Y=1.32
+ $X2=6.21 $Y2=1.395
r210 20 22 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.235 $Y=1.32
+ $X2=6.235 $Y2=0.74
r211 16 46 18.8402 $w=1.65e-07 $l=7.98436e-08 $layer=POLY_cond $X=6.2 $Y=1.47
+ $X2=6.21 $Y2=1.395
r212 16 18 361.5 $w=1.8e-07 $l=9.3e-07 $layer=POLY_cond $X=6.2 $Y=1.47 $X2=6.2
+ $Y2=2.4
r213 14 77 149.653 $w=1.8e-07 $l=3.85e-07 $layer=POLY_cond $X=4.465 $Y=2.75
+ $X2=4.465 $Y2=2.365
r214 10 44 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.45 $Y=1.015
+ $X2=4.45 $Y2=0.94
r215 10 76 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=4.45 $Y=1.015
+ $X2=4.45 $Y2=2.035
r216 7 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.265 $Y=0.865
+ $X2=4.265 $Y2=0.94
r217 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.265 $Y=0.865
+ $X2=4.265 $Y2=0.58
r218 2 67 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.33
+ $Y=1.84 $X2=5.475 $Y2=1.985
r219 2 56 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=5.33
+ $Y=1.84 $X2=5.475 $Y2=2.815
r220 1 63 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.895
+ $Y=0.37 $X2=5.04 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_2%A_670_74# 1 2 9 13 15 16 17 23 24 26 28 29
+ 33 37 38 42 44
c109 38 0 4.74009e-20 $X=3.507 $Y=2.405
c110 24 0 4.17599e-20 $X=3.665 $Y=1.795
r111 40 42 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=4.14 $Y=0.97
+ $X2=4.385 $Y2=0.97
r112 37 38 8.46257 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=3.507 $Y=2.57
+ $X2=3.507 $Y2=2.405
r113 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.9
+ $Y=1.515 $X2=4.9 $Y2=1.515
r114 31 33 6.91466 $w=3.23e-07 $l=1.95e-07 $layer=LI1_cond $X=4.897 $Y=1.71
+ $X2=4.897 $Y2=1.515
r115 30 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.47 $Y=1.795
+ $X2=4.385 $Y2=1.795
r116 29 31 7.72402 $w=1.7e-07 $l=2.00035e-07 $layer=LI1_cond $X=4.735 $Y=1.795
+ $X2=4.897 $Y2=1.71
r117 29 30 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.735 $Y=1.795
+ $X2=4.47 $Y2=1.795
r118 28 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.385 $Y=1.71
+ $X2=4.385 $Y2=1.795
r119 27 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.385 $Y=1.055
+ $X2=4.385 $Y2=0.97
r120 27 28 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.385 $Y=1.055
+ $X2=4.385 $Y2=1.71
r121 26 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=0.885
+ $X2=4.14 $Y2=0.97
r122 25 26 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.14 $Y=0.61
+ $X2=4.14 $Y2=0.885
r123 23 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=1.795
+ $X2=4.385 $Y2=1.795
r124 23 24 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.3 $Y=1.795
+ $X2=3.665 $Y2=1.795
r125 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.58 $Y=1.88
+ $X2=3.665 $Y2=1.795
r126 21 38 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.58 $Y=1.88
+ $X2=3.58 $Y2=2.405
r127 17 25 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.055 $Y=0.485
+ $X2=4.14 $Y2=0.61
r128 17 19 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=4.055 $Y=0.485
+ $X2=3.575 $Y2=0.485
r129 15 34 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=5.15 $Y=1.515
+ $X2=4.9 $Y2=1.515
r130 15 16 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.15 $Y=1.515
+ $X2=5.24 $Y2=1.515
r131 11 16 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=5.255 $Y=1.35
+ $X2=5.24 $Y2=1.515
r132 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.255 $Y=1.35
+ $X2=5.255 $Y2=0.74
r133 7 16 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=5.24 $Y=1.68
+ $X2=5.24 $Y2=1.515
r134 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.24 $Y=1.68 $X2=5.24
+ $Y2=2.4
r135 2 37 600 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=1 $X=3.38
+ $Y=1.96 $X2=3.52 $Y2=2.57
r136 1 19 182 $w=1.7e-07 $l=2.92404e-07 $layer=licon1_NDIFF $count=1 $X=3.35
+ $Y=0.37 $X2=3.575 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_2%RESET_B 3 6 8 11 13
c39 13 0 2.4962e-20 $X=5.735 $Y=1.22
r40 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.735 $Y=1.385
+ $X2=5.735 $Y2=1.55
r41 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.735 $Y=1.385
+ $X2=5.735 $Y2=1.22
r42 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.735
+ $Y=1.385 $X2=5.735 $Y2=1.385
r43 8 12 8.25398 $w=3.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6 $Y=1.365 $X2=5.735
+ $Y2=1.365
r44 6 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=5.7 $Y=2.4 $X2=5.7
+ $Y2=1.55
r45 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.645 $Y=0.74
+ $X2=5.645 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_2%A_1448_74# 1 2 9 11 13 14 18 20 22 23 24 25
+ 28 32 38 41
c68 23 0 1.27392e-19 $X=8.075 $Y=1.385
r69 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.065
+ $Y=1.385 $X2=8.065 $Y2=1.385
r70 36 41 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.545 $Y=1.385
+ $X2=7.38 $Y2=1.385
r71 36 38 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=7.545 $Y=1.385
+ $X2=8.065 $Y2=1.385
r72 32 34 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=7.38 $Y=1.985
+ $X2=7.38 $Y2=2.695
r73 30 41 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.38 $Y=1.55
+ $X2=7.38 $Y2=1.385
r74 30 32 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=7.38 $Y=1.55
+ $X2=7.38 $Y2=1.985
r75 26 41 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.38 $Y=1.22
+ $X2=7.38 $Y2=1.385
r76 26 28 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=7.38 $Y=1.22
+ $X2=7.38 $Y2=0.515
r77 23 39 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=8.075 $Y=1.385
+ $X2=8.065 $Y2=1.385
r78 23 24 7.86782 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.075 $Y=1.385
+ $X2=8.075 $Y2=1.22
r79 20 25 18.8402 $w=1.65e-07 $l=1e-07 $layer=POLY_cond $X=8.625 $Y=1.22
+ $X2=8.525 $Y2=1.22
r80 20 22 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.625 $Y=1.22
+ $X2=8.625 $Y2=0.74
r81 16 25 18.8402 $w=1.65e-07 $l=2.81425e-07 $layer=POLY_cond $X=8.615 $Y=1.46
+ $X2=8.525 $Y2=1.22
r82 16 18 365.387 $w=1.8e-07 $l=9.4e-07 $layer=POLY_cond $X=8.615 $Y=1.46
+ $X2=8.615 $Y2=2.4
r83 15 24 7.86782 $w=1.5e-07 $l=1.88812e-07 $layer=POLY_cond $X=8.23 $Y=1.295
+ $X2=8.075 $Y2=1.22
r84 14 25 6.66866 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.525 $Y=1.295
+ $X2=8.525 $Y2=1.22
r85 14 15 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=8.525 $Y=1.295
+ $X2=8.23 $Y2=1.295
r86 11 24 16.8416 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=8.155 $Y=1.22
+ $X2=8.075 $Y2=1.22
r87 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.155 $Y=1.22
+ $X2=8.155 $Y2=0.74
r88 7 24 16.8416 $w=1.8e-07 $l=5.23068e-07 $layer=POLY_cond $X=8.165 $Y=1.7
+ $X2=8.075 $Y2=1.22
r89 7 9 272.097 $w=1.8e-07 $l=7e-07 $layer=POLY_cond $X=8.165 $Y=1.7 $X2=8.165
+ $Y2=2.4
r90 2 34 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=7.245
+ $Y=1.84 $X2=7.38 $Y2=2.695
r91 2 32 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.245
+ $Y=1.84 $X2=7.38 $Y2=1.985
r92 1 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.24
+ $Y=0.37 $X2=7.38 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_2%VPWR 1 2 3 4 5 6 7 26 30 34 38 42 46 48 53
+ 54 55 57 65 70 79 83 89 92 95 104 107 111
r118 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r119 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r120 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r121 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r122 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r123 87 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r124 87 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r125 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r126 84 107 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=7.9 $Y2=3.33
r127 84 86 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=8.4 $Y2=3.33
r128 83 110 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=8.755 $Y=3.33
+ $X2=8.937 $Y2=3.33
r129 83 86 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.755 $Y=3.33
+ $X2=8.4 $Y2=3.33
r130 82 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r131 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r132 79 107 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.775 $Y=3.33
+ $X2=7.9 $Y2=3.33
r133 79 81 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.775 $Y=3.33
+ $X2=7.44 $Y2=3.33
r134 78 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r135 78 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r136 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r137 75 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.14 $Y=3.33
+ $X2=5.975 $Y2=3.33
r138 75 77 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.14 $Y=3.33
+ $X2=6.48 $Y2=3.33
r139 74 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r140 74 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r141 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r142 71 73 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=5.14 $Y=3.33
+ $X2=5.52 $Y2=3.33
r143 70 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.81 $Y=3.33
+ $X2=5.975 $Y2=3.33
r144 70 73 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.81 $Y=3.33
+ $X2=5.52 $Y2=3.33
r145 69 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r146 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r147 66 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=2.59 $Y2=3.33
r148 66 68 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=3.12 $Y2=3.33
r149 65 71 8.47627 $w=1.7e-07 $l=3.08e-07 $layer=LI1_cond $X=4.832 $Y=3.33
+ $X2=5.14 $Y2=3.33
r150 65 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r151 65 95 10.0159 $w=6.13e-07 $l=5.15e-07 $layer=LI1_cond $X=4.832 $Y=3.33
+ $X2=4.832 $Y2=2.815
r152 65 68 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=4.525 $Y=3.33
+ $X2=3.12 $Y2=3.33
r153 64 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r154 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r155 61 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r156 61 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r157 60 63 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r158 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r159 58 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.73 $Y2=3.33
r160 58 60 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=1.2 $Y2=3.33
r161 57 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.425 $Y=3.33
+ $X2=2.59 $Y2=3.33
r162 57 63 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.425 $Y=3.33
+ $X2=2.16 $Y2=3.33
r163 55 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r164 55 69 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=3.12 $Y2=3.33
r165 55 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r166 53 77 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.71 $Y=3.33
+ $X2=6.48 $Y2=3.33
r167 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.71 $Y=3.33
+ $X2=6.875 $Y2=3.33
r168 52 81 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=7.04 $Y=3.33 $X2=7.44
+ $Y2=3.33
r169 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.04 $Y=3.33
+ $X2=6.875 $Y2=3.33
r170 48 51 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=8.88 $Y=1.985
+ $X2=8.88 $Y2=2.815
r171 46 110 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.88 $Y=3.245
+ $X2=8.937 $Y2=3.33
r172 46 51 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.88 $Y=3.245
+ $X2=8.88 $Y2=2.815
r173 42 45 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=7.9 $Y=1.985
+ $X2=7.9 $Y2=2.815
r174 40 107 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=3.245
+ $X2=7.9 $Y2=3.33
r175 40 45 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.9 $Y=3.245 $X2=7.9
+ $Y2=2.815
r176 36 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.875 $Y=3.245
+ $X2=6.875 $Y2=3.33
r177 36 38 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=6.875 $Y=3.245
+ $X2=6.875 $Y2=2.68
r178 32 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.975 $Y=3.245
+ $X2=5.975 $Y2=3.33
r179 32 34 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=5.975 $Y=3.245
+ $X2=5.975 $Y2=2.78
r180 28 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=3.245
+ $X2=2.59 $Y2=3.33
r181 28 30 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.59 $Y=3.245
+ $X2=2.59 $Y2=2.985
r182 24 89 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r183 24 26 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.71
r184 7 51 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.705
+ $Y=1.84 $X2=8.84 $Y2=2.815
r185 7 48 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.705
+ $Y=1.84 $X2=8.84 $Y2=1.985
r186 6 45 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=7.795
+ $Y=1.84 $X2=7.94 $Y2=2.815
r187 6 42 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=7.795
+ $Y=1.84 $X2=7.94 $Y2=1.985
r188 5 38 600 $w=1.7e-07 $l=9.04986e-07 $layer=licon1_PDIFF $count=1 $X=6.74
+ $Y=1.84 $X2=6.875 $Y2=2.68
r189 4 34 600 $w=1.7e-07 $l=1.02835e-06 $layer=licon1_PDIFF $count=1 $X=5.79
+ $Y=1.84 $X2=5.975 $Y2=2.78
r190 3 95 600 $w=1.7e-07 $l=3.88909e-07 $layer=licon1_PDIFF $count=1 $X=4.555
+ $Y=2.54 $X2=4.83 $Y2=2.815
r191 2 30 600 $w=1.7e-07 $l=1.12966e-06 $layer=licon1_PDIFF $count=1 $X=2.37
+ $Y=1.96 $X2=2.59 $Y2=2.985
r192 1 26 600 $w=1.7e-07 $l=6.54026e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=2.12 $X2=0.73 $Y2=2.71
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_2%Q 1 2 10 11 13
c31 11 0 2.4962e-20 $X=6.425 $Y=1.82
r32 13 19 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=6.45 $Y=0.925
+ $X2=6.45 $Y2=1.13
r33 11 19 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.37 $Y=1.82 $X2=6.37
+ $Y2=1.13
r34 10 11 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.425 $Y=1.985
+ $X2=6.425 $Y2=1.82
r35 2 10 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.29
+ $Y=1.84 $X2=6.425 $Y2=1.985
r36 1 13 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=6.31
+ $Y=0.37 $X2=6.45 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_2%Q_N 1 2 12 14 15 16 23 32
r25 21 23 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=8.4 $Y=1.995 $X2=8.4
+ $Y2=2.035
r26 15 16 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=8.4 $Y=2.405 $X2=8.4
+ $Y2=2.775
r27 14 21 0.75732 $w=3.48e-07 $l=2.3e-08 $layer=LI1_cond $X=8.4 $Y=1.972 $X2=8.4
+ $Y2=1.995
r28 14 32 8.06043 $w=3.48e-07 $l=1.52e-07 $layer=LI1_cond $X=8.4 $Y=1.972
+ $X2=8.4 $Y2=1.82
r29 14 15 11.4586 $w=3.48e-07 $l=3.48e-07 $layer=LI1_cond $X=8.4 $Y=2.057
+ $X2=8.4 $Y2=2.405
r30 14 23 0.724393 $w=3.48e-07 $l=2.2e-08 $layer=LI1_cond $X=8.4 $Y=2.057
+ $X2=8.4 $Y2=2.035
r31 10 12 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=8.39 $Y=0.965 $X2=8.49
+ $Y2=0.965
r32 7 12 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.49 $Y=1.05 $X2=8.49
+ $Y2=0.965
r33 7 32 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=8.49 $Y=1.05 $X2=8.49
+ $Y2=1.82
r34 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.255
+ $Y=1.84 $X2=8.39 $Y2=1.985
r35 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.255
+ $Y=1.84 $X2=8.39 $Y2=2.815
r36 1 10 182 $w=1.7e-07 $l=6.70242e-07 $layer=licon1_NDIFF $count=1 $X=8.23
+ $Y=0.37 $X2=8.39 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_2%VGND 1 2 3 4 5 6 7 24 30 34 38 42 44 46 49
+ 50 51 53 58 66 78 82 87 93 97 103 106 109 113
r102 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r103 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r104 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r105 97 100 11.407 $w=5.38e-07 $l=5.15e-07 $layer=LI1_cond $X=2.565 $Y=0
+ $X2=2.565 $Y2=0.515
r106 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r107 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r108 91 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r109 91 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r110 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r111 88 109 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.035 $Y=0
+ $X2=7.905 $Y2=0
r112 88 90 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.035 $Y=0 $X2=8.4
+ $Y2=0
r113 87 112 4.09935 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=8.745 $Y=0
+ $X2=8.932 $Y2=0
r114 87 90 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.745 $Y=0 $X2=8.4
+ $Y2=0
r115 86 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r116 86 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.96 $Y2=0
r117 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r118 83 106 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.045 $Y=0
+ $X2=6.915 $Y2=0
r119 83 85 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=7.045 $Y=0
+ $X2=7.44 $Y2=0
r120 82 109 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.775 $Y=0
+ $X2=7.905 $Y2=0
r121 82 85 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.775 $Y=0
+ $X2=7.44 $Y2=0
r122 81 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r123 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r124 78 106 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.785 $Y=0
+ $X2=6.915 $Y2=0
r125 78 80 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.785 $Y=0
+ $X2=6.48 $Y2=0
r126 77 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r127 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r128 74 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.645 $Y=0
+ $X2=4.52 $Y2=0
r129 74 76 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=4.645 $Y=0
+ $X2=5.52 $Y2=0
r130 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r131 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r132 70 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r133 69 72 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r134 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r135 67 97 7.6426 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=2.835 $Y=0 $X2=2.565
+ $Y2=0
r136 67 69 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.835 $Y=0
+ $X2=3.12 $Y2=0
r137 66 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.395 $Y=0
+ $X2=4.52 $Y2=0
r138 66 72 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.395 $Y=0
+ $X2=4.08 $Y2=0
r139 65 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r140 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r141 62 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r142 62 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r143 61 64 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r144 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r145 59 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r146 59 61 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r147 58 97 7.6426 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.565
+ $Y2=0
r148 58 64 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.295 $Y=0
+ $X2=2.16 $Y2=0
r149 56 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r150 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r151 53 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r152 53 55 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r153 51 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r154 51 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r155 51 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r156 49 76 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.695 $Y=0
+ $X2=5.52 $Y2=0
r157 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.695 $Y=0 $X2=5.86
+ $Y2=0
r158 48 80 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=6.025 $Y=0
+ $X2=6.48 $Y2=0
r159 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.025 $Y=0 $X2=5.86
+ $Y2=0
r160 44 112 3.11287 $w=2.6e-07 $l=1.09864e-07 $layer=LI1_cond $X=8.875 $Y=0.085
+ $X2=8.932 $Y2=0
r161 44 46 19.7245 $w=2.58e-07 $l=4.45e-07 $layer=LI1_cond $X=8.875 $Y=0.085
+ $X2=8.875 $Y2=0.53
r162 40 109 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.905 $Y=0.085
+ $X2=7.905 $Y2=0
r163 40 42 19.7245 $w=2.58e-07 $l=4.45e-07 $layer=LI1_cond $X=7.905 $Y=0.085
+ $X2=7.905 $Y2=0.53
r164 36 106 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.915 $Y=0.085
+ $X2=6.915 $Y2=0
r165 36 38 19.0596 $w=2.58e-07 $l=4.3e-07 $layer=LI1_cond $X=6.915 $Y=0.085
+ $X2=6.915 $Y2=0.515
r166 32 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.86 $Y=0.085
+ $X2=5.86 $Y2=0
r167 32 34 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.86 $Y=0.085
+ $X2=5.86 $Y2=0.515
r168 28 103 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.52 $Y=0.085
+ $X2=4.52 $Y2=0
r169 28 30 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=4.52 $Y=0.085
+ $X2=4.52 $Y2=0.53
r170 24 26 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=0.79 $Y=0.53
+ $X2=0.79 $Y2=0.925
r171 22 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0
r172 22 24 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0.53
r173 7 46 91 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=2 $X=8.7
+ $Y=0.37 $X2=8.84 $Y2=0.53
r174 6 42 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=7.795
+ $Y=0.37 $X2=7.94 $Y2=0.53
r175 5 38 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.74
+ $Y=0.37 $X2=6.88 $Y2=0.515
r176 4 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.72
+ $Y=0.37 $X2=5.86 $Y2=0.515
r177 3 30 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=4.34
+ $Y=0.37 $X2=4.48 $Y2=0.53
r178 2 100 182 $w=1.7e-07 $l=3.80657e-07 $layer=licon1_NDIFF $count=1 $X=2.25
+ $Y=0.37 $X2=2.565 $Y2=0.515
r179 1 26 182 $w=1.7e-07 $l=4.62088e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.56 $X2=0.79 $Y2=0.925
r180 1 24 182 $w=1.7e-07 $l=2.34521e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.56 $X2=0.79 $Y2=0.53
.ends


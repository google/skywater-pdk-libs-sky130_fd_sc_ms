* File: sky130_fd_sc_ms__a32o_1.pex.spice
* Created: Fri Aug 28 17:07:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A32O_1%A_84_48# 1 2 9 13 16 18 19 23 28 29 32 33
r93 32 33 17.1863 $w=5.88e-07 $l=5.15e-07 $layer=LI1_cond $X=2.715 $Y=0.725
+ $X2=2.2 $Y2=0.725
r94 29 37 40.6969 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.587 $Y=1.465
+ $X2=0.587 $Y2=1.63
r95 29 36 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=0.587 $Y=1.465
+ $X2=0.587 $Y2=1.3
r96 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.465 $X2=0.59 $Y2=1.465
r97 23 25 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.06 $Y=1.97
+ $X2=3.06 $Y2=2.65
r98 21 23 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.06 $Y=1.89 $X2=3.06
+ $Y2=1.97
r99 20 28 14.7616 $w=2.81e-07 $l=4.22493e-07 $layer=LI1_cond $X=0.795 $Y=1.805
+ $X2=0.61 $Y2=1.465
r100 19 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.895 $Y=1.805
+ $X2=3.06 $Y2=1.89
r101 19 20 137.005 $w=1.68e-07 $l=2.1e-06 $layer=LI1_cond $X=2.895 $Y=1.805
+ $X2=0.795 $Y2=1.805
r102 18 33 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=0.795 $Y=0.935
+ $X2=2.2 $Y2=0.935
r103 16 28 9.05323 $w=2.81e-07 $l=2.09105e-07 $layer=LI1_cond $X=0.71 $Y=1.3
+ $X2=0.61 $Y2=1.465
r104 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.71 $Y=1.02
+ $X2=0.795 $Y2=0.935
r105 15 16 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.71 $Y=1.02
+ $X2=0.71 $Y2=1.3
r106 13 37 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.515 $Y=2.4
+ $X2=0.515 $Y2=1.63
r107 9 36 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=0.74
+ $X2=0.495 $Y2=1.3
r108 2 25 400 $w=1.7e-07 $l=8.97747e-07 $layer=licon1_PDIFF $count=1 $X=2.875
+ $Y=1.84 $X2=3.06 $Y2=2.65
r109 2 23 400 $w=1.7e-07 $l=2.41402e-07 $layer=licon1_PDIFF $count=1 $X=2.875
+ $Y=1.84 $X2=3.06 $Y2=1.97
r110 1 32 45.5 $w=1.7e-07 $l=5.48954e-07 $layer=licon1_NDIFF $count=4 $X=2.225
+ $Y=0.47 $X2=2.715 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_1%A3 3 7 8 11 13
c37 13 0 9.95713e-20 $X=1.13 $Y=1.22
c38 8 0 9.8332e-20 $X=1.2 $Y=1.295
r39 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.385
+ $X2=1.13 $Y2=1.55
r40 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.385
+ $X2=1.13 $Y2=1.22
r41 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.385 $X2=1.13 $Y2=1.385
r42 8 12 2.96342 $w=3.48e-07 $l=9e-08 $layer=LI1_cond $X=1.14 $Y=1.295 $X2=1.14
+ $Y2=1.385
r43 7 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.22 $Y=0.79 $X2=1.22
+ $Y2=1.22
r44 3 14 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=1.145 $Y=2.34
+ $X2=1.145 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_1%A2 3 7 8 11 13
c31 13 0 1.83337e-19 $X=1.67 $Y=1.22
c32 8 0 2.09874e-19 $X=1.68 $Y=1.295
r33 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.67 $Y=1.385
+ $X2=1.67 $Y2=1.55
r34 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.67 $Y=1.385
+ $X2=1.67 $Y2=1.22
r35 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.67
+ $Y=1.385 $X2=1.67 $Y2=1.385
r36 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.67 $Y=1.295 $X2=1.67
+ $Y2=1.385
r37 7 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.61 $Y=0.79 $X2=1.61
+ $Y2=1.22
r38 3 14 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=1.595 $Y=2.34
+ $X2=1.595 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_1%A1 1 3 6 8 15
c33 8 0 1.47811e-19 $X=2.16 $Y=1.295
c34 1 0 2.02667e-19 $X=2.15 $Y=1.22
r35 13 15 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=2.21 $Y=1.385
+ $X2=2.335 $Y2=1.385
r36 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.21
+ $Y=1.385 $X2=2.21 $Y2=1.385
r37 10 13 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.15 $Y=1.385 $X2=2.21
+ $Y2=1.385
r38 8 14 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.21 $Y=1.295 $X2=2.21
+ $Y2=1.385
r39 4 15 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.335 $Y=1.55
+ $X2=2.335 $Y2=1.385
r40 4 6 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=2.335 $Y=1.55
+ $X2=2.335 $Y2=2.34
r41 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.22
+ $X2=2.15 $Y2=1.385
r42 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.15 $Y=1.22 $X2=2.15
+ $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_1%B1 3 7 8 11 12 13
c32 13 0 6.28053e-20 $X=2.84 $Y=1.22
c33 12 0 9.23649e-20 $X=2.84 $Y=1.385
r34 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=1.385
+ $X2=2.84 $Y2=1.55
r35 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=1.385
+ $X2=2.84 $Y2=1.22
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.84
+ $Y=1.385 $X2=2.84 $Y2=1.385
r37 8 12 6.40246 $w=3.58e-07 $l=2e-07 $layer=LI1_cond $X=2.64 $Y=1.37 $X2=2.84
+ $Y2=1.37
r38 7 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.93 $Y=0.79 $X2=2.93
+ $Y2=1.22
r39 3 14 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=2.785 $Y=2.34
+ $X2=2.785 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_1%B2 3 6 8 11 13
r24 11 14 39.5669 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.432 $Y=1.385
+ $X2=3.432 $Y2=1.55
r25 11 13 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.432 $Y=1.385
+ $X2=3.432 $Y2=1.22
r26 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.455
+ $Y=1.385 $X2=3.455 $Y2=1.385
r27 8 12 4.91483 $w=3.38e-07 $l=1.45e-07 $layer=LI1_cond $X=3.6 $Y=1.38
+ $X2=3.455 $Y2=1.38
r28 6 14 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=3.335 $Y=2.34
+ $X2=3.335 $Y2=1.55
r29 3 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.32 $Y=0.79 $X2=3.32
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_1%X 1 2 11 14 15 16 17 28
r25 21 28 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.265 $Y=0.95
+ $X2=0.265 $Y2=0.925
r26 17 30 8.03084 $w=3.58e-07 $l=1.5e-07 $layer=LI1_cond $X=0.265 $Y=0.98
+ $X2=0.265 $Y2=1.13
r27 17 21 0.960369 $w=3.58e-07 $l=3e-08 $layer=LI1_cond $X=0.265 $Y=0.98
+ $X2=0.265 $Y2=0.95
r28 17 28 0.960369 $w=3.58e-07 $l=3e-08 $layer=LI1_cond $X=0.265 $Y=0.895
+ $X2=0.265 $Y2=0.925
r29 16 17 12.1647 $w=3.58e-07 $l=3.8e-07 $layer=LI1_cond $X=0.265 $Y=0.515
+ $X2=0.265 $Y2=0.895
r30 15 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.17 $Y=1.82 $X2=0.17
+ $Y2=1.13
r31 14 15 8.53881 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.27 $Y=1.985
+ $X2=0.27 $Y2=1.82
r32 9 14 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=0.27 $Y=2.005 $X2=0.27
+ $Y2=1.985
r33 9 11 25.2292 $w=3.68e-07 $l=8.1e-07 $layer=LI1_cond $X=0.27 $Y=2.005
+ $X2=0.27 $Y2=2.815
r34 2 14 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.29 $Y2=1.985
r35 2 11 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.29 $Y2=2.815
r36 1 16 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_1%VPWR 1 2 9 15 18 19 20 22 35 36 39
r44 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r46 33 36 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r47 32 35 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r48 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 30 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r51 27 39 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=0.82 $Y2=3.33
r52 27 29 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.015 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r55 22 39 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.82 $Y2=3.33
r56 22 24 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.24 $Y2=3.33
r57 20 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r58 20 30 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r59 18 29 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.8 $Y=3.33 $X2=1.68
+ $Y2=3.33
r60 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.8 $Y=3.33
+ $X2=1.965 $Y2=3.33
r61 17 32 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.13 $Y=3.33 $X2=2.16
+ $Y2=3.33
r62 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.13 $Y=3.33
+ $X2=1.965 $Y2=3.33
r63 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.965 $Y=3.245
+ $X2=1.965 $Y2=3.33
r64 13 15 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.965 $Y=3.245
+ $X2=1.965 $Y2=2.565
r65 9 12 17.4344 $w=3.88e-07 $l=5.9e-07 $layer=LI1_cond $X=0.82 $Y=2.225
+ $X2=0.82 $Y2=2.815
r66 7 39 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=3.245 $X2=0.82
+ $Y2=3.33
r67 7 12 12.7064 $w=3.88e-07 $l=4.3e-07 $layer=LI1_cond $X=0.82 $Y=3.245
+ $X2=0.82 $Y2=2.815
r68 2 15 600 $w=1.7e-07 $l=8.53595e-07 $layer=licon1_PDIFF $count=1 $X=1.685
+ $Y=1.84 $X2=1.965 $Y2=2.565
r69 1 12 600 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.84 $X2=0.79 $Y2=2.815
r70 1 9 600 $w=1.7e-07 $l=4.92494e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.84 $X2=0.85 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_1%A_247_368# 1 2 3 12 14 15 16 17 20 25
r40 20 23 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.56 $Y=1.985
+ $X2=3.56 $Y2=2.695
r41 18 23 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=3.56 $Y=2.905
+ $X2=3.56 $Y2=2.695
r42 16 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.395 $Y=2.99
+ $X2=3.56 $Y2=2.905
r43 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.395 $Y=2.99
+ $X2=2.725 $Y2=2.99
r44 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.56 $Y=2.905
+ $X2=2.725 $Y2=2.99
r45 14 27 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=2.23 $X2=2.56
+ $Y2=2.145
r46 14 15 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.56 $Y=2.23
+ $X2=2.56 $Y2=2.905
r47 13 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.535 $Y=2.145
+ $X2=1.37 $Y2=2.145
r48 12 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=2.145
+ $X2=2.56 $Y2=2.145
r49 12 13 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2.395 $Y=2.145
+ $X2=1.535 $Y2=2.145
r50 3 23 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=1.84 $X2=3.56 $Y2=2.695
r51 3 20 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=1.84 $X2=3.56 $Y2=1.985
r52 2 27 300 $w=1.7e-07 $l=4.01871e-07 $layer=licon1_PDIFF $count=2 $X=2.425
+ $Y=1.84 $X2=2.56 $Y2=2.18
r53 1 25 300 $w=1.7e-07 $l=4.01871e-07 $layer=licon1_PDIFF $count=2 $X=1.235
+ $Y=1.84 $X2=1.37 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_MS__A32O_1%VGND 1 2 11 13 15 17 19 28 32
r38 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r39 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r41 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r42 23 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r43 22 25 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r44 22 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r45 20 28 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=1.05 $Y=0 $X2=0.85
+ $Y2=0
r46 20 22 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.05 $Y=0 $X2=1.2
+ $Y2=0
r47 19 31 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.37 $Y=0 $X2=3.605
+ $Y2=0
r48 19 25 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.37 $Y=0 $X2=3.12
+ $Y2=0
r49 17 26 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=3.12
+ $Y2=0
r50 17 23 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r51 13 31 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=3.535 $Y=0.085
+ $X2=3.605 $Y2=0
r52 13 15 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=3.535 $Y=0.085
+ $X2=3.535 $Y2=0.615
r53 9 28 1.46811 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=0.085 $X2=0.85
+ $Y2=0
r54 9 11 13.2531 $w=3.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.85 $Y=0.085
+ $X2=0.85 $Y2=0.545
r55 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.395
+ $Y=0.47 $X2=3.535 $Y2=0.615
r56 1 11 182 $w=1.7e-07 $l=3.56931e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.85 $Y2=0.545
.ends


* File: sky130_fd_sc_ms__nand4b_2.pxi.spice
* Created: Wed Sep  2 12:14:38 2020
* 
x_PM_SKY130_FD_SC_MS__NAND4B_2%A_N N_A_N_M1010_g N_A_N_M1008_g A_N A_N
+ N_A_N_c_94_n N_A_N_c_95_n PM_SKY130_FD_SC_MS__NAND4B_2%A_N
x_PM_SKY130_FD_SC_MS__NAND4B_2%A_27_74# N_A_27_74#_M1010_s N_A_27_74#_M1008_s
+ N_A_27_74#_M1011_g N_A_27_74#_M1002_g N_A_27_74#_M1016_g N_A_27_74#_M1015_g
+ N_A_27_74#_c_126_n N_A_27_74#_c_127_n N_A_27_74#_c_128_n N_A_27_74#_c_134_n
+ N_A_27_74#_c_135_n N_A_27_74#_c_136_n N_A_27_74#_c_129_n N_A_27_74#_c_130_n
+ N_A_27_74#_c_131_n PM_SKY130_FD_SC_MS__NAND4B_2%A_27_74#
x_PM_SKY130_FD_SC_MS__NAND4B_2%B N_B_M1001_g N_B_M1012_g N_B_M1007_g N_B_M1017_g
+ B N_B_c_211_n N_B_c_212_n PM_SKY130_FD_SC_MS__NAND4B_2%B
x_PM_SKY130_FD_SC_MS__NAND4B_2%C N_C_M1009_g N_C_M1000_g N_C_M1014_g N_C_M1006_g
+ C C N_C_c_272_n PM_SKY130_FD_SC_MS__NAND4B_2%C
x_PM_SKY130_FD_SC_MS__NAND4B_2%D N_D_c_330_n N_D_M1004_g N_D_M1003_g N_D_c_327_n
+ N_D_M1013_g N_D_M1005_g D D D PM_SKY130_FD_SC_MS__NAND4B_2%D
x_PM_SKY130_FD_SC_MS__NAND4B_2%VPWR N_VPWR_M1008_d N_VPWR_M1016_s N_VPWR_M1017_s
+ N_VPWR_M1014_s N_VPWR_M1013_s N_VPWR_c_373_n N_VPWR_c_374_n N_VPWR_c_375_n
+ N_VPWR_c_376_n N_VPWR_c_377_n N_VPWR_c_378_n N_VPWR_c_379_n N_VPWR_c_380_n
+ VPWR N_VPWR_c_381_n N_VPWR_c_382_n N_VPWR_c_383_n N_VPWR_c_384_n
+ N_VPWR_c_385_n N_VPWR_c_386_n N_VPWR_c_387_n N_VPWR_c_372_n
+ PM_SKY130_FD_SC_MS__NAND4B_2%VPWR
x_PM_SKY130_FD_SC_MS__NAND4B_2%Y N_Y_M1002_s N_Y_M1011_d N_Y_M1012_d N_Y_M1009_d
+ N_Y_M1004_d N_Y_c_456_n N_Y_c_450_n N_Y_c_461_n N_Y_c_447_n N_Y_c_451_n
+ N_Y_c_478_n N_Y_c_452_n N_Y_c_497_n N_Y_c_512_n N_Y_c_453_n N_Y_c_448_n
+ N_Y_c_454_n N_Y_c_501_n Y Y PM_SKY130_FD_SC_MS__NAND4B_2%Y
x_PM_SKY130_FD_SC_MS__NAND4B_2%VGND N_VGND_M1010_d N_VGND_M1003_s N_VGND_c_549_n
+ N_VGND_c_550_n VGND N_VGND_c_551_n N_VGND_c_552_n N_VGND_c_553_n
+ N_VGND_c_554_n N_VGND_c_555_n N_VGND_c_556_n PM_SKY130_FD_SC_MS__NAND4B_2%VGND
x_PM_SKY130_FD_SC_MS__NAND4B_2%A_225_74# N_A_225_74#_M1002_d N_A_225_74#_M1015_d
+ N_A_225_74#_M1007_d N_A_225_74#_c_605_n N_A_225_74#_c_606_n
+ N_A_225_74#_c_607_n N_A_225_74#_c_619_n PM_SKY130_FD_SC_MS__NAND4B_2%A_225_74#
x_PM_SKY130_FD_SC_MS__NAND4B_2%A_490_74# N_A_490_74#_M1001_s N_A_490_74#_M1000_s
+ N_A_490_74#_c_642_n N_A_490_74#_c_648_n N_A_490_74#_c_643_n
+ PM_SKY130_FD_SC_MS__NAND4B_2%A_490_74#
x_PM_SKY130_FD_SC_MS__NAND4B_2%A_719_123# N_A_719_123#_M1000_d
+ N_A_719_123#_M1006_d N_A_719_123#_M1005_d N_A_719_123#_c_669_n
+ N_A_719_123#_c_670_n N_A_719_123#_c_671_n N_A_719_123#_c_672_n
+ N_A_719_123#_c_673_n N_A_719_123#_c_674_n N_A_719_123#_c_675_n
+ N_A_719_123#_c_676_n PM_SKY130_FD_SC_MS__NAND4B_2%A_719_123#
cc_1 VNB N_A_N_M1010_g 0.0318449f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_2 VNB N_A_N_M1008_g 0.0132343f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=2.34
cc_3 VNB N_A_N_c_94_n 0.0245924f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.345
cc_4 VNB N_A_N_c_95_n 0.0688576f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.345
cc_5 VNB N_A_27_74#_M1002_g 0.0266096f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.345
cc_6 VNB N_A_27_74#_M1015_g 0.0239157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_27_74#_c_126_n 0.0203664f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.345
cc_8 VNB N_A_27_74#_c_127_n 0.0105263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_74#_c_128_n 0.00949248f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_74#_c_129_n 0.00567489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_74#_c_130_n 0.00646829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_74#_c_131_n 0.0382628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B_M1001_g 0.0255964f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.69
cc_14 VNB N_B_M1007_g 0.0293822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_c_211_n 0.00465678f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.345
cc_16 VNB N_B_c_212_n 0.0553778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_C_M1000_g 0.023676f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=2.34
cc_18 VNB N_C_M1006_g 0.0200129f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.345
cc_19 VNB C 0.00377768f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.345
cc_20 VNB N_C_c_272_n 0.0575497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_D_M1003_g 0.0202431f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=2.34
cc_22 VNB N_D_c_327_n 0.0367312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_D_M1005_g 0.028245f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB D 0.0203907f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.345
cc_25 VNB N_VPWR_c_372_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_447_n 0.00841801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_448_n 0.00418682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB Y 0.0025475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_549_n 0.0100536f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_30 VNB N_VGND_c_550_n 0.0069637f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.345
cc_31 VNB N_VGND_c_551_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.345
cc_32 VNB N_VGND_c_552_n 0.0979637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_553_n 0.0183664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_554_n 0.332581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_555_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_556_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_225_74#_c_605_n 0.00846754f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_38 VNB N_A_225_74#_c_606_n 0.00194367f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.345
cc_39 VNB N_A_225_74#_c_607_n 0.00305483f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.345
cc_40 VNB N_A_490_74#_c_642_n 0.0219302f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=2.34
cc_41 VNB N_A_490_74#_c_643_n 0.00366476f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.345
cc_42 VNB N_A_719_123#_c_669_n 0.00392221f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_43 VNB N_A_719_123#_c_670_n 0.00551296f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.345
cc_44 VNB N_A_719_123#_c_671_n 0.00461713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_719_123#_c_672_n 0.00210056f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=1.345
cc_46 VNB N_A_719_123#_c_673_n 0.00323568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_719_123#_c_674_n 0.0131055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_719_123#_c_675_n 0.0220272f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.345
cc_49 VNB N_A_719_123#_c_676_n 0.00178419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VPB N_A_N_M1008_g 0.0281055f $X=-0.19 $Y=1.66 $X2=0.895 $Y2=2.34
cc_51 VPB N_A_27_74#_M1011_g 0.0233878f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_52 VPB N_A_27_74#_M1016_g 0.0247322f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=1.345
cc_53 VPB N_A_27_74#_c_134_n 0.0415136f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_A_27_74#_c_135_n 0.00256945f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_27_74#_c_136_n 0.0094432f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_27_74#_c_130_n 0.00300058f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_A_27_74#_c_131_n 0.00594884f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_B_M1012_g 0.0246086f $X=-0.19 $Y=1.66 $X2=0.895 $Y2=2.34
cc_59 VPB N_B_M1017_g 0.0221105f $X=-0.19 $Y=1.66 $X2=0.82 $Y2=1.345
cc_60 VPB N_B_c_211_n 0.00720696f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.345
cc_61 VPB N_B_c_212_n 0.0149393f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_C_M1009_g 0.0218585f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.69
cc_63 VPB N_C_M1014_g 0.0232614f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB C 0.00454411f $X=-0.19 $Y=1.66 $X2=0.895 $Y2=1.345
cc_65 VPB N_C_c_272_n 0.00732482f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_D_c_330_n 0.0180839f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.18
cc_67 VPB N_D_c_327_n 0.0103086f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_D_M1013_g 0.0246339f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_69 VPB D 0.0148561f $X=-0.19 $Y=1.66 $X2=0.895 $Y2=1.345
cc_70 VPB N_VPWR_c_373_n 0.0103004f $X=-0.19 $Y=1.66 $X2=0.895 $Y2=1.345
cc_71 VPB N_VPWR_c_374_n 0.0110015f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_375_n 0.00899828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_376_n 0.00987189f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_377_n 0.0113253f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_378_n 0.0508384f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_379_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_380_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_381_n 0.0332141f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_382_n 0.0175344f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_383_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_384_n 0.0199677f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_385_n 0.00613202f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_386_n 0.0114188f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_387_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_372_n 0.0884445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_86 VPB N_Y_c_450_n 0.00225166f $X=-0.19 $Y=1.66 $X2=0.895 $Y2=1.345
cc_87 VPB N_Y_c_451_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_Y_c_452_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_Y_c_453_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_Y_c_454_n 0.00262024f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB Y 0.00124879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 N_A_N_M1008_g N_A_27_74#_M1011_g 0.0153253f $X=0.895 $Y=2.34 $X2=0 $Y2=0
cc_93 N_A_N_c_95_n N_A_27_74#_M1002_g 0.00377133f $X=0.895 $Y=1.345 $X2=0 $Y2=0
cc_94 N_A_N_M1010_g N_A_27_74#_c_126_n 0.00264672f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_95 N_A_N_M1010_g N_A_27_74#_c_127_n 0.0143914f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_96 N_A_N_c_94_n N_A_27_74#_c_127_n 0.0415659f $X=0.82 $Y=1.345 $X2=0 $Y2=0
cc_97 N_A_N_c_95_n N_A_27_74#_c_127_n 0.00988866f $X=0.895 $Y=1.345 $X2=0 $Y2=0
cc_98 N_A_N_c_94_n N_A_27_74#_c_128_n 0.0204809f $X=0.82 $Y=1.345 $X2=0 $Y2=0
cc_99 N_A_N_c_95_n N_A_27_74#_c_128_n 0.00115581f $X=0.895 $Y=1.345 $X2=0 $Y2=0
cc_100 N_A_N_M1008_g N_A_27_74#_c_134_n 0.0144222f $X=0.895 $Y=2.34 $X2=0 $Y2=0
cc_101 N_A_N_M1008_g N_A_27_74#_c_135_n 0.0131281f $X=0.895 $Y=2.34 $X2=0 $Y2=0
cc_102 N_A_N_c_94_n N_A_27_74#_c_135_n 0.010678f $X=0.82 $Y=1.345 $X2=0 $Y2=0
cc_103 N_A_N_M1008_g N_A_27_74#_c_136_n 0.00411429f $X=0.895 $Y=2.34 $X2=0 $Y2=0
cc_104 N_A_N_c_94_n N_A_27_74#_c_136_n 0.0276947f $X=0.82 $Y=1.345 $X2=0 $Y2=0
cc_105 N_A_N_c_95_n N_A_27_74#_c_136_n 0.00724507f $X=0.895 $Y=1.345 $X2=0 $Y2=0
cc_106 N_A_N_M1010_g N_A_27_74#_c_129_n 0.0037584f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_107 N_A_N_c_94_n N_A_27_74#_c_129_n 0.013468f $X=0.82 $Y=1.345 $X2=0 $Y2=0
cc_108 N_A_N_c_95_n N_A_27_74#_c_129_n 5.96187e-19 $X=0.895 $Y=1.345 $X2=0 $Y2=0
cc_109 N_A_N_c_94_n N_A_27_74#_c_130_n 0.013971f $X=0.82 $Y=1.345 $X2=0 $Y2=0
cc_110 N_A_N_c_95_n N_A_27_74#_c_130_n 0.00529992f $X=0.895 $Y=1.345 $X2=0 $Y2=0
cc_111 N_A_N_c_95_n N_A_27_74#_c_131_n 0.0153253f $X=0.895 $Y=1.345 $X2=0 $Y2=0
cc_112 N_A_N_M1008_g N_VPWR_c_373_n 0.00777258f $X=0.895 $Y=2.34 $X2=0 $Y2=0
cc_113 N_A_N_M1008_g N_VPWR_c_381_n 0.00567889f $X=0.895 $Y=2.34 $X2=0 $Y2=0
cc_114 N_A_N_M1008_g N_VPWR_c_372_n 0.00610055f $X=0.895 $Y=2.34 $X2=0 $Y2=0
cc_115 N_A_N_M1010_g N_VGND_c_549_n 0.0115915f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_116 N_A_N_M1010_g N_VGND_c_551_n 0.00383152f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_117 N_A_N_M1010_g N_VGND_c_554_n 0.00387625f $X=0.495 $Y=0.69 $X2=0 $Y2=0
cc_118 N_A_N_M1010_g N_A_225_74#_c_605_n 6.17645e-19 $X=0.495 $Y=0.69 $X2=0
+ $Y2=0
cc_119 N_A_27_74#_M1015_g N_B_M1001_g 0.0334156f $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_120 N_A_27_74#_M1016_g N_B_M1012_g 0.0119814f $X=1.885 $Y=2.4 $X2=0 $Y2=0
cc_121 N_A_27_74#_M1016_g N_B_c_211_n 0.00332618f $X=1.885 $Y=2.4 $X2=0 $Y2=0
cc_122 N_A_27_74#_c_130_n N_B_c_211_n 0.017469f $X=1.555 $Y=1.515 $X2=0 $Y2=0
cc_123 N_A_27_74#_c_131_n N_B_c_211_n 0.0040727f $X=1.945 $Y=1.515 $X2=0 $Y2=0
cc_124 N_A_27_74#_c_130_n N_B_c_212_n 2.0756e-19 $X=1.555 $Y=1.515 $X2=0 $Y2=0
cc_125 N_A_27_74#_c_131_n N_B_c_212_n 0.0181293f $X=1.945 $Y=1.515 $X2=0 $Y2=0
cc_126 N_A_27_74#_c_135_n N_VPWR_M1008_d 0.00119058f $X=1.155 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_127 N_A_27_74#_c_130_n N_VPWR_M1008_d 0.00147181f $X=1.555 $Y=1.515 $X2=-0.19
+ $Y2=-0.245
cc_128 N_A_27_74#_M1011_g N_VPWR_c_373_n 0.0162707f $X=1.435 $Y=2.4 $X2=0 $Y2=0
cc_129 N_A_27_74#_M1016_g N_VPWR_c_373_n 6.15067e-19 $X=1.885 $Y=2.4 $X2=0 $Y2=0
cc_130 N_A_27_74#_c_134_n N_VPWR_c_373_n 0.0278269f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_131 N_A_27_74#_c_135_n N_VPWR_c_373_n 0.00915704f $X=1.155 $Y=1.765 $X2=0
+ $Y2=0
cc_132 N_A_27_74#_c_130_n N_VPWR_c_373_n 0.0135852f $X=1.555 $Y=1.515 $X2=0
+ $Y2=0
cc_133 N_A_27_74#_M1016_g N_VPWR_c_374_n 0.00256578f $X=1.885 $Y=2.4 $X2=0 $Y2=0
cc_134 N_A_27_74#_c_134_n N_VPWR_c_381_n 0.00975961f $X=0.67 $Y=1.985 $X2=0
+ $Y2=0
cc_135 N_A_27_74#_M1011_g N_VPWR_c_382_n 0.00475445f $X=1.435 $Y=2.4 $X2=0 $Y2=0
cc_136 N_A_27_74#_M1016_g N_VPWR_c_382_n 0.005209f $X=1.885 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A_27_74#_M1011_g N_VPWR_c_372_n 0.00938661f $X=1.435 $Y=2.4 $X2=0 $Y2=0
cc_138 N_A_27_74#_M1016_g N_VPWR_c_372_n 0.00984248f $X=1.885 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A_27_74#_c_134_n N_VPWR_c_372_n 0.0111753f $X=0.67 $Y=1.985 $X2=0 $Y2=0
cc_140 N_A_27_74#_M1016_g N_Y_c_456_n 0.00562475f $X=1.885 $Y=2.4 $X2=0 $Y2=0
cc_141 N_A_27_74#_c_130_n N_Y_c_456_n 0.0126667f $X=1.555 $Y=1.515 $X2=0 $Y2=0
cc_142 N_A_27_74#_c_131_n N_Y_c_456_n 7.0902e-19 $X=1.945 $Y=1.515 $X2=0 $Y2=0
cc_143 N_A_27_74#_M1011_g N_Y_c_450_n 2.47199e-19 $X=1.435 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A_27_74#_M1016_g N_Y_c_450_n 0.0160616f $X=1.885 $Y=2.4 $X2=0 $Y2=0
cc_145 N_A_27_74#_M1016_g N_Y_c_461_n 0.0188784f $X=1.885 $Y=2.4 $X2=0 $Y2=0
cc_146 N_A_27_74#_M1015_g N_Y_c_447_n 0.012995f $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A_27_74#_M1002_g N_Y_c_448_n 0.00727448f $X=1.485 $Y=0.74 $X2=0 $Y2=0
cc_148 N_A_27_74#_M1015_g N_Y_c_448_n 0.00682377f $X=1.945 $Y=0.74 $X2=0 $Y2=0
cc_149 N_A_27_74#_c_127_n N_Y_c_448_n 0.0119985f $X=1.155 $Y=0.925 $X2=0 $Y2=0
cc_150 N_A_27_74#_c_129_n N_Y_c_448_n 0.0108039f $X=1.24 $Y=1.35 $X2=0 $Y2=0
cc_151 N_A_27_74#_c_130_n N_Y_c_448_n 0.0147728f $X=1.555 $Y=1.515 $X2=0 $Y2=0
cc_152 N_A_27_74#_c_131_n N_Y_c_448_n 0.00248968f $X=1.945 $Y=1.515 $X2=0 $Y2=0
cc_153 N_A_27_74#_c_127_n N_VGND_M1010_d 0.00425898f $X=1.155 $Y=0.925 $X2=-0.19
+ $Y2=-0.245
cc_154 N_A_27_74#_M1002_g N_VGND_c_549_n 0.0032818f $X=1.485 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A_27_74#_c_126_n N_VGND_c_549_n 0.0121972f $X=0.28 $Y=0.68 $X2=0 $Y2=0
cc_156 N_A_27_74#_c_127_n N_VGND_c_549_n 0.0215034f $X=1.155 $Y=0.925 $X2=0
+ $Y2=0
cc_157 N_A_27_74#_c_126_n N_VGND_c_551_n 0.0110419f $X=0.28 $Y=0.68 $X2=0 $Y2=0
cc_158 N_A_27_74#_M1002_g N_VGND_c_552_n 0.00291649f $X=1.485 $Y=0.74 $X2=0
+ $Y2=0
cc_159 N_A_27_74#_M1015_g N_VGND_c_552_n 0.00291649f $X=1.945 $Y=0.74 $X2=0
+ $Y2=0
cc_160 N_A_27_74#_M1002_g N_VGND_c_554_n 0.00364413f $X=1.485 $Y=0.74 $X2=0
+ $Y2=0
cc_161 N_A_27_74#_M1015_g N_VGND_c_554_n 0.00359511f $X=1.945 $Y=0.74 $X2=0
+ $Y2=0
cc_162 N_A_27_74#_c_126_n N_VGND_c_554_n 0.00915013f $X=0.28 $Y=0.68 $X2=0 $Y2=0
cc_163 N_A_27_74#_c_127_n N_VGND_c_554_n 0.0144197f $X=1.155 $Y=0.925 $X2=0
+ $Y2=0
cc_164 N_A_27_74#_c_127_n N_A_225_74#_M1002_d 0.00509711f $X=1.155 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_165 N_A_27_74#_c_129_n N_A_225_74#_M1002_d 0.00174945f $X=1.24 $Y=1.35
+ $X2=-0.19 $Y2=-0.245
cc_166 N_A_27_74#_M1002_g N_A_225_74#_c_605_n 0.0154696f $X=1.485 $Y=0.74 $X2=0
+ $Y2=0
cc_167 N_A_27_74#_M1015_g N_A_225_74#_c_605_n 0.0122685f $X=1.945 $Y=0.74 $X2=0
+ $Y2=0
cc_168 N_A_27_74#_c_127_n N_A_225_74#_c_605_n 0.0148275f $X=1.155 $Y=0.925 $X2=0
+ $Y2=0
cc_169 N_B_M1017_g N_C_M1009_g 0.020343f $X=3.15 $Y=2.4 $X2=0 $Y2=0
cc_170 N_B_c_212_n C 0.00336533f $X=3.15 $Y=1.515 $X2=0 $Y2=0
cc_171 N_B_c_212_n N_C_c_272_n 0.0150236f $X=3.15 $Y=1.515 $X2=0 $Y2=0
cc_172 N_B_M1012_g N_VPWR_c_374_n 0.00263334f $X=2.7 $Y=2.4 $X2=0 $Y2=0
cc_173 N_B_M1017_g N_VPWR_c_375_n 0.00209996f $X=3.15 $Y=2.4 $X2=0 $Y2=0
cc_174 N_B_M1012_g N_VPWR_c_379_n 0.005209f $X=2.7 $Y=2.4 $X2=0 $Y2=0
cc_175 N_B_M1017_g N_VPWR_c_379_n 0.005209f $X=3.15 $Y=2.4 $X2=0 $Y2=0
cc_176 N_B_M1012_g N_VPWR_c_372_n 0.00984248f $X=2.7 $Y=2.4 $X2=0 $Y2=0
cc_177 N_B_M1017_g N_VPWR_c_372_n 0.00982576f $X=3.15 $Y=2.4 $X2=0 $Y2=0
cc_178 N_B_M1012_g N_Y_c_461_n 0.0192154f $X=2.7 $Y=2.4 $X2=0 $Y2=0
cc_179 N_B_c_211_n N_Y_c_461_n 0.0420661f $X=2.425 $Y=1.515 $X2=0 $Y2=0
cc_180 N_B_c_212_n N_Y_c_461_n 0.00171572f $X=3.15 $Y=1.515 $X2=0 $Y2=0
cc_181 N_B_M1001_g N_Y_c_447_n 0.0112328f $X=2.375 $Y=0.74 $X2=0 $Y2=0
cc_182 N_B_M1007_g N_Y_c_447_n 0.0133177f $X=2.965 $Y=0.74 $X2=0 $Y2=0
cc_183 N_B_c_211_n N_Y_c_447_n 0.042165f $X=2.425 $Y=1.515 $X2=0 $Y2=0
cc_184 N_B_c_212_n N_Y_c_447_n 0.0102469f $X=3.15 $Y=1.515 $X2=0 $Y2=0
cc_185 N_B_M1012_g N_Y_c_451_n 0.0166517f $X=2.7 $Y=2.4 $X2=0 $Y2=0
cc_186 N_B_M1017_g N_Y_c_451_n 0.0125032f $X=3.15 $Y=2.4 $X2=0 $Y2=0
cc_187 N_B_M1017_g N_Y_c_478_n 0.00346523f $X=3.15 $Y=2.4 $X2=0 $Y2=0
cc_188 N_B_M1017_g N_Y_c_452_n 5.04845e-19 $X=3.15 $Y=2.4 $X2=0 $Y2=0
cc_189 N_B_M1001_g N_Y_c_448_n 9.39477e-19 $X=2.375 $Y=0.74 $X2=0 $Y2=0
cc_190 N_B_M1012_g N_Y_c_454_n 0.00794088f $X=2.7 $Y=2.4 $X2=0 $Y2=0
cc_191 N_B_M1017_g N_Y_c_454_n 0.0151455f $X=3.15 $Y=2.4 $X2=0 $Y2=0
cc_192 N_B_c_212_n N_Y_c_454_n 0.00316115f $X=3.15 $Y=1.515 $X2=0 $Y2=0
cc_193 N_B_M1001_g Y 7.76767e-19 $X=2.375 $Y=0.74 $X2=0 $Y2=0
cc_194 N_B_M1012_g Y 0.00160954f $X=2.7 $Y=2.4 $X2=0 $Y2=0
cc_195 N_B_M1007_g Y 0.00655125f $X=2.965 $Y=0.74 $X2=0 $Y2=0
cc_196 N_B_M1017_g Y 0.00408417f $X=3.15 $Y=2.4 $X2=0 $Y2=0
cc_197 N_B_c_211_n Y 0.0166916f $X=2.425 $Y=1.515 $X2=0 $Y2=0
cc_198 N_B_c_212_n Y 0.0206134f $X=3.15 $Y=1.515 $X2=0 $Y2=0
cc_199 N_B_M1001_g N_VGND_c_552_n 0.00324657f $X=2.375 $Y=0.74 $X2=0 $Y2=0
cc_200 N_B_M1007_g N_VGND_c_552_n 0.00278271f $X=2.965 $Y=0.74 $X2=0 $Y2=0
cc_201 N_B_M1001_g N_VGND_c_554_n 0.00412223f $X=2.375 $Y=0.74 $X2=0 $Y2=0
cc_202 N_B_M1007_g N_VGND_c_554_n 0.00359811f $X=2.965 $Y=0.74 $X2=0 $Y2=0
cc_203 N_B_M1001_g N_A_225_74#_c_606_n 0.00739353f $X=2.375 $Y=0.74 $X2=0 $Y2=0
cc_204 N_B_M1007_g N_A_225_74#_c_606_n 9.2292e-19 $X=2.965 $Y=0.74 $X2=0 $Y2=0
cc_205 N_B_M1001_g N_A_225_74#_c_607_n 3.34639e-19 $X=2.375 $Y=0.74 $X2=0 $Y2=0
cc_206 N_B_M1007_g N_A_225_74#_c_607_n 0.00257863f $X=2.965 $Y=0.74 $X2=0 $Y2=0
cc_207 N_B_c_212_n N_A_225_74#_c_607_n 7.68732e-19 $X=3.15 $Y=1.515 $X2=0 $Y2=0
cc_208 N_B_M1001_g N_A_225_74#_c_619_n 0.00982687f $X=2.375 $Y=0.74 $X2=0 $Y2=0
cc_209 N_B_M1007_g N_A_225_74#_c_619_n 0.00850118f $X=2.965 $Y=0.74 $X2=0 $Y2=0
cc_210 N_B_M1007_g N_A_490_74#_c_642_n 0.0120769f $X=2.965 $Y=0.74 $X2=0 $Y2=0
cc_211 N_B_M1001_g N_A_490_74#_c_643_n 0.00416113f $X=2.375 $Y=0.74 $X2=0 $Y2=0
cc_212 N_B_M1007_g N_A_719_123#_c_669_n 0.00139553f $X=2.965 $Y=0.74 $X2=0 $Y2=0
cc_213 N_B_M1007_g N_A_719_123#_c_671_n 0.00312109f $X=2.965 $Y=0.74 $X2=0 $Y2=0
cc_214 N_C_M1006_g N_D_M1003_g 0.011802f $X=4.385 $Y=0.79 $X2=0 $Y2=0
cc_215 N_C_M1014_g N_D_c_327_n 0.0281892f $X=4.15 $Y=2.4 $X2=0 $Y2=0
cc_216 C N_D_c_327_n 3.14196e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_217 N_C_c_272_n N_D_c_327_n 0.0153027f $X=4.15 $Y=1.515 $X2=0 $Y2=0
cc_218 C D 0.0279008f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_219 N_C_c_272_n D 0.00810695f $X=4.15 $Y=1.515 $X2=0 $Y2=0
cc_220 N_C_M1009_g N_VPWR_c_375_n 0.00349714f $X=3.7 $Y=2.4 $X2=0 $Y2=0
cc_221 N_C_M1014_g N_VPWR_c_376_n 0.0103864f $X=4.15 $Y=2.4 $X2=0 $Y2=0
cc_222 N_C_M1009_g N_VPWR_c_383_n 0.005209f $X=3.7 $Y=2.4 $X2=0 $Y2=0
cc_223 N_C_M1014_g N_VPWR_c_383_n 0.005209f $X=4.15 $Y=2.4 $X2=0 $Y2=0
cc_224 N_C_M1009_g N_VPWR_c_372_n 0.00982576f $X=3.7 $Y=2.4 $X2=0 $Y2=0
cc_225 N_C_M1014_g N_VPWR_c_372_n 0.00984648f $X=4.15 $Y=2.4 $X2=0 $Y2=0
cc_226 N_C_M1000_g N_Y_c_447_n 5.99596e-19 $X=3.955 $Y=0.79 $X2=0 $Y2=0
cc_227 N_C_M1009_g N_Y_c_451_n 5.04845e-19 $X=3.7 $Y=2.4 $X2=0 $Y2=0
cc_228 N_C_M1009_g N_Y_c_478_n 0.0134293f $X=3.7 $Y=2.4 $X2=0 $Y2=0
cc_229 C N_Y_c_478_n 0.0187969f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_230 N_C_c_272_n N_Y_c_478_n 3.60552e-19 $X=4.15 $Y=1.515 $X2=0 $Y2=0
cc_231 N_C_M1009_g N_Y_c_452_n 0.0120365f $X=3.7 $Y=2.4 $X2=0 $Y2=0
cc_232 N_C_M1014_g N_Y_c_452_n 0.0132828f $X=4.15 $Y=2.4 $X2=0 $Y2=0
cc_233 N_C_M1014_g N_Y_c_497_n 0.0151731f $X=4.15 $Y=2.4 $X2=0 $Y2=0
cc_234 C N_Y_c_497_n 0.00762725f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_235 N_C_c_272_n N_Y_c_497_n 0.00565523f $X=4.15 $Y=1.515 $X2=0 $Y2=0
cc_236 N_C_M1014_g N_Y_c_453_n 8.8199e-19 $X=4.15 $Y=2.4 $X2=0 $Y2=0
cc_237 N_C_M1009_g N_Y_c_501_n 8.84614e-19 $X=3.7 $Y=2.4 $X2=0 $Y2=0
cc_238 N_C_M1014_g N_Y_c_501_n 8.84614e-19 $X=4.15 $Y=2.4 $X2=0 $Y2=0
cc_239 C N_Y_c_501_n 0.0235495f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_240 N_C_c_272_n N_Y_c_501_n 5.48413e-19 $X=4.15 $Y=1.515 $X2=0 $Y2=0
cc_241 N_C_M1009_g Y 0.00112035f $X=3.7 $Y=2.4 $X2=0 $Y2=0
cc_242 N_C_M1000_g Y 0.00367138f $X=3.955 $Y=0.79 $X2=0 $Y2=0
cc_243 C Y 0.0265053f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_244 N_C_c_272_n Y 3.90559e-19 $X=4.15 $Y=1.515 $X2=0 $Y2=0
cc_245 N_C_M1006_g N_VGND_c_550_n 4.25532e-19 $X=4.385 $Y=0.79 $X2=0 $Y2=0
cc_246 N_C_M1000_g N_VGND_c_552_n 8.94875e-19 $X=3.955 $Y=0.79 $X2=0 $Y2=0
cc_247 N_C_M1006_g N_VGND_c_552_n 0.00465842f $X=4.385 $Y=0.79 $X2=0 $Y2=0
cc_248 N_C_M1006_g N_VGND_c_554_n 0.00441603f $X=4.385 $Y=0.79 $X2=0 $Y2=0
cc_249 N_C_M1000_g N_A_490_74#_c_642_n 0.011917f $X=3.955 $Y=0.79 $X2=0 $Y2=0
cc_250 N_C_M1006_g N_A_490_74#_c_642_n 0.00409781f $X=4.385 $Y=0.79 $X2=0 $Y2=0
cc_251 N_C_M1000_g N_A_490_74#_c_648_n 0.00944526f $X=3.955 $Y=0.79 $X2=0 $Y2=0
cc_252 N_C_M1006_g N_A_490_74#_c_648_n 0.00370415f $X=4.385 $Y=0.79 $X2=0 $Y2=0
cc_253 N_C_M1000_g N_A_719_123#_c_670_n 0.0140147f $X=3.955 $Y=0.79 $X2=0 $Y2=0
cc_254 N_C_M1006_g N_A_719_123#_c_670_n 0.0183977f $X=4.385 $Y=0.79 $X2=0 $Y2=0
cc_255 C N_A_719_123#_c_670_n 0.0285914f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_256 N_C_c_272_n N_A_719_123#_c_670_n 0.00452889f $X=4.15 $Y=1.515 $X2=0 $Y2=0
cc_257 C N_A_719_123#_c_671_n 0.0212141f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_258 N_C_c_272_n N_A_719_123#_c_671_n 0.00663695f $X=4.15 $Y=1.515 $X2=0 $Y2=0
cc_259 N_C_M1006_g N_A_719_123#_c_672_n 3.98786e-19 $X=4.385 $Y=0.79 $X2=0 $Y2=0
cc_260 N_D_c_330_n N_VPWR_c_376_n 0.0105406f $X=4.8 $Y=1.77 $X2=0 $Y2=0
cc_261 N_D_M1013_g N_VPWR_c_378_n 0.00525902f $X=5.25 $Y=2.4 $X2=0 $Y2=0
cc_262 D N_VPWR_c_378_n 0.0226229f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_263 N_D_c_330_n N_VPWR_c_384_n 0.005209f $X=4.8 $Y=1.77 $X2=0 $Y2=0
cc_264 N_D_M1013_g N_VPWR_c_384_n 0.005209f $X=5.25 $Y=2.4 $X2=0 $Y2=0
cc_265 N_D_c_330_n N_VPWR_c_372_n 0.009842f $X=4.8 $Y=1.77 $X2=0 $Y2=0
cc_266 N_D_M1013_g N_VPWR_c_372_n 0.00985353f $X=5.25 $Y=2.4 $X2=0 $Y2=0
cc_267 N_D_c_330_n N_Y_c_452_n 8.94462e-19 $X=4.8 $Y=1.77 $X2=0 $Y2=0
cc_268 N_D_c_330_n N_Y_c_497_n 0.0138429f $X=4.8 $Y=1.77 $X2=0 $Y2=0
cc_269 D N_Y_c_497_n 0.0299481f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_270 N_D_c_330_n N_Y_c_512_n 8.84614e-19 $X=4.8 $Y=1.77 $X2=0 $Y2=0
cc_271 N_D_c_327_n N_Y_c_512_n 5.54777e-19 $X=5.25 $Y=1.68 $X2=0 $Y2=0
cc_272 N_D_M1013_g N_Y_c_512_n 0.00242423f $X=5.25 $Y=2.4 $X2=0 $Y2=0
cc_273 D N_Y_c_512_n 0.0235495f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_274 N_D_c_330_n N_Y_c_453_n 0.0129471f $X=4.8 $Y=1.77 $X2=0 $Y2=0
cc_275 N_D_M1013_g N_Y_c_453_n 0.0107114f $X=5.25 $Y=2.4 $X2=0 $Y2=0
cc_276 N_D_M1003_g N_VGND_c_550_n 0.00804216f $X=4.815 $Y=0.79 $X2=0 $Y2=0
cc_277 N_D_M1005_g N_VGND_c_550_n 0.00985076f $X=5.265 $Y=0.79 $X2=0 $Y2=0
cc_278 N_D_M1003_g N_VGND_c_552_n 0.00449979f $X=4.815 $Y=0.79 $X2=0 $Y2=0
cc_279 N_D_M1005_g N_VGND_c_553_n 0.00522181f $X=5.265 $Y=0.79 $X2=0 $Y2=0
cc_280 N_D_M1003_g N_VGND_c_554_n 0.00445136f $X=4.815 $Y=0.79 $X2=0 $Y2=0
cc_281 N_D_M1005_g N_VGND_c_554_n 0.00515793f $X=5.265 $Y=0.79 $X2=0 $Y2=0
cc_282 N_D_M1003_g N_A_490_74#_c_642_n 3.29564e-19 $X=4.815 $Y=0.79 $X2=0 $Y2=0
cc_283 D N_A_719_123#_c_670_n 0.00483207f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_284 N_D_M1003_g N_A_719_123#_c_672_n 3.99083e-19 $X=4.815 $Y=0.79 $X2=0 $Y2=0
cc_285 N_D_M1003_g N_A_719_123#_c_673_n 0.0148218f $X=4.815 $Y=0.79 $X2=0 $Y2=0
cc_286 N_D_c_327_n N_A_719_123#_c_673_n 0.00293928f $X=5.25 $Y=1.68 $X2=0 $Y2=0
cc_287 N_D_M1005_g N_A_719_123#_c_673_n 0.0154779f $X=5.265 $Y=0.79 $X2=0 $Y2=0
cc_288 D N_A_719_123#_c_673_n 0.0544516f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_289 D N_A_719_123#_c_674_n 0.0216404f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_290 N_D_M1005_g N_A_719_123#_c_675_n 0.0015993f $X=5.265 $Y=0.79 $X2=0 $Y2=0
cc_291 D N_A_719_123#_c_676_n 0.017132f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_292 N_VPWR_c_373_n N_Y_c_450_n 0.0315621f $X=1.205 $Y=2.105 $X2=0 $Y2=0
cc_293 N_VPWR_c_374_n N_Y_c_450_n 0.0260414f $X=2.475 $Y=2.455 $X2=0 $Y2=0
cc_294 N_VPWR_c_382_n N_Y_c_450_n 0.0120948f $X=1.995 $Y=3.33 $X2=0 $Y2=0
cc_295 N_VPWR_c_372_n N_Y_c_450_n 0.00994292f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_296 N_VPWR_M1016_s N_Y_c_461_n 0.0134289f $X=1.975 $Y=1.84 $X2=0 $Y2=0
cc_297 N_VPWR_c_374_n N_Y_c_461_n 0.0423878f $X=2.475 $Y=2.455 $X2=0 $Y2=0
cc_298 N_VPWR_c_374_n N_Y_c_451_n 0.0267545f $X=2.475 $Y=2.455 $X2=0 $Y2=0
cc_299 N_VPWR_c_375_n N_Y_c_451_n 0.0266809f $X=3.425 $Y=2.415 $X2=0 $Y2=0
cc_300 N_VPWR_c_379_n N_Y_c_451_n 0.0144623f $X=3.26 $Y=3.33 $X2=0 $Y2=0
cc_301 N_VPWR_c_372_n N_Y_c_451_n 0.0118344f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_302 N_VPWR_M1017_s N_Y_c_478_n 0.0106571f $X=3.24 $Y=1.84 $X2=0 $Y2=0
cc_303 N_VPWR_c_375_n N_Y_c_478_n 0.0208278f $X=3.425 $Y=2.415 $X2=0 $Y2=0
cc_304 N_VPWR_c_375_n N_Y_c_452_n 0.0266809f $X=3.425 $Y=2.415 $X2=0 $Y2=0
cc_305 N_VPWR_c_376_n N_Y_c_452_n 0.0424978f $X=4.485 $Y=2.41 $X2=0 $Y2=0
cc_306 N_VPWR_c_383_n N_Y_c_452_n 0.0144623f $X=4.32 $Y=3.33 $X2=0 $Y2=0
cc_307 N_VPWR_c_372_n N_Y_c_452_n 0.0118344f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_308 N_VPWR_M1014_s N_Y_c_497_n 0.00980226f $X=4.24 $Y=1.84 $X2=0 $Y2=0
cc_309 N_VPWR_c_376_n N_Y_c_497_n 0.0266856f $X=4.485 $Y=2.41 $X2=0 $Y2=0
cc_310 N_VPWR_c_376_n N_Y_c_453_n 0.0455581f $X=4.485 $Y=2.41 $X2=0 $Y2=0
cc_311 N_VPWR_c_378_n N_Y_c_453_n 0.0330049f $X=5.475 $Y=2.115 $X2=0 $Y2=0
cc_312 N_VPWR_c_384_n N_Y_c_453_n 0.0144623f $X=5.36 $Y=3.33 $X2=0 $Y2=0
cc_313 N_VPWR_c_372_n N_Y_c_453_n 0.0118344f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_314 N_Y_c_447_n N_A_225_74#_M1015_d 0.00176461f $X=3.005 $Y=1.095 $X2=0 $Y2=0
cc_315 N_Y_c_447_n N_A_225_74#_M1007_d 0.00300606f $X=3.005 $Y=1.095 $X2=0 $Y2=0
cc_316 N_Y_M1002_s N_A_225_74#_c_605_n 0.00211578f $X=1.56 $Y=0.37 $X2=0 $Y2=0
cc_317 N_Y_c_447_n N_A_225_74#_c_605_n 0.00459468f $X=3.005 $Y=1.095 $X2=0 $Y2=0
cc_318 N_Y_c_448_n N_A_225_74#_c_605_n 0.0187497f $X=1.715 $Y=0.965 $X2=0 $Y2=0
cc_319 N_Y_c_447_n N_A_225_74#_c_606_n 0.0149311f $X=3.005 $Y=1.095 $X2=0 $Y2=0
cc_320 N_Y_c_447_n N_A_225_74#_c_619_n 0.0540678f $X=3.005 $Y=1.095 $X2=0 $Y2=0
cc_321 N_Y_c_447_n N_A_490_74#_M1001_s 0.00391227f $X=3.005 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_322 N_Y_c_447_n N_A_719_123#_c_671_n 0.00962672f $X=3.005 $Y=1.095 $X2=0
+ $Y2=0
cc_323 N_VGND_c_549_n N_A_225_74#_c_605_n 0.0198879f $X=0.71 $Y=0.55 $X2=0 $Y2=0
cc_324 N_VGND_c_552_n N_A_225_74#_c_605_n 0.039681f $X=4.865 $Y=0 $X2=0 $Y2=0
cc_325 N_VGND_c_554_n N_A_225_74#_c_605_n 0.0333579f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_326 N_VGND_c_552_n N_A_225_74#_c_606_n 0.0107387f $X=4.865 $Y=0 $X2=0 $Y2=0
cc_327 N_VGND_c_554_n N_A_225_74#_c_606_n 0.00894442f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_328 N_VGND_c_552_n N_A_225_74#_c_619_n 0.00237563f $X=4.865 $Y=0 $X2=0 $Y2=0
cc_329 N_VGND_c_554_n N_A_225_74#_c_619_n 0.00539332f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_330 N_VGND_c_550_n N_A_490_74#_c_642_n 0.00485382f $X=5.03 $Y=0.58 $X2=0
+ $Y2=0
cc_331 N_VGND_c_552_n N_A_490_74#_c_642_n 0.0231371f $X=4.865 $Y=0 $X2=0 $Y2=0
cc_332 N_VGND_c_554_n N_A_490_74#_c_642_n 0.0127322f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_333 N_VGND_c_552_n N_A_490_74#_c_643_n 0.0966814f $X=4.865 $Y=0 $X2=0 $Y2=0
cc_334 N_VGND_c_554_n N_A_490_74#_c_643_n 0.0558053f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_335 N_VGND_c_550_n N_A_719_123#_c_672_n 0.0142351f $X=5.03 $Y=0.58 $X2=0
+ $Y2=0
cc_336 N_VGND_c_552_n N_A_719_123#_c_672_n 0.00698151f $X=4.865 $Y=0 $X2=0 $Y2=0
cc_337 N_VGND_c_554_n N_A_719_123#_c_672_n 0.00673015f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_338 N_VGND_M1003_s N_A_719_123#_c_673_n 0.00200085f $X=4.89 $Y=0.42 $X2=0
+ $Y2=0
cc_339 N_VGND_c_550_n N_A_719_123#_c_673_n 0.017643f $X=5.03 $Y=0.58 $X2=0 $Y2=0
cc_340 N_VGND_c_550_n N_A_719_123#_c_675_n 0.0125364f $X=5.03 $Y=0.58 $X2=0
+ $Y2=0
cc_341 N_VGND_c_553_n N_A_719_123#_c_675_n 0.00920966f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_342 N_VGND_c_554_n N_A_719_123#_c_675_n 0.00887807f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_343 N_A_225_74#_c_619_n N_A_490_74#_M1001_s 0.00727678f $X=3.015 $Y=0.717
+ $X2=-0.19 $Y2=-0.245
cc_344 N_A_225_74#_M1007_d N_A_490_74#_c_642_n 0.00226585f $X=3.04 $Y=0.37 $X2=0
+ $Y2=0
cc_345 N_A_225_74#_c_607_n N_A_490_74#_c_642_n 0.0191024f $X=3.18 $Y=0.715 $X2=0
+ $Y2=0
cc_346 N_A_225_74#_c_619_n N_A_490_74#_c_642_n 0.00570513f $X=3.015 $Y=0.717
+ $X2=0 $Y2=0
cc_347 N_A_225_74#_c_606_n N_A_490_74#_c_643_n 0.00599132f $X=2.2 $Y=0.49 $X2=0
+ $Y2=0
cc_348 N_A_225_74#_c_619_n N_A_490_74#_c_643_n 0.0232532f $X=3.015 $Y=0.717
+ $X2=0 $Y2=0
cc_349 N_A_225_74#_c_607_n N_A_719_123#_c_669_n 0.0167582f $X=3.18 $Y=0.715
+ $X2=0 $Y2=0
cc_350 N_A_490_74#_c_642_n N_A_719_123#_M1000_d 0.00206713f $X=4.005 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_351 N_A_490_74#_c_642_n N_A_719_123#_c_669_n 0.0187376f $X=4.005 $Y=0.34
+ $X2=0 $Y2=0
cc_352 N_A_490_74#_M1000_s N_A_719_123#_c_670_n 0.00178571f $X=4.03 $Y=0.42
+ $X2=0 $Y2=0
cc_353 N_A_490_74#_c_642_n N_A_719_123#_c_670_n 0.00356278f $X=4.005 $Y=0.34
+ $X2=0 $Y2=0
cc_354 N_A_490_74#_c_648_n N_A_719_123#_c_670_n 0.0171301f $X=4.17 $Y=0.58 $X2=0
+ $Y2=0
cc_355 N_A_490_74#_c_642_n N_A_719_123#_c_672_n 0.00178319f $X=4.005 $Y=0.34
+ $X2=0 $Y2=0

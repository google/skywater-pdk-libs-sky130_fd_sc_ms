* File: sky130_fd_sc_ms__a41oi_1.pex.spice
* Created: Fri Aug 28 17:09:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A41OI_1%B1 3 7 9 13 16
r26 15 16 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.465
+ $X2=0.505 $Y2=1.465
r27 12 15 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.27 $Y=1.465
+ $X2=0.495 $Y2=1.465
r28 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r29 9 13 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.27 $Y=1.665 $X2=0.27
+ $Y2=1.465
r30 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.465
r31 5 7 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.74
r32 1 16 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=1.465
r33 1 3 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A41OI_1%A4 3 7 9 15 16
r38 14 16 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=1.17 $Y=1.515
+ $X2=1.31 $Y2=1.515
r39 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.515 $X2=1.17 $Y2=1.515
r40 11 14 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.515
+ $X2=1.17 $Y2=1.515
r41 9 15 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.17 $Y=1.665
+ $X2=1.17 $Y2=1.515
r42 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.31 $Y=1.35
+ $X2=1.31 $Y2=1.515
r43 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.31 $Y=1.35 $X2=1.31
+ $Y2=0.74
r44 1 11 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.68
+ $X2=1.005 $Y2=1.515
r45 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.005 $Y=1.68
+ $X2=1.005 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A41OI_1%A3 3 7 9 12 13
r35 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=1.515
+ $X2=1.79 $Y2=1.68
r36 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=1.515
+ $X2=1.79 $Y2=1.35
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.79
+ $Y=1.515 $X2=1.79 $Y2=1.515
r38 9 13 4.43247 $w=3.88e-07 $l=1.5e-07 $layer=LI1_cond $X=1.76 $Y=1.665
+ $X2=1.76 $Y2=1.515
r39 7 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.845 $Y=2.4
+ $X2=1.845 $Y2=1.68
r40 3 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.7 $Y=0.74 $X2=1.7
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__A41OI_1%A2 3 7 9 12
c35 7 0 6.15358e-20 $X=2.295 $Y=2.4
r36 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.36 $Y=1.515
+ $X2=2.36 $Y2=1.68
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.36 $Y=1.515
+ $X2=2.36 $Y2=1.35
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.36
+ $Y=1.515 $X2=2.36 $Y2=1.515
r39 9 13 7.50428 $w=4.28e-07 $l=2.8e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.36 $Y2=1.565
r40 7 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.295 $Y=2.4
+ $X2=2.295 $Y2=1.68
r41 3 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.27 $Y=0.74 $X2=2.27
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__A41OI_1%A1 3 7 9 15 16
c27 16 0 6.15358e-20 $X=3.09 $Y=1.465
r28 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.465 $X2=3.09 $Y2=1.465
r29 13 15 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=2.855 $Y=1.465
+ $X2=3.09 $Y2=1.465
r30 11 13 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.84 $Y=1.465
+ $X2=2.855 $Y2=1.465
r31 9 16 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.09 $Y=1.665 $X2=3.09
+ $Y2=1.465
r32 5 13 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.855 $Y=1.63
+ $X2=2.855 $Y2=1.465
r33 5 7 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=2.855 $Y=1.63
+ $X2=2.855 $Y2=2.4
r34 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=1.3 $X2=2.84
+ $Y2=1.465
r35 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.84 $Y=1.3 $X2=2.84
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A41OI_1%Y 1 2 3 12 16 18 19 22 32 34
r54 32 34 32.8196 $w=2.28e-07 $l=6.55e-07 $layer=LI1_cond $X=0.72 $Y=1.95
+ $X2=0.72 $Y2=1.295
r55 29 32 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=0.28 $Y=2.035
+ $X2=0.72 $Y2=2.035
r56 27 34 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.72 $Y=1.13
+ $X2=0.72 $Y2=1.295
r57 20 22 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.055 $Y=0.96
+ $X2=3.055 $Y2=0.515
r58 19 27 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.835 $Y=1.045
+ $X2=0.72 $Y2=1.045
r59 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.89 $Y=1.045
+ $X2=3.055 $Y2=0.96
r60 18 19 134.07 $w=1.68e-07 $l=2.055e-06 $layer=LI1_cond $X=2.89 $Y=1.045
+ $X2=0.835 $Y2=1.045
r61 16 29 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.28 $Y=2.815
+ $X2=0.28 $Y2=2.12
r62 10 27 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=0.28 $Y=1.045
+ $X2=0.72 $Y2=1.045
r63 10 12 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.28 $Y=0.96
+ $X2=0.28 $Y2=0.515
r64 3 29 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.035
r65 3 16 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r66 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.915
+ $Y=0.37 $X2=3.055 $Y2=0.515
r67 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A41OI_1%A_119_368# 1 2 3 12 13 16 18 21
r39 16 23 3.46012 $w=3.3e-07 $l=1.7e-07 $layer=LI1_cond $X=3.08 $Y=2.29 $X2=3.08
+ $Y2=2.12
r40 16 18 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=3.08 $Y=2.29
+ $X2=3.08 $Y2=2.815
r41 13 21 18.5174 $w=3.4e-07 $l=5.73738e-07 $layer=LI1_cond $X=1.275 $Y=2.12
+ $X2=0.78 $Y2=2.29
r42 13 15 26.9468 $w=3.38e-07 $l=7.95e-07 $layer=LI1_cond $X=1.275 $Y=2.12
+ $X2=2.07 $Y2=2.12
r43 12 23 3.35835 $w=3.4e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=2.12
+ $X2=3.08 $Y2=2.12
r44 12 15 28.6416 $w=3.38e-07 $l=8.45e-07 $layer=LI1_cond $X=2.915 $Y=2.12
+ $X2=2.07 $Y2=2.12
r45 3 23 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=2.945
+ $Y=1.84 $X2=3.08 $Y2=2.035
r46 3 18 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.945
+ $Y=1.84 $X2=3.08 $Y2=2.815
r47 2 15 600 $w=1.7e-07 $l=3.40881e-07 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=1.84 $X2=2.07 $Y2=2.12
r48 1 21 300 $w=1.7e-07 $l=6.20645e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.78 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_MS__A41OI_1%VPWR 1 2 9 11 13 18 25 26 31 34
r37 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 29 31 12.18 $w=6.11e-07 $l=6.1e-07 $layer=LI1_cond $X=1.45 $Y=2.72 $X2=1.45
+ $Y2=3.33
r39 26 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 23 34 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.745 $Y=3.33
+ $X2=2.575 $Y2=3.33
r42 23 25 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.745 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 22 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 19 31 8.43407 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=1.45 $Y2=3.33
r46 19 21 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 18 34 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.405 $Y=3.33
+ $X2=2.575 $Y2=3.33
r48 18 21 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.405 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 15 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 13 31 8.43407 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=1.45 $Y2=3.33
r51 13 15 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 11 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 11 16 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 11 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 7 34 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.575 $Y=3.245
+ $X2=2.575 $Y2=3.33
r56 7 9 21.0151 $w=3.38e-07 $l=6.2e-07 $layer=LI1_cond $X=2.575 $Y=3.245
+ $X2=2.575 $Y2=2.625
r57 2 9 600 $w=1.7e-07 $l=8.74857e-07 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=1.84 $X2=2.575 $Y2=2.625
r58 1 29 300 $w=1.7e-07 $l=1.11194e-06 $layer=licon1_PDIFF $count=2 $X=1.095
+ $Y=1.84 $X2=1.62 $Y2=2.72
.ends

.subckt PM_SKY130_FD_SC_MS__A41OI_1%VGND 1 4 6 13 14
r22 19 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r23 13 14 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r24 11 13 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=1.26 $Y=0 $X2=3.12
+ $Y2=0
r25 9 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r26 8 9 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r27 6 23 9.55008 $w=6.43e-07 $l=5.15e-07 $layer=LI1_cond $X=0.937 $Y=0 $X2=0.937
+ $Y2=0.515
r28 6 11 8.78548 $w=1.7e-07 $l=3.23e-07 $layer=LI1_cond $X=0.937 $Y=0 $X2=1.26
+ $Y2=0
r29 6 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r30 6 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r31 6 8 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r32 4 14 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r33 4 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r34 1 23 91 $w=1.7e-07 $l=5.93085e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=1.095 $Y2=0.515
.ends


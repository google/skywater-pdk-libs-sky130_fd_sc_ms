* File: sky130_fd_sc_ms__nand4b_4.spice
* Created: Wed Sep  2 12:14:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nand4b_4.pex.spice"
.subckt sky130_fd_sc_ms__nand4b_4  VNB VPB A_N B C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1023 N_VGND_M1023_d N_A_N_M1023_g N_A_27_158#_M1023_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.19515 AS=0.1962 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_A_225_74#_M1005_d N_A_27_158#_M1005_g N_Y_M1005_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1962 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75003.2 A=0.111 P=1.78 MULT=1
MM1011 N_A_225_74#_M1011_d N_A_27_158#_M1011_g N_Y_M1005_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75002.8 A=0.111 P=1.78 MULT=1
MM1024 N_A_225_74#_M1011_d N_A_27_158#_M1024_g N_Y_M1024_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75002.3 A=0.111 P=1.78 MULT=1
MM1025 N_A_225_74#_M1025_d N_A_27_158#_M1025_g N_Y_M1024_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75001.9 A=0.111 P=1.78 MULT=1
MM1003 N_A_225_74#_M1025_d N_B_M1003_g N_A_656_74#_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.9 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1009 N_A_225_74#_M1009_d N_B_M1009_g N_A_656_74#_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.3 SB=75001 A=0.111 P=1.78 MULT=1
MM1019 N_A_225_74#_M1009_d N_B_M1019_g N_A_656_74#_M1019_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.8 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1021 N_A_225_74#_M1021_d N_B_M1021_g N_A_656_74#_M1019_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.19515 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75003.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_656_74#_M1000_d N_C_M1000_g N_A_1025_158#_M1000_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1962 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75003.3 A=0.111 P=1.78 MULT=1
MM1008 N_A_656_74#_M1000_d N_C_M1008_g N_A_1025_158#_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75002.9 A=0.111 P=1.78 MULT=1
MM1013 N_A_656_74#_M1013_d N_C_M1013_g N_A_1025_158#_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.10915 AS=0.1036 PD=1.035 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1026 N_A_656_74#_M1013_d N_C_M1026_g N_A_1025_158#_M1026_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.10915 AS=0.1036 PD=1.035 PS=1.02 NRD=2.424 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75002 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_D_M1001_g N_A_1025_158#_M1026_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1001_d N_D_M1007_g N_A_1025_158#_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.4
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1014_d N_D_M1014_g N_A_1025_158#_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.14615 AS=0.1036 PD=1.135 PS=1.02 NRD=3.24 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1014_d N_D_M1015_g N_A_1025_158#_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.14615 AS=0.2109 PD=1.135 PS=2.05 NRD=15.396 NRS=0 M=1 R=4.93333
+ SA=75003.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1018 N_A_27_158#_M1018_d N_A_N_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.2772 PD=1.11 PS=2.34 NRD=0 NRS=10.5395 M=1 R=4.66667 SA=90000.2
+ SB=90007.9 A=0.1512 P=2.04 MULT=1
MM1022 N_A_27_158#_M1018_d N_A_N_M1022_g N_VPWR_M1022_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.1614 PD=1.11 PS=1.26429 NRD=0 NRS=18.7544 M=1 R=4.66667
+ SA=90000.7 SB=90007.4 A=0.1512 P=2.04 MULT=1
MM1002 N_Y_M1002_d N_A_27_158#_M1002_g N_VPWR_M1022_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3808 AS=0.2152 PD=1.8 PS=1.68571 NRD=0 NRS=0 M=1 R=6.22222 SA=90001
+ SB=90006.9 A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1002_d N_A_27_158#_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3808 AS=0.7168 PD=1.8 PS=2.4 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.8
+ SB=90006 A=0.2016 P=2.6 MULT=1
MM1016 N_Y_M1016_d N_B_M1016_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.7168 PD=1.39 PS=2.4 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.3 SB=90004.6
+ A=0.2016 P=2.6 MULT=1
MM1020 N_Y_M1016_d N_B_M1020_g N_VPWR_M1020_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.5964 PD=1.39 PS=2.185 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.7 SB=90004.1
+ A=0.2016 P=2.6 MULT=1
MM1012 N_VPWR_M1020_s N_C_M1012_g N_Y_M1012_s VPB PSHORT L=0.18 W=1.12 AD=0.5964
+ AS=0.364 PD=2.185 PS=1.77 NRD=0 NRS=0 M=1 R=6.22222 SA=90005 SB=90002.9
+ A=0.2016 P=2.6 MULT=1
MM1017 N_VPWR_M1017_d N_C_M1017_g N_Y_M1012_s VPB PSHORT L=0.18 W=1.12 AD=0.6384
+ AS=0.364 PD=2.26 PS=1.77 NRD=0 NRS=0 M=1 R=6.22222 SA=90005.8 SB=90002
+ A=0.2016 P=2.6 MULT=1
MM1006 N_Y_M1006_d N_D_M1006_g N_VPWR_M1017_d VPB PSHORT L=0.18 W=1.12 AD=0.1624
+ AS=0.6384 PD=1.41 PS=2.26 NRD=2.6201 NRS=0 M=1 R=6.22222 SA=90007.1 SB=90000.7
+ A=0.2016 P=2.6 MULT=1
MM1010 N_Y_M1006_d N_D_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.18 W=1.12 AD=0.1624
+ AS=0.3696 PD=1.41 PS=2.9 NRD=0 NRS=0 M=1 R=6.22222 SA=90007.6 SB=90000.2
+ A=0.2016 P=2.6 MULT=1
DX27_noxref VNB VPB NWDIODE A=17.67 P=22.72
c_75 VNB 0 7.64129e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__nand4b_4.pxi.spice"
*
.ends
*
*

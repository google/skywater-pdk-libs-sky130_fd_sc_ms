* File: sky130_fd_sc_ms__or4b_1.pex.spice
* Created: Wed Sep  2 12:29:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__OR4B_1%D_N 3 5 7 9 13
r34 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.405
+ $Y=1.615 $X2=0.405 $Y2=1.615
r35 9 13 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.405 $Y2=1.615
r36 5 12 34.0194 $w=3.43e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.51 $Y=1.78
+ $X2=0.42 $Y2=1.615
r37 5 7 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=0.51 $Y=1.78 $X2=0.51
+ $Y2=2.54
r38 1 12 38.7084 $w=3.43e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.42 $Y2=1.615
r39 1 3 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.495 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_1%A_27_74# 1 2 9 11 13 15 18 22 24 25 26 27 29
+ 31 34
r69 34 35 36.5941 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=0.975 $Y=1.69
+ $X2=0.975 $Y2=1.58
r70 32 34 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=0.975 $Y=1.745
+ $X2=0.975 $Y2=1.69
r71 31 33 13.2509 $w=2.67e-07 $l=2.9e-07 $layer=LI1_cond $X=0.975 $Y=1.745
+ $X2=0.975 $Y2=2.035
r72 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.745 $X2=0.975 $Y2=1.745
r73 29 31 9.14344 $w=2.67e-07 $l=2.0106e-07 $layer=LI1_cond $X=0.895 $Y=1.58
+ $X2=0.975 $Y2=1.745
r74 28 29 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.895 $Y=1.28
+ $X2=0.895 $Y2=1.58
r75 26 33 3.37873 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.81 $Y=2.035
+ $X2=0.975 $Y2=2.035
r76 26 27 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.81 $Y=2.035
+ $X2=0.45 $Y2=2.035
r77 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.81 $Y=1.195
+ $X2=0.895 $Y2=1.28
r78 24 25 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.81 $Y=1.195
+ $X2=0.445 $Y2=1.195
r79 20 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.285 $Y=2.12
+ $X2=0.45 $Y2=2.035
r80 20 22 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.285 $Y=2.12
+ $X2=0.285 $Y2=2.265
r81 16 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.11
+ $X2=0.445 $Y2=1.195
r82 16 18 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.28 $Y=1.11
+ $X2=0.28 $Y2=0.645
r83 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.705 $Y=1.765
+ $X2=1.705 $Y2=2.34
r84 12 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=1.69
+ $X2=0.975 $Y2=1.69
r85 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.615 $Y=1.69
+ $X2=1.705 $Y2=1.765
r86 11 12 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.615 $Y=1.69
+ $X2=1.14 $Y2=1.69
r87 9 35 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=1.065 $Y=0.645
+ $X2=1.065 $Y2=1.58
r88 2 22 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.14
+ $Y=2.12 $X2=0.285 $Y2=2.265
r89 1 18 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_1%C 3 7 8 9 13 14 15
r33 13 16 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.05 $Y=1.21
+ $X2=2.05 $Y2=1.375
r34 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.05 $Y=1.21
+ $X2=2.05 $Y2=1.045
r35 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.05
+ $Y=1.21 $X2=2.05 $Y2=1.21
r36 8 9 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.08 $Y=1.295 $X2=2.08
+ $Y2=1.665
r37 8 14 2.51173 $w=3.88e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=1.295
+ $X2=2.08 $Y2=1.21
r38 7 15 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.14 $Y=0.645 $X2=2.14
+ $Y2=1.045
r39 3 16 375.105 $w=1.8e-07 $l=9.65e-07 $layer=POLY_cond $X=2.125 $Y=2.34
+ $X2=2.125 $Y2=1.375
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_1%B 3 7 9 10 14
r33 14 17 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.62 $Y=1.345
+ $X2=2.62 $Y2=1.51
r34 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.62 $Y=1.345
+ $X2=2.62 $Y2=1.18
r35 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.62 $Y=1.295
+ $X2=2.62 $Y2=1.665
r36 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.62
+ $Y=1.345 $X2=2.62 $Y2=1.345
r37 7 16 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.71 $Y=0.645
+ $X2=2.71 $Y2=1.18
r38 3 17 322.629 $w=1.8e-07 $l=8.3e-07 $layer=POLY_cond $X=2.545 $Y=2.34
+ $X2=2.545 $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_1%A 3 7 9 12 13
c43 7 0 7.34258e-20 $X=3.14 $Y=0.645
c44 3 0 1.18964e-19 $X=3.085 $Y=2.34
r45 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.16 $Y=1.515
+ $X2=3.16 $Y2=1.68
r46 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.16 $Y=1.515
+ $X2=3.16 $Y2=1.35
r47 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.16
+ $Y=1.515 $X2=3.16 $Y2=1.515
r48 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.16 $Y=1.665
+ $X2=3.16 $Y2=1.515
r49 7 14 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=3.14 $Y=0.645 $X2=3.14
+ $Y2=1.35
r50 3 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.085 $Y=2.34
+ $X2=3.085 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_1%A_228_74# 1 2 3 12 16 18 19 22 26 28 30 33 35
+ 36 40 45
r107 45 48 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=1.465
+ $X2=3.73 $Y2=1.63
r108 45 47 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=1.465
+ $X2=3.73 $Y2=1.3
r109 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.73
+ $Y=1.465 $X2=3.73 $Y2=1.465
r110 35 44 9.00568 $w=2.92e-07 $l=2.14942e-07 $layer=LI1_cond $X=3.58 $Y=1.63
+ $X2=3.695 $Y2=1.465
r111 35 36 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.58 $Y=1.63
+ $X2=3.58 $Y2=1.95
r112 34 41 3.08766 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.125 $Y=1.095
+ $X2=2.955 $Y2=1.095
r113 33 44 15.4589 $w=2.92e-07 $l=4.59238e-07 $layer=LI1_cond $X=3.495 $Y=1.095
+ $X2=3.695 $Y2=1.465
r114 33 34 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.495 $Y=1.095
+ $X2=3.125 $Y2=1.095
r115 30 41 12.4049 $w=3.65e-07 $l=3.43439e-07 $layer=LI1_cond $X=2.942 $Y=0.758
+ $X2=2.955 $Y2=1.095
r116 30 32 3.77699 $w=3.65e-07 $l=1.13e-07 $layer=LI1_cond $X=2.942 $Y=0.758
+ $X2=2.942 $Y2=0.645
r117 29 40 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.645 $Y=2.035
+ $X2=1.48 $Y2=2.035
r118 28 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.495 $Y=2.035
+ $X2=3.58 $Y2=1.95
r119 28 29 120.695 $w=1.68e-07 $l=1.85e-06 $layer=LI1_cond $X=3.495 $Y=2.035
+ $X2=1.645 $Y2=2.035
r120 24 38 3.40825 $w=3.3e-07 $l=2.65e-07 $layer=LI1_cond $X=1.645 $Y=0.71
+ $X2=1.38 $Y2=0.71
r121 24 26 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.645 $Y=0.71
+ $X2=1.925 $Y2=0.71
r122 20 40 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.48 $Y=2.12
+ $X2=1.48 $Y2=2.035
r123 20 22 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=1.48 $Y=2.12
+ $X2=1.48 $Y2=2.695
r124 19 40 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.48 $Y=1.95
+ $X2=1.48 $Y2=2.035
r125 18 38 3.40825 $w=3.3e-07 $l=2.09105e-07 $layer=LI1_cond $X=1.48 $Y=0.875
+ $X2=1.38 $Y2=0.71
r126 18 19 37.5417 $w=3.28e-07 $l=1.075e-06 $layer=LI1_cond $X=1.48 $Y=0.875
+ $X2=1.48 $Y2=1.95
r127 16 47 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.785 $Y=0.74
+ $X2=3.785 $Y2=1.3
r128 12 48 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=3.775 $Y=2.4
+ $X2=3.775 $Y2=1.63
r129 3 40 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.335
+ $Y=1.84 $X2=1.48 $Y2=1.985
r130 3 22 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.335
+ $Y=1.84 $X2=1.48 $Y2=2.695
r131 2 32 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.785
+ $Y=0.37 $X2=2.925 $Y2=0.645
r132 1 38 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=1.14
+ $Y=0.37 $X2=1.28 $Y2=0.71
r133 1 26 182 $w=1.7e-07 $l=9.39747e-07 $layer=licon1_NDIFF $count=1 $X=1.14
+ $Y=0.37 $X2=1.925 $Y2=0.71
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_1%VPWR 1 2 9 13 18 19 20 22 35 36 39
r42 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r44 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r45 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 30 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 29 32 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r49 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=3.33
+ $X2=0.785 $Y2=3.33
r50 27 29 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.95 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=3.33
+ $X2=0.785 $Y2=3.33
r54 22 24 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.62 $Y=3.33
+ $X2=0.24 $Y2=3.33
r55 20 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 20 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r57 18 32 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.335 $Y=3.33
+ $X2=3.12 $Y2=3.33
r58 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.335 $Y=3.33
+ $X2=3.5 $Y2=3.33
r59 17 35 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.665 $Y=3.33
+ $X2=4.08 $Y2=3.33
r60 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.665 $Y=3.33
+ $X2=3.5 $Y2=3.33
r61 13 16 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.5 $Y=2.455 $X2=3.5
+ $Y2=2.815
r62 11 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.5 $Y=3.245 $X2=3.5
+ $Y2=3.33
r63 11 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.5 $Y=3.245 $X2=3.5
+ $Y2=2.815
r64 7 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=3.245
+ $X2=0.785 $Y2=3.33
r65 7 9 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=0.785 $Y=3.245
+ $X2=0.785 $Y2=2.455
r66 2 16 600 $w=1.7e-07 $l=1.12583e-06 $layer=licon1_PDIFF $count=1 $X=3.175
+ $Y=1.84 $X2=3.5 $Y2=2.815
r67 2 13 600 $w=1.7e-07 $l=7.60329e-07 $layer=licon1_PDIFF $count=1 $X=3.175
+ $Y=1.84 $X2=3.5 $Y2=2.455
r68 1 9 300 $w=1.7e-07 $l=4.17373e-07 $layer=licon1_PDIFF $count=2 $X=0.6
+ $Y=2.12 $X2=0.785 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_1%X 1 2 9 13 14 15 16 23 33
c28 14 0 1.18964e-19 $X=3.995 $Y=1.95
c29 13 0 7.34258e-20 $X=4.035 $Y=1.13
r30 21 23 0.432166 $w=3.98e-07 $l=1.5e-08 $layer=LI1_cond $X=4.035 $Y=2.02
+ $X2=4.035 $Y2=2.035
r31 15 16 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=4.035 $Y=2.405
+ $X2=4.035 $Y2=2.775
r32 14 21 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=4.035 $Y=1.985
+ $X2=4.035 $Y2=2.02
r33 14 33 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=4.035 $Y=1.985
+ $X2=4.035 $Y2=1.82
r34 14 15 9.65171 $w=3.98e-07 $l=3.35e-07 $layer=LI1_cond $X=4.035 $Y=2.07
+ $X2=4.035 $Y2=2.405
r35 14 23 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=4.035 $Y=2.07
+ $X2=4.035 $Y2=2.035
r36 13 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.15 $Y=1.13 $X2=4.15
+ $Y2=1.82
r37 7 13 9.656 $w=3.98e-07 $l=2e-07 $layer=LI1_cond $X=4.035 $Y=0.93 $X2=4.035
+ $Y2=1.13
r38 7 9 11.9566 $w=3.98e-07 $l=4.15e-07 $layer=LI1_cond $X=4.035 $Y=0.93
+ $X2=4.035 $Y2=0.515
r39 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.865
+ $Y=1.84 $X2=4 $Y2=1.985
r40 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.865
+ $Y=1.84 $X2=4 $Y2=2.815
r41 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.86
+ $Y=0.37 $X2=4 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__OR4B_1%VGND 1 2 3 12 16 20 23 24 26 27 28 30 46 47
+ 50
r54 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r55 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r56 44 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r57 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r58 38 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r59 37 40 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r60 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r61 35 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.78
+ $Y2=0
r62 35 37 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r63 33 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r64 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r65 30 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.78
+ $Y2=0
r66 30 32 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.24
+ $Y2=0
r67 28 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r68 28 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r69 28 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r70 26 43 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.295 $Y=0 $X2=3.12
+ $Y2=0
r71 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=0 $X2=3.46
+ $Y2=0
r72 25 46 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.625 $Y=0 $X2=4.08
+ $Y2=0
r73 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.625 $Y=0 $X2=3.46
+ $Y2=0
r74 23 40 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.26 $Y=0 $X2=2.16
+ $Y2=0
r75 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=0 $X2=2.425
+ $Y2=0
r76 22 43 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.59 $Y=0 $X2=3.12
+ $Y2=0
r77 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.59 $Y=0 $X2=2.425
+ $Y2=0
r78 18 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=0.085
+ $X2=3.46 $Y2=0
r79 18 20 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=3.46 $Y=0.085
+ $X2=3.46 $Y2=0.595
r80 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=0.085
+ $X2=2.425 $Y2=0
r81 14 16 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=2.425 $Y=0.085
+ $X2=2.425 $Y2=0.61
r82 10 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r83 10 12 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.645
r84 3 20 182 $w=1.7e-07 $l=3.39338e-07 $layer=licon1_NDIFF $count=1 $X=3.215
+ $Y=0.37 $X2=3.46 $Y2=0.595
r85 2 16 182 $w=1.7e-07 $l=3.28634e-07 $layer=licon1_NDIFF $count=1 $X=2.215
+ $Y=0.37 $X2=2.425 $Y2=0.61
r86 1 12 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.645
.ends


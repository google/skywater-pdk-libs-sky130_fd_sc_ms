* File: sky130_fd_sc_ms__nor3_2.spice
* Created: Wed Sep  2 12:16:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nor3_2.pex.spice"
.subckt sky130_fd_sc_ms__nor3_2  VNB VPB C B A Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_C_M1006_g N_Y_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.32745 AS=0.2109 PD=1.625 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.8 A=0.111 P=1.78 MULT=1
MM1008 N_Y_M1008_d N_B_M1008_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.74 AD=0.1295
+ AS=0.32745 PD=1.09 PS=1.625 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75000.8 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g N_Y_M1008_d VNB NLOWVT L=0.15 W=0.74 AD=0.2627
+ AS=0.1295 PD=2.19 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.7 SB=75000.3
+ A=0.111 P=1.78 MULT=1
MM1000 N_A_27_368#_M1000_d N_C_M1000_g N_Y_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.1792 PD=2.8 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.2
+ SB=90002.5 A=0.2016 P=2.6 MULT=1
MM1002 N_A_27_368#_M1002_d N_C_M1002_g N_Y_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.7
+ SB=90002 A=0.2016 P=2.6 MULT=1
MM1001 N_A_309_368#_M1001_d N_B_M1001_g N_A_27_368#_M1002_d VPB PSHORT L=0.18
+ W=1.12 AD=0.168 AS=0.1512 PD=1.42 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1003 N_A_309_368#_M1001_d N_A_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.168 AS=0.1624 PD=1.42 PS=1.41 NRD=4.3931 NRS=2.6201 M=1 R=6.22222
+ SA=90001.6 SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1005 N_A_309_368#_M1005_d N_A_M1005_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1624 PD=1.39 PS=1.41 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.1
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1004 N_A_309_368#_M1005_d N_B_M1004_g N_A_27_368#_M1004_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX9_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__nor3_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__nor4b_4.spice
* Created: Fri Aug 28 17:50:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nor4b_4.pex.spice"
.subckt sky130_fd_sc_ms__nor4b_4  VNB VPB D_N C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_D_N_M1010_g N_A_47_88#_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.10915 AS=0.31115 PD=1.035 PS=2.85 NRD=2.424 NRS=0 M=1 R=4.93333
+ SA=75000.3 SB=75008.8 A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_A_47_88#_M1002_g N_VGND_M1010_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1332 AS=0.10915 PD=1.1 PS=1.035 NRD=12.972 NRS=0 M=1 R=4.93333 SA=75000.8
+ SB=75008.4 A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1002_d N_A_47_88#_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1332 AS=0.1295 PD=1.1 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.3
+ SB=75007.8 A=0.111 P=1.78 MULT=1
MM1011 N_Y_M1011_d N_A_47_88#_M1011_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.8
+ SB=75007.3 A=0.111 P=1.78 MULT=1
MM1028 N_Y_M1011_d N_A_47_88#_M1028_g N_VGND_M1028_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75002.2
+ SB=75006.9 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1028_s N_C_M1006_g N_Y_M1006_s VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75002.8 SB=75006.3
+ A=0.111 P=1.78 MULT=1
MM1025 N_VGND_M1025_d N_C_M1025_g N_Y_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.30525 AS=0.1036 PD=1.565 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.2
+ SB=75005.9 A=0.111 P=1.78 MULT=1
MM1030 N_VGND_M1025_d N_C_M1030_g N_Y_M1030_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.30525 AS=0.1036 PD=1.565 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.2
+ SB=75004.9 A=0.111 P=1.78 MULT=1
MM1034 N_VGND_M1034_d N_C_M1034_g N_Y_M1030_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.28305 AS=0.1036 PD=1.505 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.6
+ SB=75004.5 A=0.111 P=1.78 MULT=1
MM1004 N_Y_M1004_d N_B_M1004_g N_VGND_M1034_d VNB NLOWVT L=0.15 W=0.74 AD=0.1295
+ AS=0.28305 PD=1.09 PS=1.505 NRD=0 NRS=0 M=1 R=4.93333 SA=75005.6 SB=75003.6
+ A=0.111 P=1.78 MULT=1
MM1008 N_Y_M1004_d N_B_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74 AD=0.1295
+ AS=0.1295 PD=1.09 PS=1.09 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75006.1 SB=75003.1
+ A=0.111 P=1.78 MULT=1
MM1009 N_Y_M1009_d N_B_M1009_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75006.6 SB=75002.6
+ A=0.111 P=1.78 MULT=1
MM1019 N_Y_M1009_d N_B_M1019_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.16465 PD=1.02 PS=1.185 NRD=0 NRS=12.972 M=1 R=4.93333 SA=75007 SB=75002.2
+ A=0.111 P=1.78 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.16465 PD=1.02 PS=1.185 NRD=0 NRS=13.776 M=1 R=4.93333 SA=75007.6
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1007 N_Y_M1005_d N_A_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75008 SB=75001.1
+ A=0.111 P=1.78 MULT=1
MM1015 N_Y_M1015_d N_A_M1015_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75008.4 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1029 N_Y_M1015_d N_A_M1029_g N_VGND_M1029_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75008.9 SB=75000.3
+ A=0.111 P=1.78 MULT=1
MM1012 N_A_47_88#_M1012_d N_D_N_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.2352 PD=1.11 PS=2.24 NRD=0 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.6 A=0.1512 P=2.04 MULT=1
MM1013 N_A_47_88#_M1012_d N_D_N_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.2352 PD=1.11 PS=2.24 NRD=0 NRS=0 M=1 R=4.66667 SA=90000.6
+ SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1022 N_Y_M1022_d N_A_47_88#_M1022_g N_A_319_368#_M1022_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003.5 A=0.2016 P=2.6 MULT=1
MM1024 N_Y_M1022_d N_A_47_88#_M1024_g N_A_319_368#_M1024_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=2.6201 M=1 R=6.22222
+ SA=90000.6 SB=90003.1 A=0.2016 P=2.6 MULT=1
MM1026 N_Y_M1026_d N_A_47_88#_M1026_g N_A_319_368#_M1024_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=4.3931 M=1 R=6.22222
+ SA=90001.1 SB=90002.6 A=0.2016 P=2.6 MULT=1
MM1027 N_Y_M1026_d N_A_47_88#_M1027_g N_A_319_368#_M1027_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.6 SB=90002.1 A=0.2016 P=2.6 MULT=1
MM1000 N_A_781_368#_M1000_d N_C_M1000_g N_A_319_368#_M1027_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90002 SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1001 N_A_781_368#_M1000_d N_C_M1001_g N_A_319_368#_M1001_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1792 AS=0.1932 PD=1.44 PS=1.465 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90002.5 SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1031 N_A_781_368#_M1031_d N_C_M1031_g N_A_319_368#_M1001_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1652 AS=0.1932 PD=1.415 PS=1.465 NRD=3.5066 NRS=3.5066 M=1
+ R=6.22222 SA=90003.1 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1032 N_A_781_368#_M1031_d N_C_M1032_g N_A_319_368#_M1032_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1652 AS=0.3136 PD=1.415 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90003.5 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1014 N_A_781_368#_M1014_d N_B_M1014_g N_A_1191_368#_M1014_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1792 AS=0.3136 PD=1.44 PS=2.8 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90003.4 A=0.2016 P=2.6 MULT=1
MM1016 N_A_781_368#_M1014_d N_B_M1016_g N_A_1191_368#_M1016_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90000.7 SB=90002.9 A=0.2016 P=2.6 MULT=1
MM1017 N_A_781_368#_M1017_d N_B_M1017_g N_A_1191_368#_M1016_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.2 SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1018 N_A_781_368#_M1017_d N_B_M1018_g N_A_1191_368#_M1018_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.6 SB=90002 A=0.2016 P=2.6 MULT=1
MM1020 N_VPWR_M1020_d N_A_M1020_g N_A_1191_368#_M1018_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.1
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1021 N_VPWR_M1020_d N_A_M1021_g N_A_1191_368#_M1021_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.5
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1023 N_VPWR_M1023_d N_A_M1023_g N_A_1191_368#_M1021_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1033 N_VPWR_M1023_d N_A_M1033_g N_A_1191_368#_M1033_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.4
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX35_noxref VNB VPB NWDIODE A=19.4556 P=24.64
*
.include "sky130_fd_sc_ms__nor4b_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__nand2_2.pex.spice
* Created: Fri Aug 28 17:41:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NAND2_2%B 3 7 11 15 17 18 28
c39 15 0 8.01953e-20 $X=0.975 $Y=0.74
c40 11 0 1.53462e-19 $X=0.96 $Y=2.4
r41 27 28 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.96 $Y=1.515
+ $X2=0.975 $Y2=1.515
r42 25 27 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.77 $Y=1.515
+ $X2=0.96 $Y2=1.515
r43 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.77
+ $Y=1.515 $X2=0.77 $Y2=1.515
r44 23 25 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=0.51 $Y=1.515
+ $X2=0.77 $Y2=1.515
r45 21 23 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.515
+ $X2=0.51 $Y2=1.515
r46 18 26 11.5244 $w=4.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=0.77 $Y2=1.565
r47 17 26 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=0.72 $Y=1.565 $X2=0.77
+ $Y2=1.565
r48 13 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.35
+ $X2=0.975 $Y2=1.515
r49 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.975 $Y=1.35
+ $X2=0.975 $Y2=0.74
r50 9 27 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.68
+ $X2=0.96 $Y2=1.515
r51 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.96 $Y=1.68 $X2=0.96
+ $Y2=2.4
r52 5 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.68
+ $X2=0.51 $Y2=1.515
r53 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.51 $Y=1.68 $X2=0.51
+ $Y2=2.4
r54 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.515
r55 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NAND2_2%A 3 7 11 15 17 24 26
c45 11 0 1.47716e-19 $X=1.87 $Y=2.4
c46 7 0 1.50498e-19 $X=1.42 $Y=2.4
r47 25 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.87 $Y=1.515
+ $X2=1.885 $Y2=1.515
r48 23 25 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=1.65 $Y=1.515
+ $X2=1.87 $Y2=1.515
r49 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.65
+ $Y=1.515 $X2=1.65 $Y2=1.515
r50 21 23 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=1.42 $Y=1.515
+ $X2=1.65 $Y2=1.515
r51 19 21 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.405 $Y=1.515
+ $X2=1.42 $Y2=1.515
r52 17 24 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.65 $Y=1.665
+ $X2=1.65 $Y2=1.515
r53 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.885 $Y=1.35
+ $X2=1.885 $Y2=1.515
r54 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.885 $Y=1.35
+ $X2=1.885 $Y2=0.74
r55 9 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.87 $Y=1.68
+ $X2=1.87 $Y2=1.515
r56 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.87 $Y=1.68 $X2=1.87
+ $Y2=2.4
r57 5 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=1.68
+ $X2=1.42 $Y2=1.515
r58 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.42 $Y=1.68 $X2=1.42
+ $Y2=2.4
r59 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.35
+ $X2=1.405 $Y2=1.515
r60 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.405 $Y=1.35
+ $X2=1.405 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NAND2_2%VPWR 1 2 3 10 12 18 20 22 24 26 31 40 44
r39 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 35 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r43 32 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.35 $Y=3.33
+ $X2=1.185 $Y2=3.33
r44 32 34 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.35 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 31 43 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=1.93 $Y=3.33
+ $X2=2.165 $Y2=3.33
r46 31 34 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.93 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 30 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 27 37 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.37 $Y=3.33
+ $X2=0.185 $Y2=3.33
r50 27 29 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.37 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 26 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.02 $Y=3.33
+ $X2=1.185 $Y2=3.33
r52 26 29 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.02 $Y=3.33 $X2=0.72
+ $Y2=3.33
r53 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 24 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r56 20 43 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=2.095 $Y=3.245
+ $X2=2.165 $Y2=3.33
r57 20 22 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.095 $Y=3.245
+ $X2=2.095 $Y2=2.455
r58 16 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=3.245
+ $X2=1.185 $Y2=3.33
r59 16 18 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.185 $Y=3.245
+ $X2=1.185 $Y2=2.455
r60 12 15 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=0.245 $Y=1.985
+ $X2=0.245 $Y2=2.815
r61 10 37 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.245 $Y=3.245
+ $X2=0.185 $Y2=3.33
r62 10 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.245 $Y=3.245
+ $X2=0.245 $Y2=2.815
r63 3 22 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.96
+ $Y=1.84 $X2=2.095 $Y2=2.455
r64 2 18 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.05
+ $Y=1.84 $X2=1.185 $Y2=2.455
r65 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.815
r66 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__NAND2_2%Y 1 2 3 10 12 14 18 22 24 26 27 31 34 35
c46 27 0 8.01953e-20 $X=1.785 $Y=1.095
c47 22 0 2.98213e-19 $X=1.645 $Y=2.815
c48 12 0 1.53462e-19 $X=0.735 $Y=2.815
r49 34 35 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=1.295
+ $X2=2.16 $Y2=1.665
r50 33 35 14.2803 $w=2.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.16 $Y=1.95
+ $X2=2.16 $Y2=1.665
r51 32 34 5.76222 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.16 $Y=1.18
+ $X2=2.16 $Y2=1.295
r52 26 32 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.045 $Y=1.095
+ $X2=2.16 $Y2=1.18
r53 26 27 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.045 $Y=1.095
+ $X2=1.785 $Y2=1.095
r54 25 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=2.035
+ $X2=1.645 $Y2=2.035
r55 24 33 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.045 $Y=2.035
+ $X2=2.16 $Y2=1.95
r56 24 25 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.045 $Y=2.035
+ $X2=1.73 $Y2=2.035
r57 20 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=2.12
+ $X2=1.645 $Y2=2.035
r58 20 22 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.645 $Y=2.12
+ $X2=1.645 $Y2=2.815
r59 16 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.62 $Y=1.01
+ $X2=1.785 $Y2=1.095
r60 16 18 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.62 $Y=1.01
+ $X2=1.62 $Y2=0.86
r61 15 29 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.82 $Y=2.035
+ $X2=0.695 $Y2=2.035
r62 14 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.56 $Y=2.035
+ $X2=1.645 $Y2=2.035
r63 14 15 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.56 $Y=2.035
+ $X2=0.82 $Y2=2.035
r64 10 29 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=2.12
+ $X2=0.695 $Y2=2.035
r65 10 12 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=0.695 $Y=2.12
+ $X2=0.695 $Y2=2.815
r66 3 31 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.51
+ $Y=1.84 $X2=1.645 $Y2=2.115
r67 3 22 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.51
+ $Y=1.84 $X2=1.645 $Y2=2.815
r68 2 29 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.84 $X2=0.735 $Y2=2.115
r69 2 12 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.84 $X2=0.735 $Y2=2.815
r70 1 18 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=1.48
+ $Y=0.37 $X2=1.62 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__NAND2_2%A_27_74# 1 2 3 12 14 15 20 21 24
r34 22 24 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.12 $Y=0.425
+ $X2=2.12 $Y2=0.595
r35 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.955 $Y=0.34
+ $X2=2.12 $Y2=0.425
r36 20 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.955 $Y=0.34
+ $X2=1.275 $Y2=0.34
r37 17 19 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.19 $Y=1.01
+ $X2=1.19 $Y2=0.515
r38 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.19 $Y=0.425
+ $X2=1.275 $Y2=0.34
r39 16 19 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.19 $Y=0.425 $X2=1.19
+ $Y2=0.515
r40 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.105 $Y=1.095
+ $X2=1.19 $Y2=1.01
r41 14 15 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.105 $Y=1.095
+ $X2=0.365 $Y2=1.095
r42 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.365 $Y2=1.095
r43 10 12 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.24 $Y=1.01
+ $X2=0.24 $Y2=0.515
r44 3 24 182 $w=1.7e-07 $l=2.94321e-07 $layer=licon1_NDIFF $count=1 $X=1.96
+ $Y=0.37 $X2=2.12 $Y2=0.595
r45 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.05
+ $Y=0.37 $X2=1.19 $Y2=0.515
r46 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__NAND2_2%VGND 1 6 8 10 20 21 24
r25 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r26 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r27 17 20 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r28 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r29 15 17 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r30 13 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r31 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r32 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r33 10 12 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r34 8 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r35 8 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r36 8 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r37 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0
r38 4 6 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0.595
r39 1 6 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.595
.ends


* File: sky130_fd_sc_ms__o2bb2a_2.pex.spice
* Created: Wed Sep  2 12:24:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O2BB2A_2%B1 3 5 7 9 13
r26 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.405
+ $Y=1.615 $X2=0.405 $Y2=1.615
r27 9 13 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.405 $Y2=1.615
r28 5 12 34.0194 $w=3.43e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.51 $Y=1.78
+ $X2=0.42 $Y2=1.615
r29 5 7 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=0.51 $Y=1.78 $X2=0.51
+ $Y2=2.46
r30 1 12 38.7084 $w=3.43e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.42 $Y2=1.615
r31 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2A_2%B2 3 7 9 12
c32 3 0 1.42739e-19 $X=0.93 $Y=2.46
r33 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.615
+ $X2=0.975 $Y2=1.78
r34 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.615
+ $X2=0.975 $Y2=1.45
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.615 $X2=0.975 $Y2=1.615
r36 9 13 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=0.975 $Y2=1.615
r37 7 14 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.925 $Y=0.74
+ $X2=0.925 $Y2=1.45
r38 3 15 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=0.93 $Y=2.46 $X2=0.93
+ $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2A_2%A_270_48# 1 2 9 13 18 19 20 21 23 27 30 31
+ 32
c73 30 0 1.41594e-19 $X=1.62 $Y=1.615
r74 34 36 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.425 $Y=1.615
+ $X2=1.44 $Y2=1.615
r75 31 36 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.62 $Y=1.615
+ $X2=1.44 $Y2=1.615
r76 30 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.62 $Y=1.615
+ $X2=1.62 $Y2=1.78
r77 30 32 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.62 $Y=1.615
+ $X2=1.62 $Y2=1.45
r78 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.62
+ $Y=1.615 $X2=1.62 $Y2=1.615
r79 25 27 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.21 $Y=1.135
+ $X2=2.21 $Y2=0.81
r80 21 23 26.2757 $w=2.48e-07 $l=5.7e-07 $layer=LI1_cond $X=1.785 $Y=2.1
+ $X2=2.355 $Y2=2.1
r81 19 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.045 $Y=1.22
+ $X2=2.21 $Y2=1.135
r82 19 20 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.045 $Y=1.22
+ $X2=1.785 $Y2=1.22
r83 18 21 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.7 $Y=1.975
+ $X2=1.785 $Y2=2.1
r84 18 33 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=1.975
+ $X2=1.7 $Y2=1.78
r85 15 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.7 $Y=1.305
+ $X2=1.785 $Y2=1.22
r86 15 32 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.7 $Y=1.305
+ $X2=1.7 $Y2=1.45
r87 11 36 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.44 $Y=1.78
+ $X2=1.44 $Y2=1.615
r88 11 13 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=1.44 $Y=1.78
+ $X2=1.44 $Y2=2.46
r89 7 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.45
+ $X2=1.425 $Y2=1.615
r90 7 9 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.425 $Y=1.45
+ $X2=1.425 $Y2=0.74
r91 2 23 600 $w=1.7e-07 $l=2.52785e-07 $layer=licon1_PDIFF $count=1 $X=2.175
+ $Y=1.965 $X2=2.355 $Y2=2.14
r92 1 27 182 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_NDIFF $count=1 $X=2.065
+ $Y=0.37 $X2=2.21 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2A_2%A2_N 3 7 9 12 14 17 19
c48 19 0 1.41594e-19 $X=2.16 $Y=1.475
r49 17 20 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=1.64
+ $X2=2.16 $Y2=1.805
r50 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.16 $Y=1.64
+ $X2=2.16 $Y2=1.475
r51 14 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.16
+ $Y=1.64 $X2=2.16 $Y2=1.64
r52 10 12 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=2.25 $Y=1.16
+ $X2=2.425 $Y2=1.16
r53 7 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.425 $Y=1.085
+ $X2=2.425 $Y2=1.16
r54 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.425 $Y=1.085
+ $X2=2.425 $Y2=0.69
r55 5 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.25 $Y=1.235
+ $X2=2.25 $Y2=1.16
r56 5 19 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.25 $Y=1.235
+ $X2=2.25 $Y2=1.475
r57 3 20 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=2.085 $Y=2.385
+ $X2=2.085 $Y2=1.805
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2A_2%A1_N 3 7 9 16
c42 9 0 1.85545e-19 $X=2.64 $Y=1.665
c43 7 0 1.63062e-19 $X=2.815 $Y=0.69
r44 14 16 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=2.7 $Y=1.64
+ $X2=2.815 $Y2=1.64
r45 11 14 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.64
+ $X2=2.7 $Y2=1.64
r46 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.7 $Y=1.64
+ $X2=2.7 $Y2=1.64
r47 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.815 $Y=1.475
+ $X2=2.815 $Y2=1.64
r48 5 7 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=2.815 $Y=1.475
+ $X2=2.815 $Y2=0.69
r49 1 11 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.805
+ $X2=2.625 $Y2=1.64
r50 1 3 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=2.625 $Y=1.805
+ $X2=2.625 $Y2=2.385
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2A_2%A_204_392# 1 2 9 13 17 21 25 29 31 35 37 38
+ 40 41 42 43 44 45 55
c126 55 0 1.85545e-19 $X=3.815 $Y=1.47
c127 25 0 1.42739e-19 $X=1.215 $Y=2.115
r128 54 55 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=3.81 $Y=1.47
+ $X2=3.815 $Y2=1.47
r129 53 54 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.38 $Y=1.47
+ $X2=3.81 $Y2=1.47
r130 52 53 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.365 $Y=1.47
+ $X2=3.38 $Y2=1.47
r131 49 52 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=3.265 $Y=1.47
+ $X2=3.365 $Y2=1.47
r132 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.265
+ $Y=1.47 $X2=3.265 $Y2=1.47
r133 43 48 9.03377 $w=2.85e-07 $l=2.03912e-07 $layer=LI1_cond $X=3.17 $Y=1.635
+ $X2=3.257 $Y2=1.47
r134 43 44 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=3.17 $Y=1.635
+ $X2=3.17 $Y2=2.395
r135 41 48 10.7018 $w=2.85e-07 $l=3.24808e-07 $layer=LI1_cond $X=3.085 $Y=1.22
+ $X2=3.257 $Y2=1.47
r136 41 42 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.085 $Y=1.22
+ $X2=2.715 $Y2=1.22
r137 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.63 $Y=1.135
+ $X2=2.715 $Y2=1.22
r138 39 40 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.63 $Y=0.425
+ $X2=2.63 $Y2=1.135
r139 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.545 $Y=0.34
+ $X2=2.63 $Y2=0.425
r140 37 38 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.545 $Y=0.34
+ $X2=1.805 $Y2=0.34
r141 33 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.64 $Y=0.425
+ $X2=1.805 $Y2=0.34
r142 33 35 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=1.64 $Y=0.425
+ $X2=1.64 $Y2=0.495
r143 32 45 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.38 $Y=2.48
+ $X2=1.215 $Y2=2.48
r144 31 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.085 $Y=2.48
+ $X2=3.17 $Y2=2.395
r145 31 32 111.235 $w=1.68e-07 $l=1.705e-06 $layer=LI1_cond $X=3.085 $Y=2.48
+ $X2=1.38 $Y2=2.48
r146 27 45 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=2.565
+ $X2=1.215 $Y2=2.48
r147 27 29 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.215 $Y=2.565
+ $X2=1.215 $Y2=2.815
r148 23 45 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=2.395
+ $X2=1.215 $Y2=2.48
r149 23 25 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.215 $Y=2.395
+ $X2=1.215 $Y2=2.115
r150 19 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.81 $Y=1.305
+ $X2=3.81 $Y2=1.47
r151 19 21 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=3.81 $Y=1.305
+ $X2=3.81 $Y2=0.74
r152 15 55 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.815 $Y=1.635
+ $X2=3.815 $Y2=1.47
r153 15 17 297.363 $w=1.8e-07 $l=7.65e-07 $layer=POLY_cond $X=3.815 $Y=1.635
+ $X2=3.815 $Y2=2.4
r154 11 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.38 $Y=1.305
+ $X2=3.38 $Y2=1.47
r155 11 13 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=3.38 $Y=1.305
+ $X2=3.38 $Y2=0.74
r156 7 52 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.365 $Y=1.635
+ $X2=3.365 $Y2=1.47
r157 7 9 297.363 $w=1.8e-07 $l=7.65e-07 $layer=POLY_cond $X=3.365 $Y=1.635
+ $X2=3.365 $Y2=2.4
r158 2 29 400 $w=1.7e-07 $l=9.47497e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.96 $X2=1.215 $Y2=2.815
r159 2 25 400 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.96 $X2=1.215 $Y2=2.115
r160 1 35 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.5
+ $Y=0.37 $X2=1.64 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2A_2%VPWR 1 2 3 4 13 15 21 25 27 29 33 35 40 45
+ 54 57 61
c54 15 0 1.42909e-19 $X=0.285 $Y=2.115
r55 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r56 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r59 49 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r60 49 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r61 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r62 46 57 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=3.22 $Y=3.33
+ $X2=2.995 $Y2=3.33
r63 46 48 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.22 $Y=3.33 $X2=3.6
+ $Y2=3.33
r64 45 60 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=3.955 $Y=3.33
+ $X2=4.137 $Y2=3.33
r65 45 48 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.955 $Y=3.33
+ $X2=3.6 $Y2=3.33
r66 44 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r67 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r68 41 54 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=1.94 $Y=3.33
+ $X2=1.762 $Y2=3.33
r69 41 43 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.94 $Y=3.33 $X2=2.64
+ $Y2=3.33
r70 40 57 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=2.77 $Y=3.33
+ $X2=2.995 $Y2=3.33
r71 40 43 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.77 $Y=3.33
+ $X2=2.64 $Y2=3.33
r72 39 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r73 39 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r74 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r75 36 51 4.72267 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.45 $Y=3.33
+ $X2=0.225 $Y2=3.33
r76 36 38 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=0.45 $Y=3.33 $X2=1.2
+ $Y2=3.33
r77 35 54 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=1.585 $Y=3.33
+ $X2=1.762 $Y2=3.33
r78 35 38 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.585 $Y=3.33
+ $X2=1.2 $Y2=3.33
r79 33 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r80 33 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r81 29 32 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=4.08 $Y=1.985
+ $X2=4.08 $Y2=2.815
r82 27 60 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.08 $Y=3.245
+ $X2=4.137 $Y2=3.33
r83 27 32 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=4.08 $Y=3.245
+ $X2=4.08 $Y2=2.815
r84 23 57 1.79621 $w=4.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=3.245
+ $X2=2.995 $Y2=3.33
r85 23 25 9.16993 $w=4.48e-07 $l=3.45e-07 $layer=LI1_cond $X=2.995 $Y=3.245
+ $X2=2.995 $Y2=2.9
r86 19 54 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.762 $Y=3.245
+ $X2=1.762 $Y2=3.33
r87 19 21 11.1998 $w=3.53e-07 $l=3.45e-07 $layer=LI1_cond $X=1.762 $Y=3.245
+ $X2=1.762 $Y2=2.9
r88 15 18 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.285 $Y=2.115
+ $X2=0.285 $Y2=2.815
r89 13 51 3.0435 $w=3.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.285 $Y=3.245
+ $X2=0.225 $Y2=3.33
r90 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.285 $Y=3.245
+ $X2=0.285 $Y2=2.815
r91 4 32 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=1.84 $X2=4.04 $Y2=2.815
r92 4 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.905
+ $Y=1.84 $X2=4.04 $Y2=1.985
r93 3 25 600 $w=1.7e-07 $l=1.06584e-06 $layer=licon1_PDIFF $count=1 $X=2.715
+ $Y=1.965 $X2=2.995 $Y2=2.9
r94 2 21 600 $w=1.7e-07 $l=1.04871e-06 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.96 $X2=1.76 $Y2=2.9
r95 1 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.96 $X2=0.285 $Y2=2.815
r96 1 15 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.96 $X2=0.285 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2A_2%X 1 2 9 13 14 15 16 23 32
c33 9 0 1.63062e-19 $X=3.595 $Y=0.515
r34 21 23 1.43638 $w=3.43e-07 $l=4.3e-08 $layer=LI1_cond $X=3.597 $Y=1.992
+ $X2=3.597 $Y2=2.035
r35 15 16 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=3.597 $Y=2.405
+ $X2=3.597 $Y2=2.775
r36 14 21 0.701487 $w=3.43e-07 $l=2.1e-08 $layer=LI1_cond $X=3.597 $Y=1.971
+ $X2=3.597 $Y2=1.992
r37 14 32 8.01174 $w=3.43e-07 $l=1.51e-07 $layer=LI1_cond $X=3.597 $Y=1.971
+ $X2=3.597 $Y2=1.82
r38 14 15 11.658 $w=3.43e-07 $l=3.49e-07 $layer=LI1_cond $X=3.597 $Y=2.056
+ $X2=3.597 $Y2=2.405
r39 14 23 0.701487 $w=3.43e-07 $l=2.1e-08 $layer=LI1_cond $X=3.597 $Y=2.056
+ $X2=3.597 $Y2=2.035
r40 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.685 $Y=1.13
+ $X2=3.685 $Y2=1.82
r41 7 13 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=3.6 $Y=0.96 $X2=3.6
+ $Y2=1.13
r42 7 9 15.0834 $w=3.38e-07 $l=4.45e-07 $layer=LI1_cond $X=3.6 $Y=0.96 $X2=3.6
+ $Y2=0.515
r43 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.455
+ $Y=1.84 $X2=3.59 $Y2=1.985
r44 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.455
+ $Y=1.84 $X2=3.59 $Y2=2.815
r45 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.455
+ $Y=0.37 $X2=3.595 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2A_2%A_27_74# 1 2 9 11 12 15
c26 12 0 1.42909e-19 $X=0.365 $Y=1.195
r27 13 15 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=1.18 $Y=1.11
+ $X2=1.18 $Y2=0.515
r28 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.055 $Y=1.195
+ $X2=1.18 $Y2=1.11
r29 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.055 $Y=1.195
+ $X2=0.365 $Y2=1.195
r30 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.24 $Y=1.11
+ $X2=0.365 $Y2=1.195
r31 7 9 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=0.24 $Y=1.11 $X2=0.24
+ $Y2=0.515
r32 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1 $Y=0.37
+ $X2=1.14 $Y2=0.515
r33 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O2BB2A_2%VGND 1 2 3 12 16 18 20 22 24 29 37 43 46 50
r51 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r52 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r53 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r54 41 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r55 41 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r56 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r57 38 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.05
+ $Y2=0
r58 38 40 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.6
+ $Y2=0
r59 37 49 3.99177 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.94 $Y=0 $X2=4.13
+ $Y2=0
r60 37 40 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.94 $Y=0 $X2=3.6
+ $Y2=0
r61 36 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r62 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r63 33 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r64 32 35 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r65 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r66 30 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r67 30 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r68 29 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=3.05
+ $Y2=0
r69 29 35 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=2.64
+ $Y2=0
r70 27 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r71 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r72 24 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r73 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r74 22 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r75 22 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r76 18 49 3.1514 $w=2.5e-07 $l=1.12916e-07 $layer=LI1_cond $X=4.065 $Y=0.085
+ $X2=4.13 $Y2=0
r77 18 20 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=4.065 $Y=0.085
+ $X2=4.065 $Y2=0.515
r78 14 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.05 $Y=0.085
+ $X2=3.05 $Y2=0
r79 14 16 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.05 $Y=0.085
+ $X2=3.05 $Y2=0.495
r80 10 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0
r81 10 12 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.71 $Y=0.085
+ $X2=0.71 $Y2=0.495
r82 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.885
+ $Y=0.37 $X2=4.025 $Y2=0.515
r83 2 16 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=2.89
+ $Y=0.37 $X2=3.05 $Y2=0.495
r84 1 12 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.495
.ends


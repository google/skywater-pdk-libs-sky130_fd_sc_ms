* File: sky130_fd_sc_ms__a31oi_2.pxi.spice
* Created: Fri Aug 28 17:07:32 2020
* 
x_PM_SKY130_FD_SC_MS__A31OI_2%A3 N_A3_M1002_g N_A3_c_75_n N_A3_M1006_g
+ N_A3_M1011_g N_A3_M1004_g N_A3_c_77_n N_A3_c_78_n N_A3_c_79_n A3 N_A3_c_80_n
+ N_A3_c_81_n N_A3_c_82_n PM_SKY130_FD_SC_MS__A31OI_2%A3
x_PM_SKY130_FD_SC_MS__A31OI_2%A2 N_A2_M1007_g N_A2_M1003_g N_A2_M1012_g
+ N_A2_M1008_g A2 A2 N_A2_c_160_n N_A2_c_161_n PM_SKY130_FD_SC_MS__A31OI_2%A2
x_PM_SKY130_FD_SC_MS__A31OI_2%B1 N_B1_M1009_g N_B1_c_215_n N_B1_M1001_g
+ N_B1_M1013_g B1 N_B1_c_218_n PM_SKY130_FD_SC_MS__A31OI_2%B1
x_PM_SKY130_FD_SC_MS__A31OI_2%A1 N_A1_M1000_g N_A1_M1010_g N_A1_M1005_g
+ N_A1_M1014_g A1 N_A1_c_264_n PM_SKY130_FD_SC_MS__A31OI_2%A1
x_PM_SKY130_FD_SC_MS__A31OI_2%A_27_368# N_A_27_368#_M1002_d N_A_27_368#_M1003_s
+ N_A_27_368#_M1004_d N_A_27_368#_M1013_s N_A_27_368#_M1014_s
+ N_A_27_368#_c_313_n N_A_27_368#_c_314_n N_A_27_368#_c_324_n
+ N_A_27_368#_c_315_n N_A_27_368#_c_327_n N_A_27_368#_c_330_n
+ N_A_27_368#_c_333_n N_A_27_368#_c_316_n N_A_27_368#_c_317_n
+ N_A_27_368#_c_380_p N_A_27_368#_c_347_n N_A_27_368#_c_318_n
+ N_A_27_368#_c_319_n N_A_27_368#_c_341_n PM_SKY130_FD_SC_MS__A31OI_2%A_27_368#
x_PM_SKY130_FD_SC_MS__A31OI_2%VPWR N_VPWR_M1002_s N_VPWR_M1008_d N_VPWR_M1010_d
+ N_VPWR_c_383_n N_VPWR_c_384_n N_VPWR_c_385_n VPWR N_VPWR_c_386_n
+ N_VPWR_c_387_n N_VPWR_c_388_n N_VPWR_c_389_n N_VPWR_c_382_n N_VPWR_c_391_n
+ N_VPWR_c_392_n N_VPWR_c_393_n PM_SKY130_FD_SC_MS__A31OI_2%VPWR
x_PM_SKY130_FD_SC_MS__A31OI_2%Y N_Y_M1001_d N_Y_M1005_s N_Y_M1009_d N_Y_c_449_n
+ N_Y_c_439_n N_Y_c_446_n N_Y_c_447_n N_Y_c_440_n N_Y_c_441_n N_Y_c_442_n
+ N_Y_c_443_n N_Y_c_444_n Y Y PM_SKY130_FD_SC_MS__A31OI_2%Y
x_PM_SKY130_FD_SC_MS__A31OI_2%VGND N_VGND_M1006_d N_VGND_M1011_d N_VGND_c_503_n
+ N_VGND_c_504_n N_VGND_c_505_n VGND N_VGND_c_506_n N_VGND_c_507_n
+ N_VGND_c_508_n N_VGND_c_509_n PM_SKY130_FD_SC_MS__A31OI_2%VGND
x_PM_SKY130_FD_SC_MS__A31OI_2%A_114_74# N_A_114_74#_M1006_s N_A_114_74#_M1012_d
+ N_A_114_74#_c_554_n N_A_114_74#_c_549_n N_A_114_74#_c_550_n
+ N_A_114_74#_c_551_n PM_SKY130_FD_SC_MS__A31OI_2%A_114_74#
x_PM_SKY130_FD_SC_MS__A31OI_2%A_200_74# N_A_200_74#_M1007_s N_A_200_74#_M1000_d
+ N_A_200_74#_c_579_n N_A_200_74#_c_589_n N_A_200_74#_c_581_n
+ PM_SKY130_FD_SC_MS__A31OI_2%A_200_74#
cc_1 VNB N_A3_M1002_g 0.0093723f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A3_c_75_n 0.0180369f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_3 VNB N_A3_M1004_g 0.00642655f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_4 VNB N_A3_c_77_n 0.013953f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.175
cc_5 VNB N_A3_c_78_n 0.00327939f $X=-0.19 $Y=-0.245 $X2=1.95 $Y2=1.175
cc_6 VNB N_A3_c_79_n 0.0322354f $X=-0.19 $Y=-0.245 $X2=1.95 $Y2=1.385
cc_7 VNB N_A3_c_80_n 0.059187f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.385
cc_8 VNB N_A3_c_81_n 0.0176884f $X=-0.19 $Y=-0.245 $X2=1.95 $Y2=1.22
cc_9 VNB N_A3_c_82_n 0.00919567f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.175
cc_10 VNB N_A2_M1007_g 0.0225868f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_11 VNB N_A2_M1012_g 0.0233616f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.55
cc_12 VNB N_A2_c_160_n 0.00687509f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_13 VNB N_A2_c_161_n 0.0373512f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_14 VNB N_B1_M1009_g 0.00604014f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_15 VNB N_B1_c_215_n 0.0204105f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.22
cc_16 VNB N_B1_M1013_g 0.00617181f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.74
cc_17 VNB B1 0.00737967f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_18 VNB N_B1_c_218_n 0.053602f $X=-0.19 $Y=-0.245 $X2=1.95 $Y2=1.385
cc_19 VNB N_A1_M1000_g 0.0235927f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_20 VNB N_A1_M1005_g 0.0288415f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.55
cc_21 VNB A1 0.0129671f $X=-0.19 $Y=-0.245 $X2=1.95 $Y2=1.175
cc_22 VNB N_A1_c_264_n 0.0422277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_382_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_439_n 0.00508054f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=1.175
cc_25 VNB N_Y_c_440_n 0.00282314f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_26 VNB N_Y_c_441_n 0.0126098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_442_n 0.0162516f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_28 VNB N_Y_c_443_n 0.00170724f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_29 VNB N_Y_c_444_n 9.8643e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB Y 0.025175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_503_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_32 VNB N_VGND_c_504_n 0.0322848f $X=-0.19 $Y=-0.245 $X2=1.925 $Y2=0.74
cc_33 VNB N_VGND_c_505_n 0.00888639f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_34 VNB N_VGND_c_506_n 0.0397672f $X=-0.19 $Y=-0.245 $X2=1.95 $Y2=1.175
cc_35 VNB N_VGND_c_507_n 0.0474546f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.385
cc_36 VNB N_VGND_c_508_n 0.249272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_509_n 0.00631417f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_38 VNB N_A_114_74#_c_549_n 0.00304663f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.55
cc_39 VNB N_A_114_74#_c_550_n 0.00203753f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_40 VNB N_A_114_74#_c_551_n 0.00239627f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=2.4
cc_41 VPB N_A3_M1002_g 0.0307449f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_42 VPB N_A3_M1004_g 0.023618f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_43 VPB N_A2_M1003_g 0.0206667f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_44 VPB N_A2_M1008_g 0.0218499f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=1.175
cc_45 VPB N_A2_c_160_n 0.00850739f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_46 VPB N_A2_c_161_n 0.00570124f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_47 VPB N_B1_M1009_g 0.02154f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_48 VPB N_B1_M1013_g 0.0212445f $X=-0.19 $Y=1.66 $X2=1.925 $Y2=0.74
cc_49 VPB N_A1_M1010_g 0.0207441f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_50 VPB N_A1_M1014_g 0.0267725f $X=-0.19 $Y=1.66 $X2=1.785 $Y2=1.175
cc_51 VPB A1 0.0110833f $X=-0.19 $Y=1.66 $X2=1.95 $Y2=1.175
cc_52 VPB N_A1_c_264_n 0.0047762f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_A_27_368#_c_313_n 0.0139723f $X=-0.19 $Y=1.66 $X2=0.435 $Y2=1.175
cc_54 VPB N_A_27_368#_c_314_n 0.033959f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_A_27_368#_c_315_n 0.00275632f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_27_368#_c_316_n 0.00558777f $X=-0.19 $Y=1.66 $X2=1.95 $Y2=1.385
cc_57 VPB N_A_27_368#_c_317_n 0.00167433f $X=-0.19 $Y=1.66 $X2=1.95 $Y2=1.22
cc_58 VPB N_A_27_368#_c_318_n 0.0117346f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_27_368#_c_319_n 0.030564f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_383_n 0.00396467f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=2.4
cc_61 VPB N_VPWR_c_384_n 0.00845772f $X=-0.19 $Y=1.66 $X2=0.435 $Y2=1.175
cc_62 VPB N_VPWR_c_385_n 0.00396467f $X=-0.19 $Y=1.66 $X2=1.95 $Y2=1.385
cc_63 VPB N_VPWR_c_386_n 0.0180274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_387_n 0.0194914f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.385
cc_65 VPB N_VPWR_c_388_n 0.038009f $X=-0.19 $Y=1.66 $X2=1.95 $Y2=1.55
cc_66 VPB N_VPWR_c_389_n 0.017793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_382_n 0.0649226f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_391_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_392_n 0.0047791f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_393_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_Y_c_446_n 0.006074f $X=-0.19 $Y=1.66 $X2=1.95 $Y2=1.385
cc_72 VPB N_Y_c_447_n 0.00223855f $X=-0.19 $Y=1.66 $X2=1.95 $Y2=1.385
cc_73 VPB N_Y_c_440_n 5.82959e-19 $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_74 N_A3_c_75_n N_A2_M1007_g 0.014776f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_75 N_A3_c_77_n N_A2_M1007_g 0.0126743f $X=1.785 $Y=1.175 $X2=0 $Y2=0
cc_76 N_A3_c_80_n N_A2_M1007_g 0.0154884f $X=0.505 $Y=1.385 $X2=0 $Y2=0
cc_77 N_A3_c_82_n N_A2_M1007_g 9.30523e-19 $X=0.27 $Y=1.175 $X2=0 $Y2=0
cc_78 N_A3_M1002_g N_A2_M1003_g 0.0190654f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_79 N_A3_c_77_n N_A2_M1012_g 0.0108498f $X=1.785 $Y=1.175 $X2=0 $Y2=0
cc_80 N_A3_c_78_n N_A2_M1012_g 6.94001e-19 $X=1.95 $Y=1.175 $X2=0 $Y2=0
cc_81 N_A3_c_79_n N_A2_M1012_g 0.00596063f $X=1.95 $Y=1.385 $X2=0 $Y2=0
cc_82 N_A3_c_81_n N_A2_M1012_g 0.0288704f $X=1.95 $Y=1.22 $X2=0 $Y2=0
cc_83 N_A3_M1004_g N_A2_c_160_n 0.00140212f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_84 N_A3_c_77_n N_A2_c_160_n 0.070864f $X=1.785 $Y=1.175 $X2=0 $Y2=0
cc_85 N_A3_c_78_n N_A2_c_160_n 0.0072012f $X=1.95 $Y=1.175 $X2=0 $Y2=0
cc_86 N_A3_c_79_n N_A2_c_160_n 4.37274e-19 $X=1.95 $Y=1.385 $X2=0 $Y2=0
cc_87 N_A3_c_80_n N_A2_c_160_n 0.00889759f $X=0.505 $Y=1.385 $X2=0 $Y2=0
cc_88 N_A3_c_82_n N_A2_c_160_n 0.010034f $X=0.27 $Y=1.175 $X2=0 $Y2=0
cc_89 N_A3_M1004_g N_A2_c_161_n 0.0314611f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_90 N_A3_c_77_n N_A2_c_161_n 0.00572896f $X=1.785 $Y=1.175 $X2=0 $Y2=0
cc_91 N_A3_c_78_n N_A2_c_161_n 7.61756e-19 $X=1.95 $Y=1.175 $X2=0 $Y2=0
cc_92 N_A3_c_79_n N_A2_c_161_n 0.0113878f $X=1.95 $Y=1.385 $X2=0 $Y2=0
cc_93 N_A3_c_80_n N_A2_c_161_n 0.0190654f $X=0.505 $Y=1.385 $X2=0 $Y2=0
cc_94 N_A3_M1004_g N_B1_M1009_g 0.0241657f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_95 N_A3_c_78_n N_B1_c_215_n 0.00203659f $X=1.95 $Y=1.175 $X2=0 $Y2=0
cc_96 N_A3_c_81_n N_B1_c_215_n 0.025977f $X=1.95 $Y=1.22 $X2=0 $Y2=0
cc_97 N_A3_c_78_n B1 0.0251424f $X=1.95 $Y=1.175 $X2=0 $Y2=0
cc_98 N_A3_c_79_n B1 0.00114566f $X=1.95 $Y=1.385 $X2=0 $Y2=0
cc_99 N_A3_c_78_n N_B1_c_218_n 0.00131409f $X=1.95 $Y=1.175 $X2=0 $Y2=0
cc_100 N_A3_c_79_n N_B1_c_218_n 0.0212469f $X=1.95 $Y=1.385 $X2=0 $Y2=0
cc_101 N_A3_M1002_g N_A_27_368#_c_313_n 8.13654e-19 $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_102 N_A3_c_80_n N_A_27_368#_c_313_n 0.00187045f $X=0.505 $Y=1.385 $X2=0 $Y2=0
cc_103 N_A3_c_82_n N_A_27_368#_c_313_n 0.0153227f $X=0.27 $Y=1.175 $X2=0 $Y2=0
cc_104 N_A3_M1002_g N_A_27_368#_c_314_n 0.00147311f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_105 N_A3_M1002_g N_A_27_368#_c_324_n 0.0193419f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A3_c_82_n N_A_27_368#_c_324_n 0.00167764f $X=0.27 $Y=1.175 $X2=0 $Y2=0
cc_107 N_A3_M1004_g N_A_27_368#_c_315_n 6.3785e-19 $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_108 N_A3_M1004_g N_A_27_368#_c_327_n 0.0143954f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_109 N_A3_c_78_n N_A_27_368#_c_327_n 0.0075155f $X=1.95 $Y=1.175 $X2=0 $Y2=0
cc_110 N_A3_c_79_n N_A_27_368#_c_327_n 2.83709e-19 $X=1.95 $Y=1.385 $X2=0 $Y2=0
cc_111 N_A3_M1004_g N_A_27_368#_c_330_n 0.00113798f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_112 N_A3_c_78_n N_A_27_368#_c_330_n 0.00287038f $X=1.95 $Y=1.175 $X2=0 $Y2=0
cc_113 N_A3_c_79_n N_A_27_368#_c_330_n 2.41155e-19 $X=1.95 $Y=1.385 $X2=0 $Y2=0
cc_114 N_A3_M1004_g N_A_27_368#_c_333_n 0.0103322f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_115 N_A3_M1004_g N_A_27_368#_c_317_n 0.00341623f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_116 N_A3_M1002_g N_VPWR_c_383_n 0.016085f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_117 N_A3_M1004_g N_VPWR_c_384_n 0.00137311f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A3_M1002_g N_VPWR_c_386_n 0.00460063f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A3_M1004_g N_VPWR_c_388_n 0.00517089f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A3_M1002_g N_VPWR_c_382_n 0.00912296f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_121 N_A3_M1004_g N_VPWR_c_382_n 0.00977577f $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_122 N_A3_M1004_g N_Y_c_449_n 2.17386e-19 $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_123 N_A3_M1004_g N_Y_c_447_n 7.99388e-19 $X=1.955 $Y=2.4 $X2=0 $Y2=0
cc_124 N_A3_c_82_n N_VGND_M1006_d 0.0024932f $X=0.27 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_125 N_A3_c_78_n N_VGND_M1011_d 9.04723e-19 $X=1.95 $Y=1.175 $X2=0 $Y2=0
cc_126 N_A3_c_75_n N_VGND_c_504_n 0.00620694f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_127 N_A3_c_80_n N_VGND_c_504_n 0.00142564f $X=0.505 $Y=1.385 $X2=0 $Y2=0
cc_128 N_A3_c_82_n N_VGND_c_504_n 0.0217072f $X=0.27 $Y=1.175 $X2=0 $Y2=0
cc_129 N_A3_c_81_n N_VGND_c_505_n 0.00276164f $X=1.95 $Y=1.22 $X2=0 $Y2=0
cc_130 N_A3_c_75_n N_VGND_c_506_n 0.00430908f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_131 N_A3_c_81_n N_VGND_c_506_n 0.00328473f $X=1.95 $Y=1.22 $X2=0 $Y2=0
cc_132 N_A3_c_75_n N_VGND_c_508_n 0.00819438f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_133 N_A3_c_81_n N_VGND_c_508_n 0.00428654f $X=1.95 $Y=1.22 $X2=0 $Y2=0
cc_134 N_A3_c_77_n N_A_114_74#_M1006_s 0.00176461f $X=1.785 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_135 N_A3_c_77_n N_A_114_74#_M1012_d 0.00247441f $X=1.785 $Y=1.175 $X2=0 $Y2=0
cc_136 N_A3_c_75_n N_A_114_74#_c_554_n 0.00572319f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_137 N_A3_c_77_n N_A_114_74#_c_554_n 0.0170465f $X=1.785 $Y=1.175 $X2=0 $Y2=0
cc_138 N_A3_c_77_n N_A_114_74#_c_549_n 0.00270072f $X=1.785 $Y=1.175 $X2=0 $Y2=0
cc_139 N_A3_c_75_n N_A_114_74#_c_550_n 0.00332137f $X=0.495 $Y=1.22 $X2=0 $Y2=0
cc_140 N_A3_c_81_n N_A_114_74#_c_551_n 0.00514425f $X=1.95 $Y=1.22 $X2=0 $Y2=0
cc_141 N_A3_c_77_n N_A_200_74#_M1007_s 0.00251484f $X=1.785 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_142 N_A3_c_77_n N_A_200_74#_c_579_n 0.0447587f $X=1.785 $Y=1.175 $X2=0 $Y2=0
cc_143 N_A3_c_81_n N_A_200_74#_c_579_n 5.08337e-19 $X=1.95 $Y=1.22 $X2=0 $Y2=0
cc_144 N_A3_c_78_n N_A_200_74#_c_581_n 0.0161066f $X=1.95 $Y=1.175 $X2=0 $Y2=0
cc_145 N_A3_c_79_n N_A_200_74#_c_581_n 7.09629e-19 $X=1.95 $Y=1.385 $X2=0 $Y2=0
cc_146 N_A3_c_81_n N_A_200_74#_c_581_n 0.0128917f $X=1.95 $Y=1.22 $X2=0 $Y2=0
cc_147 N_A2_M1003_g N_A_27_368#_c_324_n 0.0145835f $X=0.965 $Y=2.4 $X2=0 $Y2=0
cc_148 N_A2_c_160_n N_A_27_368#_c_324_n 0.030672f $X=1.38 $Y=1.515 $X2=0 $Y2=0
cc_149 N_A2_M1008_g N_A_27_368#_c_315_n 0.0121719f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_150 N_A2_M1008_g N_A_27_368#_c_327_n 0.0131783f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_151 N_A2_c_160_n N_A_27_368#_c_327_n 0.0107289f $X=1.38 $Y=1.515 $X2=0 $Y2=0
cc_152 N_A2_M1008_g N_A_27_368#_c_333_n 5.94347e-19 $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_153 N_A2_M1008_g N_A_27_368#_c_341_n 8.84614e-19 $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_154 N_A2_c_160_n N_A_27_368#_c_341_n 0.0238144f $X=1.38 $Y=1.515 $X2=0 $Y2=0
cc_155 N_A2_c_161_n N_A_27_368#_c_341_n 8.00284e-19 $X=1.425 $Y=1.515 $X2=0
+ $Y2=0
cc_156 N_A2_M1003_g N_VPWR_c_383_n 0.0117265f $X=0.965 $Y=2.4 $X2=0 $Y2=0
cc_157 N_A2_M1008_g N_VPWR_c_383_n 6.92187e-19 $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_158 N_A2_M1008_g N_VPWR_c_384_n 0.00306788f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_159 N_A2_M1003_g N_VPWR_c_387_n 0.00490827f $X=0.965 $Y=2.4 $X2=0 $Y2=0
cc_160 N_A2_M1008_g N_VPWR_c_387_n 0.005209f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_161 N_A2_M1003_g N_VPWR_c_382_n 0.00969162f $X=0.965 $Y=2.4 $X2=0 $Y2=0
cc_162 N_A2_M1008_g N_VPWR_c_382_n 0.00983226f $X=1.455 $Y=2.4 $X2=0 $Y2=0
cc_163 N_A2_M1007_g N_VGND_c_506_n 0.00278247f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A2_M1012_g N_VGND_c_506_n 0.00278271f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A2_M1007_g N_VGND_c_508_n 0.00354182f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A2_M1012_g N_VGND_c_508_n 0.00354798f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A2_M1007_g N_A_114_74#_c_554_n 0.0070131f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_168 N_A2_M1012_g N_A_114_74#_c_554_n 6.39115e-19 $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A2_M1007_g N_A_114_74#_c_549_n 0.00848669f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A2_M1012_g N_A_114_74#_c_549_n 0.00929356f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A2_M1007_g N_A_114_74#_c_550_n 0.00184341f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A2_M1012_g N_A_114_74#_c_551_n 4.46617e-19 $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A2_M1012_g N_A_200_74#_c_579_n 0.00405243f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A2_M1012_g N_A_200_74#_c_581_n 0.00838479f $X=1.425 $Y=0.74 $X2=0 $Y2=0
cc_175 N_B1_c_215_n N_A1_M1000_g 0.0101821f $X=2.495 $Y=1.22 $X2=0 $Y2=0
cc_176 B1 N_A1_M1000_g 4.7522e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_177 N_B1_c_218_n N_A1_M1000_g 0.0155192f $X=2.865 $Y=1.385 $X2=0 $Y2=0
cc_178 N_B1_M1013_g N_A1_c_264_n 0.0193104f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_179 N_B1_c_218_n N_A1_c_264_n 0.00227531f $X=2.865 $Y=1.385 $X2=0 $Y2=0
cc_180 N_B1_M1009_g N_A_27_368#_c_316_n 0.0140316f $X=2.415 $Y=2.4 $X2=0 $Y2=0
cc_181 N_B1_M1013_g N_A_27_368#_c_316_n 0.0139924f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_182 N_B1_M1009_g N_VPWR_c_388_n 0.00333926f $X=2.415 $Y=2.4 $X2=0 $Y2=0
cc_183 N_B1_M1013_g N_VPWR_c_388_n 0.00333926f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_184 N_B1_M1009_g N_VPWR_c_382_n 0.00422893f $X=2.415 $Y=2.4 $X2=0 $Y2=0
cc_185 N_B1_M1013_g N_VPWR_c_382_n 0.00423254f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_186 N_B1_M1009_g N_Y_c_449_n 0.010868f $X=2.415 $Y=2.4 $X2=0 $Y2=0
cc_187 N_B1_M1013_g N_Y_c_449_n 0.0113362f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_188 N_B1_c_215_n N_Y_c_439_n 0.00610484f $X=2.495 $Y=1.22 $X2=0 $Y2=0
cc_189 N_B1_M1013_g N_Y_c_446_n 0.0131722f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_190 B1 N_Y_c_446_n 0.0138047f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_191 N_B1_c_218_n N_Y_c_446_n 2.7493e-19 $X=2.865 $Y=1.385 $X2=0 $Y2=0
cc_192 N_B1_M1009_g N_Y_c_447_n 0.00535352f $X=2.415 $Y=2.4 $X2=0 $Y2=0
cc_193 N_B1_M1013_g N_Y_c_447_n 0.00228619f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_194 B1 N_Y_c_447_n 0.0279189f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_195 N_B1_c_218_n N_Y_c_447_n 7.12326e-19 $X=2.865 $Y=1.385 $X2=0 $Y2=0
cc_196 N_B1_M1013_g N_Y_c_440_n 0.00342019f $X=2.865 $Y=2.4 $X2=0 $Y2=0
cc_197 B1 N_Y_c_440_n 0.0230017f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_198 N_B1_c_218_n N_Y_c_440_n 0.00185038f $X=2.865 $Y=1.385 $X2=0 $Y2=0
cc_199 N_B1_c_215_n N_Y_c_443_n 0.00178324f $X=2.495 $Y=1.22 $X2=0 $Y2=0
cc_200 B1 N_Y_c_443_n 0.00727246f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_201 N_B1_c_218_n N_Y_c_443_n 2.85775e-19 $X=2.865 $Y=1.385 $X2=0 $Y2=0
cc_202 N_B1_c_215_n N_VGND_c_505_n 0.00277948f $X=2.495 $Y=1.22 $X2=0 $Y2=0
cc_203 N_B1_c_215_n N_VGND_c_507_n 0.00328098f $X=2.495 $Y=1.22 $X2=0 $Y2=0
cc_204 N_B1_c_215_n N_VGND_c_508_n 0.00430037f $X=2.495 $Y=1.22 $X2=0 $Y2=0
cc_205 N_B1_c_215_n N_A_200_74#_c_581_n 0.014466f $X=2.495 $Y=1.22 $X2=0 $Y2=0
cc_206 B1 N_A_200_74#_c_581_n 0.0348692f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_207 N_B1_c_218_n N_A_200_74#_c_581_n 0.00274718f $X=2.865 $Y=1.385 $X2=0
+ $Y2=0
cc_208 N_A1_M1010_g N_A_27_368#_c_316_n 0.00108516f $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_209 N_A1_M1010_g N_A_27_368#_c_347_n 0.0179051f $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_210 N_A1_M1014_g N_A_27_368#_c_347_n 0.0126733f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_211 A1 N_A_27_368#_c_347_n 0.0176603f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_212 N_A1_c_264_n N_A_27_368#_c_347_n 4.64269e-19 $X=3.755 $Y=1.515 $X2=0
+ $Y2=0
cc_213 N_A1_M1010_g N_A_27_368#_c_318_n 5.24523e-19 $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_214 N_A1_M1014_g N_A_27_368#_c_318_n 0.00433757f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_215 A1 N_A_27_368#_c_318_n 0.0249167f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_216 N_A1_M1014_g N_A_27_368#_c_319_n 4.78926e-19 $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_217 N_A1_M1010_g N_VPWR_c_385_n 0.0104008f $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_218 N_A1_M1014_g N_VPWR_c_385_n 0.0140619f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_219 N_A1_M1010_g N_VPWR_c_388_n 0.00460063f $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_220 N_A1_M1014_g N_VPWR_c_389_n 0.00460063f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_221 N_A1_M1010_g N_VPWR_c_382_n 0.00909121f $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_222 N_A1_M1014_g N_VPWR_c_382_n 0.00912296f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_223 N_A1_M1010_g N_Y_c_449_n 5.42856e-19 $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_224 N_A1_M1010_g N_Y_c_446_n 0.00640365f $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_225 N_A1_M1014_g N_Y_c_446_n 5.97673e-19 $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_226 A1 N_Y_c_446_n 0.00526544f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_227 N_A1_M1000_g N_Y_c_440_n 0.00240171f $X=3.31 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A1_M1010_g N_Y_c_440_n 7.81836e-19 $X=3.365 $Y=2.4 $X2=0 $Y2=0
cc_229 N_A1_M1005_g N_Y_c_440_n 4.99051e-19 $X=3.755 $Y=0.74 $X2=0 $Y2=0
cc_230 A1 N_Y_c_440_n 0.0221538f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_231 N_A1_c_264_n N_Y_c_440_n 0.0119664f $X=3.755 $Y=1.515 $X2=0 $Y2=0
cc_232 N_A1_M1000_g N_Y_c_441_n 0.00709202f $X=3.31 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A1_M1005_g N_Y_c_441_n 0.0127318f $X=3.755 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A1_M1000_g N_Y_c_442_n 0.00571032f $X=3.31 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A1_M1005_g N_Y_c_442_n 0.0139134f $X=3.755 $Y=0.74 $X2=0 $Y2=0
cc_236 A1 N_Y_c_442_n 0.055637f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_237 N_A1_c_264_n N_Y_c_442_n 0.00582464f $X=3.755 $Y=1.515 $X2=0 $Y2=0
cc_238 N_A1_M1000_g N_Y_c_443_n 0.00471824f $X=3.31 $Y=0.74 $X2=0 $Y2=0
cc_239 N_A1_M1000_g N_Y_c_444_n 0.00605333f $X=3.31 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A1_M1005_g N_Y_c_444_n 4.69291e-19 $X=3.755 $Y=0.74 $X2=0 $Y2=0
cc_241 N_A1_M1000_g N_VGND_c_507_n 0.00278271f $X=3.31 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A1_M1005_g N_VGND_c_507_n 0.00278271f $X=3.755 $Y=0.74 $X2=0 $Y2=0
cc_243 N_A1_M1000_g N_VGND_c_508_n 0.0035626f $X=3.31 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A1_M1005_g N_VGND_c_508_n 0.00357451f $X=3.755 $Y=0.74 $X2=0 $Y2=0
cc_245 N_A1_M1005_g N_A_200_74#_c_589_n 0.00338709f $X=3.755 $Y=0.74 $X2=0 $Y2=0
cc_246 N_A1_M1000_g N_A_200_74#_c_581_n 0.0105179f $X=3.31 $Y=0.74 $X2=0 $Y2=0
cc_247 N_A_27_368#_c_324_n N_VPWR_M1002_s 0.00353353f $X=1.065 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_248 N_A_27_368#_c_327_n N_VPWR_M1008_d 0.00950071f $X=2.015 $Y=2.035 $X2=0
+ $Y2=0
cc_249 N_A_27_368#_c_347_n N_VPWR_M1010_d 0.00354527f $X=3.875 $Y=2.145 $X2=0
+ $Y2=0
cc_250 N_A_27_368#_c_314_n N_VPWR_c_383_n 0.0234083f $X=0.28 $Y=2.4 $X2=0 $Y2=0
cc_251 N_A_27_368#_c_324_n N_VPWR_c_383_n 0.0170777f $X=1.065 $Y=2.035 $X2=0
+ $Y2=0
cc_252 N_A_27_368#_c_315_n N_VPWR_c_383_n 0.0266809f $X=1.23 $Y=2.815 $X2=0
+ $Y2=0
cc_253 N_A_27_368#_c_315_n N_VPWR_c_384_n 0.0234083f $X=1.23 $Y=2.815 $X2=0
+ $Y2=0
cc_254 N_A_27_368#_c_327_n N_VPWR_c_384_n 0.0167599f $X=2.015 $Y=2.035 $X2=0
+ $Y2=0
cc_255 N_A_27_368#_c_317_n N_VPWR_c_384_n 0.0117278f $X=2.275 $Y=2.99 $X2=0
+ $Y2=0
cc_256 N_A_27_368#_c_316_n N_VPWR_c_385_n 0.0117236f $X=2.975 $Y=2.99 $X2=0
+ $Y2=0
cc_257 N_A_27_368#_c_347_n N_VPWR_c_385_n 0.0170259f $X=3.875 $Y=2.145 $X2=0
+ $Y2=0
cc_258 N_A_27_368#_c_319_n N_VPWR_c_385_n 0.022534f $X=4.04 $Y=2.465 $X2=0 $Y2=0
cc_259 N_A_27_368#_c_314_n N_VPWR_c_386_n 0.011066f $X=0.28 $Y=2.4 $X2=0 $Y2=0
cc_260 N_A_27_368#_c_315_n N_VPWR_c_387_n 0.014549f $X=1.23 $Y=2.815 $X2=0 $Y2=0
cc_261 N_A_27_368#_c_316_n N_VPWR_c_388_n 0.0640326f $X=2.975 $Y=2.99 $X2=0
+ $Y2=0
cc_262 N_A_27_368#_c_317_n N_VPWR_c_388_n 0.0185331f $X=2.275 $Y=2.99 $X2=0
+ $Y2=0
cc_263 N_A_27_368#_c_319_n N_VPWR_c_389_n 0.0124046f $X=4.04 $Y=2.465 $X2=0
+ $Y2=0
cc_264 N_A_27_368#_c_314_n N_VPWR_c_382_n 0.00915947f $X=0.28 $Y=2.4 $X2=0 $Y2=0
cc_265 N_A_27_368#_c_315_n N_VPWR_c_382_n 0.0119743f $X=1.23 $Y=2.815 $X2=0
+ $Y2=0
cc_266 N_A_27_368#_c_316_n N_VPWR_c_382_n 0.0355545f $X=2.975 $Y=2.99 $X2=0
+ $Y2=0
cc_267 N_A_27_368#_c_317_n N_VPWR_c_382_n 0.00997093f $X=2.275 $Y=2.99 $X2=0
+ $Y2=0
cc_268 N_A_27_368#_c_319_n N_VPWR_c_382_n 0.0102675f $X=4.04 $Y=2.465 $X2=0
+ $Y2=0
cc_269 N_A_27_368#_c_316_n N_Y_M1009_d 0.00165831f $X=2.975 $Y=2.99 $X2=0 $Y2=0
cc_270 N_A_27_368#_c_316_n N_Y_c_449_n 0.0159318f $X=2.975 $Y=2.99 $X2=0 $Y2=0
cc_271 N_A_27_368#_M1013_s N_Y_c_446_n 0.0022023f $X=2.955 $Y=1.84 $X2=0 $Y2=0
cc_272 N_A_27_368#_c_380_p N_Y_c_446_n 0.01719f $X=3.115 $Y=2.23 $X2=0 $Y2=0
cc_273 N_A_27_368#_c_347_n N_Y_c_446_n 0.00449434f $X=3.875 $Y=2.145 $X2=0 $Y2=0
cc_274 N_Y_c_439_n N_VGND_c_505_n 0.0183769f $X=3.098 $Y=0.417 $X2=0 $Y2=0
cc_275 N_Y_c_439_n N_VGND_c_507_n 0.0867817f $X=3.098 $Y=0.417 $X2=0 $Y2=0
cc_276 N_Y_c_441_n N_VGND_c_507_n 0.0236566f $X=3.875 $Y=0.34 $X2=0 $Y2=0
cc_277 N_Y_c_439_n N_VGND_c_508_n 0.0489046f $X=3.098 $Y=0.417 $X2=0 $Y2=0
cc_278 N_Y_c_441_n N_VGND_c_508_n 0.0128296f $X=3.875 $Y=0.34 $X2=0 $Y2=0
cc_279 N_Y_c_441_n N_A_200_74#_M1000_d 0.00226893f $X=3.875 $Y=0.34 $X2=0 $Y2=0
cc_280 N_Y_c_442_n N_A_200_74#_M1000_d 0.00192876f $X=3.875 $Y=1.175 $X2=0 $Y2=0
cc_281 N_Y_c_441_n N_A_200_74#_c_589_n 0.0104832f $X=3.875 $Y=0.34 $X2=0 $Y2=0
cc_282 N_Y_M1001_d N_A_200_74#_c_581_n 0.0190703f $X=2.57 $Y=0.37 $X2=0 $Y2=0
cc_283 N_Y_c_439_n N_A_200_74#_c_581_n 0.0440008f $X=3.098 $Y=0.417 $X2=0 $Y2=0
cc_284 N_Y_c_441_n N_A_200_74#_c_581_n 0.00438711f $X=3.875 $Y=0.34 $X2=0 $Y2=0
cc_285 N_Y_c_442_n N_A_200_74#_c_581_n 0.018569f $X=3.875 $Y=1.175 $X2=0 $Y2=0
cc_286 N_Y_c_443_n N_A_200_74#_c_581_n 0.00867519f $X=3.335 $Y=1.175 $X2=0 $Y2=0
cc_287 N_VGND_c_506_n N_A_114_74#_c_549_n 0.0423335f $X=2.045 $Y=0 $X2=0 $Y2=0
cc_288 N_VGND_c_508_n N_A_114_74#_c_549_n 0.0239357f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_289 N_VGND_c_504_n N_A_114_74#_c_550_n 0.0112234f $X=0.28 $Y=0.725 $X2=0
+ $Y2=0
cc_290 N_VGND_c_506_n N_A_114_74#_c_550_n 0.0234416f $X=2.045 $Y=0 $X2=0 $Y2=0
cc_291 N_VGND_c_508_n N_A_114_74#_c_550_n 0.0125934f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_292 N_VGND_c_505_n N_A_114_74#_c_551_n 0.0169378f $X=2.21 $Y=0.495 $X2=0
+ $Y2=0
cc_293 N_VGND_c_506_n N_A_114_74#_c_551_n 0.0221892f $X=2.045 $Y=0 $X2=0 $Y2=0
cc_294 N_VGND_c_508_n N_A_114_74#_c_551_n 0.0124106f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_295 N_VGND_M1011_d N_A_200_74#_c_581_n 0.0127148f $X=2 $Y=0.37 $X2=0 $Y2=0
cc_296 N_VGND_c_505_n N_A_200_74#_c_581_n 0.0240865f $X=2.21 $Y=0.495 $X2=0
+ $Y2=0
cc_297 N_VGND_c_506_n N_A_200_74#_c_581_n 0.00192411f $X=2.045 $Y=0 $X2=0 $Y2=0
cc_298 N_VGND_c_507_n N_A_200_74#_c_581_n 0.00190416f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_299 N_VGND_c_508_n N_A_200_74#_c_581_n 0.0114772f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_300 N_A_114_74#_c_549_n N_A_200_74#_M1007_s 0.00251484f $X=1.545 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_301 N_A_114_74#_c_549_n N_A_200_74#_c_579_n 0.0185727f $X=1.545 $Y=0.34 $X2=0
+ $Y2=0
cc_302 N_A_114_74#_M1012_d N_A_200_74#_c_581_n 0.00494481f $X=1.5 $Y=0.37 $X2=0
+ $Y2=0
cc_303 N_A_114_74#_c_549_n N_A_200_74#_c_581_n 0.00440728f $X=1.545 $Y=0.34
+ $X2=0 $Y2=0
cc_304 N_A_114_74#_c_551_n N_A_200_74#_c_581_n 0.0191402f $X=1.71 $Y=0.34 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__clkinv_4.pxi.spice
* Created: Fri Aug 28 17:20:04 2020
* 
x_PM_SKY130_FD_SC_MS__CLKINV_4%A N_A_M1002_g N_A_c_55_n N_A_M1000_g N_A_M1003_g
+ N_A_M1004_g N_A_M1001_g N_A_M1005_g N_A_M1006_g N_A_M1008_g N_A_M1007_g
+ N_A_M1009_g A A A A A N_A_c_61_n N_A_c_62_n PM_SKY130_FD_SC_MS__CLKINV_4%A
x_PM_SKY130_FD_SC_MS__CLKINV_4%VPWR N_VPWR_M1002_s N_VPWR_M1003_s N_VPWR_M1005_s
+ N_VPWR_M1007_s N_VPWR_c_163_n N_VPWR_c_164_n N_VPWR_c_165_n N_VPWR_c_166_n
+ N_VPWR_c_167_n N_VPWR_c_168_n N_VPWR_c_169_n N_VPWR_c_170_n VPWR
+ N_VPWR_c_171_n N_VPWR_c_172_n N_VPWR_c_173_n N_VPWR_c_162_n
+ PM_SKY130_FD_SC_MS__CLKINV_4%VPWR
x_PM_SKY130_FD_SC_MS__CLKINV_4%Y N_Y_M1000_d N_Y_M1008_d N_Y_M1002_d N_Y_M1004_d
+ N_Y_M1006_d N_Y_c_215_n N_Y_c_216_n N_Y_c_225_n N_Y_c_239_n N_Y_c_242_n
+ N_Y_c_226_n N_Y_c_217_n N_Y_c_253_n N_Y_c_218_n N_Y_c_227_n N_Y_c_219_n
+ N_Y_c_228_n N_Y_c_220_n N_Y_c_221_n N_Y_c_275_n N_Y_c_222_n N_Y_c_283_n Y
+ PM_SKY130_FD_SC_MS__CLKINV_4%Y
x_PM_SKY130_FD_SC_MS__CLKINV_4%VGND N_VGND_M1000_s N_VGND_M1001_s N_VGND_M1009_s
+ N_VGND_c_322_n N_VGND_c_323_n N_VGND_c_324_n VGND N_VGND_c_325_n
+ N_VGND_c_326_n N_VGND_c_327_n N_VGND_c_328_n N_VGND_c_329_n
+ PM_SKY130_FD_SC_MS__CLKINV_4%VGND
cc_1 VNB N_A_c_55_n 0.0114828f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.605
cc_2 VNB N_A_M1000_g 0.0533591f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=0.61
cc_3 VNB N_A_M1001_g 0.0463332f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.61
cc_4 VNB N_A_M1008_g 0.0390581f $X=-0.19 $Y=-0.245 $X2=2.365 $Y2=0.61
cc_5 VNB N_A_M1009_g 0.0454945f $X=-0.19 $Y=-0.245 $X2=2.82 $Y2=0.61
cc_6 VNB A 0.00410794f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.58
cc_7 VNB N_A_c_61_n 0.0113652f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.515
cc_8 VNB N_A_c_62_n 0.102332f $X=-0.19 $Y=-0.245 $X2=2.82 $Y2=1.515
cc_9 VNB N_VPWR_c_162_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.515
cc_10 VNB N_Y_c_215_n 0.0207859f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_11 VNB N_Y_c_216_n 0.00997995f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.35
cc_12 VNB N_Y_c_217_n 0.00961836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_Y_c_218_n 0.0047561f $X=-0.19 $Y=-0.245 $X2=2.805 $Y2=2.4
cc_14 VNB N_Y_c_219_n 0.015358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_Y_c_220_n 0.0110787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_Y_c_221_n 0.00940303f $X=-0.19 $Y=-0.245 $X2=0.94 $Y2=1.515
cc_17 VNB N_Y_c_222_n 0.00245776f $X=-0.19 $Y=-0.245 $X2=1.03 $Y2=1.515
cc_18 VNB Y 0.0243509f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.515
cc_19 VNB N_VGND_c_322_n 0.0138293f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.4
cc_20 VNB N_VGND_c_323_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_324_n 0.0348923f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.4
cc_22 VNB N_VGND_c_325_n 0.0299922f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.61
cc_23 VNB N_VGND_c_326_n 0.0188284f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=2.4
cc_24 VNB N_VGND_c_327_n 0.0542217f $X=-0.19 $Y=-0.245 $X2=2.365 $Y2=1.35
cc_25 VNB N_VGND_c_328_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_329_n 0.214061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VPB N_A_M1002_g 0.0238151f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_28 VPB N_A_c_55_n 9.52843e-19 $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.605
cc_29 VPB N_A_M1003_g 0.0204945f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_30 VPB N_A_M1004_g 0.020498f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_31 VPB N_A_M1005_g 0.0210675f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_32 VPB N_A_M1006_g 0.0210641f $X=-0.19 $Y=1.66 $X2=2.355 $Y2=2.4
cc_33 VPB N_A_M1007_g 0.0224075f $X=-0.19 $Y=1.66 $X2=2.805 $Y2=2.4
cc_34 VPB A 0.0135485f $X=-0.19 $Y=1.66 $X2=2.555 $Y2=1.58
cc_35 VPB N_A_c_61_n 0.00314639f $X=-0.19 $Y=1.66 $X2=0.865 $Y2=1.515
cc_36 VPB N_A_c_62_n 0.0165362f $X=-0.19 $Y=1.66 $X2=2.82 $Y2=1.515
cc_37 VPB N_VPWR_c_163_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.4
cc_38 VPB N_VPWR_c_164_n 0.0376858f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=1.68
cc_39 VPB N_VPWR_c_165_n 0.00797179f $X=-0.19 $Y=1.66 $X2=1.795 $Y2=1.35
cc_40 VPB N_VPWR_c_166_n 0.0081889f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.68
cc_41 VPB N_VPWR_c_167_n 0.0121909f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=2.4
cc_42 VPB N_VPWR_c_168_n 0.0384698f $X=-0.19 $Y=1.66 $X2=2.355 $Y2=1.68
cc_43 VPB N_VPWR_c_169_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_170_n 0.00324402f $X=-0.19 $Y=1.66 $X2=2.365 $Y2=1.35
cc_45 VPB N_VPWR_c_171_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_172_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_173_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_162_n 0.0608616f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.515
cc_49 VPB N_Y_c_215_n 0.00618364f $X=-0.19 $Y=1.66 $X2=1.405 $Y2=2.4
cc_50 VPB N_Y_c_225_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_Y_c_226_n 0.00231613f $X=-0.19 $Y=1.66 $X2=2.355 $Y2=2.4
cc_52 VPB N_Y_c_227_n 0.00231613f $X=-0.19 $Y=1.66 $X2=2.82 $Y2=0.61
cc_53 VPB N_Y_c_228_n 0.00707089f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_54 VPB Y 0.013063f $X=-0.19 $Y=1.66 $X2=1.855 $Y2=1.515
cc_55 N_A_M1002_g N_VPWR_c_164_n 0.00501904f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_56 N_A_M1003_g N_VPWR_c_165_n 0.0027763f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_57 N_A_M1004_g N_VPWR_c_165_n 0.0027763f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_58 N_A_M1005_g N_VPWR_c_166_n 0.00306788f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_59 N_A_M1006_g N_VPWR_c_166_n 0.00187311f $X=2.355 $Y=2.4 $X2=0 $Y2=0
cc_60 N_A_M1007_g N_VPWR_c_168_n 0.00394849f $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_61 N_A_M1002_g N_VPWR_c_169_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_62 N_A_M1003_g N_VPWR_c_169_n 0.005209f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_63 N_A_M1004_g N_VPWR_c_171_n 0.005209f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_64 N_A_M1005_g N_VPWR_c_171_n 0.005209f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_65 N_A_M1006_g N_VPWR_c_172_n 0.005209f $X=2.355 $Y=2.4 $X2=0 $Y2=0
cc_66 N_A_M1007_g N_VPWR_c_172_n 0.005209f $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_67 N_A_M1002_g N_VPWR_c_162_n 0.00986008f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_68 N_A_M1003_g N_VPWR_c_162_n 0.00982266f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_69 N_A_M1004_g N_VPWR_c_162_n 0.00982266f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_70 N_A_M1005_g N_VPWR_c_162_n 0.00982754f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_71 N_A_M1006_g N_VPWR_c_162_n 0.00982082f $X=2.355 $Y=2.4 $X2=0 $Y2=0
cc_72 N_A_M1007_g N_VPWR_c_162_n 0.00985497f $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_73 N_A_M1002_g N_Y_c_215_n 0.00869982f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_74 N_A_c_55_n N_Y_c_215_n 0.00534776f $X=0.595 $Y=1.605 $X2=0 $Y2=0
cc_75 N_A_M1000_g N_Y_c_215_n 0.00442873f $X=0.94 $Y=0.61 $X2=0 $Y2=0
cc_76 N_A_M1003_g N_Y_c_215_n 6.43615e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_77 A N_Y_c_215_n 0.0344967f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_78 N_A_c_62_n N_Y_c_215_n 6.94144e-19 $X=2.82 $Y=1.515 $X2=0 $Y2=0
cc_79 N_A_M1002_g N_Y_c_225_n 0.01694f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_80 N_A_M1003_g N_Y_c_225_n 0.0121623f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_81 N_A_M1004_g N_Y_c_225_n 6.51317e-19 $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_82 N_A_M1003_g N_Y_c_239_n 0.012931f $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_83 N_A_M1004_g N_Y_c_239_n 0.012931f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_84 N_A_c_62_n N_Y_c_239_n 4.90767e-19 $X=2.82 $Y=1.515 $X2=0 $Y2=0
cc_85 N_A_M1002_g N_Y_c_242_n 0.0191578f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_86 N_A_M1003_g N_Y_c_242_n 9.43996e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_87 A N_Y_c_242_n 0.0582742f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_88 N_A_c_61_n N_Y_c_242_n 4.9731e-19 $X=0.865 $Y=1.515 $X2=0 $Y2=0
cc_89 N_A_M1003_g N_Y_c_226_n 6.50516e-19 $X=0.955 $Y=2.4 $X2=0 $Y2=0
cc_90 N_A_M1004_g N_Y_c_226_n 0.0120549f $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_91 N_A_M1005_g N_Y_c_226_n 0.012298f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_92 N_A_M1006_g N_Y_c_226_n 6.3785e-19 $X=2.355 $Y=2.4 $X2=0 $Y2=0
cc_93 N_A_M1001_g N_Y_c_217_n 0.0118691f $X=1.795 $Y=0.61 $X2=0 $Y2=0
cc_94 N_A_M1008_g N_Y_c_217_n 0.0118691f $X=2.365 $Y=0.61 $X2=0 $Y2=0
cc_95 N_A_c_62_n N_Y_c_217_n 0.00577492f $X=2.82 $Y=1.515 $X2=0 $Y2=0
cc_96 N_A_M1005_g N_Y_c_253_n 0.0132272f $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_97 N_A_M1006_g N_Y_c_253_n 0.0132272f $X=2.355 $Y=2.4 $X2=0 $Y2=0
cc_98 A N_Y_c_253_n 0.0431694f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_99 N_A_c_62_n N_Y_c_253_n 7.63416e-19 $X=2.82 $Y=1.515 $X2=0 $Y2=0
cc_100 N_A_M1001_g N_Y_c_218_n 6.22763e-19 $X=1.795 $Y=0.61 $X2=0 $Y2=0
cc_101 N_A_M1008_g N_Y_c_218_n 0.0110981f $X=2.365 $Y=0.61 $X2=0 $Y2=0
cc_102 N_A_M1009_g N_Y_c_218_n 0.00547196f $X=2.82 $Y=0.61 $X2=0 $Y2=0
cc_103 N_A_M1005_g N_Y_c_227_n 6.10838e-19 $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_104 N_A_M1006_g N_Y_c_227_n 0.0118128f $X=2.355 $Y=2.4 $X2=0 $Y2=0
cc_105 N_A_M1007_g N_Y_c_227_n 0.016185f $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A_M1009_g N_Y_c_219_n 0.0187429f $X=2.82 $Y=0.61 $X2=0 $Y2=0
cc_107 A N_Y_c_219_n 6.95742e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_108 N_A_M1007_g N_Y_c_228_n 0.0187429f $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_109 A N_Y_c_228_n 6.95742e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_110 N_A_c_55_n N_Y_c_220_n 0.00579235f $X=0.595 $Y=1.605 $X2=0 $Y2=0
cc_111 N_A_M1000_g N_Y_c_220_n 0.0130527f $X=0.94 $Y=0.61 $X2=0 $Y2=0
cc_112 A N_Y_c_220_n 0.144874f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_113 N_A_c_61_n N_Y_c_220_n 0.00118654f $X=0.865 $Y=1.515 $X2=0 $Y2=0
cc_114 N_A_M1000_g N_Y_c_221_n 0.0256826f $X=0.94 $Y=0.61 $X2=0 $Y2=0
cc_115 N_A_M1001_g N_Y_c_221_n 0.0162981f $X=1.795 $Y=0.61 $X2=0 $Y2=0
cc_116 N_A_M1008_g N_Y_c_221_n 6.05295e-19 $X=2.365 $Y=0.61 $X2=0 $Y2=0
cc_117 N_A_c_62_n N_Y_c_221_n 0.0137608f $X=2.82 $Y=1.515 $X2=0 $Y2=0
cc_118 N_A_M1004_g N_Y_c_275_n 8.84614e-19 $X=1.405 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A_M1005_g N_Y_c_275_n 8.84614e-19 $X=1.855 $Y=2.4 $X2=0 $Y2=0
cc_120 A N_Y_c_275_n 0.0235495f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_121 N_A_c_62_n N_Y_c_275_n 5.51595e-19 $X=2.82 $Y=1.515 $X2=0 $Y2=0
cc_122 N_A_M1008_g N_Y_c_222_n 0.00294386f $X=2.365 $Y=0.61 $X2=0 $Y2=0
cc_123 N_A_M1009_g N_Y_c_222_n 0.00218126f $X=2.82 $Y=0.61 $X2=0 $Y2=0
cc_124 A N_Y_c_222_n 0.028235f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_125 N_A_c_62_n N_Y_c_222_n 0.00305f $X=2.82 $Y=1.515 $X2=0 $Y2=0
cc_126 N_A_M1006_g N_Y_c_283_n 8.84614e-19 $X=2.355 $Y=2.4 $X2=0 $Y2=0
cc_127 N_A_M1007_g N_Y_c_283_n 8.84614e-19 $X=2.805 $Y=2.4 $X2=0 $Y2=0
cc_128 A N_Y_c_283_n 0.0235495f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_129 N_A_c_62_n N_Y_c_283_n 5.54777e-19 $X=2.82 $Y=1.515 $X2=0 $Y2=0
cc_130 N_A_M1009_g Y 0.0249699f $X=2.82 $Y=0.61 $X2=0 $Y2=0
cc_131 A Y 0.0261103f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_132 N_A_M1001_g N_VGND_c_322_n 0.00651086f $X=1.795 $Y=0.61 $X2=0 $Y2=0
cc_133 N_A_M1008_g N_VGND_c_322_n 0.00473938f $X=2.365 $Y=0.61 $X2=0 $Y2=0
cc_134 N_A_M1009_g N_VGND_c_324_n 0.00492488f $X=2.82 $Y=0.61 $X2=0 $Y2=0
cc_135 N_A_M1000_g N_VGND_c_325_n 0.0053111f $X=0.94 $Y=0.61 $X2=0 $Y2=0
cc_136 N_A_M1001_g N_VGND_c_325_n 0.0053111f $X=1.795 $Y=0.61 $X2=0 $Y2=0
cc_137 N_A_M1008_g N_VGND_c_326_n 0.00530655f $X=2.365 $Y=0.61 $X2=0 $Y2=0
cc_138 N_A_M1009_g N_VGND_c_326_n 0.0055601f $X=2.82 $Y=0.61 $X2=0 $Y2=0
cc_139 N_A_M1000_g N_VGND_c_327_n 0.012091f $X=0.94 $Y=0.61 $X2=0 $Y2=0
cc_140 N_A_M1000_g N_VGND_c_329_n 0.00536257f $X=0.94 $Y=0.61 $X2=0 $Y2=0
cc_141 N_A_M1001_g N_VGND_c_329_n 0.00536257f $X=1.795 $Y=0.61 $X2=0 $Y2=0
cc_142 N_A_M1008_g N_VGND_c_329_n 0.00536257f $X=2.365 $Y=0.61 $X2=0 $Y2=0
cc_143 N_A_M1009_g N_VGND_c_329_n 0.00536257f $X=2.82 $Y=0.61 $X2=0 $Y2=0
cc_144 N_VPWR_M1002_s N_Y_c_215_n 0.00446915f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_145 N_VPWR_c_164_n N_Y_c_225_n 0.0234083f $X=0.28 $Y=2.455 $X2=0 $Y2=0
cc_146 N_VPWR_c_165_n N_Y_c_225_n 0.0233699f $X=1.18 $Y=2.455 $X2=0 $Y2=0
cc_147 N_VPWR_c_169_n N_Y_c_225_n 0.0144623f $X=1.095 $Y=3.33 $X2=0 $Y2=0
cc_148 N_VPWR_c_162_n N_Y_c_225_n 0.0118344f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_149 N_VPWR_M1003_s N_Y_c_239_n 0.00314376f $X=1.045 $Y=1.84 $X2=0 $Y2=0
cc_150 N_VPWR_c_165_n N_Y_c_239_n 0.0126919f $X=1.18 $Y=2.455 $X2=0 $Y2=0
cc_151 N_VPWR_M1002_s N_Y_c_242_n 0.00882858f $X=0.135 $Y=1.84 $X2=0 $Y2=0
cc_152 N_VPWR_c_164_n N_Y_c_242_n 0.00752987f $X=0.28 $Y=2.455 $X2=0 $Y2=0
cc_153 N_VPWR_c_165_n N_Y_c_226_n 0.0233699f $X=1.18 $Y=2.455 $X2=0 $Y2=0
cc_154 N_VPWR_c_166_n N_Y_c_226_n 0.0234083f $X=2.08 $Y=2.455 $X2=0 $Y2=0
cc_155 N_VPWR_c_171_n N_Y_c_226_n 0.0144623f $X=1.995 $Y=3.33 $X2=0 $Y2=0
cc_156 N_VPWR_c_162_n N_Y_c_226_n 0.0118344f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_157 N_VPWR_M1005_s N_Y_c_253_n 0.00410979f $X=1.945 $Y=1.84 $X2=0 $Y2=0
cc_158 N_VPWR_c_166_n N_Y_c_253_n 0.0167599f $X=2.08 $Y=2.455 $X2=0 $Y2=0
cc_159 N_VPWR_c_166_n N_Y_c_227_n 0.0266484f $X=2.08 $Y=2.455 $X2=0 $Y2=0
cc_160 N_VPWR_c_168_n N_Y_c_227_n 0.0266809f $X=3.08 $Y=2.455 $X2=0 $Y2=0
cc_161 N_VPWR_c_172_n N_Y_c_227_n 0.0144623f $X=2.915 $Y=3.33 $X2=0 $Y2=0
cc_162 N_VPWR_c_162_n N_Y_c_227_n 0.0118344f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_163 N_VPWR_M1007_s N_Y_c_228_n 0.0063718f $X=2.895 $Y=1.84 $X2=0 $Y2=0
cc_164 N_VPWR_c_168_n N_Y_c_228_n 0.0249562f $X=3.08 $Y=2.455 $X2=0 $Y2=0
cc_165 N_VPWR_M1007_s Y 0.00217208f $X=2.895 $Y=1.84 $X2=0 $Y2=0
cc_166 N_Y_c_217_n N_VGND_c_322_n 0.0277029f $X=2.415 $Y=1.095 $X2=0 $Y2=0
cc_167 N_Y_c_218_n N_VGND_c_322_n 0.0188413f $X=2.58 $Y=0.61 $X2=0 $Y2=0
cc_168 N_Y_c_221_n N_VGND_c_322_n 0.0169695f $X=1.745 $Y=0.817 $X2=0 $Y2=0
cc_169 N_Y_c_218_n N_VGND_c_324_n 0.0193875f $X=2.58 $Y=0.61 $X2=0 $Y2=0
cc_170 N_Y_c_219_n N_VGND_c_324_n 0.0290296f $X=3.005 $Y=1.095 $X2=0 $Y2=0
cc_171 N_Y_c_221_n N_VGND_c_325_n 0.0210518f $X=1.745 $Y=0.817 $X2=0 $Y2=0
cc_172 N_Y_c_218_n N_VGND_c_326_n 0.012991f $X=2.58 $Y=0.61 $X2=0 $Y2=0
cc_173 N_Y_c_216_n N_VGND_c_327_n 0.0103794f $X=0.435 $Y=1.095 $X2=0 $Y2=0
cc_174 N_Y_c_220_n N_VGND_c_327_n 0.0207787f $X=0.99 $Y=0.817 $X2=0 $Y2=0
cc_175 N_Y_c_218_n N_VGND_c_329_n 0.0118717f $X=2.58 $Y=0.61 $X2=0 $Y2=0
cc_176 N_Y_c_221_n N_VGND_c_329_n 0.0259639f $X=1.745 $Y=0.817 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__a32oi_1.pxi.spice
* Created: Fri Aug 28 17:08:37 2020
* 
x_PM_SKY130_FD_SC_MS__A32OI_1%B2 N_B2_M1003_g N_B2_c_52_n N_B2_M1005_g B2
+ N_B2_c_54_n PM_SKY130_FD_SC_MS__A32OI_1%B2
x_PM_SKY130_FD_SC_MS__A32OI_1%B1 N_B1_c_75_n N_B1_M1000_g N_B1_M1002_g B1
+ N_B1_c_78_n PM_SKY130_FD_SC_MS__A32OI_1%B1
x_PM_SKY130_FD_SC_MS__A32OI_1%A1 N_A1_M1006_g N_A1_c_108_n N_A1_M1008_g A1
+ N_A1_c_110_n PM_SKY130_FD_SC_MS__A32OI_1%A1
x_PM_SKY130_FD_SC_MS__A32OI_1%A2 N_A2_M1009_g N_A2_M1004_g A2 A2 A2 N_A2_c_142_n
+ N_A2_c_143_n PM_SKY130_FD_SC_MS__A32OI_1%A2
x_PM_SKY130_FD_SC_MS__A32OI_1%A3 N_A3_M1001_g N_A3_M1007_g A3 N_A3_c_182_n
+ N_A3_c_183_n PM_SKY130_FD_SC_MS__A32OI_1%A3
x_PM_SKY130_FD_SC_MS__A32OI_1%A_27_368# N_A_27_368#_M1003_s N_A_27_368#_M1002_d
+ N_A_27_368#_M1004_d N_A_27_368#_c_207_n N_A_27_368#_c_208_n
+ N_A_27_368#_c_209_n N_A_27_368#_c_220_n N_A_27_368#_c_221_n
+ N_A_27_368#_c_222_n N_A_27_368#_c_210_n N_A_27_368#_c_211_n
+ N_A_27_368#_c_228_n PM_SKY130_FD_SC_MS__A32OI_1%A_27_368#
x_PM_SKY130_FD_SC_MS__A32OI_1%Y N_Y_M1000_d N_Y_M1003_d N_Y_c_257_n N_Y_c_271_n
+ N_Y_c_258_n N_Y_c_259_n N_Y_c_261_n Y N_Y_c_263_n
+ PM_SKY130_FD_SC_MS__A32OI_1%Y
x_PM_SKY130_FD_SC_MS__A32OI_1%VPWR N_VPWR_M1006_d N_VPWR_M1007_d N_VPWR_c_310_n
+ N_VPWR_c_311_n VPWR N_VPWR_c_312_n N_VPWR_c_313_n N_VPWR_c_314_n
+ N_VPWR_c_309_n PM_SKY130_FD_SC_MS__A32OI_1%VPWR
x_PM_SKY130_FD_SC_MS__A32OI_1%VGND N_VGND_M1005_s N_VGND_M1001_d N_VGND_c_348_n
+ N_VGND_c_349_n N_VGND_c_350_n N_VGND_c_351_n VGND N_VGND_c_352_n
+ N_VGND_c_353_n PM_SKY130_FD_SC_MS__A32OI_1%VGND
cc_1 VNB N_B2_M1003_g 0.00952444f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_B2_c_52_n 0.0199632f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.22
cc_3 VNB B2 0.00806923f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_B2_c_54_n 0.058145f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.385
cc_5 VNB N_B1_c_75_n 0.0229989f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.55
cc_6 VNB N_B1_M1002_g 0.0069754f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.74
cc_7 VNB B1 0.00758946f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_B1_c_78_n 0.0415823f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.385
cc_9 VNB N_A1_M1006_g 0.00798022f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_10 VNB N_A1_c_108_n 0.0231454f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.22
cc_11 VNB A1 0.00429394f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_12 VNB N_A1_c_110_n 0.0417548f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.385
cc_13 VNB N_A2_M1004_g 0.00736631f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.74
cc_14 VNB A2 0.00819917f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_15 VNB N_A2_c_142_n 0.0306202f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.385
cc_16 VNB N_A2_c_143_n 0.0174586f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.295
cc_17 VNB N_A3_M1007_g 0.00936933f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.74
cc_18 VNB A3 0.0219295f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_19 VNB N_A3_c_182_n 0.0350799f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_20 VNB N_A3_c_183_n 0.0223315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_257_n 0.0100996f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_22 VNB N_Y_c_258_n 0.00159849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_259_n 0.00778594f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.385
cc_24 VNB N_VPWR_c_309_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_348_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.74
cc_26 VNB N_VGND_c_349_n 0.0377474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_350_n 0.0128247f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.385
cc_28 VNB N_VGND_c_351_n 0.0344702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_352_n 0.0649785f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.295
cc_30 VNB N_VGND_c_353_n 0.215051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VPB N_B2_M1003_g 0.0298002f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_32 VPB N_B1_M1002_g 0.0231154f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.74
cc_33 VPB N_A1_M1006_g 0.0259112f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_34 VPB N_A2_M1004_g 0.0255463f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.74
cc_35 VPB N_A3_M1007_g 0.0285741f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.74
cc_36 VPB N_A_27_368#_c_207_n 0.0434878f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.385
cc_37 VPB N_A_27_368#_c_208_n 0.00629259f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_A_27_368#_c_209_n 0.00965867f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.295
cc_39 VPB N_A_27_368#_c_210_n 0.0100338f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A_27_368#_c_211_n 0.00229053f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_Y_c_257_n 0.00132726f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_42 VPB N_Y_c_261_n 0.00461959f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 VPB Y 0.0101374f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.385
cc_44 VPB N_Y_c_263_n 0.00893879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_310_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=0.74
cc_46 VPB N_VPWR_c_311_n 0.0564405f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_312_n 0.042496f $X=-0.19 $Y=1.66 $X2=0.52 $Y2=1.385
cc_48 VPB N_VPWR_c_313_n 0.0183219f $X=-0.19 $Y=1.66 $X2=0.28 $Y2=1.385
cc_49 VPB N_VPWR_c_314_n 0.0185351f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_309_n 0.0574653f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 N_B2_c_52_n N_B1_c_75_n 0.0321121f $X=0.52 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_52 N_B2_M1003_g N_B1_M1002_g 0.0278996f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_53 N_B2_c_54_n N_B1_c_78_n 0.0321121f $X=0.52 $Y=1.385 $X2=0 $Y2=0
cc_54 N_B2_M1003_g N_A_27_368#_c_207_n 0.0157774f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_55 B2 N_A_27_368#_c_207_n 0.0196739f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_56 N_B2_c_54_n N_A_27_368#_c_207_n 0.00223706f $X=0.52 $Y=1.385 $X2=0 $Y2=0
cc_57 N_B2_M1003_g N_A_27_368#_c_208_n 0.0118818f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_58 N_B2_M1003_g N_A_27_368#_c_209_n 0.00291251f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_59 N_B2_c_52_n N_Y_c_257_n 0.00939186f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_60 B2 N_Y_c_257_n 0.0279669f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_61 N_B2_c_52_n N_Y_c_258_n 0.00269193f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_62 N_B2_M1003_g N_Y_c_261_n 0.00356709f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_63 N_B2_M1003_g N_VPWR_c_312_n 0.00333896f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_64 N_B2_M1003_g N_VPWR_c_309_n 0.00426993f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_65 N_B2_c_52_n N_VGND_c_349_n 0.00533858f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_66 B2 N_VGND_c_349_n 0.0263177f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_67 N_B2_c_54_n N_VGND_c_349_n 0.00216978f $X=0.52 $Y=1.385 $X2=0 $Y2=0
cc_68 N_B2_c_52_n N_VGND_c_352_n 0.00460063f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_69 N_B2_c_52_n N_VGND_c_353_n 0.00910551f $X=0.52 $Y=1.22 $X2=0 $Y2=0
cc_70 N_B1_M1002_g N_A1_M1006_g 0.0279432f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_71 B1 A1 0.0253469f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_72 N_B1_c_78_n A1 3.96911e-19 $X=1.12 $Y=1.385 $X2=0 $Y2=0
cc_73 B1 N_A1_c_110_n 0.0020937f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_74 N_B1_c_78_n N_A1_c_110_n 0.0178871f $X=1.12 $Y=1.385 $X2=0 $Y2=0
cc_75 N_B1_M1002_g N_A_27_368#_c_207_n 7.65597e-19 $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_76 N_B1_M1002_g N_A_27_368#_c_208_n 0.0145636f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_77 N_B1_c_75_n N_Y_c_257_n 0.00474996f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_78 N_B1_M1002_g N_Y_c_257_n 0.00377659f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_79 B1 N_Y_c_257_n 0.0279522f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_80 N_B1_M1002_g N_Y_c_271_n 0.0138833f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_81 N_B1_c_75_n N_Y_c_259_n 0.0228512f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_82 B1 N_Y_c_259_n 0.0284419f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_83 N_B1_c_78_n N_Y_c_259_n 0.00194618f $X=1.12 $Y=1.385 $X2=0 $Y2=0
cc_84 N_B1_M1002_g N_Y_c_261_n 0.00337881f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_85 N_B1_c_78_n N_Y_c_261_n 0.00387084f $X=1.12 $Y=1.385 $X2=0 $Y2=0
cc_86 N_B1_M1002_g Y 5.4014e-19 $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_87 N_B1_M1002_g N_Y_c_263_n 0.01399f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_88 B1 N_Y_c_263_n 0.0268776f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_89 N_B1_c_78_n N_Y_c_263_n 0.0013394f $X=1.12 $Y=1.385 $X2=0 $Y2=0
cc_90 N_B1_M1002_g N_VPWR_c_312_n 0.00333926f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_91 N_B1_M1002_g N_VPWR_c_309_n 0.00424688f $X=1.005 $Y=2.4 $X2=0 $Y2=0
cc_92 N_B1_c_75_n N_VGND_c_352_n 0.00291649f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_93 N_B1_c_75_n N_VGND_c_353_n 0.0036383f $X=0.91 $Y=1.22 $X2=0 $Y2=0
cc_94 N_A1_M1006_g N_A2_M1004_g 0.0200156f $X=1.615 $Y=2.4 $X2=0 $Y2=0
cc_95 N_A1_c_108_n A2 0.0118388f $X=1.88 $Y=1.22 $X2=0 $Y2=0
cc_96 A1 A2 0.0277288f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_97 N_A1_c_110_n N_A2_c_142_n 0.033517f $X=1.88 $Y=1.385 $X2=0 $Y2=0
cc_98 N_A1_c_108_n N_A2_c_143_n 0.033517f $X=1.88 $Y=1.22 $X2=0 $Y2=0
cc_99 A1 N_A2_c_143_n 3.10488e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_100 N_A1_M1006_g N_A_27_368#_c_208_n 0.00184533f $X=1.615 $Y=2.4 $X2=0 $Y2=0
cc_101 N_A1_M1006_g N_A_27_368#_c_220_n 0.00539532f $X=1.615 $Y=2.4 $X2=0 $Y2=0
cc_102 N_A1_M1006_g N_A_27_368#_c_221_n 0.00724838f $X=1.615 $Y=2.4 $X2=0 $Y2=0
cc_103 N_A1_M1006_g N_A_27_368#_c_222_n 0.0155765f $X=1.615 $Y=2.4 $X2=0 $Y2=0
cc_104 N_A1_M1006_g N_Y_c_271_n 7.22837e-19 $X=1.615 $Y=2.4 $X2=0 $Y2=0
cc_105 N_A1_c_108_n N_Y_c_259_n 0.00905028f $X=1.88 $Y=1.22 $X2=0 $Y2=0
cc_106 A1 N_Y_c_259_n 0.0237588f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_107 N_A1_c_110_n N_Y_c_259_n 0.0017926f $X=1.88 $Y=1.385 $X2=0 $Y2=0
cc_108 N_A1_M1006_g Y 0.0193405f $X=1.615 $Y=2.4 $X2=0 $Y2=0
cc_109 N_A1_c_110_n Y 0.00573163f $X=1.88 $Y=1.385 $X2=0 $Y2=0
cc_110 N_A1_M1006_g N_Y_c_263_n 0.00603417f $X=1.615 $Y=2.4 $X2=0 $Y2=0
cc_111 A1 N_Y_c_263_n 0.0257356f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_112 N_A1_M1006_g N_VPWR_c_312_n 0.00461464f $X=1.615 $Y=2.4 $X2=0 $Y2=0
cc_113 N_A1_M1006_g N_VPWR_c_314_n 0.0091917f $X=1.615 $Y=2.4 $X2=0 $Y2=0
cc_114 N_A1_M1006_g N_VPWR_c_309_n 0.00462294f $X=1.615 $Y=2.4 $X2=0 $Y2=0
cc_115 N_A1_c_108_n N_VGND_c_352_n 0.00433162f $X=1.88 $Y=1.22 $X2=0 $Y2=0
cc_116 N_A1_c_108_n N_VGND_c_353_n 0.00822327f $X=1.88 $Y=1.22 $X2=0 $Y2=0
cc_117 N_A2_M1004_g N_A3_M1007_g 0.0230682f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_118 A2 A3 0.0223908f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_119 N_A2_c_142_n A3 0.00121116f $X=2.36 $Y=1.385 $X2=0 $Y2=0
cc_120 A2 N_A3_c_182_n 4.18785e-19 $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_121 N_A2_c_142_n N_A3_c_182_n 0.017626f $X=2.36 $Y=1.385 $X2=0 $Y2=0
cc_122 A2 N_A3_c_183_n 0.00950494f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_123 N_A2_c_143_n N_A3_c_183_n 0.0241574f $X=2.36 $Y=1.22 $X2=0 $Y2=0
cc_124 N_A2_M1004_g N_A_27_368#_c_222_n 0.0153941f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_125 N_A2_M1004_g N_A_27_368#_c_210_n 0.0125697f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_126 A2 N_A_27_368#_c_210_n 0.0035131f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_127 N_A2_c_142_n N_A_27_368#_c_210_n 2.15726e-19 $X=2.36 $Y=1.385 $X2=0 $Y2=0
cc_128 N_A2_M1004_g N_A_27_368#_c_211_n 2.69566e-19 $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_129 N_A2_M1004_g N_A_27_368#_c_228_n 0.00121691f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_130 A2 N_Y_c_259_n 0.0401943f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_131 N_A2_c_143_n N_Y_c_259_n 9.06958e-19 $X=2.36 $Y=1.22 $X2=0 $Y2=0
cc_132 N_A2_M1004_g Y 0.00652513f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_133 A2 Y 0.0202848f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_134 N_A2_c_142_n Y 5.97934e-19 $X=2.36 $Y=1.385 $X2=0 $Y2=0
cc_135 N_A2_M1004_g N_VPWR_c_313_n 0.00461464f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_136 N_A2_M1004_g N_VPWR_c_314_n 0.0093231f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A2_M1004_g N_VPWR_c_309_n 0.00460921f $X=2.405 $Y=2.4 $X2=0 $Y2=0
cc_138 A2 N_VGND_c_351_n 0.025354f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_139 N_A2_c_143_n N_VGND_c_351_n 0.00141413f $X=2.36 $Y=1.22 $X2=0 $Y2=0
cc_140 A2 N_VGND_c_352_n 0.0132057f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_141 N_A2_c_143_n N_VGND_c_352_n 0.00303293f $X=2.36 $Y=1.22 $X2=0 $Y2=0
cc_142 A2 N_VGND_c_353_n 0.0159188f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_143 N_A2_c_143_n N_VGND_c_353_n 0.00372643f $X=2.36 $Y=1.22 $X2=0 $Y2=0
cc_144 A2 A_391_74# 0.00780801f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_145 A2 A_469_74# 0.0100426f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_146 N_A3_M1007_g N_A_27_368#_c_210_n 0.00729209f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_147 A3 N_A_27_368#_c_210_n 0.00161008f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_148 N_A3_M1007_g N_A_27_368#_c_211_n 0.00682235f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_149 N_A3_M1007_g N_A_27_368#_c_228_n 0.00213632f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_150 N_A3_M1007_g N_VPWR_c_311_n 0.00517389f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_151 A3 N_VPWR_c_311_n 0.014999f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_152 N_A3_c_182_n N_VPWR_c_311_n 0.00218096f $X=2.93 $Y=1.385 $X2=0 $Y2=0
cc_153 N_A3_M1007_g N_VPWR_c_313_n 0.005209f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_154 N_A3_M1007_g N_VPWR_c_314_n 4.26462e-19 $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_155 N_A3_M1007_g N_VPWR_c_309_n 0.00986118f $X=2.855 $Y=2.4 $X2=0 $Y2=0
cc_156 A3 N_VGND_c_351_n 0.0259407f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_157 N_A3_c_182_n N_VGND_c_351_n 0.0011179f $X=2.93 $Y=1.385 $X2=0 $Y2=0
cc_158 N_A3_c_183_n N_VGND_c_351_n 0.0159756f $X=2.93 $Y=1.22 $X2=0 $Y2=0
cc_159 N_A3_c_183_n N_VGND_c_352_n 0.00383152f $X=2.93 $Y=1.22 $X2=0 $Y2=0
cc_160 N_A3_c_183_n N_VGND_c_353_n 0.00758792f $X=2.93 $Y=1.22 $X2=0 $Y2=0
cc_161 N_A_27_368#_c_208_n N_Y_M1003_d 0.00218982f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_162 N_A_27_368#_c_208_n N_Y_c_271_n 0.0177084f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_163 N_A_27_368#_c_207_n N_Y_c_261_n 0.00352479f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_164 N_A_27_368#_c_220_n Y 0.0073333f $X=1.28 $Y=2.49 $X2=0 $Y2=0
cc_165 N_A_27_368#_c_222_n Y 0.0470968f $X=2.465 $Y=2.405 $X2=0 $Y2=0
cc_166 N_A_27_368#_c_210_n Y 0.0121588f $X=2.63 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A_27_368#_M1002_d N_Y_c_263_n 0.00383831f $X=1.095 $Y=1.84 $X2=0 $Y2=0
cc_168 N_A_27_368#_c_220_n N_Y_c_263_n 0.0228277f $X=1.28 $Y=2.49 $X2=0 $Y2=0
cc_169 N_A_27_368#_c_222_n N_Y_c_263_n 0.00288953f $X=2.465 $Y=2.405 $X2=0 $Y2=0
cc_170 N_A_27_368#_c_222_n N_VPWR_M1006_d 0.0128113f $X=2.465 $Y=2.405 $X2=-0.19
+ $Y2=1.66
cc_171 N_A_27_368#_c_210_n N_VPWR_c_311_n 0.0171158f $X=2.63 $Y=1.985 $X2=0
+ $Y2=0
cc_172 N_A_27_368#_c_211_n N_VPWR_c_311_n 0.0163859f $X=2.63 $Y=2.815 $X2=0
+ $Y2=0
cc_173 N_A_27_368#_c_208_n N_VPWR_c_312_n 0.0658009f $X=1.115 $Y=2.99 $X2=0
+ $Y2=0
cc_174 N_A_27_368#_c_209_n N_VPWR_c_312_n 0.0235185f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_175 N_A_27_368#_c_211_n N_VPWR_c_313_n 0.0123179f $X=2.63 $Y=2.815 $X2=0
+ $Y2=0
cc_176 N_A_27_368#_c_208_n N_VPWR_c_314_n 0.011907f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_177 N_A_27_368#_c_221_n N_VPWR_c_314_n 0.0158718f $X=1.28 $Y=2.815 $X2=0
+ $Y2=0
cc_178 N_A_27_368#_c_222_n N_VPWR_c_314_n 0.0437071f $X=2.465 $Y=2.405 $X2=0
+ $Y2=0
cc_179 N_A_27_368#_c_211_n N_VPWR_c_314_n 0.0141508f $X=2.63 $Y=2.815 $X2=0
+ $Y2=0
cc_180 N_A_27_368#_c_208_n N_VPWR_c_309_n 0.036511f $X=1.115 $Y=2.99 $X2=0 $Y2=0
cc_181 N_A_27_368#_c_209_n N_VPWR_c_309_n 0.0126877f $X=0.445 $Y=2.99 $X2=0
+ $Y2=0
cc_182 N_A_27_368#_c_222_n N_VPWR_c_309_n 0.0123109f $X=2.465 $Y=2.405 $X2=0
+ $Y2=0
cc_183 N_A_27_368#_c_211_n N_VPWR_c_309_n 0.0101276f $X=2.63 $Y=2.815 $X2=0
+ $Y2=0
cc_184 N_A_27_368#_c_228_n N_VPWR_c_309_n 0.00170101f $X=2.63 $Y=2.405 $X2=0
+ $Y2=0
cc_185 Y N_VPWR_M1006_d 0.0117635f $X=2.075 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_186 N_Y_c_258_n N_VGND_c_349_n 0.0284176f $X=0.785 $Y=0.68 $X2=0 $Y2=0
cc_187 N_Y_c_258_n N_VGND_c_352_n 0.00758556f $X=0.785 $Y=0.68 $X2=0 $Y2=0
cc_188 N_Y_c_259_n N_VGND_c_352_n 0.0457898f $X=1.665 $Y=0.495 $X2=0 $Y2=0
cc_189 N_Y_c_258_n N_VGND_c_353_n 0.00627867f $X=0.785 $Y=0.68 $X2=0 $Y2=0
cc_190 N_Y_c_259_n N_VGND_c_353_n 0.037678f $X=1.665 $Y=0.495 $X2=0 $Y2=0

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a32oi_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 VPWR A2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 a_27_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 a_1313_74# A2 a_868_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VPWR A3 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X4 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_27_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X6 VPWR A3 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 a_27_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 Y B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X9 a_27_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X10 a_27_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X11 a_27_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X12 a_27_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X13 a_868_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 Y A1 a_868_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 a_27_368# B1 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X16 VGND B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 VPWR A1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X18 VPWR A1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X19 a_1313_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 a_27_368# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X21 Y A1 a_868_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 a_1313_74# A2 a_868_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 Y B1 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 a_1313_74# A3 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 a_27_368# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X26 VPWR A2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X27 Y B1 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X28 VGND B2 a_27_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X29 a_868_74# A2 a_1313_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X30 a_868_74# A2 a_1313_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X31 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X32 a_27_74# B1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X33 VGND A3 a_1313_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X34 Y B2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X35 Y B2 a_27_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X36 a_27_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X37 a_868_74# A1 Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X38 a_27_368# A3 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X39 VGND A3 a_1313_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

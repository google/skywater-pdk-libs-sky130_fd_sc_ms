* NGSPICE file created from sky130_fd_sc_ms__dlrtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__dlrtp_2 D GATE RESET_B VGND VNB VPB VPWR Q
M1000 a_759_508# a_347_98# a_646_74# VPB pshort w=420000u l=180000u
+  ad=2.121e+11p pd=1.85e+06u as=3.115e+11p ps=2.71e+06u
M1001 VGND a_235_74# a_347_98# VNB nlowvt w=740000u l=150000u
+  ad=1.38725e+12p pd=1.126e+07u as=2.701e+11p ps=2.21e+06u
M1002 VPWR D a_27_392# VPB pshort w=840000u l=180000u
+  ad=2.11845e+12p pd=1.561e+07u as=2.352e+11p ps=2.24e+06u
M1003 a_568_74# a_27_392# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1004 a_646_74# a_347_98# a_568_74# VNB nlowvt w=640000u l=150000u
+  ad=3.21575e+11p pd=2.36e+06u as=0p ps=0u
M1005 VGND RESET_B a_1060_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.776e+11p ps=1.96e+06u
M1006 Q a_832_55# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.146e+11p pd=2.06e+06u as=0p ps=0u
M1007 VPWR a_235_74# a_347_98# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1008 Q a_832_55# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.192e+11p pd=2.81e+06u as=0p ps=0u
M1009 a_832_55# a_646_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1010 VPWR RESET_B a_832_55# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_832_55# a_759_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND D a_27_392# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1013 VPWR a_832_55# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_568_392# a_27_392# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1015 a_235_74# GATE VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1016 a_646_74# a_235_74# a_568_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1060_74# a_646_74# a_832_55# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1018 VGND a_832_55# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_784_81# a_235_74# a_646_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1020 VGND a_832_55# a_784_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_235_74# GATE VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
.ends


* File: sky130_fd_sc_ms__dfrtp_4.pex.spice
* Created: Fri Aug 28 17:23:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DFRTP_4%D 2 4 7 11 13 14 15 16 21 22 25
r36 25 27 35.4289 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.42 $Y=1.845
+ $X2=0.42 $Y2=2.01
r37 25 26 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.845 $X2=0.385 $Y2=1.845
r38 21 23 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.42 $Y=1.165
+ $X2=0.42 $Y2=1
r39 21 22 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.165 $X2=0.385 $Y2=1.165
r40 16 26 5.61447 $w=3.88e-07 $l=1.9e-07 $layer=LI1_cond $X=0.32 $Y=2.035
+ $X2=0.32 $Y2=1.845
r41 15 26 5.31897 $w=3.88e-07 $l=1.8e-07 $layer=LI1_cond $X=0.32 $Y=1.665
+ $X2=0.32 $Y2=1.845
r42 14 15 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.32 $Y=1.295
+ $X2=0.32 $Y2=1.665
r43 14 22 3.84148 $w=3.88e-07 $l=1.3e-07 $layer=LI1_cond $X=0.32 $Y=1.295
+ $X2=0.32 $Y2=1.165
r44 11 23 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.545 $Y=0.6 $X2=0.545
+ $Y2=1
r45 7 13 155.484 $w=1.8e-07 $l=4e-07 $layer=POLY_cond $X=0.5 $Y=2.75 $X2=0.5
+ $Y2=2.35
r46 4 13 34.6974 $w=2.1e-07 $l=1.05e-07 $layer=POLY_cond $X=0.515 $Y=2.245
+ $X2=0.515 $Y2=2.35
r47 4 27 74.2101 $w=2.1e-07 $l=2.35e-07 $layer=POLY_cond $X=0.515 $Y=2.245
+ $X2=0.515 $Y2=2.01
r48 2 25 4.86635 $w=4e-07 $l=3.5e-08 $layer=POLY_cond $X=0.42 $Y=1.81 $X2=0.42
+ $Y2=1.845
r49 1 21 4.86635 $w=4e-07 $l=3.5e-08 $layer=POLY_cond $X=0.42 $Y=1.2 $X2=0.42
+ $Y2=1.165
r50 1 2 84.8135 $w=4e-07 $l=6.1e-07 $layer=POLY_cond $X=0.42 $Y=1.2 $X2=0.42
+ $Y2=1.81
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_4%CLK 3 6 7 10 12 13
c47 7 0 1.60579e-19 $X=2.16 $Y=1.665
r48 10 13 59.925 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=1.93 $Y=1.61
+ $X2=1.93 $Y2=1.885
r49 10 12 52.3316 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=1.93 $Y=1.61 $X2=1.93
+ $Y2=1.41
r50 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.93
+ $Y=1.61 $X2=1.93 $Y2=1.61
r51 7 11 6.00857 $w=4.67e-07 $l=2.3e-07 $layer=LI1_cond $X=2.16 $Y=1.545
+ $X2=1.93 $Y2=1.545
r52 6 12 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.95 $Y=0.965
+ $X2=1.95 $Y2=1.41
r53 3 13 174.056 $w=1.8e-07 $l=6.5e-07 $layer=POLY_cond $X=1.945 $Y=2.535
+ $X2=1.945 $Y2=1.885
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_4%A_497_395# 1 2 7 9 11 13 15 17 19 20 21 24
+ 27 32 33 35 37 41 45 46 52 55 59 65 68 78
c198 52 0 1.60579e-19 $X=3.355 $Y=1.725
c199 46 0 1.63369e-19 $X=2.78 $Y=0.415
c200 41 0 9.26151e-20 $X=7.905 $Y=2.14
c201 33 0 1.29851e-19 $X=4.305 $Y=0.415
c202 15 0 1.85309e-19 $X=3.985 $Y=0.9
c203 13 0 3.29442e-19 $X=3.985 $Y=1.385
c204 7 0 1.00854e-19 $X=3.42 $Y=1.89
r205 67 68 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=7.905 $Y=1.18
+ $X2=8.19 $Y2=1.18
r206 65 74 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.71 $Y=1.18 $X2=7.71
+ $Y2=1.27
r207 64 67 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=7.71 $Y=1.18
+ $X2=7.905 $Y2=1.18
r208 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.71
+ $Y=1.18 $X2=7.71 $Y2=1.18
r209 59 61 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.48 $Y=0.34
+ $X2=5.48 $Y2=0.625
r210 55 57 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.39 $Y=0.415
+ $X2=4.39 $Y2=0.625
r211 53 70 8.81707 $w=3.28e-07 $l=6e-08 $layer=POLY_cond $X=3.355 $Y=1.725
+ $X2=3.355 $Y2=1.665
r212 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.355
+ $Y=1.725 $X2=3.355 $Y2=1.725
r213 49 50 7.30169 $w=4.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=0.72
+ $X2=2.78 $Y2=0.805
r214 46 49 7.76179 $w=4.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.78 $Y=0.415
+ $X2=2.78 $Y2=0.72
r215 45 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.19 $Y=1.015
+ $X2=8.19 $Y2=1.18
r216 44 45 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.19 $Y=0.425
+ $X2=8.19 $Y2=1.015
r217 42 78 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=7.905 $Y=2.14
+ $X2=8.06 $Y2=2.14
r218 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.905
+ $Y=2.14 $X2=7.905 $Y2=2.14
r219 39 67 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=7.905 $Y=1.345
+ $X2=7.905 $Y2=1.18
r220 39 41 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=7.905 $Y=1.345
+ $X2=7.905 $Y2=2.14
r221 38 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=0.34
+ $X2=5.48 $Y2=0.34
r222 37 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.105 $Y=0.34
+ $X2=8.19 $Y2=0.425
r223 37 38 165.711 $w=1.68e-07 $l=2.54e-06 $layer=LI1_cond $X=8.105 $Y=0.34
+ $X2=5.565 $Y2=0.34
r224 36 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.475 $Y=0.625
+ $X2=4.39 $Y2=0.625
r225 35 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=0.625
+ $X2=5.48 $Y2=0.625
r226 35 36 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=5.395 $Y=0.625
+ $X2=4.475 $Y2=0.625
r227 34 46 6.76998 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.015 $Y=0.415
+ $X2=2.78 $Y2=0.415
r228 33 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.305 $Y=0.415
+ $X2=4.39 $Y2=0.415
r229 33 34 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=4.305 $Y=0.415
+ $X2=3.015 $Y2=0.415
r230 32 52 9.25877 $w=4.22e-07 $l=2.91033e-07 $layer=LI1_cond $X=2.93 $Y=1.56
+ $X2=3.15 $Y2=1.725
r231 32 50 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.93 $Y=1.56
+ $X2=2.93 $Y2=0.805
r232 27 52 10.3209 $w=4.22e-07 $l=4.86142e-07 $layer=LI1_cond $X=2.845 $Y=2.082
+ $X2=3.15 $Y2=1.725
r233 27 29 9.42908 $w=2.73e-07 $l=2.25e-07 $layer=LI1_cond $X=2.845 $Y=2.082
+ $X2=2.62 $Y2=2.082
r234 22 78 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.06 $Y=2.305
+ $X2=8.06 $Y2=2.14
r235 22 24 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=8.06 $Y=2.305
+ $X2=8.06 $Y2=2.675
r236 20 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.545 $Y=1.27
+ $X2=7.71 $Y2=1.27
r237 20 21 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=7.545 $Y=1.27
+ $X2=7.185 $Y2=1.27
r238 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.11 $Y=1.195
+ $X2=7.185 $Y2=1.27
r239 17 19 146.207 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=7.11 $Y=1.195
+ $X2=7.11 $Y2=0.74
r240 13 26 71.6325 $w=1.96e-07 $l=3.06268e-07 $layer=POLY_cond $X=3.985 $Y=1.385
+ $X2=3.93 $Y2=1.665
r241 13 15 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=3.985 $Y=1.385
+ $X2=3.985 $Y2=0.9
r242 12 70 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.52 $Y=1.665
+ $X2=3.355 $Y2=1.665
r243 11 26 9.11062 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=3.8 $Y=1.665
+ $X2=3.93 $Y2=1.665
r244 11 12 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.8 $Y=1.665
+ $X2=3.52 $Y2=1.665
r245 7 53 33.9886 $w=3.28e-07 $l=1.94808e-07 $layer=POLY_cond $X=3.42 $Y=1.89
+ $X2=3.355 $Y2=1.725
r246 7 9 246.831 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=3.42 $Y=1.89
+ $X2=3.42 $Y2=2.525
r247 2 29 600 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=1 $X=2.485
+ $Y=1.975 $X2=2.62 $Y2=2.135
r248 1 49 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=2.545
+ $Y=0.595 $X2=2.71 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_4%A_834_355# 1 2 9 13 17 18 21 23 24 26 30 35
c90 35 0 1.49998e-19 $X=6.45 $Y=2.125
c91 30 0 1.42689e-20 $X=5.735 $Y=0.885
c92 24 0 5.02509e-20 $X=6.325 $Y=0.885
c93 21 0 3.05298e-19 $X=4.57 $Y=0.965
c94 13 0 1.36289e-19 $X=4.375 $Y=0.9
r95 29 31 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=5.9 $Y=0.885
+ $X2=6.24 $Y2=0.885
r96 29 30 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.9 $Y=0.885
+ $X2=5.735 $Y2=0.885
r97 24 31 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=6.325 $Y=0.885
+ $X2=6.24 $Y2=0.885
r98 24 26 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=6.325 $Y=0.885
+ $X2=6.825 $Y2=0.885
r99 23 35 8.20383 $w=2.93e-07 $l=2.1e-07 $layer=LI1_cond $X=6.24 $Y=2.087
+ $X2=6.45 $Y2=2.087
r100 22 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.24 $Y=1.05
+ $X2=6.24 $Y2=0.885
r101 22 23 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=6.24 $Y=1.05
+ $X2=6.24 $Y2=1.94
r102 21 30 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=4.57 $Y=0.965
+ $X2=5.735 $Y2=0.965
r103 18 39 39.9775 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=1.94
+ $X2=4.37 $Y2=2.105
r104 18 38 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=1.94
+ $X2=4.37 $Y2=1.775
r105 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.405
+ $Y=1.94 $X2=4.405 $Y2=1.94
r106 15 21 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=4.437 $Y=1.05
+ $X2=4.57 $Y2=0.965
r107 15 17 38.7047 $w=2.63e-07 $l=8.9e-07 $layer=LI1_cond $X=4.437 $Y=1.05
+ $X2=4.437 $Y2=1.94
r108 13 38 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=4.375 $Y=0.9
+ $X2=4.375 $Y2=1.775
r109 9 39 163.258 $w=1.8e-07 $l=4.2e-07 $layer=POLY_cond $X=4.26 $Y=2.525
+ $X2=4.26 $Y2=2.105
r110 2 35 600 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=6.315
+ $Y=1.96 $X2=6.45 $Y2=2.125
r111 1 29 182 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_NDIFF $count=1 $X=5.76
+ $Y=0.37 $X2=5.9 $Y2=0.885
r112 1 26 91 $w=1.7e-07 $l=1.29719e-06 $layer=licon1_NDIFF $count=2 $X=5.76
+ $Y=0.37 $X2=6.825 $Y2=0.885
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_4%RESET_B 4 6 9 11 12 16 19 22 25 29 33 36 37
+ 38 39 40 43 45 46 48 51 55 56 59 63
c230 55 0 1.15254e-19 $X=1.155 $Y=1.295
c231 51 0 1.66354e-20 $X=5.25 $Y=1.835
c232 43 0 1.36553e-19 $X=5.52 $Y=2.035
c233 40 0 1.63054e-19 $X=5.665 $Y=2.035
c234 36 0 1.42689e-20 $X=4.87 $Y=1.835
c235 19 0 1.24602e-19 $X=4.87 $Y=2.525
c236 11 0 1.19989e-19 $X=4.69 $Y=0.18
r237 63 66 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.975 $Y=2.11
+ $X2=8.975 $Y2=2.275
r238 63 65 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.975 $Y=2.11
+ $X2=8.975 $Y2=1.945
r239 59 61 41.3282 $w=4.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.975
+ $X2=1.09 $Y2=2.14
r240 59 60 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.975 $X2=1.155 $Y2=1.975
r241 56 60 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.155 $Y=1.295
+ $X2=1.155 $Y2=1.975
r242 55 57 47.2161 $w=4.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.295
+ $X2=1.09 $Y2=1.13
r243 55 56 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.295 $X2=1.155 $Y2=1.295
r244 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.25
+ $Y=1.835 $X2=5.25 $Y2=1.835
r245 48 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.035
+ $X2=1.2 $Y2=2.035
r246 46 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.975
+ $Y=2.11 $X2=8.975 $Y2=2.11
r247 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=2.035
+ $X2=8.88 $Y2=2.035
r248 43 52 7.17647 $w=4.48e-07 $l=2.7e-07 $layer=LI1_cond $X=5.52 $Y=1.895
+ $X2=5.25 $Y2=1.895
r249 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=2.035
+ $X2=5.52 $Y2=2.035
r250 40 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=2.035
+ $X2=5.52 $Y2=2.035
r251 39 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.735 $Y=2.035
+ $X2=8.88 $Y2=2.035
r252 39 40 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=8.735 $Y=2.035
+ $X2=5.665 $Y2=2.035
r253 38 48 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=2.035
+ $X2=1.2 $Y2=2.035
r254 37 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=2.035
+ $X2=5.52 $Y2=2.035
r255 37 38 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=5.375 $Y=2.035
+ $X2=1.345 $Y2=2.035
r256 35 51 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=4.96 $Y=1.835
+ $X2=5.25 $Y2=1.835
r257 35 36 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.96 $Y=1.835
+ $X2=4.87 $Y2=1.835
r258 31 33 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=4.765 $Y=1.26
+ $X2=4.885 $Y2=1.26
r259 29 65 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=9.06 $Y=0.615
+ $X2=9.06 $Y2=1.945
r260 25 66 155.484 $w=1.8e-07 $l=4e-07 $layer=POLY_cond $X=9.02 $Y=2.675
+ $X2=9.02 $Y2=2.275
r261 22 36 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=4.885 $Y=1.67
+ $X2=4.87 $Y2=1.835
r262 21 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.885 $Y=1.335
+ $X2=4.885 $Y2=1.26
r263 21 22 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=4.885 $Y=1.335
+ $X2=4.885 $Y2=1.67
r264 17 36 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=4.87 $Y=2
+ $X2=4.87 $Y2=1.835
r265 17 19 204.073 $w=1.8e-07 $l=5.25e-07 $layer=POLY_cond $X=4.87 $Y=2 $X2=4.87
+ $Y2=2.525
r266 14 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.765 $Y=1.185
+ $X2=4.765 $Y2=1.26
r267 14 16 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.765 $Y=1.185
+ $X2=4.765 $Y2=0.9
r268 13 16 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=4.765 $Y=0.255
+ $X2=4.765 $Y2=0.9
r269 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.69 $Y=0.18
+ $X2=4.765 $Y2=0.255
r270 11 12 1886.98 $w=1.5e-07 $l=3.68e-06 $layer=POLY_cond $X=4.69 $Y=0.18
+ $X2=1.01 $Y2=0.18
r271 9 61 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=0.95 $Y=2.75
+ $X2=0.95 $Y2=2.14
r272 6 59 7.8587 $w=4.6e-07 $l=6.5e-08 $layer=POLY_cond $X=1.09 $Y=1.91 $X2=1.09
+ $Y2=1.975
r273 5 55 7.8587 $w=4.6e-07 $l=6.5e-08 $layer=POLY_cond $X=1.09 $Y=1.36 $X2=1.09
+ $Y2=1.295
r274 5 6 66.4967 $w=4.6e-07 $l=5.5e-07 $layer=POLY_cond $X=1.09 $Y=1.36 $X2=1.09
+ $Y2=1.91
r275 4 57 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.935 $Y=0.6
+ $X2=0.935 $Y2=1.13
r276 1 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.935 $Y=0.255
+ $X2=1.01 $Y2=0.18
r277 1 4 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=0.935 $Y=0.255
+ $X2=0.935 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_4%A_303_395# 1 2 7 9 10 12 14 15 16 17 18 19
+ 21 24 26 29 30 32 34 38 40 43 47 50 51 54 55 57 58 64 65 73
c226 65 0 1.73349e-19 $X=5.56 $Y=2.375
c227 64 0 2.80152e-19 $X=5.56 $Y=2.375
c228 55 0 1.15254e-19 $X=1.665 $Y=1.055
c229 54 0 1.35587e-19 $X=6.87 $Y=2.405
c230 50 0 1.00854e-19 $X=2.56 $Y=1.435
c231 43 0 1.63369e-19 $X=1.69 $Y=0.715
c232 24 0 1.93874e-19 $X=3.87 $Y=2.525
c233 17 0 9.3565e-20 $X=3.41 $Y=1.26
r234 71 84 37.5066 $w=3.02e-07 $l=2.35e-07 $layer=POLY_cond $X=6.66 $Y=1.425
+ $X2=6.66 $Y2=1.66
r235 70 73 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=6.66 $Y=1.425
+ $X2=6.87 $Y2=1.425
r236 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.66
+ $Y=1.425 $X2=6.66 $Y2=1.425
r237 65 79 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=5.56 $Y=2.375
+ $X2=5.385 $Y2=2.375
r238 64 67 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=5.56 $Y=2.375
+ $X2=5.56 $Y2=2.49
r239 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.56
+ $Y=2.375 $X2=5.56 $Y2=2.375
r240 62 78 33.258 $w=5e-07 $l=3.45e-07 $layer=POLY_cond $X=2.56 $Y=1.535
+ $X2=2.905 $Y2=1.535
r241 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.56
+ $Y=1.61 $X2=2.56 $Y2=1.61
r242 57 58 9.31166 $w=3.48e-07 $l=1.9e-07 $layer=LI1_cond $X=1.63 $Y=2.135
+ $X2=1.63 $Y2=1.945
r243 53 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.87 $Y=1.59
+ $X2=6.87 $Y2=1.425
r244 53 54 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=6.87 $Y=1.59
+ $X2=6.87 $Y2=2.405
r245 52 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.725 $Y=2.49
+ $X2=5.56 $Y2=2.49
r246 51 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.785 $Y=2.49
+ $X2=6.87 $Y2=2.405
r247 51 52 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=6.785 $Y=2.49
+ $X2=5.725 $Y2=2.49
r248 50 61 9.28261 $w=2.3e-07 $l=1.75e-07 $layer=LI1_cond $X=2.56 $Y=1.435
+ $X2=2.56 $Y2=1.61
r249 49 50 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.56 $Y=1.14
+ $X2=2.56 $Y2=1.435
r250 48 55 3.3845 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=1.875 $Y=1.055
+ $X2=1.665 $Y2=1.055
r251 47 49 9.71848 $w=1.44e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.445 $Y=1.055
+ $X2=2.56 $Y2=1.14
r252 47 48 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.445 $Y=1.055
+ $X2=1.875 $Y2=1.055
r253 45 55 3.19717 $w=2.95e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.54 $Y=1.14
+ $X2=1.665 $Y2=1.055
r254 45 58 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.54 $Y=1.14
+ $X2=1.54 $Y2=1.945
r255 41 55 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=0.97
+ $X2=1.665 $Y2=1.055
r256 41 43 6.99698 $w=4.18e-07 $l=2.55e-07 $layer=LI1_cond $X=1.665 $Y=0.97
+ $X2=1.665 $Y2=0.715
r257 36 38 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=8.16 $Y=1.585
+ $X2=8.16 $Y2=0.615
r258 35 84 19.1248 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.825 $Y=1.66
+ $X2=6.66 $Y2=1.66
r259 34 36 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.085 $Y=1.66
+ $X2=8.16 $Y2=1.585
r260 34 35 646.085 $w=1.5e-07 $l=1.26e-06 $layer=POLY_cond $X=8.085 $Y=1.66
+ $X2=6.825 $Y2=1.66
r261 30 84 19.7735 $w=3.02e-07 $l=8.21584e-08 $layer=POLY_cond $X=6.675 $Y=1.735
+ $X2=6.66 $Y2=1.66
r262 30 32 281.815 $w=1.8e-07 $l=7.25e-07 $layer=POLY_cond $X=6.675 $Y=1.735
+ $X2=6.675 $Y2=2.46
r263 28 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.385 $Y=2.54
+ $X2=5.385 $Y2=2.375
r264 28 29 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=5.385 $Y=2.54
+ $X2=5.385 $Y2=3.075
r265 27 40 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.96 $Y=3.15 $X2=3.87
+ $Y2=3.15
r266 26 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.31 $Y=3.15
+ $X2=5.385 $Y2=3.075
r267 26 27 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=5.31 $Y=3.15
+ $X2=3.96 $Y2=3.15
r268 22 40 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.87 $Y=3.075
+ $X2=3.87 $Y2=3.15
r269 22 24 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=3.87 $Y=3.075
+ $X2=3.87 $Y2=2.525
r270 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.485 $Y=1.185
+ $X2=3.485 $Y2=0.9
r271 18 78 37.1056 $w=5e-07 $l=3.2749e-07 $layer=POLY_cond $X=3.02 $Y=1.26
+ $X2=2.905 $Y2=1.535
r272 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.41 $Y=1.26
+ $X2=3.485 $Y2=1.185
r273 17 18 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.41 $Y=1.26
+ $X2=3.02 $Y2=1.26
r274 15 40 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.78 $Y=3.15 $X2=3.87
+ $Y2=3.15
r275 15 16 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.78 $Y=3.15 $X2=2.98
+ $Y2=3.15
r276 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.905 $Y=3.075
+ $X2=2.98 $Y2=3.15
r277 13 78 31.4081 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.905 $Y=1.885
+ $X2=2.905 $Y2=1.535
r278 13 14 610.191 $w=1.5e-07 $l=1.19e-06 $layer=POLY_cond $X=2.905 $Y=1.885
+ $X2=2.905 $Y2=3.075
r279 10 62 8.676 $w=5e-07 $l=9e-08 $layer=POLY_cond $X=2.47 $Y=1.535 $X2=2.56
+ $Y2=1.535
r280 10 75 7.23 $w=5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.47 $Y=1.535 $X2=2.395
+ $Y2=1.535
r281 10 12 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.47 $Y=1.41
+ $X2=2.47 $Y2=0.965
r282 7 75 26.863 $w=1.8e-07 $l=3.5e-07 $layer=POLY_cond $X=2.395 $Y=1.885
+ $X2=2.395 $Y2=1.535
r283 7 9 174.056 $w=1.8e-07 $l=6.5e-07 $layer=POLY_cond $X=2.395 $Y=1.885
+ $X2=2.395 $Y2=2.535
r284 2 57 600 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_PDIFF $count=1 $X=1.515
+ $Y=1.975 $X2=1.64 $Y2=2.135
r285 1 43 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.545
+ $Y=0.59 $X2=1.69 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_4%A_702_463# 1 2 3 10 12 15 17 19 20 21 27 28
+ 31 32 34 38 41 42 43
c138 31 0 1.38915e-19 $X=4.83 $Y=2.295
c139 27 0 9.3565e-20 $X=4.05 $Y=2.4
c140 21 0 1.30745e-19 $X=6.225 $Y=1.73
c141 19 0 2.99607e-19 $X=5.76 $Y=1.385
c142 15 0 5.50928e-20 $X=6.225 $Y=1.82
r143 43 45 8.354 $w=3.87e-07 $l=2.65e-07 $layer=LI1_cond $X=4.83 $Y=2.525
+ $X2=5.095 $Y2=2.525
r144 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.82
+ $Y=1.385 $X2=5.82 $Y2=1.385
r145 32 34 37.2486 $w=2.78e-07 $l=9.05e-07 $layer=LI1_cond $X=4.915 $Y=1.36
+ $X2=5.82 $Y2=1.36
r146 31 43 5.57805 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=4.83 $Y=2.295
+ $X2=4.83 $Y2=2.525
r147 30 32 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=4.83 $Y=1.5
+ $X2=4.915 $Y2=1.36
r148 30 31 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=4.83 $Y=1.5
+ $X2=4.83 $Y2=2.295
r149 28 43 6.57826 $w=3.87e-07 $l=1.03078e-07 $layer=LI1_cond $X=4.745 $Y=2.485
+ $X2=4.83 $Y2=2.525
r150 28 42 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=4.745 $Y=2.485
+ $X2=4.23 $Y2=2.485
r151 27 42 9.01544 $w=3.73e-07 $l=1.8e-07 $layer=LI1_cond $X=4.05 $Y=2.587
+ $X2=4.23 $Y2=2.587
r152 27 41 2.80732 $w=3.73e-07 $l=8.5e-08 $layer=LI1_cond $X=4.05 $Y=2.587
+ $X2=3.965 $Y2=2.587
r153 26 38 11.3867 $w=3e-07 $l=3.62767e-07 $layer=LI1_cond $X=4.05 $Y=1.05
+ $X2=3.77 $Y2=0.86
r154 26 27 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=4.05 $Y=1.05
+ $X2=4.05 $Y2=2.4
r155 24 41 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=3.645 $Y=2.61
+ $X2=3.965 $Y2=2.61
r156 20 35 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=6.135 $Y=1.385
+ $X2=5.82 $Y2=1.385
r157 19 35 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=5.76 $Y=1.385
+ $X2=5.82 $Y2=1.385
r158 15 21 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.225 $Y=1.82
+ $X2=6.225 $Y2=1.73
r159 15 17 248.774 $w=1.8e-07 $l=6.4e-07 $layer=POLY_cond $X=6.225 $Y=1.82
+ $X2=6.225 $Y2=2.46
r160 13 20 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=6.21 $Y=1.55
+ $X2=6.135 $Y2=1.385
r161 13 21 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=6.21 $Y=1.55
+ $X2=6.21 $Y2=1.73
r162 10 19 17.4878 $w=4.41e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.685 $Y=1.22
+ $X2=5.76 $Y2=1.385
r163 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.685 $Y=1.22
+ $X2=5.685 $Y2=0.74
r164 3 45 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=4.96
+ $Y=2.315 $X2=5.095 $Y2=2.525
r165 2 24 600 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_PDIFF $count=1 $X=3.51
+ $Y=2.315 $X2=3.645 $Y2=2.61
r166 1 38 182 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.69 $X2=3.77 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_4%A_1678_395# 1 2 9 15 17 18 19 22 23 24 27 30
+ 31 35 40 42
c122 40 0 1.63846e-19 $X=9.395 $Y=2.675
c123 30 0 1.27304e-19 $X=9.86 $Y=1.875
c124 23 0 1.26767e-19 $X=9.775 $Y=1.96
c125 17 0 9.26151e-20 $X=8.492 $Y=1.975
r126 38 40 3.90026 $w=4.58e-07 $l=1.5e-07 $layer=LI1_cond $X=9.245 $Y=2.675
+ $X2=9.395 $Y2=2.675
r127 35 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.61 $Y=1.2
+ $X2=8.61 $Y2=1.365
r128 35 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.61 $Y=1.2
+ $X2=8.61 $Y2=1.035
r129 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.61
+ $Y=1.2 $X2=8.61 $Y2=1.2
r130 31 34 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=8.61 $Y=1.12 $X2=8.61
+ $Y2=1.2
r131 29 42 3.70735 $w=2.5e-07 $l=1.75425e-07 $layer=LI1_cond $X=9.86 $Y=1.205
+ $X2=9.722 $Y2=1.12
r132 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.86 $Y=1.205
+ $X2=9.86 $Y2=1.875
r133 25 42 3.70735 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.665 $Y=1.035
+ $X2=9.722 $Y2=1.12
r134 25 27 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=9.665 $Y=1.035
+ $X2=9.665 $Y2=0.615
r135 23 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.775 $Y=1.96
+ $X2=9.86 $Y2=1.875
r136 23 24 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.775 $Y=1.96
+ $X2=9.48 $Y2=1.96
r137 22 40 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=9.395 $Y=2.445
+ $X2=9.395 $Y2=2.675
r138 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.395 $Y=2.045
+ $X2=9.48 $Y2=1.96
r139 21 22 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=9.395 $Y=2.045
+ $X2=9.395 $Y2=2.445
r140 20 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.775 $Y=1.12
+ $X2=8.61 $Y2=1.12
r141 19 42 2.76166 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=9.5 $Y=1.12
+ $X2=9.722 $Y2=1.12
r142 19 20 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=9.5 $Y=1.12
+ $X2=8.775 $Y2=1.12
r143 17 18 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=8.492 $Y=1.975
+ $X2=8.492 $Y2=2.125
r144 17 45 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.52 $Y=1.975
+ $X2=8.52 $Y2=1.365
r145 15 44 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=8.55 $Y=0.615
+ $X2=8.55 $Y2=1.035
r146 9 18 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=8.48 $Y=2.675
+ $X2=8.48 $Y2=2.125
r147 2 38 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=9.11
+ $Y=2.465 $X2=9.245 $Y2=2.675
r148 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.525
+ $Y=0.405 $X2=9.665 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_4%A_1353_392# 1 2 9 13 15 19 21 25 28 31 32 33
+ 34 35 36 37 40 42 47 48 49 55 56
c163 47 0 9.99956e-20 $X=8.325 $Y=2.475
c164 35 0 1.07146e-19 $X=10.475 $Y=1.335
c165 25 0 2.54071e-19 $X=10.425 $Y=2.465
c166 19 0 1.63846e-19 $X=9.975 $Y=2.465
r167 62 63 24.9528 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.51 $Y=1.63
+ $X2=9.51 $Y2=1.705
r168 56 62 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.51 $Y=1.54 $X2=9.51
+ $Y2=1.63
r169 56 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.51 $Y=1.54
+ $X2=9.51 $Y2=1.375
r170 55 58 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=9.475 $Y=1.54
+ $X2=9.475 $Y2=1.62
r171 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.51
+ $Y=1.54 $X2=9.51 $Y2=1.54
r172 48 58 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.345 $Y=1.62
+ $X2=9.475 $Y2=1.62
r173 48 49 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=9.345 $Y=1.62 $X2=8.41
+ $Y2=1.62
r174 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.325 $Y=1.705
+ $X2=8.41 $Y2=1.62
r175 46 47 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=8.325 $Y=1.705
+ $X2=8.325 $Y2=2.475
r176 43 51 2.79691 $w=3.3e-07 $l=1.03e-07 $layer=LI1_cond $X=7.33 $Y=2.64
+ $X2=7.227 $Y2=2.64
r177 43 45 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=7.33 $Y=2.64
+ $X2=7.835 $Y2=2.64
r178 42 47 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.24 $Y=2.64
+ $X2=8.325 $Y2=2.475
r179 42 45 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=8.24 $Y=2.64
+ $X2=7.835 $Y2=2.64
r180 38 53 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.33 $Y=0.72
+ $X2=7.245 $Y2=0.72
r181 38 40 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=7.33 $Y=0.72
+ $X2=7.77 $Y2=0.72
r182 37 51 4.96927 $w=1.7e-07 $l=1.73767e-07 $layer=LI1_cond $X=7.245 $Y=2.475
+ $X2=7.227 $Y2=2.64
r183 36 53 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.245 $Y=0.845
+ $X2=7.245 $Y2=0.72
r184 36 37 106.342 $w=1.68e-07 $l=1.63e-06 $layer=LI1_cond $X=7.245 $Y=0.845
+ $X2=7.245 $Y2=2.475
r185 34 35 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=10.475 $Y=1.185
+ $X2=10.475 $Y2=1.335
r186 31 34 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=10.51 $Y=0.74
+ $X2=10.51 $Y2=1.185
r187 28 33 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=10.44 $Y=1.555
+ $X2=10.425 $Y2=1.63
r188 28 35 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=10.44 $Y=1.555
+ $X2=10.44 $Y2=1.335
r189 23 33 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=10.425 $Y=1.705
+ $X2=10.425 $Y2=1.63
r190 23 25 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=10.425 $Y=1.705
+ $X2=10.425 $Y2=2.465
r191 22 32 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=10.065 $Y=1.63
+ $X2=9.975 $Y2=1.63
r192 21 33 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=10.335 $Y=1.63
+ $X2=10.425 $Y2=1.63
r193 21 22 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=10.335 $Y=1.63
+ $X2=10.065 $Y2=1.63
r194 17 32 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.975 $Y=1.705
+ $X2=9.975 $Y2=1.63
r195 17 19 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=9.975 $Y=1.705
+ $X2=9.975 $Y2=2.465
r196 16 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.675 $Y=1.63
+ $X2=9.51 $Y2=1.63
r197 15 32 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.885 $Y=1.63
+ $X2=9.975 $Y2=1.63
r198 15 16 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=9.885 $Y=1.63
+ $X2=9.675 $Y2=1.63
r199 13 63 377.048 $w=1.8e-07 $l=9.7e-07 $layer=POLY_cond $X=9.47 $Y=2.675
+ $X2=9.47 $Y2=1.705
r200 9 61 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=9.45 $Y=0.615
+ $X2=9.45 $Y2=1.375
r201 2 51 600 $w=1.7e-07 $l=8.88144e-07 $layer=licon1_PDIFF $count=1 $X=6.765
+ $Y=1.96 $X2=7.245 $Y2=2.64
r202 2 45 600 $w=1.7e-07 $l=1.36839e-06 $layer=licon1_PDIFF $count=1 $X=6.765
+ $Y=1.96 $X2=7.835 $Y2=2.64
r203 1 53 182 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_NDIFF $count=1 $X=7.185
+ $Y=0.37 $X2=7.325 $Y2=0.68
r204 1 40 182 $w=1.7e-07 $l=7.23585e-07 $layer=licon1_NDIFF $count=1 $X=7.185
+ $Y=0.37 $X2=7.77 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_4%A_2013_409# 1 2 9 12 15 19 21 22 25 29 33 37
+ 41 45 47 48 51 58 61 63 70
c126 25 0 1.38275e-19 $X=12.025 $Y=0.74
r127 64 65 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=11.425 $Y=1.465
+ $X2=11.5 $Y2=1.465
r128 59 68 66.9444 $w=1.98e-07 $l=2.75e-07 $layer=POLY_cond $X=12.075 $Y=1.48
+ $X2=12.35 $Y2=1.48
r129 59 66 12.1717 $w=1.98e-07 $l=5e-08 $layer=POLY_cond $X=12.075 $Y=1.48
+ $X2=12.025 $Y2=1.48
r130 58 59 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=12.075
+ $Y=1.465 $X2=12.075 $Y2=1.465
r131 56 64 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=11.395 $Y=1.465
+ $X2=11.425 $Y2=1.465
r132 56 63 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.395 $Y=1.465
+ $X2=11.23 $Y2=1.465
r133 55 58 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=11.395 $Y=1.465
+ $X2=12.075 $Y2=1.465
r134 55 56 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=11.395
+ $Y=1.465 $X2=11.395 $Y2=1.465
r135 53 61 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=10.89 $Y=1.465
+ $X2=10.725 $Y2=1.465
r136 53 55 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=10.89 $Y=1.465
+ $X2=11.395 $Y2=1.465
r137 49 61 0.364692 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=10.725 $Y=1.3
+ $X2=10.725 $Y2=1.465
r138 49 51 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=10.725 $Y=1.3
+ $X2=10.725 $Y2=0.515
r139 47 61 6.46576 $w=2.5e-07 $l=2.0106e-07 $layer=LI1_cond $X=10.56 $Y=1.545
+ $X2=10.725 $Y2=1.465
r140 47 48 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=10.56 $Y=1.545
+ $X2=10.365 $Y2=1.545
r141 43 48 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.24 $Y=1.63
+ $X2=10.365 $Y2=1.545
r142 43 45 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=10.24 $Y=1.63
+ $X2=10.24 $Y2=2.19
r143 39 70 37.7323 $w=1.98e-07 $l=1.55e-07 $layer=POLY_cond $X=12.955 $Y=1.48
+ $X2=12.8 $Y2=1.48
r144 39 41 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=12.955 $Y=1.48
+ $X2=12.955 $Y2=0.74
r145 35 70 5.10115 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=12.8 $Y=1.63
+ $X2=12.8 $Y2=1.48
r146 35 37 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=12.8 $Y=1.63
+ $X2=12.8 $Y2=2.4
r147 31 70 66.9444 $w=1.98e-07 $l=2.75e-07 $layer=POLY_cond $X=12.525 $Y=1.48
+ $X2=12.8 $Y2=1.48
r148 31 68 42.601 $w=1.98e-07 $l=1.75e-07 $layer=POLY_cond $X=12.525 $Y=1.48
+ $X2=12.35 $Y2=1.48
r149 31 33 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=12.525 $Y=1.48
+ $X2=12.525 $Y2=0.74
r150 27 68 5.10115 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=12.35 $Y=1.63
+ $X2=12.35 $Y2=1.48
r151 27 29 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=12.35 $Y=1.63
+ $X2=12.35 $Y2=2.4
r152 23 66 9.34494 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=12.025 $Y=1.3
+ $X2=12.025 $Y2=1.48
r153 23 25 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=12.025 $Y=1.3
+ $X2=12.025 $Y2=0.74
r154 22 65 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=11.575 $Y=1.465
+ $X2=11.5 $Y2=1.465
r155 21 66 18.6067 $w=3.3e-07 $l=8.21584e-08 $layer=POLY_cond $X=11.95 $Y=1.465
+ $X2=12.025 $Y2=1.48
r156 21 22 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=11.95 $Y=1.465
+ $X2=11.575 $Y2=1.465
r157 17 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.5 $Y=1.3
+ $X2=11.5 $Y2=1.465
r158 17 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.5 $Y=1.3
+ $X2=11.5 $Y2=0.74
r159 13 64 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=11.425 $Y=1.63
+ $X2=11.425 $Y2=1.465
r160 13 15 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=11.425 $Y=1.63
+ $X2=11.425 $Y2=2.4
r161 12 63 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=11.02 $Y=1.555
+ $X2=11.23 $Y2=1.555
r162 7 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=10.93 $Y=1.63
+ $X2=11.02 $Y2=1.555
r163 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=10.93 $Y=1.63
+ $X2=10.93 $Y2=2.4
r164 2 45 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=10.065
+ $Y=2.045 $X2=10.2 $Y2=2.19
r165 1 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.585
+ $Y=0.37 $X2=10.725 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_4%VPWR 1 2 3 4 5 6 7 8 9 10 31 33 37 41 45 49
+ 53 57 61 65 67 69 74 75 77 78 80 81 82 84 89 94 102 120 124 133 136 139 142
+ 145 149
c170 149 0 2.33512e-20 $X=13.2 $Y=3.33
c171 61 0 1.07146e-19 $X=10.7 $Y=2.19
r172 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r173 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r174 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r175 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r176 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r177 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r178 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r179 128 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r180 128 146 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=11.76 $Y2=3.33
r181 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r182 125 145 13.7128 $w=1.7e-07 $l=3.53e-07 $layer=LI1_cond $X=12.24 $Y=3.33
+ $X2=11.887 $Y2=3.33
r183 125 127 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r184 124 148 4.57341 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=12.91 $Y=3.33
+ $X2=13.175 $Y2=3.33
r185 124 127 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=12.91 $Y=3.33
+ $X2=12.72 $Y2=3.33
r186 123 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r187 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r188 120 145 13.7128 $w=1.7e-07 $l=3.52e-07 $layer=LI1_cond $X=11.535 $Y=3.33
+ $X2=11.887 $Y2=3.33
r189 120 122 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.535 $Y=3.33
+ $X2=11.28 $Y2=3.33
r190 119 123 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r191 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r192 116 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r193 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r194 113 116 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r195 112 113 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r196 110 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r197 109 112 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=8.4 $Y2=3.33
r198 109 110 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r199 107 142 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=6.165 $Y=3.33
+ $X2=5.997 $Y2=3.33
r200 107 109 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.165 $Y=3.33
+ $X2=6.48 $Y2=3.33
r201 106 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r202 106 140 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r203 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r204 103 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.73 $Y=3.33
+ $X2=4.565 $Y2=3.33
r205 103 105 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.73 $Y=3.33
+ $X2=5.52 $Y2=3.33
r206 102 142 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=5.83 $Y=3.33
+ $X2=5.997 $Y2=3.33
r207 102 105 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.83 $Y=3.33
+ $X2=5.52 $Y2=3.33
r208 101 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r209 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r210 98 101 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r211 98 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r212 97 100 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r213 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r214 95 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=2.17 $Y2=3.33
r215 95 97 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=2.64 $Y2=3.33
r216 94 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.4 $Y=3.33
+ $X2=4.565 $Y2=3.33
r217 94 100 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.4 $Y=3.33
+ $X2=4.08 $Y2=3.33
r218 93 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r219 93 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r220 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r221 90 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.34 $Y=3.33
+ $X2=1.175 $Y2=3.33
r222 90 92 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.34 $Y=3.33
+ $X2=1.68 $Y2=3.33
r223 89 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=3.33
+ $X2=2.17 $Y2=3.33
r224 89 92 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.005 $Y=3.33
+ $X2=1.68 $Y2=3.33
r225 88 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r226 88 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r227 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r228 85 130 4.01803 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.36 $Y=3.33
+ $X2=0.18 $Y2=3.33
r229 85 87 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.36 $Y=3.33
+ $X2=0.72 $Y2=3.33
r230 84 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.01 $Y=3.33
+ $X2=1.175 $Y2=3.33
r231 84 87 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.01 $Y=3.33
+ $X2=0.72 $Y2=3.33
r232 82 113 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=8.4 $Y2=3.33
r233 82 110 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=6.48 $Y2=3.33
r234 80 118 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=10.535 $Y=3.33
+ $X2=10.32 $Y2=3.33
r235 80 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.535 $Y=3.33
+ $X2=10.7 $Y2=3.33
r236 79 122 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=10.865 $Y=3.33
+ $X2=11.28 $Y2=3.33
r237 79 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.865 $Y=3.33
+ $X2=10.7 $Y2=3.33
r238 77 115 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=9.65 $Y=3.33
+ $X2=9.36 $Y2=3.33
r239 77 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.65 $Y=3.33
+ $X2=9.775 $Y2=3.33
r240 76 118 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=9.9 $Y=3.33
+ $X2=10.32 $Y2=3.33
r241 76 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.9 $Y=3.33
+ $X2=9.775 $Y2=3.33
r242 74 112 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.58 $Y=3.33
+ $X2=8.4 $Y2=3.33
r243 74 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.58 $Y=3.33
+ $X2=8.745 $Y2=3.33
r244 73 115 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=8.91 $Y=3.33
+ $X2=9.36 $Y2=3.33
r245 73 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.91 $Y=3.33
+ $X2=8.745 $Y2=3.33
r246 69 72 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=13.075 $Y=2.115
+ $X2=13.075 $Y2=2.815
r247 67 148 3.19276 $w=3.3e-07 $l=1.36015e-07 $layer=LI1_cond $X=13.075 $Y=3.245
+ $X2=13.175 $Y2=3.33
r248 67 72 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.075 $Y=3.245
+ $X2=13.075 $Y2=2.815
r249 63 145 2.87722 $w=7.05e-07 $l=8.5e-08 $layer=LI1_cond $X=11.887 $Y=3.245
+ $X2=11.887 $Y2=3.33
r250 63 65 15.9477 $w=7.03e-07 $l=9.4e-07 $layer=LI1_cond $X=11.887 $Y=3.245
+ $X2=11.887 $Y2=2.305
r251 59 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.7 $Y=3.245
+ $X2=10.7 $Y2=3.33
r252 59 61 36.8433 $w=3.28e-07 $l=1.055e-06 $layer=LI1_cond $X=10.7 $Y=3.245
+ $X2=10.7 $Y2=2.19
r253 55 78 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.775 $Y=3.245
+ $X2=9.775 $Y2=3.33
r254 55 57 26.2757 $w=2.48e-07 $l=5.7e-07 $layer=LI1_cond $X=9.775 $Y=3.245
+ $X2=9.775 $Y2=2.675
r255 51 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.745 $Y=3.245
+ $X2=8.745 $Y2=3.33
r256 51 53 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=8.745 $Y=3.245
+ $X2=8.745 $Y2=2.675
r257 47 142 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=5.997 $Y=3.245
+ $X2=5.997 $Y2=3.33
r258 47 49 14.2765 $w=3.33e-07 $l=4.15e-07 $layer=LI1_cond $X=5.997 $Y=3.245
+ $X2=5.997 $Y2=2.83
r259 43 139 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=3.245
+ $X2=4.565 $Y2=3.33
r260 43 45 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=4.565 $Y=3.245
+ $X2=4.565 $Y2=2.825
r261 39 136 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=3.33
r262 39 41 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=2.815
r263 35 133 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.175 $Y=3.245
+ $X2=1.175 $Y2=3.33
r264 35 37 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.175 $Y=3.245
+ $X2=1.175 $Y2=2.815
r265 31 130 3.12513 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.235 $Y=3.245
+ $X2=0.18 $Y2=3.33
r266 31 33 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.235 $Y=3.245
+ $X2=0.235 $Y2=2.75
r267 10 72 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=12.89
+ $Y=1.84 $X2=13.075 $Y2=2.815
r268 10 69 400 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=1 $X=12.89
+ $Y=1.84 $X2=13.075 $Y2=2.115
r269 9 65 150 $w=1.7e-07 $l=8.04581e-07 $layer=licon1_PDIFF $count=4 $X=11.515
+ $Y=1.84 $X2=12.12 $Y2=2.305
r270 8 61 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=10.515
+ $Y=2.045 $X2=10.7 $Y2=2.19
r271 7 57 600 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_PDIFF $count=1 $X=9.56
+ $Y=2.465 $X2=9.735 $Y2=2.675
r272 6 53 600 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_PDIFF $count=1 $X=8.57
+ $Y=2.465 $X2=8.745 $Y2=2.675
r273 5 49 600 $w=1.7e-07 $l=2.41402e-07 $layer=licon1_PDIFF $count=1 $X=5.81
+ $Y=2.7 $X2=5.995 $Y2=2.83
r274 4 45 600 $w=1.7e-07 $l=6.08071e-07 $layer=licon1_PDIFF $count=1 $X=4.35
+ $Y=2.315 $X2=4.565 $Y2=2.825
r275 3 41 600 $w=1.7e-07 $l=9.04986e-07 $layer=licon1_PDIFF $count=1 $X=2.035
+ $Y=1.975 $X2=2.17 $Y2=2.815
r276 2 37 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.04
+ $Y=2.54 $X2=1.175 $Y2=2.815
r277 1 33 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.275 $Y2=2.75
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_4%A_37_78# 1 2 3 4 13 17 20 21 25 27 29 30 32
+ 34 38 40
c117 29 0 1.35567e-19 $X=3.625 $Y=1.305
r118 40 42 4.00386 $w=2.59e-07 $l=8.5e-08 $layer=LI1_cond $X=3.195 $Y=2.475
+ $X2=3.195 $Y2=2.56
r119 39 40 13.4247 $w=2.59e-07 $l=2.85e-07 $layer=LI1_cond $X=3.195 $Y=2.19
+ $X2=3.195 $Y2=2.475
r120 34 36 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.33 $Y=0.6
+ $X2=0.33 $Y2=0.745
r121 31 32 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=3.71 $Y=1.39
+ $X2=3.71 $Y2=2.105
r122 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.625 $Y=1.305
+ $X2=3.71 $Y2=1.39
r123 29 30 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.625 $Y=1.305
+ $X2=3.435 $Y2=1.305
r124 28 39 3.20129 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.36 $Y=2.19
+ $X2=3.195 $Y2=2.19
r125 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.625 $Y=2.19
+ $X2=3.71 $Y2=2.105
r126 27 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.625 $Y=2.19
+ $X2=3.36 $Y2=2.19
r127 23 30 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.31 $Y=1.22
+ $X2=3.435 $Y2=1.305
r128 23 25 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=3.31 $Y=1.22
+ $X2=3.31 $Y2=0.9
r129 22 38 2.36881 $w=1.7e-07 $l=3.46771e-07 $layer=LI1_cond $X=0.885 $Y=2.475
+ $X2=0.56 $Y2=2.52
r130 21 40 3.20129 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.03 $Y=2.475
+ $X2=3.195 $Y2=2.475
r131 21 22 139.941 $w=1.68e-07 $l=2.145e-06 $layer=LI1_cond $X=3.03 $Y=2.475
+ $X2=0.885 $Y2=2.475
r132 20 38 4.06715 $w=2.25e-07 $l=2.67208e-07 $layer=LI1_cond $X=0.77 $Y=2.39
+ $X2=0.56 $Y2=2.52
r133 19 20 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=0.77 $Y=0.83
+ $X2=0.77 $Y2=2.39
r134 15 38 4.06715 $w=2.25e-07 $l=1.77482e-07 $layer=LI1_cond $X=0.7 $Y=2.605
+ $X2=0.56 $Y2=2.52
r135 15 17 8.64332 $w=2.78e-07 $l=2.1e-07 $layer=LI1_cond $X=0.7 $Y=2.605
+ $X2=0.7 $Y2=2.815
r136 14 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.495 $Y=0.745
+ $X2=0.33 $Y2=0.745
r137 13 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.685 $Y=0.745
+ $X2=0.77 $Y2=0.83
r138 13 14 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.685 $Y=0.745
+ $X2=0.495 $Y2=0.745
r139 4 42 600 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_PDIFF $count=1 $X=3.055
+ $Y=2.315 $X2=3.195 $Y2=2.56
r140 3 17 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=2.54 $X2=0.725 $Y2=2.815
r141 2 25 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=3.145
+ $Y=0.69 $X2=3.27 $Y2=0.9
r142 1 34 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.39 $X2=0.33 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_4%Q 1 2 3 4 15 19 20 21 23 25 29 35 38 41 42
c71 42 0 1.38275e-19 $X=13.2 $Y=1.665
r72 44 45 2.94971 $w=5.17e-07 $l=1.25e-07 $layer=LI1_cond $X=12.575 $Y=1.62
+ $X2=12.7 $Y2=1.62
r73 42 45 11.7988 $w=5.17e-07 $l=5e-07 $layer=LI1_cond $X=13.2 $Y=1.62 $X2=12.7
+ $Y2=1.62
r74 38 45 5.00057 $w=2.5e-07 $l=3.5e-07 $layer=LI1_cond $X=12.7 $Y=1.27 $X2=12.7
+ $Y2=1.62
r75 37 41 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=12.7 $Y=1.13
+ $X2=12.7 $Y2=1.005
r76 37 38 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=12.7 $Y=1.13
+ $X2=12.7 $Y2=1.27
r77 33 41 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=12.7 $Y=0.88
+ $X2=12.7 $Y2=1.005
r78 33 35 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=12.7 $Y=0.88
+ $X2=12.7 $Y2=0.515
r79 29 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=12.575 $Y=1.985
+ $X2=12.575 $Y2=2.815
r80 27 44 3.36414 $w=3.3e-07 $l=3.5e-07 $layer=LI1_cond $X=12.575 $Y=1.97
+ $X2=12.575 $Y2=1.62
r81 27 29 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=12.575 $Y=1.97
+ $X2=12.575 $Y2=1.985
r82 26 40 3.87155 $w=2.5e-07 $l=1.58e-07 $layer=LI1_cond $X=11.91 $Y=1.005
+ $X2=11.752 $Y2=1.005
r83 25 41 1.34256 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=12.575 $Y=1.005
+ $X2=12.7 $Y2=1.005
r84 25 26 30.655 $w=2.48e-07 $l=6.65e-07 $layer=LI1_cond $X=12.575 $Y=1.005
+ $X2=11.91 $Y2=1.005
r85 21 40 3.06294 $w=3.15e-07 $l=1.25e-07 $layer=LI1_cond $X=11.752 $Y=0.88
+ $X2=11.752 $Y2=1.005
r86 21 23 12.8049 $w=3.13e-07 $l=3.5e-07 $layer=LI1_cond $X=11.752 $Y=0.88
+ $X2=11.752 $Y2=0.53
r87 19 44 9.81494 $w=5.17e-07 $l=3.37565e-07 $layer=LI1_cond $X=12.41 $Y=1.885
+ $X2=12.575 $Y2=1.62
r88 19 20 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=12.41 $Y=1.885
+ $X2=11.365 $Y2=1.885
r89 15 17 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=11.2 $Y=1.985
+ $X2=11.2 $Y2=2.815
r90 13 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.2 $Y=1.97
+ $X2=11.365 $Y2=1.885
r91 13 15 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=11.2 $Y=1.97
+ $X2=11.2 $Y2=1.985
r92 4 31 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=12.44
+ $Y=1.84 $X2=12.575 $Y2=2.815
r93 4 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=12.44
+ $Y=1.84 $X2=12.575 $Y2=1.985
r94 3 17 400 $w=1.7e-07 $l=1.06119e-06 $layer=licon1_PDIFF $count=1 $X=11.02
+ $Y=1.84 $X2=11.2 $Y2=2.815
r95 3 15 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=11.02
+ $Y=1.84 $X2=11.2 $Y2=1.985
r96 2 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.6
+ $Y=0.37 $X2=12.74 $Y2=0.515
r97 1 40 182 $w=1.7e-07 $l=6.81249e-07 $layer=licon1_NDIFF $count=1 $X=11.575
+ $Y=0.37 $X2=11.76 $Y2=0.965
r98 1 23 182 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=1 $X=11.575
+ $Y=0.37 $X2=11.76 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTP_4%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 49 51
+ 54 55 57 58 59 65 69 77 89 93 98 104 108 114 117 120 124
c141 124 0 6.43803e-21 $X=13.2 $Y=0
r142 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r143 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r144 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r145 114 115 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r146 108 111 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=5.06 $Y=0
+ $X2=5.06 $Y2=0.285
r147 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r148 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r149 102 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r150 102 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r151 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r152 99 120 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=12.405 $Y=0
+ $X2=12.242 $Y2=0
r153 99 101 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.405 $Y=0
+ $X2=12.72 $Y2=0
r154 98 123 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=13.005 $Y=0
+ $X2=13.222 $Y2=0
r155 98 101 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=13.005 $Y=0
+ $X2=12.72 $Y2=0
r156 97 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r157 97 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r158 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r159 94 117 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.41 $Y=0
+ $X2=11.265 $Y2=0
r160 94 96 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=11.41 $Y=0
+ $X2=11.76 $Y2=0
r161 93 120 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=12.08 $Y=0
+ $X2=12.242 $Y2=0
r162 93 96 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=12.08 $Y=0 $X2=11.76
+ $Y2=0
r163 92 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r164 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r165 89 117 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.12 $Y=0
+ $X2=11.265 $Y2=0
r166 89 91 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=11.12 $Y=0 $X2=10.8
+ $Y2=0
r167 88 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=10.8
+ $Y2=0
r168 88 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=8.88 $Y2=0
r169 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r170 85 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.955 $Y=0
+ $X2=8.79 $Y2=0
r171 85 87 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=8.955 $Y=0 $X2=9.84
+ $Y2=0
r172 84 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r173 83 84 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r174 81 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=5.04 $Y2=0
r175 80 83 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=8.4
+ $Y2=0
r176 80 81 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r177 78 108 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.225 $Y=0
+ $X2=5.06 $Y2=0
r178 78 80 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.225 $Y=0 $X2=5.52
+ $Y2=0
r179 77 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.625 $Y=0
+ $X2=8.79 $Y2=0
r180 77 83 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=8.625 $Y=0 $X2=8.4
+ $Y2=0
r181 76 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.04 $Y2=0
r182 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r183 73 76 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.56 $Y2=0
r184 73 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=2.16 $Y2=0
r185 72 75 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r186 72 73 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r187 70 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=0
+ $X2=2.21 $Y2=0
r188 70 72 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.375 $Y=0
+ $X2=2.64 $Y2=0
r189 69 108 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.895 $Y=0
+ $X2=5.06 $Y2=0
r190 69 75 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.895 $Y=0
+ $X2=4.56 $Y2=0
r191 68 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r192 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r193 65 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.045 $Y=0
+ $X2=2.21 $Y2=0
r194 65 67 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.045 $Y=0
+ $X2=1.68 $Y2=0
r195 63 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r196 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r197 59 84 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=6.72 $Y=0 $X2=8.4
+ $Y2=0
r198 59 81 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=6.72 $Y=0 $X2=5.52
+ $Y2=0
r199 57 87 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=9.84 $Y2=0
r200 57 58 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=10.252 $Y2=0
r201 56 91 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=10.39 $Y=0 $X2=10.8
+ $Y2=0
r202 56 58 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=10.39 $Y=0
+ $X2=10.252 $Y2=0
r203 54 62 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.72
+ $Y2=0
r204 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.065 $Y=0 $X2=1.15
+ $Y2=0
r205 53 67 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.235 $Y=0
+ $X2=1.68 $Y2=0
r206 53 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.15
+ $Y2=0
r207 49 123 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=13.17 $Y=0.085
+ $X2=13.222 $Y2=0
r208 49 51 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.17 $Y=0.085
+ $X2=13.17 $Y2=0.515
r209 45 120 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=12.242 $Y=0.085
+ $X2=12.242 $Y2=0
r210 45 47 15.7796 $w=3.23e-07 $l=4.45e-07 $layer=LI1_cond $X=12.242 $Y=0.085
+ $X2=12.242 $Y2=0.53
r211 41 117 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=11.265 $Y=0.085
+ $X2=11.265 $Y2=0
r212 41 43 17.684 $w=2.88e-07 $l=4.45e-07 $layer=LI1_cond $X=11.265 $Y=0.085
+ $X2=11.265 $Y2=0.53
r213 37 58 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=10.252 $Y=0.085
+ $X2=10.252 $Y2=0
r214 37 39 18.02 $w=2.73e-07 $l=4.3e-07 $layer=LI1_cond $X=10.252 $Y=0.085
+ $X2=10.252 $Y2=0.515
r215 33 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.79 $Y=0.085
+ $X2=8.79 $Y2=0
r216 33 35 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=8.79 $Y=0.085
+ $X2=8.79 $Y2=0.615
r217 29 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.21 $Y=0.085
+ $X2=2.21 $Y2=0
r218 29 31 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=2.21 $Y=0.085
+ $X2=2.21 $Y2=0.715
r219 25 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0
r220 25 27 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0.6
r221 8 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.03
+ $Y=0.37 $X2=13.17 $Y2=0.515
r222 7 47 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=12.1
+ $Y=0.37 $X2=12.24 $Y2=0.53
r223 6 43 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=11.14
+ $Y=0.37 $X2=11.285 $Y2=0.53
r224 5 39 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=10.08
+ $Y=0.37 $X2=10.225 $Y2=0.515
r225 4 35 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=8.625
+ $Y=0.405 $X2=8.79 $Y2=0.615
r226 3 111 182 $w=1.7e-07 $l=5.03115e-07 $layer=licon1_NDIFF $count=1 $X=4.84
+ $Y=0.69 $X2=5.06 $Y2=0.285
r227 2 31 182 $w=1.7e-07 $l=2.37539e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.595 $X2=2.21 $Y2=0.715
r228 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.01
+ $Y=0.39 $X2=1.15 $Y2=0.6
.ends


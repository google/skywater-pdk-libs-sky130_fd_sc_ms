* File: sky130_fd_sc_ms__dlrtp_1.spice
* Created: Fri Aug 28 17:28:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dlrtp_1.pex.spice"
.subckt sky130_fd_sc_ms__dlrtp_1  VNB VPB D GATE RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1017 N_VGND_M1017_d N_D_M1017_g N_A_27_424#_M1017_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.125093 AS=0.15675 PD=1.00194 PS=1.67 NRD=34.356 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1007 N_A_219_424#_M1007_d N_GATE_M1007_g N_VGND_M1017_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.168307 PD=2.05 PS=1.34806 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_A_219_424#_M1012_g N_A_363_74#_M1012_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.136954 AS=0.32225 PD=1.17971 PS=2.64 NRD=4.86 NRS=61.692 M=1
+ R=4.93333 SA=75000.3 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1018 A_565_74# N_A_27_424#_M1018_g N_VGND_M1012_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.118446 PD=0.88 PS=1.02029 NRD=12.18 NRS=9.372 M=1 R=4.26667
+ SA=75000.8 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1019 N_A_643_74#_M1019_d N_A_363_74#_M1019_g A_565_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.175517 AS=0.0768 PD=1.35245 PS=0.88 NRD=11.244 NRS=12.18 M=1
+ R=4.26667 SA=75001.2 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1010 A_769_74# N_A_219_424#_M1010_g N_A_643_74#_M1019_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.115183 PD=0.66 PS=0.887547 NRD=18.564 NRS=41.424 M=1
+ R=2.8 SA=75001.8 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_817_48#_M1011_g A_769_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 A_1045_74# N_A_643_74#_M1015_g N_A_817_48#_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1009 N_VGND_M1009_d N_RESET_B_M1009_g A_1045_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1332 AS=0.0888 PD=1.1 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75000.6
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1014 N_Q_M1014_d N_A_817_48#_M1014_g N_VGND_M1009_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1332 PD=2.05 PS=1.1 NRD=0 NRS=12.972 M=1 R=4.93333 SA=75001.1
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1008 N_VPWR_M1008_d N_D_M1008_g N_A_27_424#_M1008_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1344 AS=0.2352 PD=1.16 PS=2.24 NRD=10.5395 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.9 A=0.1512 P=2.04 MULT=1
MM1006 N_A_219_424#_M1006_d N_GATE_M1006_g N_VPWR_M1008_d VPB PSHORT L=0.18
+ W=0.84 AD=0.42675 AS=0.1344 PD=2.84 PS=1.16 NRD=29.3136 NRS=0 M=1 R=4.66667
+ SA=90000.7 SB=90000.4 A=0.1512 P=2.04 MULT=1
MM1001 N_VPWR_M1001_d N_A_219_424#_M1001_g N_A_363_74#_M1001_s VPB PSHORT L=0.18
+ W=0.84 AD=0.17713 AS=0.2352 PD=1.27826 PS=2.24 NRD=24.625 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90002.1 A=0.1512 P=2.04 MULT=1
MM1016 A_571_392# N_A_27_424#_M1016_g N_VPWR_M1001_d VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.21087 PD=1.24 PS=1.52174 NRD=12.7853 NRS=3.9203 M=1 R=5.55556
+ SA=90000.7 SB=90001.9 A=0.18 P=2.36 MULT=1
MM1000 N_A_643_74#_M1000_d N_A_219_424#_M1000_g A_571_392# VPB PSHORT L=0.18 W=1
+ AD=0.219366 AS=0.12 PD=1.90845 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556
+ SA=90001.1 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1005 A_762_508# N_A_363_74#_M1005_g N_A_643_74#_M1000_d VPB PSHORT L=0.18
+ W=0.42 AD=0.09975 AS=0.0921338 PD=0.895 PS=0.801549 NRD=85.5965 NRS=39.8531
+ M=1 R=2.33333 SA=90001.5 SB=90002.7 A=0.0756 P=1.2 MULT=1
MM1013 N_VPWR_M1013_d N_A_817_48#_M1013_g A_762_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.114938 AS=0.09975 PD=0.934648 PS=0.895 NRD=70.3487 NRS=85.5965 M=1
+ R=2.33333 SA=90002.2 SB=90002 A=0.0756 P=1.2 MULT=1
MM1003 N_A_817_48#_M1003_d N_A_643_74#_M1003_g N_VPWR_M1013_d VPB PSHORT L=0.18
+ W=1 AD=0.16 AS=0.273662 PD=1.32 PS=2.22535 NRD=8.8453 NRS=29.55 M=1 R=5.55556
+ SA=90001.3 SB=90001.3 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_RESET_B_M1002_g N_A_817_48#_M1003_d VPB PSHORT L=0.18
+ W=1 AD=0.20283 AS=0.16 PD=1.43396 PS=1.32 NRD=8.8453 NRS=0 M=1 R=5.55556
+ SA=90001.8 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1004 N_Q_M1004_d N_A_817_48#_M1004_g N_VPWR_M1002_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.22717 PD=2.8 PS=1.60604 NRD=0 NRS=13.1793 M=1 R=6.22222
+ SA=90002.2 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX20_noxref VNB VPB NWDIODE A=12.9966 P=18.16
c_858 A_571_392# 0 1.45332e-19 $X=2.855 $Y=1.96
c_959 A_565_74# 0 5.47968e-20 $X=2.825 $Y=0.37
*
.include "sky130_fd_sc_ms__dlrtp_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__a2bb2oi_4.spice
* Created: Fri Aug 28 17:05:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a2bb2oi_4.pex.spice"
.subckt sky130_fd_sc_ms__a2bb2oi_4  VNB VPB A2_N A1_N B2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* B2	B2
* A1_N	A1_N
* A2_N	A2_N
* VPB	VPB
* VNB	VNB
MM1027 N_A_117_392#_M1027_d N_A2_N_M1027_g N_VGND_M1027_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.4 A=0.111 P=1.78 MULT=1
MM1006 N_VGND_M1006_d N_A1_N_M1006_g N_A_117_392#_M1027_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1184 AS=0.1036 PD=1.06 PS=1.02 NRD=3.24 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75002 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1006_d N_A_117_392#_M1003_g N_Y_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1184 AS=0.1036 PD=1.06 PS=1.02 NRD=3.24 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A_117_392#_M1004_g N_Y_M1003_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1004_d N_A_117_392#_M1014_g N_Y_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1028 N_VGND_M1028_d N_A_117_392#_M1028_g N_Y_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.4
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_Y_M1001_d N_B2_M1001_g N_A_914_74#_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1961 PD=1.02 PS=2.01 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75003.2 A=0.111 P=1.78 MULT=1
MM1009 N_Y_M1001_d N_B2_M1009_g N_A_914_74#_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75002.8 A=0.111 P=1.78 MULT=1
MM1012 N_Y_M1012_d N_B2_M1012_g N_A_914_74#_M1009_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1013 N_Y_M1012_d N_B2_M1013_g N_A_914_74#_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1000 N_A_914_74#_M1013_s N_B1_M1000_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.9
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1011 N_A_914_74#_M1011_d N_B1_M1011_g N_VGND_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.3
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1025 N_A_914_74#_M1011_d N_B1_M1025_g N_VGND_M1025_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1029 N_A_914_74#_M1029_d N_B1_M1029_g N_VGND_M1025_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.1036 PD=2.01 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1017 N_A_117_392#_M1017_d N_A2_N_M1017_g N_A_29_392#_M1017_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.5 A=0.18 P=2.36 MULT=1
MM1018 N_A_117_392#_M1017_d N_A2_N_M1018_g N_A_29_392#_M1018_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.6
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1020 N_VPWR_M1020_d N_A1_N_M1020_g N_A_29_392#_M1018_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.135 PD=1.27 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.1
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1022 N_VPWR_M1020_d N_A1_N_M1022_g N_A_29_392#_M1022_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.26 PD=1.27 PS=2.52 NRD=0 NRS=0 M=1 R=5.55556 SA=90001.5
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1015 N_Y_M1015_d N_A_117_392#_M1015_g N_A_539_368#_M1015_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90005.1 A=0.2016 P=2.6 MULT=1
MM1021 N_Y_M1015_d N_A_117_392#_M1021_g N_A_539_368#_M1021_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90004.7 A=0.2016 P=2.6 MULT=1
MM1023 N_Y_M1023_d N_A_117_392#_M1023_g N_A_539_368#_M1021_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.1 SB=90004.2 A=0.2016 P=2.6 MULT=1
MM1024 N_Y_M1023_d N_A_117_392#_M1024_g N_A_539_368#_M1024_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.5 SB=90003.8 A=0.2016 P=2.6 MULT=1
MM1002 N_A_539_368#_M1024_s N_B2_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90003.3 A=0.2016 P=2.6 MULT=1
MM1005 N_A_539_368#_M1005_d N_B2_M1005_g N_VPWR_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.4
+ SB=90002.9 A=0.2016 P=2.6 MULT=1
MM1007 N_A_539_368#_M1005_d N_B2_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.9
+ SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1026 N_A_539_368#_M1026_d N_B2_M1026_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.3
+ SB=90002 A=0.2016 P=2.6 MULT=1
MM1008 N_VPWR_M1008_d N_B1_M1008_g N_A_539_368#_M1026_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.8
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1010 N_VPWR_M1008_d N_B1_M1010_g N_A_539_368#_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.2
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1016 N_VPWR_M1016_d N_B1_M1016_g N_A_539_368#_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.7
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1019 N_VPWR_M1016_d N_B1_M1019_g N_A_539_368#_M1019_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2912 PD=1.39 PS=2.76 NRD=0 NRS=0 M=1 R=6.22222 SA=90005.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX30_noxref VNB VPB NWDIODE A=16.7772 P=21.76
*
.include "sky130_fd_sc_ms__a2bb2oi_4.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__nor4bb_1.pex.spice
* Created: Wed Sep  2 12:17:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NOR4BB_1%C_N 3 5 7 8 13
r26 13 14 33.7665 $w=3.64e-07 $l=2.55e-07 $layer=POLY_cond $X=0.505 $Y=1.415
+ $X2=0.76 $Y2=1.415
r27 11 13 31.1181 $w=3.64e-07 $l=2.35e-07 $layer=POLY_cond $X=0.27 $Y=1.415
+ $X2=0.505 $Y2=1.415
r28 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.385 $X2=0.27 $Y2=1.385
r29 8 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.27 $Y=1.295 $X2=0.27
+ $Y2=1.385
r30 5 14 23.572 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=0.76 $Y=1.22 $X2=0.76
+ $Y2=1.415
r31 5 7 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.76 $Y=1.22 $X2=0.76
+ $Y2=0.835
r32 1 13 19.2285 $w=1.8e-07 $l=1.95e-07 $layer=POLY_cond $X=0.505 $Y=1.61
+ $X2=0.505 $Y2=1.415
r33 1 3 252.661 $w=1.8e-07 $l=6.5e-07 $layer=POLY_cond $X=0.505 $Y=1.61
+ $X2=0.505 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4BB_1%A 3 7 9 10 15 18
r42 17 18 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=1.395 $Y=1.515
+ $X2=1.49 $Y2=1.515
r43 14 17 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=1.24 $Y=1.515
+ $X2=1.395 $Y2=1.515
r44 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.24
+ $Y=1.515 $X2=1.24 $Y2=1.515
r45 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.24 $Y=1.665
+ $X2=1.24 $Y2=2.035
r46 9 15 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.24 $Y=1.665
+ $X2=1.24 $Y2=1.515
r47 5 18 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.49 $Y=1.68
+ $X2=1.49 $Y2=1.515
r48 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.49 $Y=1.68 $X2=1.49
+ $Y2=2.4
r49 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.395 $Y=1.35
+ $X2=1.395 $Y2=1.515
r50 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.395 $Y=1.35
+ $X2=1.395 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4BB_1%B 3 7 9 15 16
c36 7 0 3.40843e-20 $X=1.91 $Y=2.4
r37 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.08
+ $Y=1.515 $X2=2.08 $Y2=1.515
r38 13 15 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=1.91 $Y=1.515
+ $X2=2.08 $Y2=1.515
r39 11 13 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.895 $Y=1.515
+ $X2=1.91 $Y2=1.515
r40 9 16 4.80185 $w=3.58e-07 $l=1.5e-07 $layer=LI1_cond $X=2.095 $Y=1.665
+ $X2=2.095 $Y2=1.515
r41 5 13 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.91 $Y=1.68
+ $X2=1.91 $Y2=1.515
r42 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.91 $Y=1.68 $X2=1.91
+ $Y2=2.4
r43 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=1.35
+ $X2=1.895 $Y2=1.515
r44 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.895 $Y=1.35
+ $X2=1.895 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4BB_1%A_27_112# 1 2 9 13 15 20 24 25 27 28 30 32
+ 33
c102 24 0 3.40843e-20 $X=2.65 $Y=1.515
r103 32 34 11.9608 $w=6.58e-07 $l=6.6e-07 $layer=LI1_cond $X=0.445 $Y=1.985
+ $X2=0.445 $Y2=2.645
r104 32 33 10.5469 $w=6.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=1.985
+ $X2=0.445 $Y2=1.82
r105 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.71 $Y=1.89
+ $X2=3.71 $Y2=2.56
r106 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.625 $Y=1.805
+ $X2=3.71 $Y2=1.89
r107 27 28 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=3.625 $Y=1.805
+ $X2=2.815 $Y2=1.805
r108 25 38 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.65 $Y=1.515
+ $X2=2.65 $Y2=1.68
r109 25 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.65 $Y=1.515
+ $X2=2.65 $Y2=1.35
r110 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.65
+ $Y=1.515 $X2=2.65 $Y2=1.515
r111 22 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.65 $Y=1.72
+ $X2=2.815 $Y2=1.805
r112 22 24 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=2.65 $Y=1.72
+ $X2=2.65 $Y2=1.515
r113 21 34 8.93547 $w=1.7e-07 $l=3.3e-07 $layer=LI1_cond $X=0.775 $Y=2.645
+ $X2=0.445 $Y2=2.645
r114 20 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.625 $Y=2.645
+ $X2=3.71 $Y2=2.56
r115 20 21 185.936 $w=1.68e-07 $l=2.85e-06 $layer=LI1_cond $X=3.625 $Y=2.645
+ $X2=0.775 $Y2=2.645
r116 18 33 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=0.69 $Y=1.01
+ $X2=0.69 $Y2=1.82
r117 15 18 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.605 $Y=0.845
+ $X2=0.69 $Y2=1.01
r118 15 17 2.21818 $w=3.3e-07 $l=6e-08 $layer=LI1_cond $X=0.605 $Y=0.845
+ $X2=0.545 $Y2=0.845
r119 13 37 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.74 $Y=0.74
+ $X2=2.74 $Y2=1.35
r120 9 38 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.575 $Y=2.4
+ $X2=2.575 $Y2=1.68
r121 2 32 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
r122 1 17 182 $w=1.7e-07 $l=5.33807e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.56 $X2=0.545 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4BB_1%A_611_244# 1 2 10 11 13 14 15 17 20 24 28
+ 33 36 37 38 43
c75 37 0 1.67721e-19 $X=4.52 $Y=1.175
c76 36 0 1.14509e-19 $X=3.74 $Y=1.32
c77 17 0 1.84713e-19 $X=3.665 $Y=3.035
r78 39 41 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=3.145 $Y=1.385
+ $X2=3.24 $Y2=1.385
r79 34 43 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.575 $Y=1.385
+ $X2=3.665 $Y2=1.385
r80 34 41 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=3.575 $Y=1.385
+ $X2=3.24 $Y2=1.385
r81 33 36 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.575 $Y=1.32
+ $X2=3.74 $Y2=1.32
r82 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.575
+ $Y=1.385 $X2=3.575 $Y2=1.385
r83 30 37 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.6 $Y=1.26
+ $X2=4.52 $Y2=1.175
r84 30 38 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.6 $Y=1.26 $X2=4.6
+ $Y2=2.1
r85 28 38 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.52 $Y=2.265
+ $X2=4.52 $Y2=2.1
r86 22 37 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.52 $Y=1.09 $X2=4.52
+ $Y2=1.175
r87 22 24 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=4.52 $Y=1.09
+ $X2=4.52 $Y2=0.835
r88 20 37 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.355 $Y=1.175
+ $X2=4.52 $Y2=1.175
r89 20 36 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.355 $Y=1.175
+ $X2=3.74 $Y2=1.175
r90 16 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.665 $Y=1.55
+ $X2=3.665 $Y2=1.385
r91 16 17 761.457 $w=1.5e-07 $l=1.485e-06 $layer=POLY_cond $X=3.665 $Y=1.55
+ $X2=3.665 $Y2=3.035
r92 14 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.59 $Y=3.11
+ $X2=3.665 $Y2=3.035
r93 14 15 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=3.59 $Y=3.11
+ $X2=3.235 $Y2=3.11
r94 11 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.24 $Y=1.22
+ $X2=3.24 $Y2=1.385
r95 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.24 $Y=1.22 $X2=3.24
+ $Y2=0.74
r96 8 15 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.145 $Y=3.035
+ $X2=3.235 $Y2=3.11
r97 8 10 246.831 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=3.145 $Y=3.035
+ $X2=3.145 $Y2=2.4
r98 7 39 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.145 $Y=1.55
+ $X2=3.145 $Y2=1.385
r99 7 10 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.145 $Y=1.55
+ $X2=3.145 $Y2=2.4
r100 2 28 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=4.385
+ $Y=2.12 $X2=4.52 $Y2=2.265
r101 1 24 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=4.38
+ $Y=0.56 $X2=4.52 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4BB_1%D_N 1 3 7 9 13
c33 13 0 1.84713e-19 $X=4.18 $Y=1.615
c34 1 0 2.8223e-19 $X=4.295 $Y=1.87
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.18
+ $Y=1.615 $X2=4.18 $Y2=1.615
r36 9 13 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=4.08 $Y=1.615 $X2=4.18
+ $Y2=1.615
r37 5 12 38.571 $w=3.25e-07 $l=2.11069e-07 $layer=POLY_cond $X=4.305 $Y=1.45
+ $X2=4.2 $Y2=1.615
r38 5 7 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=4.305 $Y=1.45
+ $X2=4.305 $Y2=0.835
r39 1 12 47.3393 $w=3.25e-07 $l=2.98747e-07 $layer=POLY_cond $X=4.295 $Y=1.87
+ $X2=4.2 $Y2=1.615
r40 1 3 260.435 $w=1.8e-07 $l=6.7e-07 $layer=POLY_cond $X=4.295 $Y=1.87
+ $X2=4.295 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4BB_1%VPWR 1 2 11 13 15 25 26 29 37 39
r40 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r41 35 37 9.14549 $w=5.13e-07 $l=1.45e-07 $layer=LI1_cond $X=1.2 $Y=3.157
+ $X2=1.345 $Y2=3.157
r42 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r43 33 35 0.464496 $w=5.13e-07 $l=2e-08 $layer=LI1_cond $X=1.18 $Y=3.157 $X2=1.2
+ $Y2=3.157
r44 30 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r45 29 33 10.6834 $w=5.13e-07 $l=4.6e-07 $layer=LI1_cond $X=0.72 $Y=3.157
+ $X2=1.18 $Y2=3.157
r46 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 26 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r48 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r49 23 39 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=4.185 $Y=3.33
+ $X2=4.075 $Y2=3.33
r50 23 25 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.185 $Y=3.33
+ $X2=4.56 $Y2=3.33
r51 22 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r52 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r53 19 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r54 18 21 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r55 18 37 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=1.345 $Y2=3.33
r56 18 19 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 15 39 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.965 $Y=3.33
+ $X2=4.075 $Y2=3.33
r58 15 21 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.965 $Y=3.33
+ $X2=3.6 $Y2=3.33
r59 13 22 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=3.6
+ $Y2=3.33
r60 13 19 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=1.68 $Y2=3.33
r61 9 39 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.075 $Y=3.245
+ $X2=4.075 $Y2=3.33
r62 9 11 51.3361 $w=2.18e-07 $l=9.8e-07 $layer=LI1_cond $X=4.075 $Y=3.245
+ $X2=4.075 $Y2=2.265
r63 2 11 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=3.945
+ $Y=2.12 $X2=4.07 $Y2=2.265
r64 1 33 300 $w=1.7e-07 $l=1.40743e-06 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=1.18 $Y2=2.985
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4BB_1%Y 1 2 3 12 15 16 18 20 23 25 28
r61 25 28 1.22927 $w=3.73e-07 $l=4e-08 $layer=LI1_cond $X=3.047 $Y=0.555
+ $X2=3.047 $Y2=0.515
r62 24 25 9.98784 $w=3.73e-07 $l=3.25e-07 $layer=LI1_cond $X=3.047 $Y=0.88
+ $X2=3.047 $Y2=0.555
r63 21 23 2.76166 $w=1.7e-07 $l=1.83916e-07 $layer=LI1_cond $X=1.775 $Y=0.965
+ $X2=1.61 $Y2=1.005
r64 20 24 8.1532 $w=1.7e-07 $l=2.2553e-07 $layer=LI1_cond $X=2.86 $Y=0.965
+ $X2=3.047 $Y2=0.88
r65 20 21 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=2.86 $Y=0.965
+ $X2=1.775 $Y2=0.965
r66 16 18 56.7491 $w=3.28e-07 $l=1.625e-06 $layer=LI1_cond $X=1.745 $Y=2.225
+ $X2=3.37 $Y2=2.225
r67 15 16 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.66 $Y=2.06
+ $X2=1.745 $Y2=2.225
r68 14 23 3.70735 $w=2.5e-07 $l=1.47902e-07 $layer=LI1_cond $X=1.66 $Y=1.13
+ $X2=1.61 $Y2=1.005
r69 14 15 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=1.66 $Y=1.13
+ $X2=1.66 $Y2=2.06
r70 10 23 3.70735 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.61 $Y=0.88
+ $X2=1.61 $Y2=1.005
r71 10 12 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.61 $Y=0.88
+ $X2=1.61 $Y2=0.515
r72 3 18 600 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=1 $X=3.235
+ $Y=1.84 $X2=3.37 $Y2=2.225
r73 2 28 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=2.815
+ $Y=0.37 $X2=3.025 $Y2=0.515
r74 1 23 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.47
+ $Y=0.37 $X2=1.61 $Y2=0.965
r75 1 12 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.47
+ $Y=0.37 $X2=1.61 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__NOR4BB_1%VGND 1 2 3 12 18 21 22 23 33 40 41 46 49 51
r56 52 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r57 51 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r58 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r59 48 49 11.2171 $w=7.63e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=0.297
+ $X2=2.69 $Y2=0.297
r60 44 48 5.70678 $w=7.63e-07 $l=3.65e-07 $layer=LI1_cond $X=2.16 $Y=0.297
+ $X2=2.525 $Y2=0.297
r61 44 46 11.9988 $w=7.63e-07 $l=2.15e-07 $layer=LI1_cond $X=2.16 $Y=0.297
+ $X2=1.945 $Y2=0.297
r62 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r63 41 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r64 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r65 38 51 14.3545 $w=1.7e-07 $l=3.85e-07 $layer=LI1_cond $X=4.175 $Y=0 $X2=3.79
+ $Y2=0
r66 38 40 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.175 $Y=0 $X2=4.56
+ $Y2=0
r67 37 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r68 36 49 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=2.69
+ $Y2=0
r69 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r70 33 51 14.3545 $w=1.7e-07 $l=3.85e-07 $layer=LI1_cond $X=3.405 $Y=0 $X2=3.79
+ $Y2=0
r71 33 36 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.405 $Y=0 $X2=3.12
+ $Y2=0
r72 32 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r73 31 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=1.945
+ $Y2=0
r74 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r75 27 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r76 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r77 23 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r78 23 45 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r79 21 26 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.72
+ $Y2=0
r80 21 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.11
+ $Y2=0
r81 20 31 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.275 $Y=0 $X2=1.68
+ $Y2=0
r82 20 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.275 $Y=0 $X2=1.11
+ $Y2=0
r83 16 51 3.05715 $w=7.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.79 $Y=0.085
+ $X2=3.79 $Y2=0
r84 16 18 6.36873 $w=7.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.79 $Y=0.085
+ $X2=3.79 $Y2=0.495
r85 12 14 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.11 $Y=0.515
+ $X2=1.11 $Y2=0.965
r86 10 22 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.11 $Y=0.085
+ $X2=1.11 $Y2=0
r87 10 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.11 $Y=0.085
+ $X2=1.11 $Y2=0.515
r88 3 18 45.5 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_NDIFF $count=4 $X=3.315
+ $Y=0.37 $X2=4.01 $Y2=0.495
r89 2 48 91 $w=1.7e-07 $l=6.23298e-07 $layer=licon1_NDIFF $count=2 $X=1.97
+ $Y=0.37 $X2=2.525 $Y2=0.515
r90 1 14 182 $w=1.7e-07 $l=5.24786e-07 $layer=licon1_NDIFF $count=1 $X=0.835
+ $Y=0.56 $X2=1.11 $Y2=0.965
r91 1 12 182 $w=1.7e-07 $l=2.96648e-07 $layer=licon1_NDIFF $count=1 $X=0.835
+ $Y=0.56 $X2=1.11 $Y2=0.515
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__o211ai_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__o211ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 0.435000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.550000 1.165000 1.630000 ;
        RECT 0.605000 1.630000 0.835000 2.890000 ;
        RECT 0.665000 1.300000 1.165000 1.550000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.405000 1.300000 1.795000 1.630000 ;
        RECT 1.565000 0.440000 1.795000 1.300000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.975000 1.180000 2.305000 1.550000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.377200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.125000 1.800000 2.770000 1.970000 ;
        RECT 1.125000 1.970000 1.455000 2.980000 ;
        RECT 2.045000 0.440000 2.770000 1.010000 ;
        RECT 2.205000 1.970000 2.770000 2.980000 ;
        RECT 2.595000 1.010000 2.770000 1.800000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.115000  1.950000 0.365000 3.245000 ;
      RECT 0.135000  0.350000 0.465000 0.960000 ;
      RECT 0.135000  0.960000 1.395000 1.130000 ;
      RECT 0.635000  0.085000 0.965000 0.780000 ;
      RECT 1.145000  0.350000 1.395000 0.960000 ;
      RECT 1.705000  2.140000 2.035000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_ms__o211ai_1
END LIBRARY

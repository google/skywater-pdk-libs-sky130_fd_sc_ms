* File: sky130_fd_sc_ms__nor3_1.spice
* Created: Wed Sep  2 12:15:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nor3_1.pex.spice"
.subckt sky130_fd_sc_ms__nor3_1  VNB VPB A B C VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_Y_M1003_d N_A_M1003_g N_VGND_M1003_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0.396 M=1 R=4.93333 SA=75000.2 SB=75001.1
+ A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_B_M1004_g N_Y_M1003_d VNB NLOWVT L=0.15 W=0.74 AD=0.1295
+ AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1002 N_Y_M1002_d N_C_M1002_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1001 A_117_368# N_A_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1.12 AD=0.1344
+ AS=0.3024 PD=1.36 PS=2.78 NRD=11.426 NRS=0 M=1 R=6.22222 SA=90000.2 SB=90001.1
+ A=0.2016 P=2.6 MULT=1
MM1005 A_201_368# N_B_M1005_g A_117_368# VPB PSHORT L=0.18 W=1.12 AD=0.1848
+ AS=0.1344 PD=1.45 PS=1.36 NRD=19.3454 NRS=11.426 M=1 R=6.22222 SA=90000.6
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1000 N_Y_M1000_d N_C_M1000_g A_201_368# VPB PSHORT L=0.18 W=1.12 AD=0.3024
+ AS=0.1848 PD=2.78 PS=1.45 NRD=0 NRS=19.3454 M=1 R=6.22222 SA=90001.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.278 P=8.32
*
.include "sky130_fd_sc_ms__nor3_1.pxi.spice"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_701_463# a_299_387# a_791_463# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X1 a_1471_493# a_1518_203# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X2 a_1518_203# a_1266_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X3 VGND a_1266_74# a_1867_409# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X4 a_299_387# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_833_400# a_493_387# a_1266_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 a_299_387# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 VGND a_701_463# a_833_400# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 Q a_1867_409# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X9 a_791_463# a_833_400# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X10 Q a_1867_409# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X11 VGND RESET_B a_1656_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X12 a_30_78# a_493_387# a_701_463# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X13 a_1656_81# a_1266_74# a_1518_203# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X14 VPWR RESET_B a_1518_203# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X15 a_894_138# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X16 a_30_78# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X17 VPWR a_701_463# a_833_400# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X18 VPWR RESET_B a_701_463# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X19 VPWR a_299_387# a_493_387# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X20 VPWR a_1266_74# a_1867_409# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X21 a_117_78# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X22 a_30_78# D a_117_78# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X23 a_30_78# a_299_387# a_701_463# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X24 a_833_400# a_299_387# a_1266_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X25 VGND a_299_387# a_493_387# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X26 a_701_463# a_493_387# a_821_138# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X27 a_1476_81# a_1518_203# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X28 a_1266_74# a_493_387# a_1471_493# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X29 a_821_138# a_833_400# a_894_138# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X30 VPWR D a_30_78# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X31 a_1266_74# a_299_387# a_1476_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
.ends

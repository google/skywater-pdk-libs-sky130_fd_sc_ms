* File: sky130_fd_sc_ms__fa_4.pxi.spice
* Created: Wed Sep  2 12:09:18 2020
* 
x_PM_SKY130_FD_SC_MS__FA_4%B N_B_M1017_g N_B_M1030_g N_B_M1026_g N_B_M1029_g
+ N_B_M1033_g N_B_M1012_g N_B_M1031_g N_B_M1039_g N_B_c_193_n N_B_c_204_n
+ N_B_c_216_p N_B_c_292_p N_B_c_194_n N_B_c_195_n N_B_c_222_p N_B_c_207_n
+ N_B_c_196_n N_B_c_316_p N_B_c_209_n B B N_B_c_198_n N_B_c_199_n
+ PM_SKY130_FD_SC_MS__FA_4%B
x_PM_SKY130_FD_SC_MS__FA_4%CIN N_CIN_M1001_g N_CIN_M1027_g N_CIN_M1032_g
+ N_CIN_M1006_g N_CIN_M1009_g N_CIN_M1028_g N_CIN_c_422_n N_CIN_c_423_n
+ N_CIN_c_424_n N_CIN_c_425_n N_CIN_c_426_n N_CIN_c_427_n N_CIN_c_428_n
+ N_CIN_c_429_n CIN N_CIN_c_430_n N_CIN_c_431_n N_CIN_c_432_n N_CIN_c_433_n
+ N_CIN_c_434_n N_CIN_c_435_n PM_SKY130_FD_SC_MS__FA_4%CIN
x_PM_SKY130_FD_SC_MS__FA_4%A_418_74# N_A_418_74#_M1001_d N_A_418_74#_M1027_d
+ N_A_418_74#_M1016_g N_A_418_74#_M1013_g N_A_418_74#_M1000_g
+ N_A_418_74#_M1011_g N_A_418_74#_M1019_g N_A_418_74#_M1014_g
+ N_A_418_74#_M1021_g N_A_418_74#_M1025_g N_A_418_74#_M1023_g
+ N_A_418_74#_M1037_g N_A_418_74#_c_590_n N_A_418_74#_c_685_p
+ N_A_418_74#_c_614_n N_A_418_74#_c_617_n N_A_418_74#_c_619_n
+ N_A_418_74#_c_651_n N_A_418_74#_c_591_n N_A_418_74#_c_621_n
+ N_A_418_74#_c_657_n N_A_418_74#_c_592_n N_A_418_74#_c_593_n
+ N_A_418_74#_c_628_n N_A_418_74#_c_696_p N_A_418_74#_c_629_n
+ N_A_418_74#_c_594_n N_A_418_74#_c_595_n N_A_418_74#_c_777_p
+ N_A_418_74#_c_630_n N_A_418_74#_c_634_n N_A_418_74#_c_637_n
+ N_A_418_74#_c_660_n N_A_418_74#_c_606_n N_A_418_74#_c_641_n
+ N_A_418_74#_c_644_n N_A_418_74#_c_596_n N_A_418_74#_c_597_n
+ N_A_418_74#_c_598_n N_A_418_74#_c_599_n PM_SKY130_FD_SC_MS__FA_4%A_418_74#
x_PM_SKY130_FD_SC_MS__FA_4%A N_A_M1003_g N_A_M1034_g N_A_c_889_n N_A_c_890_n
+ N_A_c_878_n N_A_M1005_g N_A_M1035_g N_A_c_892_n N_A_M1015_g N_A_c_880_n
+ N_A_M1004_g N_A_c_894_n N_A_M1002_g N_A_c_883_n N_A_M1018_g N_A_c_884_n
+ N_A_c_898_n N_A_c_885_n N_A_c_899_n A A N_A_c_887_n PM_SKY130_FD_SC_MS__FA_4%A
x_PM_SKY130_FD_SC_MS__FA_4%A_1024_74# N_A_1024_74#_M1016_d N_A_1024_74#_M1013_d
+ N_A_1024_74#_M1007_g N_A_1024_74#_M1022_g N_A_1024_74#_M1008_g
+ N_A_1024_74#_M1024_g N_A_1024_74#_M1010_g N_A_1024_74#_M1036_g
+ N_A_1024_74#_M1020_g N_A_1024_74#_M1038_g N_A_1024_74#_c_1053_n
+ N_A_1024_74#_c_1056_n N_A_1024_74#_c_1059_n N_A_1024_74#_c_1040_n
+ N_A_1024_74#_c_1048_n N_A_1024_74#_c_1041_n N_A_1024_74#_c_1050_n
+ N_A_1024_74#_c_1064_n N_A_1024_74#_c_1077_n N_A_1024_74#_c_1065_n
+ N_A_1024_74#_c_1067_n N_A_1024_74#_c_1042_n N_A_1024_74#_c_1043_n
+ PM_SKY130_FD_SC_MS__FA_4%A_1024_74#
x_PM_SKY130_FD_SC_MS__FA_4%A_27_392# N_A_27_392#_M1003_s N_A_27_392#_M1017_d
+ N_A_27_392#_c_1193_n N_A_27_392#_c_1194_n N_A_27_392#_c_1202_n
+ N_A_27_392#_c_1203_n N_A_27_392#_c_1195_n N_A_27_392#_c_1196_n
+ PM_SKY130_FD_SC_MS__FA_4%A_27_392#
x_PM_SKY130_FD_SC_MS__FA_4%VPWR N_VPWR_M1003_d N_VPWR_M1005_d N_VPWR_M1012_d
+ N_VPWR_M1018_d N_VPWR_M1008_s N_VPWR_M1020_s N_VPWR_M1019_d N_VPWR_M1023_d
+ N_VPWR_c_1242_n N_VPWR_c_1243_n N_VPWR_c_1244_n N_VPWR_c_1245_n
+ N_VPWR_c_1246_n N_VPWR_c_1247_n N_VPWR_c_1248_n N_VPWR_c_1249_n
+ N_VPWR_c_1250_n N_VPWR_c_1251_n N_VPWR_c_1252_n VPWR N_VPWR_c_1253_n
+ N_VPWR_c_1254_n N_VPWR_c_1255_n N_VPWR_c_1256_n N_VPWR_c_1257_n
+ N_VPWR_c_1258_n N_VPWR_c_1259_n N_VPWR_c_1260_n N_VPWR_c_1261_n
+ N_VPWR_c_1262_n N_VPWR_c_1263_n N_VPWR_c_1264_n N_VPWR_c_1241_n
+ PM_SKY130_FD_SC_MS__FA_4%VPWR
x_PM_SKY130_FD_SC_MS__FA_4%A_740_347# N_A_740_347#_M1006_d N_A_740_347#_M1004_d
+ N_A_740_347#_c_1390_n N_A_740_347#_c_1394_n N_A_740_347#_c_1386_n
+ N_A_740_347#_c_1387_n PM_SKY130_FD_SC_MS__FA_4%A_740_347#
x_PM_SKY130_FD_SC_MS__FA_4%SUM N_SUM_M1022_s N_SUM_M1036_s N_SUM_M1007_d
+ N_SUM_M1010_d N_SUM_c_1426_n N_SUM_c_1427_n N_SUM_c_1423_n N_SUM_c_1454_n
+ N_SUM_c_1424_n N_SUM_c_1425_n SUM SUM SUM SUM PM_SKY130_FD_SC_MS__FA_4%SUM
x_PM_SKY130_FD_SC_MS__FA_4%COUT N_COUT_M1011_d N_COUT_M1025_d N_COUT_M1000_s
+ N_COUT_M1021_s N_COUT_c_1488_n N_COUT_c_1489_n N_COUT_c_1484_n N_COUT_c_1490_n
+ N_COUT_c_1506_n N_COUT_c_1485_n N_COUT_c_1486_n N_COUT_c_1487_n
+ N_COUT_c_1521_n COUT COUT COUT COUT N_COUT_c_1491_n COUT
+ PM_SKY130_FD_SC_MS__FA_4%COUT
x_PM_SKY130_FD_SC_MS__FA_4%A_27_74# N_A_27_74#_M1034_s N_A_27_74#_M1030_d
+ N_A_27_74#_c_1553_n N_A_27_74#_c_1554_n N_A_27_74#_c_1557_n
+ N_A_27_74#_c_1555_n PM_SKY130_FD_SC_MS__FA_4%A_27_74#
x_PM_SKY130_FD_SC_MS__FA_4%VGND N_VGND_M1034_d N_VGND_M1035_d N_VGND_M1033_d
+ N_VGND_M1002_d N_VGND_M1024_d N_VGND_M1038_d N_VGND_M1014_s N_VGND_M1037_s
+ N_VGND_c_1585_n N_VGND_c_1586_n N_VGND_c_1587_n N_VGND_c_1588_n
+ N_VGND_c_1589_n N_VGND_c_1590_n N_VGND_c_1591_n N_VGND_c_1592_n VGND
+ N_VGND_c_1593_n N_VGND_c_1594_n N_VGND_c_1595_n N_VGND_c_1596_n
+ N_VGND_c_1597_n N_VGND_c_1598_n N_VGND_c_1599_n N_VGND_c_1600_n
+ N_VGND_c_1601_n N_VGND_c_1602_n N_VGND_c_1603_n N_VGND_c_1604_n
+ PM_SKY130_FD_SC_MS__FA_4%VGND
x_PM_SKY130_FD_SC_MS__FA_4%A_734_74# N_A_734_74#_M1032_d N_A_734_74#_M1015_d
+ N_A_734_74#_c_1734_n N_A_734_74#_c_1732_n N_A_734_74#_c_1733_n
+ PM_SKY130_FD_SC_MS__FA_4%A_734_74#
cc_1 VNB N_B_M1030_g 0.0209127f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=0.74
cc_2 VNB N_B_M1026_g 0.0210869f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=0.74
cc_3 VNB N_B_M1033_g 0.0203825f $X=-0.19 $Y=-0.245 $X2=4.025 $Y2=0.74
cc_4 VNB N_B_M1039_g 0.0183203f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=0.74
cc_5 VNB N_B_c_193_n 0.00309095f $X=-0.19 $Y=-0.245 $X2=1.665 $Y2=1.417
cc_6 VNB N_B_c_194_n 8.09421e-19 $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.41
cc_7 VNB N_B_c_195_n 0.0248536f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.41
cc_8 VNB N_B_c_196_n 0.0265504f $X=-0.19 $Y=-0.245 $X2=4.115 $Y2=1.41
cc_9 VNB B 0.00826485f $X=-0.19 $Y=-0.245 $X2=6.395 $Y2=1.58
cc_10 VNB N_B_c_198_n 0.0397424f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=1.41
cc_11 VNB N_B_c_199_n 0.0217419f $X=-0.19 $Y=-0.245 $X2=6.175 $Y2=1.41
cc_12 VNB N_CIN_M1032_g 0.019466f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=0.74
cc_13 VNB N_CIN_c_422_n 0.0025906f $X=-0.19 $Y=-0.245 $X2=6.1 $Y2=1.575
cc_14 VNB N_CIN_c_423_n 0.0232814f $X=-0.19 $Y=-0.245 $X2=6.1 $Y2=2.235
cc_15 VNB N_CIN_c_424_n 0.0071807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_CIN_c_425_n 0.00290723f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=1.245
cc_17 VNB N_CIN_c_426_n 0.018935f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=0.74
cc_18 VNB N_CIN_c_427_n 0.00298431f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=0.74
cc_19 VNB N_CIN_c_428_n 0.00460694f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.41
cc_20 VNB N_CIN_c_429_n 0.00274216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_CIN_c_430_n 0.0307256f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.745
cc_22 VNB N_CIN_c_431_n 0.018815f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.41
cc_23 VNB N_CIN_c_432_n 0.0293303f $X=-0.19 $Y=-0.245 $X2=4.115 $Y2=1.41
cc_24 VNB N_CIN_c_433_n 0.0178512f $X=-0.19 $Y=-0.245 $X2=4.115 $Y2=1.41
cc_25 VNB N_CIN_c_434_n 0.00310764f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=2.035
cc_26 VNB N_CIN_c_435_n 0.00361772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_418_74#_M1000_g 5.11652e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_418_74#_M1011_g 0.0209667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_418_74#_M1019_g 4.96731e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_418_74#_M1014_g 0.0185701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_418_74#_M1021_g 4.9443e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_418_74#_M1025_g 0.0182888f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.41
cc_33 VNB N_A_418_74#_M1023_g 7.19436e-19 $X=-0.19 $Y=-0.245 $X2=2.48 $Y2=2.035
cc_34 VNB N_A_418_74#_M1037_g 0.0251724f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.41
cc_35 VNB N_A_418_74#_c_590_n 0.00500716f $X=-0.19 $Y=-0.245 $X2=3.95 $Y2=1.83
cc_36 VNB N_A_418_74#_c_591_n 0.00333942f $X=-0.19 $Y=-0.245 $X2=5.915 $Y2=1.58
cc_37 VNB N_A_418_74#_c_592_n 0.00802253f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=1.41
cc_38 VNB N_A_418_74#_c_593_n 9.82756e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_418_74#_c_594_n 0.00296963f $X=-0.19 $Y=-0.245 $X2=4.115 $Y2=1.575
cc_40 VNB N_A_418_74#_c_595_n 0.00392926f $X=-0.19 $Y=-0.245 $X2=6.175 $Y2=1.41
cc_41 VNB N_A_418_74#_c_596_n 0.00879717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_418_74#_c_597_n 0.0276885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_418_74#_c_598_n 0.0177385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_418_74#_c_599_n 0.104376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_M1003_g 0.00400194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_M1034_g 0.0277073f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=0.74
cc_47 VNB N_A_c_878_n 0.005061f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=0.74
cc_48 VNB N_A_M1005_g 0.0110176f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=2.235
cc_49 VNB N_A_c_880_n 0.00549706f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=2.235
cc_50 VNB N_A_M1004_g 0.0140582f $X=-0.19 $Y=-0.245 $X2=6.1 $Y2=2.235
cc_51 VNB N_A_M1002_g 0.0403652f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=0.74
cc_52 VNB N_A_c_883_n 0.00252311f $X=-0.19 $Y=-0.245 $X2=1.665 $Y2=1.417
cc_53 VNB N_A_c_884_n 0.0161869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_c_885_n 0.0169826f $X=-0.19 $Y=-0.245 $X2=1.75 $Y2=1.95
cc_55 VNB A 0.0194965f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.41
cc_56 VNB N_A_c_887_n 0.0599934f $X=-0.19 $Y=-0.245 $X2=4.115 $Y2=1.41
cc_57 VNB N_A_1024_74#_M1022_g 0.0221413f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=1.575
cc_58 VNB N_A_1024_74#_M1024_g 0.0217363f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=1.575
cc_59 VNB N_A_1024_74#_M1036_g 0.0210584f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=1.245
cc_60 VNB N_A_1024_74#_M1038_g 0.0220203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1024_74#_c_1040_n 0.00361783f $X=-0.19 $Y=-0.245 $X2=4.115
+ $Y2=1.41
cc_62 VNB N_A_1024_74#_c_1041_n 3.03738e-19 $X=-0.19 $Y=-0.245 $X2=5.915
+ $Y2=1.58
cc_63 VNB N_A_1024_74#_c_1042_n 0.0029978f $X=-0.19 $Y=-0.245 $X2=6.175 $Y2=1.41
cc_64 VNB N_A_1024_74#_c_1043_n 0.0833164f $X=-0.19 $Y=-0.245 $X2=6.175
+ $Y2=1.575
cc_65 VNB N_VPWR_c_1241_n 0.462217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_SUM_c_1423_n 0.00586669f $X=-0.19 $Y=-0.245 $X2=4.025 $Y2=1.245
cc_67 VNB N_SUM_c_1424_n 0.00234369f $X=-0.19 $Y=-0.245 $X2=4.06 $Y2=2.235
cc_68 VNB N_SUM_c_1425_n 0.00137885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_COUT_c_1484_n 0.00220089f $X=-0.19 $Y=-0.245 $X2=4.025 $Y2=0.74
cc_70 VNB N_COUT_c_1485_n 0.00123375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_COUT_c_1486_n 0.00229206f $X=-0.19 $Y=-0.245 $X2=6.1 $Y2=2.235
cc_72 VNB N_COUT_c_1487_n 0.00154258f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=0.74
cc_73 VNB N_A_27_74#_c_1553_n 0.00249128f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=0.74
cc_74 VNB N_A_27_74#_c_1554_n 0.0306363f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=2.235
cc_75 VNB N_A_27_74#_c_1555_n 0.00162437f $X=-0.19 $Y=-0.245 $X2=4.025 $Y2=0.74
cc_76 VNB N_VGND_c_1585_n 0.00574325f $X=-0.19 $Y=-0.245 $X2=6.1 $Y2=2.235
cc_77 VNB N_VGND_c_1586_n 0.00546039f $X=-0.19 $Y=-0.245 $X2=6.115 $Y2=0.74
cc_78 VNB N_VGND_c_1587_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=1.665 $Y2=1.417
cc_79 VNB N_VGND_c_1588_n 0.0471419f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=1.41
cc_80 VNB N_VGND_c_1589_n 0.0556692f $X=-0.19 $Y=-0.245 $X2=1.75 $Y2=1.575
cc_81 VNB N_VGND_c_1590_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=1.75 $Y2=1.95
cc_82 VNB N_VGND_c_1591_n 0.0133472f $X=-0.19 $Y=-0.245 $X2=2.48 $Y2=2.035
cc_83 VNB N_VGND_c_1592_n 0.0178103f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=2.035
cc_84 VNB N_VGND_c_1593_n 0.0547728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1594_n 0.0185379f $X=-0.19 $Y=-0.245 $X2=4.115 $Y2=1.41
cc_86 VNB N_VGND_c_1595_n 0.0185379f $X=-0.19 $Y=-0.245 $X2=6.175 $Y2=1.41
cc_87 VNB N_VGND_c_1596_n 0.0175388f $X=-0.19 $Y=-0.245 $X2=6 $Y2=1.575
cc_88 VNB N_VGND_c_1597_n 0.0174844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1598_n 0.0185699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1599_n 0.01914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1600_n 0.0153962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1601_n 0.0170767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1602_n 0.015362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1603_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1604_n 0.579257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_734_74#_c_1732_n 0.00205545f $X=-0.19 $Y=-0.245 $X2=2.585 $Y2=0.74
cc_97 VNB N_A_734_74#_c_1733_n 0.00203932f $X=-0.19 $Y=-0.245 $X2=2.6 $Y2=2.235
cc_98 VPB N_B_M1017_g 0.0217243f $X=-0.19 $Y=1.66 $X2=1.155 $Y2=2.235
cc_99 VPB N_B_M1029_g 0.0180821f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=2.235
cc_100 VPB N_B_M1012_g 0.0185879f $X=-0.19 $Y=1.66 $X2=4.06 $Y2=2.235
cc_101 VPB N_B_M1031_g 0.0187565f $X=-0.19 $Y=1.66 $X2=6.1 $Y2=2.235
cc_102 VPB N_B_c_204_n 0.00259536f $X=-0.19 $Y=1.66 $X2=1.75 $Y2=1.95
cc_103 VPB N_B_c_194_n 0.00277573f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=1.41
cc_104 VPB N_B_c_195_n 0.00560327f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=1.41
cc_105 VPB N_B_c_207_n 0.00344703f $X=-0.19 $Y=1.66 $X2=4.115 $Y2=1.41
cc_106 VPB N_B_c_196_n 0.0056223f $X=-0.19 $Y=1.66 $X2=4.115 $Y2=1.41
cc_107 VPB N_B_c_209_n 0.00127169f $X=-0.19 $Y=1.66 $X2=4.62 $Y2=1.805
cc_108 VPB B 0.0111341f $X=-0.19 $Y=1.66 $X2=5.915 $Y2=1.58
cc_109 VPB B 0.00292356f $X=-0.19 $Y=1.66 $X2=6.395 $Y2=1.58
cc_110 VPB N_B_c_198_n 0.0174804f $X=-0.19 $Y=1.66 $X2=1.585 $Y2=1.41
cc_111 VPB N_B_c_199_n 0.0054384f $X=-0.19 $Y=1.66 $X2=6.175 $Y2=1.41
cc_112 VPB N_CIN_M1027_g 0.0212926f $X=-0.19 $Y=1.66 $X2=1.585 $Y2=0.74
cc_113 VPB N_CIN_M1006_g 0.0198206f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=2.235
cc_114 VPB N_CIN_M1009_g 0.0211116f $X=-0.19 $Y=1.66 $X2=4.025 $Y2=0.74
cc_115 VPB N_CIN_c_422_n 0.00192839f $X=-0.19 $Y=1.66 $X2=6.1 $Y2=1.575
cc_116 VPB N_CIN_c_423_n 0.00471211f $X=-0.19 $Y=1.66 $X2=6.1 $Y2=2.235
cc_117 VPB N_CIN_c_434_n 0.00278862f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=2.035
cc_118 VPB N_CIN_c_435_n 4.02791e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_418_74#_M1013_g 0.0214796f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_418_74#_M1000_g 0.0234399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_418_74#_M1019_g 0.0228127f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_418_74#_M1021_g 0.0227905f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_418_74#_M1023_g 0.0274184f $X=-0.19 $Y=1.66 $X2=2.48 $Y2=2.035
cc_124 VPB N_A_418_74#_c_590_n 0.00142531f $X=-0.19 $Y=1.66 $X2=3.95 $Y2=1.83
cc_125 VPB N_A_418_74#_c_606_n 0.00217873f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_M1003_g 0.0328377f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_c_889_n 0.17793f $X=-0.19 $Y=1.66 $X2=2.585 $Y2=1.245
cc_128 VPB N_A_c_890_n 0.0143041f $X=-0.19 $Y=1.66 $X2=2.585 $Y2=0.74
cc_129 VPB N_A_M1005_g 0.0376301f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=2.235
cc_130 VPB N_A_c_892_n 0.0915019f $X=-0.19 $Y=1.66 $X2=4.025 $Y2=0.74
cc_131 VPB N_A_M1004_g 0.0383822f $X=-0.19 $Y=1.66 $X2=6.1 $Y2=2.235
cc_132 VPB N_A_c_894_n 0.154052f $X=-0.19 $Y=1.66 $X2=6.1 $Y2=2.235
cc_133 VPB N_A_M1002_g 0.00127901f $X=-0.19 $Y=1.66 $X2=6.115 $Y2=0.74
cc_134 VPB N_A_c_883_n 0.00364873f $X=-0.19 $Y=1.66 $X2=1.665 $Y2=1.417
cc_135 VPB N_A_M1018_g 0.0281783f $X=-0.19 $Y=1.66 $X2=1.51 $Y2=1.41
cc_136 VPB N_A_c_898_n 0.0087959f $X=-0.19 $Y=1.66 $X2=1.75 $Y2=1.575
cc_137 VPB N_A_c_899_n 0.0087959f $X=-0.19 $Y=1.66 $X2=2.48 $Y2=2.035
cc_138 VPB A 0.0114306f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=1.41
cc_139 VPB N_A_c_887_n 0.00515871f $X=-0.19 $Y=1.66 $X2=4.115 $Y2=1.41
cc_140 VPB N_A_1024_74#_M1007_g 0.0232745f $X=-0.19 $Y=1.66 $X2=2.585 $Y2=1.245
cc_141 VPB N_A_1024_74#_M1008_g 0.0223736f $X=-0.19 $Y=1.66 $X2=4.025 $Y2=1.245
cc_142 VPB N_A_1024_74#_M1010_g 0.0223369f $X=-0.19 $Y=1.66 $X2=6.1 $Y2=1.575
cc_143 VPB N_A_1024_74#_M1020_g 0.022202f $X=-0.19 $Y=1.66 $X2=1.665 $Y2=1.417
cc_144 VPB N_A_1024_74#_c_1048_n 0.00294257f $X=-0.19 $Y=1.66 $X2=4.115 $Y2=1.41
cc_145 VPB N_A_1024_74#_c_1041_n 7.08103e-19 $X=-0.19 $Y=1.66 $X2=5.915 $Y2=1.58
cc_146 VPB N_A_1024_74#_c_1050_n 0.00262534f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_1024_74#_c_1043_n 0.0101968f $X=-0.19 $Y=1.66 $X2=6.175 $Y2=1.575
cc_148 VPB N_A_27_392#_c_1193_n 0.0146163f $X=-0.19 $Y=1.66 $X2=1.585 $Y2=0.74
cc_149 VPB N_A_27_392#_c_1194_n 0.0301301f $X=-0.19 $Y=1.66 $X2=2.585 $Y2=1.245
cc_150 VPB N_A_27_392#_c_1195_n 0.00249638f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=2.235
cc_151 VPB N_A_27_392#_c_1196_n 0.0103364f $X=-0.19 $Y=1.66 $X2=4.025 $Y2=0.74
cc_152 VPB N_VPWR_c_1242_n 0.00768987f $X=-0.19 $Y=1.66 $X2=6.115 $Y2=1.245
cc_153 VPB N_VPWR_c_1243_n 0.00532246f $X=-0.19 $Y=1.66 $X2=1.665 $Y2=1.417
cc_154 VPB N_VPWR_c_1244_n 0.00573745f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_1245_n 0.0102279f $X=-0.19 $Y=1.66 $X2=1.835 $Y2=2.035
cc_156 VPB N_VPWR_c_1246_n 0.00884785f $X=-0.19 $Y=1.66 $X2=3.95 $Y2=1.83
cc_157 VPB N_VPWR_c_1247_n 0.018624f $X=-0.19 $Y=1.66 $X2=4.115 $Y2=1.41
cc_158 VPB N_VPWR_c_1248_n 0.00884785f $X=-0.19 $Y=1.66 $X2=4.115 $Y2=1.817
cc_159 VPB N_VPWR_c_1249_n 0.012247f $X=-0.19 $Y=1.66 $X2=6.395 $Y2=1.58
cc_160 VPB N_VPWR_c_1250_n 0.0586854f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_1251_n 0.0634767f $X=-0.19 $Y=1.66 $X2=1.585 $Y2=1.41
cc_162 VPB N_VPWR_c_1252_n 0.00436868f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_1253_n 0.0175187f $X=-0.19 $Y=1.66 $X2=6.175 $Y2=1.245
cc_164 VPB N_VPWR_c_1254_n 0.0664038f $X=-0.19 $Y=1.66 $X2=6 $Y2=1.575
cc_165 VPB N_VPWR_c_1255_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_1256_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_1257_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_1258_n 0.0195713f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_1259_n 0.0212973f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_1260_n 0.00530087f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_1261_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_1262_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_1263_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_1264_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_1241_n 0.0740968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_740_347#_c_1386_n 0.00290549f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=1.575
cc_177 VPB N_A_740_347#_c_1387_n 0.00219575f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_SUM_c_1426_n 0.00117235f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=1.575
cc_179 VPB N_SUM_c_1427_n 0.00231613f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=2.235
cc_180 VPB N_SUM_c_1425_n 0.00160343f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB SUM 0.00231613f $X=-0.19 $Y=1.66 $X2=1.75 $Y2=1.575
cc_182 VPB N_COUT_c_1488_n 0.00224287f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=1.575
cc_183 VPB N_COUT_c_1489_n 0.00231613f $X=-0.19 $Y=1.66 $X2=2.6 $Y2=2.235
cc_184 VPB N_COUT_c_1490_n 0.00249468f $X=-0.19 $Y=1.66 $X2=4.06 $Y2=1.575
cc_185 VPB N_COUT_c_1491_n 0.00214167f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=1.41
cc_186 VPB COUT 0.00231613f $X=-0.19 $Y=1.66 $X2=2.645 $Y2=1.41
cc_187 N_B_M1029_g N_CIN_M1027_g 0.0431055f $X=2.6 $Y=2.235 $X2=0 $Y2=0
cc_188 N_B_c_204_n N_CIN_M1027_g 0.00513554f $X=1.75 $Y=1.95 $X2=0 $Y2=0
cc_189 N_B_c_216_p N_CIN_M1027_g 0.0132486f $X=2.48 $Y=2.035 $X2=0 $Y2=0
cc_190 N_B_c_194_n N_CIN_M1027_g 5.73116e-19 $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_191 N_B_c_195_n N_CIN_M1027_g 0.00129392f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_192 N_B_c_198_n N_CIN_M1027_g 7.23203e-19 $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_193 N_B_M1033_g N_CIN_M1032_g 0.0293113f $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_194 N_B_M1012_g N_CIN_M1006_g 0.025979f $X=4.06 $Y=2.235 $X2=0 $Y2=0
cc_195 N_B_c_222_p N_CIN_M1006_g 0.016421f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_196 N_B_c_207_n N_CIN_M1006_g 0.00343576f $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_197 B N_CIN_M1009_g 0.0119567f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_198 B N_CIN_M1009_g 0.00453099f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_199 N_B_c_199_n N_CIN_M1009_g 0.0589212f $X=6.175 $Y=1.41 $X2=0 $Y2=0
cc_200 N_B_c_207_n N_CIN_c_422_n 0.0194879f $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_201 N_B_c_196_n N_CIN_c_422_n 0.00108757f $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_202 N_B_c_222_p N_CIN_c_423_n 0.00234121f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_203 N_B_c_207_n N_CIN_c_423_n 4.68399e-19 $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_204 N_B_c_196_n N_CIN_c_423_n 0.0214173f $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_205 N_B_M1026_g N_CIN_c_424_n 0.00166151f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_206 N_B_c_216_p N_CIN_c_424_n 0.00534188f $X=2.48 $Y=2.035 $X2=0 $Y2=0
cc_207 N_B_c_194_n N_CIN_c_424_n 0.025012f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_208 N_B_c_195_n N_CIN_c_424_n 0.00263938f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_209 N_B_c_222_p N_CIN_c_424_n 0.00606814f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_210 N_B_M1026_g N_CIN_c_425_n 7.01969e-19 $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_211 N_B_c_193_n N_CIN_c_425_n 0.00117817f $X=1.665 $Y=1.417 $X2=0 $Y2=0
cc_212 N_B_c_216_p N_CIN_c_425_n 0.00191142f $X=2.48 $Y=2.035 $X2=0 $Y2=0
cc_213 N_B_c_194_n N_CIN_c_425_n 0.0013005f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_214 N_B_c_195_n N_CIN_c_425_n 6.81723e-19 $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_215 N_B_M1033_g N_CIN_c_426_n 0.00157687f $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_216 N_B_c_222_p N_CIN_c_426_n 0.00740196f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_217 N_B_c_207_n N_CIN_c_426_n 0.0245256f $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_218 N_B_c_196_n N_CIN_c_426_n 0.00277849f $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_219 N_B_c_209_n N_CIN_c_426_n 0.00815389f $X=4.62 $Y=1.805 $X2=0 $Y2=0
cc_220 B N_CIN_c_426_n 0.0132686f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_221 N_B_M1026_g N_CIN_c_427_n 6.4019e-19 $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_222 N_B_c_194_n N_CIN_c_427_n 0.00130776f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_223 N_B_c_195_n N_CIN_c_427_n 6.86607e-19 $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_224 N_B_c_222_p N_CIN_c_427_n 0.00247813f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_225 B N_CIN_c_428_n 0.00350418f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_226 B N_CIN_c_428_n 9.68406e-19 $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_227 N_B_M1039_g N_CIN_c_429_n 3.61499e-19 $X=6.115 $Y=0.74 $X2=0 $Y2=0
cc_228 B N_CIN_c_429_n 0.0222605f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_229 B N_CIN_c_429_n 0.0224776f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_230 N_B_c_199_n N_CIN_c_429_n 3.67751e-19 $X=6.175 $Y=1.41 $X2=0 $Y2=0
cc_231 N_B_M1026_g N_CIN_c_430_n 0.00136863f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_232 N_B_c_193_n N_CIN_c_430_n 0.00218231f $X=1.665 $Y=1.417 $X2=0 $Y2=0
cc_233 N_B_c_216_p N_CIN_c_430_n 0.0021066f $X=2.48 $Y=2.035 $X2=0 $Y2=0
cc_234 N_B_c_194_n N_CIN_c_430_n 4.64676e-19 $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_235 N_B_c_195_n N_CIN_c_430_n 0.0197774f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_236 N_B_c_198_n N_CIN_c_430_n 0.0141766f $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_237 N_B_M1030_g N_CIN_c_431_n 0.0288887f $X=1.585 $Y=0.74 $X2=0 $Y2=0
cc_238 N_B_M1026_g N_CIN_c_431_n 0.0240859f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_239 B N_CIN_c_432_n 0.00451129f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_240 B N_CIN_c_432_n 0.00187682f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_241 N_B_c_199_n N_CIN_c_432_n 0.0190182f $X=6.175 $Y=1.41 $X2=0 $Y2=0
cc_242 N_B_M1039_g N_CIN_c_433_n 0.0538055f $X=6.115 $Y=0.74 $X2=0 $Y2=0
cc_243 N_B_M1030_g N_CIN_c_434_n 3.51335e-19 $X=1.585 $Y=0.74 $X2=0 $Y2=0
cc_244 N_B_M1026_g N_CIN_c_434_n 0.00105583f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_245 N_B_M1029_g N_CIN_c_434_n 5.5793e-19 $X=2.6 $Y=2.235 $X2=0 $Y2=0
cc_246 N_B_c_193_n N_CIN_c_434_n 0.0243757f $X=1.665 $Y=1.417 $X2=0 $Y2=0
cc_247 N_B_c_204_n N_CIN_c_434_n 0.0140408f $X=1.75 $Y=1.95 $X2=0 $Y2=0
cc_248 N_B_c_216_p N_CIN_c_434_n 0.0131999f $X=2.48 $Y=2.035 $X2=0 $Y2=0
cc_249 N_B_c_194_n N_CIN_c_434_n 0.0317858f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_250 N_B_c_195_n N_CIN_c_434_n 0.00163291f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_251 N_B_c_198_n N_CIN_c_434_n 4.09781e-19 $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_252 N_B_M1026_g N_CIN_c_435_n 8.34658e-19 $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_253 N_B_c_194_n N_CIN_c_435_n 0.0223381f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_254 N_B_c_195_n N_CIN_c_435_n 0.00176431f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_255 N_B_c_222_p N_CIN_c_435_n 0.0460084f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_256 N_B_c_216_p N_A_418_74#_M1027_d 0.00476167f $X=2.48 $Y=2.035 $X2=0 $Y2=0
cc_257 B N_A_418_74#_M1013_g 0.016725f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_258 N_B_M1017_g N_A_418_74#_c_590_n 0.00665518f $X=1.155 $Y=2.235 $X2=0 $Y2=0
cc_259 N_B_M1030_g N_A_418_74#_c_590_n 0.00442274f $X=1.585 $Y=0.74 $X2=0 $Y2=0
cc_260 N_B_c_193_n N_A_418_74#_c_590_n 0.0232015f $X=1.665 $Y=1.417 $X2=0 $Y2=0
cc_261 N_B_c_204_n N_A_418_74#_c_590_n 0.0054586f $X=1.75 $Y=1.95 $X2=0 $Y2=0
cc_262 N_B_c_198_n N_A_418_74#_c_590_n 0.0120428f $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_263 N_B_M1017_g N_A_418_74#_c_614_n 0.0110718f $X=1.155 $Y=2.235 $X2=0 $Y2=0
cc_264 N_B_c_204_n N_A_418_74#_c_614_n 0.00250585f $X=1.75 $Y=1.95 $X2=0 $Y2=0
cc_265 N_B_c_292_p N_A_418_74#_c_614_n 0.0138309f $X=1.835 $Y=2.035 $X2=0 $Y2=0
cc_266 N_B_c_216_p N_A_418_74#_c_617_n 0.0223331f $X=2.48 $Y=2.035 $X2=0 $Y2=0
cc_267 N_B_c_292_p N_A_418_74#_c_617_n 0.0137412f $X=1.835 $Y=2.035 $X2=0 $Y2=0
cc_268 N_B_M1017_g N_A_418_74#_c_619_n 0.00392884f $X=1.155 $Y=2.235 $X2=0 $Y2=0
cc_269 N_B_M1026_g N_A_418_74#_c_591_n 0.00341585f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_270 N_B_M1033_g N_A_418_74#_c_621_n 0.0110518f $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_271 N_B_c_222_p N_A_418_74#_c_621_n 0.00159983f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_272 N_B_c_207_n N_A_418_74#_c_621_n 0.0184553f $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_273 N_B_c_196_n N_A_418_74#_c_621_n 0.00310854f $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_274 N_B_c_209_n N_A_418_74#_c_621_n 0.0032782f $X=4.62 $Y=1.805 $X2=0 $Y2=0
cc_275 B N_A_418_74#_c_621_n 0.00298874f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_276 N_B_M1039_g N_A_418_74#_c_592_n 0.0102703f $X=6.115 $Y=0.74 $X2=0 $Y2=0
cc_277 N_B_M1039_g N_A_418_74#_c_628_n 0.00376916f $X=6.115 $Y=0.74 $X2=0 $Y2=0
cc_278 N_B_M1039_g N_A_418_74#_c_629_n 0.00295923f $X=6.115 $Y=0.74 $X2=0 $Y2=0
cc_279 N_B_M1017_g N_A_418_74#_c_630_n 0.0148813f $X=1.155 $Y=2.235 $X2=0 $Y2=0
cc_280 N_B_c_193_n N_A_418_74#_c_630_n 0.0110357f $X=1.665 $Y=1.417 $X2=0 $Y2=0
cc_281 N_B_c_204_n N_A_418_74#_c_630_n 0.0133105f $X=1.75 $Y=1.95 $X2=0 $Y2=0
cc_282 N_B_c_198_n N_A_418_74#_c_630_n 0.00568662f $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_283 N_B_M1030_g N_A_418_74#_c_634_n 0.0124111f $X=1.585 $Y=0.74 $X2=0 $Y2=0
cc_284 N_B_c_193_n N_A_418_74#_c_634_n 0.0208902f $X=1.665 $Y=1.417 $X2=0 $Y2=0
cc_285 N_B_c_198_n N_A_418_74#_c_634_n 0.00862669f $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_286 N_B_c_193_n N_A_418_74#_c_637_n 0.0124459f $X=1.665 $Y=1.417 $X2=0 $Y2=0
cc_287 N_B_M1029_g N_A_418_74#_c_606_n 0.0114661f $X=2.6 $Y=2.235 $X2=0 $Y2=0
cc_288 N_B_c_216_p N_A_418_74#_c_606_n 0.0144089f $X=2.48 $Y=2.035 $X2=0 $Y2=0
cc_289 N_B_c_316_p N_A_418_74#_c_606_n 0.00234595f $X=2.645 $Y=1.83 $X2=0 $Y2=0
cc_290 N_B_M1026_g N_A_418_74#_c_641_n 0.0133548f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_291 N_B_c_194_n N_A_418_74#_c_641_n 0.0122929f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_292 N_B_c_195_n N_A_418_74#_c_641_n 8.31105e-19 $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_293 N_B_M1033_g N_A_418_74#_c_644_n 3.88992e-19 $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_294 N_B_c_207_n N_A_418_74#_c_596_n 0.00547767f $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_295 B N_A_418_74#_c_596_n 0.0242486f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_296 B N_A_418_74#_c_597_n 0.00105083f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_297 N_B_M1017_g N_A_M1003_g 0.0223878f $X=1.155 $Y=2.235 $X2=0 $Y2=0
cc_298 N_B_M1017_g N_A_c_889_n 0.0106216f $X=1.155 $Y=2.235 $X2=0 $Y2=0
cc_299 N_B_M1029_g N_A_c_889_n 0.0123594f $X=2.6 $Y=2.235 $X2=0 $Y2=0
cc_300 N_B_M1026_g N_A_c_878_n 0.00188318f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_301 N_B_c_194_n N_A_c_878_n 4.83088e-19 $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_302 N_B_c_195_n N_A_c_878_n 0.0212349f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_303 N_B_M1029_g N_A_M1005_g 0.0468834f $X=2.6 $Y=2.235 $X2=0 $Y2=0
cc_304 N_B_c_194_n N_A_M1005_g 0.0039036f $X=2.645 $Y=1.41 $X2=0 $Y2=0
cc_305 N_B_c_222_p N_A_M1005_g 0.0167804f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_306 N_B_c_316_p N_A_M1005_g 0.00109021f $X=2.645 $Y=1.83 $X2=0 $Y2=0
cc_307 N_B_M1012_g N_A_c_892_n 0.0123594f $X=4.06 $Y=2.235 $X2=0 $Y2=0
cc_308 N_B_c_207_n N_A_c_880_n 0.00146089f $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_309 N_B_c_196_n N_A_c_880_n 0.0169501f $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_310 N_B_M1012_g N_A_M1004_g 0.0320637f $X=4.06 $Y=2.235 $X2=0 $Y2=0
cc_311 N_B_c_207_n N_A_M1004_g 0.00330365f $X=4.115 $Y=1.41 $X2=0 $Y2=0
cc_312 N_B_c_209_n N_A_M1004_g 0.00788898f $X=4.62 $Y=1.805 $X2=0 $Y2=0
cc_313 B N_A_M1004_g 0.00774307f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_314 N_B_M1031_g N_A_c_894_n 0.0124996f $X=6.1 $Y=2.235 $X2=0 $Y2=0
cc_315 N_B_M1031_g N_A_M1002_g 0.0451757f $X=6.1 $Y=2.235 $X2=0 $Y2=0
cc_316 N_B_M1039_g N_A_M1002_g 0.0321719f $X=6.115 $Y=0.74 $X2=0 $Y2=0
cc_317 B N_A_M1002_g 0.00394145f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_318 N_B_c_199_n N_A_M1002_g 0.019873f $X=6.175 $Y=1.41 $X2=0 $Y2=0
cc_319 B N_A_c_883_n 0.00268989f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_320 B N_A_M1018_g 0.00338754f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_321 N_B_M1026_g N_A_c_884_n 0.0295343f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_322 N_B_M1033_g N_A_c_885_n 0.0260938f $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_323 N_B_c_198_n A 0.00205068f $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_324 N_B_c_198_n N_A_c_887_n 0.0157952f $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_325 B N_A_1024_74#_M1013_d 0.00218982f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_326 N_B_M1031_g N_A_1024_74#_c_1053_n 0.0165938f $X=6.1 $Y=2.235 $X2=0 $Y2=0
cc_327 B N_A_1024_74#_c_1053_n 0.0201202f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_328 B N_A_1024_74#_c_1053_n 0.014429f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_329 N_B_M1039_g N_A_1024_74#_c_1056_n 0.00801378f $X=6.115 $Y=0.74 $X2=0
+ $Y2=0
cc_330 B N_A_1024_74#_c_1056_n 0.00823733f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_331 N_B_c_199_n N_A_1024_74#_c_1056_n 0.00329274f $X=6.175 $Y=1.41 $X2=0
+ $Y2=0
cc_332 B N_A_1024_74#_c_1059_n 0.0105533f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_333 B N_A_1024_74#_c_1040_n 0.00244385f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_334 B N_A_1024_74#_c_1048_n 0.00554056f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_335 N_B_M1031_g N_A_1024_74#_c_1050_n 0.00247959f $X=6.1 $Y=2.235 $X2=0 $Y2=0
cc_336 B N_A_1024_74#_c_1050_n 0.0190369f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_337 N_B_M1039_g N_A_1024_74#_c_1064_n 9.8919e-19 $X=6.115 $Y=0.74 $X2=0 $Y2=0
cc_338 N_B_M1039_g N_A_1024_74#_c_1065_n 0.00623463f $X=6.115 $Y=0.74 $X2=0
+ $Y2=0
cc_339 B N_A_1024_74#_c_1065_n 0.0290034f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_340 N_B_M1031_g N_A_1024_74#_c_1067_n 0.00312726f $X=6.1 $Y=2.235 $X2=0 $Y2=0
cc_341 B N_A_1024_74#_c_1067_n 0.0135032f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_342 N_B_c_199_n N_A_1024_74#_c_1067_n 3.81675e-19 $X=6.175 $Y=1.41 $X2=0
+ $Y2=0
cc_343 B N_A_1024_74#_c_1042_n 0.0140535f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_344 N_B_c_204_n N_A_27_392#_M1017_d 0.00657631f $X=1.75 $Y=1.95 $X2=0 $Y2=0
cc_345 N_B_c_216_p N_A_27_392#_M1017_d 0.00704391f $X=2.48 $Y=2.035 $X2=0 $Y2=0
cc_346 N_B_c_292_p N_A_27_392#_M1017_d 0.00509404f $X=1.835 $Y=2.035 $X2=0 $Y2=0
cc_347 N_B_M1017_g N_A_27_392#_c_1193_n 5.90871e-19 $X=1.155 $Y=2.235 $X2=0
+ $Y2=0
cc_348 N_B_M1017_g N_A_27_392#_c_1194_n 2.41803e-19 $X=1.155 $Y=2.235 $X2=0
+ $Y2=0
cc_349 N_B_M1017_g N_A_27_392#_c_1202_n 0.00691045f $X=1.155 $Y=2.235 $X2=0
+ $Y2=0
cc_350 N_B_M1017_g N_A_27_392#_c_1203_n 0.0144496f $X=1.155 $Y=2.235 $X2=0 $Y2=0
cc_351 N_B_M1017_g N_A_27_392#_c_1195_n 0.0045331f $X=1.155 $Y=2.235 $X2=0 $Y2=0
cc_352 N_B_M1017_g N_A_27_392#_c_1196_n 0.0122477f $X=1.155 $Y=2.235 $X2=0 $Y2=0
cc_353 N_B_c_222_p N_VPWR_M1005_d 0.00417829f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_354 N_B_c_209_n N_VPWR_M1012_d 0.00647789f $X=4.62 $Y=1.805 $X2=0 $Y2=0
cc_355 N_B_M1017_g N_VPWR_c_1242_n 0.00132436f $X=1.155 $Y=2.235 $X2=0 $Y2=0
cc_356 N_B_M1029_g N_VPWR_c_1243_n 0.00282337f $X=2.6 $Y=2.235 $X2=0 $Y2=0
cc_357 N_B_c_222_p N_VPWR_c_1243_n 0.0189268f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_358 N_B_c_316_p N_VPWR_c_1243_n 0.00111625f $X=2.645 $Y=1.83 $X2=0 $Y2=0
cc_359 N_B_M1012_g N_VPWR_c_1244_n 0.00408953f $X=4.06 $Y=2.235 $X2=0 $Y2=0
cc_360 N_B_M1029_g N_VPWR_c_1241_n 0.00112709f $X=2.6 $Y=2.235 $X2=0 $Y2=0
cc_361 N_B_M1012_g N_VPWR_c_1241_n 0.00112709f $X=4.06 $Y=2.235 $X2=0 $Y2=0
cc_362 N_B_M1031_g N_VPWR_c_1241_n 0.00112709f $X=6.1 $Y=2.235 $X2=0 $Y2=0
cc_363 N_B_c_222_p A_538_347# 0.00827664f $X=3.95 $Y=1.83 $X2=-0.19 $Y2=-0.245
cc_364 N_B_c_316_p A_538_347# 0.00279189f $X=2.645 $Y=1.83 $X2=-0.19 $Y2=-0.245
cc_365 N_B_c_222_p N_A_740_347#_M1006_d 0.00458324f $X=3.95 $Y=1.83 $X2=-0.19
+ $Y2=-0.245
cc_366 B N_A_740_347#_M1004_d 0.00232187f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_367 N_B_M1012_g N_A_740_347#_c_1390_n 0.0132612f $X=4.06 $Y=2.235 $X2=0 $Y2=0
cc_368 N_B_c_196_n N_A_740_347#_c_1390_n 3.72861e-19 $X=4.115 $Y=1.41 $X2=0
+ $Y2=0
cc_369 N_B_c_209_n N_A_740_347#_c_1390_n 0.0376356f $X=4.62 $Y=1.805 $X2=0 $Y2=0
cc_370 B N_A_740_347#_c_1390_n 0.00601209f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_371 B N_A_740_347#_c_1394_n 0.0171173f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_372 N_B_M1012_g N_A_740_347#_c_1387_n 0.00909377f $X=4.06 $Y=2.235 $X2=0
+ $Y2=0
cc_373 N_B_c_222_p N_A_740_347#_c_1387_n 0.014917f $X=3.95 $Y=1.83 $X2=0 $Y2=0
cc_374 N_B_c_209_n N_A_740_347#_c_1387_n 0.00248731f $X=4.62 $Y=1.805 $X2=0
+ $Y2=0
cc_375 B A_1144_347# 0.00145989f $X=5.915 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_376 B A_1144_347# 4.20571e-19 $X=6.395 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_377 B A_1238_347# 0.00209298f $X=6.395 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_378 N_B_M1030_g N_A_27_74#_c_1553_n 0.0150217f $X=1.585 $Y=0.74 $X2=0 $Y2=0
cc_379 N_B_c_198_n N_A_27_74#_c_1557_n 7.61274e-19 $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_380 N_B_M1026_g N_VGND_c_1585_n 0.00200275f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_381 N_B_M1030_g N_VGND_c_1589_n 0.00291649f $X=1.585 $Y=0.74 $X2=0 $Y2=0
cc_382 N_B_M1026_g N_VGND_c_1589_n 0.00461464f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_383 N_B_M1033_g N_VGND_c_1591_n 0.00220663f $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_384 N_B_M1033_g N_VGND_c_1592_n 0.00316493f $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_385 N_B_M1039_g N_VGND_c_1593_n 0.00278271f $X=6.115 $Y=0.74 $X2=0 $Y2=0
cc_386 N_B_M1030_g N_VGND_c_1599_n 0.00383588f $X=1.585 $Y=0.74 $X2=0 $Y2=0
cc_387 N_B_M1030_g N_VGND_c_1604_n 0.00364217f $X=1.585 $Y=0.74 $X2=0 $Y2=0
cc_388 N_B_M1026_g N_VGND_c_1604_n 0.0046687f $X=2.585 $Y=0.74 $X2=0 $Y2=0
cc_389 N_B_M1033_g N_VGND_c_1604_n 0.00393316f $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_390 N_B_M1039_g N_VGND_c_1604_n 0.00353931f $X=6.115 $Y=0.74 $X2=0 $Y2=0
cc_391 N_B_M1033_g N_A_734_74#_c_1734_n 0.00936301f $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_392 N_B_M1033_g N_A_734_74#_c_1732_n 0.00573013f $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_393 N_B_M1033_g N_A_734_74#_c_1733_n 8.6409e-19 $X=4.025 $Y=0.74 $X2=0 $Y2=0
cc_394 N_CIN_M1009_g N_A_418_74#_M1013_g 0.0241134f $X=5.63 $Y=2.235 $X2=0 $Y2=0
cc_395 N_CIN_M1027_g N_A_418_74#_c_614_n 0.00451566f $X=2.15 $Y=2.235 $X2=0
+ $Y2=0
cc_396 N_CIN_M1027_g N_A_418_74#_c_617_n 0.011867f $X=2.15 $Y=2.235 $X2=0 $Y2=0
cc_397 N_CIN_c_425_n N_A_418_74#_c_651_n 8.8084e-19 $X=2.305 $Y=1.295 $X2=0
+ $Y2=0
cc_398 N_CIN_c_431_n N_A_418_74#_c_651_n 0.0139672f $X=2.105 $Y=1.22 $X2=0 $Y2=0
cc_399 N_CIN_c_434_n N_A_418_74#_c_651_n 0.00689032f $X=2.16 $Y=1.295 $X2=0
+ $Y2=0
cc_400 N_CIN_c_431_n N_A_418_74#_c_591_n 0.00305832f $X=2.105 $Y=1.22 $X2=0
+ $Y2=0
cc_401 N_CIN_M1032_g N_A_418_74#_c_621_n 0.0102982f $X=3.595 $Y=0.74 $X2=0 $Y2=0
cc_402 N_CIN_c_423_n N_A_418_74#_c_621_n 0.00114091f $X=3.575 $Y=1.41 $X2=0
+ $Y2=0
cc_403 N_CIN_c_433_n N_A_418_74#_c_657_n 0.00343696f $X=5.635 $Y=1.22 $X2=0
+ $Y2=0
cc_404 N_CIN_c_433_n N_A_418_74#_c_592_n 0.0109994f $X=5.635 $Y=1.22 $X2=0 $Y2=0
cc_405 N_CIN_c_431_n N_A_418_74#_c_637_n 0.00235187f $X=2.105 $Y=1.22 $X2=0
+ $Y2=0
cc_406 N_CIN_c_424_n N_A_418_74#_c_660_n 0.00798157f $X=2.975 $Y=1.295 $X2=0
+ $Y2=0
cc_407 N_CIN_c_425_n N_A_418_74#_c_660_n 0.00288269f $X=2.305 $Y=1.295 $X2=0
+ $Y2=0
cc_408 N_CIN_c_430_n N_A_418_74#_c_660_n 9.09478e-19 $X=2.105 $Y=1.385 $X2=0
+ $Y2=0
cc_409 N_CIN_c_434_n N_A_418_74#_c_660_n 0.0098023f $X=2.16 $Y=1.295 $X2=0 $Y2=0
cc_410 N_CIN_M1027_g N_A_418_74#_c_606_n 0.0121124f $X=2.15 $Y=2.235 $X2=0 $Y2=0
cc_411 N_CIN_c_422_n N_A_418_74#_c_641_n 0.00659689f $X=3.575 $Y=1.41 $X2=0
+ $Y2=0
cc_412 N_CIN_c_424_n N_A_418_74#_c_641_n 0.0153931f $X=2.975 $Y=1.295 $X2=0
+ $Y2=0
cc_413 N_CIN_c_426_n N_A_418_74#_c_641_n 0.00299186f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_414 N_CIN_c_427_n N_A_418_74#_c_641_n 0.00799415f $X=3.265 $Y=1.295 $X2=0
+ $Y2=0
cc_415 N_CIN_c_435_n N_A_418_74#_c_641_n 0.0111957f $X=3.215 $Y=1.377 $X2=0
+ $Y2=0
cc_416 N_CIN_M1032_g N_A_418_74#_c_644_n 0.00631936f $X=3.595 $Y=0.74 $X2=0
+ $Y2=0
cc_417 N_CIN_c_422_n N_A_418_74#_c_644_n 0.0185241f $X=3.575 $Y=1.41 $X2=0 $Y2=0
cc_418 N_CIN_c_423_n N_A_418_74#_c_644_n 0.0018054f $X=3.575 $Y=1.41 $X2=0 $Y2=0
cc_419 N_CIN_c_426_n N_A_418_74#_c_644_n 0.0441427f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_420 N_CIN_c_426_n N_A_418_74#_c_596_n 0.0310488f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_421 N_CIN_c_428_n N_A_418_74#_c_596_n 0.0027738f $X=5.52 $Y=1.295 $X2=0 $Y2=0
cc_422 N_CIN_c_429_n N_A_418_74#_c_596_n 0.0267617f $X=5.52 $Y=1.295 $X2=0 $Y2=0
cc_423 N_CIN_c_432_n N_A_418_74#_c_596_n 4.59775e-19 $X=5.635 $Y=1.385 $X2=0
+ $Y2=0
cc_424 N_CIN_c_433_n N_A_418_74#_c_596_n 0.00293705f $X=5.635 $Y=1.22 $X2=0
+ $Y2=0
cc_425 N_CIN_c_426_n N_A_418_74#_c_597_n 0.0013891f $X=5.375 $Y=1.295 $X2=0
+ $Y2=0
cc_426 N_CIN_c_429_n N_A_418_74#_c_597_n 9.45146e-19 $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_427 N_CIN_c_432_n N_A_418_74#_c_597_n 0.0214172f $X=5.635 $Y=1.385 $X2=0
+ $Y2=0
cc_428 N_CIN_c_433_n N_A_418_74#_c_598_n 0.0134862f $X=5.635 $Y=1.22 $X2=0 $Y2=0
cc_429 N_CIN_M1027_g N_A_c_889_n 0.0120239f $X=2.15 $Y=2.235 $X2=0 $Y2=0
cc_430 N_CIN_c_423_n N_A_c_878_n 0.0213683f $X=3.575 $Y=1.41 $X2=0 $Y2=0
cc_431 N_CIN_c_435_n N_A_c_878_n 0.00270838f $X=3.215 $Y=1.377 $X2=0 $Y2=0
cc_432 N_CIN_M1006_g N_A_M1005_g 0.0224824f $X=3.61 $Y=2.235 $X2=0 $Y2=0
cc_433 N_CIN_c_435_n N_A_M1005_g 0.0107649f $X=3.215 $Y=1.377 $X2=0 $Y2=0
cc_434 N_CIN_M1006_g N_A_c_892_n 0.0123594f $X=3.61 $Y=2.235 $X2=0 $Y2=0
cc_435 N_CIN_c_426_n N_A_c_880_n 0.00251789f $X=5.375 $Y=1.295 $X2=0 $Y2=0
cc_436 N_CIN_c_426_n N_A_M1004_g 0.00369614f $X=5.375 $Y=1.295 $X2=0 $Y2=0
cc_437 N_CIN_M1009_g N_A_c_894_n 0.0123594f $X=5.63 $Y=2.235 $X2=0 $Y2=0
cc_438 N_CIN_M1032_g N_A_c_884_n 0.0241987f $X=3.595 $Y=0.74 $X2=0 $Y2=0
cc_439 N_CIN_c_427_n N_A_c_884_n 0.00140441f $X=3.265 $Y=1.295 $X2=0 $Y2=0
cc_440 N_CIN_c_435_n N_A_c_884_n 0.00117185f $X=3.215 $Y=1.377 $X2=0 $Y2=0
cc_441 N_CIN_M1009_g N_A_1024_74#_c_1053_n 0.0127807f $X=5.63 $Y=2.235 $X2=0
+ $Y2=0
cc_442 N_CIN_M1009_g N_A_1024_74#_c_1050_n 0.0122495f $X=5.63 $Y=2.235 $X2=0
+ $Y2=0
cc_443 N_CIN_c_428_n N_A_1024_74#_c_1064_n 0.00673868f $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_444 N_CIN_c_429_n N_A_1024_74#_c_1064_n 0.0151874f $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_445 N_CIN_c_432_n N_A_1024_74#_c_1064_n 0.00107034f $X=5.635 $Y=1.385 $X2=0
+ $Y2=0
cc_446 N_CIN_c_433_n N_A_1024_74#_c_1064_n 0.00623624f $X=5.635 $Y=1.22 $X2=0
+ $Y2=0
cc_447 N_CIN_c_429_n N_A_1024_74#_c_1077_n 0.00504528f $X=5.52 $Y=1.295 $X2=0
+ $Y2=0
cc_448 N_CIN_c_433_n N_A_1024_74#_c_1077_n 0.0102416f $X=5.635 $Y=1.22 $X2=0
+ $Y2=0
cc_449 N_CIN_c_433_n N_A_1024_74#_c_1065_n 0.00111404f $X=5.635 $Y=1.22 $X2=0
+ $Y2=0
cc_450 N_CIN_M1027_g N_A_27_392#_c_1196_n 0.00778168f $X=2.15 $Y=2.235 $X2=0
+ $Y2=0
cc_451 N_CIN_M1006_g N_VPWR_c_1243_n 0.00212303f $X=3.61 $Y=2.235 $X2=0 $Y2=0
cc_452 N_CIN_M1027_g N_VPWR_c_1241_n 0.00112709f $X=2.15 $Y=2.235 $X2=0 $Y2=0
cc_453 N_CIN_M1006_g N_VPWR_c_1241_n 0.00112709f $X=3.61 $Y=2.235 $X2=0 $Y2=0
cc_454 N_CIN_M1009_g N_VPWR_c_1241_n 0.00112709f $X=5.63 $Y=2.235 $X2=0 $Y2=0
cc_455 N_CIN_M1006_g N_A_740_347#_c_1387_n 0.00889371f $X=3.61 $Y=2.235 $X2=0
+ $Y2=0
cc_456 N_CIN_c_431_n N_A_27_74#_c_1553_n 0.00409096f $X=2.105 $Y=1.22 $X2=0
+ $Y2=0
cc_457 N_CIN_M1032_g N_VGND_c_1585_n 0.00193337f $X=3.595 $Y=0.74 $X2=0 $Y2=0
cc_458 N_CIN_c_431_n N_VGND_c_1589_n 0.00433162f $X=2.105 $Y=1.22 $X2=0 $Y2=0
cc_459 N_CIN_M1032_g N_VGND_c_1592_n 0.00461464f $X=3.595 $Y=0.74 $X2=0 $Y2=0
cc_460 N_CIN_c_433_n N_VGND_c_1593_n 0.00278271f $X=5.635 $Y=1.22 $X2=0 $Y2=0
cc_461 N_CIN_M1032_g N_VGND_c_1604_n 0.00804222f $X=3.595 $Y=0.74 $X2=0 $Y2=0
cc_462 N_CIN_c_431_n N_VGND_c_1604_n 0.0044836f $X=2.105 $Y=1.22 $X2=0 $Y2=0
cc_463 N_CIN_c_433_n N_VGND_c_1604_n 0.00354203f $X=5.635 $Y=1.22 $X2=0 $Y2=0
cc_464 N_A_418_74#_c_630_n N_A_M1003_g 0.00288058f $X=1.41 $Y=1.83 $X2=0 $Y2=0
cc_465 N_A_418_74#_c_590_n N_A_M1034_g 0.00398634f $X=1.09 $Y=1.745 $X2=0 $Y2=0
cc_466 N_A_418_74#_c_685_p N_A_M1034_g 0.00328708f $X=1.175 $Y=1.005 $X2=0 $Y2=0
cc_467 N_A_418_74#_c_617_n N_A_c_889_n 0.00154558f $X=2.21 $Y=2.375 $X2=0 $Y2=0
cc_468 N_A_418_74#_c_606_n N_A_c_889_n 0.00549911f $X=2.375 $Y=2.375 $X2=0 $Y2=0
cc_469 N_A_418_74#_c_606_n N_A_M1005_g 0.00141635f $X=2.375 $Y=2.375 $X2=0 $Y2=0
cc_470 N_A_418_74#_c_596_n N_A_c_880_n 0.00253264f $X=5.095 $Y=1.005 $X2=0 $Y2=0
cc_471 N_A_418_74#_c_597_n N_A_c_880_n 0.0208244f $X=5.095 $Y=1.385 $X2=0 $Y2=0
cc_472 N_A_418_74#_c_598_n N_A_c_880_n 0.00165443f $X=5.095 $Y=1.22 $X2=0 $Y2=0
cc_473 N_A_418_74#_M1013_g N_A_M1004_g 0.0243146f $X=5.13 $Y=2.235 $X2=0 $Y2=0
cc_474 N_A_418_74#_M1013_g N_A_c_894_n 0.0123594f $X=5.13 $Y=2.235 $X2=0 $Y2=0
cc_475 N_A_418_74#_c_592_n N_A_M1002_g 0.00209511f $X=6.255 $Y=0.34 $X2=0 $Y2=0
cc_476 N_A_418_74#_c_628_n N_A_M1002_g 0.00349056f $X=6.34 $Y=0.58 $X2=0 $Y2=0
cc_477 N_A_418_74#_c_696_p N_A_M1002_g 0.012131f $X=8.965 $Y=0.665 $X2=0 $Y2=0
cc_478 N_A_418_74#_c_641_n N_A_c_884_n 0.0122961f $X=3.385 $Y=0.965 $X2=0 $Y2=0
cc_479 N_A_418_74#_c_644_n N_A_c_884_n 0.00216961f $X=3.555 $Y=0.965 $X2=0 $Y2=0
cc_480 N_A_418_74#_c_621_n N_A_c_885_n 0.0127763f $X=4.93 $Y=1.005 $X2=0 $Y2=0
cc_481 N_A_418_74#_c_657_n N_A_c_885_n 9.47922e-19 $X=5.17 $Y=0.92 $X2=0 $Y2=0
cc_482 N_A_418_74#_c_593_n N_A_c_885_n 3.23044e-19 $X=5.255 $Y=0.34 $X2=0 $Y2=0
cc_483 N_A_418_74#_c_596_n N_A_c_885_n 0.00165995f $X=5.095 $Y=1.005 $X2=0 $Y2=0
cc_484 N_A_418_74#_c_598_n N_A_c_885_n 0.0249033f $X=5.095 $Y=1.22 $X2=0 $Y2=0
cc_485 N_A_418_74#_c_590_n A 0.0422556f $X=1.09 $Y=1.745 $X2=0 $Y2=0
cc_486 N_A_418_74#_c_630_n A 0.00291428f $X=1.41 $Y=1.83 $X2=0 $Y2=0
cc_487 N_A_418_74#_c_590_n N_A_c_887_n 9.1952e-19 $X=1.09 $Y=1.745 $X2=0 $Y2=0
cc_488 N_A_418_74#_c_657_n N_A_1024_74#_M1016_d 0.00532706f $X=5.17 $Y=0.92
+ $X2=-0.19 $Y2=-0.245
cc_489 N_A_418_74#_c_592_n N_A_1024_74#_M1016_d 0.0087698f $X=6.255 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_490 N_A_418_74#_c_596_n N_A_1024_74#_M1016_d 0.00250765f $X=5.095 $Y=1.005
+ $X2=-0.19 $Y2=-0.245
cc_491 N_A_418_74#_c_696_p N_A_1024_74#_M1022_g 0.0136954f $X=8.965 $Y=0.665
+ $X2=0 $Y2=0
cc_492 N_A_418_74#_c_696_p N_A_1024_74#_M1024_g 0.0120977f $X=8.965 $Y=0.665
+ $X2=0 $Y2=0
cc_493 N_A_418_74#_c_696_p N_A_1024_74#_M1036_g 0.0120967f $X=8.965 $Y=0.665
+ $X2=0 $Y2=0
cc_494 N_A_418_74#_M1000_g N_A_1024_74#_M1020_g 0.00966283f $X=9.085 $Y=2.4
+ $X2=0 $Y2=0
cc_495 N_A_418_74#_M1011_g N_A_1024_74#_M1038_g 0.021129f $X=9.255 $Y=0.78 $X2=0
+ $Y2=0
cc_496 N_A_418_74#_c_696_p N_A_1024_74#_M1038_g 0.0156149f $X=8.965 $Y=0.665
+ $X2=0 $Y2=0
cc_497 N_A_418_74#_c_594_n N_A_1024_74#_M1038_g 0.00692925f $X=9.05 $Y=1.32
+ $X2=0 $Y2=0
cc_498 N_A_418_74#_c_595_n N_A_1024_74#_M1038_g 0.0017339f $X=9.135 $Y=1.485
+ $X2=0 $Y2=0
cc_499 N_A_418_74#_c_599_n N_A_1024_74#_M1038_g 0.00877228f $X=10.485 $Y=1.485
+ $X2=0 $Y2=0
cc_500 N_A_418_74#_c_592_n N_A_1024_74#_c_1056_n 0.00321187f $X=6.255 $Y=0.34
+ $X2=0 $Y2=0
cc_501 N_A_418_74#_c_696_p N_A_1024_74#_c_1056_n 0.0396142f $X=8.965 $Y=0.665
+ $X2=0 $Y2=0
cc_502 N_A_418_74#_c_629_n N_A_1024_74#_c_1056_n 0.0134799f $X=6.425 $Y=0.665
+ $X2=0 $Y2=0
cc_503 N_A_418_74#_c_696_p N_A_1024_74#_c_1041_n 0.00424675f $X=8.965 $Y=0.665
+ $X2=0 $Y2=0
cc_504 N_A_418_74#_M1013_g N_A_1024_74#_c_1050_n 4.63834e-19 $X=5.13 $Y=2.235
+ $X2=0 $Y2=0
cc_505 N_A_418_74#_c_657_n N_A_1024_74#_c_1064_n 0.0242712f $X=5.17 $Y=0.92
+ $X2=0 $Y2=0
cc_506 N_A_418_74#_c_592_n N_A_1024_74#_c_1064_n 0.0138888f $X=6.255 $Y=0.34
+ $X2=0 $Y2=0
cc_507 N_A_418_74#_c_629_n N_A_1024_74#_c_1064_n 0.0047823f $X=6.425 $Y=0.665
+ $X2=0 $Y2=0
cc_508 N_A_418_74#_c_596_n N_A_1024_74#_c_1064_n 0.00751744f $X=5.095 $Y=1.005
+ $X2=0 $Y2=0
cc_509 N_A_418_74#_c_598_n N_A_1024_74#_c_1064_n 0.0012068f $X=5.095 $Y=1.22
+ $X2=0 $Y2=0
cc_510 N_A_418_74#_c_592_n N_A_1024_74#_c_1077_n 0.00892235f $X=6.255 $Y=0.34
+ $X2=0 $Y2=0
cc_511 N_A_418_74#_c_596_n N_A_1024_74#_c_1065_n 0.00253405f $X=5.095 $Y=1.005
+ $X2=0 $Y2=0
cc_512 N_A_418_74#_c_696_p N_A_1024_74#_c_1043_n 2.94247e-19 $X=8.965 $Y=0.665
+ $X2=0 $Y2=0
cc_513 N_A_418_74#_c_595_n N_A_1024_74#_c_1043_n 0.00159647f $X=9.135 $Y=1.485
+ $X2=0 $Y2=0
cc_514 N_A_418_74#_c_599_n N_A_1024_74#_c_1043_n 0.00966283f $X=10.485 $Y=1.485
+ $X2=0 $Y2=0
cc_515 N_A_418_74#_c_614_n N_A_27_392#_M1017_d 0.0110843f $X=1.41 $Y=2.29 $X2=0
+ $Y2=0
cc_516 N_A_418_74#_c_617_n N_A_27_392#_M1017_d 0.0185537f $X=2.21 $Y=2.375 $X2=0
+ $Y2=0
cc_517 N_A_418_74#_c_619_n N_A_27_392#_M1017_d 0.00460616f $X=1.495 $Y=2.375
+ $X2=0 $Y2=0
cc_518 N_A_418_74#_c_630_n N_A_27_392#_M1017_d 0.00555537f $X=1.41 $Y=1.83 $X2=0
+ $Y2=0
cc_519 N_A_418_74#_c_614_n N_A_27_392#_c_1202_n 0.0133617f $X=1.41 $Y=2.29 $X2=0
+ $Y2=0
cc_520 N_A_418_74#_c_630_n N_A_27_392#_c_1202_n 0.00690066f $X=1.41 $Y=1.83
+ $X2=0 $Y2=0
cc_521 N_A_418_74#_c_614_n N_A_27_392#_c_1203_n 0.00238694f $X=1.41 $Y=2.29
+ $X2=0 $Y2=0
cc_522 N_A_418_74#_c_619_n N_A_27_392#_c_1203_n 0.0134181f $X=1.495 $Y=2.375
+ $X2=0 $Y2=0
cc_523 N_A_418_74#_c_617_n N_A_27_392#_c_1196_n 0.038786f $X=2.21 $Y=2.375 $X2=0
+ $Y2=0
cc_524 N_A_418_74#_c_619_n N_A_27_392#_c_1196_n 0.0142344f $X=1.495 $Y=2.375
+ $X2=0 $Y2=0
cc_525 N_A_418_74#_c_606_n N_A_27_392#_c_1196_n 0.00479707f $X=2.375 $Y=2.375
+ $X2=0 $Y2=0
cc_526 N_A_418_74#_c_630_n N_VPWR_M1003_d 0.00249008f $X=1.41 $Y=1.83 $X2=-0.19
+ $Y2=-0.245
cc_527 N_A_418_74#_c_606_n N_VPWR_c_1243_n 0.011746f $X=2.375 $Y=2.375 $X2=0
+ $Y2=0
cc_528 N_A_418_74#_M1013_g N_VPWR_c_1244_n 6.00163e-19 $X=5.13 $Y=2.235 $X2=0
+ $Y2=0
cc_529 N_A_418_74#_M1000_g N_VPWR_c_1247_n 0.00361832f $X=9.085 $Y=2.4 $X2=0
+ $Y2=0
cc_530 N_A_418_74#_c_595_n N_VPWR_c_1247_n 8.43278e-19 $X=9.135 $Y=1.485 $X2=0
+ $Y2=0
cc_531 N_A_418_74#_M1019_g N_VPWR_c_1248_n 0.00356597f $X=9.535 $Y=2.4 $X2=0
+ $Y2=0
cc_532 N_A_418_74#_M1021_g N_VPWR_c_1248_n 0.00371548f $X=10.035 $Y=2.4 $X2=0
+ $Y2=0
cc_533 N_A_418_74#_M1023_g N_VPWR_c_1250_n 0.0064857f $X=10.485 $Y=2.4 $X2=0
+ $Y2=0
cc_534 N_A_418_74#_c_606_n N_VPWR_c_1251_n 0.00721197f $X=2.375 $Y=2.375 $X2=0
+ $Y2=0
cc_535 N_A_418_74#_M1000_g N_VPWR_c_1257_n 0.005209f $X=9.085 $Y=2.4 $X2=0 $Y2=0
cc_536 N_A_418_74#_M1019_g N_VPWR_c_1257_n 0.005209f $X=9.535 $Y=2.4 $X2=0 $Y2=0
cc_537 N_A_418_74#_M1021_g N_VPWR_c_1258_n 0.005209f $X=10.035 $Y=2.4 $X2=0
+ $Y2=0
cc_538 N_A_418_74#_M1023_g N_VPWR_c_1258_n 0.0050957f $X=10.485 $Y=2.4 $X2=0
+ $Y2=0
cc_539 N_A_418_74#_M1013_g N_VPWR_c_1241_n 0.00112709f $X=5.13 $Y=2.235 $X2=0
+ $Y2=0
cc_540 N_A_418_74#_M1000_g N_VPWR_c_1241_n 0.0098216f $X=9.085 $Y=2.4 $X2=0
+ $Y2=0
cc_541 N_A_418_74#_M1019_g N_VPWR_c_1241_n 0.00982754f $X=9.535 $Y=2.4 $X2=0
+ $Y2=0
cc_542 N_A_418_74#_M1021_g N_VPWR_c_1241_n 0.00982082f $X=10.035 $Y=2.4 $X2=0
+ $Y2=0
cc_543 N_A_418_74#_M1023_g N_VPWR_c_1241_n 0.00949482f $X=10.485 $Y=2.4 $X2=0
+ $Y2=0
cc_544 N_A_418_74#_c_606_n N_VPWR_c_1241_n 0.00886293f $X=2.375 $Y=2.375 $X2=0
+ $Y2=0
cc_545 N_A_418_74#_M1013_g N_A_740_347#_c_1394_n 0.00235607f $X=5.13 $Y=2.235
+ $X2=0 $Y2=0
cc_546 N_A_418_74#_M1013_g N_A_740_347#_c_1386_n 0.00656212f $X=5.13 $Y=2.235
+ $X2=0 $Y2=0
cc_547 N_A_418_74#_c_696_p N_SUM_M1022_s 0.00437807f $X=8.965 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_548 N_A_418_74#_c_696_p N_SUM_M1036_s 0.00437412f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_549 N_A_418_74#_c_696_p N_SUM_c_1423_n 0.0576451f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_550 N_A_418_74#_c_696_p N_SUM_c_1424_n 0.0170377f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_551 N_A_418_74#_c_594_n N_SUM_c_1424_n 0.011264f $X=9.05 $Y=1.32 $X2=0 $Y2=0
cc_552 N_A_418_74#_M1000_g N_SUM_c_1425_n 7.98897e-19 $X=9.085 $Y=2.4 $X2=0
+ $Y2=0
cc_553 N_A_418_74#_c_594_n N_SUM_c_1425_n 0.00593841f $X=9.05 $Y=1.32 $X2=0
+ $Y2=0
cc_554 N_A_418_74#_c_595_n N_SUM_c_1425_n 0.0134827f $X=9.135 $Y=1.485 $X2=0
+ $Y2=0
cc_555 N_A_418_74#_c_599_n N_SUM_c_1425_n 2.94226e-19 $X=10.485 $Y=1.485 $X2=0
+ $Y2=0
cc_556 N_A_418_74#_M1000_g N_COUT_c_1488_n 0.00258023f $X=9.085 $Y=2.4 $X2=0
+ $Y2=0
cc_557 N_A_418_74#_M1019_g N_COUT_c_1488_n 0.00112087f $X=9.535 $Y=2.4 $X2=0
+ $Y2=0
cc_558 N_A_418_74#_c_777_p N_COUT_c_1488_n 0.0275631f $X=9.84 $Y=1.485 $X2=0
+ $Y2=0
cc_559 N_A_418_74#_c_599_n N_COUT_c_1488_n 0.00245159f $X=10.485 $Y=1.485 $X2=0
+ $Y2=0
cc_560 N_A_418_74#_M1000_g N_COUT_c_1489_n 0.0122358f $X=9.085 $Y=2.4 $X2=0
+ $Y2=0
cc_561 N_A_418_74#_M1019_g N_COUT_c_1489_n 0.014321f $X=9.535 $Y=2.4 $X2=0 $Y2=0
cc_562 N_A_418_74#_M1021_g N_COUT_c_1489_n 6.73979e-19 $X=10.035 $Y=2.4 $X2=0
+ $Y2=0
cc_563 N_A_418_74#_M1011_g N_COUT_c_1484_n 0.00852713f $X=9.255 $Y=0.78 $X2=0
+ $Y2=0
cc_564 N_A_418_74#_M1014_g N_COUT_c_1484_n 3.13308e-19 $X=9.685 $Y=0.78 $X2=0
+ $Y2=0
cc_565 N_A_418_74#_M1019_g N_COUT_c_1490_n 0.0132272f $X=9.535 $Y=2.4 $X2=0
+ $Y2=0
cc_566 N_A_418_74#_M1021_g N_COUT_c_1490_n 0.0152762f $X=10.035 $Y=2.4 $X2=0
+ $Y2=0
cc_567 N_A_418_74#_c_777_p N_COUT_c_1490_n 0.0354452f $X=9.84 $Y=1.485 $X2=0
+ $Y2=0
cc_568 N_A_418_74#_c_599_n N_COUT_c_1490_n 0.00367077f $X=10.485 $Y=1.485 $X2=0
+ $Y2=0
cc_569 N_A_418_74#_M1014_g N_COUT_c_1506_n 0.0122129f $X=9.685 $Y=0.78 $X2=0
+ $Y2=0
cc_570 N_A_418_74#_M1025_g N_COUT_c_1506_n 0.0129763f $X=10.115 $Y=0.78 $X2=0
+ $Y2=0
cc_571 N_A_418_74#_c_777_p N_COUT_c_1506_n 0.0250701f $X=9.84 $Y=1.485 $X2=0
+ $Y2=0
cc_572 N_A_418_74#_c_599_n N_COUT_c_1506_n 0.00261635f $X=10.485 $Y=1.485 $X2=0
+ $Y2=0
cc_573 N_A_418_74#_M1011_g N_COUT_c_1485_n 0.00211285f $X=9.255 $Y=0.78 $X2=0
+ $Y2=0
cc_574 N_A_418_74#_c_777_p N_COUT_c_1485_n 0.0178863f $X=9.84 $Y=1.485 $X2=0
+ $Y2=0
cc_575 N_A_418_74#_c_599_n N_COUT_c_1485_n 0.00272398f $X=10.485 $Y=1.485 $X2=0
+ $Y2=0
cc_576 N_A_418_74#_M1014_g N_COUT_c_1486_n 6.05373e-19 $X=9.685 $Y=0.78 $X2=0
+ $Y2=0
cc_577 N_A_418_74#_M1025_g N_COUT_c_1486_n 0.00849808f $X=10.115 $Y=0.78 $X2=0
+ $Y2=0
cc_578 N_A_418_74#_M1037_g N_COUT_c_1486_n 4.03226e-19 $X=10.545 $Y=0.78 $X2=0
+ $Y2=0
cc_579 N_A_418_74#_M1014_g N_COUT_c_1487_n 8.24123e-19 $X=9.685 $Y=0.78 $X2=0
+ $Y2=0
cc_580 N_A_418_74#_M1025_g N_COUT_c_1487_n 0.00456448f $X=10.115 $Y=0.78 $X2=0
+ $Y2=0
cc_581 N_A_418_74#_M1037_g N_COUT_c_1487_n 0.00407331f $X=10.545 $Y=0.78 $X2=0
+ $Y2=0
cc_582 N_A_418_74#_c_777_p N_COUT_c_1487_n 0.0151308f $X=9.84 $Y=1.485 $X2=0
+ $Y2=0
cc_583 N_A_418_74#_c_599_n N_COUT_c_1487_n 0.0209301f $X=10.485 $Y=1.485 $X2=0
+ $Y2=0
cc_584 N_A_418_74#_M1025_g N_COUT_c_1521_n 3.84191e-19 $X=10.115 $Y=0.78 $X2=0
+ $Y2=0
cc_585 N_A_418_74#_M1021_g N_COUT_c_1491_n 0.00607039f $X=10.035 $Y=2.4 $X2=0
+ $Y2=0
cc_586 N_A_418_74#_M1023_g N_COUT_c_1491_n 0.0114116f $X=10.485 $Y=2.4 $X2=0
+ $Y2=0
cc_587 N_A_418_74#_c_777_p N_COUT_c_1491_n 0.0066008f $X=9.84 $Y=1.485 $X2=0
+ $Y2=0
cc_588 N_A_418_74#_c_599_n N_COUT_c_1491_n 0.0108916f $X=10.485 $Y=1.485 $X2=0
+ $Y2=0
cc_589 N_A_418_74#_M1019_g COUT 6.41635e-19 $X=9.535 $Y=2.4 $X2=0 $Y2=0
cc_590 N_A_418_74#_M1021_g COUT 0.0137444f $X=10.035 $Y=2.4 $X2=0 $Y2=0
cc_591 N_A_418_74#_M1023_g COUT 0.0140068f $X=10.485 $Y=2.4 $X2=0 $Y2=0
cc_592 N_A_418_74#_c_651_n N_A_27_74#_M1030_d 0.00228734f $X=2.135 $Y=0.925
+ $X2=0 $Y2=0
cc_593 N_A_418_74#_c_637_n N_A_27_74#_M1030_d 0.00356839f $X=1.835 $Y=0.965
+ $X2=0 $Y2=0
cc_594 N_A_418_74#_c_591_n N_A_27_74#_c_1553_n 0.0140589f $X=2.3 $Y=0.515 $X2=0
+ $Y2=0
cc_595 N_A_418_74#_c_634_n N_A_27_74#_c_1553_n 0.00782456f $X=1.665 $Y=0.965
+ $X2=0 $Y2=0
cc_596 N_A_418_74#_c_637_n N_A_27_74#_c_1553_n 0.0142648f $X=1.835 $Y=0.965
+ $X2=0 $Y2=0
cc_597 N_A_418_74#_c_685_p N_A_27_74#_c_1554_n 0.00503853f $X=1.175 $Y=1.005
+ $X2=0 $Y2=0
cc_598 N_A_418_74#_c_685_p N_A_27_74#_c_1557_n 0.013831f $X=1.175 $Y=1.005 $X2=0
+ $Y2=0
cc_599 N_A_418_74#_c_634_n N_A_27_74#_c_1557_n 0.0207538f $X=1.665 $Y=0.965
+ $X2=0 $Y2=0
cc_600 N_A_418_74#_c_590_n N_VGND_M1034_d 5.28288e-19 $X=1.09 $Y=1.745 $X2=-0.19
+ $Y2=-0.245
cc_601 N_A_418_74#_c_685_p N_VGND_M1034_d 0.00604059f $X=1.175 $Y=1.005
+ $X2=-0.19 $Y2=-0.245
cc_602 N_A_418_74#_c_634_n N_VGND_M1034_d 0.00740987f $X=1.665 $Y=0.965
+ $X2=-0.19 $Y2=-0.245
cc_603 N_A_418_74#_c_641_n N_VGND_M1035_d 0.00278732f $X=3.385 $Y=0.965 $X2=0
+ $Y2=0
cc_604 N_A_418_74#_c_644_n N_VGND_M1035_d 0.00256535f $X=3.555 $Y=0.965 $X2=0
+ $Y2=0
cc_605 N_A_418_74#_c_621_n N_VGND_M1033_d 0.00849548f $X=4.93 $Y=1.005 $X2=0
+ $Y2=0
cc_606 N_A_418_74#_c_696_p N_VGND_M1002_d 0.007557f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_607 N_A_418_74#_c_696_p N_VGND_M1024_d 0.00726636f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_608 N_A_418_74#_c_696_p N_VGND_M1038_d 0.0116153f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_609 N_A_418_74#_c_594_n N_VGND_M1038_d 0.00806651f $X=9.05 $Y=1.32 $X2=0
+ $Y2=0
cc_610 N_A_418_74#_c_641_n N_VGND_c_1585_n 0.0176682f $X=3.385 $Y=0.965 $X2=0
+ $Y2=0
cc_611 N_A_418_74#_M1011_g N_VGND_c_1586_n 4.88565e-19 $X=9.255 $Y=0.78 $X2=0
+ $Y2=0
cc_612 N_A_418_74#_M1014_g N_VGND_c_1586_n 0.00879111f $X=9.685 $Y=0.78 $X2=0
+ $Y2=0
cc_613 N_A_418_74#_M1025_g N_VGND_c_1586_n 0.00176539f $X=10.115 $Y=0.78 $X2=0
+ $Y2=0
cc_614 N_A_418_74#_M1025_g N_VGND_c_1588_n 5.99782e-19 $X=10.115 $Y=0.78 $X2=0
+ $Y2=0
cc_615 N_A_418_74#_M1037_g N_VGND_c_1588_n 0.0157698f $X=10.545 $Y=0.78 $X2=0
+ $Y2=0
cc_616 N_A_418_74#_c_591_n N_VGND_c_1589_n 0.0146038f $X=2.3 $Y=0.515 $X2=0
+ $Y2=0
cc_617 N_A_418_74#_c_593_n N_VGND_c_1591_n 0.00302543f $X=5.255 $Y=0.34 $X2=0
+ $Y2=0
cc_618 N_A_418_74#_c_592_n N_VGND_c_1593_n 0.0753865f $X=6.255 $Y=0.34 $X2=0
+ $Y2=0
cc_619 N_A_418_74#_c_593_n N_VGND_c_1593_n 0.0120637f $X=5.255 $Y=0.34 $X2=0
+ $Y2=0
cc_620 N_A_418_74#_c_696_p N_VGND_c_1593_n 0.00540182f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_621 N_A_418_74#_c_598_n N_VGND_c_1593_n 0.00418685f $X=5.095 $Y=1.22 $X2=0
+ $Y2=0
cc_622 N_A_418_74#_c_696_p N_VGND_c_1594_n 0.0114147f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_623 N_A_418_74#_c_696_p N_VGND_c_1595_n 0.0114147f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_624 N_A_418_74#_M1011_g N_VGND_c_1596_n 0.00523933f $X=9.255 $Y=0.78 $X2=0
+ $Y2=0
cc_625 N_A_418_74#_M1014_g N_VGND_c_1596_n 0.00455951f $X=9.685 $Y=0.78 $X2=0
+ $Y2=0
cc_626 N_A_418_74#_M1025_g N_VGND_c_1597_n 0.00523933f $X=10.115 $Y=0.78 $X2=0
+ $Y2=0
cc_627 N_A_418_74#_M1037_g N_VGND_c_1597_n 0.00455951f $X=10.545 $Y=0.78 $X2=0
+ $Y2=0
cc_628 N_A_418_74#_c_592_n N_VGND_c_1600_n 0.00746752f $X=6.255 $Y=0.34 $X2=0
+ $Y2=0
cc_629 N_A_418_74#_c_696_p N_VGND_c_1600_n 0.0244407f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_630 N_A_418_74#_c_696_p N_VGND_c_1601_n 0.0244835f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_631 N_A_418_74#_M1011_g N_VGND_c_1602_n 0.00192643f $X=9.255 $Y=0.78 $X2=0
+ $Y2=0
cc_632 N_A_418_74#_c_696_p N_VGND_c_1602_n 0.0256831f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_633 N_A_418_74#_M1011_g N_VGND_c_1604_n 0.00533081f $X=9.255 $Y=0.78 $X2=0
+ $Y2=0
cc_634 N_A_418_74#_M1014_g N_VGND_c_1604_n 0.00447788f $X=9.685 $Y=0.78 $X2=0
+ $Y2=0
cc_635 N_A_418_74#_M1025_g N_VGND_c_1604_n 0.00533081f $X=10.115 $Y=0.78 $X2=0
+ $Y2=0
cc_636 N_A_418_74#_M1037_g N_VGND_c_1604_n 0.00447788f $X=10.545 $Y=0.78 $X2=0
+ $Y2=0
cc_637 N_A_418_74#_c_591_n N_VGND_c_1604_n 0.0121018f $X=2.3 $Y=0.515 $X2=0
+ $Y2=0
cc_638 N_A_418_74#_c_592_n N_VGND_c_1604_n 0.04278f $X=6.255 $Y=0.34 $X2=0 $Y2=0
cc_639 N_A_418_74#_c_593_n N_VGND_c_1604_n 0.00644906f $X=5.255 $Y=0.34 $X2=0
+ $Y2=0
cc_640 N_A_418_74#_c_696_p N_VGND_c_1604_n 0.0551926f $X=8.965 $Y=0.665 $X2=0
+ $Y2=0
cc_641 N_A_418_74#_c_637_n N_VGND_c_1604_n 0.00539663f $X=1.835 $Y=0.965 $X2=0
+ $Y2=0
cc_642 N_A_418_74#_c_641_n N_VGND_c_1604_n 0.0236322f $X=3.385 $Y=0.965 $X2=0
+ $Y2=0
cc_643 N_A_418_74#_c_644_n N_VGND_c_1604_n 0.00156853f $X=3.555 $Y=0.965 $X2=0
+ $Y2=0
cc_644 N_A_418_74#_c_598_n N_VGND_c_1604_n 0.0078168f $X=5.095 $Y=1.22 $X2=0
+ $Y2=0
cc_645 N_A_418_74#_c_641_n A_532_74# 0.00912043f $X=3.385 $Y=0.965 $X2=-0.19
+ $Y2=-0.245
cc_646 N_A_418_74#_c_621_n N_A_734_74#_M1032_d 0.00443657f $X=4.93 $Y=1.005
+ $X2=-0.19 $Y2=-0.245
cc_647 N_A_418_74#_c_621_n N_A_734_74#_M1015_d 0.00451688f $X=4.93 $Y=1.005
+ $X2=0 $Y2=0
cc_648 N_A_418_74#_c_621_n N_A_734_74#_c_1734_n 0.0390509f $X=4.93 $Y=1.005
+ $X2=0 $Y2=0
cc_649 N_A_418_74#_c_621_n N_A_734_74#_c_1732_n 0.0140929f $X=4.93 $Y=1.005
+ $X2=0 $Y2=0
cc_650 N_A_418_74#_c_621_n N_A_734_74#_c_1733_n 0.0140929f $X=4.93 $Y=1.005
+ $X2=0 $Y2=0
cc_651 N_A_418_74#_c_593_n N_A_734_74#_c_1733_n 0.00392045f $X=5.255 $Y=0.34
+ $X2=0 $Y2=0
cc_652 N_A_418_74#_c_592_n A_1160_74# 0.00206111f $X=6.255 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_653 N_A_418_74#_c_592_n A_1238_74# 8.72382e-19 $X=6.255 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_654 N_A_418_74#_c_628_n A_1238_74# 0.00341292f $X=6.34 $Y=0.58 $X2=-0.19
+ $Y2=-0.245
cc_655 N_A_418_74#_c_696_p A_1238_74# 0.00180488f $X=8.965 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_656 N_A_418_74#_c_629_n A_1238_74# 0.0049852f $X=6.425 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_657 N_A_M1018_g N_A_1024_74#_M1007_g 0.0148403f $X=6.64 $Y=2.34 $X2=0 $Y2=0
cc_658 N_A_M1002_g N_A_1024_74#_M1022_g 0.025914f $X=6.625 $Y=0.74 $X2=0 $Y2=0
cc_659 N_A_M1002_g N_A_1024_74#_c_1056_n 0.0149876f $X=6.625 $Y=0.74 $X2=0 $Y2=0
cc_660 N_A_M1018_g N_A_1024_74#_c_1059_n 0.0208776f $X=6.64 $Y=2.34 $X2=0 $Y2=0
cc_661 N_A_M1002_g N_A_1024_74#_c_1040_n 0.00444019f $X=6.625 $Y=0.74 $X2=0
+ $Y2=0
cc_662 N_A_c_883_n N_A_1024_74#_c_1048_n 0.00453536f $X=6.64 $Y=1.705 $X2=0
+ $Y2=0
cc_663 N_A_c_894_n N_A_1024_74#_c_1050_n 0.00614211f $X=6.55 $Y=3.15 $X2=0 $Y2=0
cc_664 N_A_M1002_g N_A_1024_74#_c_1065_n 3.84346e-19 $X=6.625 $Y=0.74 $X2=0
+ $Y2=0
cc_665 N_A_M1018_g N_A_1024_74#_c_1067_n 0.00280267f $X=6.64 $Y=2.34 $X2=0 $Y2=0
cc_666 N_A_M1002_g N_A_1024_74#_c_1042_n 0.0031874f $X=6.625 $Y=0.74 $X2=0 $Y2=0
cc_667 N_A_c_883_n N_A_1024_74#_c_1042_n 5.25256e-19 $X=6.64 $Y=1.705 $X2=0
+ $Y2=0
cc_668 N_A_M1002_g N_A_1024_74#_c_1043_n 0.00698694f $X=6.625 $Y=0.74 $X2=0
+ $Y2=0
cc_669 N_A_c_883_n N_A_1024_74#_c_1043_n 0.0148403f $X=6.64 $Y=1.705 $X2=0 $Y2=0
cc_670 N_A_M1003_g N_A_27_392#_c_1193_n 0.00407809f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_671 A N_A_27_392#_c_1193_n 0.0290526f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_672 N_A_c_887_n N_A_27_392#_c_1193_n 0.00143639f $X=0.63 $Y=1.41 $X2=0 $Y2=0
cc_673 N_A_M1003_g N_A_27_392#_c_1194_n 0.0108661f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_674 N_A_M1003_g N_A_27_392#_c_1202_n 0.0146031f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_675 A N_A_27_392#_c_1202_n 0.0184173f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_676 N_A_c_887_n N_A_27_392#_c_1202_n 7.35771e-19 $X=0.63 $Y=1.41 $X2=0 $Y2=0
cc_677 N_A_M1003_g N_A_27_392#_c_1203_n 0.00149436f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_678 N_A_c_889_n N_A_27_392#_c_1195_n 0.00262007f $X=3.02 $Y=3.15 $X2=0 $Y2=0
cc_679 N_A_c_889_n N_A_27_392#_c_1196_n 0.0177535f $X=3.02 $Y=3.15 $X2=0 $Y2=0
cc_680 A N_VPWR_M1003_d 6.98785e-19 $X=0.635 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_681 N_A_M1003_g N_VPWR_c_1242_n 0.0031197f $X=0.505 $Y=2.46 $X2=0 $Y2=0
cc_682 N_A_c_889_n N_VPWR_c_1242_n 0.0155821f $X=3.02 $Y=3.15 $X2=0 $Y2=0
cc_683 N_A_M1005_g N_VPWR_c_1243_n 0.0313955f $X=3.11 $Y=2.235 $X2=0 $Y2=0
cc_684 N_A_c_892_n N_VPWR_c_1243_n 0.0177656f $X=4.54 $Y=3.15 $X2=0 $Y2=0
cc_685 N_A_c_898_n N_VPWR_c_1243_n 0.00476669f $X=3.11 $Y=3.15 $X2=0 $Y2=0
cc_686 N_A_c_892_n N_VPWR_c_1244_n 0.021565f $X=4.54 $Y=3.15 $X2=0 $Y2=0
cc_687 N_A_M1004_g N_VPWR_c_1244_n 0.0219822f $X=4.63 $Y=2.235 $X2=0 $Y2=0
cc_688 N_A_c_899_n N_VPWR_c_1244_n 0.00477316f $X=4.63 $Y=3.15 $X2=0 $Y2=0
cc_689 N_A_M1018_g N_VPWR_c_1245_n 0.026294f $X=6.64 $Y=2.34 $X2=0 $Y2=0
cc_690 N_A_c_889_n N_VPWR_c_1251_n 0.0663415f $X=3.02 $Y=3.15 $X2=0 $Y2=0
cc_691 N_A_c_892_n N_VPWR_c_1253_n 0.0199069f $X=4.54 $Y=3.15 $X2=0 $Y2=0
cc_692 N_A_c_899_n N_VPWR_c_1254_n 0.0706703f $X=4.63 $Y=3.15 $X2=0 $Y2=0
cc_693 N_A_c_890_n N_VPWR_c_1259_n 0.00853352f $X=0.595 $Y=3.15 $X2=0 $Y2=0
cc_694 N_A_c_889_n N_VPWR_c_1241_n 0.0761827f $X=3.02 $Y=3.15 $X2=0 $Y2=0
cc_695 N_A_c_890_n N_VPWR_c_1241_n 0.011799f $X=0.595 $Y=3.15 $X2=0 $Y2=0
cc_696 N_A_c_892_n N_VPWR_c_1241_n 0.0200963f $X=4.54 $Y=3.15 $X2=0 $Y2=0
cc_697 N_A_c_894_n N_VPWR_c_1241_n 0.0846502f $X=6.55 $Y=3.15 $X2=0 $Y2=0
cc_698 N_A_c_898_n N_VPWR_c_1241_n 0.00904288f $X=3.11 $Y=3.15 $X2=0 $Y2=0
cc_699 N_A_c_899_n N_VPWR_c_1241_n 0.00904288f $X=4.63 $Y=3.15 $X2=0 $Y2=0
cc_700 N_A_M1004_g N_A_740_347#_c_1390_n 0.014943f $X=4.63 $Y=2.235 $X2=0 $Y2=0
cc_701 N_A_M1004_g N_A_740_347#_c_1386_n 3.31317e-19 $X=4.63 $Y=2.235 $X2=0
+ $Y2=0
cc_702 N_A_c_894_n N_A_740_347#_c_1386_n 0.00473258f $X=6.55 $Y=3.15 $X2=0 $Y2=0
cc_703 N_A_c_892_n N_A_740_347#_c_1387_n 0.00562388f $X=4.54 $Y=3.15 $X2=0 $Y2=0
cc_704 N_A_M1004_g N_A_740_347#_c_1387_n 7.72743e-19 $X=4.63 $Y=2.235 $X2=0
+ $Y2=0
cc_705 N_A_M1018_g N_SUM_c_1427_n 0.00102531f $X=6.64 $Y=2.34 $X2=0 $Y2=0
cc_706 N_A_M1034_g N_A_27_74#_c_1554_n 0.0205742f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_707 A N_A_27_74#_c_1554_n 0.0246165f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_708 N_A_c_887_n N_A_27_74#_c_1554_n 0.00671825f $X=0.63 $Y=1.41 $X2=0 $Y2=0
cc_709 N_A_M1034_g N_A_27_74#_c_1557_n 0.0120858f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_710 A N_A_27_74#_c_1557_n 0.0119709f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_711 N_A_c_887_n N_A_27_74#_c_1557_n 0.003838f $X=0.63 $Y=1.41 $X2=0 $Y2=0
cc_712 N_A_c_884_n N_VGND_c_1585_n 0.010869f $X=3.11 $Y=1.185 $X2=0 $Y2=0
cc_713 N_A_c_884_n N_VGND_c_1589_n 0.00383152f $X=3.11 $Y=1.185 $X2=0 $Y2=0
cc_714 N_A_c_885_n N_VGND_c_1591_n 0.0023296f $X=4.63 $Y=1.185 $X2=0 $Y2=0
cc_715 N_A_M1002_g N_VGND_c_1593_n 0.00320129f $X=6.625 $Y=0.74 $X2=0 $Y2=0
cc_716 N_A_c_885_n N_VGND_c_1593_n 0.00316493f $X=4.63 $Y=1.185 $X2=0 $Y2=0
cc_717 N_A_M1034_g N_VGND_c_1598_n 0.00316493f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_718 N_A_M1034_g N_VGND_c_1599_n 0.00608124f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_719 N_A_M1002_g N_VGND_c_1600_n 0.00253998f $X=6.625 $Y=0.74 $X2=0 $Y2=0
cc_720 N_A_M1034_g N_VGND_c_1604_n 0.00400459f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_721 N_A_M1002_g N_VGND_c_1604_n 0.00405511f $X=6.625 $Y=0.74 $X2=0 $Y2=0
cc_722 N_A_c_884_n N_VGND_c_1604_n 0.00384996f $X=3.11 $Y=1.185 $X2=0 $Y2=0
cc_723 N_A_c_885_n N_VGND_c_1604_n 0.00393316f $X=4.63 $Y=1.185 $X2=0 $Y2=0
cc_724 N_A_c_885_n N_A_734_74#_c_1734_n 0.00936301f $X=4.63 $Y=1.185 $X2=0 $Y2=0
cc_725 N_A_c_885_n N_A_734_74#_c_1732_n 8.6409e-19 $X=4.63 $Y=1.185 $X2=0 $Y2=0
cc_726 N_A_c_885_n N_A_734_74#_c_1733_n 0.0057442f $X=4.63 $Y=1.185 $X2=0 $Y2=0
cc_727 N_A_1024_74#_c_1059_n N_VPWR_M1018_d 0.00862083f $X=6.905 $Y=2.035 $X2=0
+ $Y2=0
cc_728 N_A_1024_74#_c_1048_n N_VPWR_M1018_d 0.00197943f $X=6.99 $Y=1.95 $X2=0
+ $Y2=0
cc_729 N_A_1024_74#_M1007_g N_VPWR_c_1245_n 0.00314456f $X=7.185 $Y=2.4 $X2=0
+ $Y2=0
cc_730 N_A_1024_74#_c_1059_n N_VPWR_c_1245_n 0.020778f $X=6.905 $Y=2.035 $X2=0
+ $Y2=0
cc_731 N_A_1024_74#_M1008_g N_VPWR_c_1246_n 0.00346635f $X=7.635 $Y=2.4 $X2=0
+ $Y2=0
cc_732 N_A_1024_74#_M1010_g N_VPWR_c_1246_n 0.00360947f $X=8.135 $Y=2.4 $X2=0
+ $Y2=0
cc_733 N_A_1024_74#_M1020_g N_VPWR_c_1247_n 0.00348414f $X=8.585 $Y=2.4 $X2=0
+ $Y2=0
cc_734 N_A_1024_74#_c_1043_n N_VPWR_c_1247_n 5.712e-19 $X=8.585 $Y=1.505 $X2=0
+ $Y2=0
cc_735 N_A_1024_74#_c_1050_n N_VPWR_c_1254_n 0.00749501f $X=5.405 $Y=2.145 $X2=0
+ $Y2=0
cc_736 N_A_1024_74#_M1007_g N_VPWR_c_1255_n 0.005209f $X=7.185 $Y=2.4 $X2=0
+ $Y2=0
cc_737 N_A_1024_74#_M1008_g N_VPWR_c_1255_n 0.005209f $X=7.635 $Y=2.4 $X2=0
+ $Y2=0
cc_738 N_A_1024_74#_M1010_g N_VPWR_c_1256_n 0.005209f $X=8.135 $Y=2.4 $X2=0
+ $Y2=0
cc_739 N_A_1024_74#_M1020_g N_VPWR_c_1256_n 0.005209f $X=8.585 $Y=2.4 $X2=0
+ $Y2=0
cc_740 N_A_1024_74#_M1007_g N_VPWR_c_1241_n 0.00983208f $X=7.185 $Y=2.4 $X2=0
+ $Y2=0
cc_741 N_A_1024_74#_M1008_g N_VPWR_c_1241_n 0.00982754f $X=7.635 $Y=2.4 $X2=0
+ $Y2=0
cc_742 N_A_1024_74#_M1010_g N_VPWR_c_1241_n 0.00982082f $X=8.135 $Y=2.4 $X2=0
+ $Y2=0
cc_743 N_A_1024_74#_M1020_g N_VPWR_c_1241_n 0.00982832f $X=8.585 $Y=2.4 $X2=0
+ $Y2=0
cc_744 N_A_1024_74#_c_1050_n N_VPWR_c_1241_n 0.009077f $X=5.405 $Y=2.145 $X2=0
+ $Y2=0
cc_745 N_A_1024_74#_c_1050_n N_A_740_347#_c_1386_n 0.0195141f $X=5.405 $Y=2.145
+ $X2=0 $Y2=0
cc_746 N_A_1024_74#_c_1053_n A_1144_347# 0.00856328f $X=6.255 $Y=2.145 $X2=-0.19
+ $Y2=-0.245
cc_747 N_A_1024_74#_c_1053_n A_1238_347# 8.21762e-19 $X=6.255 $Y=2.145 $X2=-0.19
+ $Y2=-0.245
cc_748 N_A_1024_74#_c_1059_n A_1238_347# 0.00373218f $X=6.905 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_749 N_A_1024_74#_c_1067_n A_1238_347# 0.0117621f $X=6.34 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_750 N_A_1024_74#_M1007_g N_SUM_c_1426_n 0.0023456f $X=7.185 $Y=2.4 $X2=0
+ $Y2=0
cc_751 N_A_1024_74#_M1008_g N_SUM_c_1426_n 8.84614e-19 $X=7.635 $Y=2.4 $X2=0
+ $Y2=0
cc_752 N_A_1024_74#_c_1041_n N_SUM_c_1426_n 0.0218858f $X=7.94 $Y=1.505 $X2=0
+ $Y2=0
cc_753 N_A_1024_74#_c_1043_n N_SUM_c_1426_n 0.00215577f $X=8.585 $Y=1.505 $X2=0
+ $Y2=0
cc_754 N_A_1024_74#_M1007_g N_SUM_c_1427_n 0.0138838f $X=7.185 $Y=2.4 $X2=0
+ $Y2=0
cc_755 N_A_1024_74#_M1008_g N_SUM_c_1427_n 0.0138483f $X=7.635 $Y=2.4 $X2=0
+ $Y2=0
cc_756 N_A_1024_74#_M1010_g N_SUM_c_1427_n 6.68421e-19 $X=8.135 $Y=2.4 $X2=0
+ $Y2=0
cc_757 N_A_1024_74#_M1022_g N_SUM_c_1423_n 0.0035804f $X=7.215 $Y=0.78 $X2=0
+ $Y2=0
cc_758 N_A_1024_74#_M1024_g N_SUM_c_1423_n 0.0120038f $X=7.645 $Y=0.78 $X2=0
+ $Y2=0
cc_759 N_A_1024_74#_M1036_g N_SUM_c_1423_n 0.0122903f $X=8.235 $Y=0.78 $X2=0
+ $Y2=0
cc_760 N_A_1024_74#_c_1056_n N_SUM_c_1423_n 0.0135437f $X=6.905 $Y=1.005 $X2=0
+ $Y2=0
cc_761 N_A_1024_74#_c_1040_n N_SUM_c_1423_n 0.00568635f $X=6.99 $Y=1.34 $X2=0
+ $Y2=0
cc_762 N_A_1024_74#_c_1041_n N_SUM_c_1423_n 0.064353f $X=7.94 $Y=1.505 $X2=0
+ $Y2=0
cc_763 N_A_1024_74#_c_1043_n N_SUM_c_1423_n 0.00871607f $X=8.585 $Y=1.505 $X2=0
+ $Y2=0
cc_764 N_A_1024_74#_M1008_g N_SUM_c_1454_n 0.0132272f $X=7.635 $Y=2.4 $X2=0
+ $Y2=0
cc_765 N_A_1024_74#_M1010_g N_SUM_c_1454_n 0.0145392f $X=8.135 $Y=2.4 $X2=0
+ $Y2=0
cc_766 N_A_1024_74#_c_1041_n N_SUM_c_1454_n 0.0344509f $X=7.94 $Y=1.505 $X2=0
+ $Y2=0
cc_767 N_A_1024_74#_c_1043_n N_SUM_c_1454_n 0.00313888f $X=8.585 $Y=1.505 $X2=0
+ $Y2=0
cc_768 N_A_1024_74#_M1036_g N_SUM_c_1424_n 0.00114171f $X=8.235 $Y=0.78 $X2=0
+ $Y2=0
cc_769 N_A_1024_74#_M1038_g N_SUM_c_1424_n 0.00537066f $X=8.665 $Y=0.78 $X2=0
+ $Y2=0
cc_770 N_A_1024_74#_M1024_g N_SUM_c_1425_n 7.63771e-19 $X=7.645 $Y=0.78 $X2=0
+ $Y2=0
cc_771 N_A_1024_74#_M1010_g N_SUM_c_1425_n 0.00428339f $X=8.135 $Y=2.4 $X2=0
+ $Y2=0
cc_772 N_A_1024_74#_M1036_g N_SUM_c_1425_n 0.00486056f $X=8.235 $Y=0.78 $X2=0
+ $Y2=0
cc_773 N_A_1024_74#_M1020_g N_SUM_c_1425_n 0.0045348f $X=8.585 $Y=2.4 $X2=0
+ $Y2=0
cc_774 N_A_1024_74#_M1038_g N_SUM_c_1425_n 0.00183896f $X=8.665 $Y=0.78 $X2=0
+ $Y2=0
cc_775 N_A_1024_74#_c_1041_n N_SUM_c_1425_n 0.0244401f $X=7.94 $Y=1.505 $X2=0
+ $Y2=0
cc_776 N_A_1024_74#_c_1043_n N_SUM_c_1425_n 0.021524f $X=8.585 $Y=1.505 $X2=0
+ $Y2=0
cc_777 N_A_1024_74#_M1010_g SUM 0.00128801f $X=8.135 $Y=2.4 $X2=0 $Y2=0
cc_778 N_A_1024_74#_M1020_g SUM 0.00204309f $X=8.585 $Y=2.4 $X2=0 $Y2=0
cc_779 N_A_1024_74#_M1008_g SUM 6.37103e-19 $X=7.635 $Y=2.4 $X2=0 $Y2=0
cc_780 N_A_1024_74#_M1010_g SUM 0.0132857f $X=8.135 $Y=2.4 $X2=0 $Y2=0
cc_781 N_A_1024_74#_M1020_g SUM 0.0124584f $X=8.585 $Y=2.4 $X2=0 $Y2=0
cc_782 N_A_1024_74#_M1038_g N_COUT_c_1484_n 9.32329e-19 $X=8.665 $Y=0.78 $X2=0
+ $Y2=0
cc_783 N_A_1024_74#_c_1056_n N_VGND_M1002_d 0.0123197f $X=6.905 $Y=1.005 $X2=0
+ $Y2=0
cc_784 N_A_1024_74#_c_1040_n N_VGND_M1002_d 0.00175048f $X=6.99 $Y=1.34 $X2=0
+ $Y2=0
cc_785 N_A_1024_74#_M1022_g N_VGND_c_1594_n 0.00414982f $X=7.215 $Y=0.78 $X2=0
+ $Y2=0
cc_786 N_A_1024_74#_M1024_g N_VGND_c_1594_n 0.00414982f $X=7.645 $Y=0.78 $X2=0
+ $Y2=0
cc_787 N_A_1024_74#_M1036_g N_VGND_c_1595_n 0.00414982f $X=8.235 $Y=0.78 $X2=0
+ $Y2=0
cc_788 N_A_1024_74#_M1038_g N_VGND_c_1595_n 0.00414982f $X=8.665 $Y=0.78 $X2=0
+ $Y2=0
cc_789 N_A_1024_74#_M1022_g N_VGND_c_1600_n 0.00378066f $X=7.215 $Y=0.78 $X2=0
+ $Y2=0
cc_790 N_A_1024_74#_M1024_g N_VGND_c_1601_n 0.00378066f $X=7.645 $Y=0.78 $X2=0
+ $Y2=0
cc_791 N_A_1024_74#_M1036_g N_VGND_c_1601_n 0.00378066f $X=8.235 $Y=0.78 $X2=0
+ $Y2=0
cc_792 N_A_1024_74#_M1038_g N_VGND_c_1602_n 0.00378066f $X=8.665 $Y=0.78 $X2=0
+ $Y2=0
cc_793 N_A_1024_74#_M1022_g N_VGND_c_1604_n 0.00533081f $X=7.215 $Y=0.78 $X2=0
+ $Y2=0
cc_794 N_A_1024_74#_M1024_g N_VGND_c_1604_n 0.00533081f $X=7.645 $Y=0.78 $X2=0
+ $Y2=0
cc_795 N_A_1024_74#_M1036_g N_VGND_c_1604_n 0.00533081f $X=8.235 $Y=0.78 $X2=0
+ $Y2=0
cc_796 N_A_1024_74#_M1038_g N_VGND_c_1604_n 0.00533081f $X=8.665 $Y=0.78 $X2=0
+ $Y2=0
cc_797 N_A_1024_74#_c_1077_n A_1160_74# 0.00308137f $X=5.915 $Y=0.965 $X2=-0.19
+ $Y2=-0.245
cc_798 N_A_1024_74#_c_1065_n A_1160_74# 0.00302066f $X=6.085 $Y=0.965 $X2=-0.19
+ $Y2=-0.245
cc_799 N_A_1024_74#_c_1056_n A_1238_74# 0.00608853f $X=6.905 $Y=1.005 $X2=-0.19
+ $Y2=-0.245
cc_800 N_A_27_392#_c_1202_n N_VPWR_M1003_d 0.0180809f $X=0.985 $Y=2.17 $X2=-0.19
+ $Y2=1.66
cc_801 N_A_27_392#_c_1203_n N_VPWR_M1003_d 0.00422093f $X=1.07 $Y=2.63 $X2=-0.19
+ $Y2=1.66
cc_802 N_A_27_392#_c_1195_n N_VPWR_M1003_d 9.96039e-19 $X=1.155 $Y=2.795
+ $X2=-0.19 $Y2=1.66
cc_803 N_A_27_392#_c_1194_n N_VPWR_c_1242_n 0.0189222f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_804 N_A_27_392#_c_1202_n N_VPWR_c_1242_n 0.0131801f $X=0.985 $Y=2.17 $X2=0
+ $Y2=0
cc_805 N_A_27_392#_c_1203_n N_VPWR_c_1242_n 0.0148533f $X=1.07 $Y=2.63 $X2=0
+ $Y2=0
cc_806 N_A_27_392#_c_1195_n N_VPWR_c_1242_n 0.0272459f $X=1.155 $Y=2.795 $X2=0
+ $Y2=0
cc_807 N_A_27_392#_c_1195_n N_VPWR_c_1251_n 0.00701426f $X=1.155 $Y=2.795 $X2=0
+ $Y2=0
cc_808 N_A_27_392#_c_1196_n N_VPWR_c_1251_n 0.0331696f $X=1.84 $Y=2.795 $X2=0
+ $Y2=0
cc_809 N_A_27_392#_c_1194_n N_VPWR_c_1259_n 0.014549f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_810 N_A_27_392#_c_1194_n N_VPWR_c_1241_n 0.0119743f $X=0.28 $Y=2.815 $X2=0
+ $Y2=0
cc_811 N_A_27_392#_c_1195_n N_VPWR_c_1241_n 0.00552059f $X=1.155 $Y=2.795 $X2=0
+ $Y2=0
cc_812 N_A_27_392#_c_1196_n N_VPWR_c_1241_n 0.0268277f $X=1.84 $Y=2.795 $X2=0
+ $Y2=0
cc_813 N_VPWR_M1012_d N_A_740_347#_c_1390_n 0.00606391f $X=4.15 $Y=1.735 $X2=0
+ $Y2=0
cc_814 N_VPWR_c_1244_n N_A_740_347#_c_1390_n 0.0246219f $X=4.37 $Y=2.59 $X2=0
+ $Y2=0
cc_815 N_VPWR_c_1244_n N_A_740_347#_c_1386_n 0.0135428f $X=4.37 $Y=2.59 $X2=0
+ $Y2=0
cc_816 N_VPWR_c_1254_n N_A_740_347#_c_1386_n 0.00747717f $X=6.795 $Y=3.33 $X2=0
+ $Y2=0
cc_817 N_VPWR_c_1241_n N_A_740_347#_c_1386_n 0.00905985f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_818 N_VPWR_c_1243_n N_A_740_347#_c_1387_n 0.0195141f $X=3.335 $Y=2.17 $X2=0
+ $Y2=0
cc_819 N_VPWR_c_1244_n N_A_740_347#_c_1387_n 0.0131962f $X=4.37 $Y=2.59 $X2=0
+ $Y2=0
cc_820 N_VPWR_c_1253_n N_A_740_347#_c_1387_n 0.00740628f $X=4.17 $Y=3.33 $X2=0
+ $Y2=0
cc_821 N_VPWR_c_1241_n N_A_740_347#_c_1387_n 0.00902643f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_822 N_VPWR_c_1245_n N_SUM_c_1427_n 0.0234083f $X=6.96 $Y=2.455 $X2=0 $Y2=0
cc_823 N_VPWR_c_1246_n N_SUM_c_1427_n 0.0270323f $X=7.86 $Y=2.345 $X2=0 $Y2=0
cc_824 N_VPWR_c_1255_n N_SUM_c_1427_n 0.0144623f $X=7.775 $Y=3.33 $X2=0 $Y2=0
cc_825 N_VPWR_c_1241_n N_SUM_c_1427_n 0.0118344f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_826 N_VPWR_M1008_s N_SUM_c_1454_n 0.0040648f $X=7.725 $Y=1.84 $X2=0 $Y2=0
cc_827 N_VPWR_c_1246_n N_SUM_c_1454_n 0.0167599f $X=7.86 $Y=2.345 $X2=0 $Y2=0
cc_828 N_VPWR_c_1247_n N_SUM_c_1425_n 0.00127217f $X=8.81 $Y=1.985 $X2=0 $Y2=0
cc_829 N_VPWR_c_1246_n SUM 0.0307758f $X=7.86 $Y=2.345 $X2=0 $Y2=0
cc_830 N_VPWR_c_1247_n SUM 0.0326001f $X=8.81 $Y=1.985 $X2=0 $Y2=0
cc_831 N_VPWR_c_1256_n SUM 0.0144623f $X=8.725 $Y=3.33 $X2=0 $Y2=0
cc_832 N_VPWR_c_1241_n SUM 0.0118344f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_833 N_VPWR_c_1247_n N_COUT_c_1488_n 0.00792222f $X=8.81 $Y=1.985 $X2=0 $Y2=0
cc_834 N_VPWR_c_1247_n N_COUT_c_1489_n 0.0378676f $X=8.81 $Y=1.985 $X2=0 $Y2=0
cc_835 N_VPWR_c_1248_n N_COUT_c_1489_n 0.0276912f $X=9.76 $Y=2.325 $X2=0 $Y2=0
cc_836 N_VPWR_c_1257_n N_COUT_c_1489_n 0.0144623f $X=9.675 $Y=3.33 $X2=0 $Y2=0
cc_837 N_VPWR_c_1241_n N_COUT_c_1489_n 0.0118344f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_838 N_VPWR_M1019_d N_COUT_c_1490_n 0.00218982f $X=9.625 $Y=1.84 $X2=0 $Y2=0
cc_839 N_VPWR_c_1248_n N_COUT_c_1490_n 0.0167599f $X=9.76 $Y=2.325 $X2=0 $Y2=0
cc_840 N_VPWR_c_1250_n N_COUT_c_1491_n 0.00725063f $X=10.71 $Y=1.985 $X2=0 $Y2=0
cc_841 N_VPWR_c_1248_n COUT 0.0316672f $X=9.76 $Y=2.325 $X2=0 $Y2=0
cc_842 N_VPWR_c_1250_n COUT 0.0348023f $X=10.71 $Y=1.985 $X2=0 $Y2=0
cc_843 N_VPWR_c_1258_n COUT 0.0148786f $X=10.625 $Y=3.33 $X2=0 $Y2=0
cc_844 N_VPWR_c_1241_n COUT 0.0121555f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_845 N_VPWR_c_1250_n N_VGND_c_1588_n 0.00906267f $X=10.71 $Y=1.985 $X2=0 $Y2=0
cc_846 N_SUM_c_1423_n N_VGND_M1024_d 0.00452945f $X=8.285 $Y=1.045 $X2=0 $Y2=0
cc_847 N_COUT_c_1506_n N_VGND_M1014_s 0.00356752f $X=10.165 $Y=1.065 $X2=0 $Y2=0
cc_848 N_COUT_c_1484_n N_VGND_c_1586_n 0.0151543f $X=9.47 $Y=0.555 $X2=0 $Y2=0
cc_849 N_COUT_c_1506_n N_VGND_c_1586_n 0.0152916f $X=10.165 $Y=1.065 $X2=0 $Y2=0
cc_850 N_COUT_c_1486_n N_VGND_c_1586_n 0.0152413f $X=10.33 $Y=0.555 $X2=0 $Y2=0
cc_851 N_COUT_c_1486_n N_VGND_c_1588_n 0.0229007f $X=10.33 $Y=0.555 $X2=0 $Y2=0
cc_852 N_COUT_c_1487_n N_VGND_c_1588_n 0.00151292f $X=10.295 $Y=1.55 $X2=0 $Y2=0
cc_853 N_COUT_c_1484_n N_VGND_c_1596_n 0.00946322f $X=9.47 $Y=0.555 $X2=0 $Y2=0
cc_854 N_COUT_c_1486_n N_VGND_c_1597_n 0.00984752f $X=10.33 $Y=0.555 $X2=0 $Y2=0
cc_855 N_COUT_c_1484_n N_VGND_c_1602_n 0.00148615f $X=9.47 $Y=0.555 $X2=0 $Y2=0
cc_856 N_COUT_c_1484_n N_VGND_c_1604_n 0.00891381f $X=9.47 $Y=0.555 $X2=0 $Y2=0
cc_857 N_COUT_c_1486_n N_VGND_c_1604_n 0.0092741f $X=10.33 $Y=0.555 $X2=0 $Y2=0
cc_858 N_A_27_74#_c_1557_n N_VGND_M1034_d 0.0262462f $X=1.325 $Y=0.55 $X2=-0.19
+ $Y2=-0.245
cc_859 N_A_27_74#_c_1555_n N_VGND_M1034_d 0.00943635f $X=1.495 $Y=0.55 $X2=-0.19
+ $Y2=-0.245
cc_860 N_A_27_74#_c_1557_n N_VGND_c_1589_n 0.003347f $X=1.325 $Y=0.55 $X2=0
+ $Y2=0
cc_861 N_A_27_74#_c_1555_n N_VGND_c_1589_n 0.0265731f $X=1.495 $Y=0.55 $X2=0
+ $Y2=0
cc_862 N_A_27_74#_c_1554_n N_VGND_c_1598_n 0.0145639f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_863 N_A_27_74#_c_1557_n N_VGND_c_1598_n 0.00294077f $X=1.325 $Y=0.55 $X2=0
+ $Y2=0
cc_864 N_A_27_74#_c_1554_n N_VGND_c_1599_n 0.00294333f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_865 N_A_27_74#_c_1557_n N_VGND_c_1599_n 0.0392999f $X=1.325 $Y=0.55 $X2=0
+ $Y2=0
cc_866 N_A_27_74#_c_1555_n N_VGND_c_1599_n 0.00517613f $X=1.495 $Y=0.55 $X2=0
+ $Y2=0
cc_867 N_A_27_74#_c_1554_n N_VGND_c_1604_n 0.0119984f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_868 N_A_27_74#_c_1557_n N_VGND_c_1604_n 0.0124477f $X=1.325 $Y=0.55 $X2=0
+ $Y2=0
cc_869 N_A_27_74#_c_1555_n N_VGND_c_1604_n 0.022248f $X=1.495 $Y=0.55 $X2=0
+ $Y2=0
cc_870 N_VGND_M1033_d N_A_734_74#_c_1734_n 0.0072679f $X=4.1 $Y=0.37 $X2=0 $Y2=0
cc_871 N_VGND_c_1591_n N_A_734_74#_c_1734_n 0.0243979f $X=4.32 $Y=0 $X2=0 $Y2=0
cc_872 N_VGND_c_1592_n N_A_734_74#_c_1734_n 0.0029521f $X=4.155 $Y=0 $X2=0 $Y2=0
cc_873 N_VGND_c_1593_n N_A_734_74#_c_1734_n 0.0029521f $X=6.755 $Y=0 $X2=0 $Y2=0
cc_874 N_VGND_c_1604_n N_A_734_74#_c_1734_n 0.011204f $X=10.8 $Y=0 $X2=0 $Y2=0
cc_875 N_VGND_c_1585_n N_A_734_74#_c_1732_n 0.00129215f $X=3.34 $Y=0.55 $X2=0
+ $Y2=0
cc_876 N_VGND_c_1591_n N_A_734_74#_c_1732_n 0.00282013f $X=4.32 $Y=0 $X2=0 $Y2=0
cc_877 N_VGND_c_1592_n N_A_734_74#_c_1732_n 0.0105866f $X=4.155 $Y=0 $X2=0 $Y2=0
cc_878 N_VGND_c_1604_n N_A_734_74#_c_1732_n 0.00888607f $X=10.8 $Y=0 $X2=0 $Y2=0
cc_879 N_VGND_c_1591_n N_A_734_74#_c_1733_n 0.00282013f $X=4.32 $Y=0 $X2=0 $Y2=0
cc_880 N_VGND_c_1593_n N_A_734_74#_c_1733_n 0.0105866f $X=6.755 $Y=0 $X2=0 $Y2=0
cc_881 N_VGND_c_1604_n N_A_734_74#_c_1733_n 0.00888607f $X=10.8 $Y=0 $X2=0 $Y2=0

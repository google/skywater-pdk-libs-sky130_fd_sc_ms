* File: sky130_fd_sc_ms__fa_4.pex.spice
* Created: Fri Aug 28 17:35:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__FA_4%B 3 7 11 15 19 23 27 31 33 39 40 41 44 45 47 51
+ 52 54 56 58 59 66 75
c232 75 0 1.67591e-19 $X=6.175 $Y=1.41
c233 59 0 1.72486e-19 $X=6.48 $Y=1.665
c234 56 0 1.26815e-19 $X=4.62 $Y=1.805
c235 51 0 6.08971e-20 $X=4.115 $Y=1.41
c236 44 0 1.16364e-19 $X=2.645 $Y=1.41
c237 33 0 2.07083e-19 $X=1.665 $Y=1.417
c238 3 0 1.28731e-19 $X=1.155 $Y=2.235
r239 75 78 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.175 $Y=1.41
+ $X2=6.175 $Y2=1.575
r240 75 77 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.175 $Y=1.41
+ $X2=6.175 $Y2=1.245
r241 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.175
+ $Y=1.41 $X2=6.175 $Y2=1.41
r242 59 76 8.49543 $w=4.38e-07 $l=3.05e-07 $layer=LI1_cond $X=6.48 $Y=1.575
+ $X2=6.175 $Y2=1.575
r243 58 76 4.87443 $w=4.38e-07 $l=1.75e-07 $layer=LI1_cond $X=6 $Y=1.575
+ $X2=6.175 $Y2=1.575
r244 56 58 72.095 $w=1.98e-07 $l=1.295e-06 $layer=LI1_cond $X=4.62 $Y=1.805
+ $X2=5.915 $Y2=1.805
r245 54 55 10.3347 $w=2.42e-07 $l=2.05e-07 $layer=LI1_cond $X=2.645 $Y=1.83
+ $X2=2.645 $Y2=2.035
r246 52 73 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.115 $Y=1.41
+ $X2=4.115 $Y2=1.575
r247 52 72 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.115 $Y=1.41
+ $X2=4.115 $Y2=1.245
r248 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.115
+ $Y=1.41 $X2=4.115 $Y2=1.41
r249 49 56 35.0057 $w=1.76e-07 $l=5.10965e-07 $layer=LI1_cond $X=4.115 $Y=1.817
+ $X2=4.62 $Y2=1.805
r250 49 51 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.115 $Y=1.745
+ $X2=4.115 $Y2=1.41
r251 48 54 2.80567 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.81 $Y=1.83
+ $X2=2.645 $Y2=1.83
r252 47 49 11.4375 $w=1.76e-07 $l=1.71377e-07 $layer=LI1_cond $X=3.95 $Y=1.83
+ $X2=4.115 $Y2=1.817
r253 47 48 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=3.95 $Y=1.83
+ $X2=2.81 $Y2=1.83
r254 45 70 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.41
+ $X2=2.645 $Y2=1.575
r255 45 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.41
+ $X2=2.645 $Y2=1.245
r256 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.645
+ $Y=1.41 $X2=2.645 $Y2=1.41
r257 42 54 4.03333 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.645 $Y=1.745
+ $X2=2.645 $Y2=1.83
r258 42 44 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.645 $Y=1.745
+ $X2=2.645 $Y2=1.41
r259 40 55 2.80567 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.48 $Y=2.035
+ $X2=2.645 $Y2=2.035
r260 40 41 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=2.48 $Y=2.035
+ $X2=1.835 $Y2=2.035
r261 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.75 $Y=1.95
+ $X2=1.835 $Y2=2.035
r262 38 39 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.75 $Y=1.575
+ $X2=1.75 $Y2=1.95
r263 36 66 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.51 $Y=1.41
+ $X2=1.585 $Y2=1.41
r264 36 63 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.51 $Y=1.41
+ $X2=1.155 $Y2=1.41
r265 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.51
+ $Y=1.41 $X2=1.51 $Y2=1.41
r266 33 38 7.64049 $w=3.15e-07 $l=1.95944e-07 $layer=LI1_cond $X=1.665 $Y=1.417
+ $X2=1.75 $Y2=1.575
r267 33 35 5.67075 $w=3.13e-07 $l=1.55e-07 $layer=LI1_cond $X=1.665 $Y=1.417
+ $X2=1.51 $Y2=1.417
r268 31 77 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.115 $Y=0.74
+ $X2=6.115 $Y2=1.245
r269 27 78 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=6.1 $Y=2.235
+ $X2=6.1 $Y2=1.575
r270 23 73 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=4.06 $Y=2.235
+ $X2=4.06 $Y2=1.575
r271 19 72 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.025 $Y=0.74
+ $X2=4.025 $Y2=1.245
r272 15 70 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.6 $Y=2.235
+ $X2=2.6 $Y2=1.575
r273 11 69 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.585 $Y=0.74
+ $X2=2.585 $Y2=1.245
r274 5 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=1.245
+ $X2=1.585 $Y2=1.41
r275 5 7 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.585 $Y=1.245
+ $X2=1.585 $Y2=0.74
r276 1 63 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=1.575
+ $X2=1.155 $Y2=1.41
r277 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.155 $Y=1.575
+ $X2=1.155 $Y2=2.235
.ends

.subckt PM_SKY130_FD_SC_MS__FA_4%CIN 3 6 10 14 18 22 25 26 28 29 30 31 36 37 39
+ 42 44 50 52 55 64
c161 37 0 9.09194e-20 $X=5.52 $Y=1.295
c162 18 0 2.27929e-19 $X=5.63 $Y=2.235
c163 10 0 1.78103e-19 $X=3.595 $Y=0.74
c164 6 0 1.64344e-19 $X=2.15 $Y=2.235
r165 50 53 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.635 $Y=1.385
+ $X2=5.635 $Y2=1.55
r166 50 52 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.635 $Y=1.385
+ $X2=5.635 $Y2=1.22
r167 42 45 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.105 $Y=1.385
+ $X2=2.105 $Y2=1.55
r168 42 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.105 $Y=1.385
+ $X2=2.105 $Y2=1.22
r169 42 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.105
+ $Y=1.385 $X2=2.105 $Y2=1.385
r170 39 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=1.295
+ $X2=2.16 $Y2=1.295
r171 37 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.635
+ $Y=1.385 $X2=5.635 $Y2=1.385
r172 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.295
+ $X2=5.52 $Y2=1.295
r173 34 64 3.27739 $w=3.93e-07 $l=9.5e-08 $layer=LI1_cond $X=3.12 $Y=1.377
+ $X2=3.215 $Y2=1.377
r174 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=1.295
+ $X2=3.12 $Y2=1.295
r175 31 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.265 $Y=1.295
+ $X2=3.12 $Y2=1.295
r176 30 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=1.295
+ $X2=5.52 $Y2=1.295
r177 30 31 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=5.375 $Y=1.295
+ $X2=3.265 $Y2=1.295
r178 29 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=1.295
+ $X2=2.16 $Y2=1.295
r179 28 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.975 $Y=1.295
+ $X2=3.12 $Y2=1.295
r180 28 29 0.829206 $w=1.4e-07 $l=6.7e-07 $layer=MET1_cond $X=2.975 $Y=1.295
+ $X2=2.305 $Y2=1.295
r181 26 48 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.575 $Y=1.41
+ $X2=3.575 $Y2=1.575
r182 26 47 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.575 $Y=1.41
+ $X2=3.575 $Y2=1.245
r183 25 64 13.1708 $w=3.13e-07 $l=3.6e-07 $layer=LI1_cond $X=3.575 $Y=1.417
+ $X2=3.215 $Y2=1.417
r184 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.575
+ $Y=1.41 $X2=3.575 $Y2=1.41
r185 22 52 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.725 $Y=0.74
+ $X2=5.725 $Y2=1.22
r186 18 53 266.266 $w=1.8e-07 $l=6.85e-07 $layer=POLY_cond $X=5.63 $Y=2.235
+ $X2=5.63 $Y2=1.55
r187 14 48 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.61 $Y=2.235
+ $X2=3.61 $Y2=1.575
r188 10 47 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.595 $Y=0.74
+ $X2=3.595 $Y2=1.245
r189 6 45 266.266 $w=1.8e-07 $l=6.85e-07 $layer=POLY_cond $X=2.15 $Y=2.235
+ $X2=2.15 $Y2=1.55
r190 3 44 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.015 $Y=0.74
+ $X2=2.015 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__FA_4%A_418_74# 1 2 9 12 16 20 24 28 32 36 40 44 47
+ 49 51 52 53 54 58 62 65 66 67 69 70 71 73 74 79 84 86 87 89 90 95 96 97 100
+ 102 112
c294 102 0 2.53523e-19 $X=5.095 $Y=1.22
c295 97 0 2.88491e-20 $X=5.095 $Y=1.005
c296 47 0 2.59206e-19 $X=1.09 $Y=1.745
c297 12 0 2.03228e-19 $X=5.13 $Y=2.235
r298 112 113 8.89846 $w=3.25e-07 $l=6e-08 $layer=POLY_cond $X=10.485 $Y=1.485
+ $X2=10.545 $Y2=1.485
r299 111 112 54.8738 $w=3.25e-07 $l=3.7e-07 $layer=POLY_cond $X=10.115 $Y=1.485
+ $X2=10.485 $Y2=1.485
r300 110 111 11.8646 $w=3.25e-07 $l=8e-08 $layer=POLY_cond $X=10.035 $Y=1.485
+ $X2=10.115 $Y2=1.485
r301 107 108 22.2462 $w=3.25e-07 $l=1.5e-07 $layer=POLY_cond $X=9.535 $Y=1.485
+ $X2=9.685 $Y2=1.485
r302 106 107 41.5262 $w=3.25e-07 $l=2.8e-07 $layer=POLY_cond $X=9.255 $Y=1.485
+ $X2=9.535 $Y2=1.485
r303 100 103 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.095 $Y=1.385
+ $X2=5.095 $Y2=1.55
r304 100 102 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.095 $Y=1.385
+ $X2=5.095 $Y2=1.22
r305 99 100 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.095
+ $Y=1.385 $X2=5.095 $Y2=1.385
r306 97 99 14.1774 $w=3.27e-07 $l=3.8e-07 $layer=LI1_cond $X=5.095 $Y=1.005
+ $X2=5.095 $Y2=1.385
r307 95 96 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=3.385 $Y=0.965
+ $X2=3.555 $Y2=0.965
r308 90 93 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.375 $Y=2.375
+ $X2=2.375 $Y2=2.455
r309 86 87 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=1.665 $Y=0.965
+ $X2=1.835 $Y2=0.965
r310 82 84 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.09 $Y=1.83
+ $X2=1.41 $Y2=1.83
r311 80 110 28.92 $w=3.25e-07 $l=1.95e-07 $layer=POLY_cond $X=9.84 $Y=1.485
+ $X2=10.035 $Y2=1.485
r312 80 108 22.9877 $w=3.25e-07 $l=1.55e-07 $layer=POLY_cond $X=9.84 $Y=1.485
+ $X2=9.685 $Y2=1.485
r313 79 80 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=9.84
+ $Y=1.485 $X2=9.84 $Y2=1.485
r314 77 106 14.0892 $w=3.25e-07 $l=9.5e-08 $layer=POLY_cond $X=9.16 $Y=1.485
+ $X2=9.255 $Y2=1.485
r315 77 104 11.1231 $w=3.25e-07 $l=7.5e-08 $layer=POLY_cond $X=9.16 $Y=1.485
+ $X2=9.085 $Y2=1.485
r316 76 79 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=9.16 $Y=1.485
+ $X2=9.84 $Y2=1.485
r317 76 77 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=9.16
+ $Y=1.485 $X2=9.16 $Y2=1.485
r318 74 76 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=9.135 $Y=1.485
+ $X2=9.16 $Y2=1.485
r319 73 74 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.05 $Y=1.32
+ $X2=9.135 $Y2=1.485
r320 72 73 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=9.05 $Y=0.75
+ $X2=9.05 $Y2=1.32
r321 70 72 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.965 $Y=0.665
+ $X2=9.05 $Y2=0.75
r322 70 71 165.711 $w=1.68e-07 $l=2.54e-06 $layer=LI1_cond $X=8.965 $Y=0.665
+ $X2=6.425 $Y2=0.665
r323 69 71 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.34 $Y=0.58
+ $X2=6.425 $Y2=0.665
r324 68 69 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=6.34 $Y=0.425
+ $X2=6.34 $Y2=0.58
r325 66 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.255 $Y=0.34
+ $X2=6.34 $Y2=0.425
r326 66 67 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=6.255 $Y=0.34
+ $X2=5.255 $Y2=0.34
r327 65 97 5.97199 $w=3.27e-07 $l=1.16619e-07 $layer=LI1_cond $X=5.17 $Y=0.92
+ $X2=5.095 $Y2=1.005
r328 64 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.17 $Y=0.425
+ $X2=5.255 $Y2=0.34
r329 64 65 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.17 $Y=0.425
+ $X2=5.17 $Y2=0.92
r330 62 97 4.5696 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.93 $Y=1.005
+ $X2=5.095 $Y2=1.005
r331 62 96 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=4.93 $Y=1.005
+ $X2=3.555 $Y2=1.005
r332 61 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=0.925
+ $X2=2.3 $Y2=0.925
r333 61 95 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.465 $Y=0.925
+ $X2=3.385 $Y2=0.925
r334 56 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=0.84 $X2=2.3
+ $Y2=0.925
r335 56 58 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.3 $Y=0.84
+ $X2=2.3 $Y2=0.515
r336 54 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=0.925
+ $X2=2.3 $Y2=0.925
r337 54 87 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.135 $Y=0.925
+ $X2=1.835 $Y2=0.925
r338 52 90 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=2.375
+ $X2=2.375 $Y2=2.375
r339 52 53 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.21 $Y=2.375
+ $X2=1.495 $Y2=2.375
r340 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.41 $Y=2.29
+ $X2=1.495 $Y2=2.375
r341 50 84 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.41 $Y=1.915
+ $X2=1.41 $Y2=1.83
r342 50 51 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.41 $Y=1.915
+ $X2=1.41 $Y2=2.29
r343 49 86 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.175 $Y=1.005
+ $X2=1.665 $Y2=1.005
r344 47 82 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.09 $Y=1.745
+ $X2=1.09 $Y2=1.83
r345 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.09 $Y=1.09
+ $X2=1.175 $Y2=1.005
r346 46 47 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.09 $Y=1.09
+ $X2=1.09 $Y2=1.745
r347 42 113 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.545 $Y=1.32
+ $X2=10.545 $Y2=1.485
r348 42 44 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=10.545 $Y=1.32
+ $X2=10.545 $Y2=0.78
r349 38 112 16.5763 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.485 $Y=1.65
+ $X2=10.485 $Y2=1.485
r350 38 40 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=10.485 $Y=1.65
+ $X2=10.485 $Y2=2.4
r351 34 111 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.115 $Y=1.32
+ $X2=10.115 $Y2=1.485
r352 34 36 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=10.115 $Y=1.32
+ $X2=10.115 $Y2=0.78
r353 30 110 16.5763 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.035 $Y=1.65
+ $X2=10.035 $Y2=1.485
r354 30 32 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=10.035 $Y=1.65
+ $X2=10.035 $Y2=2.4
r355 26 108 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.685 $Y=1.32
+ $X2=9.685 $Y2=1.485
r356 26 28 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=9.685 $Y=1.32
+ $X2=9.685 $Y2=0.78
r357 22 107 16.5763 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.535 $Y=1.65
+ $X2=9.535 $Y2=1.485
r358 22 24 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=9.535 $Y=1.65
+ $X2=9.535 $Y2=2.4
r359 18 106 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.255 $Y=1.32
+ $X2=9.255 $Y2=1.485
r360 18 20 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=9.255 $Y=1.32
+ $X2=9.255 $Y2=0.78
r361 14 104 16.5763 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.085 $Y=1.65
+ $X2=9.085 $Y2=1.485
r362 14 16 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=9.085 $Y=1.65
+ $X2=9.085 $Y2=2.4
r363 12 103 266.266 $w=1.8e-07 $l=6.85e-07 $layer=POLY_cond $X=5.13 $Y=2.235
+ $X2=5.13 $Y2=1.55
r364 9 102 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.045 $Y=0.74
+ $X2=5.045 $Y2=1.22
r365 2 93 600 $w=1.7e-07 $l=7.84602e-07 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=1.735 $X2=2.375 $Y2=2.455
r366 1 89 182 $w=1.7e-07 $l=6.51594e-07 $layer=licon1_NDIFF $count=1 $X=2.09
+ $Y=0.37 $X2=2.3 $Y2=0.925
r367 1 58 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.09
+ $Y=0.37 $X2=2.3 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__FA_4%A 4 7 9 10 11 14 17 18 22 23 26 27 31 33 36 37
+ 38 39 40 42 43 50
c160 43 0 1.28731e-19 $X=0.72 $Y=1.665
c161 36 0 6.35672e-20 $X=6.64 $Y=2.34
c162 31 0 1.30844e-19 $X=6.625 $Y=0.74
c163 14 0 1.40726e-19 $X=3.11 $Y=2.235
c164 4 0 1.6759e-19 $X=0.505 $Y=2.46
r165 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.63
+ $Y=1.41 $X2=0.63 $Y2=1.41
r166 48 50 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=0.505 $Y=1.41
+ $X2=0.63 $Y2=1.41
r167 46 48 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.505 $Y2=1.41
r168 43 51 2.01209 $w=5.33e-07 $l=9e-08 $layer=LI1_cond $X=0.72 $Y=1.512
+ $X2=0.63 $Y2=1.512
r169 42 51 8.71908 $w=5.33e-07 $l=3.9e-07 $layer=LI1_cond $X=0.24 $Y=1.512
+ $X2=0.63 $Y2=1.512
r170 34 36 285.702 $w=1.8e-07 $l=7.35e-07 $layer=POLY_cond $X=6.64 $Y=3.075
+ $X2=6.64 $Y2=2.34
r171 33 41 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.64 $Y=1.705
+ $X2=6.64 $Y2=1.615
r172 33 36 246.831 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=6.64 $Y=1.705
+ $X2=6.64 $Y2=2.34
r173 31 41 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=6.625 $Y=0.74
+ $X2=6.625 $Y2=1.615
r174 28 40 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.72 $Y=3.15 $X2=4.63
+ $Y2=3.15
r175 27 34 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.55 $Y=3.15
+ $X2=6.64 $Y2=3.075
r176 27 28 938.362 $w=1.5e-07 $l=1.83e-06 $layer=POLY_cond $X=6.55 $Y=3.15
+ $X2=4.72 $Y2=3.15
r177 24 40 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.63 $Y=3.075
+ $X2=4.63 $Y2=3.15
r178 24 26 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=4.63 $Y=3.075
+ $X2=4.63 $Y2=2.235
r179 23 39 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.63 $Y=1.275
+ $X2=4.63 $Y2=1.185
r180 23 26 373.161 $w=1.8e-07 $l=9.6e-07 $layer=POLY_cond $X=4.63 $Y=1.275
+ $X2=4.63 $Y2=2.235
r181 22 39 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.615 $Y=0.74
+ $X2=4.615 $Y2=1.185
r182 19 38 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.2 $Y=3.15 $X2=3.11
+ $Y2=3.15
r183 18 40 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.54 $Y=3.15 $X2=4.63
+ $Y2=3.15
r184 18 19 687.106 $w=1.5e-07 $l=1.34e-06 $layer=POLY_cond $X=4.54 $Y=3.15
+ $X2=3.2 $Y2=3.15
r185 17 37 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.125 $Y=0.74
+ $X2=3.125 $Y2=1.185
r186 12 38 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.11 $Y=3.075
+ $X2=3.11 $Y2=3.15
r187 12 14 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=3.11 $Y=3.075
+ $X2=3.11 $Y2=2.235
r188 11 37 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=3.11 $Y=1.275
+ $X2=3.11 $Y2=1.185
r189 11 14 373.161 $w=1.8e-07 $l=9.6e-07 $layer=POLY_cond $X=3.11 $Y=1.275
+ $X2=3.11 $Y2=2.235
r190 9 38 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.02 $Y=3.15 $X2=3.11
+ $Y2=3.15
r191 9 10 1243.46 $w=1.5e-07 $l=2.425e-06 $layer=POLY_cond $X=3.02 $Y=3.15
+ $X2=0.595 $Y2=3.15
r192 5 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.245
+ $X2=0.495 $Y2=1.41
r193 5 7 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.495 $Y=1.245
+ $X2=0.495 $Y2=0.74
r194 2 10 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=0.505 $Y=3.075
+ $X2=0.595 $Y2=3.15
r195 2 4 239.056 $w=1.8e-07 $l=6.15e-07 $layer=POLY_cond $X=0.505 $Y=3.075
+ $X2=0.505 $Y2=2.46
r196 1 48 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.575
+ $X2=0.505 $Y2=1.41
r197 1 4 344.008 $w=1.8e-07 $l=8.85e-07 $layer=POLY_cond $X=0.505 $Y=1.575
+ $X2=0.505 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__FA_4%A_1024_74# 1 2 9 13 17 21 25 29 33 37 41 45 47
+ 50 52 58 62 64 68 69 70 74 83
c157 83 0 1.43637e-19 $X=8.585 $Y=1.505
c158 74 0 7.54566e-20 $X=6.99 $Y=1.505
c159 41 0 1.67591e-19 $X=6.255 $Y=2.145
r160 83 84 11.9752 $w=3.22e-07 $l=8e-08 $layer=POLY_cond $X=8.585 $Y=1.505
+ $X2=8.665 $Y2=1.505
r161 82 83 52.3913 $w=3.22e-07 $l=3.5e-07 $layer=POLY_cond $X=8.235 $Y=1.505
+ $X2=8.585 $Y2=1.505
r162 81 82 14.9689 $w=3.22e-07 $l=1e-07 $layer=POLY_cond $X=8.135 $Y=1.505
+ $X2=8.235 $Y2=1.505
r163 78 79 1.49689 $w=3.22e-07 $l=1e-08 $layer=POLY_cond $X=7.635 $Y=1.505
+ $X2=7.645 $Y2=1.505
r164 75 76 4.49068 $w=3.22e-07 $l=3e-08 $layer=POLY_cond $X=7.185 $Y=1.505
+ $X2=7.215 $Y2=1.505
r165 70 72 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.34 $Y=2.035
+ $X2=6.34 $Y2=2.145
r166 68 69 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=5.915 $Y=0.965
+ $X2=6.085 $Y2=0.965
r167 64 66 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=5.55 $Y=0.8
+ $X2=5.55 $Y2=0.925
r168 59 81 29.1894 $w=3.22e-07 $l=1.95e-07 $layer=POLY_cond $X=7.94 $Y=1.505
+ $X2=8.135 $Y2=1.505
r169 59 79 44.1584 $w=3.22e-07 $l=2.95e-07 $layer=POLY_cond $X=7.94 $Y=1.505
+ $X2=7.645 $Y2=1.505
r170 58 59 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.94
+ $Y=1.505 $X2=7.94 $Y2=1.505
r171 56 78 56.1335 $w=3.22e-07 $l=3.75e-07 $layer=POLY_cond $X=7.26 $Y=1.505
+ $X2=7.635 $Y2=1.505
r172 56 76 6.73602 $w=3.22e-07 $l=4.5e-08 $layer=POLY_cond $X=7.26 $Y=1.505
+ $X2=7.215 $Y2=1.505
r173 55 58 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.26 $Y=1.505
+ $X2=7.94 $Y2=1.505
r174 55 56 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.26
+ $Y=1.505 $X2=7.26 $Y2=1.505
r175 53 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.075 $Y=1.505
+ $X2=6.99 $Y2=1.505
r176 53 55 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=7.075 $Y=1.505
+ $X2=7.26 $Y2=1.505
r177 51 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.99 $Y=1.67
+ $X2=6.99 $Y2=1.505
r178 51 52 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=6.99 $Y=1.67
+ $X2=6.99 $Y2=1.95
r179 50 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.99 $Y=1.34
+ $X2=6.99 $Y2=1.505
r180 49 50 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.99 $Y=1.09
+ $X2=6.99 $Y2=1.34
r181 48 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.425 $Y=2.035
+ $X2=6.34 $Y2=2.035
r182 47 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.905 $Y=2.035
+ $X2=6.99 $Y2=1.95
r183 47 48 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=6.905 $Y=2.035
+ $X2=6.425 $Y2=2.035
r184 45 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.905 $Y=1.005
+ $X2=6.99 $Y2=1.09
r185 45 69 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=6.905 $Y=1.005
+ $X2=6.085 $Y2=1.005
r186 44 66 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.675 $Y=0.925
+ $X2=5.55 $Y2=0.925
r187 44 68 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.675 $Y=0.925
+ $X2=5.915 $Y2=0.925
r188 42 62 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.57 $Y=2.145
+ $X2=5.405 $Y2=2.145
r189 41 72 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.255 $Y=2.145
+ $X2=6.34 $Y2=2.145
r190 41 42 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=6.255 $Y=2.145
+ $X2=5.57 $Y2=2.145
r191 35 84 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.665 $Y=1.34
+ $X2=8.665 $Y2=1.505
r192 35 37 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.665 $Y=1.34
+ $X2=8.665 $Y2=0.78
r193 31 83 16.3606 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.585 $Y=1.67
+ $X2=8.585 $Y2=1.505
r194 31 33 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=8.585 $Y=1.67
+ $X2=8.585 $Y2=2.4
r195 27 82 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.235 $Y=1.34
+ $X2=8.235 $Y2=1.505
r196 27 29 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.235 $Y=1.34
+ $X2=8.235 $Y2=0.78
r197 23 81 16.3606 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.135 $Y=1.67
+ $X2=8.135 $Y2=1.505
r198 23 25 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=8.135 $Y=1.67
+ $X2=8.135 $Y2=2.4
r199 19 79 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.645 $Y=1.34
+ $X2=7.645 $Y2=1.505
r200 19 21 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.645 $Y=1.34
+ $X2=7.645 $Y2=0.78
r201 15 78 16.3606 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.635 $Y=1.67
+ $X2=7.635 $Y2=1.505
r202 15 17 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=7.635 $Y=1.67
+ $X2=7.635 $Y2=2.4
r203 11 76 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.215 $Y=1.34
+ $X2=7.215 $Y2=1.505
r204 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.215 $Y=1.34
+ $X2=7.215 $Y2=0.78
r205 7 75 16.3606 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.185 $Y=1.67
+ $X2=7.185 $Y2=1.505
r206 7 9 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=7.185 $Y=1.67
+ $X2=7.185 $Y2=2.4
r207 2 62 300 $w=1.7e-07 $l=4.93913e-07 $layer=licon1_PDIFF $count=2 $X=5.22
+ $Y=1.735 $X2=5.405 $Y2=2.145
r208 1 64 182 $w=1.7e-07 $l=5.93801e-07 $layer=licon1_NDIFF $count=1 $X=5.12
+ $Y=0.37 $X2=5.51 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_MS__FA_4%A_27_392# 1 2 7 9 11 14 15 19
r48 17 19 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=1.465 $Y=2.795
+ $X2=1.84 $Y2=2.795
r49 15 17 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.155 $Y=2.795
+ $X2=1.465 $Y2=2.795
r50 14 15 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.07 $Y=2.63
+ $X2=1.155 $Y2=2.795
r51 13 14 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.07 $Y=2.255
+ $X2=1.07 $Y2=2.63
r52 12 22 4.68787 $w=1.7e-07 $l=1.96074e-07 $layer=LI1_cond $X=0.445 $Y=2.17
+ $X2=0.28 $Y2=2.102
r53 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.985 $Y=2.17
+ $X2=1.07 $Y2=2.255
r54 11 12 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=0.985 $Y=2.17
+ $X2=0.445 $Y2=2.17
r55 7 22 3.0783 $w=3.3e-07 $l=1.53e-07 $layer=LI1_cond $X=0.28 $Y=2.255 $X2=0.28
+ $Y2=2.102
r56 7 9 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.28 $Y=2.255 $X2=0.28
+ $Y2=2.815
r57 2 19 600 $w=1.7e-07 $l=1.3245e-06 $layer=licon1_PDIFF $count=1 $X=1.245
+ $Y=1.735 $X2=1.84 $Y2=2.795
r58 2 17 600 $w=1.7e-07 $l=1.16482e-06 $layer=licon1_PDIFF $count=1 $X=1.245
+ $Y=1.735 $X2=1.465 $Y2=2.795
r59 1 22 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.115
r60 1 9 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__FA_4%VPWR 1 2 3 4 5 6 7 8 29 33 37 41 47 51 57 59 61
+ 66 67 68 77 81 86 91 96 101 107 110 113 116 119 122 126
c142 3 0 6.08971e-20 $X=4.15 $Y=1.735
c143 1 0 9.16158e-20 $X=0.595 $Y=1.96
r144 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r145 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r146 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r147 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r148 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r149 110 111 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r150 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r151 105 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r152 105 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r153 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r154 102 122 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.925 $Y=3.33
+ $X2=9.8 $Y2=3.33
r155 102 104 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=9.925 $Y=3.33
+ $X2=10.32 $Y2=3.33
r156 101 125 3.95357 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=10.625 $Y=3.33
+ $X2=10.832 $Y2=3.33
r157 101 104 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.625 $Y=3.33
+ $X2=10.32 $Y2=3.33
r158 100 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r159 100 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r160 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r161 97 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.975 $Y=3.33
+ $X2=8.85 $Y2=3.33
r162 97 99 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=8.975 $Y=3.33
+ $X2=9.36 $Y2=3.33
r163 96 122 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.675 $Y=3.33
+ $X2=9.8 $Y2=3.33
r164 96 99 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.675 $Y=3.33
+ $X2=9.36 $Y2=3.33
r165 95 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r166 95 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r167 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r168 92 116 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=7.9 $Y2=3.33
r169 92 94 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=8.4 $Y2=3.33
r170 91 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.725 $Y=3.33
+ $X2=8.85 $Y2=3.33
r171 91 94 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.725 $Y=3.33
+ $X2=8.4 $Y2=3.33
r172 90 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r173 90 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r174 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r175 87 113 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.045 $Y=3.33
+ $X2=6.92 $Y2=3.33
r176 87 89 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=7.045 $Y=3.33
+ $X2=7.44 $Y2=3.33
r177 86 116 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.775 $Y=3.33
+ $X2=7.9 $Y2=3.33
r178 86 89 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.775 $Y=3.33
+ $X2=7.44 $Y2=3.33
r179 85 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r180 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r181 82 110 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=4.57 $Y=3.33 $X2=4.37
+ $Y2=3.33
r182 82 84 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=4.57 $Y=3.33
+ $X2=6.48 $Y2=3.33
r183 81 113 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.795 $Y=3.33
+ $X2=6.92 $Y2=3.33
r184 81 84 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.795 $Y=3.33
+ $X2=6.48 $Y2=3.33
r185 80 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r186 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r187 77 110 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=4.17 $Y=3.33 $X2=4.37
+ $Y2=3.33
r188 77 79 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.17 $Y=3.33 $X2=4.08
+ $Y2=3.33
r189 76 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r190 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r191 73 76 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r192 73 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r193 72 75 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r194 72 73 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r195 70 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=0.73 $Y2=3.33
r196 70 72 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.815 $Y=3.33
+ $X2=1.2 $Y2=3.33
r197 68 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r198 68 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r199 66 75 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=3.17 $Y=3.33 $X2=3.12
+ $Y2=3.33
r200 66 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.17 $Y=3.33
+ $X2=3.335 $Y2=3.33
r201 65 79 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.5 $Y=3.33
+ $X2=4.08 $Y2=3.33
r202 65 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.5 $Y=3.33
+ $X2=3.335 $Y2=3.33
r203 61 64 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=10.75 $Y=1.985
+ $X2=10.75 $Y2=2.815
r204 59 125 3.18959 $w=2.5e-07 $l=1.19143e-07 $layer=LI1_cond $X=10.75 $Y=3.245
+ $X2=10.832 $Y2=3.33
r205 59 64 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.75 $Y=3.245
+ $X2=10.75 $Y2=2.815
r206 55 122 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.8 $Y=3.245
+ $X2=9.8 $Y2=3.33
r207 55 57 42.4099 $w=2.48e-07 $l=9.2e-07 $layer=LI1_cond $X=9.8 $Y=3.245
+ $X2=9.8 $Y2=2.325
r208 51 54 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=8.85 $Y=1.985
+ $X2=8.85 $Y2=2.815
r209 49 119 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.85 $Y=3.245
+ $X2=8.85 $Y2=3.33
r210 49 54 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.85 $Y=3.245
+ $X2=8.85 $Y2=2.815
r211 45 116 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=3.245
+ $X2=7.9 $Y2=3.33
r212 45 47 41.4879 $w=2.48e-07 $l=9e-07 $layer=LI1_cond $X=7.9 $Y=3.245 $X2=7.9
+ $Y2=2.345
r213 41 44 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=6.92 $Y=2.455
+ $X2=6.92 $Y2=2.815
r214 39 113 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.92 $Y=3.245
+ $X2=6.92 $Y2=3.33
r215 39 44 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6.92 $Y=3.245
+ $X2=6.92 $Y2=2.815
r216 35 110 1.46811 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.37 $Y=3.245
+ $X2=4.37 $Y2=3.33
r217 35 37 18.8713 $w=3.98e-07 $l=6.55e-07 $layer=LI1_cond $X=4.37 $Y=3.245
+ $X2=4.37 $Y2=2.59
r218 31 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=3.245
+ $X2=3.335 $Y2=3.33
r219 31 33 37.5417 $w=3.28e-07 $l=1.075e-06 $layer=LI1_cond $X=3.335 $Y=3.245
+ $X2=3.335 $Y2=2.17
r220 27 107 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r221 27 29 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.59
r222 8 64 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.575
+ $Y=1.84 $X2=10.71 $Y2=2.815
r223 8 61 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.575
+ $Y=1.84 $X2=10.71 $Y2=1.985
r224 7 57 300 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=2 $X=9.625
+ $Y=1.84 $X2=9.76 $Y2=2.325
r225 6 54 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.675
+ $Y=1.84 $X2=8.81 $Y2=2.815
r226 6 51 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.675
+ $Y=1.84 $X2=8.81 $Y2=1.985
r227 5 47 300 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_PDIFF $count=2 $X=7.725
+ $Y=1.84 $X2=7.86 $Y2=2.345
r228 4 44 600 $w=1.7e-07 $l=1.08392e-06 $layer=licon1_PDIFF $count=1 $X=6.73
+ $Y=1.84 $X2=6.96 $Y2=2.815
r229 4 41 600 $w=1.7e-07 $l=7.20885e-07 $layer=licon1_PDIFF $count=1 $X=6.73
+ $Y=1.84 $X2=6.96 $Y2=2.455
r230 3 37 600 $w=1.7e-07 $l=9.5871e-07 $layer=licon1_PDIFF $count=1 $X=4.15
+ $Y=1.735 $X2=4.37 $Y2=2.59
r231 2 33 300 $w=1.7e-07 $l=4.97946e-07 $layer=licon1_PDIFF $count=2 $X=3.2
+ $Y=1.735 $X2=3.335 $Y2=2.17
r232 1 29 600 $w=1.7e-07 $l=6.94226e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.96 $X2=0.73 $Y2=2.59
.ends

.subckt PM_SKY130_FD_SC_MS__FA_4%A_740_347# 1 2 9 11 13 16
c30 16 0 1.40726e-19 $X=3.835 $Y=2.17
c31 13 0 1.51516e-19 $X=4.905 $Y=2.59
r32 11 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.905 $Y=2.255
+ $X2=4.905 $Y2=2.17
r33 11 13 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.905 $Y=2.255
+ $X2=4.905 $Y2=2.59
r34 10 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4 $Y=2.17 $X2=3.835
+ $Y2=2.17
r35 9 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.74 $Y=2.17
+ $X2=4.905 $Y2=2.17
r36 9 10 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=4.74 $Y=2.17 $X2=4
+ $Y2=2.17
r37 2 18 600 $w=1.7e-07 $l=5.19326e-07 $layer=licon1_PDIFF $count=1 $X=4.72
+ $Y=1.735 $X2=4.905 $Y2=2.17
r38 2 13 600 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=4.72
+ $Y=1.735 $X2=4.905 $Y2=2.59
r39 1 16 300 $w=1.7e-07 $l=4.97946e-07 $layer=licon1_PDIFF $count=2 $X=3.7
+ $Y=1.735 $X2=3.835 $Y2=2.17
.ends

.subckt PM_SKY130_FD_SC_MS__FA_4%SUM 1 2 3 4 13 15 17 21 23 24 29 30 31 38
c61 17 0 1.30844e-19 $X=8.285 $Y=1.045
c62 13 0 6.35672e-20 $X=7.41 $Y=2.01
r63 36 38 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=8.36 $Y=2.01
+ $X2=8.36 $Y2=2.035
r64 30 31 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.36 $Y=2.405
+ $X2=8.36 $Y2=2.775
r65 29 36 3.29812 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=8.36 $Y=1.925
+ $X2=8.36 $Y2=2.01
r66 29 30 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.36 $Y=2.065
+ $X2=8.36 $Y2=2.405
r67 29 38 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=8.36 $Y=2.065 $X2=8.36
+ $Y2=2.035
r68 24 29 3.29812 $w=2.85e-07 $l=1.05119e-07 $layer=LI1_cond $X=8.405 $Y=1.84
+ $X2=8.36 $Y2=1.925
r69 23 28 3.46099 $w=2.4e-07 $l=1.45774e-07 $layer=LI1_cond $X=8.405 $Y=1.17
+ $X2=8.45 $Y2=1.045
r70 23 24 32.1724 $w=2.38e-07 $l=6.7e-07 $layer=LI1_cond $X=8.405 $Y=1.17
+ $X2=8.405 $Y2=1.84
r71 22 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.575 $Y=1.925
+ $X2=7.41 $Y2=1.925
r72 21 29 3.25423 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.195 $Y=1.925
+ $X2=8.36 $Y2=1.925
r73 21 22 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=8.195 $Y=1.925
+ $X2=7.575 $Y2=1.925
r74 17 28 3.3592 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=8.285 $Y=1.045
+ $X2=8.45 $Y2=1.045
r75 17 19 39.4136 $w=2.48e-07 $l=8.55e-07 $layer=LI1_cond $X=8.285 $Y=1.045
+ $X2=7.43 $Y2=1.045
r76 13 26 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.41 $Y=2.01 $X2=7.41
+ $Y2=1.925
r77 13 15 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=7.41 $Y=2.01
+ $X2=7.41 $Y2=2.815
r78 4 29 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=8.225
+ $Y=1.84 $X2=8.36 $Y2=2.005
r79 4 31 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.225
+ $Y=1.84 $X2=8.36 $Y2=2.815
r80 3 26 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=7.275
+ $Y=1.84 $X2=7.41 $Y2=2.005
r81 3 15 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.275
+ $Y=1.84 $X2=7.41 $Y2=2.815
r82 2 28 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=8.31
+ $Y=0.41 $X2=8.45 $Y2=1.005
r83 1 19 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=7.29
+ $Y=0.41 $X2=7.43 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_MS__FA_4%COUT 1 2 3 4 13 15 19 21 23 24 27 30 33 34 35
+ 36 37 43 45
c69 43 0 9.5881e-20 $X=10.265 $Y=1.99
r70 43 45 1.52529 $w=3.38e-07 $l=4.5e-08 $layer=LI1_cond $X=10.265 $Y=1.99
+ $X2=10.265 $Y2=2.035
r71 36 37 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=10.265 $Y=2.405
+ $X2=10.265 $Y2=2.775
r72 35 43 0.944793 $w=3.4e-07 $l=2e-08 $layer=LI1_cond $X=10.265 $Y=1.97
+ $X2=10.265 $Y2=1.99
r73 35 55 2.67003 $w=2.97e-07 $l=6.5e-08 $layer=LI1_cond $X=10.265 $Y=1.97
+ $X2=10.265 $Y2=1.905
r74 35 36 11.8634 $w=3.38e-07 $l=3.5e-07 $layer=LI1_cond $X=10.265 $Y=2.055
+ $X2=10.265 $Y2=2.405
r75 35 45 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=10.265 $Y=2.055
+ $X2=10.265 $Y2=2.035
r76 34 55 9.85859 $w=2.97e-07 $l=2.4e-07 $layer=LI1_cond $X=10.265 $Y=1.665
+ $X2=10.265 $Y2=1.905
r77 30 34 4.94494 $w=2.97e-07 $l=1.29132e-07 $layer=LI1_cond $X=10.295 $Y=1.55
+ $X2=10.265 $Y2=1.665
r78 29 33 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=10.295 $Y=1.15
+ $X2=10.295 $Y2=1.065
r79 29 30 17.7299 $w=2.58e-07 $l=4e-07 $layer=LI1_cond $X=10.295 $Y=1.15
+ $X2=10.295 $Y2=1.55
r80 25 33 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=10.295 $Y=0.98
+ $X2=10.295 $Y2=1.065
r81 25 27 18.838 $w=2.58e-07 $l=4.25e-07 $layer=LI1_cond $X=10.295 $Y=0.98
+ $X2=10.295 $Y2=0.555
r82 23 33 2.90867 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.165 $Y=1.065
+ $X2=10.295 $Y2=1.065
r83 23 24 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=10.165 $Y=1.065
+ $X2=9.555 $Y2=1.065
r84 22 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.475 $Y=1.905
+ $X2=9.31 $Y2=1.905
r85 21 55 4.00195 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=10.095 $Y=1.905
+ $X2=10.265 $Y2=1.905
r86 21 22 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=10.095 $Y=1.905
+ $X2=9.475 $Y2=1.905
r87 17 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.43 $Y=0.98
+ $X2=9.555 $Y2=1.065
r88 17 19 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=9.43 $Y=0.98
+ $X2=9.43 $Y2=0.555
r89 13 32 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.31 $Y=1.99 $X2=9.31
+ $Y2=1.905
r90 13 15 28.8111 $w=3.28e-07 $l=8.25e-07 $layer=LI1_cond $X=9.31 $Y=1.99
+ $X2=9.31 $Y2=2.815
r91 4 35 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.125
+ $Y=1.84 $X2=10.26 $Y2=1.985
r92 4 37 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.125
+ $Y=1.84 $X2=10.26 $Y2=2.815
r93 3 32 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.175
+ $Y=1.84 $X2=9.31 $Y2=1.985
r94 3 15 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.175
+ $Y=1.84 $X2=9.31 $Y2=2.815
r95 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.19
+ $Y=0.41 $X2=10.33 $Y2=0.555
r96 1 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.33
+ $Y=0.41 $X2=9.47 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_MS__FA_4%A_27_74# 1 2 11 14 18 19
r32 18 19 8.64032 $w=3.18e-07 $l=1.7e-07 $layer=LI1_cond $X=1.325 $Y=0.55
+ $X2=1.495 $Y2=0.55
r33 14 16 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.28 $Y=0.515
+ $X2=0.28 $Y2=0.665
r34 11 19 10.9842 $w=3.18e-07 $l=3.05e-07 $layer=LI1_cond $X=1.8 $Y=0.51
+ $X2=1.495 $Y2=0.51
r35 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=0.665
+ $X2=0.28 $Y2=0.665
r36 8 18 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=0.445 $Y=0.665
+ $X2=1.325 $Y2=0.665
r37 2 11 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1.66 $Y=0.37
+ $X2=1.8 $Y2=0.55
r38 1 14 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__FA_4%VGND 1 2 3 4 5 6 7 8 27 31 33 35 38 39 40 41 47
+ 64 71 76 81 86 94 97 100 107 114 120 124
r146 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r147 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r148 114 117 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=8.96 $Y=0
+ $X2=8.96 $Y2=0.325
r149 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r150 107 110 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=7.94 $Y=0
+ $X2=7.94 $Y2=0.325
r151 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r152 100 103 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=6.92 $Y=0
+ $X2=6.92 $Y2=0.325
r153 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r154 96 97 11.9029 $w=4.93e-07 $l=2.65e-07 $layer=LI1_cond $X=0.89 $Y=0.162
+ $X2=1.155 $Y2=0.162
r155 92 96 4.10774 $w=4.93e-07 $l=1.7e-07 $layer=LI1_cond $X=0.72 $Y=0.162
+ $X2=0.89 $Y2=0.162
r156 92 94 7.79514 $w=4.93e-07 $l=9.5e-08 $layer=LI1_cond $X=0.72 $Y=0.162
+ $X2=0.625 $Y2=0.162
r157 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r158 90 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r159 90 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r160 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r161 87 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.985 $Y=0
+ $X2=9.86 $Y2=0
r162 87 89 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.985 $Y=0
+ $X2=10.32 $Y2=0
r163 86 123 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=10.595 $Y=0
+ $X2=10.817 $Y2=0
r164 86 89 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.595 $Y=0
+ $X2=10.32 $Y2=0
r165 85 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r166 85 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r167 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r168 82 114 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.125 $Y=0
+ $X2=8.96 $Y2=0
r169 82 84 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.125 $Y=0
+ $X2=9.36 $Y2=0
r170 81 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.735 $Y=0
+ $X2=9.86 $Y2=0
r171 81 84 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=9.735 $Y=0
+ $X2=9.36 $Y2=0
r172 80 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r173 80 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r174 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r175 77 107 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.105 $Y=0
+ $X2=7.94 $Y2=0
r176 77 79 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.105 $Y=0 $X2=8.4
+ $Y2=0
r177 76 114 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.795 $Y=0
+ $X2=8.96 $Y2=0
r178 76 79 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=8.795 $Y=0 $X2=8.4
+ $Y2=0
r179 75 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r180 75 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.96 $Y2=0
r181 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r182 72 100 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.085 $Y=0
+ $X2=6.92 $Y2=0
r183 72 74 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.085 $Y=0
+ $X2=7.44 $Y2=0
r184 71 107 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.775 $Y=0
+ $X2=7.94 $Y2=0
r185 71 74 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.775 $Y=0
+ $X2=7.44 $Y2=0
r186 70 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r187 69 70 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r188 66 69 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6.48
+ $Y2=0
r189 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r190 64 100 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.755 $Y=0
+ $X2=6.92 $Y2=0
r191 64 69 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=0
+ $X2=6.48 $Y2=0
r192 63 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r193 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r194 60 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r195 59 60 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r196 57 60 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r197 57 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r198 56 59 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r199 56 97 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.155
+ $Y2=0
r200 56 57 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r201 52 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r202 51 94 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.24 $Y=0
+ $X2=0.625 $Y2=0
r203 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r204 47 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r205 47 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r206 43 66 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.485 $Y=0 $X2=4.56
+ $Y2=0
r207 41 62 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.155 $Y=0 $X2=4.08
+ $Y2=0
r208 40 45 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.32 $Y=0 $X2=4.32
+ $Y2=0.325
r209 40 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=0 $X2=4.485
+ $Y2=0
r210 40 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.32 $Y=0 $X2=4.155
+ $Y2=0
r211 38 59 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.175 $Y=0 $X2=3.12
+ $Y2=0
r212 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.175 $Y=0 $X2=3.34
+ $Y2=0
r213 37 62 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=3.505 $Y=0
+ $X2=4.08 $Y2=0
r214 37 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.505 $Y=0 $X2=3.34
+ $Y2=0
r215 33 123 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.76 $Y=0.085
+ $X2=10.817 $Y2=0
r216 33 35 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=10.76 $Y=0.085
+ $X2=10.76 $Y2=0.555
r217 29 120 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.86 $Y=0.085
+ $X2=9.86 $Y2=0
r218 29 31 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=9.86 $Y=0.085
+ $X2=9.86 $Y2=0.645
r219 25 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.34 $Y=0.085
+ $X2=3.34 $Y2=0
r220 25 27 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.34 $Y=0.085
+ $X2=3.34 $Y2=0.55
r221 8 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.62
+ $Y=0.41 $X2=10.76 $Y2=0.555
r222 7 31 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=9.76
+ $Y=0.41 $X2=9.9 $Y2=0.645
r223 6 117 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=8.74
+ $Y=0.41 $X2=8.96 $Y2=0.325
r224 5 110 182 $w=1.7e-07 $l=2.59037e-07 $layer=licon1_NDIFF $count=1 $X=7.72
+ $Y=0.41 $X2=7.94 $Y2=0.325
r225 4 103 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=6.7
+ $Y=0.37 $X2=6.92 $Y2=0.325
r226 3 45 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=4.1
+ $Y=0.37 $X2=4.32 $Y2=0.325
r227 2 27 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.2 $Y=0.37
+ $X2=3.34 $Y2=0.55
r228 1 96 182 $w=1.7e-07 $l=3.4176e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.89 $Y2=0.325
.ends

.subckt PM_SKY130_FD_SC_MS__FA_4%A_734_74# 1 2 7 10 15
c26 15 0 1.62604e-19 $X=4.83 $Y=0.55
c27 10 0 1.78103e-19 $X=3.81 $Y=0.55
r28 15 17 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=4.79 $Y=0.55
+ $X2=4.79 $Y2=0.665
r29 10 12 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=3.85 $Y=0.55
+ $X2=3.85 $Y2=0.665
r30 8 12 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.975 $Y=0.665
+ $X2=3.85 $Y2=0.665
r31 7 17 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.665 $Y=0.665
+ $X2=4.79 $Y2=0.665
r32 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.665 $Y=0.665
+ $X2=3.975 $Y2=0.665
r33 2 15 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=4.69 $Y=0.37
+ $X2=4.83 $Y2=0.55
r34 1 10 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=3.67 $Y=0.37
+ $X2=3.81 $Y2=0.55
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfrtp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
M1000 a_1234_119# a_1037_387# a_303_464# VPB pshort w=420000u l=180000u
+  ad=2.576e+11p pd=2.93e+06u as=9.24e+11p ps=6.48e+06u
M1001 a_1320_119# a_1037_387# a_1234_119# VNB nlowvt w=420000u l=150000u
+  ad=9.87e+10p pd=1.31e+06u as=1.176e+11p ps=1.4e+06u
M1002 a_219_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=2.08418e+12p ps=1.846e+07u
M1003 VGND a_1997_272# a_1972_74# VNB nlowvt w=420000u l=150000u
+  ad=1.60052e+12p pd=1.375e+07u as=8.82e+10p ps=1.26e+06u
M1004 a_1972_74# a_835_93# a_1745_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=4.687e+11p ps=3.25e+06u
M1005 VPWR SCE a_27_88# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1006 a_1745_74# a_1037_387# a_1367_93# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1007 Q a_2402_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1008 a_312_81# a_27_88# a_225_81# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.499e+11p ps=2.87e+06u
M1009 a_303_464# D a_312_81# VNB nlowvt w=420000u l=150000u
+  ad=3.738e+11p pd=3.46e+06u as=0p ps=0u
M1010 a_1234_119# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Q a_2402_424# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1012 VGND RESET_B a_1397_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1013 a_303_464# D a_219_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1996_508# a_1037_387# a_1745_74# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=4.21675e+11p ps=3.58e+06u
M1015 a_225_81# SCD a_545_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1016 a_535_464# a_27_88# a_303_464# VPB pshort w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1017 a_1346_461# a_835_93# a_1234_119# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1018 VPWR CLK a_835_93# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1019 VPWR SCD a_535_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1397_119# a_1367_93# a_1320_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1997_272# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1022 a_1997_272# a_1745_74# a_2135_74# VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1023 a_303_464# RESET_B VPWR VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_1745_74# a_1997_272# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_545_81# SCE a_303_464# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1367_93# a_1234_119# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1027 a_2402_424# a_1745_74# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=0p ps=0u
M1028 VPWR a_1367_93# a_1346_461# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND CLK a_835_93# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.8265e+11p ps=2.43e+06u
M1030 a_1037_387# a_835_93# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1031 a_1745_74# a_835_93# a_1367_93# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1037_387# a_835_93# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.961e+11p pd=2.01e+06u as=0p ps=0u
M1033 a_1367_93# a_1234_119# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND SCE a_27_88# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1035 a_1234_119# a_835_93# a_303_464# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND RESET_B a_225_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR a_1997_272# a_1996_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_2135_74# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_2402_424# a_1745_74# VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
.ends

* File: sky130_fd_sc_ms__einvp_1.spice
* Created: Fri Aug 28 17:33:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__einvp_1.pex.spice"
.subckt sky130_fd_sc_ms__einvp_1  VNB VPB TE A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE	TE
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_TE_M1003_g N_A_44_549#_M1003_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0824069 AS=0.2604 PD=0.782069 PS=2.08 NRD=17.136 NRS=0 M=1 R=2.8
+ SA=75000.5 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 A_318_74# N_TE_M1001_g N_VGND_M1003_d VNB NLOWVT L=0.15 W=0.74 AD=0.0888
+ AS=0.145193 PD=0.98 PS=1.37793 NRD=10.536 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1002 N_Z_M1002_d N_A_M1002_g A_318_74# VNB NLOWVT L=0.15 W=0.74 AD=0.2109
+ AS=0.0888 PD=2.05 PS=0.98 NRD=0 NRS=10.536 M=1 R=4.93333 SA=75001.1 SB=75000.2
+ A=0.111 P=1.78 MULT=1
MM1005 N_VPWR_M1005_d N_TE_M1005_g N_A_44_549#_M1005_s VPB PSHORT L=0.18 W=0.42
+ AD=0.0921338 AS=0.2583 PD=0.801549 PS=2.07 NRD=37.5088 NRS=0 M=1 R=2.33333
+ SA=90000.5 SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1000 A_313_392# N_A_44_549#_M1000_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.219366 PD=1.24 PS=1.90845 NRD=12.7853 NRS=0 M=1 R=5.55556
+ SA=90000.6 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1004 N_Z_M1004_d N_A_M1004_g A_313_392# VPB PSHORT L=0.18 W=1 AD=0.28 AS=0.12
+ PD=2.56 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556 SA=90001 SB=90000.2 A=0.18
+ P=2.36 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1708 P=9.28
c_23 VNB 0 1.4658e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__einvp_1.pxi.spice"
*
.ends
*
*

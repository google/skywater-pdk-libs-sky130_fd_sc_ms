* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 X a_209_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 VPWR a_209_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X2 VGND A1 a_27_136# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 a_27_136# A1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 a_209_392# B2 a_27_136# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 VGND A2 a_27_136# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 VGND a_209_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VPWR a_209_392# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 a_519_392# B2 a_209_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X9 a_209_392# B1 a_27_136# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X10 a_27_136# B2 a_209_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X11 a_119_392# A2 a_209_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X12 a_27_136# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 a_209_392# B2 a_519_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X14 X a_209_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X15 X a_209_392# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X16 X a_209_392# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 a_209_392# A2 a_119_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X18 a_519_392# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X19 VGND a_209_392# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 VPWR B1 a_519_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X21 VPWR A1 a_119_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X22 a_27_136# B1 a_209_392# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X23 a_119_392# A1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
.ends

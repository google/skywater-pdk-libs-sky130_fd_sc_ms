* File: sky130_fd_sc_ms__nor2b_4.spice
* Created: Wed Sep  2 12:15:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nor2b_4.pex.spice"
.subckt sky130_fd_sc_ms__nor2b_4  VNB VPB A B_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B_N	B_N
* A	A
* VPB	VPB
* VNB	VNB
MM1006 N_Y_M1006_d N_A_353_323#_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.3223 PD=1.02 PS=2.57 NRD=0 NRS=61.704 M=1 R=4.93333 SA=75000.3
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1014 N_Y_M1006_d N_A_353_323#_M1014_g N_VGND_M1014_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.4097 PD=1.02 PS=1.84 NRD=0 NRS=80.856 M=1 R=4.93333 SA=75000.7
+ SB=75002.6 A=0.111 P=1.78 MULT=1
MM1003 N_Y_M1003_d N_A_M1003_g N_VGND_M1014_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.4097 PD=1.02 PS=1.84 NRD=0 NRS=80.856 M=1 R=4.93333 SA=75001.8 SB=75001.5
+ A=0.111 P=1.78 MULT=1
MM1008 N_Y_M1003_d N_A_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.2 SB=75001.1
+ A=0.111 P=1.78 MULT=1
MM1001 N_A_353_323#_M1001_d N_B_N_M1001_g N_VGND_M1008_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.518 AS=0.1036 PD=2.88 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1004 N_A_119_368#_M1004_d N_A_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90004.2 A=0.2016 P=2.6 MULT=1
MM1005 N_A_119_368#_M1004_d N_A_M1005_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90003.7 A=0.2016 P=2.6 MULT=1
MM1007 N_A_119_368#_M1007_d N_A_M1007_g N_VPWR_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90003.3 A=0.2016 P=2.6 MULT=1
MM1009 N_Y_M1009_d N_A_353_323#_M1009_g N_A_119_368#_M1007_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.5 SB=90002.8 A=0.2016 P=2.6 MULT=1
MM1010 N_Y_M1009_d N_A_353_323#_M1010_g N_A_119_368#_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1011 N_Y_M1011_d N_A_353_323#_M1011_g N_A_119_368#_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90002.4 SB=90001.9 A=0.2016 P=2.6 MULT=1
MM1013 N_Y_M1011_d N_A_353_323#_M1013_g N_A_119_368#_M1013_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90002.9 SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1012 N_A_119_368#_M1013_s N_A_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.2472 PD=1.44 PS=1.74286 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90003.4 SB=90001 A=0.2016 P=2.6 MULT=1
MM1000 N_A_353_323#_M1000_d N_B_N_M1000_g N_VPWR_M1012_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1134 AS=0.1854 PD=1.11 PS=1.30714 NRD=0 NRS=19.1484 M=1 R=4.66667
+ SA=90004 SB=90000.6 A=0.1512 P=2.04 MULT=1
MM1002 N_A_353_323#_M1000_d N_B_N_M1002_g N_VPWR_M1002_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1134 AS=0.2352 PD=1.11 PS=2.24 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90004.4 SB=90000.2 A=0.1512 P=2.04 MULT=1
DX15_noxref VNB VPB NWDIODE A=10.5276 P=15.04
*
.include "sky130_fd_sc_ms__nor2b_4.pxi.spice"
*
.ends
*
*

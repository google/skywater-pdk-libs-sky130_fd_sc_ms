* File: sky130_fd_sc_ms__dfrtp_2.spice
* Created: Wed Sep  2 12:03:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dfrtp_2.pex.spice"
.subckt sky130_fd_sc_ms__dfrtp_2  VNB VPB D CLK RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* CLK	CLK
* D	D
* VPB	VPB
* VNB	VNB
MM1028 A_117_78# N_D_M1028_g N_A_30_78#_M1028_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_RESET_B_M1012_g A_117_78# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_CLK_M1016_g N_A_306_119#_M1016_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1554 AS=0.2109 PD=1.16 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1013 N_A_493_387#_M1013_d N_A_306_119#_M1013_g N_VGND_M1016_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.198825 AS=0.1554 PD=2.05 PS=1.16 NRD=0 NRS=11.34 M=1
+ R=4.93333 SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1026 N_A_699_463#_M1026_d N_A_306_119#_M1026_g N_A_30_78#_M1026_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.7 A=0.063 P=1.14 MULT=1
MM1024 A_817_138# N_A_493_387#_M1024_g N_A_699_463#_M1026_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1008 A_895_138# N_A_837_359#_M1008_g A_817_138# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_RESET_B_M1001_g A_895_138# VNB NLOWVT L=0.15 W=0.42
+ AD=0.255829 AS=0.0504 PD=1.33241 PS=0.66 NRD=158.316 NRS=18.564 M=1 R=2.8
+ SA=75001.5 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1023 N_A_837_359#_M1023_d N_A_699_463#_M1023_g N_VGND_M1001_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.12025 AS=0.450746 PD=1.065 PS=2.34759 NRD=0 NRS=89.856 M=1
+ R=4.93333 SA=75001.7 SB=75002 A=0.111 P=1.78 MULT=1
MM1003 N_A_1271_74#_M1003_d N_A_493_387#_M1003_g N_A_837_359#_M1023_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.292172 AS=0.12025 PD=2.09241 PS=1.065 NRD=4.044 NRS=7.296
+ M=1 R=4.93333 SA=75002.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1032 A_1481_81# N_A_306_119#_M1032_g N_A_1271_74#_M1003_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.165828 PD=0.66 PS=1.18759 NRD=18.564 NRS=47.136 M=1
+ R=2.8 SA=75002.8 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_1525_212#_M1005_g A_1481_81# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0777 AS=0.0504 PD=0.79 PS=0.66 NRD=12.852 NRS=18.564 M=1 R=2.8 SA=75003.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1021 A_1663_81# N_RESET_B_M1021_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0777 PD=0.66 PS=0.79 NRD=18.564 NRS=12.852 M=1 R=2.8 SA=75003.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1022 N_A_1525_212#_M1022_d N_A_1271_74#_M1022_g A_1663_81# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1176 AS=0.0504 PD=1.4 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75004.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1020 N_A_1924_409#_M1020_d N_A_1271_74#_M1020_g N_VGND_M1020_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.2072 PD=2.05 PS=2.04 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1031 N_Q_M1031_d N_A_1924_409#_M1031_g N_VGND_M1031_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1033 N_Q_M1031_d N_A_1924_409#_M1033_g N_VGND_M1033_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2072 PD=1.02 PS=2.04 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1014 N_A_30_78#_M1014_d N_D_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=0.42
+ AD=0.0567 AS=0.1134 PD=0.69 PS=1.38 NRD=0 NRS=0 M=1 R=2.33333 SA=90000.2
+ SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1015 N_VPWR_M1015_d N_RESET_B_M1015_g N_A_30_78#_M1014_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1113 AS=0.0567 PD=1.37 PS=0.69 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1025 N_VPWR_M1025_d N_CLK_M1025_g N_A_306_119#_M1025_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2968 PD=1.39 PS=2.77 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1027 N_A_493_387#_M1027_d N_A_306_119#_M1027_g N_VPWR_M1025_d VPB PSHORT
+ L=0.18 W=1.12 AD=0.2968 AS=0.1512 PD=2.77 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1004 N_A_699_463#_M1004_d N_A_493_387#_M1004_g N_A_30_78#_M1004_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0567 AS=0.1155 PD=0.69 PS=1.39 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90001.7 A=0.0756 P=1.2 MULT=1
MM1006 A_789_463# N_A_306_119#_M1006_g N_A_699_463#_M1004_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0567 PD=0.66 PS=0.69 NRD=30.4759 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1011 N_VPWR_M1011_d N_A_837_359#_M1011_g A_789_463# VPB PSHORT L=0.18 W=0.42
+ AD=0.12865 AS=0.0504 PD=1.11 PS=0.66 NRD=39.8531 NRS=30.4759 M=1 R=2.33333
+ SA=90001.1 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1017 N_A_699_463#_M1017_d N_RESET_B_M1017_g N_VPWR_M1011_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1176 AS=0.12865 PD=1.4 PS=1.11 NRD=0 NRS=117.865 M=1 R=2.33333
+ SA=90001.7 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1000 N_A_837_359#_M1000_d N_A_699_463#_M1000_g N_VPWR_M1000_s VPB PSHORT
+ L=0.18 W=1 AD=0.169062 AS=0.28 PD=1.4 PS=2.56 NRD=8.8453 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1007 N_A_1271_74#_M1007_d N_A_306_119#_M1007_g N_A_837_359#_M1000_d VPB PSHORT
+ L=0.18 W=1 AD=0.304665 AS=0.169062 PD=2.53521 PS=1.4 NRD=7.8603 NRS=0 M=1
+ R=5.55556 SA=90000.7 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1009 A_1481_493# N_A_493_387#_M1009_g N_A_1271_74#_M1007_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.12796 PD=0.66 PS=1.06479 NRD=30.4759 NRS=0 M=1 R=2.33333
+ SA=90001.2 SB=90002.4 A=0.0756 P=1.2 MULT=1
MM1018 N_VPWR_M1018_d N_A_1525_212#_M1018_g A_1481_493# VPB PSHORT L=0.18 W=0.42
+ AD=0.0672 AS=0.0504 PD=0.74 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.33333 SA=90001.7
+ SB=90002 A=0.0756 P=1.2 MULT=1
MM1019 N_A_1525_212#_M1019_d N_RESET_B_M1019_g N_VPWR_M1018_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1113 AS=0.0672 PD=0.95 PS=0.74 NRD=58.6272 NRS=21.0987 M=1
+ R=2.33333 SA=90002.2 SB=90001.5 A=0.0756 P=1.2 MULT=1
MM1002 N_VPWR_M1002_d N_A_1271_74#_M1002_g N_A_1525_212#_M1019_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.1029 AS=0.1113 PD=0.83 PS=0.95 NRD=37.5088 NRS=58.6272 M=1
+ R=2.33333 SA=90002.9 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1010 N_A_1924_409#_M1010_d N_A_1271_74#_M1010_g N_VPWR_M1002_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2352 AS=0.2058 PD=2.24 PS=1.66 NRD=0 NRS=10.5395 M=1
+ R=4.66667 SA=90001.9 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1029 N_Q_M1029_d N_A_1924_409#_M1029_g N_VPWR_M1029_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3416 PD=1.39 PS=2.85 NRD=0 NRS=3.5066 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1030 N_Q_M1029_d N_A_1924_409#_M1030_g N_VPWR_M1030_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.7
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX34_noxref VNB VPB NWDIODE A=22.5036 P=27.76
c_117 VNB 0 8.65509e-20 $X=0 $Y=0
c_241 VPB 0 1.21261e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__dfrtp_2.pxi.spice"
*
.ends
*
*

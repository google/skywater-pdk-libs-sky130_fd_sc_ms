* File: sky130_fd_sc_ms__a41o_4.spice
* Created: Fri Aug 28 17:09:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a41o_4.pex.spice"
.subckt sky130_fd_sc_ms__a41o_4  VNB VPB B1 A1 A2 A3 A4 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1006 N_A_113_98#_M1006_d N_B1_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2072 PD=1.02 PS=2.04 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75002.7 A=0.111 P=1.78 MULT=1
MM1019 N_A_113_98#_M1006_d N_B1_M1019_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1955 PD=1.02 PS=1.43 NRD=0 NRS=33.912 M=1 R=4.93333 SA=75000.6
+ SB=75002.3 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1019_s N_A_113_98#_M1001_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1955 AS=0.1036 PD=1.43 PS=1.02 NRD=33.912 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75001.7 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1004_d N_A_113_98#_M1004_g N_X_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.193 AS=0.1036 PD=1.425 PS=1.02 NRD=33.372 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75001.3 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1004_d N_A_113_98#_M1017_g N_X_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.193 AS=0.1036 PD=1.425 PS=1.02 NRD=33.372 NRS=0 M=1 R=4.93333 SA=75002.2
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1023 N_VGND_M1023_d N_A_113_98#_M1023_g N_X_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.3495 AS=0.1036 PD=2.81 PS=1.02 NRD=67.668 NRS=0 M=1 R=4.93333 SA=75002.6
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1012 N_A_113_98#_M1012_d N_A1_M1012_g N_A_751_74#_M1012_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1013 N_A_113_98#_M1012_d N_A1_M1013_g N_A_751_74#_M1013_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1005 N_A_751_74#_M1013_s N_A2_M1005_g N_A_1010_74#_M1005_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1026 N_A_751_74#_M1026_d N_A2_M1026_g N_A_1010_74#_M1005_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2035 AS=0.1036 PD=2.03 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_A_1205_74#_M1003_d N_A3_M1003_g N_A_1010_74#_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2072 AS=0.1036 PD=2.04 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.5 A=0.111 P=1.78 MULT=1
MM1020 N_A_1205_74#_M1020_d N_A3_M1020_g N_A_1010_74#_M1003_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1002 N_A_1205_74#_M1020_d N_A4_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1015 N_A_1205_74#_M1015_d N_A4_M1015_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2072 AS=0.1036 PD=2.04 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_A_113_98#_M1000_d N_B1_M1000_g N_A_27_392#_M1000_s VPB PSHORT L=0.18
+ W=1 AD=0.16 AS=0.28 PD=1.32 PS=2.56 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1027 N_A_113_98#_M1000_d N_B1_M1027_g N_A_27_392#_M1027_s VPB PSHORT L=0.18
+ W=1 AD=0.16 AS=0.28 PD=1.32 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1021 N_X_M1021_d N_A_113_98#_M1021_g N_VPWR_M1021_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90005.4 A=0.2016 P=2.6 MULT=1
MM1022 N_X_M1021_d N_A_113_98#_M1022_g N_VPWR_M1022_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90004.9 A=0.2016 P=2.6 MULT=1
MM1024 N_X_M1024_d N_A_113_98#_M1024_g N_VPWR_M1022_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90004.5 A=0.2016 P=2.6 MULT=1
MM1025 N_X_M1024_d N_A_113_98#_M1025_g N_VPWR_M1025_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.195472 PD=1.39 PS=1.54264 NRD=0 NRS=0.8668 M=1 R=6.22222
+ SA=90001.5 SB=90004 A=0.2016 P=2.6 MULT=1
MM1016 N_VPWR_M1025_s N_A1_M1016_g N_A_27_392#_M1016_s VPB PSHORT L=0.18 W=1
+ AD=0.174528 AS=0.2325 PD=1.37736 PS=1.465 NRD=10.8153 NRS=18.715 M=1 R=5.55556
+ SA=90002.1 SB=90004 A=0.18 P=2.36 MULT=1
MM1018 N_VPWR_M1018_d N_A1_M1018_g N_A_27_392#_M1016_s VPB PSHORT L=0.18 W=1
+ AD=0.2475 AS=0.2325 PD=1.495 PS=1.465 NRD=20.685 NRS=17.73 M=1 R=5.55556
+ SA=90002.7 SB=90003.3 A=0.18 P=2.36 MULT=1
MM1011 N_A_27_392#_M1011_d N_A2_M1011_g N_VPWR_M1018_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.2475 PD=1.27 PS=1.495 NRD=0 NRS=21.67 M=1 R=5.55556 SA=90003.4
+ SB=90002.6 A=0.18 P=2.36 MULT=1
MM1014 N_A_27_392#_M1011_d N_A2_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.185 PD=1.27 PS=1.37 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90003.8
+ SB=90002.2 A=0.18 P=2.36 MULT=1
MM1008 N_A_27_392#_M1008_d N_A3_M1008_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1
+ AD=0.16 AS=0.185 PD=1.32 PS=1.37 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90004.4
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1009 N_A_27_392#_M1008_d N_A3_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1
+ AD=0.16 AS=0.16 PD=1.32 PS=1.32 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90004.9
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1007 N_A_27_392#_M1007_d N_A4_M1007_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.16 PD=1.27 PS=1.32 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90005.4
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1010 N_A_27_392#_M1007_d N_A4_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556 SA=90005.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.8844 P=20.8
c_134 VPB 0 1.25754e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__a41o_4.pxi.spice"
*
.ends
*
*

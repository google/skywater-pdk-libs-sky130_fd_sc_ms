* File: sky130_fd_sc_ms__nor4_2.spice
* Created: Wed Sep  2 12:16:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nor4_2.pex.spice"
.subckt sky130_fd_sc_ms__nor4_2  VNB VPB C D B A Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A	A
* B	B
* D	D
* C	C
* VPB	VPB
* VNB	VNB
MM1005 N_Y_M1005_d N_D_M1005_g N_VGND_M1005_s VNB NLOWVT L=0.15 W=0.74 AD=0.1184
+ AS=0.3329 PD=1.06 PS=3 NRD=6.48 NRS=4.86 M=1 R=4.93333 SA=75000.4 SB=75001.8
+ A=0.111 P=1.78 MULT=1
MM1002 N_VGND_M1002_d N_C_M1002_g N_Y_M1005_d VNB NLOWVT L=0.15 W=0.74 AD=0.1554
+ AS=0.1184 PD=1.16 PS=1.06 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.8 SB=75001.3
+ A=0.111 P=1.78 MULT=1
MM1009 N_Y_M1009_d N_B_M1009_g N_VGND_M1002_d VNB NLOWVT L=0.15 W=0.74 AD=0.1036
+ AS=0.1554 PD=1.02 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.4 SB=75000.7
+ A=0.111 P=1.78 MULT=1
MM1000 N_VGND_M1000_d N_A_M1000_g N_Y_M1009_d VNB NLOWVT L=0.15 W=0.74 AD=0.2627
+ AS=0.1036 PD=2.19 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.8 SB=75000.3
+ A=0.111 P=1.78 MULT=1
MM1001 N_A_119_368#_M1001_d N_C_M1001_g N_A_27_368#_M1001_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1596 AS=0.3136 PD=1.405 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90003.5 A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1004_d N_D_M1004_g N_A_119_368#_M1001_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1652 AS=0.1596 PD=1.415 PS=1.405 NRD=0.8668 NRS=0.8668 M=1 R=6.22222
+ SA=90000.7 SB=90003 A=0.2016 P=2.6 MULT=1
MM1006 N_Y_M1004_d N_D_M1006_g N_A_119_368#_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1652 AS=0.1512 PD=1.415 PS=1.39 NRD=1.7533 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90002.6 A=0.2016 P=2.6 MULT=1
MM1008 N_A_119_368#_M1006_s N_C_M1008_g N_A_27_368#_M1008_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.168 PD=1.39 PS=1.42 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.6
+ SB=90002.1 A=0.2016 P=2.6 MULT=1
MM1003 N_A_493_368#_M1003_d N_B_M1003_g N_A_27_368#_M1008_s VPB PSHORT L=0.18
+ W=1.12 AD=0.2016 AS=0.168 PD=1.48 PS=1.42 NRD=6.1464 NRS=4.3931 M=1 R=6.22222
+ SA=90002.1 SB=90001.6 A=0.2016 P=2.6 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g N_A_493_368#_M1003_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2016 PD=1.39 PS=1.48 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.6
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1010 N_VPWR_M1007_d N_A_M1010_g N_A_493_368#_M1010_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1011 N_A_493_368#_M1010_s N_B_M1011_g N_A_27_368#_M1011_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.5
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__nor4_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__buf_8.pxi.spice
* Created: Fri Aug 28 17:16:08 2020
* 
x_PM_SKY130_FD_SC_MS__BUF_8%A N_A_M1006_g N_A_M1001_g N_A_M1002_g N_A_M1015_g
+ N_A_M1003_g N_A_M1018_g A A A N_A_c_113_n N_A_c_114_n
+ PM_SKY130_FD_SC_MS__BUF_8%A
x_PM_SKY130_FD_SC_MS__BUF_8%A_27_74# N_A_27_74#_M1006_d N_A_27_74#_M1015_d
+ N_A_27_74#_M1001_s N_A_27_74#_M1002_s N_A_27_74#_M1000_g N_A_27_74#_M1004_g
+ N_A_27_74#_M1009_g N_A_27_74#_M1005_g N_A_27_74#_M1012_g N_A_27_74#_M1007_g
+ N_A_27_74#_M1013_g N_A_27_74#_M1008_g N_A_27_74#_M1016_g N_A_27_74#_M1010_g
+ N_A_27_74#_M1017_g N_A_27_74#_M1011_g N_A_27_74#_M1014_g N_A_27_74#_M1019_g
+ N_A_27_74#_M1020_g N_A_27_74#_M1021_g N_A_27_74#_c_193_n N_A_27_74#_c_210_n
+ N_A_27_74#_c_211_n N_A_27_74#_c_194_n N_A_27_74#_c_195_n N_A_27_74#_c_226_n
+ N_A_27_74#_c_212_n N_A_27_74#_c_196_n N_A_27_74#_c_197_n N_A_27_74#_c_238_n
+ N_A_27_74#_c_198_n N_A_27_74#_c_262_p N_A_27_74#_c_241_n N_A_27_74#_c_199_n
+ N_A_27_74#_c_200_n N_A_27_74#_c_201_n PM_SKY130_FD_SC_MS__BUF_8%A_27_74#
x_PM_SKY130_FD_SC_MS__BUF_8%VPWR N_VPWR_M1001_d N_VPWR_M1003_d N_VPWR_M1005_d
+ N_VPWR_M1008_d N_VPWR_M1011_d N_VPWR_M1021_d N_VPWR_c_418_n N_VPWR_c_419_n
+ N_VPWR_c_420_n N_VPWR_c_421_n N_VPWR_c_422_n N_VPWR_c_423_n N_VPWR_c_424_n
+ VPWR N_VPWR_c_425_n N_VPWR_c_426_n N_VPWR_c_427_n N_VPWR_c_428_n
+ N_VPWR_c_429_n N_VPWR_c_430_n N_VPWR_c_431_n N_VPWR_c_432_n N_VPWR_c_433_n
+ N_VPWR_c_434_n N_VPWR_c_417_n PM_SKY130_FD_SC_MS__BUF_8%VPWR
x_PM_SKY130_FD_SC_MS__BUF_8%X N_X_M1000_d N_X_M1012_d N_X_M1016_d N_X_M1019_d
+ N_X_M1004_s N_X_M1007_s N_X_M1010_s N_X_M1014_s N_X_c_506_n N_X_c_518_n
+ N_X_c_507_n N_X_c_508_n N_X_c_519_n N_X_c_520_n N_X_c_509_n N_X_c_521_n
+ N_X_c_510_n N_X_c_522_n N_X_c_511_n N_X_c_523_n N_X_c_512_n N_X_c_524_n
+ N_X_c_513_n N_X_c_514_n N_X_c_515_n N_X_c_526_n N_X_c_516_n N_X_c_527_n
+ N_X_c_517_n X X X X PM_SKY130_FD_SC_MS__BUF_8%X
x_PM_SKY130_FD_SC_MS__BUF_8%VGND N_VGND_M1006_s N_VGND_M1018_s N_VGND_M1009_s
+ N_VGND_M1013_s N_VGND_M1017_s N_VGND_M1020_s N_VGND_c_663_n N_VGND_c_664_n
+ N_VGND_c_665_n N_VGND_c_666_n N_VGND_c_667_n N_VGND_c_668_n N_VGND_c_669_n
+ N_VGND_c_670_n N_VGND_c_671_n N_VGND_c_672_n N_VGND_c_673_n N_VGND_c_674_n
+ N_VGND_c_675_n VGND N_VGND_c_676_n N_VGND_c_677_n N_VGND_c_678_n
+ N_VGND_c_679_n N_VGND_c_680_n N_VGND_c_681_n PM_SKY130_FD_SC_MS__BUF_8%VGND
cc_1 VNB N_A_M1006_g 0.0325279f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_M1015_g 0.0237982f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=0.74
cc_3 VNB N_A_M1018_g 0.0227248f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=0.74
cc_4 VNB N_A_c_113_n 0.0166485f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_5 VNB N_A_c_114_n 0.0568652f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.515
cc_6 VNB N_A_27_74#_M1000_g 0.0197781f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=0.74
cc_7 VNB N_A_27_74#_M1004_g 0.00164514f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=2.4
cc_8 VNB N_A_27_74#_M1009_g 0.0212166f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=0.74
cc_9 VNB N_A_27_74#_M1005_g 0.00165901f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_10 VNB N_A_27_74#_M1012_g 0.0217898f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.515
cc_11 VNB N_A_27_74#_M1007_g 0.00160182f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_12 VNB N_A_27_74#_M1013_g 0.0225551f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_13 VNB N_A_27_74#_M1008_g 0.00160182f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.515
cc_14 VNB N_A_27_74#_M1016_g 0.0225551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_74#_M1010_g 0.00160182f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_16 VNB N_A_27_74#_M1017_g 0.0225551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_74#_M1011_g 0.00158401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_74#_M1014_g 0.00159466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_74#_M1019_g 0.0225878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_74#_M1020_g 0.02608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_74#_M1021_g 0.00233655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_74#_c_193_n 0.0266107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_74#_c_194_n 0.00351687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_74#_c_195_n 0.00998227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_74#_c_196_n 0.00179731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_74#_c_197_n 0.0043023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_74#_c_198_n 4.30857e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_74#_c_199_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_74#_c_200_n 0.00335789f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_74#_c_201_n 0.196361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_417_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_X_c_506_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_33 VNB N_X_c_507_n 0.00317099f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_34 VNB N_X_c_508_n 0.00140587f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.515
cc_35 VNB N_X_c_509_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_36 VNB N_X_c_510_n 0.00311987f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_37 VNB N_X_c_511_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_X_c_512_n 0.00311987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_X_c_513_n 0.0024448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_X_c_514_n 0.00141267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_515_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_X_c_516_n 0.00230427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_X_c_517_n 0.00181295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_663_n 0.0055945f $X=-0.19 $Y=-0.245 $X2=1.4 $Y2=1.35
cc_45 VNB N_VGND_c_664_n 0.00256838f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_46 VNB N_VGND_c_665_n 0.00498656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_666_n 0.00830803f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.515
cc_48 VNB N_VGND_c_667_n 0.00831705f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.515
cc_49 VNB N_VGND_c_668_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_50 VNB N_VGND_c_669_n 0.0551405f $X=-0.19 $Y=-0.245 $X2=1.265 $Y2=1.515
cc_51 VNB N_VGND_c_670_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_671_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_53 VNB N_VGND_c_672_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_673_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.565
cc_55 VNB N_VGND_c_674_n 0.0186948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_675_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_57 VNB N_VGND_c_676_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_677_n 0.0167636f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_678_n 0.0188148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_679_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_680_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_681_n 0.322609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VPB N_A_M1001_g 0.027583f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_64 VPB N_A_M1002_g 0.0204965f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_65 VPB N_A_M1003_g 0.0213785f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=2.4
cc_66 VPB N_A_c_113_n 0.0131369f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_67 VPB N_A_c_114_n 0.00839581f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.515
cc_68 VPB N_A_27_74#_M1004_g 0.0227023f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=2.4
cc_69 VPB N_A_27_74#_M1005_g 0.0232841f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_70 VPB N_A_27_74#_M1007_g 0.0226705f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_71 VPB N_A_27_74#_M1008_g 0.0226708f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.515
cc_72 VPB N_A_27_74#_M1010_g 0.0226705f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_73 VPB N_A_27_74#_M1011_g 0.0224909f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_27_74#_M1014_g 0.0226614f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_27_74#_M1021_g 0.0275992f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_27_74#_c_210_n 0.00739392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_A_27_74#_c_211_n 0.0352219f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_27_74#_c_212_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_79 VPB N_A_27_74#_c_198_n 0.00285251f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_418_n 0.00797179f $X=-0.19 $Y=1.66 $X2=1.4 $Y2=0.74
cc_81 VPB N_VPWR_c_419_n 0.00554449f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_82 VPB N_VPWR_c_420_n 0.00884785f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.515
cc_83 VPB N_VPWR_c_421_n 0.00884785f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.515
cc_84 VPB N_VPWR_c_422_n 0.00884629f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_85 VPB N_VPWR_c_423_n 0.0120875f $X=-0.19 $Y=1.66 $X2=1.265 $Y2=1.515
cc_86 VPB N_VPWR_c_424_n 0.0645562f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=1.515
cc_87 VPB N_VPWR_c_425_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_88 VPB N_VPWR_c_426_n 0.0194914f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_427_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_428_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_429_n 0.0195592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_430_n 0.0234893f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_431_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_432_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_433_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_434_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_417_n 0.0772804f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_X_c_518_n 0.00275675f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.515
cc_99 VPB N_X_c_519_n 0.00249468f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.515
cc_100 VPB N_X_c_520_n 0.00273995f $X=-0.19 $Y=1.66 $X2=0.97 $Y2=1.515
cc_101 VPB N_X_c_521_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_102 VPB N_X_c_522_n 0.00249468f $X=-0.19 $Y=1.66 $X2=1.2 $Y2=1.565
cc_103 VPB N_X_c_523_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_X_c_524_n 0.00240456f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_X_c_514_n 8.47603e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_X_c_526_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_X_c_527_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB X 0.00181295f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB X 0.0024448f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 N_A_M1018_g N_A_27_74#_M1000_g 0.0311454f $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_111 N_A_c_114_n N_A_27_74#_M1004_g 0.0321237f $X=1.41 $Y=1.515 $X2=0 $Y2=0
cc_112 N_A_M1006_g N_A_27_74#_c_193_n 0.00159319f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_113 N_A_M1001_g N_A_27_74#_c_210_n 8.84614e-19 $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_114 N_A_c_113_n N_A_27_74#_c_210_n 0.0259449f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_115 N_A_M1001_g N_A_27_74#_c_211_n 0.0121004f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_116 N_A_M1002_g N_A_27_74#_c_211_n 6.50516e-19 $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_117 N_A_M1006_g N_A_27_74#_c_194_n 0.0139147f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_118 N_A_M1015_g N_A_27_74#_c_194_n 0.0140682f $X=0.97 $Y=0.74 $X2=0 $Y2=0
cc_119 N_A_c_113_n N_A_27_74#_c_194_n 0.0554204f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_120 N_A_c_114_n N_A_27_74#_c_194_n 0.00346768f $X=1.41 $Y=1.515 $X2=0 $Y2=0
cc_121 N_A_c_113_n N_A_27_74#_c_195_n 0.0216404f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_122 N_A_M1001_g N_A_27_74#_c_226_n 0.012931f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_123 N_A_M1002_g N_A_27_74#_c_226_n 0.012931f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_124 N_A_c_113_n N_A_27_74#_c_226_n 0.0391869f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_125 N_A_c_114_n N_A_27_74#_c_226_n 4.90767e-19 $X=1.41 $Y=1.515 $X2=0 $Y2=0
cc_126 N_A_M1001_g N_A_27_74#_c_212_n 6.50516e-19 $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_127 N_A_M1002_g N_A_27_74#_c_212_n 0.0119382f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_128 N_A_M1003_g N_A_27_74#_c_212_n 0.0120649f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_129 N_A_M1015_g N_A_27_74#_c_196_n 4.04737e-19 $X=0.97 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A_M1018_g N_A_27_74#_c_196_n 3.92313e-19 $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A_M1018_g N_A_27_74#_c_197_n 0.0135996f $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A_c_113_n N_A_27_74#_c_197_n 0.0118433f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_133 N_A_c_114_n N_A_27_74#_c_197_n 0.00103766f $X=1.41 $Y=1.515 $X2=0 $Y2=0
cc_134 N_A_M1003_g N_A_27_74#_c_238_n 0.014986f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_135 N_A_c_113_n N_A_27_74#_c_238_n 0.00580317f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_136 N_A_M1003_g N_A_27_74#_c_198_n 0.00349774f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_137 N_A_M1002_g N_A_27_74#_c_241_n 8.84614e-19 $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_138 N_A_M1003_g N_A_27_74#_c_241_n 8.84614e-19 $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_139 N_A_c_113_n N_A_27_74#_c_241_n 0.0235495f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_140 N_A_c_114_n N_A_27_74#_c_241_n 5.54777e-19 $X=1.41 $Y=1.515 $X2=0 $Y2=0
cc_141 N_A_c_113_n N_A_27_74#_c_199_n 0.0146029f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_142 N_A_c_114_n N_A_27_74#_c_199_n 0.00236901f $X=1.41 $Y=1.515 $X2=0 $Y2=0
cc_143 N_A_M1018_g N_A_27_74#_c_200_n 0.00394038f $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A_c_113_n N_A_27_74#_c_200_n 0.0341212f $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_145 N_A_c_114_n N_A_27_74#_c_200_n 0.00349774f $X=1.41 $Y=1.515 $X2=0 $Y2=0
cc_146 N_A_c_113_n N_A_27_74#_c_201_n 2.37596e-19 $X=1.265 $Y=1.515 $X2=0 $Y2=0
cc_147 N_A_c_114_n N_A_27_74#_c_201_n 0.0143466f $X=1.41 $Y=1.515 $X2=0 $Y2=0
cc_148 N_A_M1001_g N_VPWR_c_418_n 0.0027763f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_149 N_A_M1002_g N_VPWR_c_418_n 0.0027763f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_150 N_A_M1003_g N_VPWR_c_419_n 0.002979f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_151 N_A_M1002_g N_VPWR_c_425_n 0.005209f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_152 N_A_M1003_g N_VPWR_c_425_n 0.005209f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_153 N_A_M1001_g N_VPWR_c_430_n 0.005209f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_154 N_A_M1001_g N_VPWR_c_417_n 0.00986025f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_155 N_A_M1002_g N_VPWR_c_417_n 0.00982266f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_156 N_A_M1003_g N_VPWR_c_417_n 0.00982376f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_157 N_A_M1006_g N_VGND_c_663_n 0.0136079f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_158 N_A_M1015_g N_VGND_c_663_n 0.00238937f $X=0.97 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A_M1015_g N_VGND_c_664_n 4.78024e-19 $X=0.97 $Y=0.74 $X2=0 $Y2=0
cc_160 N_A_M1018_g N_VGND_c_664_n 0.010688f $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A_M1006_g N_VGND_c_676_n 0.00383152f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A_M1015_g N_VGND_c_677_n 0.00461464f $X=0.97 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A_M1018_g N_VGND_c_677_n 0.00383152f $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A_M1006_g N_VGND_c_681_n 0.00761198f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A_M1015_g N_VGND_c_681_n 0.00907982f $X=0.97 $Y=0.74 $X2=0 $Y2=0
cc_166 N_A_M1018_g N_VGND_c_681_n 0.0075754f $X=1.4 $Y=0.74 $X2=0 $Y2=0
cc_167 N_A_27_74#_c_226_n N_VPWR_M1001_d 0.00314376f $X=1.02 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_168 N_A_27_74#_c_238_n N_VPWR_M1003_d 0.00358067f $X=1.6 $Y=2.035 $X2=0 $Y2=0
cc_169 N_A_27_74#_c_198_n N_VPWR_M1003_d 0.00141518f $X=1.685 $Y=1.95 $X2=0
+ $Y2=0
cc_170 N_A_27_74#_c_211_n N_VPWR_c_418_n 0.0233699f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_171 N_A_27_74#_c_226_n N_VPWR_c_418_n 0.0126919f $X=1.02 $Y=2.035 $X2=0 $Y2=0
cc_172 N_A_27_74#_c_212_n N_VPWR_c_418_n 0.0233699f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_173 N_A_27_74#_M1004_g N_VPWR_c_419_n 0.0124987f $X=1.86 $Y=2.4 $X2=0 $Y2=0
cc_174 N_A_27_74#_M1005_g N_VPWR_c_419_n 7.12435e-19 $X=2.36 $Y=2.4 $X2=0 $Y2=0
cc_175 N_A_27_74#_c_212_n N_VPWR_c_419_n 0.0234083f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_176 N_A_27_74#_c_238_n N_VPWR_c_419_n 0.0136051f $X=1.6 $Y=2.035 $X2=0 $Y2=0
cc_177 N_A_27_74#_c_262_p N_VPWR_c_419_n 7.30215e-19 $X=4.64 $Y=1.465 $X2=0
+ $Y2=0
cc_178 N_A_27_74#_M1005_g N_VPWR_c_420_n 0.00366558f $X=2.36 $Y=2.4 $X2=0 $Y2=0
cc_179 N_A_27_74#_M1007_g N_VPWR_c_420_n 0.0038215f $X=2.86 $Y=2.4 $X2=0 $Y2=0
cc_180 N_A_27_74#_M1008_g N_VPWR_c_421_n 0.00366558f $X=3.31 $Y=2.4 $X2=0 $Y2=0
cc_181 N_A_27_74#_M1010_g N_VPWR_c_421_n 0.0038215f $X=3.81 $Y=2.4 $X2=0 $Y2=0
cc_182 N_A_27_74#_M1011_g N_VPWR_c_422_n 0.00361496f $X=4.26 $Y=2.4 $X2=0 $Y2=0
cc_183 N_A_27_74#_M1014_g N_VPWR_c_422_n 0.00385263f $X=4.745 $Y=2.4 $X2=0 $Y2=0
cc_184 N_A_27_74#_M1021_g N_VPWR_c_424_n 0.00648878f $X=5.21 $Y=2.4 $X2=0 $Y2=0
cc_185 N_A_27_74#_c_212_n N_VPWR_c_425_n 0.0144623f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_186 N_A_27_74#_M1004_g N_VPWR_c_426_n 0.00460063f $X=1.86 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A_27_74#_M1005_g N_VPWR_c_426_n 0.005209f $X=2.36 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A_27_74#_M1007_g N_VPWR_c_427_n 0.005209f $X=2.86 $Y=2.4 $X2=0 $Y2=0
cc_189 N_A_27_74#_M1008_g N_VPWR_c_427_n 0.005209f $X=3.31 $Y=2.4 $X2=0 $Y2=0
cc_190 N_A_27_74#_M1010_g N_VPWR_c_428_n 0.005209f $X=3.81 $Y=2.4 $X2=0 $Y2=0
cc_191 N_A_27_74#_M1011_g N_VPWR_c_428_n 0.005209f $X=4.26 $Y=2.4 $X2=0 $Y2=0
cc_192 N_A_27_74#_M1014_g N_VPWR_c_429_n 0.00537895f $X=4.745 $Y=2.4 $X2=0 $Y2=0
cc_193 N_A_27_74#_M1021_g N_VPWR_c_429_n 0.00515235f $X=5.21 $Y=2.4 $X2=0 $Y2=0
cc_194 N_A_27_74#_c_211_n N_VPWR_c_430_n 0.014549f $X=0.285 $Y=2.815 $X2=0 $Y2=0
cc_195 N_A_27_74#_M1004_g N_VPWR_c_417_n 0.00909043f $X=1.86 $Y=2.4 $X2=0 $Y2=0
cc_196 N_A_27_74#_M1005_g N_VPWR_c_417_n 0.00983242f $X=2.36 $Y=2.4 $X2=0 $Y2=0
cc_197 N_A_27_74#_M1007_g N_VPWR_c_417_n 0.00982082f $X=2.86 $Y=2.4 $X2=0 $Y2=0
cc_198 N_A_27_74#_M1008_g N_VPWR_c_417_n 0.00982754f $X=3.31 $Y=2.4 $X2=0 $Y2=0
cc_199 N_A_27_74#_M1010_g N_VPWR_c_417_n 0.00982082f $X=3.81 $Y=2.4 $X2=0 $Y2=0
cc_200 N_A_27_74#_M1011_g N_VPWR_c_417_n 0.00982612f $X=4.26 $Y=2.4 $X2=0 $Y2=0
cc_201 N_A_27_74#_M1014_g N_VPWR_c_417_n 0.0103679f $X=4.745 $Y=2.4 $X2=0 $Y2=0
cc_202 N_A_27_74#_M1021_g N_VPWR_c_417_n 0.00967962f $X=5.21 $Y=2.4 $X2=0 $Y2=0
cc_203 N_A_27_74#_c_211_n N_VPWR_c_417_n 0.0119743f $X=0.285 $Y=2.815 $X2=0
+ $Y2=0
cc_204 N_A_27_74#_c_212_n N_VPWR_c_417_n 0.0118344f $X=1.185 $Y=2.815 $X2=0
+ $Y2=0
cc_205 N_A_27_74#_M1000_g N_X_c_506_n 3.92313e-19 $X=1.83 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A_27_74#_M1009_g N_X_c_506_n 3.92313e-19 $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A_27_74#_M1004_g N_X_c_518_n 4.37331e-19 $X=1.86 $Y=2.4 $X2=0 $Y2=0
cc_208 N_A_27_74#_M1005_g N_X_c_518_n 0.0145412f $X=2.36 $Y=2.4 $X2=0 $Y2=0
cc_209 N_A_27_74#_M1007_g N_X_c_518_n 6.79538e-19 $X=2.86 $Y=2.4 $X2=0 $Y2=0
cc_210 N_A_27_74#_M1009_g N_X_c_507_n 0.0128315f $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_211 N_A_27_74#_M1012_g N_X_c_507_n 0.0115433f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A_27_74#_c_262_p N_X_c_507_n 0.0500092f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_213 N_A_27_74#_c_201_n N_X_c_507_n 0.00426458f $X=5.21 $Y=1.465 $X2=0 $Y2=0
cc_214 N_A_27_74#_c_262_p N_X_c_508_n 0.0143381f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_215 N_A_27_74#_c_200_n N_X_c_508_n 0.00455444f $X=1.685 $Y=1.095 $X2=0 $Y2=0
cc_216 N_A_27_74#_c_201_n N_X_c_508_n 0.00250705f $X=5.21 $Y=1.465 $X2=0 $Y2=0
cc_217 N_A_27_74#_M1005_g N_X_c_519_n 0.0132272f $X=2.36 $Y=2.4 $X2=0 $Y2=0
cc_218 N_A_27_74#_M1007_g N_X_c_519_n 0.0132272f $X=2.86 $Y=2.4 $X2=0 $Y2=0
cc_219 N_A_27_74#_c_262_p N_X_c_519_n 0.045409f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_220 N_A_27_74#_c_201_n N_X_c_519_n 0.00347377f $X=5.21 $Y=1.465 $X2=0 $Y2=0
cc_221 N_A_27_74#_M1004_g N_X_c_520_n 4.00652e-19 $X=1.86 $Y=2.4 $X2=0 $Y2=0
cc_222 N_A_27_74#_M1005_g N_X_c_520_n 0.00134395f $X=2.36 $Y=2.4 $X2=0 $Y2=0
cc_223 N_A_27_74#_c_198_n N_X_c_520_n 0.00293375f $X=1.685 $Y=1.95 $X2=0 $Y2=0
cc_224 N_A_27_74#_c_262_p N_X_c_520_n 0.0276979f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_225 N_A_27_74#_c_201_n N_X_c_520_n 0.00359665f $X=5.21 $Y=1.465 $X2=0 $Y2=0
cc_226 N_A_27_74#_M1009_g N_X_c_509_n 8.71574e-19 $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_227 N_A_27_74#_M1012_g N_X_c_509_n 0.0089455f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A_27_74#_M1013_g N_X_c_509_n 0.00916694f $X=3.19 $Y=0.74 $X2=0 $Y2=0
cc_229 N_A_27_74#_M1016_g N_X_c_509_n 6.18925e-19 $X=3.76 $Y=0.74 $X2=0 $Y2=0
cc_230 N_A_27_74#_M1005_g N_X_c_521_n 6.46654e-19 $X=2.36 $Y=2.4 $X2=0 $Y2=0
cc_231 N_A_27_74#_M1007_g N_X_c_521_n 0.0139698f $X=2.86 $Y=2.4 $X2=0 $Y2=0
cc_232 N_A_27_74#_M1008_g N_X_c_521_n 0.0145605f $X=3.31 $Y=2.4 $X2=0 $Y2=0
cc_233 N_A_27_74#_M1010_g N_X_c_521_n 6.79538e-19 $X=3.81 $Y=2.4 $X2=0 $Y2=0
cc_234 N_A_27_74#_M1013_g N_X_c_510_n 0.0118691f $X=3.19 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A_27_74#_M1016_g N_X_c_510_n 0.0118691f $X=3.76 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A_27_74#_c_262_p N_X_c_510_n 0.0493541f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_237 N_A_27_74#_c_201_n N_X_c_510_n 0.00591282f $X=5.21 $Y=1.465 $X2=0 $Y2=0
cc_238 N_A_27_74#_M1008_g N_X_c_522_n 0.0132272f $X=3.31 $Y=2.4 $X2=0 $Y2=0
cc_239 N_A_27_74#_M1010_g N_X_c_522_n 0.0132272f $X=3.81 $Y=2.4 $X2=0 $Y2=0
cc_240 N_A_27_74#_c_262_p N_X_c_522_n 0.045409f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_241 N_A_27_74#_c_201_n N_X_c_522_n 0.00327677f $X=5.21 $Y=1.465 $X2=0 $Y2=0
cc_242 N_A_27_74#_M1013_g N_X_c_511_n 6.18925e-19 $X=3.19 $Y=0.74 $X2=0 $Y2=0
cc_243 N_A_27_74#_M1016_g N_X_c_511_n 0.00916694f $X=3.76 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A_27_74#_M1017_g N_X_c_511_n 0.00916694f $X=4.19 $Y=0.74 $X2=0 $Y2=0
cc_245 N_A_27_74#_M1019_g N_X_c_511_n 6.18925e-19 $X=4.76 $Y=0.74 $X2=0 $Y2=0
cc_246 N_A_27_74#_M1008_g N_X_c_523_n 6.46654e-19 $X=3.31 $Y=2.4 $X2=0 $Y2=0
cc_247 N_A_27_74#_M1010_g N_X_c_523_n 0.0139698f $X=3.81 $Y=2.4 $X2=0 $Y2=0
cc_248 N_A_27_74#_M1011_g N_X_c_523_n 0.0145225f $X=4.26 $Y=2.4 $X2=0 $Y2=0
cc_249 N_A_27_74#_M1014_g N_X_c_523_n 6.87723e-19 $X=4.745 $Y=2.4 $X2=0 $Y2=0
cc_250 N_A_27_74#_M1017_g N_X_c_512_n 0.0118691f $X=4.19 $Y=0.74 $X2=0 $Y2=0
cc_251 N_A_27_74#_M1019_g N_X_c_512_n 0.0118144f $X=4.76 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A_27_74#_c_262_p N_X_c_512_n 0.0490309f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_253 N_A_27_74#_c_201_n N_X_c_512_n 0.00583402f $X=5.21 $Y=1.465 $X2=0 $Y2=0
cc_254 N_A_27_74#_M1011_g N_X_c_524_n 0.0131424f $X=4.26 $Y=2.4 $X2=0 $Y2=0
cc_255 N_A_27_74#_M1014_g N_X_c_524_n 0.0144547f $X=4.745 $Y=2.4 $X2=0 $Y2=0
cc_256 N_A_27_74#_c_262_p N_X_c_524_n 0.0443156f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_257 N_A_27_74#_c_201_n N_X_c_524_n 0.00280257f $X=5.21 $Y=1.465 $X2=0 $Y2=0
cc_258 N_A_27_74#_M1017_g N_X_c_513_n 6.18848e-19 $X=4.19 $Y=0.74 $X2=0 $Y2=0
cc_259 N_A_27_74#_M1019_g N_X_c_513_n 0.00918133f $X=4.76 $Y=0.74 $X2=0 $Y2=0
cc_260 N_A_27_74#_M1020_g N_X_c_513_n 0.00768946f $X=5.195 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A_27_74#_M1014_g N_X_c_514_n 0.00259597f $X=4.745 $Y=2.4 $X2=0 $Y2=0
cc_262 N_A_27_74#_M1019_g N_X_c_514_n 0.00257778f $X=4.76 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A_27_74#_M1020_g N_X_c_514_n 0.00858408f $X=5.195 $Y=0.74 $X2=0 $Y2=0
cc_264 N_A_27_74#_M1021_g N_X_c_514_n 0.0086473f $X=5.21 $Y=2.4 $X2=0 $Y2=0
cc_265 N_A_27_74#_c_262_p N_X_c_514_n 0.0249855f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_266 N_A_27_74#_c_201_n N_X_c_514_n 0.025049f $X=5.21 $Y=1.465 $X2=0 $Y2=0
cc_267 N_A_27_74#_M1012_g N_X_c_515_n 9.7541e-19 $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_268 N_A_27_74#_M1013_g N_X_c_515_n 9.7541e-19 $X=3.19 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A_27_74#_c_262_p N_X_c_515_n 0.0276081f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_270 N_A_27_74#_c_201_n N_X_c_515_n 0.00272398f $X=5.21 $Y=1.465 $X2=0 $Y2=0
cc_271 N_A_27_74#_M1007_g N_X_c_526_n 0.00135419f $X=2.86 $Y=2.4 $X2=0 $Y2=0
cc_272 N_A_27_74#_M1008_g N_X_c_526_n 0.00135419f $X=3.31 $Y=2.4 $X2=0 $Y2=0
cc_273 N_A_27_74#_c_262_p N_X_c_526_n 0.0275631f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_274 N_A_27_74#_c_201_n N_X_c_526_n 0.00245159f $X=5.21 $Y=1.465 $X2=0 $Y2=0
cc_275 N_A_27_74#_M1016_g N_X_c_516_n 9.7541e-19 $X=3.76 $Y=0.74 $X2=0 $Y2=0
cc_276 N_A_27_74#_M1017_g N_X_c_516_n 9.7541e-19 $X=4.19 $Y=0.74 $X2=0 $Y2=0
cc_277 N_A_27_74#_c_262_p N_X_c_516_n 0.0276081f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_278 N_A_27_74#_c_201_n N_X_c_516_n 0.00258594f $X=5.21 $Y=1.465 $X2=0 $Y2=0
cc_279 N_A_27_74#_M1010_g N_X_c_527_n 0.00135419f $X=3.81 $Y=2.4 $X2=0 $Y2=0
cc_280 N_A_27_74#_M1011_g N_X_c_527_n 0.00135419f $X=4.26 $Y=2.4 $X2=0 $Y2=0
cc_281 N_A_27_74#_c_262_p N_X_c_527_n 0.0275631f $X=4.64 $Y=1.465 $X2=0 $Y2=0
cc_282 N_A_27_74#_c_201_n N_X_c_527_n 0.00231354f $X=5.21 $Y=1.465 $X2=0 $Y2=0
cc_283 N_A_27_74#_M1019_g N_X_c_517_n 0.00132627f $X=4.76 $Y=0.74 $X2=0 $Y2=0
cc_284 N_A_27_74#_M1020_g N_X_c_517_n 0.00205051f $X=5.195 $Y=0.74 $X2=0 $Y2=0
cc_285 N_A_27_74#_c_201_n N_X_c_517_n 0.00150825f $X=5.21 $Y=1.465 $X2=0 $Y2=0
cc_286 N_A_27_74#_M1014_g X 0.00112654f $X=4.745 $Y=2.4 $X2=0 $Y2=0
cc_287 N_A_27_74#_M1021_g X 0.00387947f $X=5.21 $Y=2.4 $X2=0 $Y2=0
cc_288 N_A_27_74#_c_201_n X 0.00150825f $X=5.21 $Y=1.465 $X2=0 $Y2=0
cc_289 N_A_27_74#_M1011_g X 6.3296e-19 $X=4.26 $Y=2.4 $X2=0 $Y2=0
cc_290 N_A_27_74#_M1014_g X 0.0127662f $X=4.745 $Y=2.4 $X2=0 $Y2=0
cc_291 N_A_27_74#_M1021_g X 0.0140349f $X=5.21 $Y=2.4 $X2=0 $Y2=0
cc_292 N_A_27_74#_c_194_n N_VGND_M1006_s 0.00224297f $X=1.1 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_293 N_A_27_74#_c_197_n N_VGND_M1018_s 9.61034e-19 $X=1.6 $Y=1.095 $X2=0 $Y2=0
cc_294 N_A_27_74#_c_200_n N_VGND_M1018_s 0.00130977f $X=1.685 $Y=1.095 $X2=0
+ $Y2=0
cc_295 N_A_27_74#_c_193_n N_VGND_c_663_n 0.0182902f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_296 N_A_27_74#_c_194_n N_VGND_c_663_n 0.0189527f $X=1.1 $Y=1.095 $X2=0 $Y2=0
cc_297 N_A_27_74#_c_196_n N_VGND_c_663_n 0.00123668f $X=1.185 $Y=0.515 $X2=0
+ $Y2=0
cc_298 N_A_27_74#_M1000_g N_VGND_c_664_n 0.01069f $X=1.83 $Y=0.74 $X2=0 $Y2=0
cc_299 N_A_27_74#_M1009_g N_VGND_c_664_n 4.71636e-19 $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_300 N_A_27_74#_c_196_n N_VGND_c_664_n 0.0182488f $X=1.185 $Y=0.515 $X2=0
+ $Y2=0
cc_301 N_A_27_74#_c_197_n N_VGND_c_664_n 0.00731846f $X=1.6 $Y=1.095 $X2=0 $Y2=0
cc_302 N_A_27_74#_c_262_p N_VGND_c_664_n 3.19484e-19 $X=4.64 $Y=1.465 $X2=0
+ $Y2=0
cc_303 N_A_27_74#_c_200_n N_VGND_c_664_n 0.00988848f $X=1.685 $Y=1.095 $X2=0
+ $Y2=0
cc_304 N_A_27_74#_M1000_g N_VGND_c_665_n 4.56715e-19 $X=1.83 $Y=0.74 $X2=0 $Y2=0
cc_305 N_A_27_74#_M1009_g N_VGND_c_665_n 0.00956829f $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_306 N_A_27_74#_M1012_g N_VGND_c_665_n 0.00406778f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_307 N_A_27_74#_M1013_g N_VGND_c_666_n 0.00454042f $X=3.19 $Y=0.74 $X2=0 $Y2=0
cc_308 N_A_27_74#_M1016_g N_VGND_c_666_n 0.00454042f $X=3.76 $Y=0.74 $X2=0 $Y2=0
cc_309 N_A_27_74#_M1017_g N_VGND_c_667_n 0.00454042f $X=4.19 $Y=0.74 $X2=0 $Y2=0
cc_310 N_A_27_74#_M1019_g N_VGND_c_667_n 0.0045466f $X=4.76 $Y=0.74 $X2=0 $Y2=0
cc_311 N_A_27_74#_M1020_g N_VGND_c_669_n 0.0184966f $X=5.195 $Y=0.74 $X2=0 $Y2=0
cc_312 N_A_27_74#_M1000_g N_VGND_c_670_n 0.00383152f $X=1.83 $Y=0.74 $X2=0 $Y2=0
cc_313 N_A_27_74#_M1009_g N_VGND_c_670_n 0.00383152f $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_314 N_A_27_74#_M1012_g N_VGND_c_672_n 0.00434272f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_315 N_A_27_74#_M1013_g N_VGND_c_672_n 0.00434272f $X=3.19 $Y=0.74 $X2=0 $Y2=0
cc_316 N_A_27_74#_M1016_g N_VGND_c_674_n 0.00434272f $X=3.76 $Y=0.74 $X2=0 $Y2=0
cc_317 N_A_27_74#_M1017_g N_VGND_c_674_n 0.00434272f $X=4.19 $Y=0.74 $X2=0 $Y2=0
cc_318 N_A_27_74#_c_193_n N_VGND_c_676_n 0.011066f $X=0.28 $Y=0.515 $X2=0 $Y2=0
cc_319 N_A_27_74#_c_196_n N_VGND_c_677_n 0.00749631f $X=1.185 $Y=0.515 $X2=0
+ $Y2=0
cc_320 N_A_27_74#_M1019_g N_VGND_c_678_n 0.00434272f $X=4.76 $Y=0.74 $X2=0 $Y2=0
cc_321 N_A_27_74#_M1020_g N_VGND_c_678_n 0.00434272f $X=5.195 $Y=0.74 $X2=0
+ $Y2=0
cc_322 N_A_27_74#_M1000_g N_VGND_c_681_n 0.0075754f $X=1.83 $Y=0.74 $X2=0 $Y2=0
cc_323 N_A_27_74#_M1009_g N_VGND_c_681_n 0.0075754f $X=2.26 $Y=0.74 $X2=0 $Y2=0
cc_324 N_A_27_74#_M1012_g N_VGND_c_681_n 0.00820718f $X=2.76 $Y=0.74 $X2=0 $Y2=0
cc_325 N_A_27_74#_M1013_g N_VGND_c_681_n 0.00821294f $X=3.19 $Y=0.74 $X2=0 $Y2=0
cc_326 N_A_27_74#_M1016_g N_VGND_c_681_n 0.00821294f $X=3.76 $Y=0.74 $X2=0 $Y2=0
cc_327 N_A_27_74#_M1017_g N_VGND_c_681_n 0.00821294f $X=4.19 $Y=0.74 $X2=0 $Y2=0
cc_328 N_A_27_74#_M1019_g N_VGND_c_681_n 0.00821344f $X=4.76 $Y=0.74 $X2=0 $Y2=0
cc_329 N_A_27_74#_M1020_g N_VGND_c_681_n 0.00823984f $X=5.195 $Y=0.74 $X2=0
+ $Y2=0
cc_330 N_A_27_74#_c_193_n N_VGND_c_681_n 0.00915947f $X=0.28 $Y=0.515 $X2=0
+ $Y2=0
cc_331 N_A_27_74#_c_196_n N_VGND_c_681_n 0.0062048f $X=1.185 $Y=0.515 $X2=0
+ $Y2=0
cc_332 N_VPWR_c_419_n N_X_c_518_n 0.0256025f $X=1.635 $Y=2.455 $X2=0 $Y2=0
cc_333 N_VPWR_c_420_n N_X_c_518_n 0.0283501f $X=2.585 $Y=2.305 $X2=0 $Y2=0
cc_334 N_VPWR_c_426_n N_X_c_518_n 0.014549f $X=2.5 $Y=3.33 $X2=0 $Y2=0
cc_335 N_VPWR_c_417_n N_X_c_518_n 0.0119743f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_336 N_VPWR_M1005_d N_X_c_519_n 0.00218982f $X=2.45 $Y=1.84 $X2=0 $Y2=0
cc_337 N_VPWR_c_420_n N_X_c_519_n 0.0167599f $X=2.585 $Y=2.305 $X2=0 $Y2=0
cc_338 N_VPWR_c_420_n N_X_c_521_n 0.0322767f $X=2.585 $Y=2.305 $X2=0 $Y2=0
cc_339 N_VPWR_c_421_n N_X_c_521_n 0.0283501f $X=3.535 $Y=2.305 $X2=0 $Y2=0
cc_340 N_VPWR_c_427_n N_X_c_521_n 0.0144623f $X=3.45 $Y=3.33 $X2=0 $Y2=0
cc_341 N_VPWR_c_417_n N_X_c_521_n 0.0118344f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_342 N_VPWR_M1008_d N_X_c_522_n 0.00218982f $X=3.4 $Y=1.84 $X2=0 $Y2=0
cc_343 N_VPWR_c_421_n N_X_c_522_n 0.0167599f $X=3.535 $Y=2.305 $X2=0 $Y2=0
cc_344 N_VPWR_c_421_n N_X_c_523_n 0.0322767f $X=3.535 $Y=2.305 $X2=0 $Y2=0
cc_345 N_VPWR_c_422_n N_X_c_523_n 0.0283501f $X=4.485 $Y=2.305 $X2=0 $Y2=0
cc_346 N_VPWR_c_428_n N_X_c_523_n 0.0144623f $X=4.4 $Y=3.33 $X2=0 $Y2=0
cc_347 N_VPWR_c_417_n N_X_c_523_n 0.0118344f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_348 N_VPWR_M1011_d N_X_c_524_n 0.00203037f $X=4.35 $Y=1.84 $X2=0 $Y2=0
cc_349 N_VPWR_c_422_n N_X_c_524_n 0.0155395f $X=4.485 $Y=2.305 $X2=0 $Y2=0
cc_350 N_VPWR_c_424_n X 0.00634826f $X=5.435 $Y=1.985 $X2=0 $Y2=0
cc_351 N_VPWR_c_422_n X 0.0323494f $X=4.485 $Y=2.305 $X2=0 $Y2=0
cc_352 N_VPWR_c_424_n X 0.0346872f $X=5.435 $Y=1.985 $X2=0 $Y2=0
cc_353 N_VPWR_c_429_n X 0.0147153f $X=5.35 $Y=3.33 $X2=0 $Y2=0
cc_354 N_VPWR_c_417_n X 0.0120673f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_355 N_X_c_507_n N_VGND_M1009_s 0.00250873f $X=2.81 $Y=1.045 $X2=0 $Y2=0
cc_356 N_X_c_510_n N_VGND_M1013_s 0.00374767f $X=3.81 $Y=1.045 $X2=0 $Y2=0
cc_357 N_X_c_512_n N_VGND_M1017_s 0.00374767f $X=4.81 $Y=1.045 $X2=0 $Y2=0
cc_358 N_X_c_506_n N_VGND_c_664_n 0.0182488f $X=2.045 $Y=0.515 $X2=0 $Y2=0
cc_359 N_X_c_506_n N_VGND_c_665_n 0.0164567f $X=2.045 $Y=0.515 $X2=0 $Y2=0
cc_360 N_X_c_507_n N_VGND_c_665_n 0.0209867f $X=2.81 $Y=1.045 $X2=0 $Y2=0
cc_361 N_X_c_509_n N_VGND_c_665_n 0.0173003f $X=2.975 $Y=0.515 $X2=0 $Y2=0
cc_362 N_X_c_509_n N_VGND_c_666_n 0.0173003f $X=2.975 $Y=0.515 $X2=0 $Y2=0
cc_363 N_X_c_510_n N_VGND_c_666_n 0.0248957f $X=3.81 $Y=1.045 $X2=0 $Y2=0
cc_364 N_X_c_511_n N_VGND_c_666_n 0.0173003f $X=3.975 $Y=0.515 $X2=0 $Y2=0
cc_365 N_X_c_511_n N_VGND_c_667_n 0.0173003f $X=3.975 $Y=0.515 $X2=0 $Y2=0
cc_366 N_X_c_512_n N_VGND_c_667_n 0.0248957f $X=4.81 $Y=1.045 $X2=0 $Y2=0
cc_367 N_X_c_513_n N_VGND_c_667_n 0.0173384f $X=4.975 $Y=0.515 $X2=0 $Y2=0
cc_368 N_X_c_513_n N_VGND_c_669_n 0.0236943f $X=4.975 $Y=0.515 $X2=0 $Y2=0
cc_369 N_X_c_517_n N_VGND_c_669_n 0.00795492f $X=4.977 $Y=1.045 $X2=0 $Y2=0
cc_370 N_X_c_506_n N_VGND_c_670_n 0.00749631f $X=2.045 $Y=0.515 $X2=0 $Y2=0
cc_371 N_X_c_509_n N_VGND_c_672_n 0.0144922f $X=2.975 $Y=0.515 $X2=0 $Y2=0
cc_372 N_X_c_511_n N_VGND_c_674_n 0.0144922f $X=3.975 $Y=0.515 $X2=0 $Y2=0
cc_373 N_X_c_513_n N_VGND_c_678_n 0.0147153f $X=4.975 $Y=0.515 $X2=0 $Y2=0
cc_374 N_X_c_506_n N_VGND_c_681_n 0.0062048f $X=2.045 $Y=0.515 $X2=0 $Y2=0
cc_375 N_X_c_509_n N_VGND_c_681_n 0.0118826f $X=2.975 $Y=0.515 $X2=0 $Y2=0
cc_376 N_X_c_511_n N_VGND_c_681_n 0.0118826f $X=3.975 $Y=0.515 $X2=0 $Y2=0
cc_377 N_X_c_513_n N_VGND_c_681_n 0.0120673f $X=4.975 $Y=0.515 $X2=0 $Y2=0

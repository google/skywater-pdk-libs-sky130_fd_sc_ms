* File: sky130_fd_sc_ms__buf_2.spice
* Created: Wed Sep  2 11:59:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__buf_2.pex.spice"
.subckt sky130_fd_sc_ms__buf_2  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_21_260#_M1002_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_A_21_260#_M1005_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.166607 AS=0.1036 PD=1.25478 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1003 N_A_21_260#_M1003_d N_A_M1003_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.144093 PD=1.85 PS=1.08522 NRD=0 NRS=14.988 M=1 R=4.26667
+ SA=75001.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_X_M1000_d N_A_21_260#_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.7392 PD=1.39 PS=3.56 NRD=0 NRS=43.6749 M=1 R=6.22222 SA=90000.6
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1001 N_X_M1000_d N_A_21_260#_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.205298 PD=1.39 PS=1.55849 NRD=0 NRS=0 M=1 R=6.22222 SA=90001
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1004 N_A_21_260#_M1004_d N_A_M1004_g N_VPWR_M1001_s VPB PSHORT L=0.18 W=1
+ AD=0.305 AS=0.183302 PD=2.61 PS=1.39151 NRD=0.9653 NRS=16.7253 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1708 P=9.28
*
.include "sky130_fd_sc_ms__buf_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__dlxbn_1.pex.spice
* Created: Wed Sep  2 12:06:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLXBN_1%D 3 5 8 10 11 14 16
c39 8 0 1.742e-19 $X=0.675 $Y=2.54
r40 14 16 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.592 $Y=1.425
+ $X2=0.592 $Y2=1.26
r41 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.6
+ $Y=1.425 $X2=0.6 $Y2=1.425
r42 11 15 2.14223 $w=6.68e-07 $l=1.2e-07 $layer=LI1_cond $X=0.72 $Y=1.595
+ $X2=0.6 $Y2=1.595
r43 8 10 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=0.675 $Y=2.54
+ $X2=0.675 $Y2=1.93
r44 5 10 41.9095 $w=3.45e-07 $l=1.72e-07 $layer=POLY_cond $X=0.592 $Y=1.758
+ $X2=0.592 $Y2=1.93
r45 4 14 1.17081 $w=3.45e-07 $l=7e-09 $layer=POLY_cond $X=0.592 $Y=1.432
+ $X2=0.592 $Y2=1.425
r46 4 5 54.5263 $w=3.45e-07 $l=3.26e-07 $layer=POLY_cond $X=0.592 $Y=1.432
+ $X2=0.592 $Y2=1.758
r47 3 16 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.495 $Y=0.875
+ $X2=0.495 $Y2=1.26
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_1%GATE_N 3 7 9 12 13
r41 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.795
+ $X2=1.17 $Y2=1.96
r42 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.795
+ $X2=1.17 $Y2=1.63
r43 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.795 $X2=1.17 $Y2=1.795
r44 9 13 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.17 $Y=2.035 $X2=1.17
+ $Y2=1.795
r45 7 15 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=1.175 $Y=2.54
+ $X2=1.175 $Y2=1.96
r46 3 14 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=1.085 $Y=0.78
+ $X2=1.085 $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_1%A_232_82# 1 2 7 9 11 14 16 18 19 20 25 27 30
+ 36 39 44 48 49 50 54 56 58 63
c133 48 0 1.742e-19 $X=1.4 $Y=2.405
c134 16 0 1.82525e-19 $X=3.19 $Y=1.11
c135 7 0 1.72289e-19 $X=2.145 $Y=1.325
r136 54 64 39.7167 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=3.912 $Y=1.635
+ $X2=3.912 $Y2=1.8
r137 54 63 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=3.912 $Y=1.635
+ $X2=3.912 $Y2=1.47
r138 53 56 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=3.94 $Y=1.635
+ $X2=4.06 $Y2=1.635
r139 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.94
+ $Y=1.635 $X2=3.94 $Y2=1.635
r140 48 50 1.83343 $w=4.38e-07 $l=7e-08 $layer=LI1_cond $X=1.455 $Y=2.405
+ $X2=1.455 $Y2=2.475
r141 48 49 6.73996 $w=4.38e-07 $l=8.5e-08 $layer=LI1_cond $X=1.455 $Y=2.405
+ $X2=1.455 $Y2=2.32
r142 45 58 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.74 $Y=1.415
+ $X2=1.74 $Y2=1.325
r143 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.74
+ $Y=1.415 $X2=1.74 $Y2=1.415
r144 42 44 6.64871 $w=2.58e-07 $l=1.5e-07 $layer=LI1_cond $X=1.59 $Y=1.39
+ $X2=1.74 $Y2=1.39
r145 38 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.06 $Y=1.8
+ $X2=4.06 $Y2=1.635
r146 38 39 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.06 $Y=1.8 $X2=4.06
+ $Y2=2.39
r147 37 50 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=1.675 $Y=2.475
+ $X2=1.455 $Y2=2.475
r148 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.975 $Y=2.475
+ $X2=4.06 $Y2=2.39
r149 36 37 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=3.975 $Y=2.475
+ $X2=1.675 $Y2=2.475
r150 34 42 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.59 $Y=1.52
+ $X2=1.59 $Y2=1.39
r151 34 49 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=1.59 $Y=1.52 $X2=1.59
+ $Y2=2.32
r152 28 42 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=1.3 $Y=1.39
+ $X2=1.59 $Y2=1.39
r153 28 30 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.3 $Y=1.26
+ $X2=1.3 $Y2=1.005
r154 25 64 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=3.95 $Y=2.17
+ $X2=3.95 $Y2=1.8
r155 21 63 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.795 $Y=1.26
+ $X2=3.795 $Y2=1.47
r156 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.72 $Y=1.185
+ $X2=3.795 $Y2=1.26
r157 19 20 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.72 $Y=1.185
+ $X2=3.265 $Y2=1.185
r158 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.19 $Y=1.11
+ $X2=3.265 $Y2=1.185
r159 16 18 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.19 $Y=1.11
+ $X2=3.19 $Y2=0.715
r160 12 27 18.8402 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=2.235 $Y=1.4
+ $X2=2.235 $Y2=1.325
r161 12 14 380.935 $w=1.8e-07 $l=9.8e-07 $layer=POLY_cond $X=2.235 $Y=1.4
+ $X2=2.235 $Y2=2.38
r162 9 27 18.8402 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=2.22 $Y=1.25
+ $X2=2.235 $Y2=1.325
r163 9 11 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.22 $Y=1.25 $X2=2.22
+ $Y2=0.77
r164 8 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.325
+ $X2=1.74 $Y2=1.325
r165 7 27 6.66866 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.145 $Y=1.325
+ $X2=2.235 $Y2=1.325
r166 7 8 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.145 $Y=1.325
+ $X2=1.905 $Y2=1.325
r167 2 48 300 $w=1.7e-07 $l=3.45977e-07 $layer=licon1_PDIFF $count=2 $X=1.265
+ $Y=2.12 $X2=1.4 $Y2=2.405
r168 1 30 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.41 $X2=1.3 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_1%A_27_120# 1 2 9 13 19 23 24 26 32 33
c75 23 0 4.43268e-20 $X=2.7 $Y=1.415
c76 19 0 3.54814e-19 $X=2.535 $Y=0.665
c77 13 0 3.06626e-19 $X=2.8 $Y=0.715
c78 9 0 1.65096e-19 $X=2.78 $Y=2.46
r79 32 33 9.22412 $w=4.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.32 $Y=2.265
+ $X2=0.32 $Y2=2.1
r80 30 33 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=0.18 $Y=1.09
+ $X2=0.18 $Y2=2.1
r81 29 30 11.4519 $w=3.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.27 $Y=0.835
+ $X2=0.27 $Y2=1.09
r82 26 29 5.59758 $w=3.48e-07 $l=1.7e-07 $layer=LI1_cond $X=0.27 $Y=0.665
+ $X2=0.27 $Y2=0.835
r83 24 36 40.7132 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.415
+ $X2=2.705 $Y2=1.58
r84 24 35 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.415
+ $X2=2.705 $Y2=1.25
r85 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.7
+ $Y=1.415 $X2=2.7 $Y2=1.415
r86 21 23 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=2.7 $Y=0.75 $X2=2.7
+ $Y2=1.415
r87 20 26 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.445 $Y=0.665
+ $X2=0.27 $Y2=0.665
r88 19 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.535 $Y=0.665
+ $X2=2.7 $Y2=0.75
r89 19 20 136.353 $w=1.68e-07 $l=2.09e-06 $layer=LI1_cond $X=2.535 $Y=0.665
+ $X2=0.445 $Y2=0.665
r90 13 35 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.8 $Y=0.715 $X2=2.8
+ $Y2=1.25
r91 9 36 342.065 $w=1.8e-07 $l=8.8e-07 $layer=POLY_cond $X=2.78 $Y=2.46 $X2=2.78
+ $Y2=1.58
r92 2 32 300 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=2 $X=0.25
+ $Y=2.12 $X2=0.38 $Y2=2.265
r93 1 29 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.6 $X2=0.28 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_1%A_343_80# 1 2 9 13 14 19 20 21 23 24 26 27
+ 32 35 41
c100 35 0 4.43268e-20 $X=3.25 $Y=1.635
c101 26 0 6.89381e-20 $X=4.095 $Y=0.34
c102 19 0 1.48832e-19 $X=2.16 $Y=1.71
c103 14 0 1.57795e-19 $X=2.075 $Y=1.005
r104 35 38 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=1.635
+ $X2=3.25 $Y2=1.8
r105 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.25
+ $Y=1.635 $X2=3.25 $Y2=1.635
r106 32 34 3.93548 $w=4.03e-07 $l=1.3e-07 $layer=LI1_cond $X=3.12 $Y=1.845
+ $X2=3.25 $Y2=1.845
r107 30 31 4.44175 $w=4.12e-07 $l=1.5e-07 $layer=LI1_cond $X=2.01 $Y=1.965
+ $X2=2.16 $Y2=1.965
r108 27 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.095 $Y=0.34
+ $X2=4.095 $Y2=0.505
r109 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.095
+ $Y=0.34 $X2=4.095 $Y2=0.34
r110 24 26 41.027 $w=2.48e-07 $l=8.9e-07 $layer=LI1_cond $X=3.205 $Y=0.38
+ $X2=4.095 $Y2=0.38
r111 23 32 5.82385 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=3.12 $Y=1.47
+ $X2=3.12 $Y2=1.845
r112 22 24 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.12 $Y=0.505
+ $X2=3.205 $Y2=0.38
r113 22 23 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=3.12 $Y=0.505
+ $X2=3.12 $Y2=1.47
r114 21 31 2.51946 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=1.965
+ $X2=2.16 $Y2=1.965
r115 20 32 11.6947 $w=5.1e-07 $l=5.2156e-07 $layer=LI1_cond $X=2.655 $Y=1.965
+ $X2=3.12 $Y2=1.845
r116 20 21 9.61553 $w=5.08e-07 $l=4.1e-07 $layer=LI1_cond $X=2.655 $Y=1.965
+ $X2=2.245 $Y2=1.965
r117 19 31 5.95845 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=2.16 $Y=1.71
+ $X2=2.16 $Y2=1.965
r118 18 19 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.16 $Y=1.09
+ $X2=2.16 $Y2=1.71
r119 14 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.075 $Y=1.005
+ $X2=2.16 $Y2=1.09
r120 14 16 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.075 $Y=1.005
+ $X2=1.93 $Y2=1.005
r121 13 41 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.185 $Y=0.825
+ $X2=4.185 $Y2=0.505
r122 9 38 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.2 $Y=2.46 $X2=3.2
+ $Y2=1.8
r123 2 30 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=1.865
+ $Y=1.96 $X2=2.01 $Y2=2.12
r124 1 16 182 $w=1.7e-07 $l=7.04344e-07 $layer=licon1_NDIFF $count=1 $X=1.715
+ $Y=0.4 $X2=1.93 $Y2=1.005
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_1%A_863_294# 1 2 9 13 17 19 21 24 26 28 29 32
+ 34 38 40 42 47 49 50 54
c118 49 0 5.45732e-20 $X=4.48 $Y=1.635
c119 17 0 8.68138e-20 $X=6.155 $Y=2.4
c120 13 0 6.89381e-20 $X=4.575 $Y=0.825
r121 56 58 13.3156 $w=3.39e-07 $l=3.7e-07 $layer=LI1_cond $X=5.505 $Y=1.435
+ $X2=5.505 $Y2=1.805
r122 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.625
+ $Y=1.435 $X2=5.625 $Y2=1.435
r123 50 63 40.6969 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=4.482 $Y=1.635
+ $X2=4.482 $Y2=1.8
r124 50 62 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=4.482 $Y=1.635
+ $X2=4.482 $Y2=1.47
r125 49 52 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.48 $Y=1.635
+ $X2=4.48 $Y2=1.805
r126 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.48
+ $Y=1.635 $X2=4.48 $Y2=1.635
r127 47 56 8.96717 $w=3.39e-07 $l=1.79374e-07 $layer=LI1_cond $X=5.475 $Y=1.27
+ $X2=5.505 $Y2=1.435
r128 47 54 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.475 $Y=1.27
+ $X2=5.475 $Y2=0.96
r129 42 44 28.1332 $w=3.38e-07 $l=8.3e-07 $layer=LI1_cond $X=5.39 $Y=1.905
+ $X2=5.39 $Y2=2.735
r130 40 58 3.05 $w=3.4e-07 $l=1.51658e-07 $layer=LI1_cond $X=5.39 $Y=1.89
+ $X2=5.505 $Y2=1.805
r131 40 42 0.508431 $w=3.38e-07 $l=1.5e-08 $layer=LI1_cond $X=5.39 $Y=1.89
+ $X2=5.39 $Y2=1.905
r132 36 54 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=5.382 $Y=0.783
+ $X2=5.382 $Y2=0.96
r133 36 38 8.05087 $w=3.53e-07 $l=2.48e-07 $layer=LI1_cond $X=5.382 $Y=0.783
+ $X2=5.382 $Y2=0.535
r134 35 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.645 $Y=1.805
+ $X2=4.48 $Y2=1.805
r135 34 58 4.78362 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=5.22 $Y=1.805
+ $X2=5.505 $Y2=1.805
r136 34 35 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=5.22 $Y=1.805
+ $X2=4.645 $Y2=1.805
r137 32 33 2.35697 $w=4.09e-07 $l=2e-08 $layer=POLY_cond $X=6.66 $Y=1.392
+ $X2=6.68 $Y2=1.392
r138 31 32 57.7457 $w=4.09e-07 $l=4.9e-07 $layer=POLY_cond $X=6.17 $Y=1.392
+ $X2=6.66 $Y2=1.392
r139 30 31 1.76773 $w=4.09e-07 $l=1.5e-08 $layer=POLY_cond $X=6.155 $Y=1.392
+ $X2=6.17 $Y2=1.392
r140 29 57 76.939 $w=3.3e-07 $l=4.4e-07 $layer=POLY_cond $X=6.065 $Y=1.435
+ $X2=5.625 $Y2=1.435
r141 29 30 12.5452 $w=4.09e-07 $l=1.09407e-07 $layer=POLY_cond $X=6.065 $Y=1.435
+ $X2=6.155 $Y2=1.392
r142 26 33 26.4068 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.68 $Y=1.185
+ $X2=6.68 $Y2=1.392
r143 26 28 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.68 $Y=1.185
+ $X2=6.68 $Y2=0.835
r144 22 32 21.9932 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.66 $Y=1.6
+ $X2=6.66 $Y2=1.392
r145 22 24 365.387 $w=1.8e-07 $l=9.4e-07 $layer=POLY_cond $X=6.66 $Y=1.6
+ $X2=6.66 $Y2=2.54
r146 19 31 26.4068 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.17 $Y=1.185
+ $X2=6.17 $Y2=1.392
r147 19 21 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=6.17 $Y=1.185
+ $X2=6.17 $Y2=0.74
r148 15 30 21.9932 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.155 $Y=1.6
+ $X2=6.155 $Y2=1.392
r149 15 17 310.968 $w=1.8e-07 $l=8e-07 $layer=POLY_cond $X=6.155 $Y=1.6
+ $X2=6.155 $Y2=2.4
r150 13 62 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=4.575 $Y=0.825
+ $X2=4.575 $Y2=1.47
r151 9 63 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=4.435 $Y=2.17
+ $X2=4.435 $Y2=1.8
r152 2 44 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.25
+ $Y=1.76 $X2=5.385 $Y2=2.735
r153 2 42 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.25
+ $Y=1.76 $X2=5.385 $Y2=1.905
r154 1 38 91 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_NDIFF $count=2 $X=5.22
+ $Y=0.37 $X2=5.37 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_1%A_653_79# 1 2 9 12 15 16 17 19 23 27 30
c76 19 0 1.65096e-19 $X=3.53 $Y=2.135
c77 15 0 5.45732e-20 $X=3.595 $Y=2.05
r78 27 31 40.8642 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=5.07 $Y=1.385
+ $X2=5.07 $Y2=1.55
r79 27 30 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=5.07 $Y=1.385
+ $X2=5.07 $Y2=1.22
r80 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.055
+ $Y=1.385 $X2=5.055 $Y2=1.385
r81 23 26 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.055 $Y=1.215
+ $X2=5.055 $Y2=1.385
r82 20 22 8.61582 $w=5.31e-07 $l=3.75e-07 $layer=LI1_cond $X=3.595 $Y=1.012
+ $X2=3.97 $Y2=1.012
r83 17 22 9.90492 $w=5.31e-07 $l=2.7332e-07 $layer=LI1_cond $X=4.135 $Y=1.215
+ $X2=3.97 $Y2=1.012
r84 16 23 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.89 $Y=1.215
+ $X2=5.055 $Y2=1.215
r85 16 17 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4.89 $Y=1.215
+ $X2=4.135 $Y2=1.215
r86 15 19 0.716491 $w=1.7e-07 $l=1.12916e-07 $layer=LI1_cond $X=3.595 $Y=2.05
+ $X2=3.53 $Y2=2.135
r87 14 20 7.53601 $w=1.7e-07 $l=2.88e-07 $layer=LI1_cond $X=3.595 $Y=1.3
+ $X2=3.595 $Y2=1.012
r88 14 15 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=3.595 $Y=1.3
+ $X2=3.595 $Y2=2.05
r89 12 31 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=5.16 $Y=2.32
+ $X2=5.16 $Y2=1.55
r90 9 30 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.145 $Y=0.74
+ $X2=5.145 $Y2=1.22
r91 2 19 600 $w=1.7e-07 $l=3.15595e-07 $layer=licon1_PDIFF $count=1 $X=3.29
+ $Y=1.96 $X2=3.53 $Y2=2.135
r92 1 22 91 $w=1.7e-07 $l=9.19783e-07 $layer=licon1_NDIFF $count=2 $X=3.265
+ $Y=0.395 $X2=3.97 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_1%A_1350_424# 1 2 9 13 15 16 19 23 27 30
c45 30 0 8.68138e-20 $X=6.892 $Y=1.465
r46 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.335
+ $Y=1.465 $X2=7.335 $Y2=1.465
r47 25 30 1.47678 $w=3.3e-07 $l=1.73e-07 $layer=LI1_cond $X=7.065 $Y=1.465
+ $X2=6.892 $Y2=1.465
r48 25 27 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=7.065 $Y=1.465
+ $X2=7.335 $Y2=1.465
r49 21 30 5.00808 $w=3.42e-07 $l=1.65e-07 $layer=LI1_cond $X=6.892 $Y=1.63
+ $X2=6.892 $Y2=1.465
r50 21 23 21.2116 $w=3.43e-07 $l=6.35e-07 $layer=LI1_cond $X=6.892 $Y=1.63
+ $X2=6.892 $Y2=2.265
r51 17 30 5.00808 $w=3.42e-07 $l=1.65997e-07 $layer=LI1_cond $X=6.89 $Y=1.3
+ $X2=6.892 $Y2=1.465
r52 17 19 15.7614 $w=3.38e-07 $l=4.65e-07 $layer=LI1_cond $X=6.89 $Y=1.3
+ $X2=6.89 $Y2=0.835
r53 15 28 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=7.565 $Y=1.465
+ $X2=7.335 $Y2=1.465
r54 15 16 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.565 $Y=1.465
+ $X2=7.655 $Y2=1.465
r55 11 16 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=7.67 $Y=1.3
+ $X2=7.655 $Y2=1.465
r56 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=7.67 $Y=1.3 $X2=7.67
+ $Y2=0.74
r57 7 16 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.63
+ $X2=7.655 $Y2=1.465
r58 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=7.655 $Y=1.63
+ $X2=7.655 $Y2=2.4
r59 2 23 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.75
+ $Y=2.12 $X2=6.89 $Y2=2.265
r60 1 19 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=6.755
+ $Y=0.56 $X2=6.895 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_1%VPWR 1 2 3 4 5 18 22 24 28 34 38 43 44 46 47
+ 49 50 51 57 75 76 79 82
r86 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r87 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r88 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r89 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r90 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r91 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r92 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r93 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r94 67 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r95 66 69 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r96 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r97 64 82 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=5.02 $Y=3.33 $X2=4.75
+ $Y2=3.33
r98 64 66 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=5.02 $Y=3.33 $X2=5.04
+ $Y2=3.33
r99 63 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r100 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r101 60 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r102 59 62 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r103 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r104 57 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.545 $Y2=3.33
r105 57 62 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.16 $Y2=3.33
r106 55 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r107 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r108 51 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r109 51 80 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r110 49 72 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.265 $Y=3.33
+ $X2=6.96 $Y2=3.33
r111 49 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.265 $Y=3.33
+ $X2=7.39 $Y2=3.33
r112 48 75 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=7.515 $Y=3.33
+ $X2=7.92 $Y2=3.33
r113 48 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.515 $Y=3.33
+ $X2=7.39 $Y2=3.33
r114 46 69 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.3 $Y=3.33 $X2=6
+ $Y2=3.33
r115 46 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.3 $Y=3.33
+ $X2=6.425 $Y2=3.33
r116 45 72 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=6.55 $Y=3.33
+ $X2=6.96 $Y2=3.33
r117 45 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.55 $Y=3.33
+ $X2=6.425 $Y2=3.33
r118 43 54 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.735 $Y=3.33
+ $X2=0.72 $Y2=3.33
r119 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.735 $Y=3.33
+ $X2=0.9 $Y2=3.33
r120 42 59 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.2 $Y2=3.33
r121 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.9 $Y2=3.33
r122 38 41 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=7.39 $Y=1.985
+ $X2=7.39 $Y2=2.815
r123 36 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.39 $Y=3.245
+ $X2=7.39 $Y2=3.33
r124 36 41 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.39 $Y=3.245
+ $X2=7.39 $Y2=2.815
r125 32 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.425 $Y=3.245
+ $X2=6.425 $Y2=3.33
r126 32 34 45.1758 $w=2.48e-07 $l=9.8e-07 $layer=LI1_cond $X=6.425 $Y=3.245
+ $X2=6.425 $Y2=2.265
r127 28 31 12.4038 $w=5.38e-07 $l=5.6e-07 $layer=LI1_cond $X=4.75 $Y=2.175
+ $X2=4.75 $Y2=2.735
r128 26 82 2.26835 $w=5.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.75 $Y=3.245
+ $X2=4.75 $Y2=3.33
r129 26 31 11.2963 $w=5.38e-07 $l=5.1e-07 $layer=LI1_cond $X=4.75 $Y=3.245
+ $X2=4.75 $Y2=2.735
r130 25 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=3.33
+ $X2=2.545 $Y2=3.33
r131 24 82 11.8214 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=4.48 $Y=3.33
+ $X2=4.75 $Y2=3.33
r132 24 25 115.476 $w=1.68e-07 $l=1.77e-06 $layer=LI1_cond $X=4.48 $Y=3.33
+ $X2=2.71 $Y2=3.33
r133 20 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=3.245
+ $X2=2.545 $Y2=3.33
r134 20 22 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.545 $Y=3.245
+ $X2=2.545 $Y2=2.815
r135 16 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.9 $Y=3.245 $X2=0.9
+ $Y2=3.33
r136 16 18 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=0.9 $Y=3.245
+ $X2=0.9 $Y2=2.405
r137 5 41 400 $w=1.7e-07 $l=1.03797e-06 $layer=licon1_PDIFF $count=1 $X=7.3
+ $Y=1.84 $X2=7.43 $Y2=2.815
r138 5 38 400 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=7.3
+ $Y=1.84 $X2=7.43 $Y2=1.985
r139 4 34 300 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=2 $X=6.245
+ $Y=1.84 $X2=6.385 $Y2=2.265
r140 3 31 600 $w=1.7e-07 $l=9.58319e-07 $layer=licon1_PDIFF $count=1 $X=4.525
+ $Y=1.96 $X2=4.935 $Y2=2.735
r141 3 28 600 $w=1.7e-07 $l=3.14643e-07 $layer=licon1_PDIFF $count=1 $X=4.525
+ $Y=1.96 $X2=4.75 $Y2=2.175
r142 2 22 600 $w=1.7e-07 $l=9.5871e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.96 $X2=2.545 $Y2=2.815
r143 1 18 300 $w=1.7e-07 $l=3.45977e-07 $layer=licon1_PDIFF $count=2 $X=0.765
+ $Y=2.12 $X2=0.9 $Y2=2.405
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_1%Q 1 2 9 14 15 16 17 28
r36 21 28 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=5.96 $Y=0.93 $X2=5.96
+ $Y2=0.925
r37 17 30 7.28558 $w=3.38e-07 $l=1.3e-07 $layer=LI1_cond $X=5.96 $Y=0.97
+ $X2=5.96 $Y2=1.1
r38 17 21 1.35582 $w=3.38e-07 $l=4e-08 $layer=LI1_cond $X=5.96 $Y=0.97 $X2=5.96
+ $Y2=0.93
r39 17 28 1.35582 $w=3.38e-07 $l=4e-08 $layer=LI1_cond $X=5.96 $Y=0.885 $X2=5.96
+ $Y2=0.925
r40 16 17 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=5.96 $Y=0.515
+ $X2=5.96 $Y2=0.885
r41 15 30 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=6.045 $Y=1.82
+ $X2=6.045 $Y2=1.1
r42 14 15 8.52431 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=5.947 $Y=1.985
+ $X2=5.947 $Y2=1.82
r43 7 14 0.536754 $w=3.63e-07 $l=1.7e-08 $layer=LI1_cond $X=5.947 $Y=2.002
+ $X2=5.947 $Y2=1.985
r44 7 9 25.6695 $w=3.63e-07 $l=8.13e-07 $layer=LI1_cond $X=5.947 $Y=2.002
+ $X2=5.947 $Y2=2.815
r45 2 14 400 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=5.8
+ $Y=1.84 $X2=5.93 $Y2=1.985
r46 2 9 400 $w=1.7e-07 $l=1.03797e-06 $layer=licon1_PDIFF $count=1 $X=5.8
+ $Y=1.84 $X2=5.93 $Y2=2.815
r47 1 16 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.81
+ $Y=0.37 $X2=5.955 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_1%Q_N 1 2 7 8 9 10 11 12 13
r14 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=7.882 $Y=2.405
+ $X2=7.882 $Y2=2.775
r15 11 12 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=7.882 $Y=1.985
+ $X2=7.882 $Y2=2.405
r16 10 11 11.0084 $w=3.33e-07 $l=3.2e-07 $layer=LI1_cond $X=7.882 $Y=1.665
+ $X2=7.882 $Y2=1.985
r17 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=7.882 $Y=1.295
+ $X2=7.882 $Y2=1.665
r18 8 9 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=7.882 $Y=0.925
+ $X2=7.882 $Y2=1.295
r19 7 8 14.1045 $w=3.33e-07 $l=4.1e-07 $layer=LI1_cond $X=7.882 $Y=0.515
+ $X2=7.882 $Y2=0.925
r20 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.745
+ $Y=1.84 $X2=7.88 $Y2=2.815
r21 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.745
+ $Y=1.84 $X2=7.88 $Y2=1.985
r22 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.745
+ $Y=0.37 $X2=7.885 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLXBN_1%VGND 1 2 3 4 5 18 22 26 29 30 32 33 34 36 41
+ 59 65 66 70 83
r79 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r80 70 73 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.79 $Y=0 $X2=0.79
+ $Y2=0.325
r81 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r82 66 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r83 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r84 63 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.54 $Y=0 $X2=7.415
+ $Y2=0
r85 63 65 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=7.54 $Y=0 $X2=7.92
+ $Y2=0
r86 62 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r87 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r88 59 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.29 $Y=0 $X2=7.415
+ $Y2=0
r89 59 61 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.29 $Y=0 $X2=6.96
+ $Y2=0
r90 58 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r91 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r92 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r93 54 57 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=6 $Y2=0
r94 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r95 52 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r96 51 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r97 49 51 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=2.675 $Y=0
+ $X2=4.56 $Y2=0
r98 48 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r99 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r100 45 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r101 45 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r102 44 47 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r103 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r104 42 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r105 42 44 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r106 41 80 11.1804 $w=3.33e-07 $l=3.25e-07 $layer=LI1_cond $X=2.507 $Y=0
+ $X2=2.507 $Y2=0.325
r107 41 49 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.507 $Y=0
+ $X2=2.675 $Y2=0
r108 41 78 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r109 41 47 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.34 $Y=0 $X2=2.16
+ $Y2=0
r110 39 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r111 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r112 36 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r113 36 38 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0
+ $X2=0.24 $Y2=0
r114 34 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r115 34 78 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=2.64 $Y2=0
r116 32 57 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.3 $Y=0 $X2=6 $Y2=0
r117 32 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.3 $Y=0 $X2=6.425
+ $Y2=0
r118 31 61 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=6.55 $Y=0 $X2=6.96
+ $Y2=0
r119 31 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.55 $Y=0 $X2=6.425
+ $Y2=0
r120 29 51 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.705 $Y=0
+ $X2=4.56 $Y2=0
r121 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=0 $X2=4.87
+ $Y2=0
r122 28 54 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.035 $Y=0 $X2=5.04
+ $Y2=0
r123 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=0 $X2=4.87
+ $Y2=0
r124 24 83 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.415 $Y=0.085
+ $X2=7.415 $Y2=0
r125 24 26 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.415 $Y=0.085
+ $X2=7.415 $Y2=0.515
r126 20 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.425 $Y=0.085
+ $X2=6.425 $Y2=0
r127 20 22 37.1087 $w=2.48e-07 $l=8.05e-07 $layer=LI1_cond $X=6.425 $Y=0.085
+ $X2=6.425 $Y2=0.89
r128 16 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.87 $Y=0.085
+ $X2=4.87 $Y2=0
r129 16 18 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.87 $Y=0.085
+ $X2=4.87 $Y2=0.535
r130 5 26 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=7.31
+ $Y=0.37 $X2=7.455 $Y2=0.515
r131 4 22 182 $w=1.7e-07 $l=6.05475e-07 $layer=licon1_NDIFF $count=1 $X=6.245
+ $Y=0.37 $X2=6.43 $Y2=0.89
r132 3 18 91 $w=1.7e-07 $l=2.56905e-07 $layer=licon1_NDIFF $count=2 $X=4.65
+ $Y=0.615 $X2=4.87 $Y2=0.535
r133 2 80 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=2.295
+ $Y=0.4 $X2=2.505 $Y2=0.325
r134 1 73 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.6 $X2=0.79 $Y2=0.325
.ends


* File: sky130_fd_sc_ms__and3b_1.pex.spice
* Created: Fri Aug 28 17:12:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__AND3B_1%A_N 3 7 9 12 13 14 15 16 20 21
r31 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.405
+ $Y=1.275 $X2=0.405 $Y2=1.275
r32 15 16 9.58211 $w=4.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.347 $Y=1.295
+ $X2=0.347 $Y2=1.665
r33 15 21 0.517952 $w=4.43e-07 $l=2e-08 $layer=LI1_cond $X=0.347 $Y=1.295
+ $X2=0.347 $Y2=1.275
r34 13 14 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=0.495 $Y=1.78
+ $X2=0.495 $Y2=1.94
r35 12 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.405 $Y=1.615
+ $X2=0.405 $Y2=1.275
r36 12 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.405 $Y=1.615
+ $X2=0.405 $Y2=1.78
r37 11 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.405 $Y=1.11
+ $X2=0.405 $Y2=1.275
r38 7 14 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.51 $Y=2.03 $X2=0.51
+ $Y2=1.94
r39 7 9 136.567 $w=1.8e-07 $l=5.1e-07 $layer=POLY_cond $X=0.51 $Y=2.03 $X2=0.51
+ $Y2=2.54
r40 3 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.495 $Y=0.645
+ $X2=0.495 $Y2=1.11
.ends

.subckt PM_SKY130_FD_SC_MS__AND3B_1%A_114_74# 1 2 9 13 15 17 18 21 25 27 28 33
+ 34 35
c66 33 0 7.864e-20 $X=0.975 $Y=1.195
r67 34 35 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=0.86 $Y=2.1 $X2=0.86
+ $Y2=1.7
r68 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.975
+ $Y=1.195 $X2=0.975 $Y2=1.195
r69 28 35 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=0.957 $Y=1.518
+ $X2=0.957 $Y2=1.7
r70 27 32 0.870046 $w=3.65e-07 $l=8.80909e-08 $layer=LI1_cond $X=0.957 $Y=1.212
+ $X2=0.877 $Y2=1.195
r71 27 28 9.66158 $w=3.63e-07 $l=3.06e-07 $layer=LI1_cond $X=0.957 $Y=1.212
+ $X2=0.957 $Y2=1.518
r72 25 34 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.78 $Y=2.265
+ $X2=0.78 $Y2=2.1
r73 19 32 15.5822 $w=3.3e-07 $l=4.65983e-07 $layer=LI1_cond $X=0.78 $Y=0.775
+ $X2=0.877 $Y2=1.195
r74 19 21 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.78 $Y=0.775
+ $X2=0.78 $Y2=0.645
r75 15 18 18.8402 $w=1.65e-07 $l=8e-08 $layer=POLY_cond $X=1.69 $Y=1.185
+ $X2=1.61 $Y2=1.185
r76 15 17 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.69 $Y=1.185
+ $X2=1.69 $Y2=0.79
r77 11 18 18.8402 $w=1.65e-07 $l=2.81425e-07 $layer=POLY_cond $X=1.7 $Y=1.425
+ $X2=1.61 $Y2=1.185
r78 11 13 324.573 $w=1.8e-07 $l=8.35e-07 $layer=POLY_cond $X=1.7 $Y=1.425
+ $X2=1.7 $Y2=2.26
r79 10 33 19.7453 $w=1.5e-07 $l=2.00237e-07 $layer=POLY_cond $X=1.14 $Y=1.26
+ $X2=0.975 $Y2=1.182
r80 9 18 6.66866 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.61 $Y=1.26 $X2=1.61
+ $Y2=1.185
r81 9 10 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.61 $Y=1.26 $X2=1.14
+ $Y2=1.26
r82 2 25 300 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=2 $X=0.6
+ $Y=2.12 $X2=0.78 $Y2=2.265
r83 1 21 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.645
.ends

.subckt PM_SKY130_FD_SC_MS__AND3B_1%B 3 7 9 12 13
c36 13 0 1.10133e-19 $X=2.17 $Y=1.515
r37 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=1.515
+ $X2=2.17 $Y2=1.68
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=1.515
+ $X2=2.17 $Y2=1.35
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.17
+ $Y=1.515 $X2=2.17 $Y2=1.515
r40 9 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.17 $Y=1.665
+ $X2=2.17 $Y2=1.515
r41 7 15 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=2.245 $Y=2.26
+ $X2=2.245 $Y2=1.68
r42 3 14 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.08 $Y=0.79 $X2=2.08
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__AND3B_1%C 3 7 9 12 13
c34 12 0 1.69717e-19 $X=2.71 $Y=1.515
c35 7 0 1.10133e-19 $X=2.7 $Y=2.26
c36 3 0 4.57304e-20 $X=2.62 $Y=0.79
r37 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.515
+ $X2=2.71 $Y2=1.68
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.515
+ $X2=2.71 $Y2=1.35
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.71
+ $Y=1.515 $X2=2.71 $Y2=1.515
r40 9 13 4.93904 $w=3.48e-07 $l=1.5e-07 $layer=LI1_cond $X=2.7 $Y=1.665 $X2=2.7
+ $Y2=1.515
r41 7 15 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=2.7 $Y=2.26 $X2=2.7
+ $Y2=1.68
r42 3 14 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.62 $Y=0.79 $X2=2.62
+ $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__AND3B_1%A_266_94# 1 2 3 12 16 20 23 26 28 32 34 36
+ 40
c94 40 0 3.95737e-20 $X=3.25 $Y=1.465
c95 20 0 7.864e-20 $X=1.475 $Y=0.615
r96 40 43 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=1.465
+ $X2=3.25 $Y2=1.63
r97 40 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=1.465
+ $X2=3.25 $Y2=1.3
r98 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.25
+ $Y=1.465 $X2=3.25 $Y2=1.465
r99 29 34 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.64 $Y=2.035
+ $X2=1.475 $Y2=2.035
r100 28 36 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.31 $Y=2.035
+ $X2=2.475 $Y2=2.035
r101 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.31 $Y=2.035
+ $X2=1.64 $Y2=2.035
r102 27 32 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.64 $Y=1.135
+ $X2=1.475 $Y2=1.135
r103 26 39 14.2261 $w=2.83e-07 $l=4.1225e-07 $layer=LI1_cond $X=3.045 $Y=1.135
+ $X2=3.23 $Y2=1.465
r104 26 27 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=3.045 $Y=1.135
+ $X2=1.64 $Y2=1.135
r105 23 34 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.475 $Y=1.95
+ $X2=1.475 $Y2=2.035
r106 22 32 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.475 $Y=1.22
+ $X2=1.475 $Y2=1.135
r107 22 23 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=1.475 $Y=1.22
+ $X2=1.475 $Y2=1.95
r108 18 32 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.475 $Y=1.05
+ $X2=1.475 $Y2=1.135
r109 18 20 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=1.475 $Y=1.05
+ $X2=1.475 $Y2=0.615
r110 16 42 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.335 $Y=0.74
+ $X2=3.335 $Y2=1.3
r111 12 43 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=3.285 $Y=2.4
+ $X2=3.285 $Y2=1.63
r112 3 36 300 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=2 $X=2.335
+ $Y=1.84 $X2=2.475 $Y2=2.115
r113 2 34 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.33
+ $Y=1.84 $X2=1.475 $Y2=1.985
r114 1 20 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.33
+ $Y=0.47 $X2=1.475 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__AND3B_1%VPWR 1 2 3 10 12 16 20 23 24 26 27 28 41 42
c46 20 0 1.69717e-19 $X=3.01 $Y=2.115
r47 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r49 39 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r50 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 33 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r54 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r55 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 30 45 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r57 30 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 28 39 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 28 36 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 26 38 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=3.01 $Y2=3.33
r62 25 41 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.175 $Y=3.33
+ $X2=3.6 $Y2=3.33
r63 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.175 $Y=3.33
+ $X2=3.01 $Y2=3.33
r64 23 35 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.81 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.81 $Y=3.33
+ $X2=1.975 $Y2=3.33
r66 22 38 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.14 $Y=3.33 $X2=2.64
+ $Y2=3.33
r67 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.14 $Y=3.33
+ $X2=1.975 $Y2=3.33
r68 18 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.01 $Y=3.245
+ $X2=3.01 $Y2=3.33
r69 18 20 39.4624 $w=3.28e-07 $l=1.13e-06 $layer=LI1_cond $X=3.01 $Y=3.245
+ $X2=3.01 $Y2=2.115
r70 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.975 $Y=3.245
+ $X2=1.975 $Y2=3.33
r71 14 16 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.975 $Y=3.245
+ $X2=1.975 $Y2=2.455
r72 10 45 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r73 10 12 34.2241 $w=3.28e-07 $l=9.8e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.265
r74 3 20 300 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_PDIFF $count=2 $X=2.79
+ $Y=1.84 $X2=3.01 $Y2=2.115
r75 2 16 600 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=1 $X=1.79
+ $Y=1.84 $X2=1.975 $Y2=2.455
r76 1 12 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.265
.ends

.subckt PM_SKY130_FD_SC_MS__AND3B_1%X 1 2 9 13 14 15 16 23 33 34
c25 13 0 8.53041e-20 $X=3.57 $Y=1.13
r26 33 34 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=3.55 $Y=1.985
+ $X2=3.55 $Y2=1.82
r27 21 23 0.281084 $w=4.08e-07 $l=1e-08 $layer=LI1_cond $X=3.55 $Y=2.025
+ $X2=3.55 $Y2=2.035
r28 16 30 1.12433 $w=4.08e-07 $l=4e-08 $layer=LI1_cond $X=3.55 $Y=2.775 $X2=3.55
+ $Y2=2.815
r29 15 16 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=3.55 $Y=2.405
+ $X2=3.55 $Y2=2.775
r30 14 21 1.06812 $w=4.08e-07 $l=3.8e-08 $layer=LI1_cond $X=3.55 $Y=1.987
+ $X2=3.55 $Y2=2.025
r31 14 33 0.0562167 $w=4.08e-07 $l=2e-09 $layer=LI1_cond $X=3.55 $Y=1.987
+ $X2=3.55 $Y2=1.985
r32 14 15 9.36009 $w=4.08e-07 $l=3.33e-07 $layer=LI1_cond $X=3.55 $Y=2.072
+ $X2=3.55 $Y2=2.405
r33 14 23 1.04001 $w=4.08e-07 $l=3.7e-08 $layer=LI1_cond $X=3.55 $Y=2.072
+ $X2=3.55 $Y2=2.035
r34 13 34 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.67 $Y=1.13 $X2=3.67
+ $Y2=1.82
r35 7 13 9.16175 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.57 $Y=0.945
+ $X2=3.57 $Y2=1.13
r36 7 9 13.3933 $w=3.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.57 $Y=0.945 $X2=3.57
+ $Y2=0.515
r37 2 33 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.375
+ $Y=1.84 $X2=3.51 $Y2=1.985
r38 2 30 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.375
+ $Y=1.84 $X2=3.51 $Y2=2.815
r39 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.41
+ $Y=0.37 $X2=3.55 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__AND3B_1%VGND 1 2 7 9 13 15 17 24 25 31
r35 32 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r36 31 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r37 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r38 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r39 25 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r40 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r41 22 31 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=3.215 $Y=0 $X2=2.92
+ $Y2=0
r42 22 24 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.215 $Y=0 $X2=3.6
+ $Y2=0
r43 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r44 20 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r45 18 28 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r46 18 20 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r47 17 31 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=2.625 $Y=0 $X2=2.92
+ $Y2=0
r48 17 20 124.283 $w=1.68e-07 $l=1.905e-06 $layer=LI1_cond $X=2.625 $Y=0
+ $X2=0.72 $Y2=0
r49 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r50 15 21 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=0.72
+ $Y2=0
r51 11 31 2.48142 $w=5.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.92 $Y=0.085
+ $X2=2.92 $Y2=0
r52 11 13 8.31173 $w=5.88e-07 $l=4.1e-07 $layer=LI1_cond $X=2.92 $Y=0.085
+ $X2=2.92 $Y2=0.495
r53 7 28 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r54 7 9 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.28 $Y=0.085 $X2=0.28
+ $Y2=0.645
r55 2 13 91 $w=1.7e-07 $l=4.37321e-07 $layer=licon1_NDIFF $count=2 $X=2.695
+ $Y=0.47 $X2=3.12 $Y2=0.495
r56 1 9 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.645
.ends


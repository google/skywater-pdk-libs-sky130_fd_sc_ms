* File: sky130_fd_sc_ms__a2111oi_1.pxi.spice
* Created: Wed Sep  2 11:49:40 2020
* 
x_PM_SKY130_FD_SC_MS__A2111OI_1%D1 N_D1_M1007_g N_D1_M1003_g D1 N_D1_c_60_n
+ N_D1_c_61_n PM_SKY130_FD_SC_MS__A2111OI_1%D1
x_PM_SKY130_FD_SC_MS__A2111OI_1%C1 N_C1_M1004_g N_C1_M1006_g C1 N_C1_c_88_n
+ N_C1_c_89_n PM_SKY130_FD_SC_MS__A2111OI_1%C1
x_PM_SKY130_FD_SC_MS__A2111OI_1%B1 N_B1_M1005_g N_B1_M1009_g B1 N_B1_c_125_n
+ N_B1_c_126_n PM_SKY130_FD_SC_MS__A2111OI_1%B1
x_PM_SKY130_FD_SC_MS__A2111OI_1%A1 N_A1_M1008_g N_A1_M1002_g A1 N_A1_c_162_n
+ N_A1_c_163_n PM_SKY130_FD_SC_MS__A2111OI_1%A1
x_PM_SKY130_FD_SC_MS__A2111OI_1%A2 N_A2_M1001_g N_A2_M1000_g A2 N_A2_c_201_n
+ N_A2_c_202_n PM_SKY130_FD_SC_MS__A2111OI_1%A2
x_PM_SKY130_FD_SC_MS__A2111OI_1%Y N_Y_M1003_d N_Y_M1009_d N_Y_M1007_s
+ N_Y_c_228_n N_Y_c_229_n N_Y_c_230_n N_Y_c_231_n N_Y_c_232_n N_Y_c_233_n
+ N_Y_c_234_n Y Y Y PM_SKY130_FD_SC_MS__A2111OI_1%Y
x_PM_SKY130_FD_SC_MS__A2111OI_1%A_345_368# N_A_345_368#_M1005_d
+ N_A_345_368#_M1000_d N_A_345_368#_c_295_n N_A_345_368#_c_291_n
+ N_A_345_368#_c_300_n N_A_345_368#_c_292_n N_A_345_368#_c_293_n
+ PM_SKY130_FD_SC_MS__A2111OI_1%A_345_368#
x_PM_SKY130_FD_SC_MS__A2111OI_1%VPWR N_VPWR_M1008_d N_VPWR_c_322_n
+ N_VPWR_c_323_n N_VPWR_c_324_n VPWR N_VPWR_c_325_n N_VPWR_c_321_n
+ PM_SKY130_FD_SC_MS__A2111OI_1%VPWR
x_PM_SKY130_FD_SC_MS__A2111OI_1%VGND N_VGND_M1003_s N_VGND_M1006_d
+ N_VGND_M1001_d N_VGND_c_350_n N_VGND_c_351_n N_VGND_c_352_n N_VGND_c_353_n
+ N_VGND_c_354_n N_VGND_c_355_n N_VGND_c_356_n N_VGND_c_357_n N_VGND_c_358_n
+ N_VGND_c_359_n VGND N_VGND_c_360_n PM_SKY130_FD_SC_MS__A2111OI_1%VGND
cc_1 VNB N_D1_M1003_g 0.0273265f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_2 VNB N_D1_c_60_n 0.0266188f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_3 VNB N_D1_c_61_n 0.00391874f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_4 VNB N_C1_M1006_g 0.0266005f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_5 VNB N_C1_c_88_n 0.0262274f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_6 VNB N_C1_c_89_n 0.00165719f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_7 VNB N_B1_M1009_g 0.026609f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_8 VNB N_B1_c_125_n 0.0262505f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_9 VNB N_B1_c_126_n 0.00166777f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_10 VNB N_A1_M1002_g 0.0250188f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_11 VNB N_A1_c_162_n 0.0242859f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_12 VNB N_A1_c_163_n 0.00709957f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_13 VNB N_A2_M1000_g 0.00909003f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_14 VNB A2 0.0349068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_c_201_n 0.0339369f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_16 VNB N_A2_c_202_n 0.0215297f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_17 VNB N_Y_c_228_n 0.0230393f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_18 VNB N_Y_c_229_n 0.0103726f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_19 VNB N_Y_c_230_n 0.0149129f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_20 VNB N_Y_c_231_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.515
cc_21 VNB N_Y_c_232_n 0.0170798f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.665
cc_22 VNB N_Y_c_233_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_234_n 0.00677638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_321_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_350_n 0.0279165f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.515
cc_26 VNB N_VGND_c_351_n 0.00974487f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.515
cc_27 VNB N_VGND_c_352_n 0.0344702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_353_n 0.0129628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_354_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_355_n 0.0169342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_356_n 0.00788625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_357_n 0.0110534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_358_n 0.0312656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_359_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_360_n 0.227536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_D1_M1007_g 0.0257165f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=2.4
cc_37 VPB N_D1_c_60_n 0.00564702f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_38 VPB N_D1_c_61_n 0.00341338f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_39 VPB N_C1_M1004_g 0.021884f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=2.4
cc_40 VPB N_C1_c_88_n 0.00562174f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_41 VPB N_C1_c_89_n 0.00260491f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_42 VPB N_B1_M1005_g 0.0236455f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=2.4
cc_43 VPB N_B1_c_125_n 0.00561631f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_44 VPB N_B1_c_126_n 0.00200497f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_45 VPB N_A1_M1008_g 0.0222921f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=2.4
cc_46 VPB N_A1_c_162_n 0.00549634f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_47 VPB N_A1_c_163_n 0.0036192f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_48 VPB N_A2_M1000_g 0.0326315f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_49 VPB N_Y_c_228_n 0.0148016f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_50 VPB Y 0.0609165f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A_345_368#_c_291_n 0.00312968f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_52 VPB N_A_345_368#_c_292_n 0.0150854f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.515
cc_53 VPB N_A_345_368#_c_293_n 0.0358769f $X=-0.19 $Y=1.66 $X2=0.63 $Y2=1.68
cc_54 VPB N_VPWR_c_322_n 0.0067963f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_55 VPB N_VPWR_c_323_n 0.0609497f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_56 VPB N_VPWR_c_324_n 0.00689679f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_325_n 0.0236066f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_321_n 0.0739275f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 N_D1_M1007_g N_C1_M1004_g 0.0559772f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_60 N_D1_M1003_g N_C1_M1006_g 0.0195038f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_61 N_D1_c_60_n N_C1_c_88_n 0.0559772f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_62 N_D1_c_61_n N_C1_c_88_n 0.00240981f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_63 N_D1_c_60_n N_C1_c_89_n 4.95839e-19 $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_64 N_D1_c_61_n N_C1_c_89_n 0.0343047f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_65 N_D1_M1007_g N_Y_c_228_n 0.00390285f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_66 N_D1_M1003_g N_Y_c_228_n 0.00477786f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_67 N_D1_c_60_n N_Y_c_228_n 0.00739878f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_68 N_D1_c_61_n N_Y_c_228_n 0.0330212f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_69 N_D1_M1003_g N_Y_c_229_n 0.0148724f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_70 N_D1_c_60_n N_Y_c_229_n 0.00125903f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_71 N_D1_c_61_n N_Y_c_229_n 0.0279704f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_72 N_D1_M1003_g N_Y_c_231_n 3.97481e-19 $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_73 N_D1_M1007_g Y 0.0314572f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_74 N_D1_c_60_n Y 7.737e-19 $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_75 N_D1_c_61_n Y 0.0269275f $X=0.63 $Y=1.515 $X2=0 $Y2=0
cc_76 N_D1_M1007_g N_VPWR_c_323_n 0.00349978f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_77 N_D1_M1007_g N_VPWR_c_321_n 0.00433289f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_78 N_D1_M1003_g N_VGND_c_350_n 0.0127749f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_79 N_D1_M1003_g N_VGND_c_355_n 0.00383152f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_80 N_D1_M1003_g N_VGND_c_360_n 0.00757637f $X=0.72 $Y=0.74 $X2=0 $Y2=0
cc_81 N_C1_M1004_g N_B1_M1005_g 0.0448865f $X=1.095 $Y=2.4 $X2=0 $Y2=0
cc_82 N_C1_c_89_n N_B1_M1005_g 6.85212e-19 $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_83 N_C1_M1006_g N_B1_M1009_g 0.0204655f $X=1.15 $Y=0.74 $X2=0 $Y2=0
cc_84 N_C1_c_88_n N_B1_c_125_n 0.0201104f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_85 N_C1_c_89_n N_B1_c_125_n 0.00114936f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_86 N_C1_c_88_n N_B1_c_126_n 0.00114936f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_87 N_C1_c_89_n N_B1_c_126_n 0.0276388f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_88 N_C1_M1006_g N_Y_c_231_n 0.00959601f $X=1.15 $Y=0.74 $X2=0 $Y2=0
cc_89 N_C1_M1006_g N_Y_c_232_n 0.01209f $X=1.15 $Y=0.74 $X2=0 $Y2=0
cc_90 N_C1_c_88_n N_Y_c_232_n 7.68393e-19 $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_91 N_C1_c_89_n N_Y_c_232_n 0.0175347f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_92 N_C1_M1006_g N_Y_c_233_n 8.21695e-19 $X=1.15 $Y=0.74 $X2=0 $Y2=0
cc_93 N_C1_M1006_g N_Y_c_234_n 0.0015571f $X=1.15 $Y=0.74 $X2=0 $Y2=0
cc_94 N_C1_c_88_n N_Y_c_234_n 5.39598e-19 $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_95 N_C1_c_89_n N_Y_c_234_n 0.00799991f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_96 N_C1_M1004_g Y 0.0399063f $X=1.095 $Y=2.4 $X2=0 $Y2=0
cc_97 N_C1_c_88_n Y 6.54022e-19 $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_98 N_C1_c_89_n Y 0.0235098f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_99 N_C1_M1004_g N_A_345_368#_c_291_n 7.59934e-19 $X=1.095 $Y=2.4 $X2=0 $Y2=0
cc_100 N_C1_M1004_g N_VPWR_c_323_n 0.00349978f $X=1.095 $Y=2.4 $X2=0 $Y2=0
cc_101 N_C1_M1004_g N_VPWR_c_321_n 0.00429927f $X=1.095 $Y=2.4 $X2=0 $Y2=0
cc_102 N_C1_M1006_g N_VGND_c_350_n 5.17822e-19 $X=1.15 $Y=0.74 $X2=0 $Y2=0
cc_103 N_C1_M1006_g N_VGND_c_351_n 0.0053617f $X=1.15 $Y=0.74 $X2=0 $Y2=0
cc_104 N_C1_M1006_g N_VGND_c_355_n 0.00434272f $X=1.15 $Y=0.74 $X2=0 $Y2=0
cc_105 N_C1_M1006_g N_VGND_c_360_n 0.00821949f $X=1.15 $Y=0.74 $X2=0 $Y2=0
cc_106 N_B1_M1005_g N_A1_M1008_g 0.0258538f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_107 N_B1_c_126_n N_A1_M1008_g 3.38956e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_108 N_B1_M1009_g N_A1_M1002_g 0.0204481f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_109 N_B1_c_125_n N_A1_c_162_n 0.0206294f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_110 N_B1_c_126_n N_A1_c_162_n 3.80681e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_111 N_B1_M1005_g N_A1_c_163_n 2.6794e-19 $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_112 N_B1_c_125_n N_A1_c_163_n 0.00188197f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_113 N_B1_c_126_n N_A1_c_163_n 0.0347534f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_114 N_B1_M1009_g N_Y_c_231_n 8.24465e-19 $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_115 N_B1_M1009_g N_Y_c_232_n 0.0136326f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_116 N_B1_c_125_n N_Y_c_232_n 0.001245f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_117 N_B1_c_126_n N_Y_c_232_n 0.0248933f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_118 N_B1_M1009_g N_Y_c_233_n 0.00990712f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_119 N_B1_M1005_g Y 0.00974182f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_120 N_B1_M1005_g N_A_345_368#_c_295_n 0.00314634f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_121 N_B1_c_125_n N_A_345_368#_c_295_n 7.63688e-19 $X=1.71 $Y=1.515 $X2=0
+ $Y2=0
cc_122 N_B1_c_126_n N_A_345_368#_c_295_n 0.0130747f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_123 N_B1_M1005_g N_A_345_368#_c_291_n 0.014451f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_124 N_B1_M1005_g N_VPWR_c_322_n 6.73475e-19 $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_125 N_B1_M1005_g N_VPWR_c_323_n 0.005209f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_126 N_B1_M1005_g N_VPWR_c_321_n 0.00985168f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_127 N_B1_M1009_g N_VGND_c_351_n 0.00690689f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_128 N_B1_M1009_g N_VGND_c_358_n 0.00434272f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_129 N_B1_M1009_g N_VGND_c_360_n 0.00821949f $X=1.8 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A1_M1008_g N_A2_M1000_g 0.0312909f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_131 N_A1_c_163_n N_A2_M1000_g 0.00238858f $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_132 N_A1_M1002_g A2 0.00101508f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A1_c_162_n A2 6.92182e-19 $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_134 N_A1_c_163_n A2 0.013398f $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_135 N_A1_c_162_n N_A2_c_201_n 0.0210016f $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_136 N_A1_c_163_n N_A2_c_201_n 0.00113385f $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_137 N_A1_M1002_g N_A2_c_202_n 0.039902f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_138 N_A1_M1002_g N_Y_c_232_n 0.00464229f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A1_c_162_n N_Y_c_232_n 5.47418e-19 $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_140 N_A1_c_163_n N_Y_c_232_n 0.0116188f $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_141 N_A1_M1002_g N_Y_c_233_n 0.0132273f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_142 N_A1_M1008_g N_A_345_368#_c_291_n 0.00510762f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_143 N_A1_M1008_g N_A_345_368#_c_300_n 0.0171681f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A1_c_162_n N_A_345_368#_c_300_n 7.05813e-19 $X=2.25 $Y=1.515 $X2=0
+ $Y2=0
cc_145 N_A1_c_163_n N_A_345_368#_c_300_n 0.0239159f $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_146 N_A1_M1008_g N_A_345_368#_c_292_n 5.99214e-19 $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_147 N_A1_M1008_g N_A_345_368#_c_293_n 7.67392e-19 $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_148 N_A1_M1008_g N_VPWR_c_322_n 0.012948f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_149 N_A1_M1008_g N_VPWR_c_323_n 0.00460063f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_150 N_A1_M1008_g N_VPWR_c_321_n 0.00909457f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_151 N_A1_M1002_g N_VGND_c_352_n 0.00253715f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_152 N_A1_M1002_g N_VGND_c_358_n 0.00434272f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_153 N_A1_M1002_g N_VGND_c_360_n 0.00821825f $X=2.23 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A2_c_202_n N_Y_c_232_n 8.07707e-19 $X=2.79 $Y=1.22 $X2=0 $Y2=0
cc_155 N_A2_c_202_n N_Y_c_233_n 0.0019967f $X=2.79 $Y=1.22 $X2=0 $Y2=0
cc_156 N_A2_M1000_g N_A_345_368#_c_300_n 0.0146034f $X=2.715 $Y=2.4 $X2=0 $Y2=0
cc_157 A2 N_A_345_368#_c_300_n 0.00540887f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_158 N_A2_M1000_g N_A_345_368#_c_292_n 0.00407495f $X=2.715 $Y=2.4 $X2=0 $Y2=0
cc_159 A2 N_A_345_368#_c_292_n 0.0203808f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_160 N_A2_c_201_n N_A_345_368#_c_292_n 0.00330449f $X=2.79 $Y=1.385 $X2=0
+ $Y2=0
cc_161 N_A2_M1000_g N_A_345_368#_c_293_n 0.0129517f $X=2.715 $Y=2.4 $X2=0 $Y2=0
cc_162 N_A2_M1000_g N_VPWR_c_322_n 0.00741529f $X=2.715 $Y=2.4 $X2=0 $Y2=0
cc_163 N_A2_M1000_g N_VPWR_c_325_n 0.005209f $X=2.715 $Y=2.4 $X2=0 $Y2=0
cc_164 N_A2_M1000_g N_VPWR_c_321_n 0.00986635f $X=2.715 $Y=2.4 $X2=0 $Y2=0
cc_165 A2 N_VGND_c_352_n 0.0259407f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_166 N_A2_c_201_n N_VGND_c_352_n 0.0011179f $X=2.79 $Y=1.385 $X2=0 $Y2=0
cc_167 N_A2_c_202_n N_VGND_c_352_n 0.0176088f $X=2.79 $Y=1.22 $X2=0 $Y2=0
cc_168 N_A2_c_202_n N_VGND_c_358_n 0.00383152f $X=2.79 $Y=1.22 $X2=0 $Y2=0
cc_169 N_A2_c_202_n N_VGND_c_360_n 0.00757998f $X=2.79 $Y=1.22 $X2=0 $Y2=0
cc_170 Y A_159_368# 0.00433061f $X=1.115 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_171 Y A_237_368# 0.0132769f $X=1.115 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_172 Y N_A_345_368#_c_295_n 0.00791938f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_173 Y N_A_345_368#_c_291_n 0.0384991f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_174 Y N_VPWR_c_323_n 0.0517721f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_175 Y N_VPWR_c_321_n 0.0421749f $X=1.115 $Y=2.32 $X2=0 $Y2=0
cc_176 N_Y_c_229_n N_VGND_M1003_s 0.00267685f $X=0.85 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_177 N_Y_c_232_n N_VGND_M1006_d 0.00487041f $X=1.85 $Y=1.095 $X2=0 $Y2=0
cc_178 N_Y_c_229_n N_VGND_c_350_n 0.0220026f $X=0.85 $Y=1.095 $X2=0 $Y2=0
cc_179 N_Y_c_231_n N_VGND_c_350_n 0.0182902f $X=0.935 $Y=0.515 $X2=0 $Y2=0
cc_180 N_Y_c_231_n N_VGND_c_351_n 0.018437f $X=0.935 $Y=0.515 $X2=0 $Y2=0
cc_181 N_Y_c_232_n N_VGND_c_351_n 0.0314044f $X=1.85 $Y=1.095 $X2=0 $Y2=0
cc_182 N_Y_c_233_n N_VGND_c_351_n 0.0192028f $X=2.015 $Y=0.515 $X2=0 $Y2=0
cc_183 N_Y_c_233_n N_VGND_c_352_n 0.018269f $X=2.015 $Y=0.515 $X2=0 $Y2=0
cc_184 N_Y_c_231_n N_VGND_c_355_n 0.0109942f $X=0.935 $Y=0.515 $X2=0 $Y2=0
cc_185 N_Y_c_233_n N_VGND_c_358_n 0.0144922f $X=2.015 $Y=0.515 $X2=0 $Y2=0
cc_186 N_Y_c_231_n N_VGND_c_360_n 0.00904371f $X=0.935 $Y=0.515 $X2=0 $Y2=0
cc_187 N_Y_c_233_n N_VGND_c_360_n 0.0118826f $X=2.015 $Y=0.515 $X2=0 $Y2=0
cc_188 N_A_345_368#_c_300_n N_VPWR_M1008_d 0.00928873f $X=2.775 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_189 N_A_345_368#_c_291_n N_VPWR_c_322_n 0.0271521f $X=1.88 $Y=2.435 $X2=0
+ $Y2=0
cc_190 N_A_345_368#_c_300_n N_VPWR_c_322_n 0.0221812f $X=2.775 $Y=2.035 $X2=0
+ $Y2=0
cc_191 N_A_345_368#_c_293_n N_VPWR_c_322_n 0.0266947f $X=2.94 $Y=2.815 $X2=0
+ $Y2=0
cc_192 N_A_345_368#_c_291_n N_VPWR_c_323_n 0.0163338f $X=1.88 $Y=2.435 $X2=0
+ $Y2=0
cc_193 N_A_345_368#_c_293_n N_VPWR_c_325_n 0.014549f $X=2.94 $Y=2.815 $X2=0
+ $Y2=0
cc_194 N_A_345_368#_c_291_n N_VPWR_c_321_n 0.0134516f $X=1.88 $Y=2.435 $X2=0
+ $Y2=0
cc_195 N_A_345_368#_c_293_n N_VPWR_c_321_n 0.0119743f $X=2.94 $Y=2.815 $X2=0
+ $Y2=0

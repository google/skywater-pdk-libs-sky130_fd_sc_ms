* File: sky130_fd_sc_ms__and4b_4.pxi.spice
* Created: Fri Aug 28 17:14:16 2020
* 
x_PM_SKY130_FD_SC_MS__AND4B_4%A_N N_A_N_M1004_g N_A_N_M1011_g A_N N_A_N_c_145_n
+ N_A_N_c_146_n PM_SKY130_FD_SC_MS__AND4B_4%A_N
x_PM_SKY130_FD_SC_MS__AND4B_4%A_199_294# N_A_199_294#_M1013_s
+ N_A_199_294#_M1010_d N_A_199_294#_M1020_d N_A_199_294#_M1006_d
+ N_A_199_294#_M1012_s N_A_199_294#_M1001_g N_A_199_294#_M1005_g
+ N_A_199_294#_M1009_g N_A_199_294#_M1014_g N_A_199_294#_M1015_g
+ N_A_199_294#_M1022_g N_A_199_294#_M1017_g N_A_199_294#_M1025_g
+ N_A_199_294#_c_186_n N_A_199_294#_c_187_n N_A_199_294#_c_196_n
+ N_A_199_294#_c_197_n N_A_199_294#_c_247_p N_A_199_294#_c_188_n
+ N_A_199_294#_c_189_n N_A_199_294#_c_230_p N_A_199_294#_c_199_n
+ N_A_199_294#_c_208_p N_A_199_294#_c_200_n N_A_199_294#_c_190_n
+ N_A_199_294#_c_191_n PM_SKY130_FD_SC_MS__AND4B_4%A_199_294#
x_PM_SKY130_FD_SC_MS__AND4B_4%D N_D_M1003_g N_D_c_337_n N_D_c_338_n N_D_M1020_g
+ N_D_c_339_n N_D_M1007_g N_D_c_340_n N_D_M1021_g D D D N_D_c_342_n
+ PM_SKY130_FD_SC_MS__AND4B_4%D
x_PM_SKY130_FD_SC_MS__AND4B_4%C N_C_M1010_g N_C_c_396_n N_C_c_397_n N_C_M1000_g
+ N_C_c_399_n N_C_c_408_n N_C_M1024_g N_C_M1016_g N_C_c_401_n N_C_c_402_n
+ N_C_c_403_n C N_C_c_404_n N_C_c_405_n N_C_c_406_n
+ PM_SKY130_FD_SC_MS__AND4B_4%C
x_PM_SKY130_FD_SC_MS__AND4B_4%A_27_368# N_A_27_368#_M1011_s N_A_27_368#_M1004_s
+ N_A_27_368#_M1008_g N_A_27_368#_M1013_g N_A_27_368#_M1023_g
+ N_A_27_368#_M1012_g N_A_27_368#_c_483_n N_A_27_368#_c_493_n
+ N_A_27_368#_c_502_n N_A_27_368#_c_484_n N_A_27_368#_c_485_n
+ N_A_27_368#_c_530_n N_A_27_368#_c_486_n N_A_27_368#_c_487_n
+ N_A_27_368#_c_495_n N_A_27_368#_c_488_n N_A_27_368#_c_497_n
+ N_A_27_368#_c_489_n N_A_27_368#_c_490_n PM_SKY130_FD_SC_MS__AND4B_4%A_27_368#
x_PM_SKY130_FD_SC_MS__AND4B_4%B N_B_c_614_n N_B_M1006_g N_B_M1002_g N_B_c_617_n
+ N_B_c_618_n N_B_M1018_g N_B_M1019_g B N_B_c_621_n
+ PM_SKY130_FD_SC_MS__AND4B_4%B
x_PM_SKY130_FD_SC_MS__AND4B_4%VPWR N_VPWR_M1004_d N_VPWR_M1014_d N_VPWR_M1017_d
+ N_VPWR_M1003_s N_VPWR_M1024_s N_VPWR_M1008_d N_VPWR_M1018_s N_VPWR_c_679_n
+ N_VPWR_c_680_n N_VPWR_c_681_n N_VPWR_c_682_n N_VPWR_c_683_n N_VPWR_c_684_n
+ N_VPWR_c_685_n N_VPWR_c_686_n N_VPWR_c_687_n N_VPWR_c_688_n N_VPWR_c_689_n
+ N_VPWR_c_690_n N_VPWR_c_691_n VPWR N_VPWR_c_692_n N_VPWR_c_693_n
+ N_VPWR_c_694_n N_VPWR_c_695_n N_VPWR_c_696_n N_VPWR_c_697_n N_VPWR_c_678_n
+ PM_SKY130_FD_SC_MS__AND4B_4%VPWR
x_PM_SKY130_FD_SC_MS__AND4B_4%X N_X_M1005_s N_X_M1022_s N_X_M1001_s N_X_M1015_s
+ N_X_c_777_n N_X_c_772_n N_X_c_773_n X X X X X N_X_c_776_n X N_X_c_785_n
+ PM_SKY130_FD_SC_MS__AND4B_4%X
x_PM_SKY130_FD_SC_MS__AND4B_4%VGND N_VGND_M1011_d N_VGND_M1009_d N_VGND_M1025_d
+ N_VGND_M1007_d N_VGND_c_834_n N_VGND_c_835_n N_VGND_c_836_n N_VGND_c_837_n
+ N_VGND_c_838_n N_VGND_c_839_n N_VGND_c_840_n VGND N_VGND_c_841_n
+ N_VGND_c_842_n N_VGND_c_843_n N_VGND_c_844_n N_VGND_c_845_n N_VGND_c_846_n
+ N_VGND_c_847_n PM_SKY130_FD_SC_MS__AND4B_4%VGND
x_PM_SKY130_FD_SC_MS__AND4B_4%A_664_125# N_A_664_125#_M1000_d
+ N_A_664_125#_M1016_d N_A_664_125#_M1019_d N_A_664_125#_c_917_n
+ N_A_664_125#_c_918_n N_A_664_125#_c_919_n N_A_664_125#_c_920_n
+ N_A_664_125#_c_921_n N_A_664_125#_c_922_n N_A_664_125#_c_923_n
+ PM_SKY130_FD_SC_MS__AND4B_4%A_664_125#
x_PM_SKY130_FD_SC_MS__AND4B_4%A_751_125# N_A_751_125#_M1000_s
+ N_A_751_125#_M1021_s N_A_751_125#_c_977_n N_A_751_125#_c_979_n
+ N_A_751_125#_c_976_n PM_SKY130_FD_SC_MS__AND4B_4%A_751_125#
x_PM_SKY130_FD_SC_MS__AND4B_4%A_1136_125# N_A_1136_125#_M1002_s
+ N_A_1136_125#_M1023_d N_A_1136_125#_c_1000_n N_A_1136_125#_c_1001_n
+ N_A_1136_125#_c_1002_n PM_SKY130_FD_SC_MS__AND4B_4%A_1136_125#
cc_1 VNB N_A_N_M1004_g 0.00709783f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.34
cc_2 VNB A_N 0.00916222f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_A_N_c_145_n 0.0378267f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_4 VNB N_A_N_c_146_n 0.0208794f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.22
cc_5 VNB N_A_199_294#_M1001_g 0.00549559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_199_294#_M1005_g 0.0226641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_199_294#_M1009_g 0.0241832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_199_294#_M1014_g 4.87684e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_199_294#_M1015_g 5.27393e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_199_294#_M1022_g 0.0242295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_199_294#_M1017_g 4.72639e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_199_294#_M1025_g 0.0242307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_199_294#_c_186_n 0.0109969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_199_294#_c_187_n 0.00444332f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_199_294#_c_188_n 0.00296626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_199_294#_c_189_n 0.00360386f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_199_294#_c_190_n 0.00926078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_199_294#_c_191_n 0.0682349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_D_c_337_n 0.00906242f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.22
cc_20 VNB N_D_c_338_n 0.0050671f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.79
cc_21 VNB N_D_c_339_n 0.0148233f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_22 VNB N_D_c_340_n 0.0142612f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.55
cc_23 VNB D 0.010589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_D_c_342_n 0.0488567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_C_c_396_n 0.0223825f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.79
cc_26 VNB N_C_c_397_n 0.0124252f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_27 VNB N_C_M1000_g 0.0328565f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_28 VNB N_C_c_399_n 0.103403f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.22
cc_29 VNB N_C_M1016_g 0.0253364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_C_c_401_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_C_c_402_n 0.00839426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_C_c_403_n 0.0106507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_C_c_404_n 0.0356178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_C_c_405_n 0.00341194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_C_c_406_n 0.0655029f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_27_368#_M1013_g 0.0185365f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.22
cc_37 VNB N_A_27_368#_M1023_g 0.0217497f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.37
cc_38 VNB N_A_27_368#_c_483_n 0.02003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_27_368#_c_484_n 0.00244208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_27_368#_c_485_n 0.0182741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_27_368#_c_486_n 0.0170197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_27_368#_c_487_n 0.00646723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_27_368#_c_488_n 0.0297812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_27_368#_c_489_n 0.00142009f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_27_368#_c_490_n 0.021375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_B_c_614_n 0.00670072f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.55
cc_47 VNB N_B_M1006_g 0.00994453f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.34
cc_48 VNB N_B_M1002_g 0.0292859f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_49 VNB N_B_c_617_n 0.104114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_B_c_618_n 0.00962308f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.385
cc_51 VNB N_B_M1019_g 0.0363835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB B 0.00124747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_B_c_621_n 0.0188293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VPWR_c_678_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_X_c_772_n 0.00596934f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.37
cc_56 VNB N_X_c_773_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB X 0.00172508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB X 0.00280128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_X_c_776_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_834_n 0.0106049f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.37
cc_61 VNB N_VGND_c_835_n 0.02097f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.37
cc_62 VNB N_VGND_c_836_n 0.00987337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_837_n 0.0247003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_838_n 0.0102202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_839_n 0.0199677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_840_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_841_n 0.018718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_842_n 0.0356343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_843_n 0.0762007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_844_n 0.402809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_845_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_846_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_847_n 0.0043699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_664_125#_c_917_n 0.00708785f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.385
cc_75 VNB N_A_664_125#_c_918_n 0.0128721f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.55
cc_76 VNB N_A_664_125#_c_919_n 0.00493612f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.37
cc_77 VNB N_A_664_125#_c_920_n 0.00385728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_664_125#_c_921_n 0.0382876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_664_125#_c_922_n 0.00335039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_664_125#_c_923_n 0.0213365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_751_125#_c_976_n 0.00273786f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.55
cc_82 VNB N_A_1136_125#_c_1000_n 0.00255783f $X=-0.19 $Y=-0.245 $X2=0.535
+ $Y2=0.79
cc_83 VNB N_A_1136_125#_c_1001_n 0.00157665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1136_125#_c_1002_n 0.00237075f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=1.55
cc_85 VPB N_A_N_M1004_g 0.0293989f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.34
cc_86 VPB N_A_199_294#_M1001_g 0.024148f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_87 VPB N_A_199_294#_M1014_g 0.0219554f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_A_199_294#_M1015_g 0.0232935f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_89 VPB N_A_199_294#_M1017_g 0.0234502f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_90 VPB N_A_199_294#_c_196_n 0.00139365f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_91 VPB N_A_199_294#_c_197_n 0.0058507f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_92 VPB N_A_199_294#_c_189_n 0.00292216f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_93 VPB N_A_199_294#_c_199_n 0.00332675f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_A_199_294#_c_200_n 0.00854879f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_D_M1003_g 0.0228164f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.34
cc_96 VPB N_D_c_337_n 0.00914673f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=1.22
cc_97 VPB N_D_c_338_n 0.00537756f $X=-0.19 $Y=1.66 $X2=0.535 $Y2=0.79
cc_98 VPB N_D_M1020_g 0.0305685f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_99 VPB D 0.00260186f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_100 VPB N_D_c_342_n 0.0268669f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_101 VPB N_C_M1010_g 0.0293432f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.34
cc_102 VPB N_C_c_408_n 0.00639802f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.37
cc_103 VPB N_C_M1024_g 0.027971f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.37
cc_104 VPB N_C_c_402_n 0.00370107f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_C_c_404_n 0.00565389f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_C_c_405_n 0.00310957f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_27_368#_M1008_g 0.0202546f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_27_368#_M1012_g 0.0212049f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_27_368#_c_493_n 0.0153183f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_27_368#_c_486_n 0.0146378f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_27_368#_c_495_n 0.0136968f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_112 VPB N_A_27_368#_c_488_n 0.00769959f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_27_368#_c_497_n 0.0220699f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_27_368#_c_489_n 0.00172979f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_27_368#_c_490_n 0.0151523f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_B_M1006_g 0.0296565f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.34
cc_117 VPB N_B_M1018_g 0.0245934f $X=-0.19 $Y=1.66 $X2=0.585 $Y2=1.22
cc_118 VPB B 9.29746e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_B_c_621_n 0.0158279f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_679_n 0.0107372f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_680_n 0.00329267f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_681_n 0.0212593f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_682_n 0.00666636f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_683_n 0.0065007f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_684_n 0.00329222f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_685_n 0.00261656f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_686_n 0.0234846f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_687_n 0.00612764f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_688_n 0.0355792f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_689_n 0.0063829f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_690_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_691_n 0.00601668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_692_n 0.0177589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_693_n 0.017758f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_694_n 0.0276117f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_695_n 0.00656601f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_696_n 0.00641618f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_697_n 0.0387911f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_678_n 0.0801449f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_X_c_777_n 0.00647524f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.37
cc_141 VPB X 0.00154535f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 A_N N_A_199_294#_M1005_g 0.00213771f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_143 N_A_N_c_145_n N_A_199_294#_M1005_g 0.0120427f $X=0.59 $Y=1.385 $X2=0
+ $Y2=0
cc_144 N_A_N_c_146_n N_A_199_294#_M1005_g 0.0135044f $X=0.585 $Y=1.22 $X2=0
+ $Y2=0
cc_145 N_A_N_M1004_g N_A_199_294#_c_186_n 0.036549f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_146 A_N N_A_199_294#_c_186_n 5.51989e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_147 N_A_N_c_145_n N_A_199_294#_c_186_n 0.00404495f $X=0.59 $Y=1.385 $X2=0
+ $Y2=0
cc_148 N_A_N_c_146_n N_A_27_368#_c_483_n 0.00351224f $X=0.585 $Y=1.22 $X2=0
+ $Y2=0
cc_149 N_A_N_M1004_g N_A_27_368#_c_493_n 0.00816745f $X=0.505 $Y=2.34 $X2=0
+ $Y2=0
cc_150 N_A_N_M1004_g N_A_27_368#_c_502_n 0.015266f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_151 N_A_N_M1004_g N_A_27_368#_c_495_n 0.00500536f $X=0.505 $Y=2.34 $X2=0
+ $Y2=0
cc_152 A_N N_A_27_368#_c_495_n 0.00105278f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_153 A_N N_A_27_368#_c_488_n 0.0276149f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_154 N_A_N_c_145_n N_A_27_368#_c_488_n 0.0152991f $X=0.59 $Y=1.385 $X2=0 $Y2=0
cc_155 N_A_N_c_146_n N_A_27_368#_c_488_n 0.00417267f $X=0.585 $Y=1.22 $X2=0
+ $Y2=0
cc_156 N_A_N_M1004_g N_A_27_368#_c_497_n 0.00694474f $X=0.505 $Y=2.34 $X2=0
+ $Y2=0
cc_157 N_A_N_M1004_g N_VPWR_c_679_n 0.00409896f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_158 N_A_N_M1004_g N_VPWR_c_694_n 0.00567889f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_159 N_A_N_M1004_g N_VPWR_c_678_n 0.00610055f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_160 N_A_N_c_146_n X 4.11144e-19 $X=0.585 $Y=1.22 $X2=0 $Y2=0
cc_161 N_A_N_M1004_g X 0.00134903f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_162 A_N X 0.0211453f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_163 N_A_N_c_145_n X 3.30789e-19 $X=0.59 $Y=1.385 $X2=0 $Y2=0
cc_164 N_A_N_c_146_n X 2.30211e-19 $X=0.585 $Y=1.22 $X2=0 $Y2=0
cc_165 N_A_N_c_146_n N_X_c_776_n 2.11176e-19 $X=0.585 $Y=1.22 $X2=0 $Y2=0
cc_166 N_A_N_M1004_g N_X_c_785_n 0.00136573f $X=0.505 $Y=2.34 $X2=0 $Y2=0
cc_167 A_N N_VGND_c_834_n 0.0189574f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_168 N_A_N_c_145_n N_VGND_c_834_n 8.95272e-19 $X=0.59 $Y=1.385 $X2=0 $Y2=0
cc_169 N_A_N_c_146_n N_VGND_c_834_n 0.0135392f $X=0.585 $Y=1.22 $X2=0 $Y2=0
cc_170 N_A_N_c_146_n N_VGND_c_841_n 0.00421418f $X=0.585 $Y=1.22 $X2=0 $Y2=0
cc_171 N_A_N_c_146_n N_VGND_c_844_n 0.00432128f $X=0.585 $Y=1.22 $X2=0 $Y2=0
cc_172 N_A_199_294#_c_199_n N_D_M1003_g 0.00228852f $X=3.515 $Y=2.085 $X2=0
+ $Y2=0
cc_173 N_A_199_294#_c_208_p N_D_M1003_g 0.012551f $X=5.65 $Y=2.08 $X2=0 $Y2=0
cc_174 N_A_199_294#_c_208_p N_D_c_337_n 0.00431842f $X=5.65 $Y=2.08 $X2=0 $Y2=0
cc_175 N_A_199_294#_c_208_p N_D_M1020_g 0.0127436f $X=5.65 $Y=2.08 $X2=0 $Y2=0
cc_176 N_A_199_294#_c_208_p D 0.0842095f $X=5.65 $Y=2.08 $X2=0 $Y2=0
cc_177 N_A_199_294#_c_208_p N_D_c_342_n 0.0141079f $X=5.65 $Y=2.08 $X2=0 $Y2=0
cc_178 N_A_199_294#_M1017_g N_C_M1010_g 0.0395801f $X=2.575 $Y=2.4 $X2=0 $Y2=0
cc_179 N_A_199_294#_c_196_n N_C_M1010_g 0.00343539f $X=2.66 $Y=1.95 $X2=0 $Y2=0
cc_180 N_A_199_294#_c_197_n N_C_M1010_g 0.0135117f $X=3.38 $Y=2.085 $X2=0 $Y2=0
cc_181 N_A_199_294#_M1025_g N_C_c_397_n 0.0116202f $X=2.59 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A_199_294#_c_208_p N_C_M1000_g 4.85856e-19 $X=5.65 $Y=2.08 $X2=0 $Y2=0
cc_183 N_A_199_294#_c_208_p N_C_M1024_g 0.0130036f $X=5.65 $Y=2.08 $X2=0 $Y2=0
cc_184 N_A_199_294#_c_187_n N_C_c_404_n 0.00199938f $X=2.575 $Y=1.485 $X2=0
+ $Y2=0
cc_185 N_A_199_294#_c_197_n N_C_c_404_n 8.33419e-19 $X=3.38 $Y=2.085 $X2=0 $Y2=0
cc_186 N_A_199_294#_c_191_n N_C_c_404_n 0.0165214f $X=2.59 $Y=1.485 $X2=0 $Y2=0
cc_187 N_A_199_294#_M1017_g N_C_c_405_n 3.10741e-19 $X=2.575 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A_199_294#_c_187_n N_C_c_405_n 0.0253f $X=2.575 $Y=1.485 $X2=0 $Y2=0
cc_189 N_A_199_294#_c_196_n N_C_c_405_n 0.010144f $X=2.66 $Y=1.95 $X2=0 $Y2=0
cc_190 N_A_199_294#_c_197_n N_C_c_405_n 0.0260984f $X=3.38 $Y=2.085 $X2=0 $Y2=0
cc_191 N_A_199_294#_c_191_n N_C_c_405_n 3.55661e-19 $X=2.59 $Y=1.485 $X2=0 $Y2=0
cc_192 N_A_199_294#_c_187_n N_C_c_406_n 7.00615e-19 $X=2.575 $Y=1.485 $X2=0
+ $Y2=0
cc_193 N_A_199_294#_c_191_n N_C_c_406_n 0.0116202f $X=2.59 $Y=1.485 $X2=0 $Y2=0
cc_194 N_A_199_294#_c_189_n N_A_27_368#_M1008_g 0.00451766f $X=5.995 $Y=1.94
+ $X2=0 $Y2=0
cc_195 N_A_199_294#_c_230_p N_A_27_368#_M1008_g 0.00608819f $X=6.715 $Y=2.135
+ $X2=0 $Y2=0
cc_196 N_A_199_294#_c_200_n N_A_27_368#_M1008_g 0.00621526f $X=6.08 $Y=2.08
+ $X2=0 $Y2=0
cc_197 N_A_199_294#_c_188_n N_A_27_368#_M1013_g 0.0108741f $X=5.995 $Y=1.3 $X2=0
+ $Y2=0
cc_198 N_A_199_294#_c_189_n N_A_27_368#_M1013_g 0.00444636f $X=5.995 $Y=1.94
+ $X2=0 $Y2=0
cc_199 N_A_199_294#_c_188_n N_A_27_368#_M1023_g 2.63345e-19 $X=5.995 $Y=1.3
+ $X2=0 $Y2=0
cc_200 N_A_199_294#_c_189_n N_A_27_368#_M1023_g 5.77979e-19 $X=5.995 $Y=1.94
+ $X2=0 $Y2=0
cc_201 N_A_199_294#_c_189_n N_A_27_368#_M1012_g 8.11005e-19 $X=5.995 $Y=1.94
+ $X2=0 $Y2=0
cc_202 N_A_199_294#_c_230_p N_A_27_368#_M1012_g 0.0120335f $X=6.715 $Y=2.135
+ $X2=0 $Y2=0
cc_203 N_A_199_294#_M1010_d N_A_27_368#_c_502_n 0.00460877f $X=3.215 $Y=1.96
+ $X2=0 $Y2=0
cc_204 N_A_199_294#_M1020_d N_A_27_368#_c_502_n 0.0250614f $X=4.2 $Y=1.96 $X2=0
+ $Y2=0
cc_205 N_A_199_294#_M1006_d N_A_27_368#_c_502_n 0.00460877f $X=5.68 $Y=1.96
+ $X2=0 $Y2=0
cc_206 N_A_199_294#_M1012_s N_A_27_368#_c_502_n 0.00460877f $X=6.58 $Y=1.96
+ $X2=0 $Y2=0
cc_207 N_A_199_294#_M1001_g N_A_27_368#_c_502_n 0.016203f $X=1.085 $Y=2.4 $X2=0
+ $Y2=0
cc_208 N_A_199_294#_M1014_g N_A_27_368#_c_502_n 0.0130202f $X=1.535 $Y=2.4 $X2=0
+ $Y2=0
cc_209 N_A_199_294#_M1015_g N_A_27_368#_c_502_n 0.0136231f $X=2.015 $Y=2.4 $X2=0
+ $Y2=0
cc_210 N_A_199_294#_M1017_g N_A_27_368#_c_502_n 0.016684f $X=2.575 $Y=2.4 $X2=0
+ $Y2=0
cc_211 N_A_199_294#_c_197_n N_A_27_368#_c_502_n 0.238898f $X=3.38 $Y=2.085 $X2=0
+ $Y2=0
cc_212 N_A_199_294#_c_247_p N_A_27_368#_c_502_n 0.00868214f $X=2.745 $Y=2.085
+ $X2=0 $Y2=0
cc_213 N_A_199_294#_c_189_n N_A_27_368#_c_484_n 0.00543065f $X=5.995 $Y=1.94
+ $X2=0 $Y2=0
cc_214 N_A_199_294#_c_230_p N_A_27_368#_c_485_n 0.00405709f $X=6.715 $Y=2.135
+ $X2=0 $Y2=0
cc_215 N_A_199_294#_c_188_n N_A_27_368#_c_530_n 0.00867849f $X=5.995 $Y=1.3
+ $X2=0 $Y2=0
cc_216 N_A_199_294#_c_230_p N_A_27_368#_c_486_n 0.00881139f $X=6.715 $Y=2.135
+ $X2=0 $Y2=0
cc_217 N_A_199_294#_M1001_g N_A_27_368#_c_495_n 0.0019982f $X=1.085 $Y=2.4 $X2=0
+ $Y2=0
cc_218 N_A_199_294#_M1001_g N_A_27_368#_c_497_n 5.7858e-19 $X=1.085 $Y=2.4 $X2=0
+ $Y2=0
cc_219 N_A_199_294#_c_188_n N_A_27_368#_c_489_n 0.00681497f $X=5.995 $Y=1.3
+ $X2=0 $Y2=0
cc_220 N_A_199_294#_c_189_n N_A_27_368#_c_489_n 0.0240318f $X=5.995 $Y=1.94
+ $X2=0 $Y2=0
cc_221 N_A_199_294#_c_230_p N_A_27_368#_c_489_n 0.0278147f $X=6.715 $Y=2.135
+ $X2=0 $Y2=0
cc_222 N_A_199_294#_c_188_n N_A_27_368#_c_490_n 0.00265935f $X=5.995 $Y=1.3
+ $X2=0 $Y2=0
cc_223 N_A_199_294#_c_189_n N_A_27_368#_c_490_n 0.00996337f $X=5.995 $Y=1.94
+ $X2=0 $Y2=0
cc_224 N_A_199_294#_c_230_p N_A_27_368#_c_490_n 0.00223679f $X=6.715 $Y=2.135
+ $X2=0 $Y2=0
cc_225 N_A_199_294#_c_208_p N_B_M1006_g 0.0153699f $X=5.65 $Y=2.08 $X2=0 $Y2=0
cc_226 N_A_199_294#_c_200_n N_B_M1006_g 0.00327698f $X=6.08 $Y=2.08 $X2=0 $Y2=0
cc_227 N_A_199_294#_c_188_n N_B_M1002_g 0.0011858f $X=5.995 $Y=1.3 $X2=0 $Y2=0
cc_228 N_A_199_294#_c_189_n N_B_M1002_g 0.0123228f $X=5.995 $Y=1.94 $X2=0 $Y2=0
cc_229 N_A_199_294#_c_230_p N_B_M1018_g 0.00558462f $X=6.715 $Y=2.135 $X2=0
+ $Y2=0
cc_230 N_A_199_294#_c_230_p B 0.00237667f $X=6.715 $Y=2.135 $X2=0 $Y2=0
cc_231 N_A_199_294#_c_196_n N_VPWR_M1017_d 0.00138946f $X=2.66 $Y=1.95 $X2=0
+ $Y2=0
cc_232 N_A_199_294#_c_197_n N_VPWR_M1017_d 0.00947528f $X=3.38 $Y=2.085 $X2=0
+ $Y2=0
cc_233 N_A_199_294#_c_247_p N_VPWR_M1017_d 2.44056e-19 $X=2.745 $Y=2.085 $X2=0
+ $Y2=0
cc_234 N_A_199_294#_c_208_p N_VPWR_M1003_s 0.00652354f $X=5.65 $Y=2.08 $X2=0
+ $Y2=0
cc_235 N_A_199_294#_c_208_p N_VPWR_M1024_s 0.00566202f $X=5.65 $Y=2.08 $X2=0
+ $Y2=0
cc_236 N_A_199_294#_c_230_p N_VPWR_M1008_d 0.00362734f $X=6.715 $Y=2.135 $X2=0
+ $Y2=0
cc_237 N_A_199_294#_M1001_g N_VPWR_c_679_n 0.0105007f $X=1.085 $Y=2.4 $X2=0
+ $Y2=0
cc_238 N_A_199_294#_M1014_g N_VPWR_c_679_n 0.00105281f $X=1.535 $Y=2.4 $X2=0
+ $Y2=0
cc_239 N_A_199_294#_M1001_g N_VPWR_c_680_n 0.00105306f $X=1.085 $Y=2.4 $X2=0
+ $Y2=0
cc_240 N_A_199_294#_M1014_g N_VPWR_c_680_n 0.00951896f $X=1.535 $Y=2.4 $X2=0
+ $Y2=0
cc_241 N_A_199_294#_M1015_g N_VPWR_c_680_n 0.0101857f $X=2.015 $Y=2.4 $X2=0
+ $Y2=0
cc_242 N_A_199_294#_M1017_g N_VPWR_c_680_n 0.00165045f $X=2.575 $Y=2.4 $X2=0
+ $Y2=0
cc_243 N_A_199_294#_M1015_g N_VPWR_c_681_n 0.00460063f $X=2.015 $Y=2.4 $X2=0
+ $Y2=0
cc_244 N_A_199_294#_M1017_g N_VPWR_c_681_n 0.00460063f $X=2.575 $Y=2.4 $X2=0
+ $Y2=0
cc_245 N_A_199_294#_M1015_g N_VPWR_c_682_n 0.00165118f $X=2.015 $Y=2.4 $X2=0
+ $Y2=0
cc_246 N_A_199_294#_M1017_g N_VPWR_c_682_n 0.0101405f $X=2.575 $Y=2.4 $X2=0
+ $Y2=0
cc_247 N_A_199_294#_M1001_g N_VPWR_c_692_n 0.00460063f $X=1.085 $Y=2.4 $X2=0
+ $Y2=0
cc_248 N_A_199_294#_M1014_g N_VPWR_c_692_n 0.00460063f $X=1.535 $Y=2.4 $X2=0
+ $Y2=0
cc_249 N_A_199_294#_M1001_g N_VPWR_c_678_n 0.00443247f $X=1.085 $Y=2.4 $X2=0
+ $Y2=0
cc_250 N_A_199_294#_M1014_g N_VPWR_c_678_n 0.00443247f $X=1.535 $Y=2.4 $X2=0
+ $Y2=0
cc_251 N_A_199_294#_M1015_g N_VPWR_c_678_n 0.00444262f $X=2.015 $Y=2.4 $X2=0
+ $Y2=0
cc_252 N_A_199_294#_M1017_g N_VPWR_c_678_n 0.00444262f $X=2.575 $Y=2.4 $X2=0
+ $Y2=0
cc_253 N_A_199_294#_M1014_g N_X_c_777_n 0.0176399f $X=1.535 $Y=2.4 $X2=0 $Y2=0
cc_254 N_A_199_294#_M1015_g N_X_c_777_n 0.0170888f $X=2.015 $Y=2.4 $X2=0 $Y2=0
cc_255 N_A_199_294#_M1017_g N_X_c_777_n 0.00361685f $X=2.575 $Y=2.4 $X2=0 $Y2=0
cc_256 N_A_199_294#_c_187_n N_X_c_777_n 0.0725988f $X=2.575 $Y=1.485 $X2=0 $Y2=0
cc_257 N_A_199_294#_c_196_n N_X_c_777_n 0.010181f $X=2.66 $Y=1.95 $X2=0 $Y2=0
cc_258 N_A_199_294#_c_247_p N_X_c_777_n 0.0235114f $X=2.745 $Y=2.085 $X2=0 $Y2=0
cc_259 N_A_199_294#_c_190_n N_X_c_777_n 8.03946e-19 $X=1.445 $Y=1.485 $X2=0
+ $Y2=0
cc_260 N_A_199_294#_c_191_n N_X_c_777_n 0.00783942f $X=2.59 $Y=1.485 $X2=0 $Y2=0
cc_261 N_A_199_294#_M1009_g N_X_c_772_n 0.0123455f $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A_199_294#_M1022_g N_X_c_772_n 0.0133553f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_263 N_A_199_294#_M1025_g N_X_c_772_n 0.00283169f $X=2.59 $Y=0.74 $X2=0 $Y2=0
cc_264 N_A_199_294#_c_187_n N_X_c_772_n 0.0811859f $X=2.575 $Y=1.485 $X2=0 $Y2=0
cc_265 N_A_199_294#_c_191_n N_X_c_772_n 0.0101468f $X=2.59 $Y=1.485 $X2=0 $Y2=0
cc_266 N_A_199_294#_M1009_g N_X_c_773_n 8.39752e-19 $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_267 N_A_199_294#_M1022_g N_X_c_773_n 0.010036f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_268 N_A_199_294#_M1025_g N_X_c_773_n 0.00768257f $X=2.59 $Y=0.74 $X2=0 $Y2=0
cc_269 N_A_199_294#_M1005_g X 0.00437707f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_270 N_A_199_294#_M1009_g X 0.00156393f $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_271 N_A_199_294#_c_190_n X 0.00107372f $X=1.445 $Y=1.485 $X2=0 $Y2=0
cc_272 N_A_199_294#_M1001_g X 0.0081899f $X=1.085 $Y=2.4 $X2=0 $Y2=0
cc_273 N_A_199_294#_M1005_g X 0.004196f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_274 N_A_199_294#_M1009_g X 0.00389182f $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_275 N_A_199_294#_c_186_n X 0.00471673f $X=0.995 $Y=1.47 $X2=0 $Y2=0
cc_276 N_A_199_294#_c_187_n X 0.0262135f $X=2.575 $Y=1.485 $X2=0 $Y2=0
cc_277 N_A_199_294#_c_190_n X 0.00662179f $X=1.445 $Y=1.485 $X2=0 $Y2=0
cc_278 N_A_199_294#_c_191_n X 0.00527145f $X=2.59 $Y=1.485 $X2=0 $Y2=0
cc_279 N_A_199_294#_M1005_g N_X_c_776_n 0.010518f $X=1.09 $Y=0.74 $X2=0 $Y2=0
cc_280 N_A_199_294#_M1009_g N_X_c_776_n 0.00998276f $X=1.52 $Y=0.74 $X2=0 $Y2=0
cc_281 N_A_199_294#_M1022_g N_X_c_776_n 8.33931e-19 $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_282 N_A_199_294#_M1001_g N_X_c_785_n 0.0115816f $X=1.085 $Y=2.4 $X2=0 $Y2=0
cc_283 N_A_199_294#_M1005_g N_VGND_c_834_n 0.00974391f $X=1.09 $Y=0.74 $X2=0
+ $Y2=0
cc_284 N_A_199_294#_M1005_g N_VGND_c_835_n 0.00371957f $X=1.09 $Y=0.74 $X2=0
+ $Y2=0
cc_285 N_A_199_294#_M1009_g N_VGND_c_835_n 0.00434272f $X=1.52 $Y=0.74 $X2=0
+ $Y2=0
cc_286 N_A_199_294#_M1009_g N_VGND_c_836_n 0.0077868f $X=1.52 $Y=0.74 $X2=0
+ $Y2=0
cc_287 N_A_199_294#_M1022_g N_VGND_c_836_n 0.00772705f $X=2.16 $Y=0.74 $X2=0
+ $Y2=0
cc_288 N_A_199_294#_M1025_g N_VGND_c_837_n 0.00815524f $X=2.59 $Y=0.74 $X2=0
+ $Y2=0
cc_289 N_A_199_294#_c_187_n N_VGND_c_837_n 0.00294321f $X=2.575 $Y=1.485 $X2=0
+ $Y2=0
cc_290 N_A_199_294#_M1022_g N_VGND_c_839_n 0.00434272f $X=2.16 $Y=0.74 $X2=0
+ $Y2=0
cc_291 N_A_199_294#_M1025_g N_VGND_c_839_n 0.00434272f $X=2.59 $Y=0.74 $X2=0
+ $Y2=0
cc_292 N_A_199_294#_M1005_g N_VGND_c_844_n 0.00624491f $X=1.09 $Y=0.74 $X2=0
+ $Y2=0
cc_293 N_A_199_294#_M1009_g N_VGND_c_844_n 0.00822469f $X=1.52 $Y=0.74 $X2=0
+ $Y2=0
cc_294 N_A_199_294#_M1022_g N_VGND_c_844_n 0.00822693f $X=2.16 $Y=0.74 $X2=0
+ $Y2=0
cc_295 N_A_199_294#_M1025_g N_VGND_c_844_n 0.00821384f $X=2.59 $Y=0.74 $X2=0
+ $Y2=0
cc_296 N_A_199_294#_c_188_n N_A_664_125#_c_918_n 0.00159069f $X=5.995 $Y=1.3
+ $X2=0 $Y2=0
cc_297 N_A_199_294#_c_208_p N_A_664_125#_c_918_n 0.0158984f $X=5.65 $Y=2.08
+ $X2=0 $Y2=0
cc_298 N_A_199_294#_c_199_n N_A_664_125#_c_919_n 0.00175759f $X=3.515 $Y=2.085
+ $X2=0 $Y2=0
cc_299 N_A_199_294#_c_208_p N_A_664_125#_c_919_n 0.00323763f $X=5.65 $Y=2.08
+ $X2=0 $Y2=0
cc_300 N_A_199_294#_M1013_s N_A_1136_125#_c_1000_n 0.00176461f $X=6.11 $Y=0.625
+ $X2=0 $Y2=0
cc_301 N_A_199_294#_c_188_n N_A_1136_125#_c_1000_n 0.0198997f $X=5.995 $Y=1.3
+ $X2=0 $Y2=0
cc_302 N_D_c_338_n N_C_M1010_g 0.0519766f $X=3.665 $Y=1.725 $X2=0 $Y2=0
cc_303 N_D_c_338_n N_C_M1000_g 0.00883137f $X=3.665 $Y=1.725 $X2=0 $Y2=0
cc_304 N_D_c_339_n N_C_M1000_g 0.0213925f $X=4.155 $Y=1.345 $X2=0 $Y2=0
cc_305 N_D_c_339_n N_C_c_399_n 0.00852785f $X=4.155 $Y=1.345 $X2=0 $Y2=0
cc_306 N_D_c_340_n N_C_c_399_n 0.00852641f $X=4.745 $Y=1.345 $X2=0 $Y2=0
cc_307 D N_C_c_408_n 0.00488763f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_308 N_D_c_342_n N_C_c_408_n 0.00296558f $X=4.585 $Y=1.635 $X2=0 $Y2=0
cc_309 N_D_c_340_n N_C_M1016_g 0.0223678f $X=4.745 $Y=1.345 $X2=0 $Y2=0
cc_310 D N_C_c_402_n 0.00914665f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_311 N_D_c_342_n N_C_c_402_n 0.0145538f $X=4.585 $Y=1.635 $X2=0 $Y2=0
cc_312 N_D_c_340_n N_C_c_403_n 0.00502045f $X=4.745 $Y=1.345 $X2=0 $Y2=0
cc_313 D N_C_c_403_n 0.00179587f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_314 N_D_c_338_n N_C_c_404_n 0.00186082f $X=3.665 $Y=1.725 $X2=0 $Y2=0
cc_315 N_D_c_338_n N_C_c_405_n 0.00250476f $X=3.665 $Y=1.725 $X2=0 $Y2=0
cc_316 N_D_M1003_g N_A_27_368#_c_502_n 0.0135093f $X=3.575 $Y=2.46 $X2=0 $Y2=0
cc_317 N_D_M1020_g N_A_27_368#_c_502_n 0.0154419f $X=4.11 $Y=2.46 $X2=0 $Y2=0
cc_318 D N_B_c_614_n 0.00182507f $X=4.955 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_319 N_D_M1003_g N_VPWR_c_683_n 0.00486592f $X=3.575 $Y=2.46 $X2=0 $Y2=0
cc_320 N_D_M1020_g N_VPWR_c_683_n 0.0183423f $X=4.11 $Y=2.46 $X2=0 $Y2=0
cc_321 N_D_M1003_g N_VPWR_c_686_n 0.00553757f $X=3.575 $Y=2.46 $X2=0 $Y2=0
cc_322 N_D_M1020_g N_VPWR_c_688_n 0.00460063f $X=4.11 $Y=2.46 $X2=0 $Y2=0
cc_323 N_D_M1003_g N_VPWR_c_678_n 0.00535012f $X=3.575 $Y=2.46 $X2=0 $Y2=0
cc_324 N_D_M1020_g N_VPWR_c_678_n 0.0044838f $X=4.11 $Y=2.46 $X2=0 $Y2=0
cc_325 N_D_c_339_n N_VGND_c_838_n 0.00344336f $X=4.155 $Y=1.345 $X2=0 $Y2=0
cc_326 N_D_c_340_n N_VGND_c_838_n 0.00334294f $X=4.745 $Y=1.345 $X2=0 $Y2=0
cc_327 N_D_c_339_n N_VGND_c_844_n 9.49986e-19 $X=4.155 $Y=1.345 $X2=0 $Y2=0
cc_328 N_D_c_340_n N_VGND_c_844_n 9.49986e-19 $X=4.745 $Y=1.345 $X2=0 $Y2=0
cc_329 N_D_c_339_n N_A_664_125#_c_917_n 8.29779e-19 $X=4.155 $Y=1.345 $X2=0
+ $Y2=0
cc_330 N_D_c_337_n N_A_664_125#_c_918_n 0.00474719f $X=4.02 $Y=1.725 $X2=0 $Y2=0
cc_331 N_D_c_338_n N_A_664_125#_c_918_n 5.26644e-19 $X=3.665 $Y=1.725 $X2=0
+ $Y2=0
cc_332 N_D_c_339_n N_A_664_125#_c_918_n 0.0114991f $X=4.155 $Y=1.345 $X2=0 $Y2=0
cc_333 N_D_c_340_n N_A_664_125#_c_918_n 0.0112328f $X=4.745 $Y=1.345 $X2=0 $Y2=0
cc_334 D N_A_664_125#_c_918_n 0.0895722f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_335 N_D_c_342_n N_A_664_125#_c_918_n 0.00722393f $X=4.585 $Y=1.635 $X2=0
+ $Y2=0
cc_336 N_D_c_338_n N_A_664_125#_c_919_n 0.00335791f $X=3.665 $Y=1.725 $X2=0
+ $Y2=0
cc_337 N_D_c_339_n N_A_751_125#_c_977_n 0.00759913f $X=4.155 $Y=1.345 $X2=0
+ $Y2=0
cc_338 N_D_c_340_n N_A_751_125#_c_977_n 0.00813572f $X=4.745 $Y=1.345 $X2=0
+ $Y2=0
cc_339 N_D_c_339_n N_A_751_125#_c_979_n 0.00433778f $X=4.155 $Y=1.345 $X2=0
+ $Y2=0
cc_340 N_D_c_340_n N_A_751_125#_c_979_n 7.19935e-19 $X=4.745 $Y=1.345 $X2=0
+ $Y2=0
cc_341 N_D_c_339_n N_A_751_125#_c_976_n 8.5254e-19 $X=4.155 $Y=1.345 $X2=0 $Y2=0
cc_342 N_D_c_340_n N_A_751_125#_c_976_n 0.00545393f $X=4.745 $Y=1.345 $X2=0
+ $Y2=0
cc_343 N_C_M1010_g N_A_27_368#_c_502_n 0.0135265f $X=3.125 $Y=2.46 $X2=0 $Y2=0
cc_344 N_C_M1024_g N_A_27_368#_c_502_n 0.015041f $X=5.12 $Y=2.46 $X2=0 $Y2=0
cc_345 N_C_c_403_n N_B_c_614_n 0.00513299f $X=5.155 $Y=1.49 $X2=-0.19 $Y2=-0.245
cc_346 N_C_c_402_n N_B_M1006_g 0.057411f $X=5.12 $Y=1.735 $X2=0 $Y2=0
cc_347 N_C_M1016_g N_B_M1002_g 0.0138613f $X=5.175 $Y=0.945 $X2=0 $Y2=0
cc_348 N_C_c_399_n N_B_c_618_n 0.0138613f $X=5.1 $Y=0.18 $X2=0 $Y2=0
cc_349 N_C_M1010_g N_VPWR_c_682_n 0.00496468f $X=3.125 $Y=2.46 $X2=0 $Y2=0
cc_350 N_C_M1024_g N_VPWR_c_684_n 0.0184468f $X=5.12 $Y=2.46 $X2=0 $Y2=0
cc_351 N_C_M1010_g N_VPWR_c_686_n 0.00553757f $X=3.125 $Y=2.46 $X2=0 $Y2=0
cc_352 N_C_M1024_g N_VPWR_c_688_n 0.00460063f $X=5.12 $Y=2.46 $X2=0 $Y2=0
cc_353 N_C_M1010_g N_VPWR_c_678_n 0.00535191f $X=3.125 $Y=2.46 $X2=0 $Y2=0
cc_354 N_C_M1024_g N_VPWR_c_678_n 0.0044838f $X=5.12 $Y=2.46 $X2=0 $Y2=0
cc_355 N_C_c_397_n N_VGND_c_837_n 0.0213937f $X=3.245 $Y=0.18 $X2=0 $Y2=0
cc_356 N_C_c_404_n N_VGND_c_837_n 9.42658e-19 $X=3.08 $Y=1.515 $X2=0 $Y2=0
cc_357 N_C_c_405_n N_VGND_c_837_n 0.008741f $X=3.08 $Y=1.515 $X2=0 $Y2=0
cc_358 N_C_M1000_g N_VGND_c_838_n 0.00634879f $X=3.68 $Y=0.945 $X2=0 $Y2=0
cc_359 N_C_c_399_n N_VGND_c_838_n 0.025075f $X=5.1 $Y=0.18 $X2=0 $Y2=0
cc_360 N_C_M1016_g N_VGND_c_838_n 0.00659036f $X=5.175 $Y=0.945 $X2=0 $Y2=0
cc_361 N_C_c_397_n N_VGND_c_842_n 0.0372748f $X=3.245 $Y=0.18 $X2=0 $Y2=0
cc_362 N_C_c_399_n N_VGND_c_843_n 0.0196635f $X=5.1 $Y=0.18 $X2=0 $Y2=0
cc_363 N_C_c_396_n N_VGND_c_844_n 0.0116023f $X=3.605 $Y=0.18 $X2=0 $Y2=0
cc_364 N_C_c_397_n N_VGND_c_844_n 0.011445f $X=3.245 $Y=0.18 $X2=0 $Y2=0
cc_365 N_C_c_399_n N_VGND_c_844_n 0.0386483f $X=5.1 $Y=0.18 $X2=0 $Y2=0
cc_366 N_C_c_401_n N_VGND_c_844_n 0.00846253f $X=3.68 $Y=0.18 $X2=0 $Y2=0
cc_367 N_C_c_396_n N_A_664_125#_c_917_n 0.00353352f $X=3.605 $Y=0.18 $X2=0 $Y2=0
cc_368 N_C_M1000_g N_A_664_125#_c_917_n 0.00930239f $X=3.68 $Y=0.945 $X2=0 $Y2=0
cc_369 N_C_c_406_n N_A_664_125#_c_917_n 0.00523221f $X=3.08 $Y=1.35 $X2=0 $Y2=0
cc_370 N_C_M1000_g N_A_664_125#_c_918_n 0.0116916f $X=3.68 $Y=0.945 $X2=0 $Y2=0
cc_371 N_C_M1016_g N_A_664_125#_c_918_n 0.0136807f $X=5.175 $Y=0.945 $X2=0 $Y2=0
cc_372 N_C_c_403_n N_A_664_125#_c_918_n 0.00122885f $X=5.155 $Y=1.49 $X2=0 $Y2=0
cc_373 N_C_M1000_g N_A_664_125#_c_919_n 0.00248638f $X=3.68 $Y=0.945 $X2=0 $Y2=0
cc_374 N_C_c_406_n N_A_664_125#_c_919_n 0.00485899f $X=3.08 $Y=1.35 $X2=0 $Y2=0
cc_375 N_C_M1016_g N_A_664_125#_c_920_n 0.0044159f $X=5.175 $Y=0.945 $X2=0 $Y2=0
cc_376 N_C_M1016_g N_A_664_125#_c_922_n 0.00537518f $X=5.175 $Y=0.945 $X2=0
+ $Y2=0
cc_377 N_C_c_399_n N_A_751_125#_c_977_n 0.00200023f $X=5.1 $Y=0.18 $X2=0 $Y2=0
cc_378 N_C_c_399_n N_A_751_125#_c_979_n 0.00413604f $X=5.1 $Y=0.18 $X2=0 $Y2=0
cc_379 N_C_c_399_n N_A_751_125#_c_976_n 0.00367611f $X=5.1 $Y=0.18 $X2=0 $Y2=0
cc_380 N_C_M1016_g N_A_751_125#_c_976_n 0.00469613f $X=5.175 $Y=0.945 $X2=0
+ $Y2=0
cc_381 N_A_27_368#_c_490_n N_B_c_614_n 0.0162934f $X=6.465 $Y=1.635 $X2=-0.19
+ $Y2=-0.245
cc_382 N_A_27_368#_c_502_n N_B_M1006_g 0.0128792f $X=7.35 $Y=2.475 $X2=0 $Y2=0
cc_383 N_A_27_368#_c_490_n N_B_M1006_g 0.0520569f $X=6.465 $Y=1.635 $X2=0 $Y2=0
cc_384 N_A_27_368#_M1013_g N_B_M1002_g 0.0162934f $X=6.035 $Y=0.945 $X2=0 $Y2=0
cc_385 N_A_27_368#_M1013_g N_B_c_617_n 0.00737859f $X=6.035 $Y=0.945 $X2=0 $Y2=0
cc_386 N_A_27_368#_M1023_g N_B_c_617_n 0.00737859f $X=6.465 $Y=0.945 $X2=0 $Y2=0
cc_387 N_A_27_368#_M1012_g N_B_M1018_g 0.0303159f $X=6.49 $Y=2.46 $X2=0 $Y2=0
cc_388 N_A_27_368#_c_502_n N_B_M1018_g 0.0166205f $X=7.35 $Y=2.475 $X2=0 $Y2=0
cc_389 N_A_27_368#_c_486_n N_B_M1018_g 0.0148916f $X=7.435 $Y=2.39 $X2=0 $Y2=0
cc_390 N_A_27_368#_M1023_g N_B_M1019_g 0.0182961f $X=6.465 $Y=0.945 $X2=0 $Y2=0
cc_391 N_A_27_368#_c_484_n N_B_M1019_g 7.10656e-19 $X=6.59 $Y=1.47 $X2=0 $Y2=0
cc_392 N_A_27_368#_c_485_n N_B_M1019_g 0.0170156f $X=7.35 $Y=1.215 $X2=0 $Y2=0
cc_393 N_A_27_368#_c_486_n N_B_M1019_g 0.0123314f $X=7.435 $Y=2.39 $X2=0 $Y2=0
cc_394 N_A_27_368#_c_502_n B 0.00718092f $X=7.35 $Y=2.475 $X2=0 $Y2=0
cc_395 N_A_27_368#_c_485_n B 0.0246739f $X=7.35 $Y=1.215 $X2=0 $Y2=0
cc_396 N_A_27_368#_c_486_n B 0.0248009f $X=7.435 $Y=2.39 $X2=0 $Y2=0
cc_397 N_A_27_368#_c_489_n B 0.0281241f $X=6.59 $Y=1.635 $X2=0 $Y2=0
cc_398 N_A_27_368#_c_490_n B 9.04921e-19 $X=6.465 $Y=1.635 $X2=0 $Y2=0
cc_399 N_A_27_368#_c_502_n N_B_c_621_n 0.00287884f $X=7.35 $Y=2.475 $X2=0 $Y2=0
cc_400 N_A_27_368#_c_485_n N_B_c_621_n 0.00496909f $X=7.35 $Y=1.215 $X2=0 $Y2=0
cc_401 N_A_27_368#_c_489_n N_B_c_621_n 0.00117267f $X=6.59 $Y=1.635 $X2=0 $Y2=0
cc_402 N_A_27_368#_c_490_n N_B_c_621_n 0.0303159f $X=6.465 $Y=1.635 $X2=0 $Y2=0
cc_403 N_A_27_368#_c_502_n N_VPWR_M1004_d 0.0142647f $X=7.35 $Y=2.475 $X2=-0.19
+ $Y2=-0.245
cc_404 N_A_27_368#_c_502_n N_VPWR_M1014_d 0.00392025f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_405 N_A_27_368#_c_502_n N_VPWR_M1017_d 0.00546672f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_406 N_A_27_368#_c_502_n N_VPWR_M1003_s 0.00491544f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_407 N_A_27_368#_c_502_n N_VPWR_M1024_s 0.00370949f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_408 N_A_27_368#_c_502_n N_VPWR_M1008_d 0.0032036f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_409 N_A_27_368#_c_502_n N_VPWR_M1018_s 0.0229256f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_410 N_A_27_368#_c_486_n N_VPWR_M1018_s 0.0261094f $X=7.435 $Y=2.39 $X2=0
+ $Y2=0
cc_411 N_A_27_368#_c_502_n N_VPWR_c_679_n 0.0247246f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_412 N_A_27_368#_c_497_n N_VPWR_c_679_n 0.00496211f $X=0.265 $Y=2.475 $X2=0
+ $Y2=0
cc_413 N_A_27_368#_c_502_n N_VPWR_c_680_n 0.0189213f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_414 N_A_27_368#_c_502_n N_VPWR_c_682_n 0.022352f $X=7.35 $Y=2.475 $X2=0 $Y2=0
cc_415 N_A_27_368#_c_502_n N_VPWR_c_683_n 0.0211657f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_416 N_A_27_368#_M1008_g N_VPWR_c_684_n 0.00105324f $X=6.04 $Y=2.46 $X2=0
+ $Y2=0
cc_417 N_A_27_368#_c_502_n N_VPWR_c_684_n 0.0181304f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_418 N_A_27_368#_M1008_g N_VPWR_c_685_n 0.00937886f $X=6.04 $Y=2.46 $X2=0
+ $Y2=0
cc_419 N_A_27_368#_M1012_g N_VPWR_c_685_n 0.00937327f $X=6.49 $Y=2.46 $X2=0
+ $Y2=0
cc_420 N_A_27_368#_c_502_n N_VPWR_c_685_n 0.0165487f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_421 N_A_27_368#_M1008_g N_VPWR_c_690_n 0.00460063f $X=6.04 $Y=2.46 $X2=0
+ $Y2=0
cc_422 N_A_27_368#_M1012_g N_VPWR_c_693_n 0.00460063f $X=6.49 $Y=2.46 $X2=0
+ $Y2=0
cc_423 N_A_27_368#_c_497_n N_VPWR_c_694_n 0.0106591f $X=0.265 $Y=2.475 $X2=0
+ $Y2=0
cc_424 N_A_27_368#_M1012_g N_VPWR_c_697_n 0.0010519f $X=6.49 $Y=2.46 $X2=0 $Y2=0
cc_425 N_A_27_368#_c_502_n N_VPWR_c_697_n 0.0377578f $X=7.35 $Y=2.475 $X2=0
+ $Y2=0
cc_426 N_A_27_368#_M1008_g N_VPWR_c_678_n 0.00443357f $X=6.04 $Y=2.46 $X2=0
+ $Y2=0
cc_427 N_A_27_368#_M1012_g N_VPWR_c_678_n 0.00443357f $X=6.49 $Y=2.46 $X2=0
+ $Y2=0
cc_428 N_A_27_368#_c_502_n N_VPWR_c_678_n 0.159711f $X=7.35 $Y=2.475 $X2=0 $Y2=0
cc_429 N_A_27_368#_c_497_n N_VPWR_c_678_n 0.0122002f $X=0.265 $Y=2.475 $X2=0
+ $Y2=0
cc_430 N_A_27_368#_c_502_n N_X_M1001_s 0.00460662f $X=7.35 $Y=2.475 $X2=0 $Y2=0
cc_431 N_A_27_368#_c_502_n N_X_M1015_s 0.00867701f $X=7.35 $Y=2.475 $X2=0 $Y2=0
cc_432 N_A_27_368#_c_502_n N_X_c_777_n 0.0650205f $X=7.35 $Y=2.475 $X2=0 $Y2=0
cc_433 N_A_27_368#_c_502_n N_X_c_785_n 0.0135664f $X=7.35 $Y=2.475 $X2=0 $Y2=0
cc_434 N_A_27_368#_c_495_n N_X_c_785_n 0.010611f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_435 N_A_27_368#_c_483_n N_VGND_c_834_n 0.0211853f $X=0.245 $Y=0.86 $X2=0
+ $Y2=0
cc_436 N_A_27_368#_c_483_n N_VGND_c_841_n 0.0100349f $X=0.245 $Y=0.86 $X2=0
+ $Y2=0
cc_437 N_A_27_368#_c_483_n N_VGND_c_844_n 0.0109771f $X=0.245 $Y=0.86 $X2=0
+ $Y2=0
cc_438 N_A_27_368#_c_485_n N_A_664_125#_M1019_d 0.00315946f $X=7.35 $Y=1.215
+ $X2=0 $Y2=0
cc_439 N_A_27_368#_M1013_g N_A_664_125#_c_921_n 0.00116683f $X=6.035 $Y=0.945
+ $X2=0 $Y2=0
cc_440 N_A_27_368#_M1023_g N_A_664_125#_c_921_n 0.00116683f $X=6.465 $Y=0.945
+ $X2=0 $Y2=0
cc_441 N_A_27_368#_M1023_g N_A_664_125#_c_923_n 5.83127e-19 $X=6.465 $Y=0.945
+ $X2=0 $Y2=0
cc_442 N_A_27_368#_c_485_n N_A_664_125#_c_923_n 0.023263f $X=7.35 $Y=1.215 $X2=0
+ $Y2=0
cc_443 N_A_27_368#_c_485_n N_A_1136_125#_M1023_d 0.00527828f $X=7.35 $Y=1.215
+ $X2=0 $Y2=0
cc_444 N_A_27_368#_c_530_n N_A_1136_125#_M1023_d 9.89161e-19 $X=6.675 $Y=1.215
+ $X2=0 $Y2=0
cc_445 N_A_27_368#_M1013_g N_A_1136_125#_c_1000_n 0.00839754f $X=6.035 $Y=0.945
+ $X2=0 $Y2=0
cc_446 N_A_27_368#_M1023_g N_A_1136_125#_c_1000_n 0.0128612f $X=6.465 $Y=0.945
+ $X2=0 $Y2=0
cc_447 N_A_27_368#_c_530_n N_A_1136_125#_c_1000_n 0.00258843f $X=6.675 $Y=1.215
+ $X2=0 $Y2=0
cc_448 N_A_27_368#_M1023_g N_A_1136_125#_c_1002_n 0.00532016f $X=6.465 $Y=0.945
+ $X2=0 $Y2=0
cc_449 N_A_27_368#_c_485_n N_A_1136_125#_c_1002_n 0.0193536f $X=7.35 $Y=1.215
+ $X2=0 $Y2=0
cc_450 N_A_27_368#_c_530_n N_A_1136_125#_c_1002_n 0.00360032f $X=6.675 $Y=1.215
+ $X2=0 $Y2=0
cc_451 N_B_M1006_g N_VPWR_c_684_n 0.00944044f $X=5.59 $Y=2.46 $X2=0 $Y2=0
cc_452 N_B_M1006_g N_VPWR_c_685_n 0.00105361f $X=5.59 $Y=2.46 $X2=0 $Y2=0
cc_453 N_B_M1018_g N_VPWR_c_685_n 0.00105319f $X=6.94 $Y=2.46 $X2=0 $Y2=0
cc_454 N_B_M1006_g N_VPWR_c_690_n 0.00460063f $X=5.59 $Y=2.46 $X2=0 $Y2=0
cc_455 N_B_M1018_g N_VPWR_c_693_n 0.00460063f $X=6.94 $Y=2.46 $X2=0 $Y2=0
cc_456 N_B_M1018_g N_VPWR_c_697_n 0.0161887f $X=6.94 $Y=2.46 $X2=0 $Y2=0
cc_457 N_B_M1006_g N_VPWR_c_678_n 0.00443357f $X=5.59 $Y=2.46 $X2=0 $Y2=0
cc_458 N_B_M1018_g N_VPWR_c_678_n 0.00441801f $X=6.94 $Y=2.46 $X2=0 $Y2=0
cc_459 N_B_c_618_n N_VGND_c_843_n 0.0351645f $X=5.68 $Y=0.18 $X2=0 $Y2=0
cc_460 N_B_c_617_n N_VGND_c_844_n 0.0374956f $X=7.04 $Y=0.18 $X2=0 $Y2=0
cc_461 N_B_c_618_n N_VGND_c_844_n 0.00460771f $X=5.68 $Y=0.18 $X2=0 $Y2=0
cc_462 N_B_M1002_g N_A_664_125#_c_918_n 4.46128e-19 $X=5.605 $Y=0.945 $X2=0
+ $Y2=0
cc_463 N_B_M1002_g N_A_664_125#_c_920_n 0.00424861f $X=5.605 $Y=0.945 $X2=0
+ $Y2=0
cc_464 N_B_M1002_g N_A_664_125#_c_921_n 0.0151367f $X=5.605 $Y=0.945 $X2=0 $Y2=0
cc_465 N_B_c_617_n N_A_664_125#_c_921_n 0.0230464f $X=7.04 $Y=0.18 $X2=0 $Y2=0
cc_466 N_B_M1019_g N_A_664_125#_c_921_n 0.0142293f $X=7.115 $Y=0.945 $X2=0 $Y2=0
cc_467 N_B_M1019_g N_A_664_125#_c_923_n 0.013896f $X=7.115 $Y=0.945 $X2=0 $Y2=0
cc_468 N_B_M1002_g N_A_1136_125#_c_1001_n 0.00547385f $X=5.605 $Y=0.945 $X2=0
+ $Y2=0
cc_469 N_B_M1019_g N_A_1136_125#_c_1002_n 0.00345017f $X=7.115 $Y=0.945 $X2=0
+ $Y2=0
cc_470 N_VPWR_M1014_d N_X_c_777_n 0.0020349f $X=1.625 $Y=1.84 $X2=0 $Y2=0
cc_471 N_X_c_772_n N_VGND_M1009_d 0.00624639f $X=2.21 $Y=1.065 $X2=0 $Y2=0
cc_472 X N_VGND_c_834_n 0.00329614f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_473 N_X_c_776_n N_VGND_c_834_n 0.0494597f $X=1.305 $Y=0.515 $X2=0 $Y2=0
cc_474 N_X_c_776_n N_VGND_c_835_n 0.0167819f $X=1.305 $Y=0.515 $X2=0 $Y2=0
cc_475 N_X_c_772_n N_VGND_c_836_n 0.0266856f $X=2.21 $Y=1.065 $X2=0 $Y2=0
cc_476 N_X_c_773_n N_VGND_c_836_n 0.0303828f $X=2.375 $Y=0.515 $X2=0 $Y2=0
cc_477 N_X_c_776_n N_VGND_c_836_n 0.0319008f $X=1.305 $Y=0.515 $X2=0 $Y2=0
cc_478 N_X_c_772_n N_VGND_c_837_n 0.00711243f $X=2.21 $Y=1.065 $X2=0 $Y2=0
cc_479 N_X_c_773_n N_VGND_c_837_n 0.0243921f $X=2.375 $Y=0.515 $X2=0 $Y2=0
cc_480 N_X_c_773_n N_VGND_c_839_n 0.0144922f $X=2.375 $Y=0.515 $X2=0 $Y2=0
cc_481 N_X_c_773_n N_VGND_c_844_n 0.0118826f $X=2.375 $Y=0.515 $X2=0 $Y2=0
cc_482 N_X_c_776_n N_VGND_c_844_n 0.0136487f $X=1.305 $Y=0.515 $X2=0 $Y2=0
cc_483 N_VGND_c_837_n N_A_664_125#_c_917_n 0.0324343f $X=2.875 $Y=0.515 $X2=0
+ $Y2=0
cc_484 N_VGND_c_838_n N_A_664_125#_c_917_n 4.21282e-19 $X=4.45 $Y=0.535 $X2=0
+ $Y2=0
cc_485 N_VGND_c_842_n N_A_664_125#_c_917_n 0.00697755f $X=4.285 $Y=0 $X2=0 $Y2=0
cc_486 N_VGND_c_844_n N_A_664_125#_c_917_n 0.00879953f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_487 N_VGND_M1007_d N_A_664_125#_c_918_n 0.00406725f $X=4.23 $Y=0.625 $X2=0
+ $Y2=0
cc_488 N_VGND_c_843_n N_A_664_125#_c_921_n 0.131618f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_489 N_VGND_c_844_n N_A_664_125#_c_921_n 0.0695304f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_490 N_VGND_c_843_n N_A_664_125#_c_922_n 0.0121867f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_491 N_VGND_c_844_n N_A_664_125#_c_922_n 0.00660921f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_492 N_VGND_M1007_d N_A_751_125#_c_977_n 0.00687044f $X=4.23 $Y=0.625 $X2=0
+ $Y2=0
cc_493 N_VGND_c_838_n N_A_751_125#_c_977_n 0.0260575f $X=4.45 $Y=0.535 $X2=0
+ $Y2=0
cc_494 N_VGND_c_844_n N_A_751_125#_c_977_n 0.0119525f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_495 N_VGND_c_842_n N_A_751_125#_c_979_n 0.00490296f $X=4.285 $Y=0 $X2=0 $Y2=0
cc_496 N_VGND_c_844_n N_A_751_125#_c_979_n 0.00747787f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_497 N_VGND_c_838_n N_A_751_125#_c_976_n 0.00113701f $X=4.45 $Y=0.535 $X2=0
+ $Y2=0
cc_498 N_VGND_c_843_n N_A_751_125#_c_976_n 0.00663395f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_499 N_VGND_c_844_n N_A_751_125#_c_976_n 0.00851925f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_500 N_A_664_125#_c_918_n N_A_751_125#_M1000_s 0.00224844f $X=5.305 $Y=1.215
+ $X2=-0.19 $Y2=-0.245
cc_501 N_A_664_125#_c_918_n N_A_751_125#_M1021_s 0.00176461f $X=5.305 $Y=1.215
+ $X2=0 $Y2=0
cc_502 N_A_664_125#_c_918_n N_A_751_125#_c_979_n 0.0584624f $X=5.305 $Y=1.215
+ $X2=0 $Y2=0
cc_503 N_A_664_125#_c_918_n N_A_751_125#_c_976_n 0.0162105f $X=5.305 $Y=1.215
+ $X2=0 $Y2=0
cc_504 N_A_664_125#_c_920_n N_A_751_125#_c_976_n 0.0134102f $X=5.39 $Y=0.77
+ $X2=0 $Y2=0
cc_505 N_A_664_125#_c_921_n N_A_1136_125#_c_1000_n 0.0500146f $X=7.165 $Y=0.34
+ $X2=0 $Y2=0
cc_506 N_A_664_125#_c_920_n N_A_1136_125#_c_1001_n 0.0135851f $X=5.39 $Y=0.77
+ $X2=0 $Y2=0
cc_507 N_A_664_125#_c_921_n N_A_1136_125#_c_1001_n 0.0185025f $X=7.165 $Y=0.34
+ $X2=0 $Y2=0
cc_508 N_A_664_125#_c_921_n N_A_1136_125#_c_1002_n 0.0245759f $X=7.165 $Y=0.34
+ $X2=0 $Y2=0
cc_509 N_A_664_125#_c_923_n N_A_1136_125#_c_1002_n 0.0224808f $X=7.33 $Y=0.78
+ $X2=0 $Y2=0

* NGSPICE file created from sky130_fd_sc_ms__dfxtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__dfxtp_1 CLK D VGND VNB VPB VPWR Q
M1000 VPWR a_1014_424# a_1210_314# VPB pshort w=840000u l=180000u
+  ad=1.41472e+12p pd=1.248e+07u as=2.352e+11p ps=2.24e+06u
M1001 a_1168_124# a_27_74# a_1014_424# VNB nlowvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=2.362e+11p ps=2.07e+06u
M1002 a_209_368# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.553e+11p pd=2.17e+06u as=1.2645e+12p ps=1.059e+07u
M1003 a_1014_424# a_27_74# a_713_458# VPB pshort w=840000u l=180000u
+  ad=2.667e+11p pd=2.39e+06u as=4.41e+11p ps=2.73e+06u
M1004 a_713_458# a_564_463# VGND VNB nlowvt w=550000u l=150000u
+  ad=2.18125e+11p pd=2.05e+06u as=0p ps=0u
M1005 a_1121_508# a_209_368# a_1014_424# VPB pshort w=420000u l=180000u
+  ad=1.869e+11p pd=1.73e+06u as=0p ps=0u
M1006 a_1014_424# a_209_368# a_713_458# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_457_503# D VGND VNB nlowvt w=420000u l=150000u
+  ad=3.1125e+11p pd=2.43e+06u as=0p ps=0u
M1008 VGND a_1014_424# a_1210_314# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1009 VPWR CLK a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1010 a_209_368# a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1011 VPWR a_713_458# a_671_503# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1012 a_564_463# a_209_368# a_457_503# VPB pshort w=420000u l=180000u
+  ad=1.841e+11p pd=1.95e+06u as=1.841e+11p ps=1.95e+06u
M1013 Q a_1210_314# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1014 VGND a_713_458# a_731_101# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1015 a_671_503# a_27_74# a_564_463# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_731_101# a_209_368# a_564_463# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.575e+11p ps=1.73e+06u
M1017 a_564_463# a_27_74# a_457_503# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_713_458# a_564_463# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 Q a_1210_314# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1020 a_457_503# D VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_1210_314# a_1168_124# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND CLK a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1023 VPWR a_1210_314# a_1121_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends


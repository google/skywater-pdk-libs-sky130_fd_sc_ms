* File: sky130_fd_sc_ms__o31ai_4.spice
* Created: Fri Aug 28 18:03:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o31ai_4.pex.spice"
.subckt sky130_fd_sc_ms__o31ai_4  VNB VPB A1 A2 A3 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A1_M1000_g N_A_27_82#_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75007.9 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1000_d N_A1_M1007_g N_A_27_82#_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75007.4 A=0.111 P=1.78 MULT=1
MM1018 N_VGND_M1018_d N_A1_M1018_g N_A_27_82#_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75006.9 A=0.111 P=1.78 MULT=1
MM1027 N_VGND_M1018_d N_A1_M1027_g N_A_27_82#_M1027_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75006.4 A=0.111 P=1.78 MULT=1
MM1003 N_VGND_M1003_d N_A2_M1003_g N_A_27_82#_M1027_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2183 AS=0.1036 PD=1.33 PS=1.02 NRD=25.128 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75006 A=0.111 P=1.78 MULT=1
MM1004 N_VGND_M1003_d N_A2_M1004_g N_A_27_82#_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2183 AS=0.1295 PD=1.33 PS=1.09 NRD=25.128 NRS=0 M=1 R=4.93333 SA=75002.8
+ SB=75005.3 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_A2_M1010_g N_A_27_82#_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003.3
+ SB=75004.8 A=0.111 P=1.78 MULT=1
MM1015 N_VGND_M1010_d N_A2_M1015_g N_A_27_82#_M1015_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75003.7
+ SB=75004.3 A=0.111 P=1.78 MULT=1
MM1011 N_A_27_82#_M1015_s N_A3_M1011_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.3627 PD=1.02 PS=1.75 NRD=0 NRS=70.56 M=1 R=4.93333 SA=75004.2
+ SB=75003.9 A=0.111 P=1.78 MULT=1
MM1014 N_A_27_82#_M1014_d N_A3_M1014_g N_VGND_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.3627 PD=1.02 PS=1.75 NRD=0 NRS=70.56 M=1 R=4.93333 SA=75005.1
+ SB=75003 A=0.111 P=1.78 MULT=1
MM1019 N_A_27_82#_M1014_d N_A3_M1019_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.201 PD=1.02 PS=1.42 NRD=0 NRS=35.124 M=1 R=4.93333 SA=75005.5
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1026 N_A_27_82#_M1026_d N_A3_M1026_g N_VGND_M1019_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.201 PD=1.02 PS=1.42 NRD=0 NRS=35.124 M=1 R=4.93333 SA=75006.1
+ SB=75001.9 A=0.111 P=1.78 MULT=1
MM1013 N_Y_M1013_d N_B1_M1013_g N_A_27_82#_M1026_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75006.6
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1016 N_Y_M1013_d N_B1_M1016_g N_A_27_82#_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75007
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1021 N_Y_M1021_d N_B1_M1021_g N_A_27_82#_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75007.4
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1024 N_Y_M1021_d N_B1_M1024_g N_A_27_82#_M1024_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75007.9
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g N_A_28_368#_M1001_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003.8 A=0.2016 P=2.6 MULT=1
MM1002 N_VPWR_M1001_d N_A1_M1002_g N_A_28_368#_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90003.3 A=0.2016 P=2.6 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g N_A_28_368#_M1002_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90002.9 A=0.2016 P=2.6 MULT=1
MM1006 N_VPWR_M1005_d N_A1_M1006_g N_A_28_368#_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90001.6
+ SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1008 N_A_490_368#_M1008_d N_A2_M1008_g N_A_28_368#_M1006_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90002 SB=90001.9 A=0.2016 P=2.6 MULT=1
MM1009 N_A_490_368#_M1008_d N_A2_M1009_g N_A_28_368#_M1009_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1792 AS=0.3024 PD=1.44 PS=1.66 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90002.5 SB=90001.4 A=0.2016 P=2.6 MULT=1
MM1020 N_A_490_368#_M1020_d N_A2_M1020_g N_A_28_368#_M1009_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3024 PD=1.39 PS=1.66 NRD=0 NRS=37.8043 M=1 R=6.22222
+ SA=90003.3 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1023 N_A_490_368#_M1020_d N_A2_M1023_g N_A_28_368#_M1023_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90003.7 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1017 N_A_490_368#_M1017_d N_A3_M1017_g N_Y_M1017_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003.2 A=0.2016 P=2.6 MULT=1
MM1022 N_A_490_368#_M1017_d N_A3_M1022_g N_Y_M1022_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90002.8 A=0.2016 P=2.6 MULT=1
MM1025 N_A_490_368#_M1025_d N_A3_M1025_g N_Y_M1022_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90002.3 A=0.2016 P=2.6 MULT=1
MM1028 N_A_490_368#_M1025_d N_A3_M1028_g N_Y_M1028_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.5
+ SB=90001.9 A=0.2016 P=2.6 MULT=1
MM1012 N_Y_M1028_s N_B1_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.5684 PD=1.44 PS=2.135 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90001.4 A=0.2016 P=2.6 MULT=1
MM1029 N_Y_M1029_d N_B1_M1029_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.5684 PD=2.8 PS=2.135 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX30_noxref VNB VPB NWDIODE A=16.7772 P=21.76
*
.include "sky130_fd_sc_ms__o31ai_4.pxi.spice"
*
.ends
*
*

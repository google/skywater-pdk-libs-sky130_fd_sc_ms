* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfbbp_1 CLK D RESET_B SCD SCE SET_B VGND VNB VPB VPWR Q
+ Q_N
M1000 VGND a_1250_231# a_1192_96# VNB nlowvt w=420000u l=150000u
+  ad=2.22013e+12p pd=1.787e+07u as=1.61875e+11p ps=1.78e+06u
M1001 VGND a_2037_442# a_2061_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.638e+11p ps=1.62e+06u
M1002 a_877_98# a_622_98# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.516e+11p pd=2.16e+06u as=0p ps=0u
M1003 a_1881_420# a_877_98# a_1880_119# VNB nlowvt w=550000u l=150000u
+  ad=2.3445e+11p pd=2.34e+06u as=1.155e+11p ps=1.52e+06u
M1004 a_2271_74# SET_B VGND VNB nlowvt w=740000u l=150000u
+  ad=4.218e+11p pd=4.1e+06u as=0p ps=0u
M1005 Q a_2881_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1006 a_119_119# SCD VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1007 VGND RESET_B a_1625_93# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1008 VPWR a_1625_93# a_1583_379# VPB pshort w=840000u l=180000u
+  ad=2.88865e+12p pd=2.393e+07u as=2.016e+11p ps=2.16e+06u
M1009 VPWR a_1625_93# a_2387_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.1e+11p ps=2.42e+06u
M1010 VPWR SCD a_27_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=3.584e+11p ps=3.68e+06u
M1011 a_299_119# D a_197_119# VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.709e+11p ps=2.97e+06u
M1012 a_1881_420# a_622_98# a_1769_379# VPB pshort w=840000u l=180000u
+  ad=2.709e+11p pd=2.4e+06u as=3.438e+11p ps=2.85e+06u
M1013 Q_N a_2037_442# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=0p ps=0u
M1014 VPWR CLK a_622_98# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1015 a_1250_231# SET_B VPWR VPB pshort w=840000u l=180000u
+  ad=3.024e+11p pd=2.4e+06u as=0p ps=0u
M1016 VGND a_341_93# a_299_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1880_119# a_1250_231# VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_2037_442# a_2881_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1019 a_877_98# a_622_98# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1020 VPWR a_1250_231# a_1224_419# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1021 a_1250_231# a_1092_96# a_1418_125# VNB nlowvt w=550000u l=150000u
+  ad=1.54e+11p pd=1.66e+06u as=7.81e+11p ps=5.37e+06u
M1022 a_1418_125# a_1625_93# a_1250_231# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q a_2881_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1024 VPWR a_2037_442# a_1989_504# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1025 a_1418_125# SET_B VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_2061_74# a_622_98# a_1881_420# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_2037_442# a_2881_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1028 a_221_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1029 a_1092_96# a_877_98# a_197_119# VPB pshort w=640000u l=180000u
+  ad=2.167e+11p pd=2.05e+06u as=3.52e+11p ps=3.66e+06u
M1030 a_1583_379# a_1092_96# a_1250_231# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1769_379# a_1250_231# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_341_93# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.792e+11p pd=1.84e+06u as=0p ps=0u
M1033 a_197_119# SCE a_119_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1192_96# a_877_98# a_1092_96# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.47e+11p ps=1.54e+06u
M1035 a_2037_442# a_1881_420# a_2271_74# VNB nlowvt w=740000u l=150000u
+  ad=2.886e+11p pd=2.26e+06u as=0p ps=0u
M1036 Q_N a_2037_442# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1037 a_1224_419# a_622_98# a_1092_96# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1092_96# a_622_98# a_197_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_197_119# D a_221_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1989_504# a_877_98# a_1881_420# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_2387_392# a_1881_420# a_2037_442# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=3.7e+11p ps=2.74e+06u
M1042 a_27_464# a_341_93# a_197_119# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_341_93# SCE VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1044 VGND CLK a_622_98# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1045 a_2271_74# a_1625_93# a_2037_442# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 a_2037_442# SET_B VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VPWR RESET_B a_1625_93# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
.ends

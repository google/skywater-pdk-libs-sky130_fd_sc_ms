* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__clkbuf_16 A VGND VNB VPB VPWR X
X0 a_114_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X2 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X4 a_114_74# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X6 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X9 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X10 a_114_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X11 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X12 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X13 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X14 VPWR A a_114_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X16 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X17 VPWR A a_114_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X18 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X19 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X20 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X21 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X22 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X23 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X24 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X25 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X26 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X27 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X28 VPWR a_114_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X29 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X30 X a_114_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X31 a_114_74# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X32 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X33 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X34 VGND A a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X35 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X36 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X37 VGND A a_114_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X38 VGND a_114_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X39 X a_114_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
.ends

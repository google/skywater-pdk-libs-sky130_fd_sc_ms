* File: sky130_fd_sc_ms__dfrtn_1.pex.spice
* Created: Wed Sep  2 12:02:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DFRTN_1%D 2 3 5 9 13 15 20 21 22 27 28
c34 5 0 4.19395e-20 $X=0.5 $Y=2.75
r35 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.125 $X2=0.27 $Y2=1.125
r36 21 22 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.237 $Y=1.665
+ $X2=0.237 $Y2=2.035
r37 20 21 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.237 $Y=1.295
+ $X2=0.237 $Y2=1.665
r38 20 28 7.39303 $w=2.63e-07 $l=1.7e-07 $layer=LI1_cond $X=0.237 $Y=1.295
+ $X2=0.237 $Y2=1.125
r39 14 27 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.465
+ $X2=0.27 $Y2=1.125
r40 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.465
+ $X2=0.27 $Y2=1.63
r41 13 27 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=1.11
+ $X2=0.27 $Y2=1.125
r42 12 13 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.352 $Y=0.96
+ $X2=0.352 $Y2=1.11
r43 9 12 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=0.525 $Y=0.58
+ $X2=0.525 $Y2=0.96
r44 3 16 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=0.5 $Y=1.995 $X2=0.36
+ $Y2=1.995
r45 3 5 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=0.5 $Y=2.07 $X2=0.5
+ $Y2=2.75
r46 2 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.36 $Y=1.92 $X2=0.36
+ $Y2=1.995
r47 2 15 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.36 $Y=1.92 $X2=0.36
+ $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTN_1%CLK_N 1 3 4 6 7 8 9
c47 9 0 1.78864e-19 $X=1.68 $Y=1.295
c48 1 0 1.33645e-19 $X=1.915 $Y=1.66
r49 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.41 $X2=1.61 $Y2=1.41
r50 9 13 4.58497 $w=3.06e-07 $l=1.15e-07 $layer=LI1_cond $X=1.61 $Y=1.295
+ $X2=1.61 $Y2=1.41
r51 7 12 26.5718 $w=4.5e-07 $l=2.15e-07 $layer=POLY_cond $X=1.825 $Y=1.435
+ $X2=1.61 $Y2=1.435
r52 7 8 7.41388 $w=4.5e-07 $l=9e-08 $layer=POLY_cond $X=1.825 $Y=1.435 $X2=1.915
+ $Y2=1.435
r53 4 8 42.5959 $w=1.65e-07 $l=2.32379e-07 $layer=POLY_cond $X=1.93 $Y=1.21
+ $X2=1.915 $Y2=1.435
r54 4 6 151.027 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.93 $Y=1.21 $X2=1.93
+ $Y2=0.74
r55 1 8 42.5959 $w=1.65e-07 $l=2.25e-07 $layer=POLY_cond $X=1.915 $Y=1.66
+ $X2=1.915 $Y2=1.435
r56 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.915 $Y=1.66
+ $X2=1.915 $Y2=2.235
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTN_1%A_510_74# 1 2 9 13 15 19 22 23 25 27 28 32
+ 35 36 39 40 42 45 46 47 49 50 51 53 55 56 58 59 62 63 65 66 67 72
c188 72 0 1.01786e-19 $X=7.42 $Y=1.29
c189 66 0 1.94919e-19 $X=3.62 $Y=0.36
c190 62 0 1.33645e-19 $X=2.73 $Y=1.915
c191 58 0 2.79847e-19 $X=7.255 $Y=1.29
c192 56 0 2.84298e-19 $X=7.08 $Y=1.29
c193 55 0 2.21313e-20 $X=6.535 $Y=1.21
c194 42 0 4.58932e-20 $X=4.295 $Y=0.36
c195 40 0 1.27259e-19 $X=3.62 $Y=1.41
c196 36 0 8.56593e-20 $X=2.94 $Y=0.36
c197 28 0 8.64326e-20 $X=4.01 $Y=2.02
c198 22 0 1.07929e-19 $X=6.9 $Y=1.29
r199 63 65 28.4849 $w=2.63e-07 $l=6.55e-07 $layer=LI1_cond $X=2.807 $Y=1.745
+ $X2=2.807 $Y2=1.09
r200 62 63 6.23097 $w=3.73e-07 $l=1.7e-07 $layer=LI1_cond $X=2.752 $Y=1.915
+ $X2=2.752 $Y2=1.745
r201 59 72 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.255 $Y=1.29
+ $X2=7.42 $Y2=1.29
r202 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.255
+ $Y=1.29 $X2=7.255 $Y2=1.29
r203 56 67 14.2244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=7.08 $Y=1.29
+ $X2=6.75 $Y2=1.29
r204 56 58 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=7.08 $Y=1.29
+ $X2=7.255 $Y2=1.29
r205 55 67 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.535 $Y=1.21
+ $X2=6.75 $Y2=1.21
r206 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.45 $Y=1.125
+ $X2=6.535 $Y2=1.21
r207 52 53 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=6.45 $Y=0.425
+ $X2=6.45 $Y2=1.125
r208 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.365 $Y=0.34
+ $X2=6.45 $Y2=0.425
r209 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.365 $Y=0.34
+ $X2=5.695 $Y2=0.34
r210 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.61 $Y=0.425
+ $X2=5.695 $Y2=0.34
r211 48 49 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.61 $Y=0.425
+ $X2=5.61 $Y2=0.79
r212 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.525 $Y=0.875
+ $X2=5.61 $Y2=0.79
r213 46 47 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=5.525 $Y=0.875
+ $X2=4.465 $Y2=0.875
r214 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.38 $Y=0.79
+ $X2=4.465 $Y2=0.875
r215 44 45 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.38 $Y=0.465
+ $X2=4.38 $Y2=0.79
r216 43 66 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.705 $Y=0.36
+ $X2=3.62 $Y2=0.36
r217 42 44 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=4.295 $Y=0.36
+ $X2=4.38 $Y2=0.465
r218 42 43 31.1602 $w=2.08e-07 $l=5.9e-07 $layer=LI1_cond $X=4.295 $Y=0.36
+ $X2=3.705 $Y2=0.36
r219 40 70 68.4659 $w=2.64e-07 $l=3.75e-07 $layer=POLY_cond $X=3.62 $Y=1.41
+ $X2=3.995 $Y2=1.41
r220 40 68 22.822 $w=2.64e-07 $l=1.25e-07 $layer=POLY_cond $X=3.62 $Y=1.41
+ $X2=3.495 $Y2=1.41
r221 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.62
+ $Y=1.41 $X2=3.62 $Y2=1.41
r222 37 66 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.62 $Y=0.465
+ $X2=3.62 $Y2=0.36
r223 37 39 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=3.62 $Y=0.465
+ $X2=3.62 $Y2=1.41
r224 35 66 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=0.36
+ $X2=3.62 $Y2=0.36
r225 35 36 31.4242 $w=2.08e-07 $l=5.95e-07 $layer=LI1_cond $X=3.535 $Y=0.36
+ $X2=2.94 $Y2=0.36
r226 30 65 5.88737 $w=2.93e-07 $l=1.47e-07 $layer=LI1_cond $X=2.792 $Y=0.943
+ $X2=2.792 $Y2=1.09
r227 30 32 14.9622 $w=2.93e-07 $l=3.83e-07 $layer=LI1_cond $X=2.792 $Y=0.943
+ $X2=2.792 $Y2=0.56
r228 29 36 7.07071 $w=2.1e-07 $l=1.93505e-07 $layer=LI1_cond $X=2.792 $Y=0.465
+ $X2=2.94 $Y2=0.36
r229 29 32 3.71126 $w=2.93e-07 $l=9.5e-08 $layer=LI1_cond $X=2.792 $Y=0.465
+ $X2=2.792 $Y2=0.56
r230 25 27 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.675 $Y=1.125
+ $X2=7.675 $Y2=0.805
r231 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.6 $Y=1.2
+ $X2=7.675 $Y2=1.125
r232 23 72 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.6 $Y=1.2 $X2=7.42
+ $Y2=1.2
r233 22 59 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=6.9 $Y=1.29
+ $X2=7.255 $Y2=1.29
r234 17 22 18.0464 $w=4.25e-07 $l=2.05122e-07 $layer=POLY_cond $X=6.81 $Y=1.455
+ $X2=6.9 $Y2=1.29
r235 17 19 390.653 $w=1.8e-07 $l=1.005e-06 $layer=POLY_cond $X=6.81 $Y=1.455
+ $X2=6.81 $Y2=2.46
r236 13 28 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.01 $Y=2.11 $X2=4.01
+ $Y2=2.02
r237 13 15 149.653 $w=1.8e-07 $l=3.85e-07 $layer=POLY_cond $X=4.01 $Y=2.11
+ $X2=4.01 $Y2=2.495
r238 11 70 15.9823 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=1.575
+ $X2=3.995 $Y2=1.41
r239 11 28 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.995 $Y=1.575
+ $X2=3.995 $Y2=2.02
r240 7 68 15.9823 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.495 $Y=1.245
+ $X2=3.495 $Y2=1.41
r241 7 9 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=3.495 $Y=1.245
+ $X2=3.495 $Y2=0.805
r242 2 62 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=2.59
+ $Y=1.735 $X2=2.73 $Y2=1.915
r243 1 32 91 $w=1.7e-07 $l=2.65141e-07 $layer=licon1_NDIFF $count=2 $X=2.55
+ $Y=0.37 $X2=2.73 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTN_1%A_856_294# 1 2 9 13 17 18 21 27 30 31 32 34
+ 36 37
c92 36 0 2.21313e-20 $X=6.11 $Y=2.135
c93 34 0 2.66816e-19 $X=6.03 $Y=1.215
c94 13 0 4.58932e-20 $X=4.535 $Y=0.805
r95 36 38 0.373936 $w=8.33e-07 $l=5e-09 $layer=LI1_cond $X=6.282 $Y=2.135
+ $X2=6.282 $Y2=2.14
r96 36 37 11.6472 $w=8.33e-07 $l=1.65e-07 $layer=LI1_cond $X=6.282 $Y=2.135
+ $X2=6.282 $Y2=1.97
r97 31 41 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.445 $Y=1.635
+ $X2=4.445 $Y2=1.8
r98 31 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.445 $Y=1.635
+ $X2=4.445 $Y2=1.47
r99 30 32 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.445 $Y=1.635
+ $X2=4.445 $Y2=1.47
r100 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.445
+ $Y=1.635 $X2=4.445 $Y2=1.635
r101 27 38 11.3712 $w=7.08e-07 $l=6.75e-07 $layer=LI1_cond $X=6.345 $Y=2.815
+ $X2=6.345 $Y2=2.14
r102 23 34 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=5.95 $Y=1.3
+ $X2=6.03 $Y2=1.215
r103 23 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.95 $Y=1.3
+ $X2=5.95 $Y2=1.97
r104 19 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.03 $Y=1.13
+ $X2=6.03 $Y2=1.215
r105 19 21 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=6.03 $Y=1.13
+ $X2=6.03 $Y2=0.76
r106 17 34 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.865 $Y=1.215
+ $X2=6.03 $Y2=1.215
r107 17 18 81.877 $w=1.68e-07 $l=1.255e-06 $layer=LI1_cond $X=5.865 $Y=1.215
+ $X2=4.61 $Y2=1.215
r108 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.525 $Y=1.3
+ $X2=4.61 $Y2=1.215
r109 15 32 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.525 $Y=1.3
+ $X2=4.525 $Y2=1.47
r110 13 40 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=4.535 $Y=0.805
+ $X2=4.535 $Y2=1.47
r111 9 41 270.153 $w=1.8e-07 $l=6.95e-07 $layer=POLY_cond $X=4.4 $Y=2.495
+ $X2=4.4 $Y2=1.8
r112 2 36 200 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=3 $X=5.97
+ $Y=1.96 $X2=6.11 $Y2=2.135
r113 2 27 200 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=3 $X=5.97
+ $Y=1.96 $X2=6.11 $Y2=2.815
r114 1 21 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=5.89
+ $Y=0.595 $X2=6.03 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTN_1%RESET_B 3 8 9 10 13 18 21 25 27 28 29 30 35
+ 36 38 41 46 47 51 58
c215 41 0 1.78864e-19 $X=0.965 $Y=1.515
r216 51 54 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.545 $Y=1.63
+ $X2=8.545 $Y2=1.795
r217 51 53 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.545 $Y=1.63
+ $X2=8.545 $Y2=1.465
r218 46 49 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.985 $Y=1.635
+ $X2=4.985 $Y2=1.8
r219 46 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.985 $Y=1.635
+ $X2=4.985 $Y2=1.47
r220 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.985
+ $Y=1.635 $X2=4.985 $Y2=1.635
r221 42 58 6.29823 $w=4.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.965 $Y=1.565
+ $X2=1.2 $Y2=1.565
r222 41 44 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.515
+ $X2=0.965 $Y2=1.68
r223 41 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.515
+ $X2=0.965 $Y2=1.35
r224 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.965
+ $Y=1.515 $X2=0.965 $Y2=1.515
r225 38 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=1.665
+ $X2=1.2 $Y2=1.665
r226 36 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.545
+ $Y=1.63 $X2=8.545 $Y2=1.63
r227 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=1.665
+ $X2=8.4 $Y2=1.665
r228 32 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=1.665
+ $X2=5.04 $Y2=1.665
r229 30 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=1.665
+ $X2=5.04 $Y2=1.665
r230 29 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=8.4 $Y2=1.665
r231 29 30 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=8.255 $Y=1.665
+ $X2=5.185 $Y2=1.665
r232 28 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=1.665
+ $X2=1.2 $Y2=1.665
r233 27 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=1.665
+ $X2=5.04 $Y2=1.665
r234 27 28 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=4.895 $Y=1.665
+ $X2=1.345 $Y2=1.665
r235 25 54 371.218 $w=1.8e-07 $l=9.55e-07 $layer=POLY_cond $X=8.62 $Y=2.75
+ $X2=8.62 $Y2=1.795
r236 21 53 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.605 $Y=0.805
+ $X2=8.605 $Y2=1.465
r237 18 49 270.153 $w=1.8e-07 $l=6.95e-07 $layer=POLY_cond $X=4.91 $Y=2.495
+ $X2=4.91 $Y2=1.8
r238 16 18 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=4.91 $Y=3.075
+ $X2=4.91 $Y2=2.495
r239 13 48 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=4.895 $Y=0.805
+ $X2=4.895 $Y2=1.47
r240 9 16 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.82 $Y=3.15
+ $X2=4.91 $Y2=3.075
r241 9 10 1938.26 $w=1.5e-07 $l=3.78e-06 $layer=POLY_cond $X=4.82 $Y=3.15
+ $X2=1.04 $Y2=3.15
r242 8 44 415.919 $w=1.8e-07 $l=1.07e-06 $layer=POLY_cond $X=0.95 $Y=2.75
+ $X2=0.95 $Y2=1.68
r243 6 10 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=0.95 $Y=3.075
+ $X2=1.04 $Y2=3.15
r244 6 8 126.331 $w=1.8e-07 $l=3.25e-07 $layer=POLY_cond $X=0.95 $Y=3.075
+ $X2=0.95 $Y2=2.75
r245 3 43 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=0.915 $Y=0.58
+ $X2=0.915 $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTN_1%A_714_119# 1 2 3 12 16 18 19 22 25 26 27 30
+ 32 34 40
r106 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.53
+ $Y=1.635 $X2=5.53 $Y2=1.635
r107 32 34 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=5.53 $Y=2.02
+ $X2=5.53 $Y2=1.635
r108 28 32 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=5.145 $Y=2.105
+ $X2=5.53 $Y2=2.105
r109 28 30 11.3386 $w=3.08e-07 $l=3.05e-07 $layer=LI1_cond $X=5.145 $Y=2.19
+ $X2=5.145 $Y2=2.495
r110 27 39 13.9941 $w=3.4e-07 $l=4.8695e-07 $layer=LI1_cond $X=4.055 $Y=2.105
+ $X2=3.837 $Y2=2.495
r111 26 28 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.99 $Y=2.105
+ $X2=5.145 $Y2=2.105
r112 26 27 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=4.99 $Y=2.105 $X2=4.055
+ $Y2=2.105
r113 25 27 5.73712 $w=3.4e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.965 $Y=2.02
+ $X2=4.055 $Y2=2.105
r114 25 40 58.2273 $w=1.78e-07 $l=9.45e-07 $layer=LI1_cond $X=3.965 $Y=2.02
+ $X2=3.965 $Y2=1.075
r115 20 40 6.68437 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=4 $Y=0.95 $X2=4
+ $Y2=1.075
r116 20 22 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=4 $Y=0.95 $X2=4
+ $Y2=0.855
r117 18 35 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.74 $Y=1.635
+ $X2=5.53 $Y2=1.635
r118 18 19 3.90195 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=5.74 $Y=1.635
+ $X2=5.855 $Y2=1.635
r119 14 19 34.7346 $w=1.65e-07 $l=1.77059e-07 $layer=POLY_cond $X=5.88 $Y=1.8
+ $X2=5.855 $Y2=1.635
r120 14 16 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=5.88 $Y=1.8
+ $X2=5.88 $Y2=2.46
r121 10 19 34.7346 $w=1.65e-07 $l=1.83916e-07 $layer=POLY_cond $X=5.815 $Y=1.47
+ $X2=5.855 $Y2=1.635
r122 10 12 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.815 $Y=1.47
+ $X2=5.815 $Y2=0.965
r123 3 30 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=5
+ $Y=2.285 $X2=5.135 $Y2=2.495
r124 2 39 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=3.65
+ $Y=2.285 $X2=3.785 $Y2=2.495
r125 1 22 182 $w=1.7e-07 $l=5.03488e-07 $layer=licon1_NDIFF $count=1 $X=3.57
+ $Y=0.595 $X2=3.96 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTN_1%A_300_347# 1 2 7 9 10 12 14 15 16 17 18 21
+ 25 27 32 33 35 36 37 38 44 46 47 51 52 56 57 60 62 65 66
c192 60 0 1.58987e-19 $X=2.42 $Y=1.41
c193 57 0 1.21652e-19 $X=7.475 $Y=1.86
c194 16 0 8.56593e-20 $X=3.08 $Y=0.18
r195 66 77 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.345 $Y=1.635
+ $X2=6.345 $Y2=1.47
r196 65 68 3.0228 $w=3.03e-07 $l=8e-08 $layer=LI1_cond $X=6.357 $Y=1.635
+ $X2=6.357 $Y2=1.715
r197 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.345
+ $Y=1.635 $X2=6.345 $Y2=1.635
r198 61 73 5.302 $w=5e-07 $l=5.5e-08 $layer=POLY_cond $X=2.42 $Y=1.572 $X2=2.475
+ $Y2=1.572
r199 60 63 6.36939 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=1.41
+ $X2=2.325 $Y2=1.575
r200 60 62 6.18336 $w=3.58e-07 $l=1.9e-07 $layer=LI1_cond $X=2.325 $Y=1.41
+ $X2=2.325 $Y2=1.22
r201 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.42
+ $Y=1.41 $X2=2.42 $Y2=1.41
r202 56 57 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.475
+ $Y=1.86 $X2=7.475 $Y2=1.86
r203 54 56 2.76586 $w=2.48e-07 $l=6e-08 $layer=LI1_cond $X=7.435 $Y=1.8
+ $X2=7.435 $Y2=1.86
r204 53 68 4.15824 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=6.51 $Y=1.715
+ $X2=6.357 $Y2=1.715
r205 52 54 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.31 $Y=1.715
+ $X2=7.435 $Y2=1.8
r206 52 53 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=7.31 $Y=1.715
+ $X2=6.51 $Y2=1.715
r207 51 63 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=2.27 $Y=1.82
+ $X2=2.27 $Y2=1.575
r208 48 62 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.31 $Y=1.01
+ $X2=2.31 $Y2=1.22
r209 46 48 7.36389 $w=2e-07 $l=2.09105e-07 $layer=LI1_cond $X=2.145 $Y=0.91
+ $X2=2.31 $Y2=1.01
r210 46 47 15.5273 $w=1.98e-07 $l=2.8e-07 $layer=LI1_cond $X=2.145 $Y=0.91
+ $X2=1.865 $Y2=0.91
r211 42 47 7.39673 $w=2e-07 $l=2.12189e-07 $layer=LI1_cond $X=1.697 $Y=0.81
+ $X2=1.865 $Y2=0.91
r212 42 44 8.60032 $w=3.33e-07 $l=2.5e-07 $layer=LI1_cond $X=1.697 $Y=0.81
+ $X2=1.697 $Y2=0.56
r213 38 51 6.98266 $w=1.9e-07 $l=1.65831e-07 $layer=LI1_cond $X=2.145 $Y=1.915
+ $X2=2.27 $Y2=1.82
r214 38 40 27.1435 $w=1.88e-07 $l=4.65e-07 $layer=LI1_cond $X=2.145 $Y=1.915
+ $X2=1.68 $Y2=1.915
r215 37 57 40.6942 $w=4.1e-07 $l=3e-07 $layer=POLY_cond $X=7.515 $Y=2.16
+ $X2=7.515 $Y2=1.86
r216 33 37 41.944 $w=3.39e-07 $l=3.60278e-07 $layer=POLY_cond $X=7.66 $Y=2.455
+ $X2=7.515 $Y2=2.16
r217 33 35 78.9944 $w=1.8e-07 $l=2.95e-07 $layer=POLY_cond $X=7.66 $Y=2.455
+ $X2=7.66 $Y2=2.75
r218 32 77 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.255 $Y=0.965
+ $X2=6.255 $Y2=1.47
r219 29 32 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.255 $Y=0.255
+ $X2=6.255 $Y2=0.965
r220 28 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.25 $Y=0.18
+ $X2=4.175 $Y2=0.18
r221 27 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.18 $Y=0.18
+ $X2=6.255 $Y2=0.255
r222 27 28 989.638 $w=1.5e-07 $l=1.93e-06 $layer=POLY_cond $X=6.18 $Y=0.18
+ $X2=4.25 $Y2=0.18
r223 23 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.175 $Y=0.255
+ $X2=4.175 $Y2=0.18
r224 23 25 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.175 $Y=0.255
+ $X2=4.175 $Y2=0.805
r225 19 21 217.677 $w=1.8e-07 $l=5.6e-07 $layer=POLY_cond $X=3.56 $Y=1.935
+ $X2=3.56 $Y2=2.495
r226 18 75 33.2496 $w=5e-07 $l=3.23333e-07 $layer=POLY_cond $X=3.08 $Y=1.86
+ $X2=3.005 $Y2=1.572
r227 17 19 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.47 $Y=1.86
+ $X2=3.56 $Y2=1.935
r228 17 18 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.47 $Y=1.86
+ $X2=3.08 $Y2=1.86
r229 15 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.1 $Y=0.18
+ $X2=4.175 $Y2=0.18
r230 15 16 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=4.1 $Y=0.18
+ $X2=3.08 $Y2=0.18
r231 14 75 31.4081 $w=1.5e-07 $l=3.62e-07 $layer=POLY_cond $X=3.005 $Y=1.21
+ $X2=3.005 $Y2=1.572
r232 13 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.005 $Y=0.255
+ $X2=3.08 $Y2=0.18
r233 13 14 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=3.005 $Y=0.255
+ $X2=3.005 $Y2=1.21
r234 10 75 48.682 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.5 $Y=1.572
+ $X2=3.005 $Y2=1.572
r235 10 73 2.41 $w=5e-07 $l=2.5e-08 $layer=POLY_cond $X=2.5 $Y=1.572 $X2=2.475
+ $Y2=1.572
r236 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.5 $Y=1.66
+ $X2=2.5 $Y2=2.235
r237 7 73 31.4081 $w=1.5e-07 $l=3.62e-07 $layer=POLY_cond $X=2.475 $Y=1.21
+ $X2=2.475 $Y2=1.572
r238 7 9 151.027 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.475 $Y=1.21
+ $X2=2.475 $Y2=0.74
r239 2 40 600 $w=1.7e-07 $l=2.54558e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.735 $X2=1.68 $Y2=1.915
r240 1 44 91 $w=1.7e-07 $l=2.61534e-07 $layer=licon1_NDIFF $count=2 $X=1.525
+ $Y=0.37 $X2=1.695 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTN_1%A_1598_93# 1 2 9 13 15 18 22 24 27 28 32
c88 9 0 1.58195e-19 $X=8.065 $Y=0.805
r89 30 32 8.03677 $w=3.78e-07 $l=2.65e-07 $layer=LI1_cond $X=9.21 $Y=0.765
+ $X2=9.475 $Y2=0.765
r90 26 32 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.475 $Y=0.955
+ $X2=9.475 $Y2=0.765
r91 26 27 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=9.475 $Y=0.955
+ $X2=9.475 $Y2=1.965
r92 25 28 6.08426 $w=2.7e-07 $l=2.29619e-07 $layer=LI1_cond $X=9.05 $Y=2.05
+ $X2=8.865 $Y2=2.15
r93 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.39 $Y=2.05
+ $X2=9.475 $Y2=1.965
r94 24 25 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=9.39 $Y=2.05
+ $X2=9.05 $Y2=2.05
r95 20 28 0.630948 $w=3.3e-07 $l=1.94743e-07 $layer=LI1_cond $X=8.845 $Y=2.335
+ $X2=8.865 $Y2=2.15
r96 20 22 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=8.845 $Y=2.335
+ $X2=8.845 $Y2=2.75
r97 18 36 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.155 $Y=2.17
+ $X2=8.155 $Y2=2.335
r98 18 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.155 $Y=2.17
+ $X2=8.155 $Y2=2.005
r99 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.155
+ $Y=2.17 $X2=8.155 $Y2=2.17
r100 15 28 6.08426 $w=2.7e-07 $l=1.85e-07 $layer=LI1_cond $X=8.68 $Y=2.15
+ $X2=8.865 $Y2=2.15
r101 15 17 16.3522 $w=3.68e-07 $l=5.25e-07 $layer=LI1_cond $X=8.68 $Y=2.15
+ $X2=8.155 $Y2=2.15
r102 13 36 161.315 $w=1.8e-07 $l=4.15e-07 $layer=POLY_cond $X=8.08 $Y=2.75
+ $X2=8.08 $Y2=2.335
r103 9 35 615.319 $w=1.5e-07 $l=1.2e-06 $layer=POLY_cond $X=8.065 $Y=0.805
+ $X2=8.065 $Y2=2.005
r104 2 22 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=8.71
+ $Y=2.54 $X2=8.845 $Y2=2.75
r105 1 30 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=9.07
+ $Y=0.595 $X2=9.21 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTN_1%A_1266_119# 1 2 7 9 10 12 14 16 18 20 21 23
+ 25 28 32 37 39 40 45 47 49 50
c131 47 0 2.64234e-19 $X=7.815 $Y=1.21
r132 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.085
+ $Y=1.29 $X2=9.085 $Y2=1.29
r133 45 46 20.5133 $w=2.26e-07 $l=3.8e-07 $layer=LI1_cond $X=7.435 $Y=2.7
+ $X2=7.815 $Y2=2.7
r134 41 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=1.21
+ $X2=7.815 $Y2=1.21
r135 40 49 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=8.92 $Y=1.21
+ $X2=9.07 $Y2=1.21
r136 40 41 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=8.92 $Y=1.21
+ $X2=7.9 $Y2=1.21
r137 39 46 2.4068 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.815 $Y=2.535
+ $X2=7.815 $Y2=2.7
r138 38 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=1.295
+ $X2=7.815 $Y2=1.21
r139 38 39 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=7.815 $Y=1.295
+ $X2=7.815 $Y2=2.535
r140 37 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.815 $Y=1.125
+ $X2=7.815 $Y2=1.21
r141 36 37 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.815 $Y=0.955
+ $X2=7.815 $Y2=1.125
r142 32 45 1.22073 $w=3.3e-07 $l=1.75152e-07 $layer=LI1_cond $X=7.435 $Y=2.7
+ $X2=7.435 $Y2=2.7
r143 32 34 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=7.435 $Y=2.7 $X2=7.035
+ $Y2=2.7
r144 28 36 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.73 $Y=0.79
+ $X2=7.815 $Y2=0.955
r145 28 30 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=7.73 $Y=0.79
+ $X2=7.46 $Y2=0.79
r146 26 50 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=9.085 $Y=1.63
+ $X2=9.085 $Y2=1.29
r147 26 27 50.3824 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=9.085 $Y=1.63
+ $X2=9.085 $Y2=1.97
r148 24 50 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=9.085 $Y=1.275
+ $X2=9.085 $Y2=1.29
r149 24 25 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=9.085 $Y=1.275
+ $X2=9.085 $Y2=1.2
r150 21 23 122.107 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=10.03 $Y=1.125
+ $X2=10.03 $Y2=0.745
r151 18 20 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=10.04 $Y=2.045
+ $X2=10.04 $Y2=2.54
r152 17 27 18.414 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.25 $Y=1.97
+ $X2=9.085 $Y2=1.97
r153 16 18 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=9.95 $Y=1.97
+ $X2=10.04 $Y2=2.045
r154 16 17 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=9.95 $Y=1.97 $X2=9.25
+ $Y2=1.97
r155 15 25 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.25 $Y=1.2
+ $X2=9.085 $Y2=1.2
r156 14 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.955 $Y=1.2
+ $X2=10.03 $Y2=1.125
r157 14 15 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=9.955 $Y=1.2
+ $X2=9.25 $Y2=1.2
r158 10 27 19.4594 $w=2.93e-07 $l=8.21584e-08 $layer=POLY_cond $X=9.07 $Y=2.045
+ $X2=9.085 $Y2=1.97
r159 10 12 274.04 $w=1.8e-07 $l=7.05e-07 $layer=POLY_cond $X=9.07 $Y=2.045
+ $X2=9.07 $Y2=2.75
r160 7 25 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.995 $Y=1.125
+ $X2=9.085 $Y2=1.2
r161 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.995 $Y=1.125
+ $X2=8.995 $Y2=0.805
r162 2 45 600 $w=1.7e-07 $l=9.71339e-07 $layer=licon1_PDIFF $count=1 $X=6.9
+ $Y=1.96 $X2=7.435 $Y2=2.7
r163 2 34 600 $w=1.7e-07 $l=8.04674e-07 $layer=licon1_PDIFF $count=1 $X=6.9
+ $Y=1.96 $X2=7.035 $Y2=2.7
r164 1 30 91 $w=1.7e-07 $l=1.22362e-06 $layer=licon1_NDIFF $count=2 $X=6.33
+ $Y=0.595 $X2=7.46 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTN_1%A_1934_94# 1 2 9 13 14 16 20 25 28 29 32 34
r62 29 35 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.48 $Y=1.485
+ $X2=10.48 $Y2=1.65
r63 29 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.48 $Y=1.485
+ $X2=10.48 $Y2=1.32
r64 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.48
+ $Y=1.485 $X2=10.48 $Y2=1.485
r65 26 32 0.364692 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=9.98 $Y=1.485
+ $X2=9.855 $Y2=1.485
r66 26 28 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=9.98 $Y=1.485
+ $X2=10.48 $Y2=1.485
r67 25 31 1.61342 $w=2.48e-07 $l=3.5e-08 $layer=LI1_cond $X=9.855 $Y=2.27
+ $X2=9.855 $Y2=2.305
r68 22 32 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=9.855 $Y=1.65
+ $X2=9.855 $Y2=1.485
r69 22 25 28.5806 $w=2.48e-07 $l=6.2e-07 $layer=LI1_cond $X=9.855 $Y=1.65
+ $X2=9.855 $Y2=2.27
r70 18 32 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=9.855 $Y=1.32
+ $X2=9.855 $Y2=1.485
r71 18 20 26.5062 $w=2.48e-07 $l=5.75e-07 $layer=LI1_cond $X=9.855 $Y=1.32
+ $X2=9.855 $Y2=0.745
r72 14 31 6.46688 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.815 $Y=2.47
+ $X2=9.815 $Y2=2.305
r73 14 16 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=9.815 $Y=2.47
+ $X2=9.815 $Y2=2.815
r74 13 34 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=10.54 $Y=0.84
+ $X2=10.54 $Y2=1.32
r75 9 35 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=10.545 $Y=2.4
+ $X2=10.545 $Y2=1.65
r76 2 25 600 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=9.69
+ $Y=2.12 $X2=9.815 $Y2=2.27
r77 2 16 600 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_PDIFF $count=1 $X=9.69
+ $Y=2.12 $X2=9.815 $Y2=2.815
r78 1 20 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=9.67
+ $Y=0.47 $X2=9.815 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTN_1%VPWR 1 2 3 4 5 6 7 8 25 27 31 35 39 41 45 49
+ 53 57 60 61 63 64 65 67 72 77 89 98 99 105 108 111 114 117
c128 31 0 4.19395e-20 $X=1.18 $Y=2.75
r129 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r130 111 112 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r131 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r132 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r133 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r134 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r135 96 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.8 $Y2=3.33
r136 96 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r137 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r138 93 117 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.46 $Y=3.33
+ $X2=9.335 $Y2=3.33
r139 93 95 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.46 $Y=3.33
+ $X2=9.84 $Y2=3.33
r140 92 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r141 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r142 89 117 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.21 $Y=3.33
+ $X2=9.335 $Y2=3.33
r143 89 91 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.21 $Y=3.33
+ $X2=8.88 $Y2=3.33
r144 88 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r145 87 88 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r146 85 88 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=7.92 $Y2=3.33
r147 84 87 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=7.92
+ $Y2=3.33
r148 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r149 82 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.82 $Y=3.33
+ $X2=5.655 $Y2=3.33
r150 82 84 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.82 $Y=3.33 $X2=6
+ $Y2=3.33
r151 81 112 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.56 $Y2=3.33
r152 81 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r153 80 81 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r154 78 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=3.33
+ $X2=2.21 $Y2=3.33
r155 78 80 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.375 $Y=3.33
+ $X2=2.64 $Y2=3.33
r156 77 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.49 $Y=3.33
+ $X2=4.655 $Y2=3.33
r157 77 80 120.695 $w=1.68e-07 $l=1.85e-06 $layer=LI1_cond $X=4.49 $Y=3.33
+ $X2=2.64 $Y2=3.33
r158 76 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r159 76 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r160 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r161 73 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.39 $Y=3.33
+ $X2=1.225 $Y2=3.33
r162 73 75 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.39 $Y=3.33
+ $X2=1.68 $Y2=3.33
r163 72 108 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.045 $Y=3.33
+ $X2=2.21 $Y2=3.33
r164 72 75 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.045 $Y=3.33
+ $X2=1.68 $Y2=3.33
r165 71 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r166 71 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r167 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r168 68 102 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=3.33 $X2=0.22
+ $Y2=3.33
r169 68 70 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r170 67 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.06 $Y=3.33
+ $X2=1.225 $Y2=3.33
r171 67 70 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.06 $Y=3.33
+ $X2=0.72 $Y2=3.33
r172 65 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r173 65 112 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r174 65 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r175 63 95 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.15 $Y=3.33
+ $X2=9.84 $Y2=3.33
r176 63 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.15 $Y=3.33
+ $X2=10.275 $Y2=3.33
r177 62 98 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=10.4 $Y=3.33 $X2=10.8
+ $Y2=3.33
r178 62 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.4 $Y=3.33
+ $X2=10.275 $Y2=3.33
r179 60 87 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.14 $Y=3.33
+ $X2=7.92 $Y2=3.33
r180 60 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.14 $Y=3.33
+ $X2=8.305 $Y2=3.33
r181 59 91 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=8.47 $Y=3.33
+ $X2=8.88 $Y2=3.33
r182 59 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.47 $Y=3.33
+ $X2=8.305 $Y2=3.33
r183 55 64 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.275 $Y=3.245
+ $X2=10.275 $Y2=3.33
r184 55 57 45.1758 $w=2.48e-07 $l=9.8e-07 $layer=LI1_cond $X=10.275 $Y=3.245
+ $X2=10.275 $Y2=2.265
r185 51 117 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.335 $Y=3.245
+ $X2=9.335 $Y2=3.33
r186 51 53 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=9.335 $Y=3.245
+ $X2=9.335 $Y2=2.75
r187 47 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.305 $Y=3.245
+ $X2=8.305 $Y2=3.33
r188 47 49 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=8.305 $Y=3.245
+ $X2=8.305 $Y2=2.75
r189 43 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.655 $Y=3.245
+ $X2=5.655 $Y2=3.33
r190 43 45 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=5.655 $Y=3.245
+ $X2=5.655 $Y2=2.445
r191 42 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.82 $Y=3.33
+ $X2=4.655 $Y2=3.33
r192 41 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.49 $Y=3.33
+ $X2=5.655 $Y2=3.33
r193 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.49 $Y=3.33
+ $X2=4.82 $Y2=3.33
r194 37 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.655 $Y=3.245
+ $X2=4.655 $Y2=3.33
r195 37 39 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=4.655 $Y=3.245
+ $X2=4.655 $Y2=2.495
r196 33 108 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.21 $Y=3.245
+ $X2=2.21 $Y2=3.33
r197 33 35 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=2.21 $Y=3.245
+ $X2=2.21 $Y2=2.635
r198 29 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=3.245
+ $X2=1.225 $Y2=3.33
r199 29 31 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.225 $Y=3.245
+ $X2=1.225 $Y2=2.75
r200 25 102 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.22 $Y2=3.33
r201 25 27 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.275 $Y2=2.75
r202 8 57 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=10.13
+ $Y=2.12 $X2=10.315 $Y2=2.265
r203 7 53 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=9.16
+ $Y=2.54 $X2=9.295 $Y2=2.75
r204 6 49 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=8.17
+ $Y=2.54 $X2=8.305 $Y2=2.75
r205 5 45 300 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_PDIFF $count=2 $X=5.53
+ $Y=1.96 $X2=5.655 $Y2=2.445
r206 4 39 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=4.49
+ $Y=2.285 $X2=4.655 $Y2=2.495
r207 3 35 600 $w=1.7e-07 $l=9.97246e-07 $layer=licon1_PDIFF $count=1 $X=2.005
+ $Y=1.735 $X2=2.21 $Y2=2.635
r208 2 31 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.04
+ $Y=2.54 $X2=1.18 $Y2=2.75
r209 1 27 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.275 $Y2=2.75
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTN_1%A_33_74# 1 2 3 4 14 17 19 23 25 26 29 34 36
+ 38
c85 25 0 2.13692e-19 $X=3.277 $Y=2.002
c86 14 0 1.52323e-19 $X=0.625 $Y=2.18
r87 32 34 8.25044 $w=4.38e-07 $l=3.15e-07 $layer=LI1_cond $X=0.31 $Y=0.57
+ $X2=0.625 $Y2=0.57
r88 27 38 3.66998 $w=2.97e-07 $l=1.13137e-07 $layer=LI1_cond $X=3.305 $Y=2.38
+ $X2=3.277 $Y2=2.28
r89 27 29 4.90855 $w=2.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.305 $Y=2.38
+ $X2=3.305 $Y2=2.495
r90 26 38 3.66998 $w=2.97e-07 $l=1e-07 $layer=LI1_cond $X=3.277 $Y=2.18
+ $X2=3.277 $Y2=2.28
r91 25 37 6.38767 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=3.277 $Y=2.002
+ $X2=3.277 $Y2=1.84
r92 25 26 6.31184 $w=3.23e-07 $l=1.78e-07 $layer=LI1_cond $X=3.277 $Y=2.002
+ $X2=3.277 $Y2=2.18
r93 23 37 47.9416 $w=2.48e-07 $l=1.04e-06 $layer=LI1_cond $X=3.24 $Y=0.8
+ $X2=3.24 $Y2=1.84
r94 20 36 1.51883 $w=2e-07 $l=3.96863e-07 $layer=LI1_cond $X=0.89 $Y=2.28
+ $X2=0.54 $Y2=2.18
r95 19 38 2.80448 $w=2e-07 $l=1.62e-07 $layer=LI1_cond $X=3.115 $Y=2.28
+ $X2=3.277 $Y2=2.28
r96 19 20 123.386 $w=1.98e-07 $l=2.225e-06 $layer=LI1_cond $X=3.115 $Y=2.28
+ $X2=0.89 $Y2=2.28
r97 15 36 4.95952 $w=2.1e-07 $l=3.09233e-07 $layer=LI1_cond $X=0.765 $Y=2.38
+ $X2=0.54 $Y2=2.18
r98 15 17 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.765 $Y=2.38
+ $X2=0.765 $Y2=2.75
r99 14 36 4.95952 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.625 $Y=2.18
+ $X2=0.54 $Y2=2.18
r100 13 34 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.625 $Y=0.79
+ $X2=0.625 $Y2=0.57
r101 13 14 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=0.625 $Y=0.79
+ $X2=0.625 $Y2=2.18
r102 4 29 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=3.19
+ $Y=2.285 $X2=3.335 $Y2=2.495
r103 3 17 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=2.54 $X2=0.725 $Y2=2.75
r104 2 23 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=3.155
+ $Y=0.595 $X2=3.28 $Y2=0.8
r105 1 32 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=0.165
+ $Y=0.37 $X2=0.31 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTN_1%Q 1 2 9 13 14 15 16 23 32
r28 21 23 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=10.78 $Y=1.995
+ $X2=10.78 $Y2=2.035
r29 15 16 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=10.78 $Y=2.405
+ $X2=10.78 $Y2=2.775
r30 14 21 0.75732 $w=3.48e-07 $l=2.3e-08 $layer=LI1_cond $X=10.78 $Y=1.972
+ $X2=10.78 $Y2=1.995
r31 14 32 8.06043 $w=3.48e-07 $l=1.52e-07 $layer=LI1_cond $X=10.78 $Y=1.972
+ $X2=10.78 $Y2=1.82
r32 14 15 11.4586 $w=3.48e-07 $l=3.48e-07 $layer=LI1_cond $X=10.78 $Y=2.057
+ $X2=10.78 $Y2=2.405
r33 14 23 0.724393 $w=3.48e-07 $l=2.2e-08 $layer=LI1_cond $X=10.78 $Y=2.057
+ $X2=10.78 $Y2=2.035
r34 13 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.87 $Y=1.15
+ $X2=10.87 $Y2=1.82
r35 7 13 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=10.772 $Y=0.968
+ $X2=10.772 $Y2=1.15
r36 7 9 11.4613 $w=3.63e-07 $l=3.63e-07 $layer=LI1_cond $X=10.772 $Y=0.968
+ $X2=10.772 $Y2=0.605
r37 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.635
+ $Y=1.84 $X2=10.77 $Y2=1.985
r38 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.635
+ $Y=1.84 $X2=10.77 $Y2=2.815
r39 1 9 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=10.615
+ $Y=0.47 $X2=10.755 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_MS__DFRTN_1%VGND 1 2 3 4 5 18 22 26 30 34 37 38 39 45 49
+ 54 62 72 73 76 79 82 85
r109 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r110 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r111 79 80 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r112 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r113 73 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r114 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r115 70 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.41 $Y=0
+ $X2=10.285 $Y2=0
r116 70 72 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=10.41 $Y=0 $X2=10.8
+ $Y2=0
r117 69 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r118 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r119 66 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r120 66 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r121 65 68 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r122 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r123 63 82 10.4332 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=8.555 $Y=0 $X2=8.335
+ $Y2=0
r124 63 65 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.555 $Y=0
+ $X2=8.88 $Y2=0
r125 62 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.16 $Y=0
+ $X2=10.285 $Y2=0
r126 62 68 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=10.16 $Y=0 $X2=9.84
+ $Y2=0
r127 61 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r128 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r129 57 60 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=7.92
+ $Y2=0
r130 55 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.355 $Y=0 $X2=5.19
+ $Y2=0
r131 55 57 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.355 $Y=0
+ $X2=5.52 $Y2=0
r132 54 82 10.4332 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=8.115 $Y=0 $X2=8.335
+ $Y2=0
r133 54 60 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=8.115 $Y=0
+ $X2=7.92 $Y2=0
r134 53 80 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=5.04
+ $Y2=0
r135 53 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r136 52 53 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r137 50 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=0 $X2=2.2
+ $Y2=0
r138 50 52 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.365 $Y=0
+ $X2=2.64 $Y2=0
r139 49 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.025 $Y=0 $X2=5.19
+ $Y2=0
r140 49 52 155.599 $w=1.68e-07 $l=2.385e-06 $layer=LI1_cond $X=5.025 $Y=0
+ $X2=2.64 $Y2=0
r141 48 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r142 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r143 45 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=0 $X2=2.2
+ $Y2=0
r144 45 47 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.035 $Y=0
+ $X2=1.68 $Y2=0
r145 43 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r146 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r147 39 61 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=5.52 $Y=0 $X2=7.92
+ $Y2=0
r148 39 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r149 39 57 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r150 37 42 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=0
+ $X2=0.72 $Y2=0
r151 37 38 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.145
+ $Y2=0
r152 36 47 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.245 $Y=0
+ $X2=1.68 $Y2=0
r153 36 38 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.245 $Y=0 $X2=1.145
+ $Y2=0
r154 32 85 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.285 $Y=0.085
+ $X2=10.285 $Y2=0
r155 32 34 23.9708 $w=2.48e-07 $l=5.2e-07 $layer=LI1_cond $X=10.285 $Y=0.085
+ $X2=10.285 $Y2=0.605
r156 28 82 1.73497 $w=4.4e-07 $l=8.5e-08 $layer=LI1_cond $X=8.335 $Y=0.085
+ $X2=8.335 $Y2=0
r157 28 30 17.1557 $w=4.38e-07 $l=6.55e-07 $layer=LI1_cond $X=8.335 $Y=0.085
+ $X2=8.335 $Y2=0.74
r158 24 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.19 $Y=0.085
+ $X2=5.19 $Y2=0
r159 24 26 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=5.19 $Y=0.085
+ $X2=5.19 $Y2=0.535
r160 20 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=0.085 $X2=2.2
+ $Y2=0
r161 20 22 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.2 $Y=0.085
+ $X2=2.2 $Y2=0.535
r162 16 38 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=0.085
+ $X2=1.145 $Y2=0
r163 16 18 27.45 $w=1.98e-07 $l=4.95e-07 $layer=LI1_cond $X=1.145 $Y=0.085
+ $X2=1.145 $Y2=0.58
r164 5 34 91 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_NDIFF $count=2 $X=10.105
+ $Y=0.47 $X2=10.325 $Y2=0.605
r165 4 30 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=8.14
+ $Y=0.595 $X2=8.335 $Y2=0.74
r166 3 26 182 $w=1.7e-07 $l=2.48193e-07 $layer=licon1_NDIFF $count=1 $X=4.97
+ $Y=0.595 $X2=5.19 $Y2=0.535
r167 2 22 182 $w=1.7e-07 $l=2.64953e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.37 $X2=2.2 $Y2=0.535
r168 1 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.99
+ $Y=0.37 $X2=1.13 $Y2=0.58
.ends


* File: sky130_fd_sc_ms__dfstp_2.pex.spice
* Created: Wed Sep  2 12:03:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DFSTP_2%D 2 5 9 11 12 16 17 20
c33 17 0 1.14039e-19 $X=0.64 $Y=1.145
r34 20 22 39.7991 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.825
+ $X2=0.61 $Y2=1.99
r35 20 21 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.825 $X2=0.64 $Y2=1.825
r36 16 18 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.145
+ $X2=0.61 $Y2=0.98
r37 16 17 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.145 $X2=0.64 $Y2=1.145
r38 12 21 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=0.64 $Y=1.665
+ $X2=0.64 $Y2=1.825
r39 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.665
r40 11 17 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.145
r41 9 18 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.495 $Y=0.58 $X2=0.495
+ $Y2=0.98
r42 5 22 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=0.505 $Y=2.75
+ $X2=0.505 $Y2=1.99
r43 2 20 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=0.61 $Y=1.795 $X2=0.61
+ $Y2=1.825
r44 1 16 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=0.61 $Y=1.175 $X2=0.61
+ $Y2=1.145
r45 1 2 88.4142 $w=3.9e-07 $l=6.2e-07 $layer=POLY_cond $X=0.61 $Y=1.175 $X2=0.61
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_2%CLK 3 6 8 11 13
c39 11 0 9.68091e-20 $X=1.465 $Y=1.385
c40 6 0 1.14039e-19 $X=1.515 $Y=2.35
r41 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.385
+ $X2=1.465 $Y2=1.55
r42 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.385
+ $X2=1.465 $Y2=1.22
r43 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.465
+ $Y=1.385 $X2=1.465 $Y2=1.385
r44 8 12 6.69663 $w=3.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.68 $Y=1.365
+ $X2=1.465 $Y2=1.365
r45 6 14 310.968 $w=1.8e-07 $l=8e-07 $layer=POLY_cond $X=1.515 $Y=2.35 $X2=1.515
+ $Y2=1.55
r46 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.485 $Y=0.74
+ $X2=1.485 $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_2%A_398_74# 1 2 7 8 11 13 15 17 21 24 26 29 33
+ 35 36 37 38 41 48 52 53 56 57 58 60 61 62 64 66 67 68 70 71 72 76 77 81 85
c265 81 0 1.55697e-19 $X=7.455 $Y=2.215
c266 77 0 1.63034e-19 $X=6.795 $Y=1.285
c267 72 0 2.15866e-20 $X=3.77 $Y=2.325
c268 62 0 5.12754e-20 $X=5.69 $Y=2.405
c269 24 0 1.76198e-19 $X=7.53 $Y=2.75
c270 15 0 1.99877e-19 $X=3.83 $Y=1.38
c271 11 0 8.11169e-20 $X=3.005 $Y=2.49
r272 81 89 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.455 $Y=2.215
+ $X2=7.455 $Y2=2.38
r273 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.455
+ $Y=2.215 $X2=7.455 $Y2=2.215
r274 77 85 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.795 $Y=1.285
+ $X2=6.795 $Y2=1.12
r275 76 77 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.795
+ $Y=1.285 $X2=6.795 $Y2=1.285
r276 73 76 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.5 $Y=1.285
+ $X2=6.795 $Y2=1.285
r277 70 80 11.5534 $w=3.29e-07 $l=2.8058e-07 $layer=LI1_cond $X=7.575 $Y=1.98
+ $X2=7.475 $Y2=2.215
r278 69 70 99.8182 $w=1.68e-07 $l=1.53e-06 $layer=LI1_cond $X=7.575 $Y=0.45
+ $X2=7.575 $Y2=1.98
r279 67 69 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.49 $Y=0.365
+ $X2=7.575 $Y2=0.45
r280 67 68 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=7.49 $Y=0.365
+ $X2=6.585 $Y2=0.365
r281 65 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.5 $Y=1.45 $X2=6.5
+ $Y2=1.285
r282 65 66 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=6.5 $Y=1.45 $X2=6.5
+ $Y2=2.32
r283 64 73 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.5 $Y=1.12 $X2=6.5
+ $Y2=1.285
r284 63 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.5 $Y=0.45
+ $X2=6.585 $Y2=0.365
r285 63 64 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.5 $Y=0.45 $X2=6.5
+ $Y2=1.12
r286 61 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.415 $Y=2.405
+ $X2=6.5 $Y2=2.32
r287 61 62 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=6.415 $Y=2.405
+ $X2=5.69 $Y2=2.405
r288 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.605 $Y=2.49
+ $X2=5.69 $Y2=2.405
r289 59 60 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=5.605 $Y=2.49
+ $X2=5.605 $Y2=2.89
r290 57 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.52 $Y=2.975
+ $X2=5.605 $Y2=2.89
r291 57 58 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=5.52 $Y=2.975
+ $X2=4.915 $Y2=2.975
r292 56 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.83 $Y=2.89
+ $X2=4.915 $Y2=2.975
r293 55 56 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.83 $Y=2.41
+ $X2=4.83 $Y2=2.89
r294 54 72 2.45049 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.915 $Y=2.325
+ $X2=3.77 $Y2=2.325
r295 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.745 $Y=2.325
+ $X2=4.83 $Y2=2.41
r296 53 54 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=4.745 $Y=2.325
+ $X2=3.915 $Y2=2.325
r297 51 72 3.98977 $w=2.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=3.71 $Y=2.41
+ $X2=3.77 $Y2=2.325
r298 51 52 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.71 $Y=2.41
+ $X2=3.71 $Y2=2.89
r299 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.77
+ $Y=1.545 $X2=3.77 $Y2=1.545
r300 46 72 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.77 $Y=2.24
+ $X2=3.77 $Y2=2.325
r301 46 48 27.6189 $w=2.88e-07 $l=6.95e-07 $layer=LI1_cond $X=3.77 $Y=2.24
+ $X2=3.77 $Y2=1.545
r302 44 71 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=3.03 $Y=0.425
+ $X2=3.03 $Y2=1.38
r303 41 71 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.95 $Y=1.545
+ $X2=2.95 $Y2=1.38
r304 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.95
+ $Y=1.545 $X2=2.95 $Y2=1.545
r305 37 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.625 $Y=2.975
+ $X2=3.71 $Y2=2.89
r306 37 38 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=3.625 $Y=2.975
+ $X2=2.275 $Y2=2.975
r307 35 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.945 $Y=0.34
+ $X2=3.03 $Y2=0.425
r308 35 36 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.945 $Y=0.34
+ $X2=2.215 $Y2=0.34
r309 31 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.19 $Y=2.89
+ $X2=2.275 $Y2=2.975
r310 31 33 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.19 $Y=2.89
+ $X2=2.19 $Y2=2.665
r311 27 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.13 $Y=0.425
+ $X2=2.215 $Y2=0.34
r312 27 29 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.13 $Y=0.425
+ $X2=2.13 $Y2=0.515
r313 24 89 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=7.53 $Y=2.75
+ $X2=7.53 $Y2=2.38
r314 21 85 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.705 $Y=0.69
+ $X2=6.705 $Y2=1.12
r315 15 49 21.4517 $w=1.5e-07 $l=1.72337e-07 $layer=POLY_cond $X=3.83 $Y=1.38
+ $X2=3.845 $Y2=1.545
r316 15 17 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.83 $Y=1.38 $X2=3.83
+ $Y2=0.58
r317 14 42 13.4654 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.115 $Y=1.545
+ $X2=2.95 $Y2=1.545
r318 13 49 10.7258 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.755 $Y=1.545
+ $X2=3.845 $Y2=1.545
r319 13 14 111.911 $w=3.3e-07 $l=6.4e-07 $layer=POLY_cond $X=3.755 $Y=1.545
+ $X2=3.115 $Y2=1.545
r320 11 26 171.032 $w=1.8e-07 $l=4.4e-07 $layer=POLY_cond $X=3.005 $Y=2.49
+ $X2=3.005 $Y2=2.05
r321 8 26 38.198 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.885
+ $X2=2.95 $Y2=2.05
r322 7 42 13.4654 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.95 $Y=1.71
+ $X2=2.95 $Y2=1.545
r323 7 8 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=2.95 $Y=1.71
+ $X2=2.95 $Y2=1.885
r324 2 33 600 $w=1.7e-07 $l=9.4008e-07 $layer=licon1_PDIFF $count=1 $X=2.055
+ $Y=1.79 $X2=2.19 $Y2=2.665
r325 1 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.99
+ $Y=0.37 $X2=2.13 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_2%A_767_384# 1 2 9 11 12 13 15 18 21 26 31 32
+ 35 39
c78 39 0 1.05311e-20 $X=4.485 $Y=1.065
c79 31 0 1.66427e-19 $X=5.265 $Y=2.52
c80 9 0 1.89547e-19 $X=3.925 $Y=2.49
r81 31 32 10.1743 $w=2.63e-07 $l=2e-07 $layer=LI1_cond $X=5.217 $Y=2.52
+ $X2=5.217 $Y2=2.32
r82 27 39 17.4217 $w=2.49e-07 $l=9e-08 $layer=POLY_cond $X=4.575 $Y=1.065
+ $X2=4.485 $Y2=1.065
r83 26 29 12.2584 $w=4.18e-07 $l=4.2e-07 $layer=LI1_cond $X=4.575 $Y=0.9
+ $X2=4.995 $Y2=0.9
r84 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.575
+ $Y=1.065 $X2=4.575 $Y2=1.065
r85 23 32 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.17 $Y=2.07
+ $X2=5.17 $Y2=2.32
r86 21 36 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.395 $Y=1.905
+ $X2=4.395 $Y2=1.995
r87 21 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.395 $Y=1.905
+ $X2=4.395 $Y2=1.74
r88 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.395
+ $Y=1.905 $X2=4.395 $Y2=1.905
r89 18 23 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.085 $Y=1.905
+ $X2=5.17 $Y2=2.07
r90 18 20 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=5.085 $Y=1.905
+ $X2=4.395 $Y2=1.905
r91 16 39 14.627 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.485 $Y=1.23
+ $X2=4.485 $Y2=1.065
r92 16 35 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.485 $Y=1.23
+ $X2=4.485 $Y2=1.74
r93 13 39 51.2972 $w=2.49e-07 $l=3.37565e-07 $layer=POLY_cond $X=4.22 $Y=0.9
+ $X2=4.485 $Y2=1.065
r94 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.22 $Y=0.9 $X2=4.22
+ $Y2=0.58
r95 11 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.23 $Y=1.995
+ $X2=4.395 $Y2=1.995
r96 11 12 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=4.23 $Y=1.995
+ $X2=4.015 $Y2=1.995
r97 7 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.925 $Y=2.07
+ $X2=4.015 $Y2=1.995
r98 7 9 163.258 $w=1.8e-07 $l=4.2e-07 $layer=POLY_cond $X=3.925 $Y=2.07
+ $X2=3.925 $Y2=2.49
r99 2 31 600 $w=1.7e-07 $l=3e-07 $layer=licon1_PDIFF $count=1 $X=5.13 $Y=2.28
+ $X2=5.265 $Y2=2.52
r100 1 29 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=4.85
+ $Y=0.59 $X2=4.995 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_2%A_612_74# 1 2 9 13 17 21 25 29 32 34 36 38
+ 39 41 45 47 49 54 59
c133 47 0 1.63034e-19 $X=6.08 $Y=1.38
c134 39 0 1.89547e-19 $X=3.285 $Y=2.26
c135 36 0 1.05311e-20 $X=5.125 $Y=1.395
c136 32 0 1.99877e-19 $X=4.17 $Y=1.4
c137 9 0 5.12754e-20 $X=5.04 $Y=2.49
r138 58 59 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=6.255 $Y=1.38
+ $X2=6.315 $Y2=1.38
r139 48 58 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=6.08 $Y=1.38
+ $X2=6.255 $Y2=1.38
r140 47 49 5.35643 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=6.08 $Y=1.392
+ $X2=5.915 $Y2=1.392
r141 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.08
+ $Y=1.38 $X2=6.08 $Y2=1.38
r142 44 54 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=5.115 $Y=1.385
+ $X2=5.21 $Y2=1.385
r143 44 51 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.115 $Y=1.385
+ $X2=5.04 $Y2=1.385
r144 43 45 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.115 $Y=1.395
+ $X2=4.95 $Y2=1.395
r145 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.115
+ $Y=1.385 $X2=5.115 $Y2=1.385
r146 38 39 10.6751 $w=3.38e-07 $l=2.3e-07 $layer=LI1_cond $X=3.285 $Y=2.49
+ $X2=3.285 $Y2=2.26
r147 36 43 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=5.125 $Y=1.395
+ $X2=5.115 $Y2=1.395
r148 36 49 26.0123 $w=3.48e-07 $l=7.9e-07 $layer=LI1_cond $X=5.125 $Y=1.395
+ $X2=5.915 $Y2=1.395
r149 34 45 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.255 $Y=1.485
+ $X2=4.95 $Y2=1.485
r150 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.17 $Y=1.4
+ $X2=4.255 $Y2=1.485
r151 31 32 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.17 $Y=1.21
+ $X2=4.17 $Y2=1.4
r152 30 41 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=1.125
+ $X2=3.45 $Y2=1.125
r153 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.085 $Y=1.125
+ $X2=4.17 $Y2=1.21
r154 29 30 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=4.085 $Y=1.125
+ $X2=3.615 $Y2=1.125
r155 27 41 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.37 $Y=1.21
+ $X2=3.45 $Y2=1.125
r156 27 39 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=3.37 $Y=1.21
+ $X2=3.37 $Y2=2.26
r157 23 41 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.45 $Y=1.04
+ $X2=3.45 $Y2=1.125
r158 23 25 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=3.45 $Y=1.04
+ $X2=3.45 $Y2=0.585
r159 19 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.315 $Y=1.215
+ $X2=6.315 $Y2=1.38
r160 19 21 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=6.315 $Y=1.215
+ $X2=6.315 $Y2=0.69
r161 15 58 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.255 $Y=1.545
+ $X2=6.255 $Y2=1.38
r162 15 17 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=6.255 $Y=1.545
+ $X2=6.255 $Y2=2.205
r163 11 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.21 $Y=1.22
+ $X2=5.21 $Y2=1.385
r164 11 13 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=5.21 $Y=1.22
+ $X2=5.21 $Y2=0.8
r165 7 51 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.04 $Y=1.55
+ $X2=5.04 $Y2=1.385
r166 7 9 365.387 $w=1.8e-07 $l=9.4e-07 $layer=POLY_cond $X=5.04 $Y=1.55 $X2=5.04
+ $Y2=2.49
r167 2 38 600 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_PDIFF $count=1 $X=3.095
+ $Y=2.28 $X2=3.28 $Y2=2.49
r168 1 25 182 $w=1.7e-07 $l=4.85747e-07 $layer=licon1_NDIFF $count=1 $X=3.06
+ $Y=0.37 $X2=3.45 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_2%SET_B 3 7 11 15 19 20 21 22 25 27 30 31 33
c123 31 0 1.62395e-19 $X=8.565 $Y=1.645
c124 3 0 1.66427e-19 $X=5.49 $Y=2.49
r125 33 36 40.8147 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=5.577 $Y=1.955
+ $X2=5.577 $Y2=2.12
r126 33 35 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=5.577 $Y=1.955
+ $X2=5.577 $Y2=1.79
r127 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.59
+ $Y=1.955 $X2=5.59 $Y2=1.955
r128 31 44 10.8302 $w=4.13e-07 $l=3.9e-07 $layer=LI1_cond $X=8.522 $Y=1.645
+ $X2=8.522 $Y2=2.035
r129 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.565
+ $Y=1.645 $X2=8.565 $Y2=1.645
r130 27 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=2.035
+ $X2=8.4 $Y2=2.035
r131 25 34 13.125 $w=3.58e-07 $l=4.1e-07 $layer=LI1_cond $X=6 $Y=1.97 $X2=5.59
+ $Y2=1.97
r132 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=2.035 $X2=6
+ $Y2=2.035
r133 22 24 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.145 $Y=2.035
+ $X2=6 $Y2=2.035
r134 21 27 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.255 $Y=2.035
+ $X2=8.4 $Y2=2.035
r135 21 22 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=8.255 $Y=2.035
+ $X2=6.145 $Y2=2.035
r136 19 30 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.565 $Y=1.985
+ $X2=8.565 $Y2=1.645
r137 19 20 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.565 $Y=1.985
+ $X2=8.565 $Y2=2.15
r138 18 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.565 $Y=1.48
+ $X2=8.565 $Y2=1.645
r139 15 20 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=8.49 $Y=2.75 $X2=8.49
+ $Y2=2.15
r140 11 18 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=8.475 $Y=0.8
+ $X2=8.475 $Y2=1.48
r141 7 35 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=5.6 $Y=0.8 $X2=5.6
+ $Y2=1.79
r142 3 36 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=5.49 $Y=2.49
+ $X2=5.49 $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_2%A_225_74# 1 2 9 13 16 18 19 20 21 22 25 29
+ 31 36 37 38 41 44 45 46 47 49 50 51 54 58 62 65
c186 54 0 2.99812e-20 $X=1.945 $Y=1.805
c187 29 0 1.38641e-19 $X=3.505 $Y=2.49
r188 62 64 17.9907 $w=4.58e-07 $l=5e-07 $layer=LI1_cond $X=1.205 $Y=0.51
+ $X2=1.205 $Y2=1.01
r189 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.11
+ $Y=1.465 $X2=2.11 $Y2=1.465
r190 56 58 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.11 $Y=1.72
+ $X2=2.11 $Y2=1.465
r191 54 56 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.945 $Y=1.805
+ $X2=2.11 $Y2=1.72
r192 54 65 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.945 $Y=1.805
+ $X2=1.455 $Y2=1.805
r193 51 53 5.57014 $w=2.98e-07 $l=1.45e-07 $layer=LI1_cond $X=1.145 $Y=1.87
+ $X2=1.29 $Y2=1.87
r194 50 65 7.90841 $w=2.98e-07 $l=1.5e-07 $layer=LI1_cond $X=1.305 $Y=1.87
+ $X2=1.455 $Y2=1.87
r195 50 53 0.576222 $w=2.98e-07 $l=1.5e-08 $layer=LI1_cond $X=1.305 $Y=1.87
+ $X2=1.29 $Y2=1.87
r196 49 51 7.51767 $w=3e-07 $l=1.8775e-07 $layer=LI1_cond $X=1.06 $Y=1.72
+ $X2=1.145 $Y2=1.87
r197 49 64 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.06 $Y=1.72
+ $X2=1.06 $Y2=1.01
r198 45 59 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=2.41 $Y=1.465
+ $X2=2.11 $Y2=1.465
r199 45 46 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.41 $Y=1.465
+ $X2=2.485 $Y2=1.465
r200 43 59 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=2.055 $Y=1.465
+ $X2=2.11 $Y2=1.465
r201 43 44 3.90195 $w=3.3e-07 $l=1.08e-07 $layer=POLY_cond $X=2.055 $Y=1.465
+ $X2=1.947 $Y2=1.465
r202 39 41 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.37 $Y=1.66
+ $X2=7.37 $Y2=0.8
r203 37 39 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.295 $Y=1.735
+ $X2=7.37 $Y2=1.66
r204 37 38 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=7.295 $Y=1.735
+ $X2=6.85 $Y2=1.735
r205 34 36 239.056 $w=1.8e-07 $l=6.15e-07 $layer=POLY_cond $X=6.76 $Y=3.075
+ $X2=6.76 $Y2=2.46
r206 33 38 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.76 $Y=1.81
+ $X2=6.85 $Y2=1.735
r207 33 36 252.661 $w=1.8e-07 $l=6.5e-07 $layer=POLY_cond $X=6.76 $Y=1.81
+ $X2=6.76 $Y2=2.46
r208 32 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.595 $Y=3.15
+ $X2=3.505 $Y2=3.15
r209 31 34 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.67 $Y=3.15
+ $X2=6.76 $Y2=3.075
r210 31 32 1576.76 $w=1.5e-07 $l=3.075e-06 $layer=POLY_cond $X=6.67 $Y=3.15
+ $X2=3.595 $Y2=3.15
r211 27 47 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.505 $Y=3.075
+ $X2=3.505 $Y2=3.15
r212 27 29 227.395 $w=1.8e-07 $l=5.85e-07 $layer=POLY_cond $X=3.505 $Y=3.075
+ $X2=3.505 $Y2=2.49
r213 23 25 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.985 $Y=0.99
+ $X2=2.985 $Y2=0.58
r214 21 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.415 $Y=3.15
+ $X2=3.505 $Y2=3.15
r215 21 22 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=3.415 $Y=3.15
+ $X2=2.56 $Y2=3.15
r216 19 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.91 $Y=1.065
+ $X2=2.985 $Y2=0.99
r217 19 20 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=2.91 $Y=1.065
+ $X2=2.56 $Y2=1.065
r218 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.485 $Y=3.075
+ $X2=2.56 $Y2=3.15
r219 17 46 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.485 $Y=1.63
+ $X2=2.485 $Y2=1.465
r220 17 18 740.947 $w=1.5e-07 $l=1.445e-06 $layer=POLY_cond $X=2.485 $Y=1.63
+ $X2=2.485 $Y2=3.075
r221 16 46 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.485 $Y=1.3
+ $X2=2.485 $Y2=1.465
r222 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.485 $Y=1.14
+ $X2=2.56 $Y2=1.065
r223 15 16 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.485 $Y=1.14
+ $X2=2.485 $Y2=1.3
r224 11 44 34.7346 $w=1.65e-07 $l=1.73767e-07 $layer=POLY_cond $X=1.965 $Y=1.63
+ $X2=1.947 $Y2=1.465
r225 11 13 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.965 $Y=1.63
+ $X2=1.965 $Y2=2.35
r226 7 44 34.7346 $w=1.65e-07 $l=1.80291e-07 $layer=POLY_cond $X=1.915 $Y=1.3
+ $X2=1.947 $Y2=1.465
r227 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.915 $Y=1.3
+ $X2=1.915 $Y2=0.74
r228 2 53 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=1.79 $X2=1.29 $Y2=1.935
r229 1 62 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.125
+ $Y=0.37 $X2=1.27 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_2%A_1566_92# 1 2 9 12 15 18 19 22 24 25 28 32
+ 34 38
c78 18 0 1.23601e-19 $X=7.995 $Y=1.285
c79 12 0 1.62395e-19 $X=7.95 $Y=2.75
r80 30 34 3.10218 $w=3.05e-07 $l=1.09087e-07 $layer=LI1_cond $X=9.765 $Y=1.24
+ $X2=9.71 $Y2=1.155
r81 30 32 69.6076 $w=2.48e-07 $l=1.51e-06 $layer=LI1_cond $X=9.765 $Y=1.24
+ $X2=9.765 $Y2=2.75
r82 26 34 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=9.71 $Y=1.07
+ $X2=9.71 $Y2=1.155
r83 26 28 8.64332 $w=3.58e-07 $l=2.7e-07 $layer=LI1_cond $X=9.71 $Y=1.07
+ $X2=9.71 $Y2=0.8
r84 24 34 3.51065 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=9.53 $Y=1.155
+ $X2=9.71 $Y2=1.155
r85 24 25 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=9.53 $Y=1.155
+ $X2=8.145 $Y2=1.155
r86 22 38 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.995 $Y=1.965
+ $X2=7.995 $Y2=2.13
r87 21 22 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.995
+ $Y=1.965 $X2=7.995 $Y2=1.965
r88 19 22 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=7.995 $Y=1.285
+ $X2=7.995 $Y2=1.965
r89 18 21 24.8781 $w=3.13e-07 $l=6.8e-07 $layer=LI1_cond $X=7.987 $Y=1.285
+ $X2=7.987 $Y2=1.965
r90 18 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.995
+ $Y=1.285 $X2=7.995 $Y2=1.285
r91 16 25 7.64049 $w=1.7e-07 $l=1.95944e-07 $layer=LI1_cond $X=7.987 $Y=1.24
+ $X2=8.145 $Y2=1.155
r92 16 18 1.64635 $w=3.13e-07 $l=4.5e-08 $layer=LI1_cond $X=7.987 $Y=1.24
+ $X2=7.987 $Y2=1.285
r93 15 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.995 $Y=1.12
+ $X2=7.995 $Y2=1.285
r94 12 38 241 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=7.95 $Y=2.75 $X2=7.95
+ $Y2=2.13
r95 9 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.905 $Y=0.8
+ $X2=7.905 $Y2=1.12
r96 2 32 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=9.59
+ $Y=2.54 $X2=9.725 $Y2=2.75
r97 1 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.555
+ $Y=0.59 $X2=9.695 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_2%A_1356_74# 1 2 3 12 16 18 22 24 26 28 30 31
+ 35 37 38 40 41 44 46 50 51 55 61 65 71
c154 55 0 3.20959e-20 $X=7.235 $Y=1.705
c155 41 0 1.76198e-19 $X=7.93 $Y=2.435
c156 31 0 8.20619e-20 $X=10.497 $Y=1.69
r157 63 65 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=7.035 $Y=0.785
+ $X2=7.235 $Y2=0.785
r158 60 61 8.41349 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.305 $Y=2.765
+ $X2=7.47 $Y2=2.765
r159 57 60 9.64836 $w=4.28e-07 $l=3.6e-07 $layer=LI1_cond $X=6.945 $Y=2.765
+ $X2=7.305 $Y2=2.765
r160 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.305
+ $Y=1.78 $X2=9.305 $Y2=1.78
r161 48 50 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=9.305 $Y=2.32
+ $X2=9.305 $Y2=1.78
r162 47 71 6.19399 $w=2e-07 $l=1.39194e-07 $layer=LI1_cond $X=8.88 $Y=2.405
+ $X2=8.755 $Y2=2.435
r163 46 48 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.14 $Y=2.405
+ $X2=9.305 $Y2=2.32
r164 46 47 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=9.14 $Y=2.405
+ $X2=8.88 $Y2=2.405
r165 42 71 0.552779 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=8.755 $Y=2.55
+ $X2=8.755 $Y2=2.435
r166 42 44 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=8.755 $Y=2.55
+ $X2=8.755 $Y2=2.75
r167 41 69 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=7.845 $Y=2.435
+ $X2=7.845 $Y2=2.64
r168 40 71 6.19399 $w=2e-07 $l=1.25e-07 $layer=LI1_cond $X=8.63 $Y=2.435
+ $X2=8.755 $Y2=2.435
r169 40 41 35.0744 $w=2.28e-07 $l=7e-07 $layer=LI1_cond $X=8.63 $Y=2.435
+ $X2=7.93 $Y2=2.435
r170 38 69 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.76 $Y=2.64
+ $X2=7.845 $Y2=2.64
r171 38 61 17.8687 $w=1.78e-07 $l=2.9e-07 $layer=LI1_cond $X=7.76 $Y=2.64
+ $X2=7.47 $Y2=2.64
r172 37 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.235 $Y=1.62
+ $X2=7.235 $Y2=1.705
r173 36 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.235 $Y=0.95
+ $X2=7.235 $Y2=0.785
r174 36 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.235 $Y=0.95
+ $X2=7.235 $Y2=1.62
r175 33 57 3.91032 $w=2.5e-07 $l=2.15e-07 $layer=LI1_cond $X=6.945 $Y=2.55
+ $X2=6.945 $Y2=2.765
r176 33 35 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=6.945 $Y=2.55
+ $X2=6.945 $Y2=2.14
r177 32 55 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.945 $Y=1.705
+ $X2=7.235 $Y2=1.705
r178 32 35 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=6.945 $Y=1.79
+ $X2=6.945 $Y2=2.14
r179 29 51 34.6051 $w=4.5e-07 $l=2.8e-07 $layer=POLY_cond $X=9.365 $Y=2.06
+ $X2=9.365 $Y2=1.78
r180 29 30 48.4927 $w=4.5e-07 $l=2.25e-07 $layer=POLY_cond $X=9.365 $Y=2.06
+ $X2=9.365 $Y2=2.285
r181 27 51 1.85385 $w=4.5e-07 $l=1.5e-08 $layer=POLY_cond $X=9.365 $Y=1.765
+ $X2=9.365 $Y2=1.78
r182 27 28 11.1008 $w=3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.365 $Y=1.765
+ $X2=9.365 $Y2=1.69
r183 24 31 18.8402 $w=1.65e-07 $l=8.12404e-08 $layer=POLY_cond $X=10.51 $Y=1.765
+ $X2=10.497 $Y2=1.69
r184 24 26 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.51 $Y=1.765
+ $X2=10.51 $Y2=2.34
r185 20 31 18.8402 $w=1.65e-07 $l=8.74643e-08 $layer=POLY_cond $X=10.47 $Y=1.615
+ $X2=10.497 $Y2=1.69
r186 20 22 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=10.47 $Y=1.615
+ $X2=10.47 $Y2=0.79
r187 19 28 15.4994 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=9.59 $Y=1.69
+ $X2=9.365 $Y2=1.69
r188 18 31 6.66866 $w=1.5e-07 $l=1.02e-07 $layer=POLY_cond $X=10.395 $Y=1.69
+ $X2=10.497 $Y2=1.69
r189 18 19 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=10.395 $Y=1.69
+ $X2=9.59 $Y2=1.69
r190 16 30 180.75 $w=1.8e-07 $l=4.65e-07 $layer=POLY_cond $X=9.5 $Y=2.75 $X2=9.5
+ $Y2=2.285
r191 10 28 11.1008 $w=3e-07 $l=1.47817e-07 $layer=POLY_cond $X=9.48 $Y=1.615
+ $X2=9.365 $Y2=1.69
r192 10 12 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=9.48 $Y=1.615
+ $X2=9.48 $Y2=0.8
r193 3 44 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=8.58
+ $Y=2.54 $X2=8.715 $Y2=2.75
r194 2 60 600 $w=1.7e-07 $l=1.05832e-06 $layer=licon1_PDIFF $count=1 $X=6.85
+ $Y=1.96 $X2=7.305 $Y2=2.815
r195 2 35 300 $w=1.7e-07 $l=2.38118e-07 $layer=licon1_PDIFF $count=2 $X=6.85
+ $Y=1.96 $X2=6.985 $Y2=2.14
r196 1 63 182 $w=1.7e-07 $l=5.27304e-07 $layer=licon1_NDIFF $count=1 $X=6.78
+ $Y=0.37 $X2=7.035 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_2%A_2022_94# 1 2 9 13 17 21 25 29 35 38 44
c70 38 0 7.76856e-20 $X=10.27 $Y=1.465
r71 43 44 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=11.48 $Y=1.465
+ $X2=11.495 $Y2=1.465
r72 42 43 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=11.05 $Y=1.465
+ $X2=11.48 $Y2=1.465
r73 41 42 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=11.045 $Y=1.465
+ $X2=11.05 $Y2=1.465
r74 36 41 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=10.975 $Y=1.465
+ $X2=11.045 $Y2=1.465
r75 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.975
+ $Y=1.465 $X2=10.975 $Y2=1.465
r76 33 38 1.50311 $w=3.3e-07 $l=1.8e-07 $layer=LI1_cond $X=10.45 $Y=1.465
+ $X2=10.27 $Y2=1.465
r77 33 35 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=10.45 $Y=1.465
+ $X2=10.975 $Y2=1.465
r78 29 31 22.7287 $w=3.58e-07 $l=7.1e-07 $layer=LI1_cond $X=10.27 $Y=1.985
+ $X2=10.27 $Y2=2.695
r79 27 38 4.97762 $w=3.45e-07 $l=1.65e-07 $layer=LI1_cond $X=10.27 $Y=1.63
+ $X2=10.27 $Y2=1.465
r80 27 29 11.3644 $w=3.58e-07 $l=3.55e-07 $layer=LI1_cond $X=10.27 $Y=1.63
+ $X2=10.27 $Y2=1.985
r81 23 38 4.97762 $w=3.45e-07 $l=1.72337e-07 $layer=LI1_cond $X=10.255 $Y=1.3
+ $X2=10.27 $Y2=1.465
r82 23 25 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=10.255 $Y=1.3
+ $X2=10.255 $Y2=0.615
r83 19 44 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=11.495 $Y=1.63
+ $X2=11.495 $Y2=1.465
r84 19 21 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=11.495 $Y=1.63
+ $X2=11.495 $Y2=2.4
r85 15 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.48 $Y=1.3
+ $X2=11.48 $Y2=1.465
r86 15 17 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.48 $Y=1.3
+ $X2=11.48 $Y2=0.74
r87 11 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.05 $Y=1.3
+ $X2=11.05 $Y2=1.465
r88 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.05 $Y=1.3
+ $X2=11.05 $Y2=0.74
r89 7 41 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=11.045 $Y=1.63
+ $X2=11.045 $Y2=1.465
r90 7 9 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=11.045 $Y=1.63
+ $X2=11.045 $Y2=2.4
r91 2 31 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=10.14
+ $Y=1.84 $X2=10.285 $Y2=2.695
r92 2 29 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.14
+ $Y=1.84 $X2=10.285 $Y2=1.985
r93 1 25 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=10.11
+ $Y=0.47 $X2=10.255 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_2%A_27_74# 1 2 3 4 14 17 19 21 24 26 29 30 37
c70 24 0 8.11169e-20 $X=2.53 $Y=2.06
c71 21 0 1.38641e-19 $X=2.445 $Y=2.145
r72 34 37 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.53 $Y=0.76 $X2=2.69
+ $Y2=0.76
r73 30 32 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.71 $Y=2.145
+ $X2=1.71 $Y2=2.275
r74 26 28 9.71523 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=0.24 $Y=0.58
+ $X2=0.24 $Y2=0.765
r75 23 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.53 $Y=0.925
+ $X2=2.53 $Y2=0.76
r76 23 24 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=2.53 $Y=0.925
+ $X2=2.53 $Y2=2.06
r77 22 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.795 $Y=2.145
+ $X2=1.71 $Y2=2.145
r78 21 41 10.5225 $w=4e-07 $l=4.53073e-07 $layer=LI1_cond $X=2.445 $Y=2.145
+ $X2=2.695 $Y2=2.49
r79 21 24 6.71454 $w=4e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.445 $Y=2.145
+ $X2=2.53 $Y2=2.06
r80 21 22 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.445 $Y=2.145
+ $X2=1.795 $Y2=2.145
r81 20 29 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=2.275
+ $X2=0.24 $Y2=2.275
r82 19 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=2.275
+ $X2=1.71 $Y2=2.275
r83 19 20 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=1.625 $Y=2.275
+ $X2=0.365 $Y2=2.275
r84 15 29 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.36 $X2=0.24
+ $Y2=2.275
r85 15 17 17.9781 $w=2.48e-07 $l=3.9e-07 $layer=LI1_cond $X=0.24 $Y=2.36
+ $X2=0.24 $Y2=2.75
r86 14 29 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.2 $Y=2.19
+ $X2=0.24 $Y2=2.275
r87 14 28 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=0.2 $Y=2.19
+ $X2=0.2 $Y2=0.765
r88 4 41 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=2.635
+ $Y=2.28 $X2=2.78 $Y2=2.49
r89 3 17 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.28 $Y2=2.75
r90 2 37 182 $w=1.7e-07 $l=4.56782e-07 $layer=licon1_NDIFF $count=1 $X=2.545
+ $Y=0.37 $X2=2.69 $Y2=0.76
r91 1 26 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_2%VPWR 1 2 3 4 5 6 7 8 27 31 34 37 41 45 49 53
+ 55 62 65 66 67 69 74 79 84 99 103 108 114 117 120 123 126 129 133
c147 31 0 2.99812e-20 $X=1.74 $Y=2.73
r148 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r149 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r150 126 127 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r151 120 121 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r152 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r153 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r154 112 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r155 112 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r156 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r157 109 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.985 $Y=3.33
+ $X2=10.82 $Y2=3.33
r158 109 111 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.985 $Y=3.33
+ $X2=11.28 $Y2=3.33
r159 108 132 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=11.635 $Y=3.33
+ $X2=11.817 $Y2=3.33
r160 108 111 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=11.635 $Y=3.33
+ $X2=11.28 $Y2=3.33
r161 107 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r162 107 127 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.36 $Y2=3.33
r163 106 107 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r164 104 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.44 $Y=3.33
+ $X2=9.275 $Y2=3.33
r165 104 106 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=9.44 $Y=3.33
+ $X2=10.32 $Y2=3.33
r166 103 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.655 $Y=3.33
+ $X2=10.82 $Y2=3.33
r167 103 106 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=10.655 $Y=3.33
+ $X2=10.32 $Y2=3.33
r168 102 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r169 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r170 99 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.11 $Y=3.33
+ $X2=9.275 $Y2=3.33
r171 99 101 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=9.11 $Y=3.33
+ $X2=8.88 $Y2=3.33
r172 98 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r173 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r174 95 98 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.92 $Y2=3.33
r175 94 97 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=7.92 $Y2=3.33
r176 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r177 92 123 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.11 $Y=3.33
+ $X2=5.985 $Y2=3.33
r178 92 94 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.11 $Y=3.33
+ $X2=6.48 $Y2=3.33
r179 90 91 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r180 88 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r181 88 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r182 87 90 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r183 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r184 85 120 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.24 $Y=3.33
+ $X2=4.155 $Y2=3.33
r185 85 87 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.24 $Y=3.33
+ $X2=4.56 $Y2=3.33
r186 84 123 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.86 $Y=3.33
+ $X2=5.985 $Y2=3.33
r187 84 90 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.86 $Y=3.33
+ $X2=5.52 $Y2=3.33
r188 83 121 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.08 $Y2=3.33
r189 83 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r190 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r191 80 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=1.74 $Y2=3.33
r192 80 82 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.905 $Y=3.33
+ $X2=2.16 $Y2=3.33
r193 79 120 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.07 $Y=3.33
+ $X2=4.155 $Y2=3.33
r194 79 82 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=4.07 $Y=3.33
+ $X2=2.16 $Y2=3.33
r195 78 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r196 78 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r197 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r198 75 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r199 75 77 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r200 74 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.74 $Y2=3.33
r201 74 77 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.2 $Y2=3.33
r202 72 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r203 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r204 69 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r205 69 71 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r206 67 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r207 67 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r208 67 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r209 65 97 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.1 $Y=3.33
+ $X2=7.92 $Y2=3.33
r210 65 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.1 $Y=3.33
+ $X2=8.265 $Y2=3.33
r211 64 101 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=8.43 $Y=3.33
+ $X2=8.88 $Y2=3.33
r212 64 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.43 $Y=3.33
+ $X2=8.265 $Y2=3.33
r213 59 62 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.155 $Y=2.745
+ $X2=4.32 $Y2=2.745
r214 55 58 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=11.76 $Y=1.985
+ $X2=11.76 $Y2=2.815
r215 53 132 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=11.76 $Y=3.245
+ $X2=11.817 $Y2=3.33
r216 53 58 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.76 $Y=3.245
+ $X2=11.76 $Y2=2.815
r217 49 52 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=10.82 $Y=2.405
+ $X2=10.82 $Y2=2.815
r218 47 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.82 $Y=3.245
+ $X2=10.82 $Y2=3.33
r219 47 52 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.82 $Y=3.245
+ $X2=10.82 $Y2=2.815
r220 43 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.275 $Y=3.245
+ $X2=9.275 $Y2=3.33
r221 43 45 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=9.275 $Y=3.245
+ $X2=9.275 $Y2=2.78
r222 39 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.265 $Y=3.245
+ $X2=8.265 $Y2=3.33
r223 39 41 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=8.265 $Y=3.245
+ $X2=8.265 $Y2=2.81
r224 35 123 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.985 $Y=3.245
+ $X2=5.985 $Y2=3.33
r225 35 37 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=5.985 $Y=3.245
+ $X2=5.985 $Y2=2.825
r226 34 120 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.155 $Y=3.245
+ $X2=4.155 $Y2=3.33
r227 33 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.155 $Y=2.91
+ $X2=4.155 $Y2=2.745
r228 33 34 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.155 $Y=2.91
+ $X2=4.155 $Y2=3.245
r229 29 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=3.245
+ $X2=1.74 $Y2=3.33
r230 29 31 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=1.74 $Y=3.245
+ $X2=1.74 $Y2=2.73
r231 25 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r232 25 27 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.755
r233 8 58 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=11.585
+ $Y=1.84 $X2=11.72 $Y2=2.815
r234 8 55 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=11.585
+ $Y=1.84 $X2=11.72 $Y2=1.985
r235 7 52 600 $w=1.7e-07 $l=1.07941e-06 $layer=licon1_PDIFF $count=1 $X=10.6
+ $Y=1.84 $X2=10.82 $Y2=2.815
r236 7 49 600 $w=1.7e-07 $l=6.65977e-07 $layer=licon1_PDIFF $count=1 $X=10.6
+ $Y=1.84 $X2=10.82 $Y2=2.405
r237 6 45 600 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_PDIFF $count=1 $X=9.13
+ $Y=2.54 $X2=9.275 $Y2=2.78
r238 5 41 600 $w=1.7e-07 $l=3.65582e-07 $layer=licon1_PDIFF $count=1 $X=8.04
+ $Y=2.54 $X2=8.265 $Y2=2.81
r239 4 37 600 $w=1.7e-07 $l=7.04237e-07 $layer=licon1_PDIFF $count=1 $X=5.58
+ $Y=2.28 $X2=5.945 $Y2=2.825
r240 3 62 600 $w=1.7e-07 $l=5.98373e-07 $layer=licon1_PDIFF $count=1 $X=4.015
+ $Y=2.28 $X2=4.32 $Y2=2.745
r241 2 31 600 $w=1.7e-07 $l=1.00524e-06 $layer=licon1_PDIFF $count=1 $X=1.605
+ $Y=1.79 $X2=1.74 $Y2=2.73
r242 1 27 600 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=2.54 $X2=0.73 $Y2=2.755
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_2%Q 1 2 9 13 16 17 18 19 22
c39 16 0 4.37624e-21 $X=11.38 $Y=1.82
r40 19 22 0.225187 $w=3.3e-07 $l=1.55e-07 $layer=LI1_cond $X=11.31 $Y=1.985
+ $X2=11.155 $Y2=1.985
r41 18 22 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=10.8 $Y=1.985
+ $X2=11.155 $Y2=1.985
r42 16 19 6.67463 $w=2.4e-07 $l=1.96914e-07 $layer=LI1_cond $X=11.38 $Y=1.82
+ $X2=11.31 $Y2=1.985
r43 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=11.38 $Y=1.82
+ $X2=11.38 $Y2=1.13
r44 11 19 6.67463 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=11.31 $Y=2.15
+ $X2=11.31 $Y2=1.985
r45 11 13 9.29389 $w=3.08e-07 $l=2.5e-07 $layer=LI1_cond $X=11.31 $Y=2.15
+ $X2=11.31 $Y2=2.4
r46 7 17 9.06106 $w=3.63e-07 $l=1.82e-07 $layer=LI1_cond $X=11.282 $Y=0.948
+ $X2=11.282 $Y2=1.13
r47 7 9 13.6714 $w=3.63e-07 $l=4.33e-07 $layer=LI1_cond $X=11.282 $Y=0.948
+ $X2=11.282 $Y2=0.515
r48 2 19 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=11.135
+ $Y=1.84 $X2=11.27 $Y2=1.985
r49 2 13 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=11.135
+ $Y=1.84 $X2=11.27 $Y2=2.4
r50 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.125
+ $Y=0.37 $X2=11.265 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DFSTP_2%VGND 1 2 3 4 5 6 7 24 26 30 34 38 42 46 48
+ 50 52 57 65 70 78 86 92 95 98 101 111 115
c110 30 0 9.68091e-20 $X=1.7 $Y=0.495
r111 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r112 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r113 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r114 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r115 93 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r116 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r117 90 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r118 90 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r119 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r120 87 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.93 $Y=0
+ $X2=10.765 $Y2=0
r121 87 89 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=10.93 $Y=0
+ $X2=11.28 $Y2=0
r122 86 114 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=11.635 $Y=0
+ $X2=11.817 $Y2=0
r123 86 89 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=11.635 $Y=0
+ $X2=11.28 $Y2=0
r124 85 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r125 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r126 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=10.32 $Y2=0
r127 82 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r128 81 84 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=9.36 $Y=0 $X2=10.32
+ $Y2=0
r129 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r130 78 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.6 $Y=0
+ $X2=10.765 $Y2=0
r131 78 84 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.6 $Y=0 $X2=10.32
+ $Y2=0
r132 77 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r133 76 77 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r134 74 77 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r135 73 76 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r136 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r137 71 101 12.4999 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=6.245 $Y=0
+ $X2=5.947 $Y2=0
r138 71 73 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.245 $Y=0
+ $X2=6.48 $Y2=0
r139 70 108 10.5284 $w=8.33e-07 $l=7.35e-07 $layer=LI1_cond $X=8.942 $Y=0
+ $X2=8.942 $Y2=0.735
r140 70 81 10.4966 $w=1.7e-07 $l=4.18e-07 $layer=LI1_cond $X=8.942 $Y=0 $X2=9.36
+ $Y2=0
r141 70 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r142 70 76 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=8.525 $Y=0 $X2=8.4
+ $Y2=0
r143 69 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r144 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r145 66 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.6 $Y=0 $X2=4.435
+ $Y2=0
r146 66 68 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.6 $Y=0 $X2=5.52
+ $Y2=0
r147 65 101 12.4999 $w=1.7e-07 $l=2.97e-07 $layer=LI1_cond $X=5.65 $Y=0
+ $X2=5.947 $Y2=0
r148 65 68 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=5.65 $Y=0 $X2=5.52
+ $Y2=0
r149 64 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r150 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r151 61 64 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=4.08 $Y2=0
r152 61 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r153 60 63 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r154 60 61 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r155 58 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.74
+ $Y2=0
r156 58 60 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.16
+ $Y2=0
r157 57 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.27 $Y=0 $X2=4.435
+ $Y2=0
r158 57 63 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.27 $Y=0 $X2=4.08
+ $Y2=0
r159 55 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r160 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r161 52 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.67
+ $Y2=0
r162 52 54 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0
+ $X2=0.24 $Y2=0
r163 50 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r164 50 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r165 50 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r166 46 114 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=11.76 $Y=0.085
+ $X2=11.817 $Y2=0
r167 46 48 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=11.76 $Y=0.085
+ $X2=11.76 $Y2=0.515
r168 42 44 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=10.765 $Y=0.515
+ $X2=10.765 $Y2=0.965
r169 40 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.765 $Y=0.085
+ $X2=10.765 $Y2=0
r170 40 42 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.765 $Y=0.085
+ $X2=10.765 $Y2=0.515
r171 36 101 2.50116 $w=5.95e-07 $l=8.5e-08 $layer=LI1_cond $X=5.947 $Y=0.085
+ $X2=5.947 $Y2=0
r172 36 38 8.64393 $w=5.93e-07 $l=4.3e-07 $layer=LI1_cond $X=5.947 $Y=0.085
+ $X2=5.947 $Y2=0.515
r173 32 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.435 $Y=0.085
+ $X2=4.435 $Y2=0
r174 32 34 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=4.435 $Y=0.085
+ $X2=4.435 $Y2=0.53
r175 28 95 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=0.085
+ $X2=1.74 $Y2=0
r176 28 30 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=1.74 $Y=0.085
+ $X2=1.74 $Y2=0.495
r177 27 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.67
+ $Y2=0
r178 26 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.615 $Y=0 $X2=1.74
+ $Y2=0
r179 26 27 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=1.615 $Y=0
+ $X2=0.795 $Y2=0
r180 22 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0
r181 22 24 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.67 $Y=0.085
+ $X2=0.67 $Y2=0.58
r182 7 48 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=11.555
+ $Y=0.37 $X2=11.72 $Y2=0.515
r183 6 44 182 $w=1.7e-07 $l=5.94916e-07 $layer=licon1_NDIFF $count=1 $X=10.545
+ $Y=0.47 $X2=10.765 $Y2=0.965
r184 6 42 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=10.545
+ $Y=0.47 $X2=10.765 $Y2=0.515
r185 5 108 91 $w=1.7e-07 $l=7.13828e-07 $layer=licon1_NDIFF $count=2 $X=8.55
+ $Y=0.59 $X2=9.195 $Y2=0.735
r186 4 38 91 $w=1.7e-07 $l=4.40908e-07 $layer=licon1_NDIFF $count=2 $X=5.675
+ $Y=0.59 $X2=6.08 $Y2=0.515
r187 3 34 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=4.295
+ $Y=0.37 $X2=4.435 $Y2=0.53
r188 2 30 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.56
+ $Y=0.37 $X2=1.7 $Y2=0.495
r189 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.58
.ends


* File: sky130_fd_sc_ms__nor2_1.pxi.spice
* Created: Wed Sep  2 12:15:11 2020
* 
x_PM_SKY130_FD_SC_MS__NOR2_1%A N_A_M1000_g N_A_M1003_g A N_A_c_31_n N_A_c_32_n
+ PM_SKY130_FD_SC_MS__NOR2_1%A
x_PM_SKY130_FD_SC_MS__NOR2_1%B N_B_M1001_g N_B_M1002_g B N_B_c_58_n N_B_c_59_n
+ PM_SKY130_FD_SC_MS__NOR2_1%B
x_PM_SKY130_FD_SC_MS__NOR2_1%VPWR N_VPWR_M1000_s N_VPWR_c_80_n N_VPWR_c_81_n
+ VPWR N_VPWR_c_82_n N_VPWR_c_79_n PM_SKY130_FD_SC_MS__NOR2_1%VPWR
x_PM_SKY130_FD_SC_MS__NOR2_1%Y N_Y_M1003_d N_Y_M1001_d N_Y_c_97_n N_Y_c_98_n
+ N_Y_c_99_n Y Y PM_SKY130_FD_SC_MS__NOR2_1%Y
x_PM_SKY130_FD_SC_MS__NOR2_1%VGND N_VGND_M1003_s N_VGND_M1002_d N_VGND_c_123_n
+ N_VGND_c_124_n N_VGND_c_125_n N_VGND_c_126_n VGND N_VGND_c_127_n
+ N_VGND_c_128_n PM_SKY130_FD_SC_MS__NOR2_1%VGND
cc_1 VNB N_A_M1000_g 0.00188957f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A_M1003_g 0.0271489f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_3 VNB N_A_c_31_n 0.00600492f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_4 VNB N_A_c_32_n 0.0572007f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.465
cc_5 VNB N_B_M1001_g 0.00188938f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_6 VNB N_B_M1002_g 0.028217f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_7 VNB N_B_c_58_n 0.0591087f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_8 VNB N_B_c_59_n 0.00385705f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.465
cc_9 VNB N_VPWR_c_79_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.465
cc_10 VNB N_Y_c_97_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_11 VNB N_Y_c_98_n 0.00960735f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_12 VNB N_Y_c_99_n 0.0022354f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_13 VNB N_VGND_c_123_n 0.011316f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.74
cc_14 VNB N_VGND_c_124_n 0.0411496f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_15 VNB N_VGND_c_125_n 0.0120272f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_16 VNB N_VGND_c_126_n 0.0404679f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.465
cc_17 VNB N_VGND_c_127_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_128_n 0.115949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VPB N_A_M1000_g 0.0272633f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_20 VPB N_A_c_31_n 0.00716464f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_21 VPB N_B_M1001_g 0.0295056f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_22 VPB N_B_c_59_n 0.0072578f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=1.465
cc_23 VPB N_VPWR_c_80_n 0.0119967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_24 VPB N_VPWR_c_81_n 0.0487556f $X=-0.19 $Y=1.66 $X2=0.515 $Y2=0.74
cc_25 VPB N_VPWR_c_82_n 0.0288332f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_26 VPB N_VPWR_c_79_n 0.0512627f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_27 VPB N_Y_c_98_n 0.00315112f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.465
cc_28 VPB Y 0.0450983f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.465
cc_29 N_A_M1000_g N_B_M1001_g 0.0442427f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_30 N_A_M1003_g N_B_M1002_g 0.0144801f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_31 N_A_c_32_n N_B_c_58_n 0.0442427f $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_32 N_A_M1000_g N_VPWR_c_81_n 0.0184219f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_33 N_A_c_31_n N_VPWR_c_81_n 0.0256722f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_34 N_A_c_32_n N_VPWR_c_81_n 0.00146577f $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_35 N_A_M1000_g N_VPWR_c_82_n 0.00460063f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_36 N_A_M1000_g N_VPWR_c_79_n 0.00908371f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_37 N_A_M1003_g N_Y_c_97_n 0.00809519f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_38 N_A_M1003_g N_Y_c_98_n 0.00403324f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_39 N_A_c_31_n N_Y_c_98_n 0.0331382f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_40 N_A_c_32_n N_Y_c_98_n 0.00547875f $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_41 N_A_M1003_g N_Y_c_99_n 0.00278377f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_42 N_A_c_32_n N_Y_c_99_n 2.41927e-19 $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_43 N_A_M1000_g Y 2.55565e-19 $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_44 N_A_M1003_g N_VGND_c_124_n 0.00511162f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_45 N_A_c_31_n N_VGND_c_124_n 0.0215684f $X=0.29 $Y=1.465 $X2=0 $Y2=0
cc_46 N_A_c_32_n N_VGND_c_124_n 0.00196285f $X=0.515 $Y=1.465 $X2=0 $Y2=0
cc_47 N_A_M1003_g N_VGND_c_126_n 6.14817e-19 $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_48 N_A_M1003_g N_VGND_c_127_n 0.00434272f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_49 N_A_M1003_g N_VGND_c_128_n 0.00824106f $X=0.515 $Y=0.74 $X2=0 $Y2=0
cc_50 N_B_M1001_g N_VPWR_c_81_n 0.00150327f $X=0.925 $Y=2.4 $X2=0 $Y2=0
cc_51 N_B_M1001_g N_VPWR_c_82_n 0.00361596f $X=0.925 $Y=2.4 $X2=0 $Y2=0
cc_52 N_B_M1001_g N_VPWR_c_79_n 0.0044565f $X=0.925 $Y=2.4 $X2=0 $Y2=0
cc_53 N_B_M1002_g N_Y_c_97_n 0.00457569f $X=0.945 $Y=0.74 $X2=0 $Y2=0
cc_54 N_B_c_58_n N_Y_c_98_n 0.00565646f $X=1.15 $Y=1.465 $X2=0 $Y2=0
cc_55 N_B_c_59_n N_Y_c_98_n 0.0360321f $X=1.15 $Y=1.465 $X2=0 $Y2=0
cc_56 N_B_M1001_g Y 0.0353839f $X=0.925 $Y=2.4 $X2=0 $Y2=0
cc_57 N_B_c_58_n Y 0.00152065f $X=1.15 $Y=1.465 $X2=0 $Y2=0
cc_58 N_B_c_59_n Y 0.0265852f $X=1.15 $Y=1.465 $X2=0 $Y2=0
cc_59 N_B_M1002_g N_VGND_c_126_n 0.0151529f $X=0.945 $Y=0.74 $X2=0 $Y2=0
cc_60 N_B_c_58_n N_VGND_c_126_n 0.00232693f $X=1.15 $Y=1.465 $X2=0 $Y2=0
cc_61 N_B_c_59_n N_VGND_c_126_n 0.0275482f $X=1.15 $Y=1.465 $X2=0 $Y2=0
cc_62 N_B_M1002_g N_VGND_c_127_n 0.00383152f $X=0.945 $Y=0.74 $X2=0 $Y2=0
cc_63 N_B_M1002_g N_VGND_c_128_n 0.00757637f $X=0.945 $Y=0.74 $X2=0 $Y2=0
cc_64 N_VPWR_c_81_n Y 0.00262262f $X=0.28 $Y=2.115 $X2=0 $Y2=0
cc_65 N_VPWR_c_82_n Y 0.0241709f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_66 N_VPWR_c_79_n Y 0.0231171f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_67 A_119_368# Y 0.0019061f $X=0.595 $Y=1.84 $X2=1.115 $Y2=2.69
cc_68 N_Y_c_97_n N_VGND_c_124_n 0.0282134f $X=0.73 $Y=0.515 $X2=0 $Y2=0
cc_69 N_Y_c_97_n N_VGND_c_126_n 0.0294122f $X=0.73 $Y=0.515 $X2=0 $Y2=0
cc_70 N_Y_c_97_n N_VGND_c_127_n 0.0109942f $X=0.73 $Y=0.515 $X2=0 $Y2=0
cc_71 N_Y_c_97_n N_VGND_c_128_n 0.00904371f $X=0.73 $Y=0.515 $X2=0 $Y2=0

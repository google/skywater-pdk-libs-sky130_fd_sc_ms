* File: sky130_fd_sc_ms__xnor3_1.pex.spice
* Created: Wed Sep  2 12:33:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__XNOR3_1%A_81_268# 1 2 9 13 17 18 19 20 21 23 24 25
+ 27 28 29 32 35 36 37 40 45
r102 40 42 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=2.49 $Y=2.795
+ $X2=2.49 $Y2=2.99
r103 36 46 40.7727 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=1.505
+ $X2=0.58 $Y2=1.67
r104 36 45 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=1.505
+ $X2=0.58 $Y2=1.34
r105 35 38 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.605 $Y=1.505
+ $X2=0.605 $Y2=1.67
r106 35 37 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.605 $Y=1.505
+ $X2=0.605 $Y2=1.34
r107 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.505 $X2=0.59 $Y2=1.505
r108 30 32 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.5 $Y=0.425 $X2=2.5
+ $Y2=0.545
r109 28 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.335 $Y=0.34
+ $X2=2.5 $Y2=0.425
r110 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.335 $Y=0.34
+ $X2=1.665 $Y2=0.34
r111 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.58 $Y=0.425
+ $X2=1.665 $Y2=0.34
r112 26 27 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.58 $Y=0.425
+ $X2=1.58 $Y2=0.66
r113 24 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=2.99
+ $X2=2.49 $Y2=2.99
r114 24 25 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=2.325 $Y=2.99
+ $X2=1.145 $Y2=2.99
r115 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.06 $Y=2.905
+ $X2=1.145 $Y2=2.99
r116 22 23 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=1.06 $Y=2.12
+ $X2=1.06 $Y2=2.905
r117 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.975 $Y=2.035
+ $X2=1.06 $Y2=2.12
r118 20 21 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.975 $Y=2.035
+ $X2=0.785 $Y2=2.035
r119 18 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.495 $Y=0.745
+ $X2=1.58 $Y2=0.66
r120 18 19 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.495 $Y=0.745
+ $X2=0.785 $Y2=0.745
r121 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.7 $Y=1.95
+ $X2=0.785 $Y2=2.035
r122 17 38 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.7 $Y=1.95 $X2=0.7
+ $Y2=1.67
r123 14 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.7 $Y=0.83
+ $X2=0.785 $Y2=0.745
r124 14 37 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.7 $Y=0.83 $X2=0.7
+ $Y2=1.34
r125 13 45 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.495 $Y=0.86
+ $X2=0.495 $Y2=1.34
r126 9 46 283.758 $w=1.8e-07 $l=7.3e-07 $layer=POLY_cond $X=0.495 $Y=2.4
+ $X2=0.495 $Y2=1.67
r127 2 40 600 $w=1.7e-07 $l=9.26283e-07 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=1.97 $X2=2.49 $Y2=2.795
r128 1 32 91 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_NDIFF $count=2 $X=2.29
+ $Y=0.37 $X2=2.5 $Y2=0.545
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_1%C 3 6 8 10 12 14 16 18 20 21 24
c81 21 0 1.63453e-19 $X=1.16 $Y=1.35
c82 20 0 3.39391e-20 $X=1.16 $Y=1.425
r83 23 25 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.515
+ $X2=1.16 $Y2=1.68
r84 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.16
+ $Y=1.515 $X2=1.16 $Y2=1.515
r85 20 23 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.16 $Y=1.425 $X2=1.16
+ $Y2=1.515
r86 20 21 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.16 $Y=1.425
+ $X2=1.16 $Y2=1.35
r87 18 24 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.16 $Y=1.665
+ $X2=1.16 $Y2=1.515
r88 14 17 98.2126 $w=1.68e-07 $l=3.51312e-07 $layer=POLY_cond $X=2.215 $Y=1.085
+ $X2=2.192 $Y2=1.425
r89 14 16 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.215 $Y=1.085
+ $X2=2.215 $Y2=0.69
r90 10 17 44.4659 $w=1.8e-07 $l=1.68464e-07 $layer=POLY_cond $X=2.185 $Y=1.59
+ $X2=2.192 $Y2=1.425
r91 10 12 310.968 $w=1.8e-07 $l=8e-07 $layer=POLY_cond $X=2.185 $Y=1.59
+ $X2=2.185 $Y2=2.39
r92 9 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.425
+ $X2=1.16 $Y2=1.425
r93 8 17 5.52526 $w=1.5e-07 $l=9.7e-08 $layer=POLY_cond $X=2.095 $Y=1.425
+ $X2=2.192 $Y2=1.425
r94 8 9 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=2.095 $Y=1.425
+ $X2=1.325 $Y2=1.425
r95 6 25 186.581 $w=1.8e-07 $l=4.8e-07 $layer=POLY_cond $X=1.175 $Y=2.16
+ $X2=1.175 $Y2=1.68
r96 3 21 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.085 $Y=1.02
+ $X2=1.085 $Y2=1.35
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_1%A_232_162# 1 2 9 13 15 19 23 28 29 31 32 33
c89 19 0 3.39391e-20 $X=1.49 $Y=2.125
r90 32 37 40.9207 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.697 $Y=1.645
+ $X2=2.697 $Y2=1.81
r91 32 36 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.697 $Y=1.645
+ $X2=2.697 $Y2=1.48
r92 31 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.68 $Y=1.645
+ $X2=2.515 $Y2=1.645
r93 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.645 $X2=2.68 $Y2=1.645
r94 27 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=1.665
+ $X2=1.58 $Y2=1.665
r95 27 33 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=1.665 $Y=1.665
+ $X2=2.515 $Y2=1.665
r96 24 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=1.75 $X2=1.58
+ $Y2=1.665
r97 24 28 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.58 $Y=1.75 $X2=1.58
+ $Y2=1.95
r98 23 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.58 $Y=1.58 $X2=1.58
+ $Y2=1.665
r99 22 23 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.58 $Y=1.17
+ $X2=1.58 $Y2=1.58
r100 19 28 8.81775 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=1.49 $Y=2.125
+ $X2=1.49 $Y2=1.95
r101 19 21 3.48571 $w=3.5e-07 $l=1e-07 $layer=LI1_cond $X=1.49 $Y=2.125 $X2=1.49
+ $Y2=2.225
r102 15 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.495 $Y=1.085
+ $X2=1.58 $Y2=1.17
r103 15 17 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.495 $Y=1.085
+ $X2=1.3 $Y2=1.085
r104 13 37 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=2.79 $Y=2.39
+ $X2=2.79 $Y2=1.81
r105 9 36 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.715 $Y=0.69
+ $X2=2.715 $Y2=1.48
r106 2 21 600 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=1 $X=1.265
+ $Y=1.84 $X2=1.4 $Y2=2.225
r107 1 17 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.16
+ $Y=0.81 $X2=1.3 $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_1%A_786_100# 1 2 9 14 15 16 19 24 27 29 33 38
+ 40 44 45
c121 38 0 3.96032e-20 $X=4.63 $Y=1.355
c122 27 0 1.45365e-19 $X=6.095 $Y=1.395
c123 24 0 1.34101e-19 $X=6.095 $Y=1.035
c124 14 0 1.3366e-19 $X=4.97 $Y=0.925
r125 45 49 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.88 $Y=1.52
+ $X2=4.88 $Y2=1.685
r126 45 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.88 $Y=1.52
+ $X2=4.88 $Y2=1.355
r127 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.88
+ $Y=1.52 $X2=4.88 $Y2=1.52
r128 41 44 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=4.63 $Y=1.52
+ $X2=4.88 $Y2=1.52
r129 39 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.63 $Y=1.685
+ $X2=4.63 $Y2=1.52
r130 39 40 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.63 $Y=1.685
+ $X2=4.63 $Y2=1.95
r131 38 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.63 $Y=1.355
+ $X2=4.63 $Y2=1.52
r132 37 38 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.63 $Y=1.18
+ $X2=4.63 $Y2=1.355
r133 33 40 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.545 $Y=2.075
+ $X2=4.63 $Y2=1.95
r134 33 35 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=4.545 $Y=2.075
+ $X2=4.085 $Y2=2.075
r135 29 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.545 $Y=1.095
+ $X2=4.63 $Y2=1.18
r136 29 31 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=4.545 $Y=1.095
+ $X2=4.07 $Y2=1.095
r137 22 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.095 $Y=1.32
+ $X2=6.095 $Y2=1.395
r138 22 24 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.095 $Y=1.32
+ $X2=6.095 $Y2=1.035
r139 21 24 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=6.095 $Y=0.265
+ $X2=6.095 $Y2=1.035
r140 17 27 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=5.94 $Y=1.395
+ $X2=6.095 $Y2=1.395
r141 17 19 297.363 $w=1.8e-07 $l=7.65e-07 $layer=POLY_cond $X=5.94 $Y=1.47
+ $X2=5.94 $Y2=2.235
r142 15 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.02 $Y=0.19
+ $X2=6.095 $Y2=0.265
r143 15 16 499.947 $w=1.5e-07 $l=9.75e-07 $layer=POLY_cond $X=6.02 $Y=0.19
+ $X2=5.045 $Y2=0.19
r144 14 48 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.97 $Y=0.925
+ $X2=4.97 $Y2=1.355
r145 11 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.97 $Y=0.265
+ $X2=5.045 $Y2=0.19
r146 11 14 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.97 $Y=0.265
+ $X2=4.97 $Y2=0.925
r147 9 49 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=4.955 $Y=2.285
+ $X2=4.955 $Y2=1.685
r148 2 35 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=3.95
+ $Y=1.84 $X2=4.085 $Y2=2.115
r149 1 31 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=3.93
+ $Y=0.5 $X2=4.07 $Y2=1.095
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_1%B 3 5 7 9 10 11 15 18 20 22 25 28 31 32 34
+ 35 37 41
c128 32 0 1.73263e-19 $X=4.295 $Y=1.515
c129 31 0 1.2613e-19 $X=3.827 $Y=1.515
c130 25 0 1.41099e-19 $X=6.575 $Y=2.335
r131 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.21
+ $Y=1.515 $X2=4.21 $Y2=1.515
r132 37 41 2.67779 $w=6.68e-07 $l=1.5e-07 $layer=LI1_cond $X=4.04 $Y=1.665
+ $X2=4.04 $Y2=1.515
r133 33 34 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.505 $Y=1.69
+ $X2=5.505 $Y2=1.84
r134 32 40 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=4.295 $Y=1.515
+ $X2=4.21 $Y2=1.515
r135 30 40 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=3.95 $Y=1.515
+ $X2=4.21 $Y2=1.515
r136 30 31 3.90195 $w=3.3e-07 $l=1.23e-07 $layer=POLY_cond $X=3.95 $Y=1.515
+ $X2=3.827 $Y2=1.515
r137 28 36 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=6.59 $Y=0.925
+ $X2=6.59 $Y2=1.69
r138 23 25 287.645 $w=1.8e-07 $l=7.4e-07 $layer=POLY_cond $X=6.575 $Y=3.075
+ $X2=6.575 $Y2=2.335
r139 22 36 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=6.575 $Y=1.78
+ $X2=6.575 $Y2=1.69
r140 22 25 215.734 $w=1.8e-07 $l=5.55e-07 $layer=POLY_cond $X=6.575 $Y=1.78
+ $X2=6.575 $Y2=2.335
r141 21 35 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.58 $Y=3.15 $X2=5.49
+ $Y2=3.15
r142 20 23 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.485 $Y=3.15
+ $X2=6.575 $Y2=3.075
r143 20 21 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=6.485 $Y=3.15
+ $X2=5.58 $Y2=3.15
r144 18 33 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=5.535 $Y=0.925
+ $X2=5.535 $Y2=1.69
r145 15 34 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=5.49 $Y=2.235
+ $X2=5.49 $Y2=1.84
r146 13 35 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=5.49 $Y=3.075
+ $X2=5.49 $Y2=3.15
r147 13 15 326.516 $w=1.8e-07 $l=8.4e-07 $layer=POLY_cond $X=5.49 $Y=3.075
+ $X2=5.49 $Y2=2.235
r148 10 35 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.4 $Y=3.15 $X2=5.49
+ $Y2=3.15
r149 10 11 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=5.4 $Y=3.15
+ $X2=4.445 $Y2=3.15
r150 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.37 $Y=3.075
+ $X2=4.445 $Y2=3.15
r151 8 32 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.37 $Y=1.68
+ $X2=4.295 $Y2=1.515
r152 8 9 715.309 $w=1.5e-07 $l=1.395e-06 $layer=POLY_cond $X=4.37 $Y=1.68
+ $X2=4.37 $Y2=3.075
r153 5 31 34.7346 $w=1.65e-07 $l=1.78452e-07 $layer=POLY_cond $X=3.855 $Y=1.35
+ $X2=3.827 $Y2=1.515
r154 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.855 $Y=1.35
+ $X2=3.855 $Y2=0.87
r155 1 31 34.7346 $w=1.65e-07 $l=1.80748e-07 $layer=POLY_cond $X=3.86 $Y=1.68
+ $X2=3.827 $Y2=1.515
r156 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.86 $Y=1.68 $X2=3.86
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_1%A 3 7 9 12
c44 12 0 3.49804e-19 $X=7.04 $Y=1.59
c45 9 0 2.38837e-20 $X=6.96 $Y=1.665
c46 3 0 4.37781e-20 $X=7.085 $Y=0.925
r47 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.04 $Y=1.59
+ $X2=7.04 $Y2=1.755
r48 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.04 $Y=1.59
+ $X2=7.04 $Y2=1.425
r49 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.04
+ $Y=1.59 $X2=7.04 $Y2=1.59
r50 7 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=7.115 $Y=2.415
+ $X2=7.115 $Y2=1.755
r51 3 14 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=7.085 $Y=0.925
+ $X2=7.085 $Y2=1.425
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_1%A_897_54# 1 2 3 4 15 19 21 23 28 29 30 31 32
+ 33 38 42 44 51 52 53
c125 52 0 1.54564e-19 $X=7.58 $Y=1.59
c126 15 0 2.38837e-20 $X=7.65 $Y=2.415
r127 52 57 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.58 $Y=1.59
+ $X2=7.58 $Y2=1.755
r128 52 56 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.58 $Y=1.59
+ $X2=7.58 $Y2=1.425
r129 51 54 8.01359 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=7.54 $Y=1.59
+ $X2=7.54 $Y2=1.755
r130 51 53 8.01359 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=7.54 $Y=1.59
+ $X2=7.54 $Y2=1.425
r131 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.58
+ $Y=1.59 $X2=7.58 $Y2=1.59
r132 44 46 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=4.655 $Y=2.795
+ $X2=4.655 $Y2=2.99
r133 40 42 10.0285 $w=2.43e-07 $l=1.9e-07 $layer=LI1_cond $X=4.65 $Y=0.377
+ $X2=4.84 $Y2=0.377
r134 38 54 10.5499 $w=2.03e-07 $l=1.95e-07 $layer=LI1_cond $X=7.517 $Y=1.95
+ $X2=7.517 $Y2=1.755
r135 35 53 9.19734 $w=2.03e-07 $l=1.7e-07 $layer=LI1_cond $X=7.517 $Y=1.255
+ $X2=7.517 $Y2=1.425
r136 34 49 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.09 $Y=2.035
+ $X2=6.925 $Y2=2.035
r137 33 38 6.89401 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=7.415 $Y=2.035
+ $X2=7.517 $Y2=1.95
r138 33 34 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.415 $Y=2.035
+ $X2=7.09 $Y2=2.035
r139 31 35 6.89401 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=7.415 $Y=1.17
+ $X2=7.517 $Y2=1.255
r140 31 32 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=7.415 $Y=1.17
+ $X2=7.035 $Y2=1.17
r141 29 49 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.925 $Y=2.12
+ $X2=6.925 $Y2=2.035
r142 29 30 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=6.925 $Y=2.12
+ $X2=6.925 $Y2=2.905
r143 26 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.87 $Y=1.085
+ $X2=7.035 $Y2=1.17
r144 26 28 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.87 $Y=1.085
+ $X2=6.87 $Y2=0.75
r145 25 28 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=6.87 $Y=0.425
+ $X2=6.87 $Y2=0.75
r146 23 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.705 $Y=0.34
+ $X2=6.87 $Y2=0.425
r147 23 42 121.674 $w=1.68e-07 $l=1.865e-06 $layer=LI1_cond $X=6.705 $Y=0.34
+ $X2=4.84 $Y2=0.34
r148 22 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.82 $Y=2.99
+ $X2=4.655 $Y2=2.99
r149 21 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.76 $Y=2.99
+ $X2=6.925 $Y2=2.905
r150 21 22 126.567 $w=1.68e-07 $l=1.94e-06 $layer=LI1_cond $X=6.76 $Y=2.99
+ $X2=4.82 $Y2=2.99
r151 19 56 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=7.665 $Y=0.925
+ $X2=7.665 $Y2=1.425
r152 15 57 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=7.65 $Y=2.415
+ $X2=7.65 $Y2=1.755
r153 4 49 300 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_PDIFF $count=2 $X=6.665
+ $Y=1.915 $X2=6.885 $Y2=2.115
r154 3 44 600 $w=1.7e-07 $l=9.95214e-07 $layer=licon1_PDIFF $count=1 $X=4.52
+ $Y=1.865 $X2=4.655 $Y2=2.795
r155 2 28 91 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=2 $X=6.665
+ $Y=0.605 $X2=6.87 $Y2=0.75
r156 1 40 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=4.485
+ $Y=0.27 $X2=4.65 $Y2=0.415
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_1%X 1 2 9 11 15 16 17 28
c21 16 0 1.63453e-19 $X=0.24 $Y=0.555
r22 21 28 2.0808 $w=3.58e-07 $l=6.5e-08 $layer=LI1_cond $X=0.265 $Y=0.99
+ $X2=0.265 $Y2=0.925
r23 17 30 8.67109 $w=3.58e-07 $l=1.7e-07 $layer=LI1_cond $X=0.265 $Y=1 $X2=0.265
+ $Y2=1.17
r24 17 21 0.320123 $w=3.58e-07 $l=1e-08 $layer=LI1_cond $X=0.265 $Y=1 $X2=0.265
+ $Y2=0.99
r25 17 28 0.320123 $w=3.58e-07 $l=1e-08 $layer=LI1_cond $X=0.265 $Y=0.915
+ $X2=0.265 $Y2=0.925
r26 16 17 11.5244 $w=3.58e-07 $l=3.6e-07 $layer=LI1_cond $X=0.265 $Y=0.555
+ $X2=0.265 $Y2=0.915
r27 15 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.17 $Y=1.84
+ $X2=0.17 $Y2=1.17
r28 11 13 34.5733 $w=2.68e-07 $l=8.1e-07 $layer=LI1_cond $X=0.22 $Y=2.005
+ $X2=0.22 $Y2=2.815
r29 9 15 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.22 $Y=1.975
+ $X2=0.22 $Y2=1.84
r30 9 11 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=0.22 $Y=1.975 $X2=0.22
+ $Y2=2.005
r31 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.815
r32 2 11 400 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.27 $Y2=2.005
r33 1 16 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.49 $X2=0.28 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_1%VPWR 1 2 3 12 16 20 22 24 29 37 47 48 51 54
+ 57
c76 20 0 1.41099e-19 $X=7.425 $Y=2.375
r77 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r78 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r79 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r80 48 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r81 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r82 45 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.59 $Y=3.33
+ $X2=7.425 $Y2=3.33
r83 45 47 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.59 $Y=3.33
+ $X2=7.92 $Y2=3.33
r84 44 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r85 43 44 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r86 40 43 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=6.96 $Y2=3.33
r87 38 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.725 $Y=3.33
+ $X2=3.56 $Y2=3.33
r88 38 40 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.725 $Y=3.33
+ $X2=4.08 $Y2=3.33
r89 37 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.26 $Y=3.33
+ $X2=7.425 $Y2=3.33
r90 37 43 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=7.26 $Y=3.33 $X2=6.96
+ $Y2=3.33
r91 36 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r92 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r93 33 36 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r94 33 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r95 32 35 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r96 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r97 30 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=0.68 $Y2=3.33
r98 30 32 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=1.2 $Y2=3.33
r99 29 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.395 $Y=3.33
+ $X2=3.56 $Y2=3.33
r100 29 35 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.395 $Y=3.33
+ $X2=3.12 $Y2=3.33
r101 27 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r102 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r103 24 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.68 $Y2=3.33
r104 24 26 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=3.33
+ $X2=0.24 $Y2=3.33
r105 22 44 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=6.96 $Y2=3.33
r106 22 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r107 22 40 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r108 18 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.425 $Y=3.245
+ $X2=7.425 $Y2=3.33
r109 18 20 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=7.425 $Y=3.245
+ $X2=7.425 $Y2=2.375
r110 14 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.56 $Y=3.245
+ $X2=3.56 $Y2=3.33
r111 14 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.56 $Y=3.245
+ $X2=3.56 $Y2=2.875
r112 10 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=3.245
+ $X2=0.68 $Y2=3.33
r113 10 12 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=0.68 $Y=3.245
+ $X2=0.68 $Y2=2.455
r114 3 20 300 $w=1.7e-07 $l=5.59285e-07 $layer=licon1_PDIFF $count=2 $X=7.205
+ $Y=1.915 $X2=7.425 $Y2=2.375
r115 2 16 600 $w=1.7e-07 $l=1.10043e-06 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=1.84 $X2=3.56 $Y2=2.875
r116 1 12 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.84 $X2=0.72 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_1%A_363_394# 1 2 3 4 15 17 18 20 22 23 27 29
+ 33 38 39 40
c131 29 0 4.37781e-20 $X=6.255 $Y=0.68
c132 23 0 1.2613e-19 $X=5.015 $Y=2.455
r133 39 40 7.99654 $w=2.43e-07 $l=1.7e-07 $layer=LI1_cond $X=5.01 $Y=0.717
+ $X2=5.18 $Y2=0.717
r134 36 37 13.7351 $w=4.53e-07 $l=5.1e-07 $layer=LI1_cond $X=2.93 $Y=0.67
+ $X2=3.44 $Y2=0.67
r135 31 33 11.5244 $w=2.78e-07 $l=2.8e-07 $layer=LI1_cond $X=6.395 $Y=0.765
+ $X2=6.395 $Y2=1.045
r136 29 31 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=6.255 $Y=0.68
+ $X2=6.395 $Y2=0.765
r137 29 40 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=6.255 $Y=0.68
+ $X2=5.18 $Y2=0.68
r138 25 27 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=5.14 $Y=2.37
+ $X2=5.14 $Y2=2.02
r139 24 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.525 $Y=2.455
+ $X2=3.44 $Y2=2.455
r140 23 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.015 $Y=2.455
+ $X2=5.14 $Y2=2.37
r141 23 24 97.2086 $w=1.68e-07 $l=1.49e-06 $layer=LI1_cond $X=5.015 $Y=2.455
+ $X2=3.525 $Y2=2.455
r142 22 37 7.27104 $w=4.53e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.525 $Y=0.755
+ $X2=3.44 $Y2=0.67
r143 22 39 96.8824 $w=1.68e-07 $l=1.485e-06 $layer=LI1_cond $X=3.525 $Y=0.755
+ $X2=5.01 $Y2=0.755
r144 20 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=2.37
+ $X2=3.44 $Y2=2.455
r145 19 37 6.54142 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=3.44 $Y=0.97 $X2=3.44
+ $Y2=0.67
r146 19 20 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=3.44 $Y=0.97
+ $X2=3.44 $Y2=2.37
r147 17 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=2.455
+ $X2=3.44 $Y2=2.455
r148 17 18 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=3.355 $Y=2.455
+ $X2=2.125 $Y2=2.455
r149 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2 $Y=2.37
+ $X2=2.125 $Y2=2.455
r150 13 15 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=2 $Y=2.37 $X2=2
+ $Y2=2.115
r151 4 27 300 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=2 $X=5.045
+ $Y=1.865 $X2=5.18 $Y2=2.02
r152 3 15 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.815
+ $Y=1.97 $X2=1.96 $Y2=2.115
r153 2 33 182 $w=1.7e-07 $l=3.05778e-07 $layer=licon1_NDIFF $count=1 $X=6.17
+ $Y=0.825 $X2=6.375 $Y2=1.045
r154 1 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.79
+ $Y=0.37 $X2=2.93 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_1%A_371_74# 1 2 3 4 15 17 20 21 25 26 27 28 31
+ 34 37 38 44 47
c126 25 0 2.79465e-19 $X=5.52 $Y=1.41
r127 47 48 2.97244 $w=4.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=1.225
+ $X2=2.055 $Y2=1.14
r128 45 51 9.95397 $w=2.39e-07 $l=1.95e-07 $layer=LI1_cond $X=5.46 $Y=1.295
+ $X2=5.46 $Y2=1.1
r129 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.295
+ $X2=5.52 $Y2=1.295
r130 41 47 1.83343 $w=4.38e-07 $l=7e-08 $layer=LI1_cond $X=2.055 $Y=1.295
+ $X2=2.055 $Y2=1.225
r131 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=1.295
+ $X2=2.16 $Y2=1.295
r132 38 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=1.295
+ $X2=2.16 $Y2=1.295
r133 37 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=1.295
+ $X2=5.52 $Y2=1.295
r134 37 38 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=5.375 $Y=1.295
+ $X2=2.305 $Y2=1.295
r135 29 31 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.165 $Y=1.935
+ $X2=6.165 $Y2=2.195
r136 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.08 $Y=1.85
+ $X2=6.165 $Y2=1.935
r137 27 28 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=6.08 $Y=1.85
+ $X2=5.605 $Y2=1.85
r138 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.52 $Y=1.765
+ $X2=5.605 $Y2=1.85
r139 25 45 6.90437 $w=2.39e-07 $l=1.41863e-07 $layer=LI1_cond $X=5.52 $Y=1.41
+ $X2=5.46 $Y2=1.295
r140 25 26 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.52 $Y=1.41
+ $X2=5.52 $Y2=1.765
r141 21 51 2.73298 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=5.315 $Y=1.1
+ $X2=5.46 $Y2=1.1
r142 21 23 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.315 $Y=1.1
+ $X2=5.25 $Y2=1.1
r143 20 34 0.716491 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.1 $Y=2.03
+ $X2=3.015 $Y2=2.115
r144 19 20 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.1 $Y=1.31 $X2=3.1
+ $Y2=2.03
r145 18 47 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=2.275 $Y=1.225
+ $X2=2.055 $Y2=1.225
r146 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.015 $Y=1.225
+ $X2=3.1 $Y2=1.31
r147 17 18 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=3.015 $Y=1.225
+ $X2=2.275 $Y2=1.225
r148 15 48 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2 $Y=0.81 $X2=2
+ $Y2=1.14
r149 4 31 600 $w=1.7e-07 $l=3.40881e-07 $layer=licon1_PDIFF $count=1 $X=6.03
+ $Y=1.915 $X2=6.165 $Y2=2.195
r150 3 34 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.88
+ $Y=1.97 $X2=3.015 $Y2=2.115
r151 2 23 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=5.045
+ $Y=0.605 $X2=5.25 $Y2=1.1
r152 1 15 182 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_NDIFF $count=1 $X=1.855
+ $Y=0.37 $X2=2 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_1%A_1116_383# 1 2 3 4 15 17 18 19 20 22 23 25
+ 29 35 36 37 43 44 47
c115 36 0 1.54564e-19 $X=7.775 $Y=1.295
c116 22 0 1.71138e-19 $X=6.505 $Y=2.565
c117 19 0 1.78665e-19 $X=6.42 $Y=1.51
r118 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=1.295
+ $X2=7.92 $Y2=1.295
r119 40 47 7.24924 $w=3.08e-07 $l=1.95e-07 $layer=LI1_cond $X=5.93 $Y=1.295
+ $X2=5.93 $Y2=1.1
r120 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=1.295 $X2=6
+ $Y2=1.295
r121 37 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.145 $Y=1.295
+ $X2=6 $Y2=1.295
r122 36 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=1.295
+ $X2=7.92 $Y2=1.295
r123 36 37 2.01732 $w=1.4e-07 $l=1.63e-06 $layer=MET1_cond $X=7.775 $Y=1.295
+ $X2=6.145 $Y2=1.295
r124 35 44 1.92074 $w=2.38e-07 $l=4e-08 $layer=LI1_cond $X=7.955 $Y=1.255
+ $X2=7.955 $Y2=1.295
r125 33 44 42.9765 $w=2.38e-07 $l=8.95e-07 $layer=LI1_cond $X=7.955 $Y=2.19
+ $X2=7.955 $Y2=1.295
r126 31 40 4.83283 $w=3.08e-07 $l=1.3e-07 $layer=LI1_cond $X=5.93 $Y=1.425
+ $X2=5.93 $Y2=1.295
r127 27 35 6.02978 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=7.935 $Y=1.115
+ $X2=7.935 $Y2=1.255
r128 27 29 15.0229 $w=2.78e-07 $l=3.65e-07 $layer=LI1_cond $X=7.935 $Y=1.115
+ $X2=7.935 $Y2=0.75
r129 23 33 6.0629 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=7.932 $Y=2.332
+ $X2=7.932 $Y2=2.19
r130 23 25 0.930042 $w=2.83e-07 $l=2.3e-08 $layer=LI1_cond $X=7.932 $Y=2.332
+ $X2=7.932 $Y2=2.355
r131 21 22 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=6.505 $Y=1.595
+ $X2=6.505 $Y2=2.565
r132 20 31 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=6.085 $Y=1.51
+ $X2=5.93 $Y2=1.425
r133 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.42 $Y=1.51
+ $X2=6.505 $Y2=1.595
r134 19 20 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.42 $Y=1.51
+ $X2=6.085 $Y2=1.51
r135 17 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.42 $Y=2.65
+ $X2=6.505 $Y2=2.565
r136 17 18 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=6.42 $Y=2.65
+ $X2=5.88 $Y2=2.65
r137 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.715 $Y=2.565
+ $X2=5.88 $Y2=2.65
r138 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.715 $Y=2.565
+ $X2=5.715 $Y2=2.27
r139 4 25 300 $w=1.7e-07 $l=5.02991e-07 $layer=licon1_PDIFF $count=2 $X=7.74
+ $Y=1.915 $X2=7.875 $Y2=2.355
r140 3 15 600 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_PDIFF $count=1 $X=5.58
+ $Y=1.915 $X2=5.715 $Y2=2.27
r141 2 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.74
+ $Y=0.605 $X2=7.88 $Y2=0.75
r142 1 47 182 $w=1.7e-07 $l=6.07268e-07 $layer=licon1_NDIFF $count=1 $X=5.61
+ $Y=0.605 $X2=5.86 $Y2=1.1
.ends

.subckt PM_SKY130_FD_SC_MS__XNOR3_1%VGND 1 2 3 12 16 20 22 24 29 37 47 48 51 54
+ 57
r72 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r73 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r74 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r75 48 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r76 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r77 45 57 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=7.615 $Y=0 $X2=7.41
+ $Y2=0
r78 45 47 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.615 $Y=0 $X2=7.92
+ $Y2=0
r79 44 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r80 43 44 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r81 40 43 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6.96
+ $Y2=0
r82 38 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.725 $Y=0 $X2=3.56
+ $Y2=0
r83 38 40 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.725 $Y=0 $X2=4.08
+ $Y2=0
r84 37 57 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=7.205 $Y=0 $X2=7.41
+ $Y2=0
r85 37 43 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.205 $Y=0 $X2=6.96
+ $Y2=0
r86 36 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r87 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r88 33 36 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r89 33 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r90 32 35 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r91 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r92 30 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=0.79
+ $Y2=0
r93 30 32 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=0 $X2=1.2
+ $Y2=0
r94 29 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.395 $Y=0 $X2=3.56
+ $Y2=0
r95 29 35 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.395 $Y=0 $X2=3.12
+ $Y2=0
r96 27 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r97 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r98 24 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.79
+ $Y2=0
r99 24 26 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=0 $X2=0.24
+ $Y2=0
r100 22 44 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=6.96 $Y2=0
r101 22 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r102 22 40 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r103 18 57 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=7.41 $Y=0.085
+ $X2=7.41 $Y2=0
r104 18 20 18.6921 $w=4.08e-07 $l=6.65e-07 $layer=LI1_cond $X=7.41 $Y=0.085
+ $X2=7.41 $Y2=0.75
r105 14 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.56 $Y=0.085
+ $X2=3.56 $Y2=0
r106 14 16 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=3.56 $Y=0.085
+ $X2=3.56 $Y2=0.335
r107 10 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0
r108 10 12 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.79 $Y=0.085
+ $X2=0.79 $Y2=0.325
r109 3 20 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=7.16
+ $Y=0.605 $X2=7.41 $Y2=0.75
r110 2 16 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=3.415
+ $Y=0.19 $X2=3.56 $Y2=0.335
r111 1 12 182 $w=1.7e-07 $l=2.91033e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.49 $X2=0.79 $Y2=0.325
.ends


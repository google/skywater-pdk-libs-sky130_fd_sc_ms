* File: sky130_fd_sc_ms__clkbuf_16.pex.spice
* Created: Wed Sep  2 12:00:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__CLKBUF_16%A 3 7 11 15 19 23 27 31 33 34 35 36 55
c87 31 0 1.47622e-19 $X=1.86 $Y=2.4
r88 54 55 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=1.805 $Y=1.515
+ $X2=1.86 $Y2=1.515
r89 52 54 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=1.605 $Y=1.515
+ $X2=1.805 $Y2=1.515
r90 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.605
+ $Y=1.515 $X2=1.605 $Y2=1.515
r91 50 52 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.41 $Y=1.515
+ $X2=1.605 $Y2=1.515
r92 49 50 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=1.375 $Y=1.515
+ $X2=1.41 $Y2=1.515
r93 48 49 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=0.96 $Y=1.515
+ $X2=1.375 $Y2=1.515
r94 47 48 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=0.925 $Y=1.515
+ $X2=0.96 $Y2=1.515
r95 45 47 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.585 $Y=1.515
+ $X2=0.925 $Y2=1.515
r96 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.585
+ $Y=1.515 $X2=0.585 $Y2=1.515
r97 43 45 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.51 $Y=1.515
+ $X2=0.585 $Y2=1.515
r98 41 43 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.515
+ $X2=0.51 $Y2=1.515
r99 36 53 2.01008 $w=4.28e-07 $l=7.5e-08 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=1.605 $Y2=1.565
r100 35 53 10.8544 $w=4.28e-07 $l=4.05e-07 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.605 $Y2=1.565
r101 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r102 34 46 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.585 $Y2=1.565
r103 33 46 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.585 $Y2=1.565
r104 29 55 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.86 $Y=1.68
+ $X2=1.86 $Y2=1.515
r105 29 31 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.86 $Y=1.68
+ $X2=1.86 $Y2=2.4
r106 25 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.805 $Y=1.35
+ $X2=1.805 $Y2=1.515
r107 25 27 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=1.805 $Y=1.35
+ $X2=1.805 $Y2=0.58
r108 21 50 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.68
+ $X2=1.41 $Y2=1.515
r109 21 23 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.41 $Y=1.68
+ $X2=1.41 $Y2=2.4
r110 17 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=1.35
+ $X2=1.375 $Y2=1.515
r111 17 19 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=1.375 $Y=1.35
+ $X2=1.375 $Y2=0.58
r112 13 48 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.96 $Y=1.68
+ $X2=0.96 $Y2=1.515
r113 13 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.96 $Y=1.68
+ $X2=0.96 $Y2=2.4
r114 9 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=1.515
r115 9 11 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=0.925 $Y2=0.58
r116 5 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=1.68
+ $X2=0.51 $Y2=1.515
r117 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.51 $Y=1.68 $X2=0.51
+ $Y2=2.4
r118 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=1.515
r119 1 3 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__CLKBUF_16%A_114_74# 1 2 3 4 15 19 23 27 31 35 39 43
+ 47 51 55 59 63 67 71 75 79 83 87 91 95 99 103 107 111 115 119 123 127 131 135
+ 139 143 145 147 149 150 151 155 159 161 163 164 167 170 178 181 184 187 190
+ 193 195 196 251
c439 251 0 1.81624e-20 $X=9.105 $Y=1.355
r440 250 251 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=9.09 $Y=1.355
+ $X2=9.105 $Y2=1.355
r441 249 250 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=8.675 $Y=1.355
+ $X2=9.09 $Y2=1.355
r442 248 249 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=8.64 $Y=1.355
+ $X2=8.675 $Y2=1.355
r443 246 248 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=8.39 $Y=1.355
+ $X2=8.64 $Y2=1.355
r444 244 246 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=8.175 $Y=1.355
+ $X2=8.39 $Y2=1.355
r445 243 244 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=8.17 $Y=1.355
+ $X2=8.175 $Y2=1.355
r446 242 243 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=7.745 $Y=1.355
+ $X2=8.17 $Y2=1.355
r447 241 242 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=7.72 $Y=1.355
+ $X2=7.745 $Y2=1.355
r448 239 241 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=7.46 $Y=1.355
+ $X2=7.72 $Y2=1.355
r449 237 239 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=7.27 $Y=1.355
+ $X2=7.46 $Y2=1.355
r450 236 237 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=7.245 $Y=1.355
+ $X2=7.27 $Y2=1.355
r451 235 236 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=6.82 $Y=1.355
+ $X2=7.245 $Y2=1.355
r452 234 235 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=6.815 $Y=1.355
+ $X2=6.82 $Y2=1.355
r453 232 234 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=6.53 $Y=1.355
+ $X2=6.815 $Y2=1.355
r454 230 232 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=6.37 $Y=1.355
+ $X2=6.53 $Y2=1.355
r455 229 230 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=6.315 $Y=1.355
+ $X2=6.37 $Y2=1.355
r456 228 229 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=5.92 $Y=1.355
+ $X2=6.315 $Y2=1.355
r457 227 228 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=5.885 $Y=1.355
+ $X2=5.92 $Y2=1.355
r458 225 227 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=5.59 $Y=1.355
+ $X2=5.885 $Y2=1.355
r459 223 225 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=5.47 $Y=1.355
+ $X2=5.59 $Y2=1.355
r460 222 223 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=5.385 $Y=1.355
+ $X2=5.47 $Y2=1.355
r461 221 222 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=5.02 $Y=1.355
+ $X2=5.385 $Y2=1.355
r462 220 221 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=4.955 $Y=1.355
+ $X2=5.02 $Y2=1.355
r463 218 220 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=4.675 $Y=1.355
+ $X2=4.955 $Y2=1.355
r464 216 218 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=4.57 $Y=1.355
+ $X2=4.675 $Y2=1.355
r465 215 216 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=4.455 $Y=1.355
+ $X2=4.57 $Y2=1.355
r466 214 215 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=4.12 $Y=1.355
+ $X2=4.455 $Y2=1.355
r467 213 214 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=4.025 $Y=1.355
+ $X2=4.12 $Y2=1.355
r468 211 213 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=3.835 $Y=1.355
+ $X2=4.025 $Y2=1.355
r469 209 211 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.355
+ $X2=3.835 $Y2=1.355
r470 208 209 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.595 $Y=1.355
+ $X2=3.67 $Y2=1.355
r471 207 208 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=3.22 $Y=1.355
+ $X2=3.595 $Y2=1.355
r472 206 207 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=3.165 $Y=1.355
+ $X2=3.22 $Y2=1.355
r473 204 206 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=2.975 $Y=1.355
+ $X2=3.165 $Y2=1.355
r474 202 204 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=2.77 $Y=1.355
+ $X2=2.975 $Y2=1.355
r475 201 202 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=2.735 $Y=1.355
+ $X2=2.77 $Y2=1.355
r476 200 201 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=2.32 $Y=1.355
+ $X2=2.735 $Y2=1.355
r477 198 200 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.305 $Y=1.355
+ $X2=2.32 $Y2=1.355
r478 196 246 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.39
+ $Y=1.355 $X2=8.39 $Y2=1.355
r479 195 196 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.39 $Y=1.295
+ $X2=8.39 $Y2=1.295
r480 193 239 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.46
+ $Y=1.355 $X2=7.46 $Y2=1.355
r481 192 195 0.596692 $w=2.3e-07 $l=9.3e-07 $layer=MET1_cond $X=7.46 $Y=1.295
+ $X2=8.39 $Y2=1.295
r482 192 193 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.46 $Y=1.295
+ $X2=7.46 $Y2=1.295
r483 190 232 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.53
+ $Y=1.355 $X2=6.53 $Y2=1.355
r484 189 192 0.596692 $w=2.3e-07 $l=9.3e-07 $layer=MET1_cond $X=6.53 $Y=1.295
+ $X2=7.46 $Y2=1.295
r485 189 190 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.53 $Y=1.295
+ $X2=6.53 $Y2=1.295
r486 187 225 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.59
+ $Y=1.355 $X2=5.59 $Y2=1.355
r487 186 189 0.603108 $w=2.3e-07 $l=9.4e-07 $layer=MET1_cond $X=5.59 $Y=1.295
+ $X2=6.53 $Y2=1.295
r488 186 187 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.59 $Y=1.295
+ $X2=5.59 $Y2=1.295
r489 184 218 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.675
+ $Y=1.355 $X2=4.675 $Y2=1.355
r490 183 186 0.587068 $w=2.3e-07 $l=9.15e-07 $layer=MET1_cond $X=4.675 $Y=1.295
+ $X2=5.59 $Y2=1.295
r491 183 184 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.675 $Y=1.295
+ $X2=4.675 $Y2=1.295
r492 181 211 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.835
+ $Y=1.355 $X2=3.835 $Y2=1.355
r493 180 183 0.538948 $w=2.3e-07 $l=8.4e-07 $layer=MET1_cond $X=3.835 $Y=1.295
+ $X2=4.675 $Y2=1.295
r494 180 181 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.835 $Y=1.295
+ $X2=3.835 $Y2=1.295
r495 178 204 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.975
+ $Y=1.355 $X2=2.975 $Y2=1.355
r496 177 180 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=2.975 $Y=1.295
+ $X2=3.835 $Y2=1.295
r497 177 178 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.975 $Y=1.295
+ $X2=2.975 $Y2=1.295
r498 174 274 13.3619 $w=2.1e-07 $l=2.3e-07 $layer=LI1_cond $X=2.087 $Y=1.295
+ $X2=2.087 $Y2=1.065
r499 173 177 0.564612 $w=2.3e-07 $l=8.8e-07 $layer=MET1_cond $X=2.095 $Y=1.295
+ $X2=2.975 $Y2=1.295
r500 173 174 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.095 $Y=1.295
+ $X2=2.095 $Y2=1.295
r501 169 170 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.635 $Y=2.035
+ $X2=2.05 $Y2=2.035
r502 164 170 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=1.95
+ $X2=2.05 $Y2=2.035
r503 163 174 7.15932 $w=2.1e-07 $l=1.32212e-07 $layer=LI1_cond $X=2.05 $Y=1.41
+ $X2=2.087 $Y2=1.295
r504 163 164 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.05 $Y=1.41
+ $X2=2.05 $Y2=1.95
r505 162 167 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.675 $Y=1.065
+ $X2=1.55 $Y2=1.065
r506 161 274 1.9771 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=1.965 $Y=1.065
+ $X2=2.087 $Y2=1.065
r507 161 162 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.965 $Y=1.065
+ $X2=1.675 $Y2=1.065
r508 159 169 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.635 $Y=2.815
+ $X2=1.635 $Y2=2.12
r509 153 167 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=0.98
+ $X2=1.55 $Y2=1.065
r510 153 155 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=1.55 $Y=0.98
+ $X2=1.55 $Y2=0.58
r511 152 166 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.9 $Y=2.035
+ $X2=0.735 $Y2=2.035
r512 151 169 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.47 $Y=2.035
+ $X2=1.635 $Y2=2.035
r513 151 152 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.47 $Y=2.035
+ $X2=0.9 $Y2=2.035
r514 149 167 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.425 $Y=1.065
+ $X2=1.55 $Y2=1.065
r515 149 150 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.425 $Y=1.065
+ $X2=0.795 $Y2=1.065
r516 145 166 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=2.12
+ $X2=0.735 $Y2=2.035
r517 145 147 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.735 $Y=2.12
+ $X2=0.735 $Y2=2.815
r518 141 150 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.67 $Y=0.98
+ $X2=0.795 $Y2=1.065
r519 141 143 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=0.67 $Y=0.98
+ $X2=0.67 $Y2=0.58
r520 137 251 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.105 $Y=1.19
+ $X2=9.105 $Y2=1.355
r521 137 139 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.105 $Y=1.19
+ $X2=9.105 $Y2=0.58
r522 133 250 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.09 $Y=1.52
+ $X2=9.09 $Y2=1.355
r523 133 135 342.065 $w=1.8e-07 $l=8.8e-07 $layer=POLY_cond $X=9.09 $Y=1.52
+ $X2=9.09 $Y2=2.4
r524 129 249 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.675 $Y=1.19
+ $X2=8.675 $Y2=1.355
r525 129 131 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.675 $Y=1.19
+ $X2=8.675 $Y2=0.58
r526 125 248 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.64 $Y=1.52
+ $X2=8.64 $Y2=1.355
r527 125 127 342.065 $w=1.8e-07 $l=8.8e-07 $layer=POLY_cond $X=8.64 $Y=1.52
+ $X2=8.64 $Y2=2.4
r528 121 244 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.175 $Y=1.19
+ $X2=8.175 $Y2=1.355
r529 121 123 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.175 $Y=1.19
+ $X2=8.175 $Y2=0.58
r530 117 243 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.17 $Y=1.52
+ $X2=8.17 $Y2=1.355
r531 117 119 342.065 $w=1.8e-07 $l=8.8e-07 $layer=POLY_cond $X=8.17 $Y=1.52
+ $X2=8.17 $Y2=2.4
r532 113 242 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.745 $Y=1.19
+ $X2=7.745 $Y2=1.355
r533 113 115 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.745 $Y=1.19
+ $X2=7.745 $Y2=0.58
r534 109 241 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.72 $Y=1.52
+ $X2=7.72 $Y2=1.355
r535 109 111 342.065 $w=1.8e-07 $l=8.8e-07 $layer=POLY_cond $X=7.72 $Y=1.52
+ $X2=7.72 $Y2=2.4
r536 105 237 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.27 $Y=1.52
+ $X2=7.27 $Y2=1.355
r537 105 107 342.065 $w=1.8e-07 $l=8.8e-07 $layer=POLY_cond $X=7.27 $Y=1.52
+ $X2=7.27 $Y2=2.4
r538 101 236 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.245 $Y=1.19
+ $X2=7.245 $Y2=1.355
r539 101 103 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.245 $Y=1.19
+ $X2=7.245 $Y2=0.58
r540 97 234 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.815 $Y=1.19
+ $X2=6.815 $Y2=1.355
r541 97 99 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.815 $Y=1.19
+ $X2=6.815 $Y2=0.58
r542 93 235 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.82 $Y=1.52
+ $X2=6.82 $Y2=1.355
r543 93 95 342.065 $w=1.8e-07 $l=8.8e-07 $layer=POLY_cond $X=6.82 $Y=1.52
+ $X2=6.82 $Y2=2.4
r544 89 230 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.37 $Y=1.52
+ $X2=6.37 $Y2=1.355
r545 89 91 342.065 $w=1.8e-07 $l=8.8e-07 $layer=POLY_cond $X=6.37 $Y=1.52
+ $X2=6.37 $Y2=2.4
r546 85 229 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.315 $Y=1.19
+ $X2=6.315 $Y2=1.355
r547 85 87 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.315 $Y=1.19
+ $X2=6.315 $Y2=0.58
r548 81 228 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.92 $Y=1.52
+ $X2=5.92 $Y2=1.355
r549 81 83 342.065 $w=1.8e-07 $l=8.8e-07 $layer=POLY_cond $X=5.92 $Y=1.52
+ $X2=5.92 $Y2=2.4
r550 77 227 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.885 $Y=1.19
+ $X2=5.885 $Y2=1.355
r551 77 79 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.885 $Y=1.19
+ $X2=5.885 $Y2=0.58
r552 73 223 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.47 $Y=1.52
+ $X2=5.47 $Y2=1.355
r553 73 75 342.065 $w=1.8e-07 $l=8.8e-07 $layer=POLY_cond $X=5.47 $Y=1.52
+ $X2=5.47 $Y2=2.4
r554 69 222 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.385 $Y=1.19
+ $X2=5.385 $Y2=1.355
r555 69 71 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.385 $Y=1.19
+ $X2=5.385 $Y2=0.58
r556 65 221 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.02 $Y=1.52
+ $X2=5.02 $Y2=1.355
r557 65 67 342.065 $w=1.8e-07 $l=8.8e-07 $layer=POLY_cond $X=5.02 $Y=1.52
+ $X2=5.02 $Y2=2.4
r558 61 220 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.955 $Y=1.19
+ $X2=4.955 $Y2=1.355
r559 61 63 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.955 $Y=1.19
+ $X2=4.955 $Y2=0.58
r560 57 216 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.57 $Y=1.52
+ $X2=4.57 $Y2=1.355
r561 57 59 342.065 $w=1.8e-07 $l=8.8e-07 $layer=POLY_cond $X=4.57 $Y=1.52
+ $X2=4.57 $Y2=2.4
r562 53 215 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.455 $Y=1.19
+ $X2=4.455 $Y2=1.355
r563 53 55 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.455 $Y=1.19
+ $X2=4.455 $Y2=0.58
r564 49 214 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.12 $Y=1.52
+ $X2=4.12 $Y2=1.355
r565 49 51 342.065 $w=1.8e-07 $l=8.8e-07 $layer=POLY_cond $X=4.12 $Y=1.52
+ $X2=4.12 $Y2=2.4
r566 45 213 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.025 $Y=1.19
+ $X2=4.025 $Y2=1.355
r567 45 47 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.025 $Y=1.19
+ $X2=4.025 $Y2=0.58
r568 41 209 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.52
+ $X2=3.67 $Y2=1.355
r569 41 43 342.065 $w=1.8e-07 $l=8.8e-07 $layer=POLY_cond $X=3.67 $Y=1.52
+ $X2=3.67 $Y2=2.4
r570 37 208 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.595 $Y=1.19
+ $X2=3.595 $Y2=1.355
r571 37 39 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.595 $Y=1.19
+ $X2=3.595 $Y2=0.58
r572 33 207 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.22 $Y=1.52
+ $X2=3.22 $Y2=1.355
r573 33 35 342.065 $w=1.8e-07 $l=8.8e-07 $layer=POLY_cond $X=3.22 $Y=1.52
+ $X2=3.22 $Y2=2.4
r574 29 206 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=1.19
+ $X2=3.165 $Y2=1.355
r575 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.165 $Y=1.19
+ $X2=3.165 $Y2=0.58
r576 25 202 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.52
+ $X2=2.77 $Y2=1.355
r577 25 27 342.065 $w=1.8e-07 $l=8.8e-07 $layer=POLY_cond $X=2.77 $Y=1.52
+ $X2=2.77 $Y2=2.4
r578 21 201 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.735 $Y=1.19
+ $X2=2.735 $Y2=1.355
r579 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.735 $Y=1.19
+ $X2=2.735 $Y2=0.58
r580 17 200 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.32 $Y=1.52
+ $X2=2.32 $Y2=1.355
r581 17 19 342.065 $w=1.8e-07 $l=8.8e-07 $layer=POLY_cond $X=2.32 $Y=1.52
+ $X2=2.32 $Y2=2.4
r582 13 198 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=1.19
+ $X2=2.305 $Y2=1.355
r583 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.305 $Y=1.19
+ $X2=2.305 $Y2=0.58
r584 4 169 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.84 $X2=1.635 $Y2=2.115
r585 4 159 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.84 $X2=1.635 $Y2=2.815
r586 3 166 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.84 $X2=0.735 $Y2=2.115
r587 3 147 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.84 $X2=0.735 $Y2=2.815
r588 2 155 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.45
+ $Y=0.37 $X2=1.59 $Y2=0.58
r589 1 143 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__CLKBUF_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 34 36 42 46
+ 50 56 62 68 72 76 82 88 92 94 99 100 102 103 105 106 108 109 110 111 112 118
+ 135 140 145 154 157 160 163 167
r192 166 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r193 163 164 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r194 160 161 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r195 157 158 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r196 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r197 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r198 149 167 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r199 149 164 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r200 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r201 146 163 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.56 $Y=3.33
+ $X2=8.395 $Y2=3.33
r202 146 148 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.56 $Y=3.33
+ $X2=8.88 $Y2=3.33
r203 145 166 4.72267 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=9.15 $Y=3.33
+ $X2=9.375 $Y2=3.33
r204 145 148 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.15 $Y=3.33
+ $X2=8.88 $Y2=3.33
r205 144 164 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r206 144 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r207 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r208 141 160 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.66 $Y=3.33
+ $X2=7.495 $Y2=3.33
r209 141 143 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.66 $Y=3.33
+ $X2=7.92 $Y2=3.33
r210 140 163 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.23 $Y=3.33
+ $X2=8.395 $Y2=3.33
r211 140 143 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=8.23 $Y=3.33
+ $X2=7.92 $Y2=3.33
r212 139 161 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r213 139 158 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r214 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r215 136 157 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.76 $Y=3.33
+ $X2=6.595 $Y2=3.33
r216 136 138 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=6.76 $Y=3.33
+ $X2=6.96 $Y2=3.33
r217 135 160 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.33 $Y=3.33
+ $X2=7.495 $Y2=3.33
r218 135 138 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.33 $Y=3.33
+ $X2=6.96 $Y2=3.33
r219 134 158 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r220 133 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r221 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r222 128 131 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r223 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r224 125 128 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r225 125 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r226 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r227 122 154 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.25 $Y=3.33
+ $X2=2.125 $Y2=3.33
r228 122 124 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.25 $Y=3.33
+ $X2=2.64 $Y2=3.33
r229 121 155 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r230 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r231 118 154 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2 $Y=3.33
+ $X2=2.125 $Y2=3.33
r232 118 120 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2 $Y=3.33 $X2=1.68
+ $Y2=3.33
r233 117 121 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r234 117 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r235 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r236 114 151 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.37 $Y=3.33
+ $X2=0.185 $Y2=3.33
r237 114 116 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.37 $Y=3.33
+ $X2=0.72 $Y2=3.33
r238 112 134 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=5.52 $Y2=3.33
r239 112 131 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=4.56 $Y2=3.33
r240 110 133 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=5.53 $Y=3.33
+ $X2=5.52 $Y2=3.33
r241 110 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.53 $Y=3.33
+ $X2=5.695 $Y2=3.33
r242 108 130 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=4.63 $Y=3.33
+ $X2=4.56 $Y2=3.33
r243 108 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.63 $Y=3.33
+ $X2=4.795 $Y2=3.33
r244 107 133 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.96 $Y=3.33
+ $X2=5.52 $Y2=3.33
r245 107 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.96 $Y=3.33
+ $X2=4.795 $Y2=3.33
r246 105 127 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.73 $Y=3.33
+ $X2=3.6 $Y2=3.33
r247 105 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.73 $Y=3.33
+ $X2=3.895 $Y2=3.33
r248 104 130 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=4.06 $Y=3.33
+ $X2=4.56 $Y2=3.33
r249 104 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.06 $Y=3.33
+ $X2=3.895 $Y2=3.33
r250 102 124 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.83 $Y=3.33
+ $X2=2.64 $Y2=3.33
r251 102 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.83 $Y=3.33
+ $X2=2.995 $Y2=3.33
r252 101 127 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r253 101 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.16 $Y=3.33
+ $X2=2.995 $Y2=3.33
r254 99 116 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.1 $Y=3.33
+ $X2=0.72 $Y2=3.33
r255 99 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=3.33
+ $X2=1.185 $Y2=3.33
r256 98 120 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.27 $Y=3.33
+ $X2=1.68 $Y2=3.33
r257 98 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=3.33
+ $X2=1.185 $Y2=3.33
r258 94 97 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=9.315 $Y=2.115
+ $X2=9.315 $Y2=2.815
r259 92 166 3.0435 $w=3.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=9.315 $Y=3.245
+ $X2=9.375 $Y2=3.33
r260 92 97 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=9.315 $Y=3.245
+ $X2=9.315 $Y2=2.815
r261 88 91 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=8.395 $Y=2.115
+ $X2=8.395 $Y2=2.815
r262 86 163 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.395 $Y=3.245
+ $X2=8.395 $Y2=3.33
r263 86 91 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.395 $Y=3.245
+ $X2=8.395 $Y2=2.815
r264 82 85 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=7.495 $Y=2.115
+ $X2=7.495 $Y2=2.815
r265 80 160 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.495 $Y=3.245
+ $X2=7.495 $Y2=3.33
r266 80 85 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.495 $Y=3.245
+ $X2=7.495 $Y2=2.815
r267 76 79 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=6.595 $Y=2.115
+ $X2=6.595 $Y2=2.815
r268 74 157 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.595 $Y=3.245
+ $X2=6.595 $Y2=3.33
r269 74 79 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.595 $Y=3.245
+ $X2=6.595 $Y2=2.815
r270 73 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.86 $Y=3.33
+ $X2=5.695 $Y2=3.33
r271 72 157 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.43 $Y=3.33
+ $X2=6.595 $Y2=3.33
r272 72 73 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=6.43 $Y=3.33
+ $X2=5.86 $Y2=3.33
r273 68 71 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=5.695 $Y=2.115
+ $X2=5.695 $Y2=2.815
r274 66 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.695 $Y=3.245
+ $X2=5.695 $Y2=3.33
r275 66 71 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.695 $Y=3.245
+ $X2=5.695 $Y2=2.815
r276 62 65 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=4.795 $Y=2.115
+ $X2=4.795 $Y2=2.815
r277 60 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.795 $Y=3.245
+ $X2=4.795 $Y2=3.33
r278 60 65 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.795 $Y=3.245
+ $X2=4.795 $Y2=2.815
r279 56 59 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=3.895 $Y=2.115
+ $X2=3.895 $Y2=2.815
r280 54 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.895 $Y=3.245
+ $X2=3.895 $Y2=3.33
r281 54 59 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.895 $Y=3.245
+ $X2=3.895 $Y2=2.815
r282 50 53 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=2.995 $Y=2.115
+ $X2=2.995 $Y2=2.815
r283 48 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=3.245
+ $X2=2.995 $Y2=3.33
r284 48 53 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.995 $Y=3.245
+ $X2=2.995 $Y2=2.815
r285 44 154 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.125 $Y=3.245
+ $X2=2.125 $Y2=3.33
r286 44 46 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=2.125 $Y=3.245
+ $X2=2.125 $Y2=2.455
r287 40 100 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=3.245
+ $X2=1.185 $Y2=3.33
r288 40 42 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.185 $Y=3.245
+ $X2=1.185 $Y2=2.455
r289 36 39 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=0.245 $Y=2.115
+ $X2=0.245 $Y2=2.815
r290 34 151 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.245 $Y=3.245
+ $X2=0.185 $Y2=3.33
r291 34 39 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.245 $Y=3.245
+ $X2=0.245 $Y2=2.815
r292 11 97 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.18
+ $Y=1.84 $X2=9.315 $Y2=2.815
r293 11 94 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=9.18
+ $Y=1.84 $X2=9.315 $Y2=2.115
r294 10 91 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.26
+ $Y=1.84 $X2=8.395 $Y2=2.815
r295 10 88 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=8.26
+ $Y=1.84 $X2=8.395 $Y2=2.115
r296 9 85 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.36
+ $Y=1.84 $X2=7.495 $Y2=2.815
r297 9 82 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=7.36
+ $Y=1.84 $X2=7.495 $Y2=2.115
r298 8 79 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.46
+ $Y=1.84 $X2=6.595 $Y2=2.815
r299 8 76 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=6.46
+ $Y=1.84 $X2=6.595 $Y2=2.115
r300 7 71 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.56
+ $Y=1.84 $X2=5.695 $Y2=2.815
r301 7 68 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=5.56
+ $Y=1.84 $X2=5.695 $Y2=2.115
r302 6 65 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.66
+ $Y=1.84 $X2=4.795 $Y2=2.815
r303 6 62 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=4.66
+ $Y=1.84 $X2=4.795 $Y2=2.115
r304 5 59 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.76
+ $Y=1.84 $X2=3.895 $Y2=2.815
r305 5 56 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=3.76
+ $Y=1.84 $X2=3.895 $Y2=2.115
r306 4 53 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.86
+ $Y=1.84 $X2=2.995 $Y2=2.815
r307 4 50 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.86
+ $Y=1.84 $X2=2.995 $Y2=2.115
r308 3 46 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.95
+ $Y=1.84 $X2=2.085 $Y2=2.455
r309 2 42 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.05
+ $Y=1.84 $X2=1.185 $Y2=2.455
r310 1 39 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.815
r311 1 36 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.84 $X2=0.285 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__CLKBUF_16%X 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 51 55 59 65 69 73 77 79 81 85 87 91 92 95 98 101 104 106 109 116 123 130 137
+ 144 151 153 161
c252 153 0 1.65784e-19 $X=8.865 $Y=2.035
r253 158 161 6.04804 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.525 $Y=1.985
+ $X2=2.525 $Y2=2.12
r254 158 160 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.545 $Y=2.035
+ $X2=2.545 $Y2=2.035
r255 151 155 43.4785 $w=2.18e-07 $l=8.3e-07 $layer=LI1_cond $X=8.86 $Y=1.985
+ $X2=8.86 $Y2=2.815
r256 151 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.865 $Y=2.035
+ $X2=8.865 $Y2=2.035
r257 146 153 0.590276 $w=2.3e-07 $l=9.2e-07 $layer=MET1_cond $X=7.945 $Y=2.035
+ $X2=8.865 $Y2=2.035
r258 144 148 43.8355 $w=2.08e-07 $l=8.3e-07 $layer=LI1_cond $X=7.945 $Y=1.985
+ $X2=7.945 $Y2=2.815
r259 144 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.945 $Y=2.035
+ $X2=7.945 $Y2=2.035
r260 139 146 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=7.045 $Y=2.035
+ $X2=7.945 $Y2=2.035
r261 137 141 44.9047 $w=2.03e-07 $l=8.3e-07 $layer=LI1_cond $X=7.047 $Y=1.985
+ $X2=7.047 $Y2=2.815
r262 137 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.045 $Y=2.035
+ $X2=7.045 $Y2=2.035
r263 132 139 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=6.145 $Y=2.035
+ $X2=7.045 $Y2=2.035
r264 130 134 44.9047 $w=2.03e-07 $l=8.3e-07 $layer=LI1_cond $X=6.142 $Y=1.985
+ $X2=6.142 $Y2=2.815
r265 130 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.145 $Y=2.035
+ $X2=6.145 $Y2=2.035
r266 123 127 43.8355 $w=2.08e-07 $l=8.3e-07 $layer=LI1_cond $X=5.245 $Y=1.985
+ $X2=5.245 $Y2=2.815
r267 123 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.245 $Y=2.035
+ $X2=5.245 $Y2=2.035
r268 118 125 0.587068 $w=2.3e-07 $l=9.15e-07 $layer=MET1_cond $X=4.33 $Y=2.035
+ $X2=5.245 $Y2=2.035
r269 116 120 46.0273 $w=1.98e-07 $l=8.3e-07 $layer=LI1_cond $X=4.33 $Y=1.985
+ $X2=4.33 $Y2=2.815
r270 116 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.33 $Y=2.035
+ $X2=4.33 $Y2=2.035
r271 111 118 0.56782 $w=2.3e-07 $l=8.85e-07 $layer=MET1_cond $X=3.445 $Y=2.035
+ $X2=4.33 $Y2=2.035
r272 111 160 0.577444 $w=2.3e-07 $l=9e-07 $layer=MET1_cond $X=3.445 $Y=2.035
+ $X2=2.545 $Y2=2.035
r273 109 113 44.9047 $w=2.03e-07 $l=8.3e-07 $layer=LI1_cond $X=3.442 $Y=1.985
+ $X2=3.442 $Y2=2.815
r274 109 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.445 $Y=2.035
+ $X2=3.445 $Y2=2.035
r275 106 132 0.25985 $w=2.3e-07 $l=4.05e-07 $layer=MET1_cond $X=5.74 $Y=2.035
+ $X2=6.145 $Y2=2.035
r276 106 125 0.317594 $w=2.3e-07 $l=4.95e-07 $layer=MET1_cond $X=5.74 $Y=2.035
+ $X2=5.245 $Y2=2.035
r277 105 151 6.54797 $w=2.18e-07 $l=1.25e-07 $layer=LI1_cond $X=8.86 $Y=1.86
+ $X2=8.86 $Y2=1.985
r278 104 144 6.60173 $w=2.08e-07 $l=1.25e-07 $layer=LI1_cond $X=7.945 $Y=1.86
+ $X2=7.945 $Y2=1.985
r279 103 104 8.16535 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=7.922 $Y=1.69
+ $X2=7.922 $Y2=1.86
r280 101 137 6.76275 $w=2.03e-07 $l=1.25e-07 $layer=LI1_cond $X=7.047 $Y=1.86
+ $X2=7.047 $Y2=1.985
r281 100 101 8.24408 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=7.007 $Y=1.69
+ $X2=7.007 $Y2=1.86
r282 98 130 6.76275 $w=2.03e-07 $l=1.25e-07 $layer=LI1_cond $X=6.142 $Y=1.86
+ $X2=6.142 $Y2=1.985
r283 97 98 8.24408 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=6.09 $Y=1.69
+ $X2=6.09 $Y2=1.86
r284 95 123 6.60173 $w=2.08e-07 $l=1.25e-07 $layer=LI1_cond $X=5.245 $Y=1.86
+ $X2=5.245 $Y2=1.985
r285 94 95 8.62714 $w=2.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.187 $Y=1.69
+ $X2=5.187 $Y2=1.86
r286 92 116 6.93182 $w=1.98e-07 $l=1.25e-07 $layer=LI1_cond $X=4.33 $Y=1.86
+ $X2=4.33 $Y2=1.985
r287 91 92 9.70862 $w=1.98e-07 $l=1.7e-07 $layer=LI1_cond $X=4.3 $Y=1.69 $X2=4.3
+ $Y2=1.86
r288 89 91 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=4.255 $Y=0.745
+ $X2=4.255 $Y2=1.69
r289 87 89 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=4.207 $Y=0.58
+ $X2=4.207 $Y2=0.745
r290 85 109 6.76275 $w=2.03e-07 $l=1.25e-07 $layer=LI1_cond $X=3.442 $Y=1.86
+ $X2=3.442 $Y2=1.985
r291 84 85 8.82084 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=3.41 $Y=1.69
+ $X2=3.41 $Y2=1.86
r292 79 105 7.59438 $w=2.49e-07 $l=1.59922e-07 $layer=LI1_cond $X=8.85 $Y=1.705
+ $X2=8.86 $Y2=1.86
r293 79 81 51.8599 $w=2.48e-07 $l=1.125e-06 $layer=LI1_cond $X=8.85 $Y=1.705
+ $X2=8.85 $Y2=0.58
r294 77 103 51.1685 $w=2.48e-07 $l=1.11e-06 $layer=LI1_cond $X=7.92 $Y=0.58
+ $X2=7.92 $Y2=1.69
r295 73 100 51.1685 $w=2.48e-07 $l=1.11e-06 $layer=LI1_cond $X=6.99 $Y=0.58
+ $X2=6.99 $Y2=1.69
r296 69 97 51.1685 $w=2.48e-07 $l=1.11e-06 $layer=LI1_cond $X=6.06 $Y=0.58
+ $X2=6.06 $Y2=1.69
r297 65 94 55.6179 $w=2.28e-07 $l=1.11e-06 $layer=LI1_cond $X=5.14 $Y=0.58
+ $X2=5.14 $Y2=1.69
r298 59 84 56.8539 $w=2.23e-07 $l=1.11e-06 $layer=LI1_cond $X=3.387 $Y=0.58
+ $X2=3.387 $Y2=1.69
r299 55 161 14.0297 $w=2.28e-07 $l=2.8e-07 $layer=LI1_cond $X=2.545 $Y=2.4
+ $X2=2.545 $Y2=2.12
r300 51 158 59.9697 $w=2.68e-07 $l=1.405e-06 $layer=LI1_cond $X=2.525 $Y=0.58
+ $X2=2.525 $Y2=1.985
r301 16 155 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.73
+ $Y=1.84 $X2=8.865 $Y2=2.815
r302 16 151 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.73
+ $Y=1.84 $X2=8.865 $Y2=1.985
r303 15 148 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=7.81
+ $Y=1.84 $X2=7.945 $Y2=2.815
r304 15 144 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.81
+ $Y=1.84 $X2=7.945 $Y2=1.985
r305 14 141 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.91
+ $Y=1.84 $X2=7.045 $Y2=2.815
r306 14 137 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.91
+ $Y=1.84 $X2=7.045 $Y2=1.985
r307 13 134 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.01
+ $Y=1.84 $X2=6.145 $Y2=2.815
r308 13 130 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.01
+ $Y=1.84 $X2=6.145 $Y2=1.985
r309 12 127 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.11
+ $Y=1.84 $X2=5.245 $Y2=2.815
r310 12 123 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.11
+ $Y=1.84 $X2=5.245 $Y2=1.985
r311 11 120 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.21
+ $Y=1.84 $X2=4.345 $Y2=2.815
r312 11 116 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.21
+ $Y=1.84 $X2=4.345 $Y2=1.985
r313 10 113 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.31
+ $Y=1.84 $X2=3.445 $Y2=2.815
r314 10 109 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.31
+ $Y=1.84 $X2=3.445 $Y2=1.985
r315 9 158 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=1.84 $X2=2.545 $Y2=1.985
r316 9 55 300 $w=1.7e-07 $l=6.23859e-07 $layer=licon1_PDIFF $count=2 $X=2.41
+ $Y=1.84 $X2=2.545 $Y2=2.4
r317 8 81 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.75
+ $Y=0.37 $X2=8.89 $Y2=0.58
r318 7 77 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.82
+ $Y=0.37 $X2=7.96 $Y2=0.58
r319 6 73 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.89
+ $Y=0.37 $X2=7.03 $Y2=0.58
r320 5 69 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.96
+ $Y=0.37 $X2=6.1 $Y2=0.58
r321 4 65 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.03
+ $Y=0.37 $X2=5.17 $Y2=0.58
r322 3 87 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.1
+ $Y=0.37 $X2=4.24 $Y2=0.58
r323 2 59 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.24
+ $Y=0.37 $X2=3.38 $Y2=0.58
r324 1 51 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.37 $X2=2.52 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__CLKBUF_16%VGND 1 2 3 4 5 6 7 8 9 10 11 34 36 40 44
+ 48 52 54 58 62 66 70 74 76 78 81 82 84 85 87 88 89 90 91 106 111 116 121 126
+ 135 138 141 144 147 151
r167 150 151 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r168 147 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r169 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r170 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r171 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r172 135 136 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r173 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r174 130 151 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r175 130 148 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=8.4 $Y2=0
r176 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r177 127 147 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.555 $Y=0
+ $X2=8.39 $Y2=0
r178 127 129 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.555 $Y=0
+ $X2=8.88 $Y2=0
r179 126 150 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=9.155 $Y=0
+ $X2=9.377 $Y2=0
r180 126 129 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=9.155 $Y=0
+ $X2=8.88 $Y2=0
r181 125 148 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=8.4 $Y2=0
r182 125 145 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r183 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r184 122 144 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.625 $Y=0
+ $X2=7.46 $Y2=0
r185 122 124 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.625 $Y=0
+ $X2=7.92 $Y2=0
r186 121 147 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.225 $Y=0
+ $X2=8.39 $Y2=0
r187 121 124 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.225 $Y=0
+ $X2=7.92 $Y2=0
r188 120 145 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r189 120 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=6.48 $Y2=0
r190 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r191 117 141 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.695 $Y=0
+ $X2=6.53 $Y2=0
r192 117 119 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.695 $Y=0
+ $X2=6.96 $Y2=0
r193 116 144 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.295 $Y=0
+ $X2=7.46 $Y2=0
r194 116 119 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.295 $Y=0
+ $X2=6.96 $Y2=0
r195 115 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r196 115 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r197 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6
+ $Y2=0
r198 112 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.765 $Y=0
+ $X2=5.6 $Y2=0
r199 112 114 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.765 $Y=0 $X2=6
+ $Y2=0
r200 111 141 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.365 $Y=0
+ $X2=6.53 $Y2=0
r201 111 114 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.365 $Y=0 $X2=6
+ $Y2=0
r202 110 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r203 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r204 107 135 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=4.835 $Y=0
+ $X2=4.672 $Y2=0
r205 107 109 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.835 $Y=0
+ $X2=5.04 $Y2=0
r206 106 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.435 $Y=0
+ $X2=5.6 $Y2=0
r207 106 109 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.435 $Y=0
+ $X2=5.04 $Y2=0
r208 105 136 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0
+ $X2=4.56 $Y2=0
r209 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r210 102 105 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.6 $Y2=0
r211 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r212 99 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.64 $Y2=0
r213 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r214 96 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r215 96 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r216 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r217 93 132 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r218 93 95 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.72 $Y2=0
r219 91 110 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0
+ $X2=5.04 $Y2=0
r220 91 136 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0
+ $X2=4.56 $Y2=0
r221 89 104 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.67 $Y=0 $X2=3.6
+ $Y2=0
r222 89 90 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=3.67 $Y=0 $X2=3.782
+ $Y2=0
r223 87 101 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.865 $Y=0
+ $X2=2.64 $Y2=0
r224 87 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.95
+ $Y2=0
r225 86 104 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.035 $Y=0 $X2=3.6
+ $Y2=0
r226 86 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.035 $Y=0 $X2=2.95
+ $Y2=0
r227 84 98 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.855 $Y=0
+ $X2=1.68 $Y2=0
r228 84 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=2.02
+ $Y2=0
r229 83 101 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=2.185 $Y=0
+ $X2=2.64 $Y2=0
r230 83 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.185 $Y=0 $X2=2.02
+ $Y2=0
r231 81 95 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0
+ $X2=0.72 $Y2=0
r232 81 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.1
+ $Y2=0
r233 80 98 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.225 $Y=0
+ $X2=1.68 $Y2=0
r234 80 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.1
+ $Y2=0
r235 76 150 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=9.32 $Y=0.085
+ $X2=9.377 $Y2=0
r236 76 78 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=9.32 $Y=0.085
+ $X2=9.32 $Y2=0.58
r237 72 147 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.39 $Y=0.085
+ $X2=8.39 $Y2=0
r238 72 74 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.39 $Y=0.085
+ $X2=8.39 $Y2=0.515
r239 68 144 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.46 $Y=0.085
+ $X2=7.46 $Y2=0
r240 68 70 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.46 $Y=0.085
+ $X2=7.46 $Y2=0.515
r241 64 141 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.53 $Y=0.085
+ $X2=6.53 $Y2=0
r242 64 66 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.53 $Y=0.085
+ $X2=6.53 $Y2=0.515
r243 60 138 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.6 $Y=0.085
+ $X2=5.6 $Y2=0
r244 60 62 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.6 $Y=0.085
+ $X2=5.6 $Y2=0.515
r245 56 135 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=4.672 $Y=0.085
+ $X2=4.672 $Y2=0
r246 56 58 17.3753 $w=3.23e-07 $l=4.9e-07 $layer=LI1_cond $X=4.672 $Y=0.085
+ $X2=4.672 $Y2=0.575
r247 55 90 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=3.895 $Y=0
+ $X2=3.782 $Y2=0
r248 54 135 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=4.51 $Y=0 $X2=4.672
+ $Y2=0
r249 54 55 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.51 $Y=0 $X2=3.895
+ $Y2=0
r250 50 90 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=3.782 $Y=0.085
+ $X2=3.782 $Y2=0
r251 50 52 24.3294 $w=2.23e-07 $l=4.75e-07 $layer=LI1_cond $X=3.782 $Y=0.085
+ $X2=3.782 $Y2=0.56
r252 46 88 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.95 $Y=0.085
+ $X2=2.95 $Y2=0
r253 46 48 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=2.95 $Y=0.085
+ $X2=2.95 $Y2=0.515
r254 42 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0
r255 42 44 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0.58
r256 38 82 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0
r257 38 40 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.58
r258 34 132 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r259 34 36 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.58
r260 11 78 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.18
+ $Y=0.37 $X2=9.32 $Y2=0.58
r261 10 74 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=8.25
+ $Y=0.37 $X2=8.39 $Y2=0.515
r262 9 70 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.32
+ $Y=0.37 $X2=7.46 $Y2=0.515
r263 8 66 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.39
+ $Y=0.37 $X2=6.53 $Y2=0.515
r264 7 62 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.46
+ $Y=0.37 $X2=5.6 $Y2=0.515
r265 6 58 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=4.53
+ $Y=0.37 $X2=4.67 $Y2=0.575
r266 5 52 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=3.67
+ $Y=0.37 $X2=3.81 $Y2=0.56
r267 4 48 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.81
+ $Y=0.37 $X2=2.95 $Y2=0.515
r268 3 44 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.88
+ $Y=0.37 $X2=2.02 $Y2=0.58
r269 2 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.37 $X2=1.14 $Y2=0.58
r270 1 36 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdlclkp_2 CLK GATE SCE VGND VNB VPB VPWR GCLK
M1000 a_706_317# a_580_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=2.04535e+12p ps=1.691e+07u
M1001 GCLK a_1198_374# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1002 VGND CLK a_288_48# VNB nlowvt w=740000u l=150000u
+  ad=1.5071e+12p pd=1.328e+07u as=2.109e+11p ps=2.05e+06u
M1003 VPWR a_1198_374# GCLK VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_706_317# a_580_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1005 a_580_74# a_318_74# a_114_112# VPB pshort w=840000u l=180000u
+  ad=2.583e+11p pd=2.37e+06u as=4.536e+11p ps=4.44e+06u
M1006 a_318_74# a_288_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1007 VPWR a_706_317# a_711_451# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1008 a_114_112# GATE a_117_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=1.764e+11p ps=2.1e+06u
M1009 GCLK a_1198_374# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1010 VPWR CLK a_288_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.268e+11p ps=2.22e+06u
M1011 a_1198_374# a_706_317# a_1198_74# VNB nlowvt w=740000u l=150000u
+  ad=2.035e+11p pd=2.03e+06u as=1.554e+11p ps=1.9e+06u
M1012 a_318_74# a_288_48# VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1013 a_711_451# a_288_48# a_580_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND GATE a_114_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=4.8675e+11p ps=3.97e+06u
M1015 a_114_112# SCE VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1198_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_1198_374# GCLK VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_685_81# a_318_74# a_580_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.9475e+11p ps=1.85e+06u
M1019 VGND a_706_317# a_685_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_706_317# a_1198_374# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=4.85e+11p ps=2.97e+06u
M1021 a_1198_374# CLK VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_117_424# SCE VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_580_74# a_288_48# a_114_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_ms__a41o_1.pxi.spice
* Created: Fri Aug 28 17:09:04 2020
* 
x_PM_SKY130_FD_SC_MS__A41O_1%A_83_244# N_A_83_244#_M1008_d N_A_83_244#_M1010_s
+ N_A_83_244#_M1001_g N_A_83_244#_c_73_n N_A_83_244#_M1005_g N_A_83_244#_c_74_n
+ N_A_83_244#_c_75_n N_A_83_244#_c_76_n N_A_83_244#_c_82_n N_A_83_244#_c_77_n
+ N_A_83_244#_c_78_n N_A_83_244#_c_79_n N_A_83_244#_c_83_n N_A_83_244#_c_80_n
+ PM_SKY130_FD_SC_MS__A41O_1%A_83_244#
x_PM_SKY130_FD_SC_MS__A41O_1%B1 N_B1_M1010_g N_B1_M1008_g B1 N_B1_c_137_n
+ PM_SKY130_FD_SC_MS__A41O_1%B1
x_PM_SKY130_FD_SC_MS__A41O_1%A1 N_A1_M1003_g N_A1_M1011_g A1 N_A1_c_171_n
+ PM_SKY130_FD_SC_MS__A41O_1%A1
x_PM_SKY130_FD_SC_MS__A41O_1%A2 N_A2_M1000_g N_A2_M1002_g A2 A2 A2 N_A2_c_210_n
+ N_A2_c_211_n PM_SKY130_FD_SC_MS__A41O_1%A2
x_PM_SKY130_FD_SC_MS__A41O_1%A3 N_A3_M1006_g N_A3_M1004_g A3 N_A3_c_248_n
+ N_A3_c_249_n PM_SKY130_FD_SC_MS__A41O_1%A3
x_PM_SKY130_FD_SC_MS__A41O_1%A4 N_A4_c_278_n N_A4_M1009_g N_A4_M1007_g A4
+ N_A4_c_281_n PM_SKY130_FD_SC_MS__A41O_1%A4
x_PM_SKY130_FD_SC_MS__A41O_1%X N_X_M1005_s N_X_M1001_s N_X_c_303_n N_X_c_306_n
+ N_X_c_307_n N_X_c_304_n N_X_c_305_n X PM_SKY130_FD_SC_MS__A41O_1%X
x_PM_SKY130_FD_SC_MS__A41O_1%VPWR N_VPWR_M1001_d N_VPWR_M1011_d N_VPWR_M1004_d
+ N_VPWR_c_325_n N_VPWR_c_326_n N_VPWR_c_327_n N_VPWR_c_328_n N_VPWR_c_329_n
+ N_VPWR_c_330_n N_VPWR_c_331_n VPWR N_VPWR_c_332_n N_VPWR_c_324_n
+ N_VPWR_c_334_n PM_SKY130_FD_SC_MS__A41O_1%VPWR
x_PM_SKY130_FD_SC_MS__A41O_1%A_357_392# N_A_357_392#_M1010_d
+ N_A_357_392#_M1002_d N_A_357_392#_M1007_d N_A_357_392#_c_373_n
+ N_A_357_392#_c_374_n N_A_357_392#_c_375_n N_A_357_392#_c_376_n
+ N_A_357_392#_c_377_n N_A_357_392#_c_378_n N_A_357_392#_c_379_n
+ PM_SKY130_FD_SC_MS__A41O_1%A_357_392#
x_PM_SKY130_FD_SC_MS__A41O_1%VGND N_VGND_M1005_d N_VGND_M1009_d N_VGND_c_426_n
+ N_VGND_c_427_n N_VGND_c_428_n N_VGND_c_429_n N_VGND_c_430_n VGND
+ N_VGND_c_431_n N_VGND_c_432_n PM_SKY130_FD_SC_MS__A41O_1%VGND
cc_1 VNB N_A_83_244#_M1001_g 0.00769232f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_2 VNB N_A_83_244#_c_73_n 0.0215513f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.22
cc_3 VNB N_A_83_244#_c_74_n 0.0196302f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.385
cc_4 VNB N_A_83_244#_c_75_n 0.0670264f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.385
cc_5 VNB N_A_83_244#_c_76_n 0.00597917f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.33
cc_6 VNB N_A_83_244#_c_77_n 0.0124475f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.195
cc_7 VNB N_A_83_244#_c_78_n 0.00240191f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=0.515
cc_8 VNB N_A_83_244#_c_79_n 0.00286203f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.33
cc_9 VNB N_A_83_244#_c_80_n 0.00211666f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=1.95
cc_10 VNB N_B1_M1008_g 0.0304701f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.55
cc_11 VNB B1 0.00166024f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_12 VNB N_B1_c_137_n 0.0203932f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=0.74
cc_13 VNB N_A1_M1003_g 0.0299791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB A1 0.004704f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_15 VNB N_A1_c_171_n 0.0199513f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=0.74
cc_16 VNB N_A2_M1002_g 0.00642364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB A2 0.00751257f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_18 VNB N_A2_c_210_n 0.0312348f $X=-0.19 $Y=-0.245 $X2=1.095 $Y2=1.385
cc_19 VNB N_A2_c_211_n 0.0182251f $X=-0.19 $Y=-0.245 $X2=1.08 $Y2=1.33
cc_20 VNB N_A3_M1004_g 0.00667073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB A3 0.0207403f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_22 VNB N_A3_c_248_n 0.0279589f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.22
cc_23 VNB N_A3_c_249_n 0.0198625f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=0.74
cc_24 VNB N_A4_c_278_n 0.0220567f $X=-0.19 $Y=-0.245 $X2=1.815 $Y2=0.37
cc_25 VNB N_A4_M1007_g 0.00984151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB A4 0.0102f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_27 VNB N_A4_c_281_n 0.0588392f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.385
cc_28 VNB N_X_c_303_n 0.029462f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.55
cc_29 VNB N_X_c_304_n 0.00735758f $X=-0.19 $Y=-0.245 $X2=1.08 $Y2=1.33
cc_30 VNB N_X_c_305_n 0.0348735f $X=-0.19 $Y=-0.245 $X2=1.08 $Y2=1.385
cc_31 VNB N_VPWR_c_324_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_426_n 0.00944368f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.4
cc_33 VNB N_VGND_c_427_n 0.0134627f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.22
cc_34 VNB N_VGND_c_428_n 0.0344105f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=0.74
cc_35 VNB N_VGND_c_429_n 0.0343772f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.33
cc_36 VNB N_VGND_c_430_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.08 $Y2=1.33
cc_37 VNB N_VGND_c_431_n 0.0651336f $X=-0.19 $Y=-0.245 $X2=1.79 $Y2=1.195
cc_38 VNB N_VGND_c_432_n 0.284384f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=1.95
cc_39 VPB N_A_83_244#_M1001_g 0.0298763f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_40 VPB N_A_83_244#_c_82_n 0.015876f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=2.815
cc_41 VPB N_A_83_244#_c_83_n 0.00702741f $X=-0.19 $Y=1.66 $X2=1.47 $Y2=2.115
cc_42 VPB N_A_83_244#_c_80_n 0.00702583f $X=-0.19 $Y=1.66 $X2=1.39 $Y2=1.95
cc_43 VPB N_B1_M1010_g 0.0285589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB B1 0.0019308f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_45 VPB N_B1_c_137_n 0.0133245f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=0.74
cc_46 VPB N_A1_M1011_g 0.0252615f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.55
cc_47 VPB A1 0.00137127f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.4
cc_48 VPB N_A1_c_171_n 0.0130018f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=0.74
cc_49 VPB N_A2_M1002_g 0.0304432f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A3_M1004_g 0.0296902f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_A4_M1007_g 0.0386398f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_X_c_306_n 0.00878289f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=1.22
cc_53 VPB N_X_c_307_n 0.0403824f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=0.74
cc_54 VPB N_X_c_305_n 0.00790717f $X=-0.19 $Y=1.66 $X2=1.08 $Y2=1.385
cc_55 VPB N_VPWR_c_325_n 0.0269089f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.385
cc_56 VPB N_VPWR_c_326_n 0.00976734f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_327_n 0.00976275f $X=-0.19 $Y=1.66 $X2=1.39 $Y2=2.815
cc_58 VPB N_VPWR_c_328_n 0.0384309f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=1.11
cc_59 VPB N_VPWR_c_329_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=0.515
cc_60 VPB N_VPWR_c_330_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_331_n 0.00632158f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.33
cc_62 VPB N_VPWR_c_332_n 0.0204244f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_324_n 0.077656f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_334_n 0.024889f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_357_392#_c_373_n 0.00426734f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_A_357_392#_c_374_n 0.00275675f $X=-0.19 $Y=1.66 $X2=1.17 $Y2=0.74
cc_67 VPB N_A_357_392#_c_375_n 0.00793717f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.385
cc_68 VPB N_A_357_392#_c_376_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.08 $Y2=1.385
cc_69 VPB N_A_357_392#_c_377_n 0.0178871f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_357_392#_c_378_n 0.0442448f $X=-0.19 $Y=1.66 $X2=1.39 $Y2=2.815
cc_71 VPB N_A_357_392#_c_379_n 0.00999306f $X=-0.19 $Y=1.66 $X2=1.955 $Y2=0.515
cc_72 N_A_83_244#_c_82_n N_B1_M1010_g 0.00954303f $X=1.47 $Y=2.815 $X2=0 $Y2=0
cc_73 N_A_83_244#_c_83_n N_B1_M1010_g 0.00337618f $X=1.47 $Y=2.115 $X2=0 $Y2=0
cc_74 N_A_83_244#_c_80_n N_B1_M1010_g 0.00519584f $X=1.39 $Y=1.95 $X2=0 $Y2=0
cc_75 N_A_83_244#_c_73_n N_B1_M1008_g 0.0269165f $X=1.17 $Y=1.22 $X2=0 $Y2=0
cc_76 N_A_83_244#_c_77_n N_B1_M1008_g 0.014512f $X=1.79 $Y=1.195 $X2=0 $Y2=0
cc_77 N_A_83_244#_c_78_n N_B1_M1008_g 0.0106829f $X=1.955 $Y=0.515 $X2=0 $Y2=0
cc_78 N_A_83_244#_c_79_n N_B1_M1008_g 0.00397456f $X=1.23 $Y=1.33 $X2=0 $Y2=0
cc_79 N_A_83_244#_c_77_n B1 0.0243844f $X=1.79 $Y=1.195 $X2=0 $Y2=0
cc_80 N_A_83_244#_c_79_n B1 0.00843332f $X=1.23 $Y=1.33 $X2=0 $Y2=0
cc_81 N_A_83_244#_c_83_n B1 0.0124116f $X=1.47 $Y=2.115 $X2=0 $Y2=0
cc_82 N_A_83_244#_c_80_n B1 0.0172484f $X=1.39 $Y=1.95 $X2=0 $Y2=0
cc_83 N_A_83_244#_c_75_n N_B1_c_137_n 0.00529013f $X=1.095 $Y=1.385 $X2=0 $Y2=0
cc_84 N_A_83_244#_c_77_n N_B1_c_137_n 0.00125621f $X=1.79 $Y=1.195 $X2=0 $Y2=0
cc_85 N_A_83_244#_c_79_n N_B1_c_137_n 6.53316e-19 $X=1.23 $Y=1.33 $X2=0 $Y2=0
cc_86 N_A_83_244#_c_83_n N_B1_c_137_n 9.41854e-19 $X=1.47 $Y=2.115 $X2=0 $Y2=0
cc_87 N_A_83_244#_c_80_n N_B1_c_137_n 0.00515453f $X=1.39 $Y=1.95 $X2=0 $Y2=0
cc_88 N_A_83_244#_c_77_n N_A1_M1003_g 0.00496732f $X=1.79 $Y=1.195 $X2=0 $Y2=0
cc_89 N_A_83_244#_c_78_n N_A1_M1003_g 0.0131343f $X=1.955 $Y=0.515 $X2=0 $Y2=0
cc_90 N_A_83_244#_c_83_n N_A1_M1011_g 2.55989e-19 $X=1.47 $Y=2.115 $X2=0 $Y2=0
cc_91 N_A_83_244#_c_77_n A1 0.00785342f $X=1.79 $Y=1.195 $X2=0 $Y2=0
cc_92 N_A_83_244#_c_77_n N_A1_c_171_n 5.46117e-19 $X=1.79 $Y=1.195 $X2=0 $Y2=0
cc_93 N_A_83_244#_c_77_n A2 0.00747525f $X=1.79 $Y=1.195 $X2=0 $Y2=0
cc_94 N_A_83_244#_c_78_n N_A2_c_211_n 0.00111606f $X=1.955 $Y=0.515 $X2=0 $Y2=0
cc_95 N_A_83_244#_M1001_g N_X_c_306_n 0.00388688f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_96 N_A_83_244#_M1001_g N_X_c_307_n 0.0141275f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_97 N_A_83_244#_c_73_n N_X_c_304_n 0.00911848f $X=1.17 $Y=1.22 $X2=0 $Y2=0
cc_98 N_A_83_244#_c_74_n N_X_c_304_n 0.00975101f $X=0.595 $Y=1.385 $X2=0 $Y2=0
cc_99 N_A_83_244#_c_76_n N_X_c_304_n 0.045133f $X=1.145 $Y=1.33 $X2=0 $Y2=0
cc_100 N_A_83_244#_c_74_n N_X_c_305_n 0.0212801f $X=0.595 $Y=1.385 $X2=0 $Y2=0
cc_101 N_A_83_244#_c_76_n N_X_c_305_n 0.0300485f $X=1.145 $Y=1.33 $X2=0 $Y2=0
cc_102 N_A_83_244#_M1001_g N_VPWR_c_325_n 0.00649215f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_103 N_A_83_244#_c_75_n N_VPWR_c_325_n 0.00546342f $X=1.095 $Y=1.385 $X2=0
+ $Y2=0
cc_104 N_A_83_244#_c_76_n N_VPWR_c_325_n 0.0151079f $X=1.145 $Y=1.33 $X2=0 $Y2=0
cc_105 N_A_83_244#_c_80_n N_VPWR_c_325_n 0.0738739f $X=1.39 $Y=1.95 $X2=0 $Y2=0
cc_106 N_A_83_244#_c_82_n N_VPWR_c_328_n 0.0216883f $X=1.47 $Y=2.815 $X2=0 $Y2=0
cc_107 N_A_83_244#_M1001_g N_VPWR_c_324_n 0.00991141f $X=0.505 $Y=2.4 $X2=0
+ $Y2=0
cc_108 N_A_83_244#_c_82_n N_VPWR_c_324_n 0.0178836f $X=1.47 $Y=2.815 $X2=0 $Y2=0
cc_109 N_A_83_244#_M1001_g N_VPWR_c_334_n 0.005209f $X=0.505 $Y=2.4 $X2=0 $Y2=0
cc_110 N_A_83_244#_c_77_n N_A_357_392#_c_373_n 0.00756967f $X=1.79 $Y=1.195
+ $X2=0 $Y2=0
cc_111 N_A_83_244#_c_83_n N_A_357_392#_c_373_n 0.0072281f $X=1.47 $Y=2.115 $X2=0
+ $Y2=0
cc_112 N_A_83_244#_c_83_n N_A_357_392#_c_374_n 0.035031f $X=1.47 $Y=2.115 $X2=0
+ $Y2=0
cc_113 N_A_83_244#_c_79_n N_VGND_M1005_d 0.00234067f $X=1.23 $Y=1.33 $X2=-0.19
+ $Y2=-0.245
cc_114 N_A_83_244#_c_73_n N_VGND_c_426_n 0.00566111f $X=1.17 $Y=1.22 $X2=0 $Y2=0
cc_115 N_A_83_244#_c_77_n N_VGND_c_426_n 0.0246062f $X=1.79 $Y=1.195 $X2=0 $Y2=0
cc_116 N_A_83_244#_c_78_n N_VGND_c_426_n 0.0229287f $X=1.955 $Y=0.515 $X2=0
+ $Y2=0
cc_117 N_A_83_244#_c_79_n N_VGND_c_426_n 0.00166799f $X=1.23 $Y=1.33 $X2=0 $Y2=0
cc_118 N_A_83_244#_c_73_n N_VGND_c_429_n 0.00431773f $X=1.17 $Y=1.22 $X2=0 $Y2=0
cc_119 N_A_83_244#_c_78_n N_VGND_c_431_n 0.0144922f $X=1.955 $Y=0.515 $X2=0
+ $Y2=0
cc_120 N_A_83_244#_c_73_n N_VGND_c_432_n 0.00821885f $X=1.17 $Y=1.22 $X2=0 $Y2=0
cc_121 N_A_83_244#_c_78_n N_VGND_c_432_n 0.0118826f $X=1.955 $Y=0.515 $X2=0
+ $Y2=0
cc_122 N_B1_M1008_g N_A1_M1003_g 0.0249499f $X=1.74 $Y=0.74 $X2=0 $Y2=0
cc_123 N_B1_M1010_g N_A1_M1011_g 0.0134153f $X=1.695 $Y=2.46 $X2=0 $Y2=0
cc_124 B1 A1 0.0209133f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_125 N_B1_c_137_n A1 0.00114936f $X=1.65 $Y=1.615 $X2=0 $Y2=0
cc_126 B1 N_A1_c_171_n 0.00114936f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_127 N_B1_c_137_n N_A1_c_171_n 0.0201104f $X=1.65 $Y=1.615 $X2=0 $Y2=0
cc_128 N_B1_M1010_g N_VPWR_c_328_n 0.005209f $X=1.695 $Y=2.46 $X2=0 $Y2=0
cc_129 N_B1_M1010_g N_VPWR_c_324_n 0.00989063f $X=1.695 $Y=2.46 $X2=0 $Y2=0
cc_130 B1 N_A_357_392#_c_373_n 7.62703e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_131 N_B1_M1008_g N_VGND_c_426_n 0.00683336f $X=1.74 $Y=0.74 $X2=0 $Y2=0
cc_132 N_B1_M1008_g N_VGND_c_431_n 0.00434272f $X=1.74 $Y=0.74 $X2=0 $Y2=0
cc_133 N_B1_M1008_g N_VGND_c_432_n 0.0082141f $X=1.74 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A1_M1011_g N_A2_M1002_g 0.0244076f $X=2.195 $Y=2.46 $X2=0 $Y2=0
cc_135 A1 N_A2_M1002_g 0.00127608f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_136 N_A1_c_171_n N_A2_M1002_g 0.00899192f $X=2.19 $Y=1.615 $X2=0 $Y2=0
cc_137 N_A1_M1003_g A2 0.00699457f $X=2.17 $Y=0.74 $X2=0 $Y2=0
cc_138 A1 A2 0.00798656f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_139 N_A1_c_171_n A2 5.70293e-19 $X=2.19 $Y=1.615 $X2=0 $Y2=0
cc_140 N_A1_c_171_n N_A2_c_210_n 0.00625135f $X=2.19 $Y=1.615 $X2=0 $Y2=0
cc_141 N_A1_M1003_g N_A2_c_211_n 0.0435927f $X=2.17 $Y=0.74 $X2=0 $Y2=0
cc_142 N_A1_M1011_g N_VPWR_c_326_n 0.00348921f $X=2.195 $Y=2.46 $X2=0 $Y2=0
cc_143 N_A1_M1011_g N_VPWR_c_328_n 0.005209f $X=2.195 $Y=2.46 $X2=0 $Y2=0
cc_144 N_A1_M1011_g N_VPWR_c_324_n 0.00983375f $X=2.195 $Y=2.46 $X2=0 $Y2=0
cc_145 N_A1_M1011_g N_A_357_392#_c_373_n 0.00100052f $X=2.195 $Y=2.46 $X2=0
+ $Y2=0
cc_146 A1 N_A_357_392#_c_373_n 0.00910208f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_147 N_A1_c_171_n N_A_357_392#_c_373_n 6.24319e-19 $X=2.19 $Y=1.615 $X2=0
+ $Y2=0
cc_148 N_A1_M1011_g N_A_357_392#_c_374_n 0.0119151f $X=2.195 $Y=2.46 $X2=0 $Y2=0
cc_149 N_A1_M1011_g N_A_357_392#_c_375_n 0.0135588f $X=2.195 $Y=2.46 $X2=0 $Y2=0
cc_150 A1 N_A_357_392#_c_375_n 0.0159453f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_151 N_A1_c_171_n N_A_357_392#_c_375_n 4.86414e-19 $X=2.19 $Y=1.615 $X2=0
+ $Y2=0
cc_152 N_A1_M1011_g N_A_357_392#_c_379_n 0.0017003f $X=2.195 $Y=2.46 $X2=0 $Y2=0
cc_153 A1 N_A_357_392#_c_379_n 0.00193532f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_154 N_A1_M1003_g N_VGND_c_431_n 0.00434272f $X=2.17 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A1_M1003_g N_VGND_c_432_n 0.00821825f $X=2.17 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A2_M1002_g N_A3_M1004_g 0.0263975f $X=2.775 $Y=2.46 $X2=0 $Y2=0
cc_157 A2 A3 0.0223103f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_158 N_A2_c_210_n A3 0.00121006f $X=2.73 $Y=1.385 $X2=0 $Y2=0
cc_159 A2 N_A3_c_248_n 4.20157e-19 $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_160 N_A2_c_210_n N_A3_c_248_n 0.017626f $X=2.73 $Y=1.385 $X2=0 $Y2=0
cc_161 A2 N_A3_c_249_n 0.0175036f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_162 N_A2_c_211_n N_A3_c_249_n 0.0251453f $X=2.73 $Y=1.22 $X2=0 $Y2=0
cc_163 N_A2_M1002_g N_VPWR_c_326_n 0.00739211f $X=2.775 $Y=2.46 $X2=0 $Y2=0
cc_164 N_A2_M1002_g N_VPWR_c_330_n 0.005209f $X=2.775 $Y=2.46 $X2=0 $Y2=0
cc_165 N_A2_M1002_g N_VPWR_c_324_n 0.00983591f $X=2.775 $Y=2.46 $X2=0 $Y2=0
cc_166 N_A2_M1002_g N_A_357_392#_c_374_n 9.02211e-19 $X=2.775 $Y=2.46 $X2=0
+ $Y2=0
cc_167 N_A2_M1002_g N_A_357_392#_c_375_n 0.0153614f $X=2.775 $Y=2.46 $X2=0 $Y2=0
cc_168 A2 N_A_357_392#_c_375_n 0.0125729f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_169 N_A2_c_210_n N_A_357_392#_c_375_n 6.9296e-19 $X=2.73 $Y=1.385 $X2=0 $Y2=0
cc_170 N_A2_M1002_g N_A_357_392#_c_376_n 0.0124124f $X=2.775 $Y=2.46 $X2=0 $Y2=0
cc_171 N_A2_M1002_g N_A_357_392#_c_379_n 0.00877821f $X=2.775 $Y=2.46 $X2=0
+ $Y2=0
cc_172 A2 N_A_357_392#_c_379_n 0.00504036f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_173 N_A2_c_210_n N_A_357_392#_c_379_n 2.29527e-19 $X=2.73 $Y=1.385 $X2=0
+ $Y2=0
cc_174 A2 N_VGND_c_431_n 0.00999172f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_175 N_A2_c_211_n N_VGND_c_431_n 0.00303293f $X=2.73 $Y=1.22 $X2=0 $Y2=0
cc_176 A2 N_VGND_c_432_n 0.0120835f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_177 N_A2_c_211_n N_VGND_c_432_n 0.0037339f $X=2.73 $Y=1.22 $X2=0 $Y2=0
cc_178 A2 A_543_74# 0.0106871f $X=2.555 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_179 A3 N_A4_c_278_n 0.00145507f $X=3.515 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_180 N_A3_c_249_n N_A4_c_278_n 0.0301841f $X=3.3 $Y=1.22 $X2=-0.19 $Y2=-0.245
cc_181 N_A3_M1004_g N_A4_M1007_g 0.0276099f $X=3.225 $Y=2.46 $X2=0 $Y2=0
cc_182 A3 A4 0.0291227f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_183 N_A3_c_248_n A4 2.11055e-19 $X=3.3 $Y=1.385 $X2=0 $Y2=0
cc_184 A3 N_A4_c_281_n 0.00860163f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_185 N_A3_c_248_n N_A4_c_281_n 0.0182049f $X=3.3 $Y=1.385 $X2=0 $Y2=0
cc_186 N_A3_M1004_g N_VPWR_c_327_n 0.00347203f $X=3.225 $Y=2.46 $X2=0 $Y2=0
cc_187 N_A3_M1004_g N_VPWR_c_330_n 0.005209f $X=3.225 $Y=2.46 $X2=0 $Y2=0
cc_188 N_A3_M1004_g N_VPWR_c_324_n 0.00982843f $X=3.225 $Y=2.46 $X2=0 $Y2=0
cc_189 N_A3_M1004_g N_A_357_392#_c_376_n 0.0102723f $X=3.225 $Y=2.46 $X2=0 $Y2=0
cc_190 N_A3_M1004_g N_A_357_392#_c_377_n 0.0140921f $X=3.225 $Y=2.46 $X2=0 $Y2=0
cc_191 A3 N_A_357_392#_c_377_n 0.0421079f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_192 N_A3_c_248_n N_A_357_392#_c_377_n 0.00336308f $X=3.3 $Y=1.385 $X2=0 $Y2=0
cc_193 N_A3_M1004_g N_A_357_392#_c_378_n 7.34141e-19 $X=3.225 $Y=2.46 $X2=0
+ $Y2=0
cc_194 N_A3_M1004_g N_A_357_392#_c_379_n 0.00837069f $X=3.225 $Y=2.46 $X2=0
+ $Y2=0
cc_195 A3 N_A_357_392#_c_379_n 0.00233423f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_196 N_A3_c_249_n N_VGND_c_428_n 0.00352277f $X=3.3 $Y=1.22 $X2=0 $Y2=0
cc_197 N_A3_c_249_n N_VGND_c_431_n 0.00461464f $X=3.3 $Y=1.22 $X2=0 $Y2=0
cc_198 N_A3_c_249_n N_VGND_c_432_n 0.00911823f $X=3.3 $Y=1.22 $X2=0 $Y2=0
cc_199 N_A4_M1007_g N_VPWR_c_327_n 0.00879843f $X=3.795 $Y=2.46 $X2=0 $Y2=0
cc_200 N_A4_M1007_g N_VPWR_c_332_n 0.005209f $X=3.795 $Y=2.46 $X2=0 $Y2=0
cc_201 N_A4_M1007_g N_VPWR_c_324_n 0.0098699f $X=3.795 $Y=2.46 $X2=0 $Y2=0
cc_202 N_A4_M1007_g N_A_357_392#_c_377_n 0.0231322f $X=3.795 $Y=2.46 $X2=0 $Y2=0
cc_203 A4 N_A_357_392#_c_377_n 0.0255378f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_204 N_A4_c_281_n N_A_357_392#_c_377_n 0.00236651f $X=4.05 $Y=1.385 $X2=0
+ $Y2=0
cc_205 N_A4_M1007_g N_A_357_392#_c_378_n 0.0164773f $X=3.795 $Y=2.46 $X2=0 $Y2=0
cc_206 N_A4_M1007_g N_A_357_392#_c_379_n 0.00103507f $X=3.795 $Y=2.46 $X2=0
+ $Y2=0
cc_207 N_A4_c_278_n N_VGND_c_428_n 0.0199828f $X=3.78 $Y=1.22 $X2=0 $Y2=0
cc_208 A4 N_VGND_c_428_n 0.0228393f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_209 N_A4_c_281_n N_VGND_c_428_n 0.00186566f $X=4.05 $Y=1.385 $X2=0 $Y2=0
cc_210 N_A4_c_278_n N_VGND_c_431_n 0.00383152f $X=3.78 $Y=1.22 $X2=0 $Y2=0
cc_211 N_A4_c_278_n N_VGND_c_432_n 0.00758792f $X=3.78 $Y=1.22 $X2=0 $Y2=0
cc_212 N_X_c_306_n N_VPWR_c_325_n 0.0395357f $X=0.28 $Y=1.985 $X2=0 $Y2=0
cc_213 N_X_c_307_n N_VPWR_c_324_n 0.0119743f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_214 N_X_c_307_n N_VPWR_c_334_n 0.014549f $X=0.28 $Y=2.815 $X2=0 $Y2=0
cc_215 N_X_c_304_n N_VGND_c_426_n 0.0305553f $X=0.955 $Y=0.515 $X2=0 $Y2=0
cc_216 N_X_c_303_n N_VGND_c_429_n 0.0140792f $X=0.235 $Y=0.94 $X2=0 $Y2=0
cc_217 N_X_c_304_n N_VGND_c_429_n 0.044373f $X=0.955 $Y=0.515 $X2=0 $Y2=0
cc_218 N_X_c_303_n N_VGND_c_432_n 0.00916974f $X=0.235 $Y=0.94 $X2=0 $Y2=0
cc_219 N_X_c_304_n N_VGND_c_432_n 0.0290487f $X=0.955 $Y=0.515 $X2=0 $Y2=0
cc_220 N_VPWR_c_326_n N_A_357_392#_c_374_n 0.0266809f $X=2.47 $Y=2.455 $X2=0
+ $Y2=0
cc_221 N_VPWR_c_328_n N_A_357_392#_c_374_n 0.014549f $X=2.305 $Y=3.33 $X2=0
+ $Y2=0
cc_222 N_VPWR_c_324_n N_A_357_392#_c_374_n 0.0119743f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_223 N_VPWR_M1011_d N_A_357_392#_c_375_n 0.00339226f $X=2.285 $Y=1.96 $X2=0
+ $Y2=0
cc_224 N_VPWR_c_326_n N_A_357_392#_c_375_n 0.0232685f $X=2.47 $Y=2.455 $X2=0
+ $Y2=0
cc_225 N_VPWR_c_326_n N_A_357_392#_c_376_n 0.0234373f $X=2.47 $Y=2.455 $X2=0
+ $Y2=0
cc_226 N_VPWR_c_330_n N_A_357_392#_c_376_n 0.0144623f $X=3.335 $Y=3.33 $X2=0
+ $Y2=0
cc_227 N_VPWR_c_324_n N_A_357_392#_c_376_n 0.0118344f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_228 N_VPWR_c_327_n N_A_357_392#_c_377_n 0.0247884f $X=3.5 $Y=2.145 $X2=0
+ $Y2=0
cc_229 N_VPWR_c_327_n N_A_357_392#_c_378_n 0.0323086f $X=3.5 $Y=2.145 $X2=0
+ $Y2=0
cc_230 N_VPWR_c_332_n N_A_357_392#_c_378_n 0.014549f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_231 N_VPWR_c_324_n N_A_357_392#_c_378_n 0.0119743f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_232 N_VPWR_c_327_n N_A_357_392#_c_379_n 0.0352735f $X=3.5 $Y=2.145 $X2=0
+ $Y2=0

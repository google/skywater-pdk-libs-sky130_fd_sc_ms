# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__o41ai_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__o41ai_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.810000 1.350000 3.235000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 1.920000 2.295000 2.890000 ;
        RECT 2.125000 1.350000 2.525000 1.680000 ;
        RECT 2.125000 1.680000 2.295000 1.920000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 1.350000 1.955000 1.680000 ;
        RECT 1.565000 1.680000 1.795000 2.890000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055000 1.350000 1.385000 1.780000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.180000 0.435000 1.550000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.569300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.350000 0.775000 1.010000 ;
        RECT 0.605000 1.010000 0.775000 1.350000 ;
        RECT 0.605000 1.350000 0.885000 1.520000 ;
        RECT 0.715000 1.520000 0.885000 1.950000 ;
        RECT 0.715000 1.950000 1.165000 2.120000 ;
        RECT 0.835000 2.120000 1.165000 2.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.115000  1.820000 0.545000 2.650000 ;
      RECT 0.115000  2.650000 0.665000 3.245000 ;
      RECT 0.955000  0.350000 1.205000 1.010000 ;
      RECT 0.955000  1.010000 3.220000 1.180000 ;
      RECT 1.375000  0.085000 1.705000 0.840000 ;
      RECT 1.890000  0.350000 2.220000 1.010000 ;
      RECT 2.390000  0.085000 2.720000 0.840000 ;
      RECT 2.890000  0.350000 3.220000 1.010000 ;
      RECT 2.995000  1.950000 3.245000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_ms__o41ai_1
END LIBRARY

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfsbp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
M1000 VPWR a_2067_74# a_3177_368# VPB pshort w=1e+06u l=180000u
+  ad=3.4604e+12p pd=2.71e+07u as=2.8e+11p ps=2.56e+06u
M1001 VGND a_3177_368# Q VNB nlowvt w=740000u l=150000u
+  ad=2.2419e+12p pd=2.069e+07u as=2.072e+11p ps=2.04e+06u
M1002 a_1204_463# a_619_368# a_1069_81# VPB pshort w=420000u l=180000u
+  ad=1.008e+11p pd=1.32e+06u as=1.344e+11p ps=1.48e+06u
M1003 a_1789_424# a_1069_81# VPWR VPB pshort w=840000u l=180000u
+  ad=7.392e+11p pd=6.8e+06u as=0p ps=0u
M1004 Q_N a_2067_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1005 VGND a_1069_81# a_1794_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=6.208e+11p ps=5.78e+06u
M1006 a_1069_81# a_871_74# a_307_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=3.672e+11p ps=3.46e+06u
M1007 a_223_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1008 a_2501_74# a_619_368# a_2067_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=5.999e+11p ps=4.61e+06u
M1009 VPWR SCE a_27_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1010 a_2067_74# a_871_74# a_2277_455# VPB pshort w=420000u l=180000u
+  ad=4.62e+11p pd=5.02e+06u as=2.373e+11p ps=2.81e+06u
M1011 a_1794_74# a_1069_81# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_2067_74# a_3177_368# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1013 a_1567_74# a_1069_81# a_1252_376# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1014 VGND SET_B a_1567_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND SCD a_495_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1016 VPWR a_2513_258# a_2277_455# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_495_74# SCE a_307_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=4.515e+11p ps=3.83e+06u
M1018 a_2067_74# SET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1069_81# a_619_368# a_307_74# VNB nlowvt w=420000u l=150000u
+  ad=3.675e+11p pd=2.59e+06u as=0p ps=0u
M1020 a_2579_74# a_2513_258# a_2501_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1021 VGND SET_B a_2579_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Q a_3177_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q_N a_2067_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.22e+11p pd=2.08e+06u as=0p ps=0u
M1024 VGND a_1252_376# a_1274_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1025 VGND a_2067_74# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1274_81# a_871_74# a_1069_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_421_464# a_27_74# a_307_74# VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1028 a_2067_74# a_619_368# a_1789_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR a_2067_74# Q_N VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR a_1252_376# a_1204_463# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1789_424# a_619_368# a_2067_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1794_74# a_871_74# a_2067_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_307_74# D a_223_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR SET_B a_1252_376# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.554e+11p ps=1.58e+06u
M1035 a_871_74# a_619_368# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1036 VPWR CLK a_619_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1037 a_229_74# a_27_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1038 a_307_74# D a_229_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_2067_74# a_871_74# a_1794_74# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_2513_258# a_2067_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1041 VPWR SCD a_421_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 a_1252_376# a_1069_81# VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VGND CLK a_619_368# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1044 VGND SCE a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1045 VPWR a_2067_74# a_2513_258# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1046 a_871_74# a_619_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.528e+11p pd=2.87e+06u as=0p ps=0u
M1047 Q a_3177_368# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1048 VPWR a_1069_81# a_1789_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1049 VPWR a_3177_368# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

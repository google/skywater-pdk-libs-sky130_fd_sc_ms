* File: sky130_fd_sc_ms__o22a_2.pxi.spice
* Created: Fri Aug 28 17:58:20 2020
* 
x_PM_SKY130_FD_SC_MS__O22A_2%A_82_48# N_A_82_48#_M1003_d N_A_82_48#_M1008_d
+ N_A_82_48#_M1004_g N_A_82_48#_M1001_g N_A_82_48#_M1009_g N_A_82_48#_M1002_g
+ N_A_82_48#_c_76_n N_A_82_48#_c_77_n N_A_82_48#_c_89_p N_A_82_48#_c_117_p
+ N_A_82_48#_c_106_p N_A_82_48#_c_86_n N_A_82_48#_c_78_n N_A_82_48#_c_79_n
+ N_A_82_48#_c_80_n N_A_82_48#_c_81_n N_A_82_48#_c_82_n
+ PM_SKY130_FD_SC_MS__O22A_2%A_82_48#
x_PM_SKY130_FD_SC_MS__O22A_2%B1 N_B1_M1006_g N_B1_M1003_g B1 N_B1_c_171_n
+ PM_SKY130_FD_SC_MS__O22A_2%B1
x_PM_SKY130_FD_SC_MS__O22A_2%B2 N_B2_M1008_g N_B2_M1011_g B2 N_B2_c_208_n
+ N_B2_c_209_n PM_SKY130_FD_SC_MS__O22A_2%B2
x_PM_SKY130_FD_SC_MS__O22A_2%A2 N_A2_M1000_g N_A2_M1010_g A2 N_A2_c_246_n
+ PM_SKY130_FD_SC_MS__O22A_2%A2
x_PM_SKY130_FD_SC_MS__O22A_2%A1 N_A1_M1005_g N_A1_M1007_g A1 N_A1_c_281_n
+ N_A1_c_282_n PM_SKY130_FD_SC_MS__O22A_2%A1
x_PM_SKY130_FD_SC_MS__O22A_2%VPWR N_VPWR_M1001_s N_VPWR_M1002_s N_VPWR_M1005_d
+ N_VPWR_c_307_n N_VPWR_c_308_n N_VPWR_c_309_n N_VPWR_c_310_n N_VPWR_c_311_n
+ N_VPWR_c_312_n VPWR N_VPWR_c_313_n N_VPWR_c_314_n N_VPWR_c_306_n
+ PM_SKY130_FD_SC_MS__O22A_2%VPWR
x_PM_SKY130_FD_SC_MS__O22A_2%X N_X_M1004_d N_X_M1001_d N_X_c_350_n N_X_c_353_n
+ N_X_c_354_n N_X_c_351_n X PM_SKY130_FD_SC_MS__O22A_2%X
x_PM_SKY130_FD_SC_MS__O22A_2%VGND N_VGND_M1004_s N_VGND_M1009_s N_VGND_M1010_d
+ N_VGND_c_385_n N_VGND_c_386_n N_VGND_c_387_n N_VGND_c_388_n VGND
+ N_VGND_c_389_n N_VGND_c_390_n N_VGND_c_391_n N_VGND_c_392_n N_VGND_c_393_n
+ N_VGND_c_394_n PM_SKY130_FD_SC_MS__O22A_2%VGND
x_PM_SKY130_FD_SC_MS__O22A_2%A_307_74# N_A_307_74#_M1003_s N_A_307_74#_M1011_d
+ N_A_307_74#_M1007_d N_A_307_74#_c_435_n N_A_307_74#_c_436_n
+ N_A_307_74#_c_456_n N_A_307_74#_c_437_n N_A_307_74#_c_438_n
+ N_A_307_74#_c_439_n N_A_307_74#_c_440_n PM_SKY130_FD_SC_MS__O22A_2%A_307_74#
cc_1 VNB N_A_82_48#_M1004_g 0.0338946f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.74
cc_2 VNB N_A_82_48#_M1001_g 0.00231818f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.4
cc_3 VNB N_A_82_48#_M1009_g 0.0232514f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.74
cc_4 VNB N_A_82_48#_M1002_g 0.00172775f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=2.4
cc_5 VNB N_A_82_48#_c_76_n 4.10656e-19 $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=1.95
cc_6 VNB N_A_82_48#_c_77_n 0.00178028f $X=-0.19 $Y=-0.245 $X2=1.305 $Y2=1.005
cc_7 VNB N_A_82_48#_c_78_n 0.00319769f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.465
cc_8 VNB N_A_82_48#_c_79_n 0.00341558f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.3
cc_9 VNB N_A_82_48#_c_80_n 0.00372536f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=0.965
cc_10 VNB N_A_82_48#_c_81_n 0.0223221f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=0.965
cc_11 VNB N_A_82_48#_c_82_n 0.0715116f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.465
cc_12 VNB N_B1_M1003_g 0.033506f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.39
cc_13 VNB B1 0.0030524f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.74
cc_14 VNB N_B1_c_171_n 0.0258161f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.74
cc_15 VNB N_B2_M1011_g 0.0306575f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.39
cc_16 VNB N_B2_c_208_n 0.0187265f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.4
cc_17 VNB N_B2_c_209_n 0.00432046f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.4
cc_18 VNB N_A2_M1010_g 0.0311199f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.39
cc_19 VNB A2 0.00517424f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.74
cc_20 VNB N_A2_c_246_n 0.0175947f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.4
cc_21 VNB N_A1_M1005_g 0.00185507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A1_M1007_g 0.0300997f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.39
cc_23 VNB N_A1_c_281_n 0.058845f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.3
cc_24 VNB N_A1_c_282_n 0.00431187f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.74
cc_25 VNB N_VPWR_c_306_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.465
cc_26 VNB N_X_c_350_n 0.00210995f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.74
cc_27 VNB N_X_c_351_n 0.00432789f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.63
cc_28 VNB X 0.00435003f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=2.4
cc_29 VNB N_VGND_c_385_n 0.0105514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_386_n 0.0506785f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.4
cc_31 VNB N_VGND_c_387_n 0.00898285f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=0.74
cc_32 VNB N_VGND_c_388_n 0.00640205f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=2.4
cc_33 VNB N_VGND_c_389_n 0.0168951f $X=-0.19 $Y=-0.245 $X2=1.22 $Y2=1.3
cc_34 VNB N_VGND_c_390_n 0.0430142f $X=-0.19 $Y=-0.245 $X2=2.35 $Y2=2.035
cc_35 VNB N_VGND_c_391_n 0.0173909f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.63
cc_36 VNB N_VGND_c_392_n 0.234729f $X=-0.19 $Y=-0.245 $X2=2.115 $Y2=0.965
cc_37 VNB N_VGND_c_393_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.465
cc_38 VNB N_VGND_c_394_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.465
cc_39 VNB N_A_307_74#_c_435_n 0.00296475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_307_74#_c_436_n 0.00261637f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.4
cc_41 VNB N_A_307_74#_c_437_n 0.0128061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_307_74#_c_438_n 0.00950245f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.3
cc_43 VNB N_A_307_74#_c_439_n 0.0247745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_307_74#_c_440_n 0.00655754f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=2.4
cc_45 VPB N_A_82_48#_M1001_g 0.0273944f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=2.4
cc_46 VPB N_A_82_48#_M1002_g 0.0251787f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=2.4
cc_47 VPB N_A_82_48#_c_76_n 0.00302273f $X=-0.19 $Y=1.66 $X2=1.22 $Y2=1.95
cc_48 VPB N_A_82_48#_c_86_n 0.00301741f $X=-0.19 $Y=1.66 $X2=2.515 $Y2=2.775
cc_49 VPB N_B1_M1006_g 0.0233311f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB B1 0.00205071f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=0.74
cc_51 VPB N_B1_c_171_n 0.0151557f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=0.74
cc_52 VPB N_B2_M1008_g 0.0215094f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_53 VPB N_B2_c_208_n 0.00982355f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=2.4
cc_54 VPB N_B2_c_209_n 0.00404989f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=2.4
cc_55 VPB N_A2_M1000_g 0.0225926f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB A2 0.0144661f $X=-0.19 $Y=1.66 $X2=0.485 $Y2=0.74
cc_57 VPB N_A2_c_246_n 0.00982405f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=2.4
cc_58 VPB N_A1_M1005_g 0.0341513f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A1_c_282_n 0.00745299f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=0.74
cc_60 VPB N_VPWR_c_307_n 0.0128289f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_308_n 0.0679799f $X=-0.19 $Y=1.66 $X2=0.575 $Y2=2.4
cc_62 VPB N_VPWR_c_309_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=0.74
cc_63 VPB N_VPWR_c_310_n 0.0107623f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=2.4
cc_64 VPB N_VPWR_c_311_n 0.011929f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_312_n 0.0502522f $X=-0.19 $Y=1.66 $X2=1.22 $Y2=1.3
cc_66 VPB N_VPWR_c_313_n 0.0488009f $X=-0.19 $Y=1.66 $X2=1.305 $Y2=2.035
cc_67 VPB N_VPWR_c_314_n 0.0125729f $X=-0.19 $Y=1.66 $X2=2.005 $Y2=0.965
cc_68 VPB N_VPWR_c_306_n 0.0903043f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=1.465
cc_69 VPB N_X_c_353_n 0.00412671f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=1.3
cc_70 VPB N_X_c_354_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0.915 $Y2=0.74
cc_71 VPB N_X_c_351_n 0.00117649f $X=-0.19 $Y=1.66 $X2=1.025 $Y2=1.63
cc_72 N_A_82_48#_M1002_g N_B1_M1006_g 0.00810577f $X=1.025 $Y=2.4 $X2=0 $Y2=0
cc_73 N_A_82_48#_c_76_n N_B1_M1006_g 0.00297406f $X=1.22 $Y=1.95 $X2=0 $Y2=0
cc_74 N_A_82_48#_c_89_p N_B1_M1006_g 0.0189734f $X=2.35 $Y=2.035 $X2=0 $Y2=0
cc_75 N_A_82_48#_c_86_n N_B1_M1006_g 0.00269851f $X=2.515 $Y=2.775 $X2=0 $Y2=0
cc_76 N_A_82_48#_c_78_n N_B1_M1003_g 6.90513e-19 $X=1.14 $Y=1.465 $X2=0 $Y2=0
cc_77 N_A_82_48#_c_79_n N_B1_M1003_g 0.00407257f $X=1.14 $Y=1.3 $X2=0 $Y2=0
cc_78 N_A_82_48#_c_81_n N_B1_M1003_g 0.0176532f $X=2.005 $Y=0.965 $X2=0 $Y2=0
cc_79 N_A_82_48#_c_82_n N_B1_M1003_g 0.00353902f $X=1.025 $Y=1.465 $X2=0 $Y2=0
cc_80 N_A_82_48#_c_89_p B1 0.0229182f $X=2.35 $Y=2.035 $X2=0 $Y2=0
cc_81 N_A_82_48#_c_78_n B1 0.0201599f $X=1.14 $Y=1.465 $X2=0 $Y2=0
cc_82 N_A_82_48#_c_81_n B1 0.0164979f $X=2.005 $Y=0.965 $X2=0 $Y2=0
cc_83 N_A_82_48#_c_82_n B1 8.54661e-19 $X=1.025 $Y=1.465 $X2=0 $Y2=0
cc_84 N_A_82_48#_M1002_g N_B1_c_171_n 0.00271569f $X=1.025 $Y=2.4 $X2=0 $Y2=0
cc_85 N_A_82_48#_c_76_n N_B1_c_171_n 0.00103585f $X=1.22 $Y=1.95 $X2=0 $Y2=0
cc_86 N_A_82_48#_c_89_p N_B1_c_171_n 0.00123799f $X=2.35 $Y=2.035 $X2=0 $Y2=0
cc_87 N_A_82_48#_c_78_n N_B1_c_171_n 7.6891e-19 $X=1.14 $Y=1.465 $X2=0 $Y2=0
cc_88 N_A_82_48#_c_81_n N_B1_c_171_n 0.00171671f $X=2.005 $Y=0.965 $X2=0 $Y2=0
cc_89 N_A_82_48#_c_82_n N_B1_c_171_n 0.011184f $X=1.025 $Y=1.465 $X2=0 $Y2=0
cc_90 N_A_82_48#_c_89_p N_B2_M1008_g 0.0128923f $X=2.35 $Y=2.035 $X2=0 $Y2=0
cc_91 N_A_82_48#_c_106_p N_B2_M1008_g 8.84614e-19 $X=2.515 $Y=2.12 $X2=0 $Y2=0
cc_92 N_A_82_48#_c_86_n N_B2_M1008_g 0.0161086f $X=2.515 $Y=2.775 $X2=0 $Y2=0
cc_93 N_A_82_48#_c_80_n N_B2_M1011_g 0.00451145f $X=2.115 $Y=0.965 $X2=0 $Y2=0
cc_94 N_A_82_48#_c_106_p N_B2_c_208_n 7.2959e-19 $X=2.515 $Y=2.12 $X2=0 $Y2=0
cc_95 N_A_82_48#_c_80_n N_B2_c_208_n 0.00233443f $X=2.115 $Y=0.965 $X2=0 $Y2=0
cc_96 N_A_82_48#_c_89_p N_B2_c_209_n 0.0207991f $X=2.35 $Y=2.035 $X2=0 $Y2=0
cc_97 N_A_82_48#_c_106_p N_B2_c_209_n 0.0102522f $X=2.515 $Y=2.12 $X2=0 $Y2=0
cc_98 N_A_82_48#_c_80_n N_B2_c_209_n 0.0134587f $X=2.115 $Y=0.965 $X2=0 $Y2=0
cc_99 N_A_82_48#_c_86_n N_A2_M1000_g 5.53825e-19 $X=2.515 $Y=2.775 $X2=0 $Y2=0
cc_100 N_A_82_48#_c_76_n N_VPWR_M1002_s 0.00239514f $X=1.22 $Y=1.95 $X2=0 $Y2=0
cc_101 N_A_82_48#_c_89_p N_VPWR_M1002_s 0.0169622f $X=2.35 $Y=2.035 $X2=0 $Y2=0
cc_102 N_A_82_48#_c_117_p N_VPWR_M1002_s 0.00271221f $X=1.305 $Y=2.035 $X2=0
+ $Y2=0
cc_103 N_A_82_48#_M1001_g N_VPWR_c_308_n 0.00546761f $X=0.575 $Y=2.4 $X2=0 $Y2=0
cc_104 N_A_82_48#_c_82_n N_VPWR_c_308_n 0.00255704f $X=1.025 $Y=1.465 $X2=0
+ $Y2=0
cc_105 N_A_82_48#_M1001_g N_VPWR_c_309_n 0.005209f $X=0.575 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A_82_48#_M1002_g N_VPWR_c_309_n 0.005209f $X=1.025 $Y=2.4 $X2=0 $Y2=0
cc_107 N_A_82_48#_M1002_g N_VPWR_c_310_n 0.00311949f $X=1.025 $Y=2.4 $X2=0 $Y2=0
cc_108 N_A_82_48#_c_89_p N_VPWR_c_310_n 0.0344594f $X=2.35 $Y=2.035 $X2=0 $Y2=0
cc_109 N_A_82_48#_c_117_p N_VPWR_c_310_n 0.0119464f $X=1.305 $Y=2.035 $X2=0
+ $Y2=0
cc_110 N_A_82_48#_c_86_n N_VPWR_c_310_n 0.0193052f $X=2.515 $Y=2.775 $X2=0 $Y2=0
cc_111 N_A_82_48#_c_82_n N_VPWR_c_310_n 4.61822e-19 $X=1.025 $Y=1.465 $X2=0
+ $Y2=0
cc_112 N_A_82_48#_c_86_n N_VPWR_c_313_n 0.0125236f $X=2.515 $Y=2.775 $X2=0 $Y2=0
cc_113 N_A_82_48#_M1001_g N_VPWR_c_306_n 0.00985555f $X=0.575 $Y=2.4 $X2=0 $Y2=0
cc_114 N_A_82_48#_M1002_g N_VPWR_c_306_n 0.00986727f $X=1.025 $Y=2.4 $X2=0 $Y2=0
cc_115 N_A_82_48#_c_86_n N_VPWR_c_306_n 0.0117917f $X=2.515 $Y=2.775 $X2=0 $Y2=0
cc_116 N_A_82_48#_M1004_g N_X_c_350_n 0.00563952f $X=0.485 $Y=0.74 $X2=0 $Y2=0
cc_117 N_A_82_48#_M1009_g N_X_c_350_n 2.51515e-19 $X=0.915 $Y=0.74 $X2=0 $Y2=0
cc_118 N_A_82_48#_M1001_g N_X_c_353_n 0.00215936f $X=0.575 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A_82_48#_M1002_g N_X_c_353_n 0.003664f $X=1.025 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A_82_48#_c_76_n N_X_c_353_n 0.00559274f $X=1.22 $Y=1.95 $X2=0 $Y2=0
cc_121 N_A_82_48#_c_82_n N_X_c_353_n 0.0018941f $X=1.025 $Y=1.465 $X2=0 $Y2=0
cc_122 N_A_82_48#_M1001_g N_X_c_354_n 0.0127634f $X=0.575 $Y=2.4 $X2=0 $Y2=0
cc_123 N_A_82_48#_M1002_g N_X_c_354_n 0.0182659f $X=1.025 $Y=2.4 $X2=0 $Y2=0
cc_124 N_A_82_48#_M1004_g N_X_c_351_n 0.00602646f $X=0.485 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A_82_48#_M1001_g N_X_c_351_n 0.00903338f $X=0.575 $Y=2.4 $X2=0 $Y2=0
cc_126 N_A_82_48#_M1009_g N_X_c_351_n 0.0023958f $X=0.915 $Y=0.74 $X2=0 $Y2=0
cc_127 N_A_82_48#_M1002_g N_X_c_351_n 0.00150368f $X=1.025 $Y=2.4 $X2=0 $Y2=0
cc_128 N_A_82_48#_c_76_n N_X_c_351_n 0.00896365f $X=1.22 $Y=1.95 $X2=0 $Y2=0
cc_129 N_A_82_48#_c_78_n N_X_c_351_n 0.0239021f $X=1.14 $Y=1.465 $X2=0 $Y2=0
cc_130 N_A_82_48#_c_79_n N_X_c_351_n 0.00799225f $X=1.14 $Y=1.3 $X2=0 $Y2=0
cc_131 N_A_82_48#_c_82_n N_X_c_351_n 0.0202514f $X=1.025 $Y=1.465 $X2=0 $Y2=0
cc_132 N_A_82_48#_M1004_g X 0.00477711f $X=0.485 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A_82_48#_M1009_g X 0.00781845f $X=0.915 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A_82_48#_c_77_n X 0.0145044f $X=1.305 $Y=1.005 $X2=0 $Y2=0
cc_135 N_A_82_48#_c_89_p A_386_384# 0.00920959f $X=2.35 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_136 N_A_82_48#_c_77_n N_VGND_M1009_s 0.00509051f $X=1.305 $Y=1.005 $X2=0
+ $Y2=0
cc_137 N_A_82_48#_M1004_g N_VGND_c_386_n 0.00478246f $X=0.485 $Y=0.74 $X2=0
+ $Y2=0
cc_138 N_A_82_48#_M1004_g N_VGND_c_387_n 4.28647e-19 $X=0.485 $Y=0.74 $X2=0
+ $Y2=0
cc_139 N_A_82_48#_M1009_g N_VGND_c_387_n 0.00900614f $X=0.915 $Y=0.74 $X2=0
+ $Y2=0
cc_140 N_A_82_48#_c_77_n N_VGND_c_387_n 0.0112419f $X=1.305 $Y=1.005 $X2=0 $Y2=0
cc_141 N_A_82_48#_c_78_n N_VGND_c_387_n 0.00352695f $X=1.14 $Y=1.465 $X2=0 $Y2=0
cc_142 N_A_82_48#_c_82_n N_VGND_c_387_n 0.00118847f $X=1.025 $Y=1.465 $X2=0
+ $Y2=0
cc_143 N_A_82_48#_M1004_g N_VGND_c_389_n 0.00434272f $X=0.485 $Y=0.74 $X2=0
+ $Y2=0
cc_144 N_A_82_48#_M1009_g N_VGND_c_389_n 0.00383152f $X=0.915 $Y=0.74 $X2=0
+ $Y2=0
cc_145 N_A_82_48#_M1004_g N_VGND_c_392_n 0.00823683f $X=0.485 $Y=0.74 $X2=0
+ $Y2=0
cc_146 N_A_82_48#_M1009_g N_VGND_c_392_n 0.00685545f $X=0.915 $Y=0.74 $X2=0
+ $Y2=0
cc_147 N_A_82_48#_c_81_n N_A_307_74#_M1003_s 0.00296342f $X=2.005 $Y=0.965
+ $X2=-0.19 $Y2=-0.245
cc_148 N_A_82_48#_M1003_d N_A_307_74#_c_435_n 0.00262063f $X=1.96 $Y=0.37 $X2=0
+ $Y2=0
cc_149 N_A_82_48#_c_80_n N_A_307_74#_c_435_n 0.0104858f $X=2.115 $Y=0.965 $X2=0
+ $Y2=0
cc_150 N_A_82_48#_c_81_n N_A_307_74#_c_435_n 0.00476112f $X=2.005 $Y=0.965 $X2=0
+ $Y2=0
cc_151 N_A_82_48#_c_80_n N_A_307_74#_c_438_n 0.00799569f $X=2.115 $Y=0.965 $X2=0
+ $Y2=0
cc_152 N_A_82_48#_M1009_g N_A_307_74#_c_440_n 5.23807e-19 $X=0.915 $Y=0.74 $X2=0
+ $Y2=0
cc_153 N_A_82_48#_c_81_n N_A_307_74#_c_440_n 0.021503f $X=2.005 $Y=0.965 $X2=0
+ $Y2=0
cc_154 N_B1_M1006_g N_B2_M1008_g 0.0601804f $X=1.84 $Y=2.42 $X2=0 $Y2=0
cc_155 N_B1_M1003_g N_B2_M1011_g 0.0358967f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_156 B1 N_B2_c_208_n 2.82156e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_157 N_B1_c_171_n N_B2_c_208_n 0.0207707f $X=1.885 $Y=1.595 $X2=0 $Y2=0
cc_158 B1 N_B2_c_209_n 0.0283557f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_159 N_B1_c_171_n N_B2_c_209_n 0.00234411f $X=1.885 $Y=1.595 $X2=0 $Y2=0
cc_160 N_B1_M1006_g N_VPWR_c_310_n 0.0190291f $X=1.84 $Y=2.42 $X2=0 $Y2=0
cc_161 N_B1_M1006_g N_VPWR_c_313_n 0.00510822f $X=1.84 $Y=2.42 $X2=0 $Y2=0
cc_162 N_B1_M1006_g N_VPWR_c_306_n 0.00501096f $X=1.84 $Y=2.42 $X2=0 $Y2=0
cc_163 N_B1_M1003_g N_VGND_c_387_n 0.00332629f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_164 N_B1_M1003_g N_VGND_c_390_n 0.00292759f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_165 N_B1_M1003_g N_VGND_c_392_n 0.00363526f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_166 N_B1_M1003_g N_A_307_74#_c_435_n 0.0084546f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_167 N_B1_M1003_g N_A_307_74#_c_440_n 0.00558709f $X=1.885 $Y=0.74 $X2=0 $Y2=0
cc_168 N_B2_M1008_g N_A2_M1000_g 0.0126006f $X=2.29 $Y=2.42 $X2=0 $Y2=0
cc_169 N_B2_M1011_g N_A2_M1010_g 0.0286716f $X=2.345 $Y=0.74 $X2=0 $Y2=0
cc_170 N_B2_c_208_n A2 4.13796e-19 $X=2.335 $Y=1.595 $X2=0 $Y2=0
cc_171 N_B2_c_209_n A2 0.023664f $X=2.335 $Y=1.595 $X2=0 $Y2=0
cc_172 N_B2_c_208_n N_A2_c_246_n 0.0214219f $X=2.335 $Y=1.595 $X2=0 $Y2=0
cc_173 N_B2_c_209_n N_A2_c_246_n 4.14534e-19 $X=2.335 $Y=1.595 $X2=0 $Y2=0
cc_174 N_B2_M1008_g N_VPWR_c_310_n 0.00244913f $X=2.29 $Y=2.42 $X2=0 $Y2=0
cc_175 N_B2_M1008_g N_VPWR_c_313_n 0.00628513f $X=2.29 $Y=2.42 $X2=0 $Y2=0
cc_176 N_B2_M1008_g N_VPWR_c_306_n 0.00639697f $X=2.29 $Y=2.42 $X2=0 $Y2=0
cc_177 N_B2_M1011_g N_VGND_c_390_n 0.00291649f $X=2.345 $Y=0.74 $X2=0 $Y2=0
cc_178 N_B2_M1011_g N_VGND_c_392_n 0.00360203f $X=2.345 $Y=0.74 $X2=0 $Y2=0
cc_179 N_B2_M1011_g N_A_307_74#_c_435_n 0.014305f $X=2.345 $Y=0.74 $X2=0 $Y2=0
cc_180 N_B2_M1011_g N_A_307_74#_c_438_n 9.8635e-19 $X=2.345 $Y=0.74 $X2=0 $Y2=0
cc_181 N_B2_c_208_n N_A_307_74#_c_438_n 7.565e-19 $X=2.335 $Y=1.595 $X2=0 $Y2=0
cc_182 N_B2_c_209_n N_A_307_74#_c_438_n 0.00194208f $X=2.335 $Y=1.595 $X2=0
+ $Y2=0
cc_183 N_B2_M1011_g N_A_307_74#_c_440_n 6.68686e-19 $X=2.345 $Y=0.74 $X2=0 $Y2=0
cc_184 N_A2_M1000_g N_A1_M1005_g 0.0431129f $X=2.8 $Y=2.42 $X2=0 $Y2=0
cc_185 N_A2_M1010_g N_A1_M1007_g 0.0278115f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_186 N_A2_M1010_g N_A1_c_281_n 0.00558036f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_187 A2 N_A1_c_281_n 0.00287477f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_188 N_A2_c_246_n N_A1_c_281_n 0.020345f $X=2.875 $Y=1.595 $X2=0 $Y2=0
cc_189 N_A2_M1010_g N_A1_c_282_n 5.8609e-19 $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_190 A2 N_A1_c_282_n 0.0286864f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_191 N_A2_c_246_n N_A1_c_282_n 2.28512e-19 $X=2.875 $Y=1.595 $X2=0 $Y2=0
cc_192 N_A2_M1000_g N_VPWR_c_312_n 0.00506203f $X=2.8 $Y=2.42 $X2=0 $Y2=0
cc_193 N_A2_M1000_g N_VPWR_c_313_n 0.00658449f $X=2.8 $Y=2.42 $X2=0 $Y2=0
cc_194 N_A2_M1000_g N_VPWR_c_306_n 0.00639697f $X=2.8 $Y=2.42 $X2=0 $Y2=0
cc_195 N_A2_M1010_g N_VGND_c_388_n 0.00544936f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A2_M1010_g N_VGND_c_390_n 0.00433139f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_197 N_A2_M1010_g N_VGND_c_392_n 0.00817815f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_198 N_A2_M1010_g N_A_307_74#_c_436_n 0.00225753f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_199 N_A2_M1010_g N_A_307_74#_c_456_n 0.00673645f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_200 N_A2_M1010_g N_A_307_74#_c_437_n 0.0120938f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_201 A2 N_A_307_74#_c_437_n 0.0220803f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_202 N_A2_c_246_n N_A_307_74#_c_437_n 0.00245655f $X=2.875 $Y=1.595 $X2=0
+ $Y2=0
cc_203 N_A2_M1010_g N_A_307_74#_c_438_n 0.00109647f $X=2.845 $Y=0.74 $X2=0 $Y2=0
cc_204 A2 N_A_307_74#_c_438_n 0.00459921f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_205 N_A2_c_246_n N_A_307_74#_c_438_n 0.00150281f $X=2.875 $Y=1.595 $X2=0
+ $Y2=0
cc_206 N_A1_M1005_g N_VPWR_c_312_n 0.0262879f $X=3.34 $Y=2.42 $X2=0 $Y2=0
cc_207 N_A1_c_281_n N_VPWR_c_312_n 0.00152096f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_208 N_A1_c_282_n N_VPWR_c_312_n 0.0261817f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_209 N_A1_M1005_g N_VPWR_c_313_n 0.00547402f $X=3.34 $Y=2.42 $X2=0 $Y2=0
cc_210 N_A1_M1005_g N_VPWR_c_306_n 0.00536634f $X=3.34 $Y=2.42 $X2=0 $Y2=0
cc_211 N_A1_M1007_g N_VGND_c_388_n 0.012583f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_212 N_A1_M1007_g N_VGND_c_391_n 0.00383152f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_213 N_A1_M1007_g N_VGND_c_392_n 0.00761198f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A1_M1007_g N_A_307_74#_c_456_n 7.30686e-19 $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_215 N_A1_M1007_g N_A_307_74#_c_437_n 0.0171242f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A1_c_281_n N_A_307_74#_c_437_n 0.00319341f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_217 N_A1_c_282_n N_A_307_74#_c_437_n 0.0270164f $X=3.57 $Y=1.465 $X2=0 $Y2=0
cc_218 N_A1_M1007_g N_A_307_74#_c_439_n 0.00159319f $X=3.345 $Y=0.74 $X2=0 $Y2=0
cc_219 N_VPWR_c_308_n N_X_c_353_n 0.0450694f $X=0.3 $Y=1.985 $X2=0 $Y2=0
cc_220 N_VPWR_c_309_n N_X_c_354_n 0.0144623f $X=1.135 $Y=3.33 $X2=0 $Y2=0
cc_221 N_VPWR_c_310_n N_X_c_354_n 0.0267671f $X=1.615 $Y=2.41 $X2=0 $Y2=0
cc_222 N_VPWR_c_306_n N_X_c_354_n 0.0118344f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_223 N_X_c_350_n N_VGND_c_386_n 0.0300732f $X=0.7 $Y=0.515 $X2=0 $Y2=0
cc_224 N_X_c_350_n N_VGND_c_387_n 0.0113761f $X=0.7 $Y=0.515 $X2=0 $Y2=0
cc_225 N_X_c_350_n N_VGND_c_389_n 0.0112174f $X=0.7 $Y=0.515 $X2=0 $Y2=0
cc_226 N_X_c_350_n N_VGND_c_392_n 0.00922837f $X=0.7 $Y=0.515 $X2=0 $Y2=0
cc_227 X N_VGND_c_392_n 0.0025861f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_228 N_VGND_c_390_n N_A_307_74#_c_435_n 0.0247246f $X=2.965 $Y=0 $X2=0 $Y2=0
cc_229 N_VGND_c_392_n N_A_307_74#_c_435_n 0.0209615f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_230 N_VGND_c_388_n N_A_307_74#_c_436_n 0.00795492f $X=3.13 $Y=0.625 $X2=0
+ $Y2=0
cc_231 N_VGND_c_390_n N_A_307_74#_c_436_n 0.0146502f $X=2.965 $Y=0 $X2=0 $Y2=0
cc_232 N_VGND_c_392_n N_A_307_74#_c_436_n 0.0120674f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_233 N_VGND_M1010_d N_A_307_74#_c_437_n 0.00250873f $X=2.92 $Y=0.37 $X2=0
+ $Y2=0
cc_234 N_VGND_c_388_n N_A_307_74#_c_437_n 0.0209867f $X=3.13 $Y=0.625 $X2=0
+ $Y2=0
cc_235 N_VGND_c_388_n N_A_307_74#_c_439_n 0.0164982f $X=3.13 $Y=0.625 $X2=0
+ $Y2=0
cc_236 N_VGND_c_391_n N_A_307_74#_c_439_n 0.011066f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_237 N_VGND_c_392_n N_A_307_74#_c_439_n 0.00915947f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_238 N_VGND_c_387_n N_A_307_74#_c_440_n 0.0208243f $X=1.13 $Y=0.535 $X2=0
+ $Y2=0
cc_239 N_VGND_c_390_n N_A_307_74#_c_440_n 0.0139208f $X=2.965 $Y=0 $X2=0 $Y2=0
cc_240 N_VGND_c_392_n N_A_307_74#_c_440_n 0.0117508f $X=3.6 $Y=0 $X2=0 $Y2=0

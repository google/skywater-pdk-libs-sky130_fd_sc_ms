* File: sky130_fd_sc_ms__o311ai_4.pex.spice
* Created: Fri Aug 28 18:01:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O311AI_4%C1 3 5 7 8 10 13 15 17 18 19 20 22 23 24 35
r68 34 36 12.5272 $w=4.04e-07 $l=1.05e-07 $layer=POLY_cond $X=1.075 $Y=1.407
+ $X2=1.18 $Y2=1.407
r69 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.075
+ $Y=1.465 $X2=1.075 $Y2=1.465
r70 32 34 17.2995 $w=4.04e-07 $l=1.45e-07 $layer=POLY_cond $X=0.93 $Y=1.407
+ $X2=1.075 $Y2=1.407
r71 31 32 50.7054 $w=4.04e-07 $l=4.25e-07 $layer=POLY_cond $X=0.505 $Y=1.407
+ $X2=0.93 $Y2=1.407
r72 30 31 1.19307 $w=4.04e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.407
+ $X2=0.505 $Y2=1.407
r73 28 30 11.9307 $w=4.04e-07 $l=1e-07 $layer=POLY_cond $X=0.395 $Y=1.407
+ $X2=0.495 $Y2=1.407
r74 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.395
+ $Y=1.465 $X2=0.395 $Y2=1.465
r75 24 35 8.846 $w=4.78e-07 $l=3.55e-07 $layer=LI1_cond $X=0.72 $Y=1.54
+ $X2=1.075 $Y2=1.54
r76 24 29 8.09845 $w=4.78e-07 $l=3.25e-07 $layer=LI1_cond $X=0.72 $Y=1.54
+ $X2=0.395 $Y2=1.54
r77 23 29 3.86234 $w=4.78e-07 $l=1.55e-07 $layer=LI1_cond $X=0.24 $Y=1.54
+ $X2=0.395 $Y2=1.54
r78 20 22 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.79 $Y=1.185
+ $X2=1.79 $Y2=0.74
r79 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.715 $Y=1.26
+ $X2=1.79 $Y2=1.185
r80 18 19 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.715 $Y=1.26
+ $X2=1.435 $Y2=1.26
r81 15 19 28.927 $w=4.04e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.36 $Y=1.185
+ $X2=1.435 $Y2=1.26
r82 15 36 21.4752 $w=4.04e-07 $l=2.98737e-07 $layer=POLY_cond $X=1.36 $Y=1.185
+ $X2=1.18 $Y2=1.407
r83 15 17 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.36 $Y=1.185
+ $X2=1.36 $Y2=0.74
r84 11 36 21.6995 $w=1.8e-07 $l=2.23e-07 $layer=POLY_cond $X=1.18 $Y=1.63
+ $X2=1.18 $Y2=1.407
r85 11 13 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=1.18 $Y=1.63
+ $X2=1.18 $Y2=2.4
r86 8 32 26.1054 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=0.93 $Y=1.185
+ $X2=0.93 $Y2=1.407
r87 8 10 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.93 $Y=1.185
+ $X2=0.93 $Y2=0.74
r88 5 30 26.1054 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=0.495 $Y=1.185
+ $X2=0.495 $Y2=1.407
r89 5 7 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.495 $Y=1.185
+ $X2=0.495 $Y2=0.74
r90 1 31 21.6995 $w=1.8e-07 $l=2.23e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=1.407
r91 1 3 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O311AI_4%B1 1 3 4 5 6 8 11 15 19 23 25 26 27 28 41
r63 41 43 12.0836 $w=3.59e-07 $l=9e-08 $layer=POLY_cond $X=3.43 $Y=1.537
+ $X2=3.52 $Y2=1.537
r64 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.43
+ $Y=1.515 $X2=3.43 $Y2=1.515
r65 39 41 46.9916 $w=3.59e-07 $l=3.5e-07 $layer=POLY_cond $X=3.08 $Y=1.537
+ $X2=3.43 $Y2=1.537
r66 38 39 57.7326 $w=3.59e-07 $l=4.3e-07 $layer=POLY_cond $X=2.65 $Y=1.537
+ $X2=3.08 $Y2=1.537
r67 36 38 32.2228 $w=3.59e-07 $l=2.4e-07 $layer=POLY_cond $X=2.41 $Y=1.537
+ $X2=2.65 $Y2=1.537
r68 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.41
+ $Y=1.515 $X2=2.41 $Y2=1.515
r69 34 36 25.5097 $w=3.59e-07 $l=1.9e-07 $layer=POLY_cond $X=2.22 $Y=1.537
+ $X2=2.41 $Y2=1.537
r70 27 28 15.8049 $w=3.48e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.605
+ $X2=4.08 $Y2=1.605
r71 27 42 5.59758 $w=3.48e-07 $l=1.7e-07 $layer=LI1_cond $X=3.6 $Y=1.605
+ $X2=3.43 $Y2=1.605
r72 26 42 10.2074 $w=3.48e-07 $l=3.1e-07 $layer=LI1_cond $X=3.12 $Y=1.605
+ $X2=3.43 $Y2=1.605
r73 25 26 15.8049 $w=3.48e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.605
+ $X2=3.12 $Y2=1.605
r74 25 37 7.5732 $w=3.48e-07 $l=2.3e-07 $layer=LI1_cond $X=2.64 $Y=1.605
+ $X2=2.41 $Y2=1.605
r75 21 43 23.2387 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=3.52 $Y=1.35
+ $X2=3.52 $Y2=1.537
r76 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.52 $Y=1.35
+ $X2=3.52 $Y2=0.74
r77 17 39 23.2387 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=3.08 $Y=1.35
+ $X2=3.08 $Y2=1.537
r78 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.08 $Y=1.35
+ $X2=3.08 $Y2=0.74
r79 13 38 23.2387 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=2.65 $Y=1.35
+ $X2=2.65 $Y2=1.537
r80 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.65 $Y=1.35
+ $X2=2.65 $Y2=0.74
r81 9 34 23.2387 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=2.22 $Y=1.35
+ $X2=2.22 $Y2=1.537
r82 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.22 $Y=1.35 $X2=2.22
+ $Y2=0.74
r83 6 34 12.0836 $w=3.59e-07 $l=2.28613e-07 $layer=POLY_cond $X=2.13 $Y=1.725
+ $X2=2.22 $Y2=1.537
r84 6 8 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=2.13 $Y=1.725 $X2=2.13
+ $Y2=2.4
r85 4 6 28.8271 $w=3.59e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.04 $Y=1.65
+ $X2=2.13 $Y2=1.725
r86 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.04 $Y=1.65 $X2=1.77
+ $Y2=1.65
r87 1 5 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.68 $Y=1.725
+ $X2=1.77 $Y2=1.65
r88 1 3 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=1.68 $Y=1.725 $X2=1.68
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O311AI_4%A3 3 7 11 15 19 23 27 31 38 39 56 58 60 67
+ 70
c98 58 0 1.61783e-19 $X=6.24 $Y=1.515
r99 60 70 0.493904 $w=3.48e-07 $l=1.5e-08 $layer=LI1_cond $X=5.535 $Y=1.605
+ $X2=5.52 $Y2=1.605
r100 57 58 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.225 $Y=1.515
+ $X2=6.24 $Y2=1.515
r101 55 57 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=6.03 $Y=1.515
+ $X2=6.225 $Y2=1.515
r102 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.03
+ $Y=1.515 $X2=6.03 $Y2=1.515
r103 53 55 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=5.81 $Y=1.515
+ $X2=6.03 $Y2=1.515
r104 52 53 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=5.595 $Y=1.515
+ $X2=5.81 $Y2=1.515
r105 51 67 7.26255 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.35 $Y=1.605
+ $X2=5.185 $Y2=1.605
r106 50 52 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=5.35 $Y=1.515
+ $X2=5.595 $Y2=1.515
r107 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.35
+ $Y=1.515 $X2=5.35 $Y2=1.515
r108 48 50 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=5.22 $Y=1.515
+ $X2=5.35 $Y2=1.515
r109 47 48 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=5.075 $Y=1.515
+ $X2=5.22 $Y2=1.515
r110 43 45 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=4.575 $Y=1.515
+ $X2=4.79 $Y2=1.515
r111 39 56 0.987808 $w=3.48e-07 $l=3e-08 $layer=LI1_cond $X=6 $Y=1.605 $X2=6.03
+ $Y2=1.605
r112 38 70 1.15244 $w=3.48e-07 $l=3.5e-08 $layer=LI1_cond $X=5.485 $Y=1.605
+ $X2=5.52 $Y2=1.605
r113 38 51 4.44514 $w=3.48e-07 $l=1.35e-07 $layer=LI1_cond $X=5.485 $Y=1.605
+ $X2=5.35 $Y2=1.605
r114 38 39 14.1586 $w=3.48e-07 $l=4.3e-07 $layer=LI1_cond $X=5.57 $Y=1.605 $X2=6
+ $Y2=1.605
r115 38 60 1.15244 $w=3.48e-07 $l=3.5e-08 $layer=LI1_cond $X=5.57 $Y=1.605
+ $X2=5.535 $Y2=1.605
r116 36 47 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=5.01 $Y=1.515
+ $X2=5.075 $Y2=1.515
r117 36 45 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=5.01 $Y=1.515
+ $X2=4.79 $Y2=1.515
r118 35 67 9.24242 $w=2.08e-07 $l=1.75e-07 $layer=LI1_cond $X=5.01 $Y=1.535
+ $X2=5.185 $Y2=1.535
r119 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.01
+ $Y=1.515 $X2=5.01 $Y2=1.515
r120 29 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.24 $Y=1.35
+ $X2=6.24 $Y2=1.515
r121 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.24 $Y=1.35
+ $X2=6.24 $Y2=0.74
r122 25 57 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.225 $Y=1.68
+ $X2=6.225 $Y2=1.515
r123 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.225 $Y=1.68
+ $X2=6.225 $Y2=2.4
r124 21 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.81 $Y=1.35
+ $X2=5.81 $Y2=1.515
r125 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.81 $Y=1.35
+ $X2=5.81 $Y2=0.74
r126 17 52 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.595 $Y=1.68
+ $X2=5.595 $Y2=1.515
r127 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.595 $Y=1.68
+ $X2=5.595 $Y2=2.4
r128 13 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.22 $Y=1.35
+ $X2=5.22 $Y2=1.515
r129 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.22 $Y=1.35
+ $X2=5.22 $Y2=0.74
r130 9 47 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.075 $Y=1.68
+ $X2=5.075 $Y2=1.515
r131 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.075 $Y=1.68
+ $X2=5.075 $Y2=2.4
r132 5 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.79 $Y=1.35
+ $X2=4.79 $Y2=1.515
r133 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.79 $Y=1.35 $X2=4.79
+ $Y2=0.74
r134 1 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.575 $Y=1.68
+ $X2=4.575 $Y2=1.515
r135 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=4.575 $Y=1.68
+ $X2=4.575 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O311AI_4%A2 3 7 11 15 19 21 23 26 28 30 31 32 44 47
c93 28 0 5.87245e-20 $X=8.245 $Y=1.2
c94 15 0 1.36796e-19 $X=7.27 $Y=0.74
c95 11 0 9.26431e-20 $X=7.175 $Y=2.4
c96 7 0 5.58611e-20 $X=6.84 $Y=0.74
r97 47 48 9.24384 $w=3.65e-07 $l=7e-08 $layer=POLY_cond $X=8.175 $Y=1.44
+ $X2=8.245 $Y2=1.44
r98 46 47 57.4438 $w=3.65e-07 $l=4.35e-07 $layer=POLY_cond $X=7.74 $Y=1.44
+ $X2=8.175 $Y2=1.44
r99 45 46 1.98082 $w=3.65e-07 $l=1.5e-08 $layer=POLY_cond $X=7.725 $Y=1.44
+ $X2=7.74 $Y2=1.44
r100 43 45 15.1863 $w=3.65e-07 $l=1.15e-07 $layer=POLY_cond $X=7.61 $Y=1.44
+ $X2=7.725 $Y2=1.44
r101 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.61
+ $Y=1.515 $X2=7.61 $Y2=1.515
r102 38 40 32.3534 $w=3.65e-07 $l=2.45e-07 $layer=POLY_cond $X=6.93 $Y=1.44
+ $X2=7.175 $Y2=1.44
r103 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.93
+ $Y=1.515 $X2=6.93 $Y2=1.515
r104 32 44 4.55617 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.61 $Y2=1.565
r105 31 32 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.44 $Y2=1.565
r106 31 39 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=6.93 $Y2=1.565
r107 28 48 23.6381 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=8.245 $Y=1.2
+ $X2=8.245 $Y2=1.44
r108 28 30 147.813 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=8.245 $Y=1.2
+ $X2=8.245 $Y2=0.74
r109 24 47 19.2931 $w=1.8e-07 $l=2e-07 $layer=POLY_cond $X=8.175 $Y=1.64
+ $X2=8.175 $Y2=1.44
r110 24 26 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=8.175 $Y=1.64
+ $X2=8.175 $Y2=2.4
r111 21 46 23.6381 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=7.74 $Y=1.2
+ $X2=7.74 $Y2=1.44
r112 21 23 147.813 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=7.74 $Y=1.2
+ $X2=7.74 $Y2=0.74
r113 17 45 19.2931 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=7.725 $Y=1.68
+ $X2=7.725 $Y2=1.44
r114 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.725 $Y=1.68
+ $X2=7.725 $Y2=2.4
r115 13 43 44.8986 $w=3.65e-07 $l=3.4e-07 $layer=POLY_cond $X=7.27 $Y=1.44
+ $X2=7.61 $Y2=1.44
r116 13 40 12.5452 $w=3.65e-07 $l=9.5e-08 $layer=POLY_cond $X=7.27 $Y=1.44
+ $X2=7.175 $Y2=1.44
r117 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.27 $Y=1.35
+ $X2=7.27 $Y2=0.74
r118 9 40 19.2931 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=7.175 $Y=1.68
+ $X2=7.175 $Y2=1.44
r119 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.175 $Y=1.68
+ $X2=7.175 $Y2=2.4
r120 5 38 11.8849 $w=3.65e-07 $l=9e-08 $layer=POLY_cond $X=6.84 $Y=1.44 $X2=6.93
+ $Y2=1.44
r121 5 35 21.789 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=6.84 $Y=1.44
+ $X2=6.675 $Y2=1.44
r122 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.84 $Y=1.35 $X2=6.84
+ $Y2=0.74
r123 1 35 19.2931 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=6.675 $Y=1.68
+ $X2=6.675 $Y2=1.44
r124 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.675 $Y=1.68
+ $X2=6.675 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O311AI_4%A1 3 5 6 9 13 17 21 23 25 28 30 32 33 34 35
+ 49 50
c82 30 0 1.65594e-19 $X=10.545 $Y=1.2
r83 50 51 1.25195 $w=3.85e-07 $l=1e-08 $layer=POLY_cond $X=10.535 $Y=1.44
+ $X2=10.545 $Y2=1.44
r84 48 50 23.161 $w=3.85e-07 $l=1.85e-07 $layer=POLY_cond $X=10.35 $Y=1.44
+ $X2=10.535 $Y2=1.44
r85 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.35
+ $Y=1.515 $X2=10.35 $Y2=1.515
r86 46 48 31.2987 $w=3.85e-07 $l=2.5e-07 $layer=POLY_cond $X=10.1 $Y=1.44
+ $X2=10.35 $Y2=1.44
r87 45 46 1.87792 $w=3.85e-07 $l=1.5e-08 $layer=POLY_cond $X=10.085 $Y=1.44
+ $X2=10.1 $Y2=1.44
r88 44 45 56.3377 $w=3.85e-07 $l=4.5e-07 $layer=POLY_cond $X=9.635 $Y=1.44
+ $X2=10.085 $Y2=1.44
r89 42 44 38.1844 $w=3.85e-07 $l=3.05e-07 $layer=POLY_cond $X=9.33 $Y=1.44
+ $X2=9.635 $Y2=1.44
r90 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.33
+ $Y=1.515 $X2=9.33 $Y2=1.515
r91 40 42 18.1532 $w=3.85e-07 $l=1.45e-07 $layer=POLY_cond $X=9.185 $Y=1.44
+ $X2=9.33 $Y2=1.44
r92 35 49 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=10.32 $Y=1.565
+ $X2=10.35 $Y2=1.565
r93 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=9.84 $Y=1.565
+ $X2=10.32 $Y2=1.565
r94 33 34 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=9.36 $Y=1.565
+ $X2=9.84 $Y2=1.565
r95 33 43 0.80403 $w=4.28e-07 $l=3e-08 $layer=LI1_cond $X=9.36 $Y=1.565 $X2=9.33
+ $Y2=1.565
r96 30 51 24.9301 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=10.545 $Y=1.2
+ $X2=10.545 $Y2=1.44
r97 30 32 147.813 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=10.545 $Y=1.2
+ $X2=10.545 $Y2=0.74
r98 26 50 20.5538 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=10.535 $Y=1.68
+ $X2=10.535 $Y2=1.44
r99 26 28 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=10.535 $Y=1.68
+ $X2=10.535 $Y2=2.4
r100 23 46 24.9301 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=10.1 $Y=1.2
+ $X2=10.1 $Y2=1.44
r101 23 25 147.813 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=10.1 $Y=1.2
+ $X2=10.1 $Y2=0.74
r102 19 45 20.5538 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=10.085 $Y=1.68
+ $X2=10.085 $Y2=1.44
r103 19 21 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=10.085 $Y=1.68
+ $X2=10.085 $Y2=2.4
r104 15 44 20.5538 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=9.635 $Y=1.68
+ $X2=9.635 $Y2=1.44
r105 15 17 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=9.635 $Y=1.68
+ $X2=9.635 $Y2=2.4
r106 11 40 20.5538 $w=1.8e-07 $l=2.4e-07 $layer=POLY_cond $X=9.185 $Y=1.68
+ $X2=9.185 $Y2=1.44
r107 11 13 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=9.185 $Y=1.68
+ $X2=9.185 $Y2=2.4
r108 7 40 10.0156 $w=3.85e-07 $l=8e-08 $layer=POLY_cond $X=9.105 $Y=1.44
+ $X2=9.185 $Y2=1.44
r109 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.105 $Y=1.35
+ $X2=9.105 $Y2=0.74
r110 5 7 28.0374 $w=3.85e-07 $l=1.98997e-07 $layer=POLY_cond $X=9.03 $Y=1.605
+ $X2=9.105 $Y2=1.44
r111 5 6 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=9.03 $Y=1.605
+ $X2=8.75 $Y2=1.605
r112 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.675 $Y=1.53
+ $X2=8.75 $Y2=1.605
r113 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=8.675 $Y=1.53
+ $X2=8.675 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O311AI_4%VPWR 1 2 3 4 5 6 19 21 27 31 35 37 39 44 45
+ 46 56 64 69 79 88 90 93 97
r112 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r113 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r114 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r115 87 88 13.5255 $w=1.123e-06 $l=1.65e-07 $layer=LI1_cond $X=3.74 $Y=2.852
+ $X2=3.905 $Y2=2.852
r116 84 87 1.51822 $w=1.123e-06 $l=1.4e-07 $layer=LI1_cond $X=3.6 $Y=2.852
+ $X2=3.74 $Y2=2.852
r117 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r118 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r119 81 84 10.4107 $w=1.123e-06 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=2.852
+ $X2=3.6 $Y2=2.852
r120 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r121 78 81 3.09067 $w=1.123e-06 $l=2.85e-07 $layer=LI1_cond $X=2.355 $Y=2.852
+ $X2=2.64 $Y2=2.852
r122 78 79 12.9833 $w=1.123e-06 $l=1.15e-07 $layer=LI1_cond $X=2.355 $Y=2.852
+ $X2=2.24 $Y2=2.852
r123 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r124 73 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r125 73 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r126 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r127 70 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.025 $Y=3.33
+ $X2=9.86 $Y2=3.33
r128 70 72 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.025 $Y=3.33
+ $X2=10.32 $Y2=3.33
r129 69 96 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=10.675 $Y=3.33
+ $X2=10.857 $Y2=3.33
r130 69 72 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=10.675 $Y=3.33
+ $X2=10.32 $Y2=3.33
r131 68 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r132 68 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r133 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r134 65 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.125 $Y=3.33
+ $X2=8.96 $Y2=3.33
r135 65 67 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.125 $Y=3.33
+ $X2=9.36 $Y2=3.33
r136 64 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.695 $Y=3.33
+ $X2=9.86 $Y2=3.33
r137 64 67 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.695 $Y=3.33
+ $X2=9.36 $Y2=3.33
r138 63 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r139 62 63 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r140 60 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r141 59 62 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=8.4 $Y2=3.33
r142 59 88 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=3.905 $Y2=3.33
r143 59 60 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r144 56 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.795 $Y=3.33
+ $X2=8.96 $Y2=3.33
r145 56 62 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=8.795 $Y=3.33
+ $X2=8.4 $Y2=3.33
r146 55 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r147 54 79 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=2.24
+ $Y2=3.33
r148 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r149 51 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r150 51 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r151 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r152 48 75 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r153 48 50 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=1.2 $Y2=3.33
r154 46 63 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=8.4 $Y2=3.33
r155 46 60 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.08 $Y2=3.33
r156 44 50 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r157 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.24 $Y=3.33
+ $X2=1.405 $Y2=3.33
r158 43 54 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.57 $Y=3.33
+ $X2=2.16 $Y2=3.33
r159 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.57 $Y=3.33
+ $X2=1.405 $Y2=3.33
r160 39 42 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=10.8 $Y=1.985
+ $X2=10.8 $Y2=2.815
r161 37 96 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.8 $Y=3.245
+ $X2=10.857 $Y2=3.33
r162 37 42 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.8 $Y=3.245
+ $X2=10.8 $Y2=2.815
r163 33 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.86 $Y=3.245
+ $X2=9.86 $Y2=3.33
r164 33 35 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=9.86 $Y=3.245
+ $X2=9.86 $Y2=2.415
r165 29 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.96 $Y=3.245
+ $X2=8.96 $Y2=3.33
r166 29 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=8.96 $Y=3.245
+ $X2=8.96 $Y2=2.415
r167 25 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.405 $Y=3.245
+ $X2=1.405 $Y2=3.33
r168 25 27 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.405 $Y=3.245
+ $X2=1.405 $Y2=2.455
r169 21 24 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.28 $Y=2.115
+ $X2=0.28 $Y2=2.815
r170 19 75 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r171 19 24 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r172 6 42 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=10.625
+ $Y=1.84 $X2=10.76 $Y2=2.815
r173 6 39 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.625
+ $Y=1.84 $X2=10.76 $Y2=1.985
r174 5 35 300 $w=1.7e-07 $l=6.38944e-07 $layer=licon1_PDIFF $count=2 $X=9.725
+ $Y=1.84 $X2=9.86 $Y2=2.415
r175 4 31 300 $w=1.7e-07 $l=6.43428e-07 $layer=licon1_PDIFF $count=2 $X=8.815
+ $Y=1.84 $X2=8.96 $Y2=2.415
r176 3 87 120 $w=1.7e-07 $l=1.80144e-06 $layer=licon1_PDIFF $count=5 $X=2.22
+ $Y=1.84 $X2=3.74 $Y2=2.455
r177 3 78 120 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=5 $X=2.22
+ $Y=1.84 $X2=2.355 $Y2=2.455
r178 2 27 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.27
+ $Y=1.84 $X2=1.405 $Y2=2.455
r179 1 24 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r180 1 21 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__O311AI_4%Y 1 2 3 4 5 6 23 25 27 29 33 35 39 41 45 51
+ 52 54 56 58 60 61 65 67
c136 45 0 1.61783e-19 $X=6.365 $Y=2.035
r137 65 67 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=6.48 $Y=1.26
+ $X2=6.48 $Y2=1.295
r138 60 65 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.48 $Y=1.175
+ $X2=6.48 $Y2=1.26
r139 60 61 17.2866 $w=2.28e-07 $l=3.45e-07 $layer=LI1_cond $X=6.48 $Y=1.32
+ $X2=6.48 $Y2=1.665
r140 60 67 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=6.48 $Y=1.32
+ $X2=6.48 $Y2=1.295
r141 59 61 14.2803 $w=2.28e-07 $l=2.85e-07 $layer=LI1_cond $X=6.48 $Y=1.95
+ $X2=6.48 $Y2=1.665
r142 50 52 9.45624 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=1.015
+ $X2=1.74 $Y2=1.015
r143 50 51 5.30815 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=1.015
+ $X2=1.41 $Y2=1.015
r144 46 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.015 $Y=2.035
+ $X2=5.85 $Y2=2.035
r145 45 59 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=6.365 $Y=2.035
+ $X2=6.48 $Y2=1.95
r146 45 46 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=6.365 $Y=2.035
+ $X2=6.015 $Y2=2.035
r147 42 56 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=5.015 $Y=2.035
+ $X2=4.85 $Y2=1.97
r148 41 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.685 $Y=2.035
+ $X2=5.85 $Y2=2.035
r149 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.685 $Y=2.035
+ $X2=5.015 $Y2=2.035
r150 37 56 0.89609 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=4.85 $Y=2.12
+ $X2=4.85 $Y2=1.97
r151 37 39 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.85 $Y=2.12
+ $X2=4.85 $Y2=2.31
r152 36 54 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=2.07 $Y=2.035
+ $X2=1.905 $Y2=1.97
r153 35 56 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=4.685 $Y=2.035
+ $X2=4.85 $Y2=1.97
r154 35 36 170.604 $w=1.68e-07 $l=2.615e-06 $layer=LI1_cond $X=4.685 $Y=2.035
+ $X2=2.07 $Y2=2.035
r155 31 54 0.89609 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=1.905 $Y=2.12
+ $X2=1.905 $Y2=1.97
r156 31 33 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.905 $Y=2.12
+ $X2=1.905 $Y2=2.815
r157 29 60 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=6.365 $Y=1.175
+ $X2=6.48 $Y2=1.175
r158 29 52 301.738 $w=1.68e-07 $l=4.625e-06 $layer=LI1_cond $X=6.365 $Y=1.175
+ $X2=1.74 $Y2=1.175
r159 28 48 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.07 $Y=2.035
+ $X2=0.905 $Y2=2.035
r160 27 54 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=1.74 $Y=2.035
+ $X2=1.905 $Y2=1.97
r161 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.74 $Y=2.035
+ $X2=1.07 $Y2=2.035
r162 23 48 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.905 $Y=2.12
+ $X2=0.905 $Y2=2.035
r163 23 25 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.905 $Y=2.12
+ $X2=0.905 $Y2=2.815
r164 21 51 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.71 $Y=0.935
+ $X2=1.41 $Y2=0.935
r165 6 58 300 $w=1.7e-07 $l=3.47851e-07 $layer=licon1_PDIFF $count=2 $X=5.685
+ $Y=1.84 $X2=5.85 $Y2=2.115
r166 5 56 600 $w=1.7e-07 $l=2.41402e-07 $layer=licon1_PDIFF $count=1 $X=4.665
+ $Y=1.84 $X2=4.85 $Y2=1.97
r167 5 39 300 $w=1.7e-07 $l=5.54842e-07 $layer=licon1_PDIFF $count=2 $X=4.665
+ $Y=1.84 $X2=4.85 $Y2=2.31
r168 4 54 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.77
+ $Y=1.84 $X2=1.905 $Y2=1.985
r169 4 33 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.77
+ $Y=1.84 $X2=1.905 $Y2=2.815
r170 3 48 400 $w=1.7e-07 $l=4.25852e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.905 $Y2=2.115
r171 3 25 400 $w=1.7e-07 $l=1.11932e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.905 $Y2=2.815
r172 2 50 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=1.435
+ $Y=0.37 $X2=1.575 $Y2=0.95
r173 1 21 182 $w=1.7e-07 $l=6.3113e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.935
.ends

.subckt PM_SKY130_FD_SC_MS__O311AI_4%A_841_368# 1 2 3 4 5 18 20 21 24 26 30 32
+ 36 38 42 44 45 46
r74 40 42 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=8.4 $Y=2.905 $X2=8.4
+ $Y2=2.415
r75 39 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.615 $Y=2.99
+ $X2=7.45 $Y2=2.99
r76 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.235 $Y=2.99
+ $X2=8.4 $Y2=2.905
r77 38 39 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=8.235 $Y=2.99
+ $X2=7.615 $Y2=2.99
r78 34 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.45 $Y=2.905
+ $X2=7.45 $Y2=2.99
r79 34 36 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=7.45 $Y=2.905
+ $X2=7.45 $Y2=2.455
r80 33 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.615 $Y=2.99
+ $X2=6.45 $Y2=2.99
r81 32 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.285 $Y=2.99
+ $X2=7.45 $Y2=2.99
r82 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.285 $Y=2.99
+ $X2=6.615 $Y2=2.99
r83 28 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.45 $Y=2.905
+ $X2=6.45 $Y2=2.99
r84 28 30 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=6.45 $Y=2.905
+ $X2=6.45 $Y2=2.455
r85 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.515 $Y=2.99
+ $X2=5.35 $Y2=2.99
r86 26 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.285 $Y=2.99
+ $X2=6.45 $Y2=2.99
r87 26 27 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=6.285 $Y=2.99
+ $X2=5.515 $Y2=2.99
r88 22 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.35 $Y=2.905
+ $X2=5.35 $Y2=2.99
r89 22 24 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=5.35 $Y=2.905
+ $X2=5.35 $Y2=2.455
r90 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.185 $Y=2.99
+ $X2=5.35 $Y2=2.99
r91 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.185 $Y=2.99
+ $X2=4.515 $Y2=2.99
r92 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.35 $Y=2.905
+ $X2=4.515 $Y2=2.99
r93 16 18 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.35 $Y=2.905
+ $X2=4.35 $Y2=2.455
r94 5 42 300 $w=1.7e-07 $l=6.38944e-07 $layer=licon1_PDIFF $count=2 $X=8.265
+ $Y=1.84 $X2=8.4 $Y2=2.415
r95 4 36 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=7.265
+ $Y=1.84 $X2=7.45 $Y2=2.455
r96 3 30 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=6.315
+ $Y=1.84 $X2=6.45 $Y2=2.455
r97 2 24 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=5.165
+ $Y=1.84 $X2=5.35 $Y2=2.455
r98 1 18 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=4.205
+ $Y=1.84 $X2=4.35 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__O311AI_4%A_1353_368# 1 2 3 4 15 19 21 25 27 29 31 34
+ 36 38
c55 36 0 9.26431e-20 $X=7.95 $Y=2.035
r56 29 40 2.94404 $w=2.8e-07 $l=1e-07 $layer=LI1_cond $X=10.335 $Y=2.15
+ $X2=10.335 $Y2=2.05
r57 29 31 12.5534 $w=2.78e-07 $l=3.05e-07 $layer=LI1_cond $X=10.335 $Y=2.15
+ $X2=10.335 $Y2=2.455
r58 28 38 5.79383 $w=2e-07 $l=1.15e-07 $layer=LI1_cond $X=9.525 $Y=2.05 $X2=9.41
+ $Y2=2.05
r59 27 40 4.12165 $w=2e-07 $l=1.4e-07 $layer=LI1_cond $X=10.195 $Y=2.05
+ $X2=10.335 $Y2=2.05
r60 27 28 37.1545 $w=1.98e-07 $l=6.7e-07 $layer=LI1_cond $X=10.195 $Y=2.05
+ $X2=9.525 $Y2=2.05
r61 23 38 0.844453 $w=2.3e-07 $l=1e-07 $layer=LI1_cond $X=9.41 $Y=2.15 $X2=9.41
+ $Y2=2.05
r62 23 25 15.2824 $w=2.28e-07 $l=3.05e-07 $layer=LI1_cond $X=9.41 $Y=2.15
+ $X2=9.41 $Y2=2.455
r63 22 36 7.18321 $w=1.85e-07 $l=1.4e-07 $layer=LI1_cond $X=8.065 $Y=2.05
+ $X2=7.925 $Y2=2.05
r64 21 38 5.79383 $w=2e-07 $l=1.15e-07 $layer=LI1_cond $X=9.295 $Y=2.05 $X2=9.41
+ $Y2=2.05
r65 21 22 68.2091 $w=1.98e-07 $l=1.23e-06 $layer=LI1_cond $X=9.295 $Y=2.05
+ $X2=8.065 $Y2=2.05
r66 17 36 0.097681 $w=2.8e-07 $l=1e-07 $layer=LI1_cond $X=7.925 $Y=2.15
+ $X2=7.925 $Y2=2.05
r67 17 19 17.2866 $w=2.78e-07 $l=4.2e-07 $layer=LI1_cond $X=7.925 $Y=2.15
+ $X2=7.925 $Y2=2.57
r68 16 34 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.115 $Y=2.035
+ $X2=6.95 $Y2=2.035
r69 15 36 7.18321 $w=1.85e-07 $l=1.47309e-07 $layer=LI1_cond $X=7.785 $Y=2.035
+ $X2=7.925 $Y2=2.05
r70 15 16 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.785 $Y=2.035
+ $X2=7.115 $Y2=2.035
r71 4 40 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=10.175
+ $Y=1.84 $X2=10.31 $Y2=2.035
r72 4 31 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=10.175
+ $Y=1.84 $X2=10.31 $Y2=2.455
r73 3 38 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=9.275
+ $Y=1.84 $X2=9.41 $Y2=2.035
r74 3 25 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=9.275
+ $Y=1.84 $X2=9.41 $Y2=2.455
r75 2 36 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=7.815
+ $Y=1.84 $X2=7.95 $Y2=2.035
r76 2 19 600 $w=1.7e-07 $l=7.94638e-07 $layer=licon1_PDIFF $count=1 $X=7.815
+ $Y=1.84 $X2=7.95 $Y2=2.57
r77 1 34 300 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=2 $X=6.765
+ $Y=1.84 $X2=6.95 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__O311AI_4%A_27_74# 1 2 3 4 5 16 18 20 28 32
r40 30 32 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=2.865 $Y=0.835
+ $X2=3.735 $Y2=0.835
r41 28 30 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.09 $Y=0.835
+ $X2=2.865 $Y2=0.835
r42 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.005 $Y=0.75
+ $X2=2.09 $Y2=0.835
r43 25 27 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.005 $Y=0.75
+ $X2=2.005 $Y2=0.635
r44 24 27 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.005 $Y=0.6
+ $X2=2.005 $Y2=0.635
r45 21 35 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=0.475
+ $X2=0.24 $Y2=0.475
r46 21 23 35.9562 $w=2.48e-07 $l=7.8e-07 $layer=LI1_cond $X=0.365 $Y=0.475
+ $X2=1.145 $Y2=0.475
r47 20 24 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.92 $Y=0.475
+ $X2=2.005 $Y2=0.6
r48 20 23 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=1.92 $Y=0.475
+ $X2=1.145 $Y2=0.475
r49 16 35 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=0.6 $X2=0.24
+ $Y2=0.475
r50 16 18 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=0.24 $Y=0.6
+ $X2=0.24 $Y2=0.965
r51 5 32 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=3.595
+ $Y=0.37 $X2=3.735 $Y2=0.835
r52 4 30 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=2.725
+ $Y=0.37 $X2=2.865 $Y2=0.835
r53 3 27 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=1.865
+ $Y=0.37 $X2=2.005 $Y2=0.635
r54 2 23 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.37 $X2=1.145 $Y2=0.515
r55 1 35 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
r56 1 18 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_MS__O311AI_4%A_459_74# 1 2 3 4 5 6 7 8 25 32 33 34 37 39
+ 43 45 49 51 55 57 61 64 65 69 71 72 73 76 79
c149 79 0 5.87245e-20 $X=8.85 $Y=1.045
c150 73 0 1.36796e-19 $X=7.015 $Y=0.835
c151 65 0 1.65594e-19 $X=10.165 $Y=1.045
c152 51 0 5.58611e-20 $X=7.945 $Y=1.095
r153 76 77 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=8.03 $Y=1.095
+ $X2=8.03 $Y2=1.385
r154 73 74 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=7.015 $Y=0.835
+ $X2=7.015 $Y2=1.095
r155 67 69 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=10.29 $Y=0.96
+ $X2=10.29 $Y2=0.515
r156 66 79 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.975 $Y=1.045
+ $X2=8.85 $Y2=1.045
r157 65 67 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.165 $Y=1.045
+ $X2=10.29 $Y2=0.96
r158 65 66 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=10.165 $Y=1.045
+ $X2=8.975 $Y2=1.045
r159 63 79 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.85 $Y=1.13
+ $X2=8.85 $Y2=1.045
r160 63 64 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=8.85 $Y=1.13
+ $X2=8.85 $Y2=1.3
r161 59 79 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.85 $Y=0.96
+ $X2=8.85 $Y2=1.045
r162 59 61 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=8.85 $Y=0.96
+ $X2=8.85 $Y2=0.515
r163 58 77 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.115 $Y=1.385
+ $X2=8.03 $Y2=1.385
r164 57 64 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.725 $Y=1.385
+ $X2=8.85 $Y2=1.3
r165 57 58 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=8.725 $Y=1.385
+ $X2=8.115 $Y2=1.385
r166 53 76 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=8.03 $Y=1.01
+ $X2=8.03 $Y2=1.095
r167 53 55 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=8.03 $Y=1.01
+ $X2=8.03 $Y2=0.515
r168 52 74 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.14 $Y=1.095
+ $X2=7.015 $Y2=1.095
r169 51 76 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.945 $Y=1.095
+ $X2=8.03 $Y2=1.095
r170 51 52 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=7.945 $Y=1.095
+ $X2=7.14 $Y2=1.095
r171 47 73 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=7.015 $Y=0.75
+ $X2=7.015 $Y2=0.835
r172 47 49 10.833 $w=2.48e-07 $l=2.35e-07 $layer=LI1_cond $X=7.015 $Y=0.75
+ $X2=7.015 $Y2=0.515
r173 46 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.19 $Y=0.835
+ $X2=6.025 $Y2=0.835
r174 45 73 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.89 $Y=0.835
+ $X2=7.015 $Y2=0.835
r175 45 46 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=6.89 $Y=0.835
+ $X2=6.19 $Y2=0.835
r176 41 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.025 $Y=0.75
+ $X2=6.025 $Y2=0.835
r177 41 43 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=6.025 $Y=0.75
+ $X2=6.025 $Y2=0.635
r178 40 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.17 $Y=0.835
+ $X2=5.045 $Y2=0.835
r179 39 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.86 $Y=0.835
+ $X2=6.025 $Y2=0.835
r180 39 40 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.86 $Y=0.835
+ $X2=5.17 $Y2=0.835
r181 35 71 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=0.75
+ $X2=5.045 $Y2=0.835
r182 35 37 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=5.045 $Y=0.75
+ $X2=5.045 $Y2=0.635
r183 33 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.92 $Y=0.835
+ $X2=5.045 $Y2=0.835
r184 33 34 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.92 $Y=0.835
+ $X2=4.24 $Y2=0.835
r185 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.155 $Y=0.75
+ $X2=4.24 $Y2=0.835
r186 31 32 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.155 $Y=0.58
+ $X2=4.155 $Y2=0.75
r187 27 30 39.8745 $w=2.48e-07 $l=8.65e-07 $layer=LI1_cond $X=2.435 $Y=0.455
+ $X2=3.3 $Y2=0.455
r188 25 31 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.07 $Y=0.455
+ $X2=4.155 $Y2=0.58
r189 25 30 35.4952 $w=2.48e-07 $l=7.7e-07 $layer=LI1_cond $X=4.07 $Y=0.455
+ $X2=3.3 $Y2=0.455
r190 8 69 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=10.175
+ $Y=0.37 $X2=10.33 $Y2=0.515
r191 7 61 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.75
+ $Y=0.37 $X2=8.89 $Y2=0.515
r192 6 55 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=7.815
+ $Y=0.37 $X2=8.03 $Y2=0.515
r193 5 49 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.915
+ $Y=0.37 $X2=7.055 $Y2=0.515
r194 4 43 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=5.885
+ $Y=0.37 $X2=6.025 $Y2=0.635
r195 3 37 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=4.865
+ $Y=0.37 $X2=5.005 $Y2=0.635
r196 2 30 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.155
+ $Y=0.37 $X2=3.3 $Y2=0.495
r197 1 27 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.295
+ $Y=0.37 $X2=2.435 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_MS__O311AI_4%VGND 1 2 3 4 5 6 7 24 28 32 36 40 42 44 46
+ 48 56 61 66 71 81 87 90 93 96 99 104 110 113
r137 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r138 109 110 11.3568 $w=8.73e-07 $l=1.1e-07 $layer=LI1_cond $X=9.885 $Y=0.352
+ $X2=9.995 $Y2=0.352
r139 106 109 0.627429 $w=8.73e-07 $l=4.5e-08 $layer=LI1_cond $X=9.84 $Y=0.352
+ $X2=9.885 $Y2=0.352
r140 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r141 103 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r142 102 106 6.69257 $w=8.73e-07 $l=4.8e-07 $layer=LI1_cond $X=9.36 $Y=0.352
+ $X2=9.84 $Y2=0.352
r143 102 104 12.6814 $w=8.73e-07 $l=2.05e-07 $layer=LI1_cond $X=9.36 $Y=0.352
+ $X2=9.155 $Y2=0.352
r144 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r145 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r146 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r147 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r148 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r149 85 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r150 85 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=9.84 $Y2=0
r151 84 110 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=10.32 $Y=0
+ $X2=9.995 $Y2=0
r152 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r153 81 112 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=10.595 $Y=0
+ $X2=10.817 $Y2=0
r154 81 84 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.595 $Y=0
+ $X2=10.32 $Y2=0
r155 80 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r156 80 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r157 79 104 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.88 $Y=0
+ $X2=9.155 $Y2=0
r158 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r159 77 99 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.545 $Y=0 $X2=8.42
+ $Y2=0
r160 77 79 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=8.545 $Y=0
+ $X2=8.88 $Y2=0
r161 75 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r162 75 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r163 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r164 72 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.65 $Y=0 $X2=7.485
+ $Y2=0
r165 72 74 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.65 $Y=0 $X2=7.92
+ $Y2=0
r166 71 99 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.295 $Y=0 $X2=8.42
+ $Y2=0
r167 71 74 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.295 $Y=0
+ $X2=7.92 $Y2=0
r168 70 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r169 70 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r170 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r171 67 93 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.71 $Y=0 $X2=6.54
+ $Y2=0
r172 67 69 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.71 $Y=0 $X2=6.96
+ $Y2=0
r173 66 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.32 $Y=0 $X2=7.485
+ $Y2=0
r174 66 69 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=7.32 $Y=0 $X2=6.96
+ $Y2=0
r175 65 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r176 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r177 62 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.68 $Y=0 $X2=5.515
+ $Y2=0
r178 62 64 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.68 $Y=0 $X2=6
+ $Y2=0
r179 61 93 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=6.37 $Y=0 $X2=6.54
+ $Y2=0
r180 61 64 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.37 $Y=0 $X2=6
+ $Y2=0
r181 60 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r182 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r183 57 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=4.575
+ $Y2=0
r184 57 59 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=5.04
+ $Y2=0
r185 56 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.35 $Y=0 $X2=5.515
+ $Y2=0
r186 56 59 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.35 $Y=0 $X2=5.04
+ $Y2=0
r187 55 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r188 54 55 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r189 51 55 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=4.08
+ $Y2=0
r190 50 54 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=4.08
+ $Y2=0
r191 50 51 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r192 48 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.41 $Y=0 $X2=4.575
+ $Y2=0
r193 48 54 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.41 $Y=0 $X2=4.08
+ $Y2=0
r194 46 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r195 46 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r196 46 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r197 42 112 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.76 $Y=0.085
+ $X2=10.817 $Y2=0
r198 42 44 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=10.76 $Y=0.085
+ $X2=10.76 $Y2=0.515
r199 38 99 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.42 $Y=0.085
+ $X2=8.42 $Y2=0
r200 38 40 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=8.42 $Y=0.085
+ $X2=8.42 $Y2=0.515
r201 34 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.485 $Y=0.085
+ $X2=7.485 $Y2=0
r202 34 36 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=7.485 $Y=0.085
+ $X2=7.485 $Y2=0.66
r203 30 93 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=6.54 $Y=0.085
+ $X2=6.54 $Y2=0
r204 30 32 11.1855 $w=3.38e-07 $l=3.3e-07 $layer=LI1_cond $X=6.54 $Y=0.085
+ $X2=6.54 $Y2=0.415
r205 26 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.515 $Y=0.085
+ $X2=5.515 $Y2=0
r206 26 28 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=5.515 $Y=0.085
+ $X2=5.515 $Y2=0.415
r207 22 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.575 $Y=0.085
+ $X2=4.575 $Y2=0
r208 22 24 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.575 $Y=0.085
+ $X2=4.575 $Y2=0.495
r209 7 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.62
+ $Y=0.37 $X2=10.76 $Y2=0.515
r210 6 109 91 $w=1.7e-07 $l=8.22679e-07 $layer=licon1_NDIFF $count=2 $X=9.18
+ $Y=0.37 $X2=9.885 $Y2=0.625
r211 5 40 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.32
+ $Y=0.37 $X2=8.46 $Y2=0.515
r212 4 36 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=7.345
+ $Y=0.37 $X2=7.485 $Y2=0.66
r213 3 32 182 $w=1.7e-07 $l=2.46475e-07 $layer=licon1_NDIFF $count=1 $X=6.315
+ $Y=0.37 $X2=6.54 $Y2=0.415
r214 2 28 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=5.295
+ $Y=0.37 $X2=5.515 $Y2=0.415
r215 1 24 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.37 $X2=4.575 $Y2=0.495
.ends


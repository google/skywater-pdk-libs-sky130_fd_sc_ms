* File: sky130_fd_sc_ms__mux2_1.pxi.spice
* Created: Wed Sep  2 12:11:39 2020
* 
x_PM_SKY130_FD_SC_MS__MUX2_1%S N_S_M1003_g N_S_M1006_g N_S_M1011_g N_S_M1008_g
+ N_S_c_78_n N_S_c_79_n N_S_c_80_n S N_S_c_81_n PM_SKY130_FD_SC_MS__MUX2_1%S
x_PM_SKY130_FD_SC_MS__MUX2_1%A1 N_A1_M1007_g N_A1_M1005_g N_A1_c_133_n
+ N_A1_c_146_p N_A1_c_172_p N_A1_c_134_n N_A1_c_135_n A1 A1 N_A1_c_137_n
+ N_A1_c_138_n N_A1_c_162_p PM_SKY130_FD_SC_MS__MUX2_1%A1
x_PM_SKY130_FD_SC_MS__MUX2_1%A0 N_A0_M1000_g N_A0_M1002_g A0 N_A0_c_199_n
+ N_A0_c_200_n PM_SKY130_FD_SC_MS__MUX2_1%A0
x_PM_SKY130_FD_SC_MS__MUX2_1%A_27_112# N_A_27_112#_M1006_s N_A_27_112#_M1003_s
+ N_A_27_112#_M1009_g N_A_27_112#_M1004_g N_A_27_112#_c_231_n
+ N_A_27_112#_c_232_n N_A_27_112#_c_248_n N_A_27_112#_c_239_n
+ N_A_27_112#_c_240_n N_A_27_112#_c_241_n N_A_27_112#_c_233_n
+ N_A_27_112#_c_234_n N_A_27_112#_c_243_n N_A_27_112#_c_235_n
+ N_A_27_112#_c_236_n PM_SKY130_FD_SC_MS__MUX2_1%A_27_112#
x_PM_SKY130_FD_SC_MS__MUX2_1%A_304_74# N_A_304_74#_M1007_d N_A_304_74#_M1000_d
+ N_A_304_74#_M1001_g N_A_304_74#_M1010_g N_A_304_74#_c_325_n
+ N_A_304_74#_c_426_p N_A_304_74#_c_333_n N_A_304_74#_c_339_n
+ N_A_304_74#_c_353_n N_A_304_74#_c_420_p N_A_304_74#_c_360_n
+ N_A_304_74#_c_361_n N_A_304_74#_c_326_n N_A_304_74#_c_327_n
+ N_A_304_74#_c_328_n N_A_304_74#_c_342_n N_A_304_74#_c_329_n
+ N_A_304_74#_c_330_n PM_SKY130_FD_SC_MS__MUX2_1%A_304_74#
x_PM_SKY130_FD_SC_MS__MUX2_1%VPWR N_VPWR_M1003_d N_VPWR_M1004_d N_VPWR_c_433_n
+ N_VPWR_c_434_n N_VPWR_c_435_n N_VPWR_c_436_n VPWR N_VPWR_c_437_n
+ N_VPWR_c_432_n N_VPWR_c_439_n PM_SKY130_FD_SC_MS__MUX2_1%VPWR
x_PM_SKY130_FD_SC_MS__MUX2_1%X N_X_M1010_d N_X_M1001_d N_X_c_479_n N_X_c_480_n X
+ X X N_X_c_483_n N_X_c_481_n X PM_SKY130_FD_SC_MS__MUX2_1%X
x_PM_SKY130_FD_SC_MS__MUX2_1%VGND N_VGND_M1006_d N_VGND_M1009_d N_VGND_c_505_n
+ N_VGND_c_506_n N_VGND_c_507_n N_VGND_c_508_n N_VGND_c_509_n N_VGND_c_510_n
+ VGND N_VGND_c_511_n N_VGND_c_512_n N_VGND_c_513_n N_VGND_c_514_n
+ PM_SKY130_FD_SC_MS__MUX2_1%VGND
cc_1 VNB N_S_M1006_g 0.0307509f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_2 VNB N_S_M1008_g 0.0246926f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=0.74
cc_3 VNB N_S_c_78_n 0.0139974f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.515
cc_4 VNB N_S_c_79_n 0.018548f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=1.515
cc_5 VNB N_S_c_80_n 0.0111302f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.515
cc_6 VNB N_S_c_81_n 0.00177531f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.515
cc_7 VNB N_A1_M1005_g 0.0069771f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_8 VNB N_A1_c_133_n 0.00111648f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.68
cc_9 VNB N_A1_c_134_n 0.0318272f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=0.74
cc_10 VNB N_A1_c_135_n 0.00427166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB A1 0.00811709f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.515
cc_12 VNB N_A1_c_137_n 0.0189248f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.515
cc_13 VNB N_A1_c_138_n 0.0369354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A0_M1000_g 0.00973027f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.26
cc_15 VNB A0 0.00774979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A0_c_199_n 0.0277131f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=2.34
cc_17 VNB N_A0_c_200_n 0.0240239f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.35
cc_18 VNB N_A_27_112#_M1009_g 0.0298799f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.68
cc_19 VNB N_A_27_112#_M1004_g 5.50899e-19 $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.35
cc_20 VNB N_A_27_112#_c_231_n 0.0197085f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.515
cc_21 VNB N_A_27_112#_c_232_n 0.0250637f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.515
cc_22 VNB N_A_27_112#_c_233_n 3.05599e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_112#_c_234_n 0.0116048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_112#_c_235_n 0.00555683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_112#_c_236_n 0.029796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_304_74#_M1001_g 0.00184039f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.68
cc_27 VNB N_A_304_74#_M1010_g 0.0299476f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.35
cc_28 VNB N_A_304_74#_c_325_n 0.00662024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_304_74#_c_326_n 0.00440116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_304_74#_c_327_n 0.00102356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_304_74#_c_328_n 0.00294361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_304_74#_c_329_n 0.00564651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_304_74#_c_330_n 0.0351013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_432_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_X_c_479_n 0.0267746f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=1.68
cc_36 VNB N_X_c_480_n 0.014426f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.35
cc_37 VNB N_X_c_481_n 0.0248128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_505_n 0.0135512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_506_n 0.00191515f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=2.34
cc_40 VNB N_VGND_c_507_n 0.00993982f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=0.74
cc_41 VNB N_VGND_c_508_n 6.638e-19 $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.515
cc_42 VNB N_VGND_c_509_n 0.0585899f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_43 VNB N_VGND_c_510_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_511_n 0.0202692f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.515
cc_45 VNB N_VGND_c_512_n 0.0213848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_513_n 0.261293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_514_n 0.00711965f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VPB N_S_M1003_g 0.0259706f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_49 VPB N_S_M1011_g 0.0247296f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=2.34
cc_50 VPB N_S_c_78_n 8.94354e-19 $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.515
cc_51 VPB N_S_c_79_n 0.00573764f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.515
cc_52 VPB N_S_c_80_n 9.52852e-19 $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.515
cc_53 VPB N_S_c_81_n 0.00328684f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.515
cc_54 VPB N_A1_M1005_g 0.0242173f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.835
cc_55 VPB N_A0_M1000_g 0.0269517f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.26
cc_56 VPB N_A_27_112#_M1004_g 0.0238774f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=1.35
cc_57 VPB N_A_27_112#_c_232_n 0.012642f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.515
cc_58 VPB N_A_27_112#_c_239_n 0.00163287f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.515
cc_59 VPB N_A_27_112#_c_240_n 0.0525944f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_A_27_112#_c_241_n 0.00361889f $X=-0.19 $Y=1.66 $X2=0.67 $Y2=1.665
cc_61 VPB N_A_27_112#_c_233_n 0.00255506f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_62 VPB N_A_27_112#_c_243_n 0.0330491f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_A_304_74#_M1001_g 0.0306626f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.68
cc_64 VPB N_A_304_74#_c_325_n 0.00202686f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_A_304_74#_c_333_n 0.0244417f $X=-0.19 $Y=1.66 $X2=0.95 $Y2=1.515
cc_66 VPB N_VPWR_c_433_n 0.0195076f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=2.34
cc_67 VPB N_VPWR_c_434_n 0.0151577f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=0.74
cc_68 VPB N_VPWR_c_435_n 0.0550508f $X=-0.19 $Y=1.66 $X2=1.04 $Y2=1.515
cc_69 VPB N_VPWR_c_436_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_70 VPB N_VPWR_c_437_n 0.020838f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_432_n 0.0824019f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_439_n 0.0276744f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB X 0.0443119f $X=-0.19 $Y=1.66 $X2=1.055 $Y2=0.74
cc_74 VPB N_X_c_483_n 0.0169891f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_X_c_481_n 0.00782627f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 N_S_M1008_g N_A1_c_133_n 2.24893e-19 $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_77 N_S_M1008_g N_A1_c_134_n 0.0207911f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_78 N_S_M1008_g N_A1_c_135_n 3.74625e-19 $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_79 N_S_M1008_g N_A1_c_137_n 0.0476408f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_80 N_S_M1006_g N_A_27_112#_c_231_n 0.00684278f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_81 N_S_M1006_g N_A_27_112#_c_232_n 0.00602767f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_82 N_S_c_78_n N_A_27_112#_c_232_n 0.0151666f $X=0.505 $Y=1.515 $X2=0 $Y2=0
cc_83 N_S_c_81_n N_A_27_112#_c_232_n 0.026603f $X=0.67 $Y=1.515 $X2=0 $Y2=0
cc_84 N_S_M1003_g N_A_27_112#_c_248_n 0.0153348f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_85 N_S_M1011_g N_A_27_112#_c_248_n 0.0195274f $X=1.04 $Y=2.34 $X2=0 $Y2=0
cc_86 N_S_c_79_n N_A_27_112#_c_248_n 0.00155331f $X=0.95 $Y=1.515 $X2=0 $Y2=0
cc_87 N_S_c_81_n N_A_27_112#_c_248_n 0.0163099f $X=0.67 $Y=1.515 $X2=0 $Y2=0
cc_88 N_S_M1011_g N_A_27_112#_c_239_n 0.0141982f $X=1.04 $Y=2.34 $X2=0 $Y2=0
cc_89 N_S_M1011_g N_A_27_112#_c_241_n 0.00162099f $X=1.04 $Y=2.34 $X2=0 $Y2=0
cc_90 N_S_M1006_g N_A_27_112#_c_234_n 0.00498481f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_91 N_S_c_78_n N_A_27_112#_c_234_n 2.24164e-19 $X=0.505 $Y=1.515 $X2=0 $Y2=0
cc_92 N_S_M1003_g N_A_27_112#_c_243_n 0.013676f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_93 N_S_M1011_g N_A_27_112#_c_243_n 0.00108986f $X=1.04 $Y=2.34 $X2=0 $Y2=0
cc_94 N_S_M1006_g N_A_304_74#_c_325_n 0.00123241f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_95 N_S_M1011_g N_A_304_74#_c_325_n 0.00124168f $X=1.04 $Y=2.34 $X2=0 $Y2=0
cc_96 N_S_M1008_g N_A_304_74#_c_325_n 0.00908273f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_97 N_S_c_80_n N_A_304_74#_c_325_n 0.0108528f $X=1.04 $Y=1.515 $X2=0 $Y2=0
cc_98 N_S_c_81_n N_A_304_74#_c_325_n 0.0265184f $X=0.67 $Y=1.515 $X2=0 $Y2=0
cc_99 N_S_M1003_g N_A_304_74#_c_339_n 6.45041e-19 $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_100 N_S_M1011_g N_A_304_74#_c_339_n 0.0101696f $X=1.04 $Y=2.34 $X2=0 $Y2=0
cc_101 N_S_c_81_n N_A_304_74#_c_339_n 0.00503456f $X=0.67 $Y=1.515 $X2=0 $Y2=0
cc_102 N_S_M1008_g N_A_304_74#_c_342_n 0.00748628f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_103 N_S_M1003_g N_VPWR_c_433_n 0.00480121f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_104 N_S_M1011_g N_VPWR_c_433_n 0.0122409f $X=1.04 $Y=2.34 $X2=0 $Y2=0
cc_105 N_S_M1011_g N_VPWR_c_435_n 0.00492916f $X=1.04 $Y=2.34 $X2=0 $Y2=0
cc_106 N_S_M1003_g N_VPWR_c_432_n 0.00555093f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_107 N_S_M1011_g N_VPWR_c_432_n 0.00511769f $X=1.04 $Y=2.34 $X2=0 $Y2=0
cc_108 N_S_M1003_g N_VPWR_c_439_n 0.00465228f $X=0.505 $Y=2.26 $X2=0 $Y2=0
cc_109 N_S_M1006_g N_VGND_c_505_n 0.00480382f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_110 N_S_M1008_g N_VGND_c_505_n 0.006896f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_111 N_S_M1008_g N_VGND_c_506_n 0.00352246f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_112 N_S_c_79_n N_VGND_c_506_n 0.00133195f $X=0.95 $Y=1.515 $X2=0 $Y2=0
cc_113 N_S_c_81_n N_VGND_c_506_n 0.0147823f $X=0.67 $Y=1.515 $X2=0 $Y2=0
cc_114 N_S_M1008_g N_VGND_c_508_n 0.00308901f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_115 N_S_c_79_n N_VGND_c_508_n 0.00153065f $X=0.95 $Y=1.515 $X2=0 $Y2=0
cc_116 N_S_M1008_g N_VGND_c_509_n 0.00383152f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_117 N_S_M1006_g N_VGND_c_511_n 0.0043356f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_118 N_S_M1006_g N_VGND_c_513_n 0.00487769f $X=0.495 $Y=0.835 $X2=0 $Y2=0
cc_119 N_S_M1008_g N_VGND_c_513_n 0.00384101f $X=1.055 $Y=0.74 $X2=0 $Y2=0
cc_120 N_A1_M1005_g N_A0_M1000_g 0.0332707f $X=2.545 $Y=2.34 $X2=0 $Y2=0
cc_121 N_A1_c_133_n A0 0.00280644f $X=1.6 $Y=1.22 $X2=0 $Y2=0
cc_122 N_A1_c_146_p A0 0.0226197f $X=2.455 $Y=0.895 $X2=0 $Y2=0
cc_123 N_A1_c_134_n A0 4.04959e-19 $X=1.51 $Y=1.385 $X2=0 $Y2=0
cc_124 N_A1_c_135_n A0 0.0235137f $X=1.6 $Y=1.385 $X2=0 $Y2=0
cc_125 A1 A0 0.0285677f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_126 N_A1_c_138_n A0 0.00202561f $X=2.62 $Y=1.385 $X2=0 $Y2=0
cc_127 N_A1_c_146_p N_A0_c_199_n 9.7126e-19 $X=2.455 $Y=0.895 $X2=0 $Y2=0
cc_128 N_A1_c_134_n N_A0_c_199_n 0.0214266f $X=1.51 $Y=1.385 $X2=0 $Y2=0
cc_129 N_A1_c_135_n N_A0_c_199_n 0.00113394f $X=1.6 $Y=1.385 $X2=0 $Y2=0
cc_130 A1 N_A0_c_199_n 3.71725e-19 $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_131 N_A1_c_138_n N_A0_c_199_n 0.0174273f $X=2.62 $Y=1.385 $X2=0 $Y2=0
cc_132 N_A1_c_133_n N_A0_c_200_n 0.00368858f $X=1.6 $Y=1.22 $X2=0 $Y2=0
cc_133 N_A1_c_146_p N_A0_c_200_n 0.013623f $X=2.455 $Y=0.895 $X2=0 $Y2=0
cc_134 A1 N_A0_c_200_n 0.00714134f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_135 N_A1_c_137_n N_A0_c_200_n 0.0195334f $X=1.51 $Y=1.22 $X2=0 $Y2=0
cc_136 A1 N_A_27_112#_M1009_g 0.00411883f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_137 N_A1_c_138_n N_A_27_112#_M1009_g 0.0176872f $X=2.62 $Y=1.385 $X2=0 $Y2=0
cc_138 N_A1_c_162_p N_A_27_112#_M1009_g 0.0011484f $X=2.62 $Y=0.98 $X2=0 $Y2=0
cc_139 N_A1_M1005_g N_A_27_112#_c_240_n 0.0138643f $X=2.545 $Y=2.34 $X2=0 $Y2=0
cc_140 N_A1_M1005_g N_A_27_112#_c_233_n 0.0127496f $X=2.545 $Y=2.34 $X2=0 $Y2=0
cc_141 N_A1_M1005_g N_A_27_112#_c_235_n 0.00213074f $X=2.545 $Y=2.34 $X2=0 $Y2=0
cc_142 A1 N_A_27_112#_c_235_n 0.0184934f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_143 N_A1_c_138_n N_A_27_112#_c_235_n 0.00140853f $X=2.62 $Y=1.385 $X2=0 $Y2=0
cc_144 N_A1_M1005_g N_A_27_112#_c_236_n 0.0382679f $X=2.545 $Y=2.34 $X2=0 $Y2=0
cc_145 A1 N_A_27_112#_c_236_n 2.52902e-19 $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_146 N_A1_c_133_n N_A_304_74#_M1007_d 0.00178335f $X=1.6 $Y=1.22 $X2=-0.19
+ $Y2=-0.245
cc_147 N_A1_c_146_p N_A_304_74#_M1007_d 0.0138145f $X=2.455 $Y=0.895 $X2=-0.19
+ $Y2=-0.245
cc_148 N_A1_c_172_p N_A_304_74#_M1007_d 0.00115008f $X=1.685 $Y=0.895 $X2=-0.19
+ $Y2=-0.245
cc_149 N_A1_c_133_n N_A_304_74#_c_325_n 0.00640423f $X=1.6 $Y=1.22 $X2=0 $Y2=0
cc_150 N_A1_c_134_n N_A_304_74#_c_325_n 9.64054e-19 $X=1.51 $Y=1.385 $X2=0 $Y2=0
cc_151 N_A1_c_135_n N_A_304_74#_c_325_n 0.0248292f $X=1.6 $Y=1.385 $X2=0 $Y2=0
cc_152 N_A1_c_137_n N_A_304_74#_c_325_n 9.75614e-19 $X=1.51 $Y=1.22 $X2=0 $Y2=0
cc_153 N_A1_M1005_g N_A_304_74#_c_333_n 0.00272968f $X=2.545 $Y=2.34 $X2=0 $Y2=0
cc_154 N_A1_c_134_n N_A_304_74#_c_333_n 0.00798977f $X=1.51 $Y=1.385 $X2=0 $Y2=0
cc_155 N_A1_c_135_n N_A_304_74#_c_333_n 0.0255946f $X=1.6 $Y=1.385 $X2=0 $Y2=0
cc_156 N_A1_c_146_p N_A_304_74#_c_353_n 0.0469474f $X=2.455 $Y=0.895 $X2=0 $Y2=0
cc_157 N_A1_c_172_p N_A_304_74#_c_353_n 0.00879433f $X=1.685 $Y=0.895 $X2=0
+ $Y2=0
cc_158 N_A1_c_134_n N_A_304_74#_c_353_n 4.1964e-19 $X=1.51 $Y=1.385 $X2=0 $Y2=0
cc_159 N_A1_c_135_n N_A_304_74#_c_353_n 0.00424542f $X=1.6 $Y=1.385 $X2=0 $Y2=0
cc_160 N_A1_c_137_n N_A_304_74#_c_353_n 0.0157207f $X=1.51 $Y=1.22 $X2=0 $Y2=0
cc_161 N_A1_c_138_n N_A_304_74#_c_353_n 0.00101773f $X=2.62 $Y=1.385 $X2=0 $Y2=0
cc_162 N_A1_c_162_p N_A_304_74#_c_353_n 0.0267499f $X=2.62 $Y=0.98 $X2=0 $Y2=0
cc_163 N_A1_M1005_g N_A_304_74#_c_360_n 0.0120684f $X=2.545 $Y=2.34 $X2=0 $Y2=0
cc_164 N_A1_c_162_p N_A_304_74#_c_361_n 0.0137943f $X=2.62 $Y=0.98 $X2=0 $Y2=0
cc_165 A1 N_A_304_74#_c_327_n 0.0145689f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_166 N_A1_M1005_g N_VPWR_c_435_n 8.71493e-19 $X=2.545 $Y=2.34 $X2=0 $Y2=0
cc_167 N_A1_c_137_n N_VGND_c_505_n 9.47121e-19 $X=1.51 $Y=1.22 $X2=0 $Y2=0
cc_168 N_A1_c_137_n N_VGND_c_509_n 0.00296985f $X=1.51 $Y=1.22 $X2=0 $Y2=0
cc_169 N_A1_c_137_n N_VGND_c_513_n 0.00365796f $X=1.51 $Y=1.22 $X2=0 $Y2=0
cc_170 N_A1_c_146_p A_443_74# 0.00928686f $X=2.455 $Y=0.895 $X2=-0.19 $Y2=-0.245
cc_171 A1 A_443_74# 0.003907f $X=2.555 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_172 N_A1_c_162_p A_443_74# 0.00822687f $X=2.62 $Y=0.98 $X2=-0.19 $Y2=-0.245
cc_173 N_A0_M1000_g N_A_27_112#_c_248_n 0.00457265f $X=2.005 $Y=2.34 $X2=0 $Y2=0
cc_174 N_A0_M1000_g N_A_27_112#_c_239_n 0.015152f $X=2.005 $Y=2.34 $X2=0 $Y2=0
cc_175 N_A0_M1000_g N_A_27_112#_c_240_n 0.0135614f $X=2.005 $Y=2.34 $X2=0 $Y2=0
cc_176 N_A0_M1000_g N_A_304_74#_c_333_n 0.0174093f $X=2.005 $Y=2.34 $X2=0 $Y2=0
cc_177 A0 N_A_304_74#_c_333_n 0.0310181f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_178 N_A0_c_199_n N_A_304_74#_c_333_n 0.0039414f $X=2.05 $Y=1.385 $X2=0 $Y2=0
cc_179 N_A0_c_200_n N_A_304_74#_c_353_n 0.017902f $X=2.05 $Y=1.22 $X2=0 $Y2=0
cc_180 N_A0_M1000_g N_A_304_74#_c_360_n 0.040029f $X=2.005 $Y=2.34 $X2=0 $Y2=0
cc_181 N_A0_M1000_g N_VPWR_c_435_n 8.71493e-19 $X=2.005 $Y=2.34 $X2=0 $Y2=0
cc_182 N_A0_c_200_n N_VGND_c_509_n 0.00296985f $X=2.05 $Y=1.22 $X2=0 $Y2=0
cc_183 N_A0_c_200_n N_VGND_c_513_n 0.00371085f $X=2.05 $Y=1.22 $X2=0 $Y2=0
cc_184 N_A_27_112#_M1004_g N_A_304_74#_M1001_g 0.0161925f $X=3.115 $Y=2.34 $X2=0
+ $Y2=0
cc_185 N_A_27_112#_c_233_n N_A_304_74#_M1001_g 0.00108295f $X=3.04 $Y=2.905
+ $X2=0 $Y2=0
cc_186 N_A_27_112#_c_236_n N_A_304_74#_M1001_g 8.0207e-19 $X=3.19 $Y=1.485 $X2=0
+ $Y2=0
cc_187 N_A_27_112#_M1009_g N_A_304_74#_M1010_g 0.0140133f $X=3.1 $Y=0.74 $X2=0
+ $Y2=0
cc_188 N_A_27_112#_c_248_n N_A_304_74#_c_333_n 0.0108207f $X=1.15 $Y=2.145 $X2=0
+ $Y2=0
cc_189 N_A_27_112#_c_233_n N_A_304_74#_c_333_n 0.00603867f $X=3.04 $Y=2.905
+ $X2=0 $Y2=0
cc_190 N_A_27_112#_c_248_n N_A_304_74#_c_339_n 0.00947979f $X=1.15 $Y=2.145
+ $X2=0 $Y2=0
cc_191 N_A_27_112#_M1009_g N_A_304_74#_c_353_n 0.0110865f $X=3.1 $Y=0.74 $X2=0
+ $Y2=0
cc_192 N_A_27_112#_c_240_n N_A_304_74#_c_360_n 0.0229256f $X=2.955 $Y=2.99 $X2=0
+ $Y2=0
cc_193 N_A_27_112#_c_233_n N_A_304_74#_c_360_n 0.0264417f $X=3.04 $Y=2.905 $X2=0
+ $Y2=0
cc_194 N_A_27_112#_M1009_g N_A_304_74#_c_361_n 0.0123701f $X=3.1 $Y=0.74 $X2=0
+ $Y2=0
cc_195 N_A_27_112#_M1009_g N_A_304_74#_c_326_n 0.00664159f $X=3.1 $Y=0.74 $X2=0
+ $Y2=0
cc_196 N_A_27_112#_c_235_n N_A_304_74#_c_326_n 0.0170649f $X=3.19 $Y=1.485 $X2=0
+ $Y2=0
cc_197 N_A_27_112#_c_236_n N_A_304_74#_c_326_n 0.0041539f $X=3.19 $Y=1.485 $X2=0
+ $Y2=0
cc_198 N_A_27_112#_M1009_g N_A_304_74#_c_327_n 0.00567512f $X=3.1 $Y=0.74 $X2=0
+ $Y2=0
cc_199 N_A_27_112#_c_235_n N_A_304_74#_c_327_n 0.0141748f $X=3.19 $Y=1.485 $X2=0
+ $Y2=0
cc_200 N_A_27_112#_M1009_g N_A_304_74#_c_328_n 0.00279208f $X=3.1 $Y=0.74 $X2=0
+ $Y2=0
cc_201 N_A_27_112#_M1009_g N_A_304_74#_c_329_n 3.83846e-19 $X=3.1 $Y=0.74 $X2=0
+ $Y2=0
cc_202 N_A_27_112#_c_235_n N_A_304_74#_c_329_n 0.0251871f $X=3.19 $Y=1.485 $X2=0
+ $Y2=0
cc_203 N_A_27_112#_c_236_n N_A_304_74#_c_329_n 0.0010311f $X=3.19 $Y=1.485 $X2=0
+ $Y2=0
cc_204 N_A_27_112#_M1009_g N_A_304_74#_c_330_n 5.37584e-19 $X=3.1 $Y=0.74 $X2=0
+ $Y2=0
cc_205 N_A_27_112#_c_235_n N_A_304_74#_c_330_n 3.54107e-19 $X=3.19 $Y=1.485
+ $X2=0 $Y2=0
cc_206 N_A_27_112#_c_236_n N_A_304_74#_c_330_n 0.0201242f $X=3.19 $Y=1.485 $X2=0
+ $Y2=0
cc_207 N_A_27_112#_c_248_n N_VPWR_M1003_d 0.0062813f $X=1.15 $Y=2.145 $X2=-0.19
+ $Y2=-0.245
cc_208 N_A_27_112#_c_248_n N_VPWR_c_433_n 0.0217744f $X=1.15 $Y=2.145 $X2=0
+ $Y2=0
cc_209 N_A_27_112#_c_239_n N_VPWR_c_433_n 0.021319f $X=1.235 $Y=2.905 $X2=0
+ $Y2=0
cc_210 N_A_27_112#_c_241_n N_VPWR_c_433_n 0.0147692f $X=1.32 $Y=2.99 $X2=0 $Y2=0
cc_211 N_A_27_112#_c_243_n N_VPWR_c_433_n 0.0103837f $X=0.28 $Y=2.06 $X2=0 $Y2=0
cc_212 N_A_27_112#_M1004_g N_VPWR_c_434_n 0.010374f $X=3.115 $Y=2.34 $X2=0 $Y2=0
cc_213 N_A_27_112#_c_240_n N_VPWR_c_434_n 0.0147424f $X=2.955 $Y=2.99 $X2=0
+ $Y2=0
cc_214 N_A_27_112#_c_233_n N_VPWR_c_434_n 0.0803761f $X=3.04 $Y=2.905 $X2=0
+ $Y2=0
cc_215 N_A_27_112#_c_235_n N_VPWR_c_434_n 0.00497567f $X=3.19 $Y=1.485 $X2=0
+ $Y2=0
cc_216 N_A_27_112#_c_236_n N_VPWR_c_434_n 0.00137444f $X=3.19 $Y=1.485 $X2=0
+ $Y2=0
cc_217 N_A_27_112#_M1004_g N_VPWR_c_435_n 0.00311838f $X=3.115 $Y=2.34 $X2=0
+ $Y2=0
cc_218 N_A_27_112#_c_240_n N_VPWR_c_435_n 0.117416f $X=2.955 $Y=2.99 $X2=0 $Y2=0
cc_219 N_A_27_112#_c_241_n N_VPWR_c_435_n 0.0121867f $X=1.32 $Y=2.99 $X2=0 $Y2=0
cc_220 N_A_27_112#_M1004_g N_VPWR_c_432_n 0.00271136f $X=3.115 $Y=2.34 $X2=0
+ $Y2=0
cc_221 N_A_27_112#_c_240_n N_VPWR_c_432_n 0.0680683f $X=2.955 $Y=2.99 $X2=0
+ $Y2=0
cc_222 N_A_27_112#_c_241_n N_VPWR_c_432_n 0.00660921f $X=1.32 $Y=2.99 $X2=0
+ $Y2=0
cc_223 N_A_27_112#_c_243_n N_VPWR_c_432_n 0.00995531f $X=0.28 $Y=2.06 $X2=0
+ $Y2=0
cc_224 N_A_27_112#_c_243_n N_VPWR_c_439_n 0.0066444f $X=0.28 $Y=2.06 $X2=0 $Y2=0
cc_225 N_A_27_112#_c_248_n A_226_368# 0.00492277f $X=1.15 $Y=2.145 $X2=-0.19
+ $Y2=-0.245
cc_226 N_A_27_112#_c_239_n A_226_368# 0.0134064f $X=1.235 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_227 N_A_27_112#_c_233_n A_527_368# 0.0145841f $X=3.04 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_228 N_A_27_112#_M1009_g N_X_c_479_n 8.05779e-19 $X=3.1 $Y=0.74 $X2=0 $Y2=0
cc_229 N_A_27_112#_c_234_n N_VGND_c_506_n 0.0112976f $X=0.28 $Y=1.13 $X2=0 $Y2=0
cc_230 N_A_27_112#_M1009_g N_VGND_c_507_n 0.00814582f $X=3.1 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A_27_112#_c_231_n N_VGND_c_508_n 0.0112976f $X=0.28 $Y=0.835 $X2=0
+ $Y2=0
cc_232 N_A_27_112#_M1009_g N_VGND_c_509_n 0.00351724f $X=3.1 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A_27_112#_c_231_n N_VGND_c_511_n 0.0081085f $X=0.28 $Y=0.835 $X2=0
+ $Y2=0
cc_234 N_A_27_112#_M1009_g N_VGND_c_513_n 0.0055287f $X=3.1 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A_27_112#_c_231_n N_VGND_c_513_n 0.010608f $X=0.28 $Y=0.835 $X2=0 $Y2=0
cc_236 N_A_304_74#_M1001_g N_VPWR_c_434_n 0.0057579f $X=3.735 $Y=2.4 $X2=0 $Y2=0
cc_237 N_A_304_74#_c_326_n N_VPWR_c_434_n 0.00547729f $X=3.525 $Y=1.065 $X2=0
+ $Y2=0
cc_238 N_A_304_74#_c_329_n N_VPWR_c_434_n 0.00784726f $X=3.73 $Y=1.465 $X2=0
+ $Y2=0
cc_239 N_A_304_74#_c_330_n N_VPWR_c_434_n 0.0013607f $X=3.73 $Y=1.465 $X2=0
+ $Y2=0
cc_240 N_A_304_74#_M1001_g N_VPWR_c_437_n 0.005209f $X=3.735 $Y=2.4 $X2=0 $Y2=0
cc_241 N_A_304_74#_M1001_g N_VPWR_c_432_n 0.00990716f $X=3.735 $Y=2.4 $X2=0
+ $Y2=0
cc_242 N_A_304_74#_c_333_n A_226_368# 0.0230942f $X=2.065 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_243 N_A_304_74#_M1010_g N_X_c_479_n 0.0105488f $X=3.815 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A_304_74#_M1010_g N_X_c_480_n 0.00309954f $X=3.815 $Y=0.74 $X2=0 $Y2=0
cc_245 N_A_304_74#_c_326_n N_X_c_480_n 0.00664075f $X=3.525 $Y=1.065 $X2=0 $Y2=0
cc_246 N_A_304_74#_c_329_n N_X_c_480_n 0.00233746f $X=3.73 $Y=1.465 $X2=0 $Y2=0
cc_247 N_A_304_74#_M1001_g X 0.0125232f $X=3.735 $Y=2.4 $X2=0 $Y2=0
cc_248 N_A_304_74#_M1001_g N_X_c_483_n 0.00337348f $X=3.735 $Y=2.4 $X2=0 $Y2=0
cc_249 N_A_304_74#_c_329_n N_X_c_483_n 0.00754633f $X=3.73 $Y=1.465 $X2=0 $Y2=0
cc_250 N_A_304_74#_c_330_n N_X_c_483_n 0.00186529f $X=3.73 $Y=1.465 $X2=0 $Y2=0
cc_251 N_A_304_74#_M1001_g N_X_c_481_n 0.00452282f $X=3.735 $Y=2.4 $X2=0 $Y2=0
cc_252 N_A_304_74#_M1010_g N_X_c_481_n 0.00252268f $X=3.815 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A_304_74#_c_328_n N_X_c_481_n 0.005258f $X=3.61 $Y=1.3 $X2=0 $Y2=0
cc_254 N_A_304_74#_c_329_n N_X_c_481_n 0.0249903f $X=3.73 $Y=1.465 $X2=0 $Y2=0
cc_255 N_A_304_74#_c_330_n N_X_c_481_n 0.00231223f $X=3.73 $Y=1.465 $X2=0 $Y2=0
cc_256 N_A_304_74#_c_326_n N_VGND_M1009_d 0.0107009f $X=3.525 $Y=1.065 $X2=0
+ $Y2=0
cc_257 N_A_304_74#_c_325_n N_VGND_c_506_n 0.00787863f $X=1.09 $Y=1.72 $X2=0
+ $Y2=0
cc_258 N_A_304_74#_c_342_n N_VGND_c_506_n 0.0126934f $X=1.26 $Y=0.935 $X2=0
+ $Y2=0
cc_259 N_A_304_74#_M1010_g N_VGND_c_507_n 0.00795549f $X=3.815 $Y=0.74 $X2=0
+ $Y2=0
cc_260 N_A_304_74#_c_353_n N_VGND_c_507_n 0.0206009f $X=2.955 $Y=0.515 $X2=0
+ $Y2=0
cc_261 N_A_304_74#_c_361_n N_VGND_c_507_n 0.0125449f $X=3.04 $Y=0.98 $X2=0 $Y2=0
cc_262 N_A_304_74#_c_326_n N_VGND_c_507_n 0.0270533f $X=3.525 $Y=1.065 $X2=0
+ $Y2=0
cc_263 N_A_304_74#_c_330_n N_VGND_c_507_n 2.35935e-19 $X=3.73 $Y=1.465 $X2=0
+ $Y2=0
cc_264 N_A_304_74#_c_353_n N_VGND_c_509_n 0.0577426f $X=2.955 $Y=0.515 $X2=0
+ $Y2=0
cc_265 N_A_304_74#_c_420_p N_VGND_c_509_n 0.0054507f $X=1.345 $Y=0.515 $X2=0
+ $Y2=0
cc_266 N_A_304_74#_M1010_g N_VGND_c_512_n 0.00434272f $X=3.815 $Y=0.74 $X2=0
+ $Y2=0
cc_267 N_A_304_74#_M1010_g N_VGND_c_513_n 0.00827137f $X=3.815 $Y=0.74 $X2=0
+ $Y2=0
cc_268 N_A_304_74#_c_353_n N_VGND_c_513_n 0.0601803f $X=2.955 $Y=0.515 $X2=0
+ $Y2=0
cc_269 N_A_304_74#_c_420_p N_VGND_c_513_n 0.00604114f $X=1.345 $Y=0.515 $X2=0
+ $Y2=0
cc_270 N_A_304_74#_c_342_n N_VGND_c_513_n 0.00496217f $X=1.26 $Y=0.935 $X2=0
+ $Y2=0
cc_271 N_A_304_74#_c_426_p A_226_74# 3.7257e-19 $X=1.26 $Y=0.85 $X2=-0.19
+ $Y2=-0.245
cc_272 N_A_304_74#_c_420_p A_226_74# 0.00162909f $X=1.345 $Y=0.515 $X2=-0.19
+ $Y2=-0.245
cc_273 N_A_304_74#_c_342_n A_226_74# 0.00520569f $X=1.26 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_274 N_A_304_74#_c_353_n A_443_74# 0.0266902f $X=2.955 $Y=0.515 $X2=-0.19
+ $Y2=-0.245
cc_275 N_A_304_74#_c_361_n A_443_74# 0.00824479f $X=3.04 $Y=0.98 $X2=-0.19
+ $Y2=-0.245
cc_276 N_A_304_74#_c_327_n A_443_74# 0.00144215f $X=3.125 $Y=1.065 $X2=-0.19
+ $Y2=-0.245
cc_277 N_VPWR_c_437_n X 0.0194573f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_278 N_VPWR_c_432_n X 0.0160369f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_279 N_VPWR_c_434_n N_X_c_483_n 0.047026f $X=3.46 $Y=1.985 $X2=0 $Y2=0
cc_280 N_X_c_479_n N_VGND_c_507_n 0.0276686f $X=4.03 $Y=0.515 $X2=0 $Y2=0
cc_281 N_X_c_479_n N_VGND_c_512_n 0.0163488f $X=4.03 $Y=0.515 $X2=0 $Y2=0
cc_282 N_X_c_479_n N_VGND_c_513_n 0.0134757f $X=4.03 $Y=0.515 $X2=0 $Y2=0

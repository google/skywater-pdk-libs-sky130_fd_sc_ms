* File: sky130_fd_sc_ms__nand4bb_4.pxi.spice
* Created: Fri Aug 28 17:46:14 2020
* 
x_PM_SKY130_FD_SC_MS__NAND4BB_4%A_N N_A_N_c_186_n N_A_N_M1015_g N_A_N_M1018_g
+ N_A_N_c_183_n N_A_N_c_188_n N_A_N_M1016_g A_N N_A_N_c_185_n
+ PM_SKY130_FD_SC_MS__NAND4BB_4%A_N
x_PM_SKY130_FD_SC_MS__NAND4BB_4%B_N N_B_N_M1022_g N_B_N_c_230_n N_B_N_c_231_n
+ N_B_N_M1019_g N_B_N_c_234_n N_B_N_M1024_g B_N N_B_N_c_232_n
+ PM_SKY130_FD_SC_MS__NAND4BB_4%B_N
x_PM_SKY130_FD_SC_MS__NAND4BB_4%A_27_114# N_A_27_114#_M1018_s
+ N_A_27_114#_M1015_d N_A_27_114#_c_287_n N_A_27_114#_M1001_g
+ N_A_27_114#_c_303_n N_A_27_114#_M1000_g N_A_27_114#_c_288_n
+ N_A_27_114#_M1007_g N_A_27_114#_c_304_n N_A_27_114#_M1002_g
+ N_A_27_114#_c_289_n N_A_27_114#_M1011_g N_A_27_114#_c_305_n
+ N_A_27_114#_M1003_g N_A_27_114#_M1033_g N_A_27_114#_c_291_n
+ N_A_27_114#_c_292_n N_A_27_114#_c_308_n N_A_27_114#_M1006_g
+ N_A_27_114#_c_293_n N_A_27_114#_c_294_n N_A_27_114#_c_295_n
+ N_A_27_114#_c_310_n N_A_27_114#_c_311_n N_A_27_114#_c_296_n
+ N_A_27_114#_c_312_n N_A_27_114#_c_297_n N_A_27_114#_c_298_n
+ N_A_27_114#_c_299_n N_A_27_114#_c_300_n N_A_27_114#_c_301_n
+ N_A_27_114#_c_302_n PM_SKY130_FD_SC_MS__NAND4BB_4%A_27_114#
x_PM_SKY130_FD_SC_MS__NAND4BB_4%A_232_114# N_A_232_114#_M1022_d
+ N_A_232_114#_M1019_d N_A_232_114#_c_445_n N_A_232_114#_M1004_g
+ N_A_232_114#_c_446_n N_A_232_114#_c_447_n N_A_232_114#_M1010_g
+ N_A_232_114#_c_448_n N_A_232_114#_M1008_g N_A_232_114#_M1013_g
+ N_A_232_114#_c_449_n N_A_232_114#_M1014_g N_A_232_114#_M1017_g
+ N_A_232_114#_c_450_n N_A_232_114#_M1032_g N_A_232_114#_M1020_g
+ N_A_232_114#_c_451_n N_A_232_114#_c_461_n N_A_232_114#_c_462_n
+ N_A_232_114#_c_463_n N_A_232_114#_c_464_n N_A_232_114#_c_465_n
+ N_A_232_114#_c_466_n N_A_232_114#_c_452_n N_A_232_114#_c_453_n
+ N_A_232_114#_c_454_n N_A_232_114#_c_469_n N_A_232_114#_c_455_n
+ PM_SKY130_FD_SC_MS__NAND4BB_4%A_232_114#
x_PM_SKY130_FD_SC_MS__NAND4BB_4%C N_C_M1021_g N_C_M1023_g N_C_M1026_g
+ N_C_M1025_g N_C_M1027_g N_C_M1035_g N_C_M1029_g N_C_M1037_g N_C_c_641_p C
+ N_C_c_628_n N_C_c_629_n N_C_c_634_n PM_SKY130_FD_SC_MS__NAND4BB_4%C
x_PM_SKY130_FD_SC_MS__NAND4BB_4%D N_D_M1028_g N_D_M1005_g N_D_M1009_g
+ N_D_M1030_g N_D_M1012_g N_D_M1031_g N_D_M1036_g N_D_M1034_g D D D D
+ N_D_c_727_n PM_SKY130_FD_SC_MS__NAND4BB_4%D
x_PM_SKY130_FD_SC_MS__NAND4BB_4%VPWR N_VPWR_M1015_s N_VPWR_M1016_s
+ N_VPWR_M1024_s N_VPWR_M1002_d N_VPWR_M1006_d N_VPWR_M1013_s N_VPWR_M1020_s
+ N_VPWR_M1026_s N_VPWR_M1029_s N_VPWR_M1030_s N_VPWR_M1036_s N_VPWR_c_808_n
+ N_VPWR_c_809_n N_VPWR_c_810_n N_VPWR_c_811_n N_VPWR_c_812_n N_VPWR_c_813_n
+ N_VPWR_c_814_n N_VPWR_c_815_n N_VPWR_c_816_n N_VPWR_c_817_n N_VPWR_c_818_n
+ N_VPWR_c_819_n N_VPWR_c_820_n N_VPWR_c_821_n N_VPWR_c_822_n N_VPWR_c_823_n
+ N_VPWR_c_824_n N_VPWR_c_825_n N_VPWR_c_826_n VPWR N_VPWR_c_827_n
+ N_VPWR_c_828_n N_VPWR_c_829_n N_VPWR_c_830_n N_VPWR_c_831_n N_VPWR_c_832_n
+ N_VPWR_c_833_n N_VPWR_c_834_n N_VPWR_c_835_n N_VPWR_c_836_n N_VPWR_c_837_n
+ N_VPWR_c_838_n N_VPWR_c_839_n N_VPWR_c_807_n
+ PM_SKY130_FD_SC_MS__NAND4BB_4%VPWR
x_PM_SKY130_FD_SC_MS__NAND4BB_4%Y N_Y_M1001_s N_Y_M1011_s N_Y_M1000_s
+ N_Y_M1003_s N_Y_M1010_d N_Y_M1017_d N_Y_M1021_d N_Y_M1027_d N_Y_M1028_d
+ N_Y_M1031_d N_Y_c_998_n N_Y_c_1002_n N_Y_c_1168_p N_Y_c_980_n N_Y_c_983_n
+ N_Y_c_1009_n N_Y_c_984_n N_Y_c_1041_n N_Y_c_981_n N_Y_c_986_n N_Y_c_987_n
+ N_Y_c_988_n N_Y_c_1070_n N_Y_c_989_n N_Y_c_1079_n N_Y_c_990_n N_Y_c_1097_n
+ N_Y_c_1101_n N_Y_c_991_n N_Y_c_1010_n N_Y_c_996_n N_Y_c_982_n N_Y_c_1018_n
+ N_Y_c_1019_n N_Y_c_992_n N_Y_c_993_n N_Y_c_994_n N_Y_c_1109_n Y Y
+ PM_SKY130_FD_SC_MS__NAND4BB_4%Y
x_PM_SKY130_FD_SC_MS__NAND4BB_4%VGND N_VGND_M1018_d N_VGND_M1005_s
+ N_VGND_M1012_s N_VGND_c_1179_n N_VGND_c_1180_n N_VGND_c_1181_n VGND
+ N_VGND_c_1182_n N_VGND_c_1183_n N_VGND_c_1184_n N_VGND_c_1185_n
+ N_VGND_c_1186_n N_VGND_c_1187_n N_VGND_c_1188_n N_VGND_c_1189_n
+ PM_SKY130_FD_SC_MS__NAND4BB_4%VGND
x_PM_SKY130_FD_SC_MS__NAND4BB_4%A_374_74# N_A_374_74#_M1001_d
+ N_A_374_74#_M1007_d N_A_374_74#_M1033_d N_A_374_74#_M1008_s
+ N_A_374_74#_M1032_s N_A_374_74#_c_1278_n N_A_374_74#_c_1273_n
+ N_A_374_74#_c_1274_n N_A_374_74#_c_1275_n N_A_374_74#_c_1285_n
+ N_A_374_74#_c_1293_n N_A_374_74#_c_1287_n N_A_374_74#_c_1276_n
+ N_A_374_74#_c_1277_n PM_SKY130_FD_SC_MS__NAND4BB_4%A_374_74#
x_PM_SKY130_FD_SC_MS__NAND4BB_4%A_828_74# N_A_828_74#_M1004_d
+ N_A_828_74#_M1014_d N_A_828_74#_M1023_d N_A_828_74#_M1035_d
+ N_A_828_74#_c_1336_n N_A_828_74#_c_1337_n N_A_828_74#_c_1346_n
+ N_A_828_74#_c_1338_n N_A_828_74#_c_1352_n N_A_828_74#_c_1339_n
+ N_A_828_74#_c_1340_n PM_SKY130_FD_SC_MS__NAND4BB_4%A_828_74#
x_PM_SKY130_FD_SC_MS__NAND4BB_4%A_1229_74# N_A_1229_74#_M1023_s
+ N_A_1229_74#_M1025_s N_A_1229_74#_M1037_s N_A_1229_74#_M1009_d
+ N_A_1229_74#_M1034_d N_A_1229_74#_c_1387_n N_A_1229_74#_c_1388_n
+ N_A_1229_74#_c_1389_n N_A_1229_74#_c_1455_n N_A_1229_74#_c_1390_n
+ N_A_1229_74#_c_1391_n N_A_1229_74#_c_1392_n N_A_1229_74#_c_1393_n
+ N_A_1229_74#_c_1394_n N_A_1229_74#_c_1395_n N_A_1229_74#_c_1396_n
+ N_A_1229_74#_c_1397_n N_A_1229_74#_c_1398_n
+ PM_SKY130_FD_SC_MS__NAND4BB_4%A_1229_74#
cc_1 VNB N_A_N_M1018_g 0.0240966f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.94
cc_2 VNB N_A_N_c_183_n 0.0025227f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.895
cc_3 VNB A_N 0.00259701f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_A_N_c_185_n 0.0198434f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.615
cc_5 VNB N_B_N_M1022_g 0.0287863f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_6 VNB N_B_N_c_230_n 0.0109978f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.94
cc_7 VNB N_B_N_c_231_n 0.0112089f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.94
cc_8 VNB N_B_N_c_232_n 0.0257986f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_9 VNB N_A_27_114#_c_287_n 0.0202274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_114#_c_288_n 0.0171674f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.97
cc_11 VNB N_A_27_114#_c_289_n 0.0162336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_114#_M1033_g 0.0203986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_114#_c_291_n 0.0138726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_114#_c_292_n 0.100033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_114#_c_293_n 0.0152646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_114#_c_294_n 0.0106894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_114#_c_295_n 0.017588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_114#_c_296_n 0.0083148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_114#_c_297_n 0.00921485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_114#_c_298_n 0.00329688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_114#_c_299_n 0.00789124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_114#_c_300_n 0.00448773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_114#_c_301_n 0.00666148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_114#_c_302_n 0.0151117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_232_114#_c_445_n 0.014463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_232_114#_c_446_n 0.0101878f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.045
cc_27 VNB N_A_232_114#_c_447_n 0.00855598f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.54
cc_28 VNB N_A_232_114#_c_448_n 0.01378f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.97
cc_29 VNB N_A_232_114#_c_449_n 0.014886f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.45
cc_30 VNB N_A_232_114#_c_450_n 0.018169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_232_114#_c_451_n 0.00531134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_232_114#_c_452_n 0.00398754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_232_114#_c_453_n 6.33398e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_232_114#_c_454_n 0.00179663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_232_114#_c_455_n 0.10767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_C_M1021_g 4.94619e-19 $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_37 VNB N_C_M1023_g 0.0287149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_C_M1026_g 5.09034e-19 $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.54
cc_39 VNB N_C_M1025_g 0.0209341f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.97
cc_40 VNB N_C_M1027_g 5.09557e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_C_M1035_g 0.0209341f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.45
cc_42 VNB N_C_M1029_g 5.11349e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_C_M1037_g 0.0219074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_C_c_628_n 0.0971162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_C_c_629_n 0.00356294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_D_M1028_g 0.00152838f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_47 VNB N_D_M1005_g 0.0208435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_D_M1009_g 0.0203469f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.54
cc_49 VNB N_D_M1030_g 0.00130001f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.97
cc_50 VNB N_D_M1012_g 0.0212283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_D_M1031_g 0.00130001f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.45
cc_52 VNB N_D_M1036_g 0.0017572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_D_M1034_g 0.0305951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB D 0.0148545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_D_c_727_n 0.110279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VPWR_c_807_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_Y_c_980_n 0.00869888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_Y_c_981_n 0.00429846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_Y_c_982_n 0.00334121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1179_n 0.0215326f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=2.54
cc_61 VNB N_VGND_c_1180_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=0.955 $Y2=1.97
cc_62 VNB N_VGND_c_1181_n 0.00568581f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.615
cc_63 VNB N_VGND_c_1182_n 0.0194575f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.615
cc_64 VNB N_VGND_c_1183_n 0.172757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1184_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1185_n 0.0191515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1186_n 0.536444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1187_n 0.00631593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1188_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1189_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_374_74#_c_1273_n 0.00323114f $X=-0.19 $Y=-0.245 $X2=0.595
+ $Y2=1.615
cc_72 VNB N_A_374_74#_c_1274_n 0.00611261f $X=-0.19 $Y=-0.245 $X2=0.605
+ $Y2=1.615
cc_73 VNB N_A_374_74#_c_1275_n 0.00450137f $X=-0.19 $Y=-0.245 $X2=0.605
+ $Y2=1.615
cc_74 VNB N_A_374_74#_c_1276_n 0.00209585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_374_74#_c_1277_n 0.00332116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_828_74#_c_1336_n 0.00577659f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.97
cc_77 VNB N_A_828_74#_c_1337_n 0.017247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_828_74#_c_1338_n 0.00402487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_828_74#_c_1339_n 0.00129507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_828_74#_c_1340_n 0.00203124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1229_74#_c_1387_n 0.0038712f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_82 VNB N_A_1229_74#_c_1388_n 0.00307486f $X=-0.19 $Y=-0.245 $X2=0.595
+ $Y2=1.615
cc_83 VNB N_A_1229_74#_c_1389_n 0.00477062f $X=-0.19 $Y=-0.245 $X2=0.605
+ $Y2=1.615
cc_84 VNB N_A_1229_74#_c_1390_n 0.00633334f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=1.615
cc_85 VNB N_A_1229_74#_c_1391_n 0.00178889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1229_74#_c_1392_n 0.0042577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1229_74#_c_1393_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1229_74#_c_1394_n 0.0125563f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1229_74#_c_1395_n 0.02581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1229_74#_c_1396_n 0.00124819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1229_74#_c_1397_n 0.00713895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1229_74#_c_1398_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VPB N_A_N_c_186_n 0.0186787f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.045
cc_94 VPB N_A_N_c_183_n 0.0200471f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.895
cc_95 VPB N_A_N_c_188_n 0.047919f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.045
cc_96 VPB A_N 0.00149699f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_97 VPB N_B_N_M1019_g 0.0199302f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.895
cc_98 VPB N_B_N_c_234_n 0.0173724f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.54
cc_99 VPB N_B_N_c_232_n 0.0461188f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_100 VPB N_A_27_114#_c_303_n 0.02081f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.045
cc_101 VPB N_A_27_114#_c_304_n 0.0178085f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=1.97
cc_102 VPB N_A_27_114#_c_305_n 0.017317f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.615
cc_103 VPB N_A_27_114#_c_291_n 0.00600005f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_27_114#_c_292_n 0.0282512f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A_27_114#_c_308_n 0.017335f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_106 VPB N_A_27_114#_c_295_n 0.0137798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB N_A_27_114#_c_310_n 0.00571999f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_27_114#_c_311_n 0.00860392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_27_114#_c_312_n 0.00179594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_110 VPB N_A_232_114#_M1010_g 0.0208888f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB N_A_232_114#_M1013_g 0.0218729f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.615
cc_112 VPB N_A_232_114#_M1017_g 0.0212493f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 VPB N_A_232_114#_M1020_g 0.020719f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_114 VPB N_A_232_114#_c_451_n 0.00641109f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_115 VPB N_A_232_114#_c_461_n 3.95441e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_116 VPB N_A_232_114#_c_462_n 5.2859e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_117 VPB N_A_232_114#_c_463_n 0.00229053f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_A_232_114#_c_464_n 0.00366688f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_119 VPB N_A_232_114#_c_465_n 0.00267055f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_120 VPB N_A_232_114#_c_466_n 0.00310488f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_A_232_114#_c_452_n 0.00224496f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_122 VPB N_A_232_114#_c_453_n 2.94218e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_123 VPB N_A_232_114#_c_469_n 0.00351382f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_232_114#_c_455_n 0.0124461f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_C_M1021_g 0.0227204f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_126 VPB N_C_M1026_g 0.0234354f $X=-0.19 $Y=1.66 $X2=0.955 $Y2=2.54
cc_127 VPB N_C_M1027_g 0.0234552f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_C_M1029_g 0.0234486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_C_c_634_n 0.00441201f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_D_M1028_g 0.023061f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_131 VPB N_D_M1030_g 0.0214385f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.97
cc_132 VPB N_D_M1031_g 0.0214394f $X=-0.19 $Y=1.66 $X2=0.595 $Y2=1.45
cc_133 VPB N_D_M1036_g 0.0259175f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB D 0.0166328f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_808_n 0.0119967f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_809_n 0.0348831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_810_n 0.00272921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_811_n 0.00914439f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_812_n 0.00329129f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_813_n 0.0159425f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_814_n 0.0026822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_815_n 0.0173363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_816_n 0.00489191f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_817_n 0.0048755f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_818_n 0.00969617f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_819_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_820_n 0.00884785f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_821_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_822_n 0.00797179f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_823_n 0.0106521f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_824_n 0.0498587f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_825_n 0.0217466f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_826_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_827_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_828_n 0.0186092f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_829_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_830_n 0.0196495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_831_n 0.0206041f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_832_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_833_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_834_n 0.00600349f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_835_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_836_n 0.00458862f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_837_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_838_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_839_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_807_n 0.0982574f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_Y_c_983_n 0.00249203f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_Y_c_984_n 0.00229053f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_170 VPB N_Y_c_981_n 0.00252167f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_171 VPB N_Y_c_986_n 0.00179594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_Y_c_987_n 0.00990457f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_Y_c_988_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_Y_c_989_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_Y_c_990_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_Y_c_991_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_Y_c_992_n 2.04274e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_Y_c_993_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_Y_c_994_n 0.00244181f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB Y 0.00281363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 N_A_N_M1018_g N_B_N_M1022_g 0.0265012f $X=0.495 $Y=0.94 $X2=0 $Y2=0
cc_182 A_N N_B_N_M1022_g 0.00164408f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_183 N_A_N_c_185_n N_B_N_M1022_g 0.00554618f $X=0.605 $Y=1.615 $X2=0 $Y2=0
cc_184 N_A_N_c_183_n N_B_N_c_231_n 0.00554618f $X=0.595 $Y=1.895 $X2=0 $Y2=0
cc_185 N_A_N_c_188_n N_B_N_c_231_n 0.00259161f $X=0.955 $Y=2.045 $X2=0 $Y2=0
cc_186 N_A_N_c_188_n N_B_N_M1019_g 0.0118391f $X=0.955 $Y=2.045 $X2=0 $Y2=0
cc_187 N_A_N_c_183_n N_B_N_c_232_n 0.00378665f $X=0.595 $Y=1.895 $X2=0 $Y2=0
cc_188 N_A_N_c_188_n N_B_N_c_232_n 0.0118391f $X=0.955 $Y=2.045 $X2=0 $Y2=0
cc_189 N_A_N_M1018_g N_A_27_114#_c_293_n 0.00343265f $X=0.495 $Y=0.94 $X2=0
+ $Y2=0
cc_190 N_A_N_M1018_g N_A_27_114#_c_294_n 0.0059338f $X=0.495 $Y=0.94 $X2=0 $Y2=0
cc_191 N_A_N_M1018_g N_A_27_114#_c_295_n 0.0174929f $X=0.495 $Y=0.94 $X2=0 $Y2=0
cc_192 N_A_N_c_188_n N_A_27_114#_c_295_n 0.00228669f $X=0.955 $Y=2.045 $X2=0
+ $Y2=0
cc_193 A_N N_A_27_114#_c_295_n 0.0250768f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_194 N_A_N_c_186_n N_A_27_114#_c_310_n 0.0104004f $X=0.505 $Y=2.045 $X2=0
+ $Y2=0
cc_195 N_A_N_c_188_n N_A_27_114#_c_310_n 0.0153025f $X=0.955 $Y=2.045 $X2=0
+ $Y2=0
cc_196 A_N N_A_27_114#_c_310_n 0.0283597f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_197 N_A_N_M1018_g N_A_27_114#_c_296_n 0.010552f $X=0.495 $Y=0.94 $X2=0 $Y2=0
cc_198 A_N N_A_27_114#_c_296_n 0.00957008f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_199 N_A_N_c_185_n N_A_27_114#_c_296_n 0.00342578f $X=0.605 $Y=1.615 $X2=0
+ $Y2=0
cc_200 N_A_N_c_186_n N_A_27_114#_c_312_n 8.34606e-19 $X=0.505 $Y=2.045 $X2=0
+ $Y2=0
cc_201 N_A_N_c_188_n N_A_27_114#_c_312_n 8.34606e-19 $X=0.955 $Y=2.045 $X2=0
+ $Y2=0
cc_202 N_A_N_M1018_g N_A_27_114#_c_301_n 0.00422341f $X=0.495 $Y=0.94 $X2=0
+ $Y2=0
cc_203 N_A_N_M1018_g N_A_232_114#_c_451_n 5.52452e-19 $X=0.495 $Y=0.94 $X2=0
+ $Y2=0
cc_204 N_A_N_c_183_n N_A_232_114#_c_451_n 0.00266626f $X=0.595 $Y=1.895 $X2=0
+ $Y2=0
cc_205 N_A_N_c_188_n N_A_232_114#_c_451_n 0.00231886f $X=0.955 $Y=2.045 $X2=0
+ $Y2=0
cc_206 A_N N_A_232_114#_c_451_n 0.0174378f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_207 N_A_N_c_188_n N_A_232_114#_c_462_n 0.00175421f $X=0.955 $Y=2.045 $X2=0
+ $Y2=0
cc_208 N_A_N_M1018_g N_A_232_114#_c_454_n 0.0015097f $X=0.495 $Y=0.94 $X2=0
+ $Y2=0
cc_209 N_A_N_c_186_n N_VPWR_c_809_n 0.013827f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_210 N_A_N_c_188_n N_VPWR_c_809_n 5.41206e-19 $X=0.955 $Y=2.045 $X2=0 $Y2=0
cc_211 N_A_N_c_186_n N_VPWR_c_810_n 5.09586e-19 $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_212 N_A_N_c_188_n N_VPWR_c_810_n 0.0125259f $X=0.955 $Y=2.045 $X2=0 $Y2=0
cc_213 N_A_N_c_186_n N_VPWR_c_827_n 0.00460063f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_214 N_A_N_c_188_n N_VPWR_c_827_n 0.00460063f $X=0.955 $Y=2.045 $X2=0 $Y2=0
cc_215 N_A_N_c_186_n N_VPWR_c_807_n 0.00908554f $X=0.505 $Y=2.045 $X2=0 $Y2=0
cc_216 N_A_N_c_188_n N_VPWR_c_807_n 0.00908554f $X=0.955 $Y=2.045 $X2=0 $Y2=0
cc_217 N_A_N_M1018_g N_VGND_c_1179_n 0.0014541f $X=0.495 $Y=0.94 $X2=0 $Y2=0
cc_218 N_A_N_M1018_g N_VGND_c_1182_n 0.00343632f $X=0.495 $Y=0.94 $X2=0 $Y2=0
cc_219 N_A_N_M1018_g N_VGND_c_1186_n 0.00484898f $X=0.495 $Y=0.94 $X2=0 $Y2=0
cc_220 N_B_N_c_232_n N_A_27_114#_c_303_n 0.0195324f $X=1.63 $Y=1.715 $X2=0 $Y2=0
cc_221 B_N N_A_27_114#_c_292_n 0.00122321f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_222 N_B_N_c_232_n N_A_27_114#_c_292_n 0.00898345f $X=1.63 $Y=1.715 $X2=0
+ $Y2=0
cc_223 N_B_N_M1022_g N_A_27_114#_c_293_n 4.97186e-19 $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_224 N_B_N_M1022_g N_A_27_114#_c_294_n 0.00202668f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_225 N_B_N_M1022_g N_A_27_114#_c_296_n 0.017488f $X=1.085 $Y=0.94 $X2=0 $Y2=0
cc_226 N_B_N_c_232_n N_A_27_114#_c_296_n 0.00428973f $X=1.63 $Y=1.715 $X2=0
+ $Y2=0
cc_227 N_B_N_M1022_g N_A_27_114#_c_297_n 0.00403796f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_228 N_B_N_M1022_g N_A_27_114#_c_298_n 5.59728e-19 $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_229 B_N N_A_27_114#_c_298_n 0.0144744f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_230 N_B_N_c_232_n N_A_27_114#_c_298_n 0.00467287f $X=1.63 $Y=1.715 $X2=0
+ $Y2=0
cc_231 N_B_N_c_232_n N_A_27_114#_c_299_n 3.13473e-19 $X=1.63 $Y=1.715 $X2=0
+ $Y2=0
cc_232 B_N N_A_27_114#_c_302_n 0.00252998f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_233 N_B_N_c_232_n N_A_27_114#_c_302_n 0.00428347f $X=1.63 $Y=1.715 $X2=0
+ $Y2=0
cc_234 N_B_N_M1022_g N_A_232_114#_c_451_n 0.00619912f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_235 N_B_N_c_230_n N_A_232_114#_c_451_n 0.0106382f $X=1.315 $Y=1.58 $X2=0
+ $Y2=0
cc_236 N_B_N_c_231_n N_A_232_114#_c_451_n 0.002803f $X=1.16 $Y=1.58 $X2=0 $Y2=0
cc_237 B_N N_A_232_114#_c_451_n 0.024406f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_238 N_B_N_c_232_n N_A_232_114#_c_451_n 0.00557574f $X=1.63 $Y=1.715 $X2=0
+ $Y2=0
cc_239 N_B_N_c_230_n N_A_232_114#_c_461_n 5.12562e-19 $X=1.315 $Y=1.58 $X2=0
+ $Y2=0
cc_240 N_B_N_M1019_g N_A_232_114#_c_461_n 0.0187465f $X=1.405 $Y=2.54 $X2=0
+ $Y2=0
cc_241 B_N N_A_232_114#_c_461_n 0.0245203f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_242 N_B_N_M1019_g N_A_232_114#_c_463_n 8.86773e-19 $X=1.405 $Y=2.54 $X2=0
+ $Y2=0
cc_243 N_B_N_c_234_n N_A_232_114#_c_463_n 0.0133144f $X=1.855 $Y=2.055 $X2=0
+ $Y2=0
cc_244 N_B_N_c_232_n N_A_232_114#_c_464_n 0.00294147f $X=1.63 $Y=1.715 $X2=0
+ $Y2=0
cc_245 B_N N_A_232_114#_c_466_n 0.0134925f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_246 N_B_N_c_232_n N_A_232_114#_c_466_n 0.00231714f $X=1.63 $Y=1.715 $X2=0
+ $Y2=0
cc_247 N_B_N_M1022_g N_A_232_114#_c_454_n 0.00790561f $X=1.085 $Y=0.94 $X2=0
+ $Y2=0
cc_248 N_B_N_c_230_n N_A_232_114#_c_454_n 0.00604256f $X=1.315 $Y=1.58 $X2=0
+ $Y2=0
cc_249 N_B_N_c_234_n N_A_232_114#_c_469_n 0.0123092f $X=1.855 $Y=2.055 $X2=0
+ $Y2=0
cc_250 N_B_N_c_232_n N_A_232_114#_c_469_n 0.00612003f $X=1.63 $Y=1.715 $X2=0
+ $Y2=0
cc_251 N_B_N_M1019_g N_VPWR_c_810_n 0.0113019f $X=1.405 $Y=2.54 $X2=0 $Y2=0
cc_252 N_B_N_c_234_n N_VPWR_c_810_n 5.70831e-19 $X=1.855 $Y=2.055 $X2=0 $Y2=0
cc_253 N_B_N_c_234_n N_VPWR_c_811_n 0.00864366f $X=1.855 $Y=2.055 $X2=0 $Y2=0
cc_254 N_B_N_M1019_g N_VPWR_c_828_n 0.00460063f $X=1.405 $Y=2.54 $X2=0 $Y2=0
cc_255 N_B_N_c_234_n N_VPWR_c_828_n 0.005209f $X=1.855 $Y=2.055 $X2=0 $Y2=0
cc_256 N_B_N_M1019_g N_VPWR_c_807_n 0.00908554f $X=1.405 $Y=2.54 $X2=0 $Y2=0
cc_257 N_B_N_c_234_n N_VPWR_c_807_n 0.00984635f $X=1.855 $Y=2.055 $X2=0 $Y2=0
cc_258 N_B_N_c_234_n N_Y_c_996_n 2.00118e-19 $X=1.855 $Y=2.055 $X2=0 $Y2=0
cc_259 N_B_N_c_234_n Y 9.16841e-19 $X=1.855 $Y=2.055 $X2=0 $Y2=0
cc_260 N_B_N_M1022_g N_VGND_c_1179_n 0.0014541f $X=1.085 $Y=0.94 $X2=0 $Y2=0
cc_261 N_B_N_M1022_g N_VGND_c_1183_n 0.00344918f $X=1.085 $Y=0.94 $X2=0 $Y2=0
cc_262 N_B_N_M1022_g N_VGND_c_1186_n 0.00484898f $X=1.085 $Y=0.94 $X2=0 $Y2=0
cc_263 N_A_27_114#_c_296_n N_A_232_114#_M1022_d 0.00909254f $X=1.59 $Y=0.745
+ $X2=-0.19 $Y2=-0.245
cc_264 N_A_27_114#_M1033_g N_A_232_114#_c_445_n 0.0160597f $X=3.635 $Y=0.74
+ $X2=0 $Y2=0
cc_265 N_A_27_114#_c_291_n N_A_232_114#_c_447_n 0.00457802f $X=3.885 $Y=1.65
+ $X2=0 $Y2=0
cc_266 N_A_27_114#_c_292_n N_A_232_114#_c_447_n 0.0160597f $X=3.71 $Y=1.65 $X2=0
+ $Y2=0
cc_267 N_A_27_114#_c_308_n N_A_232_114#_M1010_g 0.0197354f $X=3.975 $Y=1.725
+ $X2=0 $Y2=0
cc_268 N_A_27_114#_c_310_n N_A_232_114#_c_451_n 0.00509934f $X=0.645 $Y=2.035
+ $X2=0 $Y2=0
cc_269 N_A_27_114#_c_298_n N_A_232_114#_c_451_n 0.00287569f $X=1.76 $Y=1.295
+ $X2=0 $Y2=0
cc_270 N_A_27_114#_c_310_n N_A_232_114#_c_462_n 0.00428162f $X=0.645 $Y=2.035
+ $X2=0 $Y2=0
cc_271 N_A_27_114#_c_303_n N_A_232_114#_c_463_n 8.20661e-19 $X=2.575 $Y=1.725
+ $X2=0 $Y2=0
cc_272 N_A_27_114#_c_303_n N_A_232_114#_c_464_n 0.00299721f $X=2.575 $Y=1.725
+ $X2=0 $Y2=0
cc_273 N_A_27_114#_c_303_n N_A_232_114#_c_465_n 0.0116769f $X=2.575 $Y=1.725
+ $X2=0 $Y2=0
cc_274 N_A_27_114#_c_304_n N_A_232_114#_c_465_n 0.00928655f $X=3.075 $Y=1.725
+ $X2=0 $Y2=0
cc_275 N_A_27_114#_c_305_n N_A_232_114#_c_465_n 0.00896164f $X=3.525 $Y=1.725
+ $X2=0 $Y2=0
cc_276 N_A_27_114#_c_291_n N_A_232_114#_c_465_n 0.00721007f $X=3.885 $Y=1.65
+ $X2=0 $Y2=0
cc_277 N_A_27_114#_c_292_n N_A_232_114#_c_465_n 0.0404683f $X=3.71 $Y=1.65 $X2=0
+ $Y2=0
cc_278 N_A_27_114#_c_308_n N_A_232_114#_c_465_n 0.0079737f $X=3.975 $Y=1.725
+ $X2=0 $Y2=0
cc_279 N_A_27_114#_c_299_n N_A_232_114#_c_465_n 0.0722626f $X=2.495 $Y=1.38
+ $X2=0 $Y2=0
cc_280 N_A_27_114#_c_302_n N_A_232_114#_c_465_n 8.85762e-19 $X=2.155 $Y=1.38
+ $X2=0 $Y2=0
cc_281 N_A_27_114#_c_302_n N_A_232_114#_c_466_n 0.0083714f $X=2.155 $Y=1.38
+ $X2=0 $Y2=0
cc_282 N_A_27_114#_c_291_n N_A_232_114#_c_452_n 0.00386001f $X=3.885 $Y=1.65
+ $X2=0 $Y2=0
cc_283 N_A_27_114#_c_292_n N_A_232_114#_c_452_n 0.00275733f $X=3.71 $Y=1.65
+ $X2=0 $Y2=0
cc_284 N_A_27_114#_c_296_n N_A_232_114#_c_454_n 0.0179756f $X=1.59 $Y=0.745
+ $X2=0 $Y2=0
cc_285 N_A_27_114#_c_297_n N_A_232_114#_c_454_n 0.0161513f $X=1.675 $Y=1.21
+ $X2=0 $Y2=0
cc_286 N_A_27_114#_c_298_n N_A_232_114#_c_454_n 0.0103428f $X=1.76 $Y=1.295
+ $X2=0 $Y2=0
cc_287 N_A_27_114#_c_303_n N_A_232_114#_c_469_n 0.00165165f $X=2.575 $Y=1.725
+ $X2=0 $Y2=0
cc_288 N_A_27_114#_c_302_n N_A_232_114#_c_469_n 0.0044053f $X=2.155 $Y=1.38
+ $X2=0 $Y2=0
cc_289 N_A_27_114#_c_291_n N_A_232_114#_c_455_n 0.0197354f $X=3.885 $Y=1.65
+ $X2=0 $Y2=0
cc_290 N_A_27_114#_c_292_n N_A_232_114#_c_455_n 0.00500626f $X=3.71 $Y=1.65
+ $X2=0 $Y2=0
cc_291 N_A_27_114#_c_311_n N_VPWR_M1015_s 0.00149394f $X=0.27 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_292 N_A_27_114#_c_310_n N_VPWR_c_809_n 0.0115609f $X=0.645 $Y=2.035 $X2=0
+ $Y2=0
cc_293 N_A_27_114#_c_311_n N_VPWR_c_809_n 0.0139521f $X=0.27 $Y=2.035 $X2=0
+ $Y2=0
cc_294 N_A_27_114#_c_312_n N_VPWR_c_809_n 0.0233699f $X=0.73 $Y=2.265 $X2=0
+ $Y2=0
cc_295 N_A_27_114#_c_312_n N_VPWR_c_810_n 0.0200753f $X=0.73 $Y=2.265 $X2=0
+ $Y2=0
cc_296 N_A_27_114#_c_303_n N_VPWR_c_811_n 0.00822825f $X=2.575 $Y=1.725 $X2=0
+ $Y2=0
cc_297 N_A_27_114#_c_292_n N_VPWR_c_811_n 9.12666e-19 $X=3.71 $Y=1.65 $X2=0
+ $Y2=0
cc_298 N_A_27_114#_c_303_n N_VPWR_c_812_n 6.33086e-19 $X=2.575 $Y=1.725 $X2=0
+ $Y2=0
cc_299 N_A_27_114#_c_304_n N_VPWR_c_812_n 0.0111496f $X=3.075 $Y=1.725 $X2=0
+ $Y2=0
cc_300 N_A_27_114#_c_305_n N_VPWR_c_812_n 0.0109963f $X=3.525 $Y=1.725 $X2=0
+ $Y2=0
cc_301 N_A_27_114#_c_308_n N_VPWR_c_812_n 4.5414e-19 $X=3.975 $Y=1.725 $X2=0
+ $Y2=0
cc_302 N_A_27_114#_c_305_n N_VPWR_c_813_n 0.00460063f $X=3.525 $Y=1.725 $X2=0
+ $Y2=0
cc_303 N_A_27_114#_c_308_n N_VPWR_c_813_n 0.00460063f $X=3.975 $Y=1.725 $X2=0
+ $Y2=0
cc_304 N_A_27_114#_c_305_n N_VPWR_c_814_n 4.5414e-19 $X=3.525 $Y=1.725 $X2=0
+ $Y2=0
cc_305 N_A_27_114#_c_308_n N_VPWR_c_814_n 0.0109666f $X=3.975 $Y=1.725 $X2=0
+ $Y2=0
cc_306 N_A_27_114#_c_303_n N_VPWR_c_825_n 0.00395007f $X=2.575 $Y=1.725 $X2=0
+ $Y2=0
cc_307 N_A_27_114#_c_304_n N_VPWR_c_825_n 0.00460063f $X=3.075 $Y=1.725 $X2=0
+ $Y2=0
cc_308 N_A_27_114#_c_312_n N_VPWR_c_827_n 0.00749631f $X=0.73 $Y=2.265 $X2=0
+ $Y2=0
cc_309 N_A_27_114#_c_303_n N_VPWR_c_807_n 0.00581514f $X=2.575 $Y=1.725 $X2=0
+ $Y2=0
cc_310 N_A_27_114#_c_304_n N_VPWR_c_807_n 0.00909043f $X=3.075 $Y=1.725 $X2=0
+ $Y2=0
cc_311 N_A_27_114#_c_305_n N_VPWR_c_807_n 0.00908554f $X=3.525 $Y=1.725 $X2=0
+ $Y2=0
cc_312 N_A_27_114#_c_308_n N_VPWR_c_807_n 0.00908554f $X=3.975 $Y=1.725 $X2=0
+ $Y2=0
cc_313 N_A_27_114#_c_312_n N_VPWR_c_807_n 0.0062048f $X=0.73 $Y=2.265 $X2=0
+ $Y2=0
cc_314 N_A_27_114#_c_288_n N_Y_c_998_n 0.0108071f $X=2.765 $Y=1.22 $X2=0 $Y2=0
cc_315 N_A_27_114#_c_289_n N_Y_c_998_n 0.0131525f $X=3.205 $Y=1.22 $X2=0 $Y2=0
cc_316 N_A_27_114#_c_292_n N_Y_c_998_n 7.44308e-19 $X=3.71 $Y=1.65 $X2=0 $Y2=0
cc_317 N_A_27_114#_c_300_n N_Y_c_998_n 0.0334364f $X=3 $Y=1.385 $X2=0 $Y2=0
cc_318 N_A_27_114#_c_304_n N_Y_c_1002_n 0.0142562f $X=3.075 $Y=1.725 $X2=0 $Y2=0
cc_319 N_A_27_114#_c_305_n N_Y_c_1002_n 0.0142562f $X=3.525 $Y=1.725 $X2=0 $Y2=0
cc_320 N_A_27_114#_c_292_n N_Y_c_1002_n 4.2073e-19 $X=3.71 $Y=1.65 $X2=0 $Y2=0
cc_321 N_A_27_114#_M1033_g N_Y_c_980_n 0.0126146f $X=3.635 $Y=0.74 $X2=0 $Y2=0
cc_322 N_A_27_114#_c_291_n N_Y_c_980_n 0.00667069f $X=3.885 $Y=1.65 $X2=0 $Y2=0
cc_323 N_A_27_114#_c_305_n N_Y_c_983_n 2.30273e-19 $X=3.525 $Y=1.725 $X2=0 $Y2=0
cc_324 N_A_27_114#_c_308_n N_Y_c_983_n 2.30273e-19 $X=3.975 $Y=1.725 $X2=0 $Y2=0
cc_325 N_A_27_114#_c_308_n N_Y_c_1009_n 0.0142175f $X=3.975 $Y=1.725 $X2=0 $Y2=0
cc_326 N_A_27_114#_c_292_n N_Y_c_1010_n 0.00152107f $X=3.71 $Y=1.65 $X2=0 $Y2=0
cc_327 N_A_27_114#_c_299_n N_Y_c_1010_n 0.0251547f $X=2.495 $Y=1.38 $X2=0 $Y2=0
cc_328 N_A_27_114#_c_303_n N_Y_c_996_n 0.00620796f $X=2.575 $Y=1.725 $X2=0 $Y2=0
cc_329 N_A_27_114#_c_292_n N_Y_c_996_n 7.42431e-19 $X=3.71 $Y=1.65 $X2=0 $Y2=0
cc_330 N_A_27_114#_c_289_n N_Y_c_982_n 0.00303208f $X=3.205 $Y=1.22 $X2=0 $Y2=0
cc_331 N_A_27_114#_M1033_g N_Y_c_982_n 3.32495e-19 $X=3.635 $Y=0.74 $X2=0 $Y2=0
cc_332 N_A_27_114#_c_292_n N_Y_c_982_n 0.0035988f $X=3.71 $Y=1.65 $X2=0 $Y2=0
cc_333 N_A_27_114#_c_300_n N_Y_c_982_n 0.00387326f $X=3 $Y=1.385 $X2=0 $Y2=0
cc_334 N_A_27_114#_c_292_n N_Y_c_1018_n 4.84565e-19 $X=3.71 $Y=1.65 $X2=0 $Y2=0
cc_335 N_A_27_114#_c_308_n N_Y_c_1019_n 8.87219e-19 $X=3.975 $Y=1.725 $X2=0
+ $Y2=0
cc_336 N_A_27_114#_c_303_n Y 0.0182989f $X=2.575 $Y=1.725 $X2=0 $Y2=0
cc_337 N_A_27_114#_c_304_n Y 2.6709e-19 $X=3.075 $Y=1.725 $X2=0 $Y2=0
cc_338 N_A_27_114#_c_296_n N_VGND_M1018_d 0.0124172f $X=1.59 $Y=0.745 $X2=-0.19
+ $Y2=-0.245
cc_339 N_A_27_114#_c_296_n N_VGND_c_1179_n 0.0251972f $X=1.59 $Y=0.745 $X2=0
+ $Y2=0
cc_340 N_A_27_114#_c_293_n N_VGND_c_1182_n 0.00836867f $X=0.272 $Y=0.83 $X2=0
+ $Y2=0
cc_341 N_A_27_114#_c_296_n N_VGND_c_1182_n 0.00241616f $X=1.59 $Y=0.745 $X2=0
+ $Y2=0
cc_342 N_A_27_114#_c_287_n N_VGND_c_1183_n 0.00278271f $X=2.23 $Y=1.22 $X2=0
+ $Y2=0
cc_343 N_A_27_114#_c_288_n N_VGND_c_1183_n 0.00279474f $X=2.765 $Y=1.22 $X2=0
+ $Y2=0
cc_344 N_A_27_114#_c_289_n N_VGND_c_1183_n 0.00279474f $X=3.205 $Y=1.22 $X2=0
+ $Y2=0
cc_345 N_A_27_114#_M1033_g N_VGND_c_1183_n 0.00278247f $X=3.635 $Y=0.74 $X2=0
+ $Y2=0
cc_346 N_A_27_114#_c_296_n N_VGND_c_1183_n 0.012862f $X=1.59 $Y=0.745 $X2=0
+ $Y2=0
cc_347 N_A_27_114#_c_287_n N_VGND_c_1186_n 0.00359383f $X=2.23 $Y=1.22 $X2=0
+ $Y2=0
cc_348 N_A_27_114#_c_288_n N_VGND_c_1186_n 0.00353573f $X=2.765 $Y=1.22 $X2=0
+ $Y2=0
cc_349 N_A_27_114#_c_289_n N_VGND_c_1186_n 0.00352618f $X=3.205 $Y=1.22 $X2=0
+ $Y2=0
cc_350 N_A_27_114#_M1033_g N_VGND_c_1186_n 0.00353524f $X=3.635 $Y=0.74 $X2=0
+ $Y2=0
cc_351 N_A_27_114#_c_293_n N_VGND_c_1186_n 0.0111107f $X=0.272 $Y=0.83 $X2=0
+ $Y2=0
cc_352 N_A_27_114#_c_296_n N_VGND_c_1186_n 0.0290944f $X=1.59 $Y=0.745 $X2=0
+ $Y2=0
cc_353 N_A_27_114#_c_296_n N_A_374_74#_c_1278_n 0.0141315f $X=1.59 $Y=0.745
+ $X2=0 $Y2=0
cc_354 N_A_27_114#_c_297_n N_A_374_74#_c_1278_n 0.015495f $X=1.675 $Y=1.21 $X2=0
+ $Y2=0
cc_355 N_A_27_114#_c_302_n N_A_374_74#_c_1278_n 0.013847f $X=2.155 $Y=1.38 $X2=0
+ $Y2=0
cc_356 N_A_27_114#_c_287_n N_A_374_74#_c_1273_n 0.0144073f $X=2.23 $Y=1.22 $X2=0
+ $Y2=0
cc_357 N_A_27_114#_c_288_n N_A_374_74#_c_1273_n 0.00879331f $X=2.765 $Y=1.22
+ $X2=0 $Y2=0
cc_358 N_A_27_114#_c_289_n N_A_374_74#_c_1275_n 0.00818292f $X=3.205 $Y=1.22
+ $X2=0 $Y2=0
cc_359 N_A_27_114#_M1033_g N_A_374_74#_c_1275_n 0.0102111f $X=3.635 $Y=0.74
+ $X2=0 $Y2=0
cc_360 N_A_27_114#_c_289_n N_A_374_74#_c_1285_n 5.47927e-19 $X=3.205 $Y=1.22
+ $X2=0 $Y2=0
cc_361 N_A_27_114#_M1033_g N_A_374_74#_c_1285_n 0.00468221f $X=3.635 $Y=0.74
+ $X2=0 $Y2=0
cc_362 N_A_27_114#_M1033_g N_A_374_74#_c_1287_n 0.00318514f $X=3.635 $Y=0.74
+ $X2=0 $Y2=0
cc_363 N_A_27_114#_c_287_n N_A_374_74#_c_1276_n 8.87476e-19 $X=2.23 $Y=1.22
+ $X2=0 $Y2=0
cc_364 N_A_27_114#_c_288_n N_A_374_74#_c_1276_n 0.00692257f $X=2.765 $Y=1.22
+ $X2=0 $Y2=0
cc_365 N_A_27_114#_c_289_n N_A_374_74#_c_1276_n 0.00653071f $X=3.205 $Y=1.22
+ $X2=0 $Y2=0
cc_366 N_A_27_114#_M1033_g N_A_374_74#_c_1276_n 6.08651e-19 $X=3.635 $Y=0.74
+ $X2=0 $Y2=0
cc_367 N_A_232_114#_M1020_g N_C_M1021_g 0.0192963f $X=5.825 $Y=2.4 $X2=0 $Y2=0
cc_368 N_A_232_114#_c_455_n N_C_c_628_n 0.0222482f $X=5.515 $Y=1.432 $X2=0 $Y2=0
cc_369 N_A_232_114#_c_455_n N_C_c_629_n 7.93442e-19 $X=5.515 $Y=1.432 $X2=0
+ $Y2=0
cc_370 N_A_232_114#_c_462_n N_VPWR_M1016_s 0.00260941f $X=1.295 $Y=2.135 $X2=0
+ $Y2=0
cc_371 N_A_232_114#_c_465_n N_VPWR_M1024_s 0.00537288f $X=4.145 $Y=1.805 $X2=0
+ $Y2=0
cc_372 N_A_232_114#_c_469_n N_VPWR_M1024_s 0.00274644f $X=2.05 $Y=2.135 $X2=0
+ $Y2=0
cc_373 N_A_232_114#_c_465_n N_VPWR_M1002_d 0.00166235f $X=4.145 $Y=1.805 $X2=0
+ $Y2=0
cc_374 N_A_232_114#_c_465_n N_VPWR_M1006_d 3.61809e-19 $X=4.145 $Y=1.805 $X2=0
+ $Y2=0
cc_375 N_A_232_114#_c_452_n N_VPWR_M1006_d 0.00160304f $X=4.315 $Y=1.555 $X2=0
+ $Y2=0
cc_376 N_A_232_114#_c_461_n N_VPWR_c_810_n 0.00216696f $X=1.515 $Y=2.135 $X2=0
+ $Y2=0
cc_377 N_A_232_114#_c_462_n N_VPWR_c_810_n 0.0119915f $X=1.295 $Y=2.135 $X2=0
+ $Y2=0
cc_378 N_A_232_114#_c_463_n N_VPWR_c_810_n 0.0229093f $X=1.63 $Y=2.265 $X2=0
+ $Y2=0
cc_379 N_A_232_114#_c_463_n N_VPWR_c_811_n 0.0384954f $X=1.63 $Y=2.265 $X2=0
+ $Y2=0
cc_380 N_A_232_114#_c_465_n N_VPWR_c_811_n 0.00739494f $X=4.145 $Y=1.805 $X2=0
+ $Y2=0
cc_381 N_A_232_114#_c_469_n N_VPWR_c_811_n 0.0104953f $X=2.05 $Y=2.135 $X2=0
+ $Y2=0
cc_382 N_A_232_114#_M1010_g N_VPWR_c_814_n 0.0111285f $X=4.425 $Y=2.4 $X2=0
+ $Y2=0
cc_383 N_A_232_114#_M1013_g N_VPWR_c_814_n 4.99912e-19 $X=4.875 $Y=2.4 $X2=0
+ $Y2=0
cc_384 N_A_232_114#_M1010_g N_VPWR_c_815_n 0.00460063f $X=4.425 $Y=2.4 $X2=0
+ $Y2=0
cc_385 N_A_232_114#_M1013_g N_VPWR_c_815_n 0.005209f $X=4.875 $Y=2.4 $X2=0 $Y2=0
cc_386 N_A_232_114#_M1013_g N_VPWR_c_816_n 0.00225515f $X=4.875 $Y=2.4 $X2=0
+ $Y2=0
cc_387 N_A_232_114#_M1017_g N_VPWR_c_816_n 0.0147321f $X=5.375 $Y=2.4 $X2=0
+ $Y2=0
cc_388 N_A_232_114#_M1020_g N_VPWR_c_816_n 5.72826e-19 $X=5.825 $Y=2.4 $X2=0
+ $Y2=0
cc_389 N_A_232_114#_M1017_g N_VPWR_c_817_n 5.84494e-19 $X=5.375 $Y=2.4 $X2=0
+ $Y2=0
cc_390 N_A_232_114#_M1020_g N_VPWR_c_817_n 0.0148399f $X=5.825 $Y=2.4 $X2=0
+ $Y2=0
cc_391 N_A_232_114#_c_463_n N_VPWR_c_828_n 0.0123179f $X=1.63 $Y=2.265 $X2=0
+ $Y2=0
cc_392 N_A_232_114#_M1017_g N_VPWR_c_829_n 0.00460063f $X=5.375 $Y=2.4 $X2=0
+ $Y2=0
cc_393 N_A_232_114#_M1020_g N_VPWR_c_829_n 0.00460063f $X=5.825 $Y=2.4 $X2=0
+ $Y2=0
cc_394 N_A_232_114#_M1010_g N_VPWR_c_807_n 0.00908554f $X=4.425 $Y=2.4 $X2=0
+ $Y2=0
cc_395 N_A_232_114#_M1013_g N_VPWR_c_807_n 0.00982082f $X=4.875 $Y=2.4 $X2=0
+ $Y2=0
cc_396 N_A_232_114#_M1017_g N_VPWR_c_807_n 0.00908554f $X=5.375 $Y=2.4 $X2=0
+ $Y2=0
cc_397 N_A_232_114#_M1020_g N_VPWR_c_807_n 0.00908554f $X=5.825 $Y=2.4 $X2=0
+ $Y2=0
cc_398 N_A_232_114#_c_463_n N_VPWR_c_807_n 0.0101276f $X=1.63 $Y=2.265 $X2=0
+ $Y2=0
cc_399 N_A_232_114#_c_465_n N_Y_M1000_s 0.00218982f $X=4.145 $Y=1.805 $X2=0
+ $Y2=0
cc_400 N_A_232_114#_c_465_n N_Y_M1003_s 0.00165831f $X=4.145 $Y=1.805 $X2=0
+ $Y2=0
cc_401 N_A_232_114#_c_465_n N_Y_c_1002_n 0.0356639f $X=4.145 $Y=1.805 $X2=0
+ $Y2=0
cc_402 N_A_232_114#_c_445_n N_Y_c_980_n 0.00556262f $X=4.065 $Y=1.185 $X2=0
+ $Y2=0
cc_403 N_A_232_114#_c_446_n N_Y_c_980_n 0.00428399f $X=4.335 $Y=1.26 $X2=0 $Y2=0
cc_404 N_A_232_114#_c_447_n N_Y_c_980_n 0.00395324f $X=4.14 $Y=1.26 $X2=0 $Y2=0
cc_405 N_A_232_114#_c_448_n N_Y_c_980_n 0.0055884f $X=4.495 $Y=1.185 $X2=0 $Y2=0
cc_406 N_A_232_114#_c_449_n N_Y_c_980_n 0.00599165f $X=4.925 $Y=1.185 $X2=0
+ $Y2=0
cc_407 N_A_232_114#_c_450_n N_Y_c_980_n 0.00646677f $X=5.515 $Y=1.185 $X2=0
+ $Y2=0
cc_408 N_A_232_114#_c_465_n N_Y_c_980_n 0.0208641f $X=4.145 $Y=1.805 $X2=0 $Y2=0
cc_409 N_A_232_114#_c_452_n N_Y_c_980_n 0.0131063f $X=4.315 $Y=1.555 $X2=0 $Y2=0
cc_410 N_A_232_114#_c_453_n N_Y_c_980_n 0.07199f $X=5.18 $Y=1.515 $X2=0 $Y2=0
cc_411 N_A_232_114#_c_455_n N_Y_c_980_n 0.0340321f $X=5.515 $Y=1.432 $X2=0 $Y2=0
cc_412 N_A_232_114#_M1010_g N_Y_c_1009_n 0.0141904f $X=4.425 $Y=2.4 $X2=0 $Y2=0
cc_413 N_A_232_114#_c_465_n N_Y_c_1009_n 0.0138371f $X=4.145 $Y=1.805 $X2=0
+ $Y2=0
cc_414 N_A_232_114#_c_452_n N_Y_c_1009_n 0.0104056f $X=4.315 $Y=1.555 $X2=0
+ $Y2=0
cc_415 N_A_232_114#_c_453_n N_Y_c_1009_n 0.00594509f $X=5.18 $Y=1.515 $X2=0
+ $Y2=0
cc_416 N_A_232_114#_M1010_g N_Y_c_984_n 2.00987e-19 $X=4.425 $Y=2.4 $X2=0 $Y2=0
cc_417 N_A_232_114#_M1013_g N_Y_c_984_n 0.00899841f $X=4.875 $Y=2.4 $X2=0 $Y2=0
cc_418 N_A_232_114#_M1013_g N_Y_c_1041_n 0.0142696f $X=4.875 $Y=2.4 $X2=0 $Y2=0
cc_419 N_A_232_114#_M1017_g N_Y_c_1041_n 0.0160706f $X=5.375 $Y=2.4 $X2=0 $Y2=0
cc_420 N_A_232_114#_c_453_n N_Y_c_1041_n 0.0336565f $X=5.18 $Y=1.515 $X2=0 $Y2=0
cc_421 N_A_232_114#_c_455_n N_Y_c_1041_n 0.00348259f $X=5.515 $Y=1.432 $X2=0
+ $Y2=0
cc_422 N_A_232_114#_M1017_g N_Y_c_981_n 0.0033441f $X=5.375 $Y=2.4 $X2=0 $Y2=0
cc_423 N_A_232_114#_M1020_g N_Y_c_981_n 0.0033441f $X=5.825 $Y=2.4 $X2=0 $Y2=0
cc_424 N_A_232_114#_c_453_n N_Y_c_981_n 0.0188915f $X=5.18 $Y=1.515 $X2=0 $Y2=0
cc_425 N_A_232_114#_c_455_n N_Y_c_981_n 0.0253204f $X=5.515 $Y=1.432 $X2=0 $Y2=0
cc_426 N_A_232_114#_M1017_g N_Y_c_986_n 3.62369e-19 $X=5.375 $Y=2.4 $X2=0 $Y2=0
cc_427 N_A_232_114#_M1020_g N_Y_c_986_n 3.62369e-19 $X=5.825 $Y=2.4 $X2=0 $Y2=0
cc_428 N_A_232_114#_M1020_g N_Y_c_987_n 0.0191168f $X=5.825 $Y=2.4 $X2=0 $Y2=0
cc_429 N_A_232_114#_M1020_g N_Y_c_988_n 3.09702e-19 $X=5.825 $Y=2.4 $X2=0 $Y2=0
cc_430 N_A_232_114#_c_465_n N_Y_c_996_n 0.0273822f $X=4.145 $Y=1.805 $X2=0 $Y2=0
cc_431 N_A_232_114#_c_469_n N_Y_c_996_n 0.00741551f $X=2.05 $Y=2.135 $X2=0 $Y2=0
cc_432 N_A_232_114#_c_465_n N_Y_c_982_n 0.00644065f $X=4.145 $Y=1.805 $X2=0
+ $Y2=0
cc_433 N_A_232_114#_c_465_n N_Y_c_1018_n 0.0126919f $X=4.145 $Y=1.805 $X2=0
+ $Y2=0
cc_434 N_A_232_114#_M1010_g N_Y_c_1019_n 0.00652852f $X=4.425 $Y=2.4 $X2=0 $Y2=0
cc_435 N_A_232_114#_M1013_g N_Y_c_1019_n 0.00532182f $X=4.875 $Y=2.4 $X2=0 $Y2=0
cc_436 N_A_232_114#_M1017_g N_Y_c_1019_n 0.00103221f $X=5.375 $Y=2.4 $X2=0 $Y2=0
cc_437 N_A_232_114#_c_453_n N_Y_c_1019_n 0.0211111f $X=5.18 $Y=1.515 $X2=0 $Y2=0
cc_438 N_A_232_114#_c_455_n N_Y_c_1019_n 0.00238222f $X=5.515 $Y=1.432 $X2=0
+ $Y2=0
cc_439 N_A_232_114#_M1017_g N_Y_c_992_n 6.10014e-19 $X=5.375 $Y=2.4 $X2=0 $Y2=0
cc_440 N_A_232_114#_M1020_g N_Y_c_993_n 5.23242e-19 $X=5.825 $Y=2.4 $X2=0 $Y2=0
cc_441 N_A_232_114#_c_445_n N_VGND_c_1183_n 0.00328098f $X=4.065 $Y=1.185 $X2=0
+ $Y2=0
cc_442 N_A_232_114#_c_448_n N_VGND_c_1183_n 0.00278271f $X=4.495 $Y=1.185 $X2=0
+ $Y2=0
cc_443 N_A_232_114#_c_449_n N_VGND_c_1183_n 0.00278271f $X=4.925 $Y=1.185 $X2=0
+ $Y2=0
cc_444 N_A_232_114#_c_450_n N_VGND_c_1183_n 0.00278271f $X=5.515 $Y=1.185 $X2=0
+ $Y2=0
cc_445 N_A_232_114#_c_445_n N_VGND_c_1186_n 0.00427409f $X=4.065 $Y=1.185 $X2=0
+ $Y2=0
cc_446 N_A_232_114#_c_448_n N_VGND_c_1186_n 0.00353428f $X=4.495 $Y=1.185 $X2=0
+ $Y2=0
cc_447 N_A_232_114#_c_449_n N_VGND_c_1186_n 0.00354813f $X=4.925 $Y=1.185 $X2=0
+ $Y2=0
cc_448 N_A_232_114#_c_450_n N_VGND_c_1186_n 0.00358903f $X=5.515 $Y=1.185 $X2=0
+ $Y2=0
cc_449 N_A_232_114#_c_445_n N_A_374_74#_c_1275_n 0.00120172f $X=4.065 $Y=1.185
+ $X2=0 $Y2=0
cc_450 N_A_232_114#_c_445_n N_A_374_74#_c_1293_n 0.0108788f $X=4.065 $Y=1.185
+ $X2=0 $Y2=0
cc_451 N_A_232_114#_c_446_n N_A_374_74#_c_1293_n 5.58977e-19 $X=4.335 $Y=1.26
+ $X2=0 $Y2=0
cc_452 N_A_232_114#_c_448_n N_A_374_74#_c_1293_n 0.00843174f $X=4.495 $Y=1.185
+ $X2=0 $Y2=0
cc_453 N_A_232_114#_c_449_n N_A_374_74#_c_1293_n 0.00923324f $X=4.925 $Y=1.185
+ $X2=0 $Y2=0
cc_454 N_A_232_114#_c_450_n N_A_374_74#_c_1293_n 0.00943004f $X=5.515 $Y=1.185
+ $X2=0 $Y2=0
cc_455 N_A_232_114#_c_455_n N_A_374_74#_c_1293_n 0.00196488f $X=5.515 $Y=1.432
+ $X2=0 $Y2=0
cc_456 N_A_232_114#_c_449_n N_A_374_74#_c_1277_n 7.8181e-19 $X=4.925 $Y=1.185
+ $X2=0 $Y2=0
cc_457 N_A_232_114#_c_450_n N_A_374_74#_c_1277_n 0.00496352f $X=5.515 $Y=1.185
+ $X2=0 $Y2=0
cc_458 N_A_232_114#_c_455_n N_A_374_74#_c_1277_n 0.00611361f $X=5.515 $Y=1.432
+ $X2=0 $Y2=0
cc_459 N_A_232_114#_c_445_n N_A_828_74#_c_1336_n 0.00517186f $X=4.065 $Y=1.185
+ $X2=0 $Y2=0
cc_460 N_A_232_114#_c_448_n N_A_828_74#_c_1336_n 0.0125961f $X=4.495 $Y=1.185
+ $X2=0 $Y2=0
cc_461 N_A_232_114#_c_449_n N_A_828_74#_c_1336_n 0.0163854f $X=4.925 $Y=1.185
+ $X2=0 $Y2=0
cc_462 N_A_232_114#_c_450_n N_A_828_74#_c_1337_n 0.012738f $X=5.515 $Y=1.185
+ $X2=0 $Y2=0
cc_463 N_A_232_114#_c_450_n N_A_1229_74#_c_1387_n 0.00200707f $X=5.515 $Y=1.185
+ $X2=0 $Y2=0
cc_464 N_A_232_114#_c_450_n N_A_1229_74#_c_1389_n 0.00344265f $X=5.515 $Y=1.185
+ $X2=0 $Y2=0
cc_465 N_C_M1029_g N_D_M1028_g 0.0177037f $X=7.725 $Y=2.4 $X2=0 $Y2=0
cc_466 N_C_M1037_g N_D_M1005_g 0.0127894f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_467 N_C_M1037_g D 7.06418e-19 $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_468 N_C_c_641_p D 0.00893486f $X=7.445 $Y=1.485 $X2=0 $Y2=0
cc_469 N_C_c_628_n D 0.00134811f $X=7.725 $Y=1.485 $X2=0 $Y2=0
cc_470 N_C_c_641_p N_D_c_727_n 0.00107913f $X=7.445 $Y=1.485 $X2=0 $Y2=0
cc_471 N_C_c_628_n N_D_c_727_n 0.0309149f $X=7.725 $Y=1.485 $X2=0 $Y2=0
cc_472 N_C_M1021_g N_VPWR_c_817_n 0.0034083f $X=6.275 $Y=2.4 $X2=0 $Y2=0
cc_473 N_C_M1026_g N_VPWR_c_818_n 0.00343717f $X=6.725 $Y=2.4 $X2=0 $Y2=0
cc_474 N_C_M1027_g N_VPWR_c_818_n 0.00343717f $X=7.275 $Y=2.4 $X2=0 $Y2=0
cc_475 N_C_M1027_g N_VPWR_c_819_n 0.005209f $X=7.275 $Y=2.4 $X2=0 $Y2=0
cc_476 N_C_M1029_g N_VPWR_c_819_n 0.005209f $X=7.725 $Y=2.4 $X2=0 $Y2=0
cc_477 N_C_M1029_g N_VPWR_c_820_n 0.00306788f $X=7.725 $Y=2.4 $X2=0 $Y2=0
cc_478 N_C_M1021_g N_VPWR_c_830_n 0.005209f $X=6.275 $Y=2.4 $X2=0 $Y2=0
cc_479 N_C_M1026_g N_VPWR_c_830_n 0.005209f $X=6.725 $Y=2.4 $X2=0 $Y2=0
cc_480 N_C_M1021_g N_VPWR_c_807_n 0.00982376f $X=6.275 $Y=2.4 $X2=0 $Y2=0
cc_481 N_C_M1026_g N_VPWR_c_807_n 0.00982526f $X=6.725 $Y=2.4 $X2=0 $Y2=0
cc_482 N_C_M1027_g N_VPWR_c_807_n 0.00982526f $X=7.275 $Y=2.4 $X2=0 $Y2=0
cc_483 N_C_M1029_g N_VPWR_c_807_n 0.00982832f $X=7.725 $Y=2.4 $X2=0 $Y2=0
cc_484 N_C_c_628_n N_Y_c_981_n 0.00103833f $X=7.725 $Y=1.485 $X2=0 $Y2=0
cc_485 N_C_c_629_n N_Y_c_981_n 0.0111225f $X=6.845 $Y=1.55 $X2=0 $Y2=0
cc_486 N_C_M1021_g N_Y_c_987_n 0.0138326f $X=6.275 $Y=2.4 $X2=0 $Y2=0
cc_487 N_C_c_629_n N_Y_c_987_n 0.0107119f $X=6.845 $Y=1.55 $X2=0 $Y2=0
cc_488 N_C_M1021_g N_Y_c_988_n 0.0116208f $X=6.275 $Y=2.4 $X2=0 $Y2=0
cc_489 N_C_M1026_g N_Y_c_988_n 0.0125032f $X=6.725 $Y=2.4 $X2=0 $Y2=0
cc_490 N_C_M1026_g N_Y_c_1070_n 0.0151658f $X=6.725 $Y=2.4 $X2=0 $Y2=0
cc_491 N_C_M1027_g N_Y_c_1070_n 0.0142205f $X=7.275 $Y=2.4 $X2=0 $Y2=0
cc_492 N_C_c_641_p N_Y_c_1070_n 0.0106446f $X=7.445 $Y=1.485 $X2=0 $Y2=0
cc_493 N_C_c_628_n N_Y_c_1070_n 0.00133381f $X=7.725 $Y=1.485 $X2=0 $Y2=0
cc_494 N_C_c_629_n N_Y_c_1070_n 0.00749244f $X=6.845 $Y=1.55 $X2=0 $Y2=0
cc_495 N_C_c_634_n N_Y_c_1070_n 0.0174412f $X=7.075 $Y=1.55 $X2=0 $Y2=0
cc_496 N_C_M1026_g N_Y_c_989_n 6.00071e-19 $X=6.725 $Y=2.4 $X2=0 $Y2=0
cc_497 N_C_M1027_g N_Y_c_989_n 0.0125032f $X=7.275 $Y=2.4 $X2=0 $Y2=0
cc_498 N_C_M1029_g N_Y_c_989_n 0.0127647f $X=7.725 $Y=2.4 $X2=0 $Y2=0
cc_499 N_C_M1029_g N_Y_c_1079_n 0.017729f $X=7.725 $Y=2.4 $X2=0 $Y2=0
cc_500 N_C_M1029_g N_Y_c_990_n 6.10838e-19 $X=7.725 $Y=2.4 $X2=0 $Y2=0
cc_501 N_C_M1021_g N_Y_c_993_n 0.00424108f $X=6.275 $Y=2.4 $X2=0 $Y2=0
cc_502 N_C_M1026_g N_Y_c_993_n 0.00434937f $X=6.725 $Y=2.4 $X2=0 $Y2=0
cc_503 N_C_M1027_g N_Y_c_993_n 0.00108519f $X=7.275 $Y=2.4 $X2=0 $Y2=0
cc_504 N_C_c_628_n N_Y_c_993_n 0.00245159f $X=7.725 $Y=1.485 $X2=0 $Y2=0
cc_505 N_C_c_629_n N_Y_c_993_n 0.0274034f $X=6.845 $Y=1.55 $X2=0 $Y2=0
cc_506 N_C_M1026_g N_Y_c_994_n 4.03257e-19 $X=6.725 $Y=2.4 $X2=0 $Y2=0
cc_507 N_C_M1027_g N_Y_c_994_n 0.00388509f $X=7.275 $Y=2.4 $X2=0 $Y2=0
cc_508 N_C_M1029_g N_Y_c_994_n 0.00419881f $X=7.725 $Y=2.4 $X2=0 $Y2=0
cc_509 N_C_c_641_p N_Y_c_994_n 0.0230595f $X=7.445 $Y=1.485 $X2=0 $Y2=0
cc_510 N_C_c_628_n N_Y_c_994_n 0.00239242f $X=7.725 $Y=1.485 $X2=0 $Y2=0
cc_511 N_C_M1037_g N_VGND_c_1180_n 4.98172e-19 $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_512 N_C_M1023_g N_VGND_c_1183_n 0.00278247f $X=6.505 $Y=0.74 $X2=0 $Y2=0
cc_513 N_C_M1025_g N_VGND_c_1183_n 0.00278247f $X=6.935 $Y=0.74 $X2=0 $Y2=0
cc_514 N_C_M1035_g N_VGND_c_1183_n 0.00278247f $X=7.365 $Y=0.74 $X2=0 $Y2=0
cc_515 N_C_M1037_g N_VGND_c_1183_n 0.00430908f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_516 N_C_M1023_g N_VGND_c_1186_n 0.00358425f $X=6.505 $Y=0.74 $X2=0 $Y2=0
cc_517 N_C_M1025_g N_VGND_c_1186_n 0.00353427f $X=6.935 $Y=0.74 $X2=0 $Y2=0
cc_518 N_C_M1035_g N_VGND_c_1186_n 0.00353427f $X=7.365 $Y=0.74 $X2=0 $Y2=0
cc_519 N_C_M1037_g N_VGND_c_1186_n 0.00816766f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_520 N_C_M1023_g N_A_828_74#_c_1337_n 0.00987533f $X=6.505 $Y=0.74 $X2=0 $Y2=0
cc_521 N_C_M1023_g N_A_828_74#_c_1346_n 0.0104366f $X=6.505 $Y=0.74 $X2=0 $Y2=0
cc_522 N_C_M1025_g N_A_828_74#_c_1346_n 0.00593684f $X=6.935 $Y=0.74 $X2=0 $Y2=0
cc_523 N_C_M1035_g N_A_828_74#_c_1346_n 5.63827e-19 $X=7.365 $Y=0.74 $X2=0 $Y2=0
cc_524 N_C_M1025_g N_A_828_74#_c_1338_n 0.00783479f $X=6.935 $Y=0.74 $X2=0 $Y2=0
cc_525 N_C_M1035_g N_A_828_74#_c_1338_n 0.00990232f $X=7.365 $Y=0.74 $X2=0 $Y2=0
cc_526 N_C_M1037_g N_A_828_74#_c_1338_n 0.00412426f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_527 N_C_M1025_g N_A_828_74#_c_1352_n 5.63827e-19 $X=6.935 $Y=0.74 $X2=0 $Y2=0
cc_528 N_C_M1035_g N_A_828_74#_c_1352_n 0.00593684f $X=7.365 $Y=0.74 $X2=0 $Y2=0
cc_529 N_C_M1037_g N_A_828_74#_c_1352_n 0.00473467f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_530 N_C_M1023_g N_A_828_74#_c_1340_n 0.00206753f $X=6.505 $Y=0.74 $X2=0 $Y2=0
cc_531 N_C_M1025_g N_A_828_74#_c_1340_n 0.00206753f $X=6.935 $Y=0.74 $X2=0 $Y2=0
cc_532 N_C_M1023_g N_A_1229_74#_c_1388_n 0.0119006f $X=6.505 $Y=0.74 $X2=0 $Y2=0
cc_533 N_C_M1025_g N_A_1229_74#_c_1388_n 0.0111242f $X=6.935 $Y=0.74 $X2=0 $Y2=0
cc_534 N_C_c_628_n N_A_1229_74#_c_1388_n 0.00408368f $X=7.725 $Y=1.485 $X2=0
+ $Y2=0
cc_535 N_C_c_629_n N_A_1229_74#_c_1388_n 0.0510561f $X=6.845 $Y=1.55 $X2=0 $Y2=0
cc_536 N_C_c_628_n N_A_1229_74#_c_1389_n 0.00514237f $X=7.725 $Y=1.485 $X2=0
+ $Y2=0
cc_537 N_C_c_629_n N_A_1229_74#_c_1389_n 0.0157582f $X=6.845 $Y=1.55 $X2=0 $Y2=0
cc_538 N_C_M1035_g N_A_1229_74#_c_1390_n 0.011119f $X=7.365 $Y=0.74 $X2=0 $Y2=0
cc_539 N_C_M1037_g N_A_1229_74#_c_1390_n 0.0170327f $X=7.795 $Y=0.74 $X2=0 $Y2=0
cc_540 N_C_c_641_p N_A_1229_74#_c_1390_n 0.0275868f $X=7.445 $Y=1.485 $X2=0
+ $Y2=0
cc_541 N_C_c_628_n N_A_1229_74#_c_1390_n 0.00267527f $X=7.725 $Y=1.485 $X2=0
+ $Y2=0
cc_542 N_C_M1037_g N_A_1229_74#_c_1391_n 3.92031e-19 $X=7.795 $Y=0.74 $X2=0
+ $Y2=0
cc_543 N_C_c_628_n N_A_1229_74#_c_1396_n 0.00270642f $X=7.725 $Y=1.485 $X2=0
+ $Y2=0
cc_544 N_C_c_634_n N_A_1229_74#_c_1396_n 0.0140843f $X=7.075 $Y=1.55 $X2=0 $Y2=0
cc_545 N_D_M1028_g N_VPWR_c_820_n 0.00318542f $X=8.225 $Y=2.4 $X2=0 $Y2=0
cc_546 N_D_M1028_g N_VPWR_c_821_n 0.005209f $X=8.225 $Y=2.4 $X2=0 $Y2=0
cc_547 N_D_M1030_g N_VPWR_c_821_n 0.005209f $X=8.675 $Y=2.4 $X2=0 $Y2=0
cc_548 N_D_M1030_g N_VPWR_c_822_n 0.0027763f $X=8.675 $Y=2.4 $X2=0 $Y2=0
cc_549 N_D_M1031_g N_VPWR_c_822_n 0.0027763f $X=9.125 $Y=2.4 $X2=0 $Y2=0
cc_550 N_D_M1036_g N_VPWR_c_824_n 0.00501904f $X=9.575 $Y=2.4 $X2=0 $Y2=0
cc_551 D N_VPWR_c_824_n 0.0210496f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_552 N_D_c_727_n N_VPWR_c_824_n 0.00117022f $X=9.585 $Y=1.465 $X2=0 $Y2=0
cc_553 N_D_M1031_g N_VPWR_c_831_n 0.005209f $X=9.125 $Y=2.4 $X2=0 $Y2=0
cc_554 N_D_M1036_g N_VPWR_c_831_n 0.005209f $X=9.575 $Y=2.4 $X2=0 $Y2=0
cc_555 N_D_M1028_g N_VPWR_c_807_n 0.0098216f $X=8.225 $Y=2.4 $X2=0 $Y2=0
cc_556 N_D_M1030_g N_VPWR_c_807_n 0.00982266f $X=8.675 $Y=2.4 $X2=0 $Y2=0
cc_557 N_D_M1031_g N_VPWR_c_807_n 0.00982266f $X=9.125 $Y=2.4 $X2=0 $Y2=0
cc_558 N_D_M1036_g N_VPWR_c_807_n 0.00986008f $X=9.575 $Y=2.4 $X2=0 $Y2=0
cc_559 N_D_M1028_g N_Y_c_989_n 6.3785e-19 $X=8.225 $Y=2.4 $X2=0 $Y2=0
cc_560 N_D_M1028_g N_Y_c_1079_n 0.0171084f $X=8.225 $Y=2.4 $X2=0 $Y2=0
cc_561 D N_Y_c_1079_n 0.00143862f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_562 N_D_M1028_g N_Y_c_990_n 0.0116961f $X=8.225 $Y=2.4 $X2=0 $Y2=0
cc_563 N_D_M1030_g N_Y_c_990_n 0.0119382f $X=8.675 $Y=2.4 $X2=0 $Y2=0
cc_564 N_D_M1031_g N_Y_c_990_n 6.50516e-19 $X=9.125 $Y=2.4 $X2=0 $Y2=0
cc_565 N_D_M1030_g N_Y_c_1097_n 0.012931f $X=8.675 $Y=2.4 $X2=0 $Y2=0
cc_566 N_D_M1031_g N_Y_c_1097_n 0.012931f $X=9.125 $Y=2.4 $X2=0 $Y2=0
cc_567 D N_Y_c_1097_n 0.0395816f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_568 N_D_c_727_n N_Y_c_1097_n 4.38169e-19 $X=9.585 $Y=1.465 $X2=0 $Y2=0
cc_569 N_D_M1031_g N_Y_c_1101_n 8.84614e-19 $X=9.125 $Y=2.4 $X2=0 $Y2=0
cc_570 N_D_M1036_g N_Y_c_1101_n 0.0025567f $X=9.575 $Y=2.4 $X2=0 $Y2=0
cc_571 D N_Y_c_1101_n 0.0237862f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_572 N_D_c_727_n N_Y_c_1101_n 4.97911e-19 $X=9.585 $Y=1.465 $X2=0 $Y2=0
cc_573 N_D_M1030_g N_Y_c_991_n 6.50516e-19 $X=8.675 $Y=2.4 $X2=0 $Y2=0
cc_574 N_D_M1031_g N_Y_c_991_n 0.0119382f $X=9.125 $Y=2.4 $X2=0 $Y2=0
cc_575 N_D_M1036_g N_Y_c_991_n 0.0112644f $X=9.575 $Y=2.4 $X2=0 $Y2=0
cc_576 N_D_M1028_g N_Y_c_994_n 6.08944e-19 $X=8.225 $Y=2.4 $X2=0 $Y2=0
cc_577 N_D_M1028_g N_Y_c_1109_n 8.84614e-19 $X=8.225 $Y=2.4 $X2=0 $Y2=0
cc_578 N_D_M1030_g N_Y_c_1109_n 8.84614e-19 $X=8.675 $Y=2.4 $X2=0 $Y2=0
cc_579 D N_Y_c_1109_n 0.0237862f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_580 N_D_c_727_n N_Y_c_1109_n 4.97596e-19 $X=9.585 $Y=1.465 $X2=0 $Y2=0
cc_581 N_D_M1005_g N_VGND_c_1180_n 0.0092592f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_582 N_D_M1009_g N_VGND_c_1180_n 0.00921026f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_583 N_D_M1012_g N_VGND_c_1180_n 4.56715e-19 $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_584 N_D_M1009_g N_VGND_c_1181_n 4.56715e-19 $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_585 N_D_M1012_g N_VGND_c_1181_n 0.00921984f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_586 N_D_M1034_g N_VGND_c_1181_n 0.0054497f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_587 N_D_M1005_g N_VGND_c_1183_n 0.00383152f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_588 N_D_M1009_g N_VGND_c_1184_n 0.00383152f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_589 N_D_M1012_g N_VGND_c_1184_n 0.00383152f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_590 N_D_M1034_g N_VGND_c_1185_n 0.00434272f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_591 N_D_M1005_g N_VGND_c_1186_n 0.00757637f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_592 N_D_M1009_g N_VGND_c_1186_n 0.0075754f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_593 N_D_M1012_g N_VGND_c_1186_n 0.0075754f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_594 N_D_M1034_g N_VGND_c_1186_n 0.00824376f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_595 N_D_M1005_g N_A_828_74#_c_1338_n 3.00542e-19 $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_596 N_D_M1005_g N_A_1229_74#_c_1391_n 3.92313e-19 $X=8.225 $Y=0.74 $X2=0
+ $Y2=0
cc_597 N_D_M1005_g N_A_1229_74#_c_1392_n 0.0159972f $X=8.225 $Y=0.74 $X2=0 $Y2=0
cc_598 N_D_M1009_g N_A_1229_74#_c_1392_n 0.0124847f $X=8.655 $Y=0.74 $X2=0 $Y2=0
cc_599 D N_A_1229_74#_c_1392_n 0.0395058f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_600 N_D_c_727_n N_A_1229_74#_c_1392_n 0.00281527f $X=9.585 $Y=1.465 $X2=0
+ $Y2=0
cc_601 N_D_M1009_g N_A_1229_74#_c_1393_n 3.92313e-19 $X=8.655 $Y=0.74 $X2=0
+ $Y2=0
cc_602 N_D_M1012_g N_A_1229_74#_c_1393_n 3.92313e-19 $X=9.085 $Y=0.74 $X2=0
+ $Y2=0
cc_603 N_D_M1012_g N_A_1229_74#_c_1394_n 0.0128832f $X=9.085 $Y=0.74 $X2=0 $Y2=0
cc_604 N_D_M1034_g N_A_1229_74#_c_1394_n 0.0126756f $X=9.585 $Y=0.74 $X2=0 $Y2=0
cc_605 D N_A_1229_74#_c_1394_n 0.0792081f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_606 N_D_c_727_n N_A_1229_74#_c_1394_n 0.0104362f $X=9.585 $Y=1.465 $X2=0
+ $Y2=0
cc_607 N_D_M1012_g N_A_1229_74#_c_1395_n 9.27941e-19 $X=9.085 $Y=0.74 $X2=0
+ $Y2=0
cc_608 N_D_M1034_g N_A_1229_74#_c_1395_n 0.00959678f $X=9.585 $Y=0.74 $X2=0
+ $Y2=0
cc_609 N_D_M1005_g N_A_1229_74#_c_1397_n 6.32871e-19 $X=8.225 $Y=0.74 $X2=0
+ $Y2=0
cc_610 D N_A_1229_74#_c_1398_n 0.0147161f $X=9.755 $Y=1.58 $X2=0 $Y2=0
cc_611 N_D_c_727_n N_A_1229_74#_c_1398_n 0.00246761f $X=9.585 $Y=1.465 $X2=0
+ $Y2=0
cc_612 N_VPWR_M1002_d N_Y_c_1002_n 0.00316447f $X=3.165 $Y=1.84 $X2=0 $Y2=0
cc_613 N_VPWR_c_812_n N_Y_c_1002_n 0.0170259f $X=3.3 $Y=2.495 $X2=0 $Y2=0
cc_614 N_VPWR_c_812_n N_Y_c_983_n 0.0232805f $X=3.3 $Y=2.495 $X2=0 $Y2=0
cc_615 N_VPWR_c_813_n N_Y_c_983_n 0.0105983f $X=4.035 $Y=3.33 $X2=0 $Y2=0
cc_616 N_VPWR_c_814_n N_Y_c_983_n 0.0232805f $X=4.2 $Y=2.495 $X2=0 $Y2=0
cc_617 N_VPWR_c_807_n N_Y_c_983_n 0.00847107f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_618 N_VPWR_M1006_d N_Y_c_1009_n 0.00329596f $X=4.065 $Y=1.84 $X2=0 $Y2=0
cc_619 N_VPWR_c_814_n N_Y_c_1009_n 0.0169445f $X=4.2 $Y=2.495 $X2=0 $Y2=0
cc_620 N_VPWR_c_814_n N_Y_c_984_n 0.022534f $X=4.2 $Y=2.495 $X2=0 $Y2=0
cc_621 N_VPWR_c_815_n N_Y_c_984_n 0.0123179f $X=4.985 $Y=3.33 $X2=0 $Y2=0
cc_622 N_VPWR_c_807_n N_Y_c_984_n 0.0101276f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_623 N_VPWR_M1013_s N_Y_c_1041_n 0.0040648f $X=4.965 $Y=1.84 $X2=0 $Y2=0
cc_624 N_VPWR_c_816_n N_Y_c_1041_n 0.0189268f $X=5.15 $Y=2.355 $X2=0 $Y2=0
cc_625 N_VPWR_c_816_n N_Y_c_986_n 0.0266644f $X=5.15 $Y=2.355 $X2=0 $Y2=0
cc_626 N_VPWR_c_817_n N_Y_c_986_n 0.0265275f $X=6.05 $Y=2.325 $X2=0 $Y2=0
cc_627 N_VPWR_c_829_n N_Y_c_986_n 0.00749631f $X=5.885 $Y=3.33 $X2=0 $Y2=0
cc_628 N_VPWR_c_807_n N_Y_c_986_n 0.0062048f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_629 N_VPWR_M1020_s N_Y_c_987_n 0.00165831f $X=5.915 $Y=1.84 $X2=0 $Y2=0
cc_630 N_VPWR_c_817_n N_Y_c_987_n 0.0148589f $X=6.05 $Y=2.325 $X2=0 $Y2=0
cc_631 N_VPWR_c_817_n N_Y_c_988_n 0.0276912f $X=6.05 $Y=2.325 $X2=0 $Y2=0
cc_632 N_VPWR_c_818_n N_Y_c_988_n 0.0266809f $X=7 $Y=2.455 $X2=0 $Y2=0
cc_633 N_VPWR_c_830_n N_Y_c_988_n 0.0144623f $X=6.835 $Y=3.33 $X2=0 $Y2=0
cc_634 N_VPWR_c_807_n N_Y_c_988_n 0.0118344f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_635 N_VPWR_M1026_s N_Y_c_1070_n 0.00534029f $X=6.815 $Y=1.84 $X2=0 $Y2=0
cc_636 N_VPWR_c_818_n N_Y_c_1070_n 0.0208278f $X=7 $Y=2.455 $X2=0 $Y2=0
cc_637 N_VPWR_c_818_n N_Y_c_989_n 0.0266809f $X=7 $Y=2.455 $X2=0 $Y2=0
cc_638 N_VPWR_c_819_n N_Y_c_989_n 0.0144623f $X=7.865 $Y=3.33 $X2=0 $Y2=0
cc_639 N_VPWR_c_820_n N_Y_c_989_n 0.0234083f $X=7.95 $Y=2.455 $X2=0 $Y2=0
cc_640 N_VPWR_c_807_n N_Y_c_989_n 0.0118344f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_641 N_VPWR_M1029_s N_Y_c_1079_n 0.0100499f $X=7.815 $Y=1.84 $X2=0 $Y2=0
cc_642 N_VPWR_c_820_n N_Y_c_1079_n 0.0167599f $X=7.95 $Y=2.455 $X2=0 $Y2=0
cc_643 N_VPWR_c_820_n N_Y_c_990_n 0.0266484f $X=7.95 $Y=2.455 $X2=0 $Y2=0
cc_644 N_VPWR_c_821_n N_Y_c_990_n 0.0144623f $X=8.815 $Y=3.33 $X2=0 $Y2=0
cc_645 N_VPWR_c_822_n N_Y_c_990_n 0.0233699f $X=8.9 $Y=2.455 $X2=0 $Y2=0
cc_646 N_VPWR_c_807_n N_Y_c_990_n 0.0118344f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_647 N_VPWR_M1030_s N_Y_c_1097_n 0.00315967f $X=8.765 $Y=1.84 $X2=0 $Y2=0
cc_648 N_VPWR_c_822_n N_Y_c_1097_n 0.0126919f $X=8.9 $Y=2.455 $X2=0 $Y2=0
cc_649 N_VPWR_c_822_n N_Y_c_991_n 0.0233699f $X=8.9 $Y=2.455 $X2=0 $Y2=0
cc_650 N_VPWR_c_824_n N_Y_c_991_n 0.0289761f $X=9.8 $Y=2.115 $X2=0 $Y2=0
cc_651 N_VPWR_c_831_n N_Y_c_991_n 0.0144623f $X=9.715 $Y=3.33 $X2=0 $Y2=0
cc_652 N_VPWR_c_807_n N_Y_c_991_n 0.0118344f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_653 N_VPWR_c_816_n N_Y_c_1019_n 0.0296971f $X=5.15 $Y=2.355 $X2=0 $Y2=0
cc_654 N_VPWR_c_811_n Y 0.0437222f $X=2.17 $Y=2.495 $X2=0 $Y2=0
cc_655 N_VPWR_c_812_n Y 0.0233983f $X=3.3 $Y=2.495 $X2=0 $Y2=0
cc_656 N_VPWR_c_825_n Y 0.0199376f $X=3.135 $Y=3.33 $X2=0 $Y2=0
cc_657 N_VPWR_c_807_n Y 0.015606f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_658 N_Y_c_998_n N_A_374_74#_M1007_d 0.00349797f $X=3.335 $Y=0.955 $X2=0 $Y2=0
cc_659 N_Y_c_980_n N_A_374_74#_M1033_d 0.00176461f $X=5.515 $Y=1.175 $X2=0 $Y2=0
cc_660 N_Y_c_980_n N_A_374_74#_M1008_s 0.00176891f $X=5.515 $Y=1.175 $X2=0 $Y2=0
cc_661 N_Y_c_980_n N_A_374_74#_M1032_s 7.73211e-19 $X=5.515 $Y=1.175 $X2=0 $Y2=0
cc_662 N_Y_M1001_s N_A_374_74#_c_1273_n 0.00295551f $X=2.305 $Y=0.37 $X2=0 $Y2=0
cc_663 N_Y_c_998_n N_A_374_74#_c_1273_n 0.00404257f $X=3.335 $Y=0.955 $X2=0
+ $Y2=0
cc_664 N_Y_c_1010_n N_A_374_74#_c_1273_n 0.0199719f $X=2.485 $Y=0.815 $X2=0
+ $Y2=0
cc_665 N_Y_M1011_s N_A_374_74#_c_1275_n 0.00176461f $X=3.28 $Y=0.37 $X2=0 $Y2=0
cc_666 N_Y_c_998_n N_A_374_74#_c_1275_n 0.00402702f $X=3.335 $Y=0.955 $X2=0
+ $Y2=0
cc_667 N_Y_c_1168_p N_A_374_74#_c_1275_n 0.012613f $X=3.42 $Y=0.87 $X2=0 $Y2=0
cc_668 N_Y_c_980_n N_A_374_74#_c_1275_n 0.00270072f $X=5.515 $Y=1.175 $X2=0
+ $Y2=0
cc_669 N_Y_c_980_n N_A_374_74#_c_1293_n 0.0870842f $X=5.515 $Y=1.175 $X2=0 $Y2=0
cc_670 N_Y_c_980_n N_A_374_74#_c_1287_n 0.0153817f $X=5.515 $Y=1.175 $X2=0 $Y2=0
cc_671 N_Y_c_998_n N_A_374_74#_c_1276_n 0.0165533f $X=3.335 $Y=0.955 $X2=0 $Y2=0
cc_672 N_Y_c_980_n N_A_374_74#_c_1277_n 0.00517215f $X=5.515 $Y=1.175 $X2=0
+ $Y2=0
cc_673 N_Y_c_980_n N_A_828_74#_M1004_d 0.00176891f $X=5.515 $Y=1.175 $X2=-0.19
+ $Y2=-0.245
cc_674 N_Y_c_980_n N_A_828_74#_M1014_d 0.00347389f $X=5.515 $Y=1.175 $X2=0 $Y2=0
cc_675 N_Y_c_980_n N_A_1229_74#_c_1389_n 0.0028602f $X=5.515 $Y=1.175 $X2=0
+ $Y2=0
cc_676 N_Y_c_987_n N_A_1229_74#_c_1389_n 0.0019066f $X=6.335 $Y=1.905 $X2=0
+ $Y2=0
cc_677 N_Y_c_994_n N_A_1229_74#_c_1390_n 0.00163688f $X=7.5 $Y=1.985 $X2=0 $Y2=0
cc_678 N_VGND_c_1183_n N_A_374_74#_c_1273_n 0.045537f $X=8.275 $Y=0 $X2=0 $Y2=0
cc_679 N_VGND_c_1186_n N_A_374_74#_c_1273_n 0.0257922f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_680 N_VGND_c_1183_n N_A_374_74#_c_1274_n 0.0121867f $X=8.275 $Y=0 $X2=0 $Y2=0
cc_681 N_VGND_c_1186_n N_A_374_74#_c_1274_n 0.00660921f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_682 N_VGND_c_1183_n N_A_374_74#_c_1275_n 0.051499f $X=8.275 $Y=0 $X2=0 $Y2=0
cc_683 N_VGND_c_1186_n N_A_374_74#_c_1275_n 0.0285503f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_684 N_VGND_c_1183_n N_A_374_74#_c_1293_n 0.00197884f $X=8.275 $Y=0 $X2=0
+ $Y2=0
cc_685 N_VGND_c_1186_n N_A_374_74#_c_1293_n 0.00647053f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_686 N_VGND_c_1183_n N_A_374_74#_c_1276_n 0.0226536f $X=8.275 $Y=0 $X2=0 $Y2=0
cc_687 N_VGND_c_1186_n N_A_374_74#_c_1276_n 0.0124411f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_688 N_VGND_c_1183_n N_A_828_74#_c_1336_n 0.159083f $X=8.275 $Y=0 $X2=0 $Y2=0
cc_689 N_VGND_c_1186_n N_A_828_74#_c_1336_n 0.0896859f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_690 N_VGND_c_1180_n N_A_828_74#_c_1338_n 0.0029789f $X=8.44 $Y=0.57 $X2=0
+ $Y2=0
cc_691 N_VGND_c_1183_n N_A_828_74#_c_1338_n 0.0564897f $X=8.275 $Y=0 $X2=0 $Y2=0
cc_692 N_VGND_c_1186_n N_A_828_74#_c_1338_n 0.0313161f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_693 N_VGND_c_1183_n N_A_828_74#_c_1340_n 0.0231282f $X=8.275 $Y=0 $X2=0 $Y2=0
cc_694 N_VGND_c_1186_n N_A_828_74#_c_1340_n 0.0125338f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_695 N_VGND_c_1180_n N_A_1229_74#_c_1391_n 0.0164567f $X=8.44 $Y=0.57 $X2=0
+ $Y2=0
cc_696 N_VGND_c_1183_n N_A_1229_74#_c_1391_n 0.00749631f $X=8.275 $Y=0 $X2=0
+ $Y2=0
cc_697 N_VGND_c_1186_n N_A_1229_74#_c_1391_n 0.0062048f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_698 N_VGND_M1005_s N_A_1229_74#_c_1392_n 0.00176461f $X=8.3 $Y=0.37 $X2=0
+ $Y2=0
cc_699 N_VGND_c_1180_n N_A_1229_74#_c_1392_n 0.0171619f $X=8.44 $Y=0.57 $X2=0
+ $Y2=0
cc_700 N_VGND_c_1180_n N_A_1229_74#_c_1393_n 0.0164567f $X=8.44 $Y=0.57 $X2=0
+ $Y2=0
cc_701 N_VGND_c_1181_n N_A_1229_74#_c_1393_n 0.0164567f $X=9.3 $Y=0.57 $X2=0
+ $Y2=0
cc_702 N_VGND_c_1184_n N_A_1229_74#_c_1393_n 0.00749631f $X=9.135 $Y=0 $X2=0
+ $Y2=0
cc_703 N_VGND_c_1186_n N_A_1229_74#_c_1393_n 0.0062048f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_704 N_VGND_M1012_s N_A_1229_74#_c_1394_n 0.00250873f $X=9.16 $Y=0.37 $X2=0
+ $Y2=0
cc_705 N_VGND_c_1181_n N_A_1229_74#_c_1394_n 0.0210288f $X=9.3 $Y=0.57 $X2=0
+ $Y2=0
cc_706 N_VGND_c_1181_n N_A_1229_74#_c_1395_n 0.0173003f $X=9.3 $Y=0.57 $X2=0
+ $Y2=0
cc_707 N_VGND_c_1185_n N_A_1229_74#_c_1395_n 0.0145639f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_708 N_VGND_c_1186_n N_A_1229_74#_c_1395_n 0.0119984f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_709 N_A_374_74#_c_1293_n N_A_828_74#_M1004_d 0.003292f $X=5.565 $Y=0.835
+ $X2=-0.19 $Y2=-0.245
cc_710 N_A_374_74#_c_1293_n N_A_828_74#_M1014_d 0.0070998f $X=5.565 $Y=0.835
+ $X2=0 $Y2=0
cc_711 N_A_374_74#_M1008_s N_A_828_74#_c_1336_n 0.00171274f $X=4.57 $Y=0.37
+ $X2=0 $Y2=0
cc_712 N_A_374_74#_c_1275_n N_A_828_74#_c_1336_n 0.0119071f $X=3.685 $Y=0.34
+ $X2=0 $Y2=0
cc_713 N_A_374_74#_c_1293_n N_A_828_74#_c_1336_n 0.0708016f $X=5.565 $Y=0.835
+ $X2=0 $Y2=0
cc_714 N_A_374_74#_M1032_s N_A_828_74#_c_1337_n 0.00273752f $X=5.59 $Y=0.37
+ $X2=0 $Y2=0
cc_715 N_A_374_74#_c_1293_n N_A_828_74#_c_1337_n 0.00442249f $X=5.565 $Y=0.835
+ $X2=0 $Y2=0
cc_716 N_A_374_74#_c_1277_n N_A_828_74#_c_1337_n 0.0194173f $X=5.73 $Y=0.715
+ $X2=0 $Y2=0
cc_717 N_A_374_74#_c_1277_n N_A_1229_74#_c_1387_n 0.02146f $X=5.73 $Y=0.715
+ $X2=0 $Y2=0
cc_718 N_A_828_74#_c_1337_n N_A_1229_74#_M1023_s 0.00273752f $X=6.555 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_719 N_A_828_74#_c_1338_n N_A_1229_74#_M1025_s 0.00176461f $X=7.415 $Y=0.34
+ $X2=0 $Y2=0
cc_720 N_A_828_74#_c_1337_n N_A_1229_74#_c_1387_n 0.0185632f $X=6.555 $Y=0.34
+ $X2=0 $Y2=0
cc_721 N_A_828_74#_M1023_d N_A_1229_74#_c_1388_n 0.00176461f $X=6.58 $Y=0.37
+ $X2=0 $Y2=0
cc_722 N_A_828_74#_c_1337_n N_A_1229_74#_c_1388_n 0.0031794f $X=6.555 $Y=0.34
+ $X2=0 $Y2=0
cc_723 N_A_828_74#_c_1346_n N_A_1229_74#_c_1388_n 0.0168793f $X=6.72 $Y=0.58
+ $X2=0 $Y2=0
cc_724 N_A_828_74#_c_1338_n N_A_1229_74#_c_1388_n 0.0031794f $X=7.415 $Y=0.34
+ $X2=0 $Y2=0
cc_725 N_A_828_74#_c_1338_n N_A_1229_74#_c_1455_n 0.0124395f $X=7.415 $Y=0.34
+ $X2=0 $Y2=0
cc_726 N_A_828_74#_M1035_d N_A_1229_74#_c_1390_n 0.00176461f $X=7.44 $Y=0.37
+ $X2=0 $Y2=0
cc_727 N_A_828_74#_c_1338_n N_A_1229_74#_c_1390_n 0.0031794f $X=7.415 $Y=0.34
+ $X2=0 $Y2=0
cc_728 N_A_828_74#_c_1352_n N_A_1229_74#_c_1390_n 0.0168793f $X=7.58 $Y=0.58
+ $X2=0 $Y2=0
cc_729 N_A_828_74#_c_1338_n N_A_1229_74#_c_1391_n 0.00370621f $X=7.415 $Y=0.34
+ $X2=0 $Y2=0

* File: sky130_fd_sc_ms__a2111o_4.pxi.spice
* Created: Fri Aug 28 16:55:40 2020
* 
x_PM_SKY130_FD_SC_MS__A2111O_4%A_137_260# N_A_137_260#_M1011_d
+ N_A_137_260#_M1004_s N_A_137_260#_M1009_s N_A_137_260#_M1001_d
+ N_A_137_260#_M1002_d N_A_137_260#_M1014_g N_A_137_260#_M1016_g
+ N_A_137_260#_M1003_g N_A_137_260#_M1018_g N_A_137_260#_M1010_g
+ N_A_137_260#_M1023_g N_A_137_260#_M1020_g N_A_137_260#_M1024_g
+ N_A_137_260#_c_165_n N_A_137_260#_c_166_n N_A_137_260#_c_167_n
+ N_A_137_260#_c_183_n N_A_137_260#_c_168_n N_A_137_260#_c_169_n
+ N_A_137_260#_c_170_n N_A_137_260#_c_171_n N_A_137_260#_c_172_n
+ N_A_137_260#_c_173_n N_A_137_260#_c_174_n N_A_137_260#_c_175_n
+ N_A_137_260#_c_184_n N_A_137_260#_c_176_n N_A_137_260#_c_177_n
+ N_A_137_260#_c_178_n PM_SKY130_FD_SC_MS__A2111O_4%A_137_260#
x_PM_SKY130_FD_SC_MS__A2111O_4%D1 N_D1_M1011_g N_D1_M1002_g N_D1_M1021_g
+ N_D1_M1005_g D1 N_D1_c_340_n N_D1_c_341_n PM_SKY130_FD_SC_MS__A2111O_4%D1
x_PM_SKY130_FD_SC_MS__A2111O_4%C1 N_C1_M1004_g N_C1_M1006_g N_C1_M1022_g
+ N_C1_c_398_n N_C1_M1008_g N_C1_c_399_n N_C1_c_400_n C1 C1 C1 N_C1_c_402_n
+ PM_SKY130_FD_SC_MS__A2111O_4%C1
x_PM_SKY130_FD_SC_MS__A2111O_4%B1 N_B1_c_460_n N_B1_M1009_g N_B1_c_461_n
+ N_B1_c_462_n N_B1_c_463_n N_B1_M1026_g N_B1_M1013_g N_B1_c_467_n N_B1_M1015_g
+ B1 B1 N_B1_c_465_n PM_SKY130_FD_SC_MS__A2111O_4%B1
x_PM_SKY130_FD_SC_MS__A2111O_4%A1 N_A1_M1017_g N_A1_M1001_g N_A1_M1019_g
+ N_A1_M1012_g A1 A1 N_A1_c_518_n PM_SKY130_FD_SC_MS__A2111O_4%A1
x_PM_SKY130_FD_SC_MS__A2111O_4%A2 N_A2_M1000_g N_A2_M1007_g N_A2_M1025_g
+ N_A2_M1027_g A2 A2 N_A2_c_572_n PM_SKY130_FD_SC_MS__A2111O_4%A2
x_PM_SKY130_FD_SC_MS__A2111O_4%VPWR N_VPWR_M1014_s N_VPWR_M1016_s N_VPWR_M1023_s
+ N_VPWR_M1017_d N_VPWR_M1000_s N_VPWR_c_613_n N_VPWR_c_614_n N_VPWR_c_615_n
+ N_VPWR_c_616_n N_VPWR_c_617_n N_VPWR_c_618_n N_VPWR_c_619_n N_VPWR_c_620_n
+ N_VPWR_c_621_n N_VPWR_c_622_n N_VPWR_c_623_n VPWR N_VPWR_c_624_n
+ N_VPWR_c_625_n N_VPWR_c_626_n N_VPWR_c_612_n N_VPWR_c_628_n N_VPWR_c_629_n
+ PM_SKY130_FD_SC_MS__A2111O_4%VPWR
x_PM_SKY130_FD_SC_MS__A2111O_4%X N_X_M1003_s N_X_M1020_s N_X_M1014_d N_X_M1018_d
+ N_X_c_712_n N_X_c_713_n N_X_c_719_n N_X_c_720_n N_X_c_721_n N_X_c_722_n
+ N_X_c_714_n N_X_c_715_n N_X_c_723_n N_X_c_716_n N_X_c_724_n N_X_c_717_n X X
+ PM_SKY130_FD_SC_MS__A2111O_4%X
x_PM_SKY130_FD_SC_MS__A2111O_4%A_549_392# N_A_549_392#_M1002_s
+ N_A_549_392#_M1005_s N_A_549_392#_M1008_s N_A_549_392#_c_788_n
+ N_A_549_392#_c_789_n N_A_549_392#_c_790_n N_A_549_392#_c_791_n
+ N_A_549_392#_c_792_n N_A_549_392#_c_793_n N_A_549_392#_c_794_n
+ PM_SKY130_FD_SC_MS__A2111O_4%A_549_392#
x_PM_SKY130_FD_SC_MS__A2111O_4%A_817_392# N_A_817_392#_M1006_d
+ N_A_817_392#_M1013_d N_A_817_392#_c_834_n N_A_817_392#_c_835_n
+ N_A_817_392#_c_836_n PM_SKY130_FD_SC_MS__A2111O_4%A_817_392#
x_PM_SKY130_FD_SC_MS__A2111O_4%A_1013_392# N_A_1013_392#_M1013_s
+ N_A_1013_392#_M1015_s N_A_1013_392#_M1019_s N_A_1013_392#_M1025_d
+ N_A_1013_392#_c_859_n N_A_1013_392#_c_860_n N_A_1013_392#_c_861_n
+ N_A_1013_392#_c_862_n N_A_1013_392#_c_863_n N_A_1013_392#_c_864_n
+ N_A_1013_392#_c_865_n N_A_1013_392#_c_866_n N_A_1013_392#_c_867_n
+ N_A_1013_392#_c_868_n PM_SKY130_FD_SC_MS__A2111O_4%A_1013_392#
x_PM_SKY130_FD_SC_MS__A2111O_4%VGND N_VGND_M1003_d N_VGND_M1010_d N_VGND_M1024_d
+ N_VGND_M1021_s N_VGND_M1022_d N_VGND_M1026_d N_VGND_M1007_s N_VGND_c_912_n
+ N_VGND_c_913_n N_VGND_c_914_n N_VGND_c_915_n N_VGND_c_916_n N_VGND_c_917_n
+ N_VGND_c_918_n N_VGND_c_919_n N_VGND_c_920_n N_VGND_c_921_n N_VGND_c_922_n
+ N_VGND_c_923_n N_VGND_c_924_n VGND N_VGND_c_925_n N_VGND_c_926_n
+ N_VGND_c_927_n N_VGND_c_928_n N_VGND_c_929_n N_VGND_c_930_n N_VGND_c_931_n
+ N_VGND_c_932_n N_VGND_c_933_n N_VGND_c_934_n PM_SKY130_FD_SC_MS__A2111O_4%VGND
x_PM_SKY130_FD_SC_MS__A2111O_4%A_1210_74# N_A_1210_74#_M1001_s
+ N_A_1210_74#_M1012_s N_A_1210_74#_M1027_d N_A_1210_74#_c_1026_n
+ N_A_1210_74#_c_1027_n N_A_1210_74#_c_1028_n N_A_1210_74#_c_1029_n
+ N_A_1210_74#_c_1030_n N_A_1210_74#_c_1031_n
+ PM_SKY130_FD_SC_MS__A2111O_4%A_1210_74#
cc_1 VNB N_A_137_260#_M1014_g 0.00167481f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=2.4
cc_2 VNB N_A_137_260#_M1016_g 0.00154188f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.4
cc_3 VNB N_A_137_260#_M1003_g 0.0246266f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=0.74
cc_4 VNB N_A_137_260#_M1018_g 0.00154301f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=2.4
cc_5 VNB N_A_137_260#_M1010_g 0.0209331f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=0.74
cc_6 VNB N_A_137_260#_M1023_g 0.00243969f $X=-0.19 $Y=-0.245 $X2=2.125 $Y2=2.4
cc_7 VNB N_A_137_260#_M1020_g 0.0209331f $X=-0.19 $Y=-0.245 $X2=2.145 $Y2=0.74
cc_8 VNB N_A_137_260#_M1024_g 0.021412f $X=-0.19 $Y=-0.245 $X2=2.575 $Y2=0.74
cc_9 VNB N_A_137_260#_c_165_n 0.0133831f $X=-0.19 $Y=-0.245 $X2=3.045 $Y2=1.465
cc_10 VNB N_A_137_260#_c_166_n 0.00206705f $X=-0.19 $Y=-0.245 $X2=3.265
+ $Y2=0.515
cc_11 VNB N_A_137_260#_c_167_n 0.00164495f $X=-0.19 $Y=-0.245 $X2=3.13 $Y2=1.3
cc_12 VNB N_A_137_260#_c_168_n 0.00791729f $X=-0.19 $Y=-0.245 $X2=4.05 $Y2=1.005
cc_13 VNB N_A_137_260#_c_169_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=4.135
+ $Y2=0.515
cc_14 VNB N_A_137_260#_c_170_n 0.00917015f $X=-0.19 $Y=-0.245 $X2=4.92 $Y2=1.195
cc_15 VNB N_A_137_260#_c_171_n 0.003224f $X=-0.19 $Y=-0.245 $X2=5.005 $Y2=0.515
cc_16 VNB N_A_137_260#_c_172_n 0.0166742f $X=-0.19 $Y=-0.245 $X2=6.51 $Y2=1.195
cc_17 VNB N_A_137_260#_c_173_n 9.35553e-19 $X=-0.19 $Y=-0.245 $X2=6.605 $Y2=0.79
cc_18 VNB N_A_137_260#_c_174_n 0.00256255f $X=-0.19 $Y=-0.245 $X2=3.197
+ $Y2=1.005
cc_19 VNB N_A_137_260#_c_175_n 2.54259e-19 $X=-0.19 $Y=-0.245 $X2=3.13 $Y2=1.465
cc_20 VNB N_A_137_260#_c_176_n 0.00425475f $X=-0.19 $Y=-0.245 $X2=4.135
+ $Y2=1.005
cc_21 VNB N_A_137_260#_c_177_n 0.00159638f $X=-0.19 $Y=-0.245 $X2=5.005
+ $Y2=1.195
cc_22 VNB N_A_137_260#_c_178_n 0.126542f $X=-0.19 $Y=-0.245 $X2=2.575 $Y2=1.465
cc_23 VNB N_D1_M1011_g 0.0243515f $X=-0.19 $Y=-0.245 $X2=4.865 $Y2=0.37
cc_24 VNB N_D1_M1002_g 0.00424565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_D1_M1021_g 0.0233084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_D1_M1005_g 0.00307356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_D1_c_340_n 0.00521187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_D1_c_341_n 0.039576f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=1.3
cc_29 VNB N_C1_M1004_g 0.0328076f $X=-0.19 $Y=-0.245 $X2=4.865 $Y2=0.37
cc_30 VNB N_C1_c_398_n 0.0162228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_C1_c_399_n 0.0149068f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=2.4
cc_32 VNB N_C1_c_400_n 0.00789277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB C1 0.00771653f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.4
cc_34 VNB N_C1_c_402_n 0.0350532f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=2.4
cc_35 VNB N_B1_c_460_n 0.0150917f $X=-0.19 $Y=-0.245 $X2=3.125 $Y2=0.37
cc_36 VNB N_B1_c_461_n 0.0151763f $X=-0.19 $Y=-0.245 $X2=6.465 $Y2=0.37
cc_37 VNB N_B1_c_462_n 0.00874277f $X=-0.19 $Y=-0.245 $X2=3.185 $Y2=1.96
cc_38 VNB N_B1_c_463_n 0.019199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB B1 0.00301796f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=2.4
cc_40 VNB N_B1_c_465_n 0.0972644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A1_M1001_g 0.0384872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A1_M1012_g 0.0324852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB A1 0.00484998f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=2.4
cc_44 VNB N_A1_c_518_n 0.0274267f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=0.74
cc_45 VNB N_A2_M1000_g 0.00347224f $X=-0.19 $Y=-0.245 $X2=4.865 $Y2=0.37
cc_46 VNB N_A2_M1007_g 0.0233949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A2_M1025_g 0.00418093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A2_M1027_g 0.0324492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB A2 0.0203442f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=2.4
cc_50 VNB N_A2_c_572_n 0.0436682f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=1.63
cc_51 VNB N_VPWR_c_612_n 0.342803f $X=-0.19 $Y=-0.245 $X2=5.005 $Y2=1.11
cc_52 VNB N_X_c_712_n 0.0153235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_X_c_713_n 0.0316066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_X_c_714_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_X_c_715_n 0.00423905f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=2.4
cc_56 VNB N_X_c_716_n 0.00206666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_X_c_717_n 0.00178779f $X=-0.19 $Y=-0.245 $X2=2.575 $Y2=1.3
cc_58 VNB X 0.0359196f $X=-0.19 $Y=-0.245 $X2=2.575 $Y2=0.74
cc_59 VNB N_VGND_c_912_n 0.0254564f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=1.3
cc_60 VNB N_VGND_c_913_n 0.0065212f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=1.63
cc_61 VNB N_VGND_c_914_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=1.675 $Y2=2.4
cc_62 VNB N_VGND_c_915_n 0.00424579f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=0.74
cc_63 VNB N_VGND_c_916_n 0.0182548f $X=-0.19 $Y=-0.245 $X2=2.125 $Y2=1.63
cc_64 VNB N_VGND_c_917_n 0.00266729f $X=-0.19 $Y=-0.245 $X2=2.145 $Y2=1.3
cc_65 VNB N_VGND_c_918_n 0.00250542f $X=-0.19 $Y=-0.245 $X2=2.575 $Y2=1.3
cc_66 VNB N_VGND_c_919_n 0.0158756f $X=-0.19 $Y=-0.245 $X2=3.045 $Y2=1.465
cc_67 VNB N_VGND_c_920_n 0.00396467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_921_n 0.0309422f $X=-0.19 $Y=-0.245 $X2=2.485 $Y2=1.465
cc_69 VNB N_VGND_c_922_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=3.197 $Y2=0.92
cc_70 VNB N_VGND_c_923_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=3.197 $Y2=0.515
cc_71 VNB N_VGND_c_924_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=3.265 $Y2=0.515
cc_72 VNB N_VGND_c_925_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=4.135 $Y2=0.92
cc_73 VNB N_VGND_c_926_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=4.22 $Y2=1.195
cc_74 VNB N_VGND_c_927_n 0.0440384f $X=-0.19 $Y=-0.245 $X2=6.51 $Y2=1.195
cc_75 VNB N_VGND_c_928_n 0.0169136f $X=-0.19 $Y=-0.245 $X2=3.13 $Y2=1.465
cc_76 VNB N_VGND_c_929_n 0.481891f $X=-0.19 $Y=-0.245 $X2=3.13 $Y2=2.035
cc_77 VNB N_VGND_c_930_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=3.32 $Y2=2.115
cc_78 VNB N_VGND_c_931_n 0.00622543f $X=-0.19 $Y=-0.245 $X2=4.135 $Y2=1.195
cc_79 VNB N_VGND_c_932_n 0.00622543f $X=-0.19 $Y=-0.245 $X2=0.775 $Y2=1.465
cc_80 VNB N_VGND_c_933_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=1.465
cc_81 VNB N_VGND_c_934_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=1.465
cc_82 VNB N_A_1210_74#_c_1026_n 0.00750863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1210_74#_c_1027_n 0.00445625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1210_74#_c_1028_n 0.00514874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1210_74#_c_1029_n 0.0137881f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=1.63
cc_86 VNB N_A_1210_74#_c_1030_n 0.00403069f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.4
cc_87 VNB N_A_1210_74#_c_1031_n 0.0237116f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=1.3
cc_88 VPB N_A_137_260#_M1014_g 0.023995f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=2.4
cc_89 VPB N_A_137_260#_M1016_g 0.0220553f $X=-0.19 $Y=1.66 $X2=1.225 $Y2=2.4
cc_90 VPB N_A_137_260#_M1018_g 0.0220607f $X=-0.19 $Y=1.66 $X2=1.675 $Y2=2.4
cc_91 VPB N_A_137_260#_M1023_g 0.0280079f $X=-0.19 $Y=1.66 $X2=2.125 $Y2=2.4
cc_92 VPB N_A_137_260#_c_183_n 0.00254988f $X=-0.19 $Y=1.66 $X2=3.13 $Y2=1.95
cc_93 VPB N_A_137_260#_c_184_n 0.00413741f $X=-0.19 $Y=1.66 $X2=3.32 $Y2=2.115
cc_94 VPB N_D1_M1002_g 0.0352353f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_95 VPB N_D1_M1005_g 0.0271824f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_96 VPB N_D1_c_340_n 0.00444206f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_97 VPB N_C1_M1006_g 0.021783f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_98 VPB N_C1_M1008_g 0.0289924f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=1.63
cc_99 VPB C1 0.00729028f $X=-0.19 $Y=1.66 $X2=1.225 $Y2=2.4
cc_100 VPB N_C1_c_402_n 0.0187919f $X=-0.19 $Y=1.66 $X2=1.675 $Y2=2.4
cc_101 VPB N_B1_M1013_g 0.0290075f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_102 VPB N_B1_c_467_n 0.0168666f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_103 VPB B1 0.00389013f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=2.4
cc_104 VPB N_B1_c_465_n 0.0210569f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_105 VPB N_A1_M1017_g 0.0221751f $X=-0.19 $Y=1.66 $X2=4.865 $Y2=0.37
cc_106 VPB N_A1_M1019_g 0.0221991f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_107 VPB A1 0.00274353f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=2.4
cc_108 VPB N_A1_c_518_n 0.0142792f $X=-0.19 $Y=1.66 $X2=1.285 $Y2=0.74
cc_109 VPB N_A2_M1000_g 0.0283022f $X=-0.19 $Y=1.66 $X2=4.865 $Y2=0.37
cc_110 VPB N_A2_M1025_g 0.0386589f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_111 VPB A2 0.0104325f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=2.4
cc_112 VPB N_VPWR_c_613_n 0.0433927f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=2.4
cc_113 VPB N_VPWR_c_614_n 0.00797179f $X=-0.19 $Y=1.66 $X2=1.225 $Y2=2.4
cc_114 VPB N_VPWR_c_615_n 0.0228338f $X=-0.19 $Y=1.66 $X2=1.285 $Y2=0.74
cc_115 VPB N_VPWR_c_616_n 0.00329129f $X=-0.19 $Y=1.66 $X2=1.715 $Y2=1.3
cc_116 VPB N_VPWR_c_617_n 0.0048755f $X=-0.19 $Y=1.66 $X2=2.125 $Y2=1.63
cc_117 VPB N_VPWR_c_618_n 0.0143948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_619_n 0.0047828f $X=-0.19 $Y=1.66 $X2=2.145 $Y2=1.3
cc_119 VPB N_VPWR_c_620_n 0.0206041f $X=-0.19 $Y=1.66 $X2=2.145 $Y2=0.74
cc_120 VPB N_VPWR_c_621_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_622_n 0.0206041f $X=-0.19 $Y=1.66 $X2=2.575 $Y2=0.74
cc_122 VPB N_VPWR_c_623_n 0.0047828f $X=-0.19 $Y=1.66 $X2=2.575 $Y2=0.74
cc_123 VPB N_VPWR_c_624_n 0.0908814f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_625_n 0.0164337f $X=-0.19 $Y=1.66 $X2=4.05 $Y2=1.005
cc_125 VPB N_VPWR_c_626_n 0.0197879f $X=-0.19 $Y=1.66 $X2=4.22 $Y2=1.195
cc_126 VPB N_VPWR_c_612_n 0.112304f $X=-0.19 $Y=1.66 $X2=5.005 $Y2=1.11
cc_127 VPB N_VPWR_c_628_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_629_n 0.00458862f $X=-0.19 $Y=1.66 $X2=6.64 $Y2=1.11
cc_129 VPB N_X_c_719_n 5.16931e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_X_c_720_n 0.019883f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=1.63
cc_131 VPB N_X_c_721_n 0.00231613f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_X_c_722_n 0.00443716f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_X_c_723_n 0.00231613f $X=-0.19 $Y=1.66 $X2=1.715 $Y2=0.74
cc_134 VPB N_X_c_724_n 0.00227186f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB X 0.008875f $X=-0.19 $Y=1.66 $X2=2.575 $Y2=0.74
cc_136 VPB N_A_549_392#_c_788_n 0.00614299f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_549_392#_c_789_n 0.00192243f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_549_392#_c_790_n 0.00405878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_549_392#_c_791_n 0.00686911f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=2.4
cc_140 VPB N_A_549_392#_c_792_n 0.00596394f $X=-0.19 $Y=1.66 $X2=1.225 $Y2=2.4
cc_141 VPB N_A_549_392#_c_793_n 0.00583793f $X=-0.19 $Y=1.66 $X2=1.285 $Y2=0.74
cc_142 VPB N_A_549_392#_c_794_n 0.00196551f $X=-0.19 $Y=1.66 $X2=1.675 $Y2=1.63
cc_143 VPB N_A_817_392#_c_834_n 0.0177304f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_144 VPB N_A_817_392#_c_835_n 0.00135364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_A_817_392#_c_836_n 0.00224287f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=1.63
cc_146 VPB N_A_1013_392#_c_859_n 0.00582476f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_A_1013_392#_c_860_n 0.00452282f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=2.4
cc_148 VPB N_A_1013_392#_c_861_n 0.00391099f $X=-0.19 $Y=1.66 $X2=0.775 $Y2=2.4
cc_149 VPB N_A_1013_392#_c_862_n 0.00212972f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_1013_392#_c_863_n 0.00336455f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_151 VPB N_A_1013_392#_c_864_n 0.00179594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_152 VPB N_A_1013_392#_c_865_n 0.00393558f $X=-0.19 $Y=1.66 $X2=1.675 $Y2=2.4
cc_153 VPB N_A_1013_392#_c_866_n 0.0106487f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_1013_392#_c_867_n 0.0358769f $X=-0.19 $Y=1.66 $X2=1.715 $Y2=0.74
cc_155 VPB N_A_1013_392#_c_868_n 0.00159638f $X=-0.19 $Y=1.66 $X2=2.125 $Y2=2.4
cc_156 N_A_137_260#_M1024_g N_D1_M1011_g 0.00920717f $X=2.575 $Y=0.74 $X2=0
+ $Y2=0
cc_157 N_A_137_260#_c_166_n N_D1_M1011_g 0.0088411f $X=3.265 $Y=0.515 $X2=0
+ $Y2=0
cc_158 N_A_137_260#_c_167_n N_D1_M1011_g 0.00468003f $X=3.13 $Y=1.3 $X2=0 $Y2=0
cc_159 N_A_137_260#_c_174_n N_D1_M1011_g 0.00383016f $X=3.197 $Y=1.005 $X2=0
+ $Y2=0
cc_160 N_A_137_260#_c_165_n N_D1_M1002_g 0.00201f $X=3.045 $Y=1.465 $X2=0 $Y2=0
cc_161 N_A_137_260#_c_183_n N_D1_M1002_g 0.0147167f $X=3.13 $Y=1.95 $X2=0 $Y2=0
cc_162 N_A_137_260#_c_175_n N_D1_M1002_g 6.56895e-19 $X=3.13 $Y=1.465 $X2=0
+ $Y2=0
cc_163 N_A_137_260#_c_184_n N_D1_M1002_g 0.0113289f $X=3.32 $Y=2.115 $X2=0 $Y2=0
cc_164 N_A_137_260#_c_167_n N_D1_M1021_g 0.00341074f $X=3.13 $Y=1.3 $X2=0 $Y2=0
cc_165 N_A_137_260#_c_168_n N_D1_M1021_g 0.013218f $X=4.05 $Y=1.005 $X2=0 $Y2=0
cc_166 N_A_137_260#_c_183_n N_D1_M1005_g 0.00362807f $X=3.13 $Y=1.95 $X2=0 $Y2=0
cc_167 N_A_137_260#_c_167_n N_D1_c_340_n 0.00282261f $X=3.13 $Y=1.3 $X2=0 $Y2=0
cc_168 N_A_137_260#_c_183_n N_D1_c_340_n 0.0118515f $X=3.13 $Y=1.95 $X2=0 $Y2=0
cc_169 N_A_137_260#_c_168_n N_D1_c_340_n 0.0254454f $X=4.05 $Y=1.005 $X2=0 $Y2=0
cc_170 N_A_137_260#_c_175_n N_D1_c_340_n 0.0266866f $X=3.13 $Y=1.465 $X2=0 $Y2=0
cc_171 N_A_137_260#_c_184_n N_D1_c_340_n 0.00156971f $X=3.32 $Y=2.115 $X2=0
+ $Y2=0
cc_172 N_A_137_260#_c_176_n N_D1_c_340_n 9.88457e-19 $X=4.135 $Y=1.005 $X2=0
+ $Y2=0
cc_173 N_A_137_260#_c_165_n N_D1_c_341_n 0.00928659f $X=3.045 $Y=1.465 $X2=0
+ $Y2=0
cc_174 N_A_137_260#_c_167_n N_D1_c_341_n 0.00170063f $X=3.13 $Y=1.3 $X2=0 $Y2=0
cc_175 N_A_137_260#_c_168_n N_D1_c_341_n 5.56426e-19 $X=4.05 $Y=1.005 $X2=0
+ $Y2=0
cc_176 N_A_137_260#_c_174_n N_D1_c_341_n 0.00468078f $X=3.197 $Y=1.005 $X2=0
+ $Y2=0
cc_177 N_A_137_260#_c_175_n N_D1_c_341_n 0.00872384f $X=3.13 $Y=1.465 $X2=0
+ $Y2=0
cc_178 N_A_137_260#_c_184_n N_D1_c_341_n 0.00292383f $X=3.32 $Y=2.115 $X2=0
+ $Y2=0
cc_179 N_A_137_260#_c_178_n N_D1_c_341_n 0.0165426f $X=2.575 $Y=1.465 $X2=0
+ $Y2=0
cc_180 N_A_137_260#_c_168_n N_C1_M1004_g 0.016344f $X=4.05 $Y=1.005 $X2=0 $Y2=0
cc_181 N_A_137_260#_c_176_n N_C1_M1004_g 0.00443494f $X=4.135 $Y=1.005 $X2=0
+ $Y2=0
cc_182 N_A_137_260#_c_170_n N_C1_c_398_n 0.00385041f $X=4.92 $Y=1.195 $X2=0
+ $Y2=0
cc_183 N_A_137_260#_c_169_n N_C1_c_399_n 0.00126475f $X=4.135 $Y=0.515 $X2=0
+ $Y2=0
cc_184 N_A_137_260#_c_170_n N_C1_c_400_n 0.0102868f $X=4.92 $Y=1.195 $X2=0 $Y2=0
cc_185 N_A_137_260#_c_176_n N_C1_c_400_n 0.00150966f $X=4.135 $Y=1.005 $X2=0
+ $Y2=0
cc_186 N_A_137_260#_c_168_n C1 0.00353585f $X=4.05 $Y=1.005 $X2=0 $Y2=0
cc_187 N_A_137_260#_c_170_n C1 0.0532268f $X=4.92 $Y=1.195 $X2=0 $Y2=0
cc_188 N_A_137_260#_c_172_n C1 0.00511502f $X=6.51 $Y=1.195 $X2=0 $Y2=0
cc_189 N_A_137_260#_c_176_n C1 0.014169f $X=4.135 $Y=1.005 $X2=0 $Y2=0
cc_190 N_A_137_260#_c_177_n C1 0.0150362f $X=5.005 $Y=1.195 $X2=0 $Y2=0
cc_191 N_A_137_260#_c_170_n N_C1_c_402_n 0.00439029f $X=4.92 $Y=1.195 $X2=0
+ $Y2=0
cc_192 N_A_137_260#_c_176_n N_C1_c_402_n 0.00315045f $X=4.135 $Y=1.005 $X2=0
+ $Y2=0
cc_193 N_A_137_260#_c_171_n N_B1_c_460_n 0.00202516f $X=5.005 $Y=0.515 $X2=-0.19
+ $Y2=-0.245
cc_194 N_A_137_260#_c_170_n N_B1_c_461_n 0.00376958f $X=4.92 $Y=1.195 $X2=0
+ $Y2=0
cc_195 N_A_137_260#_c_171_n N_B1_c_461_n 0.00385868f $X=5.005 $Y=0.515 $X2=0
+ $Y2=0
cc_196 N_A_137_260#_c_172_n N_B1_c_461_n 0.00376958f $X=6.51 $Y=1.195 $X2=0
+ $Y2=0
cc_197 N_A_137_260#_c_177_n N_B1_c_461_n 0.00459246f $X=5.005 $Y=1.195 $X2=0
+ $Y2=0
cc_198 N_A_137_260#_c_170_n N_B1_c_462_n 0.0114299f $X=4.92 $Y=1.195 $X2=0 $Y2=0
cc_199 N_A_137_260#_c_171_n N_B1_c_463_n 0.00202516f $X=5.005 $Y=0.515 $X2=0
+ $Y2=0
cc_200 N_A_137_260#_c_172_n B1 0.0521987f $X=6.51 $Y=1.195 $X2=0 $Y2=0
cc_201 N_A_137_260#_c_172_n N_B1_c_465_n 0.0468409f $X=6.51 $Y=1.195 $X2=0 $Y2=0
cc_202 N_A_137_260#_c_172_n N_A1_M1001_g 0.0128558f $X=6.51 $Y=1.195 $X2=0 $Y2=0
cc_203 N_A_137_260#_c_173_n N_A1_M1001_g 0.00268505f $X=6.605 $Y=0.79 $X2=0
+ $Y2=0
cc_204 N_A_137_260#_c_172_n N_A1_M1012_g 0.00567167f $X=6.51 $Y=1.195 $X2=0
+ $Y2=0
cc_205 N_A_137_260#_c_173_n N_A1_M1012_g 0.00661126f $X=6.605 $Y=0.79 $X2=0
+ $Y2=0
cc_206 N_A_137_260#_c_172_n A1 0.0380613f $X=6.51 $Y=1.195 $X2=0 $Y2=0
cc_207 N_A_137_260#_c_172_n N_A1_c_518_n 0.00526706f $X=6.51 $Y=1.195 $X2=0
+ $Y2=0
cc_208 N_A_137_260#_c_172_n N_A2_M1007_g 7.22688e-19 $X=6.51 $Y=1.195 $X2=0
+ $Y2=0
cc_209 N_A_137_260#_c_172_n A2 6.93463e-19 $X=6.51 $Y=1.195 $X2=0 $Y2=0
cc_210 N_A_137_260#_M1014_g N_VPWR_c_613_n 0.00742848f $X=0.775 $Y=2.4 $X2=0
+ $Y2=0
cc_211 N_A_137_260#_M1016_g N_VPWR_c_614_n 0.00329146f $X=1.225 $Y=2.4 $X2=0
+ $Y2=0
cc_212 N_A_137_260#_M1018_g N_VPWR_c_614_n 0.00329146f $X=1.675 $Y=2.4 $X2=0
+ $Y2=0
cc_213 N_A_137_260#_M1023_g N_VPWR_c_615_n 0.00649184f $X=2.125 $Y=2.4 $X2=0
+ $Y2=0
cc_214 N_A_137_260#_c_165_n N_VPWR_c_615_n 0.0192372f $X=3.045 $Y=1.465 $X2=0
+ $Y2=0
cc_215 N_A_137_260#_c_183_n N_VPWR_c_615_n 0.00409461f $X=3.13 $Y=1.95 $X2=0
+ $Y2=0
cc_216 N_A_137_260#_c_184_n N_VPWR_c_615_n 0.00557583f $X=3.32 $Y=2.115 $X2=0
+ $Y2=0
cc_217 N_A_137_260#_c_178_n N_VPWR_c_615_n 0.00629085f $X=2.575 $Y=1.465 $X2=0
+ $Y2=0
cc_218 N_A_137_260#_M1014_g N_VPWR_c_620_n 0.005209f $X=0.775 $Y=2.4 $X2=0 $Y2=0
cc_219 N_A_137_260#_M1016_g N_VPWR_c_620_n 0.005209f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_220 N_A_137_260#_M1018_g N_VPWR_c_622_n 0.005209f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_221 N_A_137_260#_M1023_g N_VPWR_c_622_n 0.005209f $X=2.125 $Y=2.4 $X2=0 $Y2=0
cc_222 N_A_137_260#_M1014_g N_VPWR_c_612_n 0.00986649f $X=0.775 $Y=2.4 $X2=0
+ $Y2=0
cc_223 N_A_137_260#_M1016_g N_VPWR_c_612_n 0.00982266f $X=1.225 $Y=2.4 $X2=0
+ $Y2=0
cc_224 N_A_137_260#_M1018_g N_VPWR_c_612_n 0.00982266f $X=1.675 $Y=2.4 $X2=0
+ $Y2=0
cc_225 N_A_137_260#_M1023_g N_VPWR_c_612_n 0.00987399f $X=2.125 $Y=2.4 $X2=0
+ $Y2=0
cc_226 N_A_137_260#_M1003_g N_X_c_712_n 0.0145305f $X=1.285 $Y=0.74 $X2=0 $Y2=0
cc_227 N_A_137_260#_c_165_n N_X_c_712_n 0.040362f $X=3.045 $Y=1.465 $X2=0 $Y2=0
cc_228 N_A_137_260#_c_178_n N_X_c_712_n 0.0143954f $X=2.575 $Y=1.465 $X2=0 $Y2=0
cc_229 N_A_137_260#_M1014_g N_X_c_719_n 0.0166718f $X=0.775 $Y=2.4 $X2=0 $Y2=0
cc_230 N_A_137_260#_M1014_g N_X_c_721_n 0.019068f $X=0.775 $Y=2.4 $X2=0 $Y2=0
cc_231 N_A_137_260#_M1016_g N_X_c_721_n 0.0143027f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_232 N_A_137_260#_M1018_g N_X_c_721_n 6.97946e-19 $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_233 N_A_137_260#_M1016_g N_X_c_722_n 0.012931f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_234 N_A_137_260#_M1018_g N_X_c_722_n 0.0142852f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_235 N_A_137_260#_M1023_g N_X_c_722_n 0.00373265f $X=2.125 $Y=2.4 $X2=0 $Y2=0
cc_236 N_A_137_260#_c_165_n N_X_c_722_n 0.0692143f $X=3.045 $Y=1.465 $X2=0 $Y2=0
cc_237 N_A_137_260#_c_178_n N_X_c_722_n 0.00439036f $X=2.575 $Y=1.465 $X2=0
+ $Y2=0
cc_238 N_A_137_260#_M1003_g N_X_c_714_n 3.97481e-19 $X=1.285 $Y=0.74 $X2=0 $Y2=0
cc_239 N_A_137_260#_M1010_g N_X_c_714_n 0.00845522f $X=1.715 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A_137_260#_M1020_g N_X_c_714_n 5.68006e-19 $X=2.145 $Y=0.74 $X2=0 $Y2=0
cc_241 N_A_137_260#_M1010_g N_X_c_715_n 0.0111034f $X=1.715 $Y=0.74 $X2=0 $Y2=0
cc_242 N_A_137_260#_M1020_g N_X_c_715_n 0.0120709f $X=2.145 $Y=0.74 $X2=0 $Y2=0
cc_243 N_A_137_260#_M1024_g N_X_c_715_n 2.99675e-19 $X=2.575 $Y=0.74 $X2=0 $Y2=0
cc_244 N_A_137_260#_c_165_n N_X_c_715_n 0.0598052f $X=3.045 $Y=1.465 $X2=0 $Y2=0
cc_245 N_A_137_260#_c_167_n N_X_c_715_n 8.27816e-19 $X=3.13 $Y=1.3 $X2=0 $Y2=0
cc_246 N_A_137_260#_c_178_n N_X_c_715_n 0.00470952f $X=2.575 $Y=1.465 $X2=0
+ $Y2=0
cc_247 N_A_137_260#_M1016_g N_X_c_723_n 6.97946e-19 $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_248 N_A_137_260#_M1018_g N_X_c_723_n 0.0143027f $X=1.675 $Y=2.4 $X2=0 $Y2=0
cc_249 N_A_137_260#_M1023_g N_X_c_723_n 0.0137261f $X=2.125 $Y=2.4 $X2=0 $Y2=0
cc_250 N_A_137_260#_M1010_g N_X_c_716_n 5.68006e-19 $X=1.715 $Y=0.74 $X2=0 $Y2=0
cc_251 N_A_137_260#_M1020_g N_X_c_716_n 0.00845522f $X=2.145 $Y=0.74 $X2=0 $Y2=0
cc_252 N_A_137_260#_M1024_g N_X_c_716_n 3.97481e-19 $X=2.575 $Y=0.74 $X2=0 $Y2=0
cc_253 N_A_137_260#_M1014_g N_X_c_724_n 0.00169578f $X=0.775 $Y=2.4 $X2=0 $Y2=0
cc_254 N_A_137_260#_M1016_g N_X_c_724_n 0.00135419f $X=1.225 $Y=2.4 $X2=0 $Y2=0
cc_255 N_A_137_260#_c_165_n N_X_c_724_n 0.0247465f $X=3.045 $Y=1.465 $X2=0 $Y2=0
cc_256 N_A_137_260#_c_178_n N_X_c_724_n 0.00209661f $X=2.575 $Y=1.465 $X2=0
+ $Y2=0
cc_257 N_A_137_260#_M1010_g N_X_c_717_n 9.7541e-19 $X=1.715 $Y=0.74 $X2=0 $Y2=0
cc_258 N_A_137_260#_c_165_n N_X_c_717_n 0.0209731f $X=3.045 $Y=1.465 $X2=0 $Y2=0
cc_259 N_A_137_260#_c_178_n N_X_c_717_n 0.0025465f $X=2.575 $Y=1.465 $X2=0 $Y2=0
cc_260 N_A_137_260#_M1003_g X 0.00443048f $X=1.285 $Y=0.74 $X2=0 $Y2=0
cc_261 N_A_137_260#_c_165_n X 0.0234845f $X=3.045 $Y=1.465 $X2=0 $Y2=0
cc_262 N_A_137_260#_c_178_n X 0.0186941f $X=2.575 $Y=1.465 $X2=0 $Y2=0
cc_263 N_A_137_260#_c_165_n N_A_549_392#_c_788_n 0.00954247f $X=3.045 $Y=1.465
+ $X2=0 $Y2=0
cc_264 N_A_137_260#_M1002_d N_A_549_392#_c_789_n 0.00165831f $X=3.185 $Y=1.96
+ $X2=0 $Y2=0
cc_265 N_A_137_260#_c_184_n N_A_549_392#_c_789_n 0.0117822f $X=3.32 $Y=2.115
+ $X2=0 $Y2=0
cc_266 N_A_137_260#_c_184_n N_A_549_392#_c_791_n 0.00585912f $X=3.32 $Y=2.115
+ $X2=0 $Y2=0
cc_267 N_A_137_260#_c_172_n N_A_817_392#_c_834_n 0.00663421f $X=6.51 $Y=1.195
+ $X2=0 $Y2=0
cc_268 N_A_137_260#_c_172_n N_A_1013_392#_c_862_n 0.00193826f $X=6.51 $Y=1.195
+ $X2=0 $Y2=0
cc_269 N_A_137_260#_c_172_n N_A_1013_392#_c_863_n 0.00292842f $X=6.51 $Y=1.195
+ $X2=0 $Y2=0
cc_270 N_A_137_260#_c_168_n N_VGND_M1021_s 0.00187091f $X=4.05 $Y=1.005 $X2=0
+ $Y2=0
cc_271 N_A_137_260#_M1003_g N_VGND_c_912_n 0.0112604f $X=1.285 $Y=0.74 $X2=0
+ $Y2=0
cc_272 N_A_137_260#_M1010_g N_VGND_c_912_n 5.04273e-19 $X=1.715 $Y=0.74 $X2=0
+ $Y2=0
cc_273 N_A_137_260#_M1010_g N_VGND_c_913_n 0.0017512f $X=1.715 $Y=0.74 $X2=0
+ $Y2=0
cc_274 N_A_137_260#_M1020_g N_VGND_c_913_n 0.0017512f $X=2.145 $Y=0.74 $X2=0
+ $Y2=0
cc_275 N_A_137_260#_M1020_g N_VGND_c_914_n 0.00434272f $X=2.145 $Y=0.74 $X2=0
+ $Y2=0
cc_276 N_A_137_260#_M1024_g N_VGND_c_914_n 0.00383152f $X=2.575 $Y=0.74 $X2=0
+ $Y2=0
cc_277 N_A_137_260#_M1020_g N_VGND_c_915_n 5.77606e-19 $X=2.145 $Y=0.74 $X2=0
+ $Y2=0
cc_278 N_A_137_260#_M1024_g N_VGND_c_915_n 0.0112827f $X=2.575 $Y=0.74 $X2=0
+ $Y2=0
cc_279 N_A_137_260#_c_165_n N_VGND_c_915_n 0.0133944f $X=3.045 $Y=1.465 $X2=0
+ $Y2=0
cc_280 N_A_137_260#_c_166_n N_VGND_c_915_n 0.0430526f $X=3.265 $Y=0.515 $X2=0
+ $Y2=0
cc_281 N_A_137_260#_c_174_n N_VGND_c_915_n 0.0088844f $X=3.197 $Y=1.005 $X2=0
+ $Y2=0
cc_282 N_A_137_260#_c_166_n N_VGND_c_916_n 0.013284f $X=3.265 $Y=0.515 $X2=0
+ $Y2=0
cc_283 N_A_137_260#_c_166_n N_VGND_c_917_n 0.0151524f $X=3.265 $Y=0.515 $X2=0
+ $Y2=0
cc_284 N_A_137_260#_c_168_n N_VGND_c_917_n 0.0179755f $X=4.05 $Y=1.005 $X2=0
+ $Y2=0
cc_285 N_A_137_260#_c_169_n N_VGND_c_917_n 0.0150888f $X=4.135 $Y=0.515 $X2=0
+ $Y2=0
cc_286 N_A_137_260#_c_169_n N_VGND_c_918_n 0.0219298f $X=4.135 $Y=0.515 $X2=0
+ $Y2=0
cc_287 N_A_137_260#_c_170_n N_VGND_c_918_n 0.0223605f $X=4.92 $Y=1.195 $X2=0
+ $Y2=0
cc_288 N_A_137_260#_c_171_n N_VGND_c_918_n 0.0219298f $X=5.005 $Y=0.515 $X2=0
+ $Y2=0
cc_289 N_A_137_260#_c_171_n N_VGND_c_919_n 0.0218329f $X=5.005 $Y=0.515 $X2=0
+ $Y2=0
cc_290 N_A_137_260#_c_172_n N_VGND_c_919_n 0.0232912f $X=6.51 $Y=1.195 $X2=0
+ $Y2=0
cc_291 N_A_137_260#_M1003_g N_VGND_c_923_n 0.00383152f $X=1.285 $Y=0.74 $X2=0
+ $Y2=0
cc_292 N_A_137_260#_M1010_g N_VGND_c_923_n 0.00434272f $X=1.715 $Y=0.74 $X2=0
+ $Y2=0
cc_293 N_A_137_260#_c_169_n N_VGND_c_925_n 0.00749631f $X=4.135 $Y=0.515 $X2=0
+ $Y2=0
cc_294 N_A_137_260#_c_171_n N_VGND_c_926_n 0.00749631f $X=5.005 $Y=0.515 $X2=0
+ $Y2=0
cc_295 N_A_137_260#_M1003_g N_VGND_c_929_n 0.0075754f $X=1.285 $Y=0.74 $X2=0
+ $Y2=0
cc_296 N_A_137_260#_M1010_g N_VGND_c_929_n 0.00820284f $X=1.715 $Y=0.74 $X2=0
+ $Y2=0
cc_297 N_A_137_260#_M1020_g N_VGND_c_929_n 0.00820284f $X=2.145 $Y=0.74 $X2=0
+ $Y2=0
cc_298 N_A_137_260#_M1024_g N_VGND_c_929_n 0.0075754f $X=2.575 $Y=0.74 $X2=0
+ $Y2=0
cc_299 N_A_137_260#_c_166_n N_VGND_c_929_n 0.0108098f $X=3.265 $Y=0.515 $X2=0
+ $Y2=0
cc_300 N_A_137_260#_c_169_n N_VGND_c_929_n 0.0062048f $X=4.135 $Y=0.515 $X2=0
+ $Y2=0
cc_301 N_A_137_260#_c_171_n N_VGND_c_929_n 0.0062048f $X=5.005 $Y=0.515 $X2=0
+ $Y2=0
cc_302 N_A_137_260#_c_172_n N_A_1210_74#_c_1026_n 0.0243671f $X=6.51 $Y=1.195
+ $X2=0 $Y2=0
cc_303 N_A_137_260#_M1001_d N_A_1210_74#_c_1027_n 0.00176461f $X=6.465 $Y=0.37
+ $X2=0 $Y2=0
cc_304 N_A_137_260#_c_172_n N_A_1210_74#_c_1027_n 0.00338623f $X=6.51 $Y=1.195
+ $X2=0 $Y2=0
cc_305 N_A_137_260#_c_173_n N_A_1210_74#_c_1027_n 0.0143564f $X=6.605 $Y=0.79
+ $X2=0 $Y2=0
cc_306 N_A_137_260#_c_173_n N_A_1210_74#_c_1030_n 0.0094371f $X=6.605 $Y=0.79
+ $X2=0 $Y2=0
cc_307 N_D1_M1021_g N_C1_M1004_g 0.026984f $X=3.48 $Y=0.69 $X2=0 $Y2=0
cc_308 N_D1_c_340_n N_C1_M1004_g 0.00541691f $X=3.47 $Y=1.425 $X2=0 $Y2=0
cc_309 N_D1_c_341_n N_C1_M1004_g 0.0105371f $X=3.48 $Y=1.425 $X2=0 $Y2=0
cc_310 N_D1_c_340_n C1 0.0205928f $X=3.47 $Y=1.425 $X2=0 $Y2=0
cc_311 N_D1_c_341_n C1 3.19228e-19 $X=3.48 $Y=1.425 $X2=0 $Y2=0
cc_312 N_D1_M1005_g N_C1_c_402_n 0.0345419f $X=3.545 $Y=2.46 $X2=0 $Y2=0
cc_313 N_D1_c_340_n N_C1_c_402_n 0.00144306f $X=3.47 $Y=1.425 $X2=0 $Y2=0
cc_314 N_D1_M1002_g N_VPWR_c_615_n 0.0107358f $X=3.095 $Y=2.46 $X2=0 $Y2=0
cc_315 N_D1_M1002_g N_VPWR_c_624_n 0.00333896f $X=3.095 $Y=2.46 $X2=0 $Y2=0
cc_316 N_D1_M1005_g N_VPWR_c_624_n 0.00333896f $X=3.545 $Y=2.46 $X2=0 $Y2=0
cc_317 N_D1_M1002_g N_VPWR_c_612_n 0.00427818f $X=3.095 $Y=2.46 $X2=0 $Y2=0
cc_318 N_D1_M1005_g N_VPWR_c_612_n 0.00422796f $X=3.545 $Y=2.46 $X2=0 $Y2=0
cc_319 N_D1_M1002_g N_A_549_392#_c_788_n 0.00937704f $X=3.095 $Y=2.46 $X2=0
+ $Y2=0
cc_320 N_D1_M1005_g N_A_549_392#_c_788_n 5.73047e-19 $X=3.545 $Y=2.46 $X2=0
+ $Y2=0
cc_321 N_D1_M1002_g N_A_549_392#_c_789_n 0.0116345f $X=3.095 $Y=2.46 $X2=0 $Y2=0
cc_322 N_D1_M1005_g N_A_549_392#_c_789_n 0.0116345f $X=3.545 $Y=2.46 $X2=0 $Y2=0
cc_323 N_D1_M1002_g N_A_549_392#_c_790_n 0.00291744f $X=3.095 $Y=2.46 $X2=0
+ $Y2=0
cc_324 N_D1_M1002_g N_A_549_392#_c_791_n 6.86096e-19 $X=3.095 $Y=2.46 $X2=0
+ $Y2=0
cc_325 N_D1_M1005_g N_A_549_392#_c_791_n 0.0130586f $X=3.545 $Y=2.46 $X2=0 $Y2=0
cc_326 N_D1_c_340_n N_A_549_392#_c_791_n 0.00966158f $X=3.47 $Y=1.425 $X2=0
+ $Y2=0
cc_327 N_D1_M1005_g N_A_549_392#_c_794_n 0.001916f $X=3.545 $Y=2.46 $X2=0 $Y2=0
cc_328 N_D1_M1011_g N_VGND_c_915_n 0.0034789f $X=3.05 $Y=0.69 $X2=0 $Y2=0
cc_329 N_D1_M1011_g N_VGND_c_916_n 0.00371957f $X=3.05 $Y=0.69 $X2=0 $Y2=0
cc_330 N_D1_M1021_g N_VGND_c_916_n 0.00383152f $X=3.48 $Y=0.69 $X2=0 $Y2=0
cc_331 N_D1_M1011_g N_VGND_c_917_n 4.71027e-19 $X=3.05 $Y=0.69 $X2=0 $Y2=0
cc_332 N_D1_M1021_g N_VGND_c_917_n 0.00870112f $X=3.48 $Y=0.69 $X2=0 $Y2=0
cc_333 N_D1_M1011_g N_VGND_c_929_n 0.00619993f $X=3.05 $Y=0.69 $X2=0 $Y2=0
cc_334 N_D1_M1021_g N_VGND_c_929_n 0.0075754f $X=3.48 $Y=0.69 $X2=0 $Y2=0
cc_335 N_C1_c_399_n N_B1_c_460_n 0.00859538f $X=4.36 $Y=1.085 $X2=-0.19
+ $Y2=-0.245
cc_336 N_C1_c_400_n N_B1_c_460_n 0.00368377f $X=4.36 $Y=1.235 $X2=-0.19
+ $Y2=-0.245
cc_337 N_C1_c_398_n N_B1_c_462_n 0.00368377f $X=4.37 $Y=1.45 $X2=0 $Y2=0
cc_338 C1 N_B1_c_462_n 0.00293335f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_339 C1 B1 0.0219368f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_340 C1 N_B1_c_465_n 0.00464261f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_341 N_C1_c_402_n N_B1_c_465_n 0.00337788f $X=4.445 $Y=1.615 $X2=0 $Y2=0
cc_342 N_C1_M1006_g N_VPWR_c_624_n 0.00333896f $X=3.995 $Y=2.46 $X2=0 $Y2=0
cc_343 N_C1_M1008_g N_VPWR_c_624_n 0.00333896f $X=4.445 $Y=2.46 $X2=0 $Y2=0
cc_344 N_C1_M1006_g N_VPWR_c_612_n 0.00422796f $X=3.995 $Y=2.46 $X2=0 $Y2=0
cc_345 N_C1_M1008_g N_VPWR_c_612_n 0.00427818f $X=4.445 $Y=2.46 $X2=0 $Y2=0
cc_346 N_C1_M1006_g N_A_549_392#_c_791_n 0.0141336f $X=3.995 $Y=2.46 $X2=0 $Y2=0
cc_347 N_C1_M1008_g N_A_549_392#_c_791_n 6.83772e-19 $X=4.445 $Y=2.46 $X2=0
+ $Y2=0
cc_348 N_C1_c_402_n N_A_549_392#_c_791_n 0.00239721f $X=4.445 $Y=1.615 $X2=0
+ $Y2=0
cc_349 N_C1_M1006_g N_A_549_392#_c_792_n 0.0116345f $X=3.995 $Y=2.46 $X2=0 $Y2=0
cc_350 N_C1_M1008_g N_A_549_392#_c_792_n 0.014552f $X=4.445 $Y=2.46 $X2=0 $Y2=0
cc_351 N_C1_M1006_g N_A_549_392#_c_793_n 5.73047e-19 $X=3.995 $Y=2.46 $X2=0
+ $Y2=0
cc_352 N_C1_M1008_g N_A_549_392#_c_793_n 0.00892729f $X=4.445 $Y=2.46 $X2=0
+ $Y2=0
cc_353 N_C1_M1006_g N_A_549_392#_c_794_n 0.001916f $X=3.995 $Y=2.46 $X2=0 $Y2=0
cc_354 N_C1_M1008_g N_A_817_392#_c_834_n 0.0164637f $X=4.445 $Y=2.46 $X2=0 $Y2=0
cc_355 C1 N_A_817_392#_c_834_n 0.0653606f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_356 N_C1_c_402_n N_A_817_392#_c_834_n 0.00201785f $X=4.445 $Y=1.615 $X2=0
+ $Y2=0
cc_357 C1 N_A_817_392#_c_835_n 0.0143383f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_358 N_C1_c_402_n N_A_817_392#_c_835_n 0.00233326f $X=4.445 $Y=1.615 $X2=0
+ $Y2=0
cc_359 N_C1_M1008_g N_A_1013_392#_c_861_n 5.8775e-19 $X=4.445 $Y=2.46 $X2=0
+ $Y2=0
cc_360 N_C1_M1004_g N_VGND_c_917_n 0.0084935f $X=3.92 $Y=0.69 $X2=0 $Y2=0
cc_361 N_C1_c_399_n N_VGND_c_917_n 4.44652e-19 $X=4.36 $Y=1.085 $X2=0 $Y2=0
cc_362 N_C1_M1004_g N_VGND_c_918_n 4.95643e-19 $X=3.92 $Y=0.69 $X2=0 $Y2=0
cc_363 N_C1_c_399_n N_VGND_c_918_n 0.010382f $X=4.36 $Y=1.085 $X2=0 $Y2=0
cc_364 N_C1_M1004_g N_VGND_c_925_n 0.00383152f $X=3.92 $Y=0.69 $X2=0 $Y2=0
cc_365 N_C1_c_399_n N_VGND_c_925_n 0.00383152f $X=4.36 $Y=1.085 $X2=0 $Y2=0
cc_366 N_C1_M1004_g N_VGND_c_929_n 0.0075754f $X=3.92 $Y=0.69 $X2=0 $Y2=0
cc_367 N_C1_c_399_n N_VGND_c_929_n 0.0075754f $X=4.36 $Y=1.085 $X2=0 $Y2=0
cc_368 N_B1_c_465_n N_A1_M1017_g 0.015189f $X=5.57 $Y=1.615 $X2=0 $Y2=0
cc_369 N_B1_c_465_n N_A1_M1001_g 0.0128102f $X=5.57 $Y=1.615 $X2=0 $Y2=0
cc_370 B1 A1 0.0293403f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_371 N_B1_c_465_n A1 2.76139e-19 $X=5.57 $Y=1.615 $X2=0 $Y2=0
cc_372 B1 N_A1_c_518_n 0.00295361f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_373 N_B1_c_465_n N_A1_c_518_n 0.0135315f $X=5.57 $Y=1.615 $X2=0 $Y2=0
cc_374 N_B1_M1013_g N_VPWR_c_624_n 0.00333926f $X=5.415 $Y=2.46 $X2=0 $Y2=0
cc_375 N_B1_c_467_n N_VPWR_c_624_n 0.00333926f $X=5.865 $Y=1.87 $X2=0 $Y2=0
cc_376 N_B1_M1013_g N_VPWR_c_612_n 0.0042782f $X=5.415 $Y=2.46 $X2=0 $Y2=0
cc_377 N_B1_c_467_n N_VPWR_c_612_n 0.00422798f $X=5.865 $Y=1.87 $X2=0 $Y2=0
cc_378 N_B1_M1013_g N_A_549_392#_c_792_n 5.81668e-19 $X=5.415 $Y=2.46 $X2=0
+ $Y2=0
cc_379 N_B1_M1013_g N_A_817_392#_c_834_n 0.0162693f $X=5.415 $Y=2.46 $X2=0 $Y2=0
cc_380 B1 N_A_817_392#_c_834_n 0.00496499f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_381 N_B1_M1013_g N_A_817_392#_c_836_n 0.0156043f $X=5.415 $Y=2.46 $X2=0 $Y2=0
cc_382 N_B1_c_467_n N_A_817_392#_c_836_n 0.0117517f $X=5.865 $Y=1.87 $X2=0 $Y2=0
cc_383 B1 N_A_817_392#_c_836_n 0.0275631f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_384 N_B1_c_465_n N_A_817_392#_c_836_n 0.00243055f $X=5.57 $Y=1.615 $X2=0
+ $Y2=0
cc_385 N_B1_M1013_g N_A_1013_392#_c_860_n 0.01495f $X=5.415 $Y=2.46 $X2=0 $Y2=0
cc_386 N_B1_c_467_n N_A_1013_392#_c_860_n 0.0137017f $X=5.865 $Y=1.87 $X2=0
+ $Y2=0
cc_387 B1 N_A_1013_392#_c_862_n 0.00973077f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_388 N_B1_c_460_n N_VGND_c_918_n 0.010382f $X=4.79 $Y=1.09 $X2=0 $Y2=0
cc_389 N_B1_c_463_n N_VGND_c_918_n 5.01309e-19 $X=5.22 $Y=1.09 $X2=0 $Y2=0
cc_390 N_B1_c_460_n N_VGND_c_919_n 5.01478e-19 $X=4.79 $Y=1.09 $X2=0 $Y2=0
cc_391 N_B1_c_463_n N_VGND_c_919_n 0.0114363f $X=5.22 $Y=1.09 $X2=0 $Y2=0
cc_392 N_B1_c_465_n N_VGND_c_919_n 0.00807492f $X=5.57 $Y=1.615 $X2=0 $Y2=0
cc_393 N_B1_c_460_n N_VGND_c_926_n 0.00383152f $X=4.79 $Y=1.09 $X2=0 $Y2=0
cc_394 N_B1_c_463_n N_VGND_c_926_n 0.00383152f $X=5.22 $Y=1.09 $X2=0 $Y2=0
cc_395 N_B1_c_460_n N_VGND_c_929_n 0.0075754f $X=4.79 $Y=1.09 $X2=0 $Y2=0
cc_396 N_B1_c_463_n N_VGND_c_929_n 0.0075754f $X=5.22 $Y=1.09 $X2=0 $Y2=0
cc_397 N_A1_c_518_n N_A2_M1000_g 0.0332031f $X=6.765 $Y=1.615 $X2=0 $Y2=0
cc_398 N_A1_M1012_g N_A2_M1007_g 0.0164018f $X=6.82 $Y=0.69 $X2=0 $Y2=0
cc_399 N_A1_M1012_g A2 9.03234e-19 $X=6.82 $Y=0.69 $X2=0 $Y2=0
cc_400 A1 A2 0.0291962f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_401 N_A1_c_518_n A2 2.41572e-19 $X=6.765 $Y=1.615 $X2=0 $Y2=0
cc_402 N_A1_M1012_g N_A2_c_572_n 0.010226f $X=6.82 $Y=0.69 $X2=0 $Y2=0
cc_403 A1 N_A2_c_572_n 0.0027659f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_404 N_A1_M1017_g N_VPWR_c_616_n 0.0123989f $X=6.315 $Y=2.46 $X2=0 $Y2=0
cc_405 N_A1_M1019_g N_VPWR_c_616_n 0.0130751f $X=6.765 $Y=2.46 $X2=0 $Y2=0
cc_406 N_A1_M1019_g N_VPWR_c_617_n 5.43099e-19 $X=6.765 $Y=2.46 $X2=0 $Y2=0
cc_407 N_A1_M1017_g N_VPWR_c_624_n 0.00460063f $X=6.315 $Y=2.46 $X2=0 $Y2=0
cc_408 N_A1_M1019_g N_VPWR_c_625_n 0.00460063f $X=6.765 $Y=2.46 $X2=0 $Y2=0
cc_409 N_A1_M1017_g N_VPWR_c_612_n 0.00908665f $X=6.315 $Y=2.46 $X2=0 $Y2=0
cc_410 N_A1_M1019_g N_VPWR_c_612_n 0.00908665f $X=6.765 $Y=2.46 $X2=0 $Y2=0
cc_411 N_A1_M1017_g N_A_1013_392#_c_860_n 0.00101073f $X=6.315 $Y=2.46 $X2=0
+ $Y2=0
cc_412 N_A1_M1017_g N_A_1013_392#_c_863_n 0.0150739f $X=6.315 $Y=2.46 $X2=0
+ $Y2=0
cc_413 N_A1_M1019_g N_A_1013_392#_c_863_n 0.0143228f $X=6.765 $Y=2.46 $X2=0
+ $Y2=0
cc_414 A1 N_A_1013_392#_c_863_n 0.0456455f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_415 N_A1_c_518_n N_A_1013_392#_c_863_n 0.0024356f $X=6.765 $Y=1.615 $X2=0
+ $Y2=0
cc_416 A1 N_A_1013_392#_c_868_n 0.0150385f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_417 N_A1_M1012_g N_VGND_c_920_n 3.24085e-19 $X=6.82 $Y=0.69 $X2=0 $Y2=0
cc_418 N_A1_M1001_g N_VGND_c_927_n 0.00282582f $X=6.39 $Y=0.69 $X2=0 $Y2=0
cc_419 N_A1_M1012_g N_VGND_c_927_n 0.00282606f $X=6.82 $Y=0.69 $X2=0 $Y2=0
cc_420 N_A1_M1001_g N_VGND_c_929_n 0.00359239f $X=6.39 $Y=0.69 $X2=0 $Y2=0
cc_421 N_A1_M1012_g N_VGND_c_929_n 0.00354344f $X=6.82 $Y=0.69 $X2=0 $Y2=0
cc_422 N_A1_M1001_g N_A_1210_74#_c_1026_n 0.00667566f $X=6.39 $Y=0.69 $X2=0
+ $Y2=0
cc_423 N_A1_M1012_g N_A_1210_74#_c_1026_n 4.5114e-19 $X=6.82 $Y=0.69 $X2=0 $Y2=0
cc_424 N_A1_M1001_g N_A_1210_74#_c_1027_n 0.00828071f $X=6.39 $Y=0.69 $X2=0
+ $Y2=0
cc_425 N_A1_M1012_g N_A_1210_74#_c_1027_n 0.0119714f $X=6.82 $Y=0.69 $X2=0 $Y2=0
cc_426 N_A1_M1001_g N_A_1210_74#_c_1028_n 0.00224648f $X=6.39 $Y=0.69 $X2=0
+ $Y2=0
cc_427 N_A1_M1012_g N_A_1210_74#_c_1030_n 6.58764e-19 $X=6.82 $Y=0.69 $X2=0
+ $Y2=0
cc_428 A1 N_A_1210_74#_c_1030_n 0.006568f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_429 N_A2_M1000_g N_VPWR_c_616_n 5.41206e-19 $X=7.215 $Y=2.46 $X2=0 $Y2=0
cc_430 N_A2_M1000_g N_VPWR_c_617_n 0.0124151f $X=7.215 $Y=2.46 $X2=0 $Y2=0
cc_431 N_A2_M1025_g N_VPWR_c_617_n 0.002979f $X=7.665 $Y=2.46 $X2=0 $Y2=0
cc_432 N_A2_M1000_g N_VPWR_c_625_n 0.00460063f $X=7.215 $Y=2.46 $X2=0 $Y2=0
cc_433 N_A2_M1025_g N_VPWR_c_626_n 0.005209f $X=7.665 $Y=2.46 $X2=0 $Y2=0
cc_434 N_A2_M1000_g N_VPWR_c_612_n 0.00908665f $X=7.215 $Y=2.46 $X2=0 $Y2=0
cc_435 N_A2_M1025_g N_VPWR_c_612_n 0.00985972f $X=7.665 $Y=2.46 $X2=0 $Y2=0
cc_436 N_A2_M1000_g N_A_1013_392#_c_865_n 0.0180264f $X=7.215 $Y=2.46 $X2=0
+ $Y2=0
cc_437 N_A2_M1025_g N_A_1013_392#_c_865_n 0.012931f $X=7.665 $Y=2.46 $X2=0 $Y2=0
cc_438 A2 N_A_1013_392#_c_865_n 0.0377365f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_439 N_A2_c_572_n N_A_1013_392#_c_865_n 4.03951e-19 $X=7.68 $Y=1.425 $X2=0
+ $Y2=0
cc_440 N_A2_M1025_g N_A_1013_392#_c_866_n 0.00108119f $X=7.665 $Y=2.46 $X2=0
+ $Y2=0
cc_441 A2 N_A_1013_392#_c_866_n 0.028078f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_442 N_A2_M1000_g N_A_1013_392#_c_867_n 6.74232e-19 $X=7.215 $Y=2.46 $X2=0
+ $Y2=0
cc_443 N_A2_M1025_g N_A_1013_392#_c_867_n 0.0122988f $X=7.665 $Y=2.46 $X2=0
+ $Y2=0
cc_444 N_A2_M1007_g N_VGND_c_920_n 0.00825457f $X=7.25 $Y=0.69 $X2=0 $Y2=0
cc_445 N_A2_M1027_g N_VGND_c_920_n 0.0116536f $X=7.68 $Y=0.69 $X2=0 $Y2=0
cc_446 N_A2_M1007_g N_VGND_c_927_n 0.00383152f $X=7.25 $Y=0.69 $X2=0 $Y2=0
cc_447 N_A2_M1027_g N_VGND_c_928_n 0.00383152f $X=7.68 $Y=0.69 $X2=0 $Y2=0
cc_448 N_A2_M1007_g N_VGND_c_929_n 0.00757637f $X=7.25 $Y=0.69 $X2=0 $Y2=0
cc_449 N_A2_M1027_g N_VGND_c_929_n 0.00761145f $X=7.68 $Y=0.69 $X2=0 $Y2=0
cc_450 N_A2_M1007_g N_A_1210_74#_c_1027_n 7.00191e-19 $X=7.25 $Y=0.69 $X2=0
+ $Y2=0
cc_451 N_A2_M1007_g N_A_1210_74#_c_1029_n 0.0151262f $X=7.25 $Y=0.69 $X2=0 $Y2=0
cc_452 N_A2_M1027_g N_A_1210_74#_c_1029_n 0.0138099f $X=7.68 $Y=0.69 $X2=0 $Y2=0
cc_453 A2 N_A_1210_74#_c_1029_n 0.0639085f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_454 N_A2_c_572_n N_A_1210_74#_c_1029_n 0.00443556f $X=7.68 $Y=1.425 $X2=0
+ $Y2=0
cc_455 N_A2_M1027_g N_A_1210_74#_c_1031_n 4.43891e-19 $X=7.68 $Y=0.69 $X2=0
+ $Y2=0
cc_456 N_VPWR_M1014_s N_X_c_720_n 0.00282209f $X=0.425 $Y=1.84 $X2=0 $Y2=0
cc_457 N_VPWR_c_613_n N_X_c_720_n 0.021957f $X=0.55 $Y=2.305 $X2=0 $Y2=0
cc_458 N_VPWR_c_613_n N_X_c_721_n 0.0283501f $X=0.55 $Y=2.305 $X2=0 $Y2=0
cc_459 N_VPWR_c_614_n N_X_c_721_n 0.0283117f $X=1.45 $Y=2.305 $X2=0 $Y2=0
cc_460 N_VPWR_c_620_n N_X_c_721_n 0.0144623f $X=1.365 $Y=3.33 $X2=0 $Y2=0
cc_461 N_VPWR_c_612_n N_X_c_721_n 0.0118344f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_462 N_VPWR_M1016_s N_X_c_722_n 0.00165831f $X=1.315 $Y=1.84 $X2=0 $Y2=0
cc_463 N_VPWR_c_614_n N_X_c_722_n 0.0126919f $X=1.45 $Y=2.305 $X2=0 $Y2=0
cc_464 N_VPWR_c_615_n N_X_c_722_n 0.0062222f $X=2.35 $Y=1.985 $X2=0 $Y2=0
cc_465 N_VPWR_c_614_n N_X_c_723_n 0.0283117f $X=1.45 $Y=2.305 $X2=0 $Y2=0
cc_466 N_VPWR_c_615_n N_X_c_723_n 0.0339179f $X=2.35 $Y=1.985 $X2=0 $Y2=0
cc_467 N_VPWR_c_622_n N_X_c_723_n 0.0144623f $X=2.265 $Y=3.33 $X2=0 $Y2=0
cc_468 N_VPWR_c_612_n N_X_c_723_n 0.0118344f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_469 N_VPWR_c_615_n N_A_549_392#_c_788_n 0.0463432f $X=2.35 $Y=1.985 $X2=0
+ $Y2=0
cc_470 N_VPWR_c_624_n N_A_549_392#_c_789_n 0.0357927f $X=6.375 $Y=3.33 $X2=0
+ $Y2=0
cc_471 N_VPWR_c_612_n N_A_549_392#_c_789_n 0.0200586f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_472 N_VPWR_c_615_n N_A_549_392#_c_790_n 0.0136295f $X=2.35 $Y=1.985 $X2=0
+ $Y2=0
cc_473 N_VPWR_c_624_n N_A_549_392#_c_790_n 0.0235512f $X=6.375 $Y=3.33 $X2=0
+ $Y2=0
cc_474 N_VPWR_c_612_n N_A_549_392#_c_790_n 0.0126924f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_475 N_VPWR_c_624_n N_A_549_392#_c_792_n 0.0593439f $X=6.375 $Y=3.33 $X2=0
+ $Y2=0
cc_476 N_VPWR_c_612_n N_A_549_392#_c_792_n 0.032751f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_477 N_VPWR_c_624_n N_A_549_392#_c_794_n 0.0234458f $X=6.375 $Y=3.33 $X2=0
+ $Y2=0
cc_478 N_VPWR_c_612_n N_A_549_392#_c_794_n 0.0125551f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_479 N_VPWR_c_616_n N_A_1013_392#_c_860_n 0.0103602f $X=6.54 $Y=2.4 $X2=0
+ $Y2=0
cc_480 N_VPWR_c_624_n N_A_1013_392#_c_860_n 0.0561733f $X=6.375 $Y=3.33 $X2=0
+ $Y2=0
cc_481 N_VPWR_c_612_n N_A_1013_392#_c_860_n 0.0312814f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_482 N_VPWR_c_624_n N_A_1013_392#_c_861_n 0.0200723f $X=6.375 $Y=3.33 $X2=0
+ $Y2=0
cc_483 N_VPWR_c_612_n N_A_1013_392#_c_861_n 0.0108858f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_484 N_VPWR_M1017_d N_A_1013_392#_c_863_n 0.00165831f $X=6.405 $Y=1.96 $X2=0
+ $Y2=0
cc_485 N_VPWR_c_616_n N_A_1013_392#_c_863_n 0.0170259f $X=6.54 $Y=2.4 $X2=0
+ $Y2=0
cc_486 N_VPWR_c_616_n N_A_1013_392#_c_864_n 0.0233699f $X=6.54 $Y=2.4 $X2=0
+ $Y2=0
cc_487 N_VPWR_c_617_n N_A_1013_392#_c_864_n 0.022423f $X=7.44 $Y=2.455 $X2=0
+ $Y2=0
cc_488 N_VPWR_c_625_n N_A_1013_392#_c_864_n 0.00749631f $X=7.275 $Y=3.33 $X2=0
+ $Y2=0
cc_489 N_VPWR_c_612_n N_A_1013_392#_c_864_n 0.0062048f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_490 N_VPWR_M1000_s N_A_1013_392#_c_865_n 0.00165831f $X=7.305 $Y=1.96 $X2=0
+ $Y2=0
cc_491 N_VPWR_c_617_n N_A_1013_392#_c_865_n 0.0148589f $X=7.44 $Y=2.455 $X2=0
+ $Y2=0
cc_492 N_VPWR_c_617_n N_A_1013_392#_c_867_n 0.0234083f $X=7.44 $Y=2.455 $X2=0
+ $Y2=0
cc_493 N_VPWR_c_626_n N_A_1013_392#_c_867_n 0.014549f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_494 N_VPWR_c_612_n N_A_1013_392#_c_867_n 0.0119743f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_495 N_X_c_712_n N_VGND_M1003_d 0.00328964f $X=1.415 $Y=1.045 $X2=-0.19
+ $Y2=-0.245
cc_496 N_X_c_715_n N_VGND_M1010_d 0.00176461f $X=2.195 $Y=1.045 $X2=0 $Y2=0
cc_497 N_X_c_712_n N_VGND_c_912_n 0.0219406f $X=1.415 $Y=1.045 $X2=0 $Y2=0
cc_498 N_X_c_714_n N_VGND_c_912_n 0.0164981f $X=1.5 $Y=0.515 $X2=0 $Y2=0
cc_499 N_X_c_714_n N_VGND_c_913_n 0.0157999f $X=1.5 $Y=0.515 $X2=0 $Y2=0
cc_500 N_X_c_715_n N_VGND_c_913_n 0.0135055f $X=2.195 $Y=1.045 $X2=0 $Y2=0
cc_501 N_X_c_716_n N_VGND_c_913_n 0.0157999f $X=2.36 $Y=0.515 $X2=0 $Y2=0
cc_502 N_X_c_716_n N_VGND_c_914_n 0.0109942f $X=2.36 $Y=0.515 $X2=0 $Y2=0
cc_503 N_X_c_716_n N_VGND_c_915_n 0.0216805f $X=2.36 $Y=0.515 $X2=0 $Y2=0
cc_504 N_X_c_714_n N_VGND_c_923_n 0.0109942f $X=1.5 $Y=0.515 $X2=0 $Y2=0
cc_505 N_X_c_714_n N_VGND_c_929_n 0.00904371f $X=1.5 $Y=0.515 $X2=0 $Y2=0
cc_506 N_X_c_716_n N_VGND_c_929_n 0.00904371f $X=2.36 $Y=0.515 $X2=0 $Y2=0
cc_507 N_A_549_392#_c_792_n N_A_817_392#_M1006_d 0.00165831f $X=4.505 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_508 N_A_549_392#_M1008_s N_A_817_392#_c_834_n 0.00286198f $X=4.535 $Y=1.96
+ $X2=0 $Y2=0
cc_509 N_A_549_392#_c_793_n N_A_817_392#_c_834_n 0.0219767f $X=4.67 $Y=2.455
+ $X2=0 $Y2=0
cc_510 N_A_549_392#_c_791_n N_A_817_392#_c_835_n 0.00599715f $X=3.77 $Y=2.115
+ $X2=0 $Y2=0
cc_511 N_A_549_392#_c_792_n N_A_817_392#_c_835_n 0.0118736f $X=4.505 $Y=2.99
+ $X2=0 $Y2=0
cc_512 N_A_549_392#_c_793_n N_A_1013_392#_c_859_n 0.0466988f $X=4.67 $Y=2.455
+ $X2=0 $Y2=0
cc_513 N_A_549_392#_c_792_n N_A_1013_392#_c_861_n 0.0147157f $X=4.505 $Y=2.99
+ $X2=0 $Y2=0
cc_514 N_A_817_392#_c_834_n N_A_1013_392#_M1013_s 0.00286198f $X=5.475 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_515 N_A_817_392#_c_834_n N_A_1013_392#_c_859_n 0.0198097f $X=5.475 $Y=2.035
+ $X2=0 $Y2=0
cc_516 N_A_817_392#_M1013_d N_A_1013_392#_c_860_n 0.00165831f $X=5.505 $Y=1.96
+ $X2=0 $Y2=0
cc_517 N_A_817_392#_c_836_n N_A_1013_392#_c_860_n 0.0159318f $X=5.64 $Y=2.115
+ $X2=0 $Y2=0
cc_518 N_A_817_392#_c_836_n N_A_1013_392#_c_862_n 0.00668359f $X=5.64 $Y=2.115
+ $X2=0 $Y2=0
cc_519 N_VGND_c_919_n N_A_1210_74#_c_1026_n 0.0219626f $X=5.435 $Y=0.515 $X2=0
+ $Y2=0
cc_520 N_VGND_c_920_n N_A_1210_74#_c_1027_n 0.00988046f $X=7.465 $Y=0.585 $X2=0
+ $Y2=0
cc_521 N_VGND_c_927_n N_A_1210_74#_c_1027_n 0.0425255f $X=7.3 $Y=0 $X2=0 $Y2=0
cc_522 N_VGND_c_929_n N_A_1210_74#_c_1027_n 0.0277484f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_523 N_VGND_c_919_n N_A_1210_74#_c_1028_n 0.00816634f $X=5.435 $Y=0.515 $X2=0
+ $Y2=0
cc_524 N_VGND_c_927_n N_A_1210_74#_c_1028_n 0.019738f $X=7.3 $Y=0 $X2=0 $Y2=0
cc_525 N_VGND_c_929_n N_A_1210_74#_c_1028_n 0.012511f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_526 N_VGND_M1007_s N_A_1210_74#_c_1029_n 0.00176461f $X=7.325 $Y=0.37 $X2=0
+ $Y2=0
cc_527 N_VGND_c_920_n N_A_1210_74#_c_1029_n 0.0170777f $X=7.465 $Y=0.585 $X2=0
+ $Y2=0
cc_528 N_VGND_c_920_n N_A_1210_74#_c_1031_n 0.0150645f $X=7.465 $Y=0.585 $X2=0
+ $Y2=0
cc_529 N_VGND_c_928_n N_A_1210_74#_c_1031_n 0.011066f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_530 N_VGND_c_929_n N_A_1210_74#_c_1031_n 0.00915947f $X=7.92 $Y=0 $X2=0 $Y2=0

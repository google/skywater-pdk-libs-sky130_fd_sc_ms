* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfxtp_4 CLK D VGND VNB VPB VPWR Q
M1000 VPWR a_1226_296# a_1144_508# VPB pshort w=420000u l=180000u
+  ad=2.2454e+12p pd=1.922e+07u as=1.869e+11p ps=1.73e+06u
M1001 Q a_1226_296# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1002 VGND a_1226_296# Q VNB nlowvt w=740000u l=150000u
+  ad=1.88282e+12p pd=1.54e+07u as=4.44e+11p ps=4.16e+06u
M1003 Q a_1226_296# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_1226_296# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_654_503# a_27_74# a_547_485# VPB pshort w=420000u l=180000u
+  ad=8.82e+10p pd=1.26e+06u as=1.6485e+11p ps=1.73e+06u
M1006 a_1144_508# a_209_368# a_1037_424# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=2.667e+11p ps=2.39e+06u
M1007 Q a_1226_296# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Q a_1226_296# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_440_503# D VPWR VPB pshort w=420000u l=180000u
+  ad=1.6485e+11p pd=1.73e+06u as=0p ps=0u
M1010 VPWR a_1226_296# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_696_458# a_547_485# VGND VNB nlowvt w=550000u l=150000u
+  ad=1.98e+11p pd=1.97e+06u as=0p ps=0u
M1012 VPWR CLK a_27_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1013 a_209_368# a_27_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1014 a_547_485# a_209_368# a_440_503# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1226_296# a_1037_424# VPWR VPB pshort w=840000u l=180000u
+  ad=2.268e+11p pd=2.22e+06u as=0p ps=0u
M1016 VGND a_696_458# a_735_102# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1017 VGND a_1226_296# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1037_424# a_27_74# a_696_458# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=4.2e+11p ps=2.68e+06u
M1019 VPWR a_1037_424# a_1226_296# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_1226_296# a_1178_124# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.323e+11p ps=1.47e+06u
M1021 a_735_102# a_209_368# a_547_485# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.51375e+11p ps=1.66e+06u
M1022 a_440_503# D VGND VNB nlowvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1023 a_547_485# a_27_74# a_440_503# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1037_424# a_209_368# a_696_458# VNB nlowvt w=550000u l=150000u
+  ad=2.152e+11p pd=1.97e+06u as=0p ps=0u
M1025 a_209_368# a_27_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.516e+11p pd=2.16e+06u as=0p ps=0u
M1026 VGND a_1037_424# a_1226_296# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1027 VPWR a_696_458# a_654_503# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND CLK a_27_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1029 a_696_458# a_547_485# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_1178_124# a_27_74# a_1037_424# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

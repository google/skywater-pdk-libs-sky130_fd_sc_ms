* File: sky130_fd_sc_ms__a211oi_4.pxi.spice
* Created: Fri Aug 28 16:57:43 2020
* 
x_PM_SKY130_FD_SC_MS__A211OI_4%A2 N_A2_M1006_g N_A2_M1003_g N_A2_M1009_g
+ N_A2_M1005_g N_A2_M1011_g N_A2_M1010_g N_A2_M1016_g N_A2_M1012_g A2 A2 A2 A2
+ A2 N_A2_c_118_n PM_SKY130_FD_SC_MS__A211OI_4%A2
x_PM_SKY130_FD_SC_MS__A211OI_4%A1 N_A1_M1000_g N_A1_M1020_g N_A1_M1008_g
+ N_A1_M1022_g N_A1_M1019_g N_A1_M1024_g N_A1_M1027_g N_A1_M1026_g A1 A1 A1
+ N_A1_c_203_n N_A1_c_198_n PM_SKY130_FD_SC_MS__A211OI_4%A1
x_PM_SKY130_FD_SC_MS__A211OI_4%B1 N_B1_M1007_g N_B1_M1013_g N_B1_M1017_g
+ N_B1_M1001_g N_B1_M1018_g N_B1_M1021_g B1 B1 B1 B1 N_B1_c_274_n
+ PM_SKY130_FD_SC_MS__A211OI_4%B1
x_PM_SKY130_FD_SC_MS__A211OI_4%C1 N_C1_M1014_g N_C1_M1002_g N_C1_M1015_g
+ N_C1_M1004_g N_C1_M1023_g N_C1_M1025_g C1 C1 C1 N_C1_c_346_n
+ PM_SKY130_FD_SC_MS__A211OI_4%C1
x_PM_SKY130_FD_SC_MS__A211OI_4%A_77_368# N_A_77_368#_M1006_s N_A_77_368#_M1009_s
+ N_A_77_368#_M1016_s N_A_77_368#_M1022_s N_A_77_368#_M1026_s
+ N_A_77_368#_M1007_d N_A_77_368#_M1017_d N_A_77_368#_c_405_n
+ N_A_77_368#_c_406_n N_A_77_368#_c_417_n N_A_77_368#_c_407_n
+ N_A_77_368#_c_424_n N_A_77_368#_c_408_n N_A_77_368#_c_434_n
+ N_A_77_368#_c_409_n N_A_77_368#_c_440_n N_A_77_368#_c_410_n
+ N_A_77_368#_c_411_n N_A_77_368#_c_493_p N_A_77_368#_c_451_n
+ N_A_77_368#_c_455_n N_A_77_368#_c_458_n N_A_77_368#_c_429_n
+ N_A_77_368#_c_432_n N_A_77_368#_c_445_n N_A_77_368#_c_412_n
+ N_A_77_368#_c_460_n PM_SKY130_FD_SC_MS__A211OI_4%A_77_368#
x_PM_SKY130_FD_SC_MS__A211OI_4%VPWR N_VPWR_M1006_d N_VPWR_M1011_d N_VPWR_M1020_d
+ N_VPWR_M1024_d N_VPWR_c_499_n N_VPWR_c_500_n N_VPWR_c_501_n N_VPWR_c_502_n
+ N_VPWR_c_503_n N_VPWR_c_504_n N_VPWR_c_505_n N_VPWR_c_506_n N_VPWR_c_507_n
+ VPWR N_VPWR_c_508_n N_VPWR_c_509_n N_VPWR_c_498_n N_VPWR_c_511_n
+ N_VPWR_c_512_n PM_SKY130_FD_SC_MS__A211OI_4%VPWR
x_PM_SKY130_FD_SC_MS__A211OI_4%A_901_368# N_A_901_368#_M1007_s
+ N_A_901_368#_M1013_s N_A_901_368#_M1021_s N_A_901_368#_M1004_s
+ N_A_901_368#_M1025_s N_A_901_368#_c_601_n N_A_901_368#_c_602_n
+ N_A_901_368#_c_603_n N_A_901_368#_c_617_n N_A_901_368#_c_604_n
+ N_A_901_368#_c_625_n N_A_901_368#_c_605_n N_A_901_368#_c_630_n
+ N_A_901_368#_c_606_n N_A_901_368#_c_607_n N_A_901_368#_c_608_n
+ N_A_901_368#_c_609_n N_A_901_368#_c_610_n
+ PM_SKY130_FD_SC_MS__A211OI_4%A_901_368#
x_PM_SKY130_FD_SC_MS__A211OI_4%Y N_Y_M1000_s N_Y_M1019_s N_Y_M1001_d N_Y_M1018_d
+ N_Y_M1015_s N_Y_M1002_d N_Y_M1023_d N_Y_c_676_n N_Y_c_677_n N_Y_c_678_n
+ N_Y_c_679_n N_Y_c_680_n N_Y_c_681_n N_Y_c_682_n N_Y_c_683_n N_Y_c_684_n
+ N_Y_c_685_n N_Y_c_718_n Y Y Y Y Y Y Y Y PM_SKY130_FD_SC_MS__A211OI_4%Y
x_PM_SKY130_FD_SC_MS__A211OI_4%A_92_74# N_A_92_74#_M1003_s N_A_92_74#_M1005_s
+ N_A_92_74#_M1012_s N_A_92_74#_M1008_d N_A_92_74#_M1027_d N_A_92_74#_c_749_n
+ N_A_92_74#_c_750_n N_A_92_74#_c_751_n N_A_92_74#_c_752_n N_A_92_74#_c_753_n
+ N_A_92_74#_c_754_n N_A_92_74#_c_755_n N_A_92_74#_c_756_n
+ PM_SKY130_FD_SC_MS__A211OI_4%A_92_74#
x_PM_SKY130_FD_SC_MS__A211OI_4%VGND N_VGND_M1003_d N_VGND_M1010_d N_VGND_M1001_s
+ N_VGND_M1014_d N_VGND_c_800_n N_VGND_c_801_n N_VGND_c_802_n N_VGND_c_803_n
+ N_VGND_c_804_n N_VGND_c_805_n N_VGND_c_806_n N_VGND_c_807_n VGND
+ N_VGND_c_808_n N_VGND_c_809_n N_VGND_c_810_n N_VGND_c_811_n N_VGND_c_812_n
+ N_VGND_c_813_n PM_SKY130_FD_SC_MS__A211OI_4%VGND
cc_1 VNB N_A2_M1003_g 0.0318708f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=0.74
cc_2 VNB N_A2_M1005_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=0.74
cc_3 VNB N_A2_M1010_g 0.0224899f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=0.74
cc_4 VNB N_A2_M1012_g 0.0230056f $X=-0.19 $Y=-0.245 $X2=2.09 $Y2=0.74
cc_5 VNB A2 0.0329433f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.58
cc_6 VNB N_A2_c_118_n 0.0729817f $X=-0.19 $Y=-0.245 $X2=2.09 $Y2=1.515
cc_7 VNB N_A1_M1000_g 0.0240886f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=2.4
cc_8 VNB N_A1_M1008_g 0.0234234f $X=-0.19 $Y=-0.245 $X2=1.185 $Y2=2.4
cc_9 VNB N_A1_M1019_g 0.0234256f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=2.4
cc_10 VNB N_A1_M1027_g 0.0328863f $X=-0.19 $Y=-0.245 $X2=2.085 $Y2=2.4
cc_11 VNB N_A1_c_198_n 0.0765962f $X=-0.19 $Y=-0.245 $X2=1.83 $Y2=1.515
cc_12 VNB N_B1_M1007_g 0.0017572f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=2.4
cc_13 VNB N_B1_M1013_g 0.00130001f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=0.74
cc_14 VNB N_B1_M1017_g 0.00130001f $X=-0.19 $Y=-0.245 $X2=1.185 $Y2=2.4
cc_15 VNB N_B1_M1001_g 0.0289588f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=0.74
cc_16 VNB N_B1_M1018_g 0.0208323f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=2.4
cc_17 VNB N_B1_M1021_g 0.00144367f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=0.74
cc_18 VNB B1 0.00922652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_c_274_n 0.103729f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.515
cc_20 VNB N_C1_M1014_g 0.0214f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=2.4
cc_21 VNB N_C1_M1015_g 0.0270575f $X=-0.19 $Y=-0.245 $X2=1.185 $Y2=2.4
cc_22 VNB C1 0.00375419f $X=-0.19 $Y=-0.245 $X2=2.085 $Y2=2.4
cc_23 VNB N_C1_c_346_n 0.0982692f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.515
cc_24 VNB N_VPWR_c_498_n 0.362705f $X=-0.19 $Y=-0.245 $X2=2.085 $Y2=1.515
cc_25 VNB N_Y_c_676_n 0.00622517f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=0.74
cc_26 VNB N_Y_c_677_n 0.0721116f $X=-0.19 $Y=-0.245 $X2=2.085 $Y2=2.4
cc_27 VNB N_Y_c_678_n 0.0252102f $X=-0.19 $Y=-0.245 $X2=2.09 $Y2=0.74
cc_28 VNB N_Y_c_679_n 0.00369528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_680_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_30 VNB N_Y_c_681_n 0.00306324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_682_n 0.109424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_683_n 0.00130318f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=1.515
cc_33 VNB N_Y_c_684_n 0.00180772f $X=-0.19 $Y=-0.245 $X2=1.185 $Y2=1.515
cc_34 VNB N_Y_c_685_n 0.00354475f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=1.515
cc_35 VNB N_A_92_74#_c_749_n 0.0270834f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=2.4
cc_36 VNB N_A_92_74#_c_750_n 0.00307486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_92_74#_c_751_n 0.00963497f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=1.35
cc_38 VNB N_A_92_74#_c_752_n 0.00178908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_92_74#_c_753_n 0.00917346f $X=-0.19 $Y=-0.245 $X2=2.085 $Y2=2.4
cc_40 VNB N_A_92_74#_c_754_n 0.0016059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_92_74#_c_755_n 0.0213494f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_42 VNB N_A_92_74#_c_756_n 0.00127131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_800_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.23 $Y2=0.74
cc_44 VNB N_VGND_c_801_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=2.4
cc_45 VNB N_VGND_c_802_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=0.74
cc_46 VNB N_VGND_c_803_n 0.00323505f $X=-0.19 $Y=-0.245 $X2=2.085 $Y2=2.4
cc_47 VNB N_VGND_c_804_n 0.0270966f $X=-0.19 $Y=-0.245 $X2=2.09 $Y2=0.74
cc_48 VNB N_VGND_c_805_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=2.09 $Y2=0.74
cc_49 VNB N_VGND_c_806_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_50 VNB N_VGND_c_807_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_51 VNB N_VGND_c_808_n 0.10229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_809_n 0.0151736f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.515
cc_53 VNB N_VGND_c_810_n 0.0437444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_811_n 0.517711f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_55 VNB N_VGND_c_812_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.565
cc_56 VNB N_VGND_c_813_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.565
cc_57 VPB N_A2_M1006_g 0.027583f $X=-0.19 $Y=1.66 $X2=0.735 $Y2=2.4
cc_58 VPB N_A2_M1009_g 0.0204953f $X=-0.19 $Y=1.66 $X2=1.185 $Y2=2.4
cc_59 VPB N_A2_M1011_g 0.0198955f $X=-0.19 $Y=1.66 $X2=1.635 $Y2=2.4
cc_60 VPB N_A2_M1016_g 0.0202413f $X=-0.19 $Y=1.66 $X2=2.085 $Y2=2.4
cc_61 VPB A2 0.0269007f $X=-0.19 $Y=1.66 $X2=2.075 $Y2=1.58
cc_62 VPB N_A2_c_118_n 0.0117905f $X=-0.19 $Y=1.66 $X2=2.09 $Y2=1.515
cc_63 VPB N_A1_M1020_g 0.0207996f $X=-0.19 $Y=1.66 $X2=0.8 $Y2=0.74
cc_64 VPB N_A1_M1022_g 0.0198928f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=0.74
cc_65 VPB N_A1_M1024_g 0.0198921f $X=-0.19 $Y=1.66 $X2=1.66 $Y2=0.74
cc_66 VPB N_A1_M1026_g 0.0243586f $X=-0.19 $Y=1.66 $X2=2.09 $Y2=0.74
cc_67 VPB N_A1_c_203_n 0.00755806f $X=-0.19 $Y=1.66 $X2=1.635 $Y2=1.515
cc_68 VPB N_A1_c_198_n 0.0119967f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=1.515
cc_69 VPB N_B1_M1007_g 0.0261598f $X=-0.19 $Y=1.66 $X2=0.735 $Y2=2.4
cc_70 VPB N_B1_M1013_g 0.0205757f $X=-0.19 $Y=1.66 $X2=0.8 $Y2=0.74
cc_71 VPB N_B1_M1017_g 0.0205757f $X=-0.19 $Y=1.66 $X2=1.185 $Y2=2.4
cc_72 VPB N_B1_M1021_g 0.0213856f $X=-0.19 $Y=1.66 $X2=1.66 $Y2=0.74
cc_73 VPB B1 0.0125597f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_C1_M1002_g 0.0197821f $X=-0.19 $Y=1.66 $X2=0.8 $Y2=0.74
cc_75 VPB N_C1_M1004_g 0.0196326f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=0.74
cc_76 VPB N_C1_M1023_g 0.0199998f $X=-0.19 $Y=1.66 $X2=1.635 $Y2=2.4
cc_77 VPB N_C1_M1025_g 0.0237797f $X=-0.19 $Y=1.66 $X2=1.66 $Y2=0.74
cc_78 VPB C1 0.00915857f $X=-0.19 $Y=1.66 $X2=2.085 $Y2=2.4
cc_79 VPB N_C1_c_346_n 0.0123877f $X=-0.19 $Y=1.66 $X2=0.735 $Y2=1.515
cc_80 VPB N_A_77_368#_c_405_n 0.0075508f $X=-0.19 $Y=1.66 $X2=1.66 $Y2=0.74
cc_81 VPB N_A_77_368#_c_406_n 0.0358769f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_82 VPB N_A_77_368#_c_407_n 0.00202354f $X=-0.19 $Y=1.66 $X2=2.09 $Y2=0.74
cc_83 VPB N_A_77_368#_c_408_n 0.00179594f $X=-0.19 $Y=1.66 $X2=1.595 $Y2=1.58
cc_84 VPB N_A_77_368#_c_409_n 0.00179594f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_85 VPB N_A_77_368#_c_410_n 0.0110178f $X=-0.19 $Y=1.66 $X2=0.81 $Y2=1.515
cc_86 VPB N_A_77_368#_c_411_n 0.0146646f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=1.515
cc_87 VPB N_A_77_368#_c_412_n 0.0125996f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_499_n 0.00732691f $X=-0.19 $Y=1.66 $X2=1.23 $Y2=0.74
cc_89 VPB N_VPWR_c_500_n 0.00271781f $X=-0.19 $Y=1.66 $X2=1.635 $Y2=2.4
cc_90 VPB N_VPWR_c_501_n 0.0164465f $X=-0.19 $Y=1.66 $X2=1.66 $Y2=1.35
cc_91 VPB N_VPWR_c_502_n 0.00261791f $X=-0.19 $Y=1.66 $X2=2.085 $Y2=1.68
cc_92 VPB N_VPWR_c_503_n 0.00329129f $X=-0.19 $Y=1.66 $X2=2.09 $Y2=1.35
cc_93 VPB N_VPWR_c_504_n 0.0274252f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_505_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.58
cc_95 VPB N_VPWR_c_506_n 0.0185253f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_96 VPB N_VPWR_c_507_n 0.00601644f $X=-0.19 $Y=1.66 $X2=1.115 $Y2=1.58
cc_97 VPB N_VPWR_c_508_n 0.0164465f $X=-0.19 $Y=1.66 $X2=0.8 $Y2=1.515
cc_98 VPB N_VPWR_c_509_n 0.115155f $X=-0.19 $Y=1.66 $X2=1.83 $Y2=1.515
cc_99 VPB N_VPWR_c_498_n 0.111674f $X=-0.19 $Y=1.66 $X2=2.085 $Y2=1.515
cc_100 VPB N_VPWR_c_511_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0.24 $Y2=1.565
cc_101 VPB N_VPWR_c_512_n 0.00601644f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.565
cc_102 VPB N_A_901_368#_c_601_n 0.00583793f $X=-0.19 $Y=1.66 $X2=1.635 $Y2=2.4
cc_103 VPB N_A_901_368#_c_602_n 0.00192243f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_104 VPB N_A_901_368#_c_603_n 0.00449764f $X=-0.19 $Y=1.66 $X2=1.66 $Y2=1.35
cc_105 VPB N_A_901_368#_c_604_n 0.00205771f $X=-0.19 $Y=1.66 $X2=2.085 $Y2=2.4
cc_106 VPB N_A_901_368#_c_605_n 0.00192243f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_107 VPB N_A_901_368#_c_606_n 0.0116218f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_108 VPB N_A_901_368#_c_607_n 0.030715f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_109 VPB N_A_901_368#_c_608_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0.81 $Y2=1.515
cc_110 VPB N_A_901_368#_c_609_n 0.00181992f $X=-0.19 $Y=1.66 $X2=0.81 $Y2=1.515
cc_111 VPB N_A_901_368#_c_610_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0.81 $Y2=1.515
cc_112 VPB N_Y_c_682_n 0.0206027f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_113 N_A2_M1012_g N_A1_M1000_g 0.019323f $X=2.09 $Y=0.74 $X2=0 $Y2=0
cc_114 N_A2_M1016_g N_A1_M1020_g 0.0148887f $X=2.085 $Y=2.4 $X2=0 $Y2=0
cc_115 A2 N_A1_c_203_n 0.0303407f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_116 N_A2_c_118_n N_A1_c_203_n 4.18021e-19 $X=2.09 $Y=1.515 $X2=0 $Y2=0
cc_117 A2 N_A1_c_198_n 0.00356993f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_118 N_A2_c_118_n N_A1_c_198_n 0.0148887f $X=2.09 $Y=1.515 $X2=0 $Y2=0
cc_119 N_A2_M1006_g N_A_77_368#_c_405_n 8.84614e-19 $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_120 A2 N_A_77_368#_c_405_n 0.0264312f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_121 N_A2_M1006_g N_A_77_368#_c_406_n 0.0125045f $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_122 N_A2_M1009_g N_A_77_368#_c_406_n 6.50516e-19 $X=1.185 $Y=2.4 $X2=0 $Y2=0
cc_123 N_A2_M1006_g N_A_77_368#_c_417_n 0.012931f $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_124 N_A2_M1009_g N_A_77_368#_c_417_n 0.012931f $X=1.185 $Y=2.4 $X2=0 $Y2=0
cc_125 A2 N_A_77_368#_c_417_n 0.0391869f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_126 N_A2_c_118_n N_A_77_368#_c_417_n 4.8724e-19 $X=2.09 $Y=1.515 $X2=0 $Y2=0
cc_127 N_A2_M1006_g N_A_77_368#_c_407_n 6.52999e-19 $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_128 N_A2_M1009_g N_A_77_368#_c_407_n 0.0120602f $X=1.185 $Y=2.4 $X2=0 $Y2=0
cc_129 N_A2_M1011_g N_A_77_368#_c_407_n 2.39324e-19 $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_130 N_A2_M1011_g N_A_77_368#_c_424_n 0.0142562f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_131 N_A2_M1016_g N_A_77_368#_c_424_n 0.0142562f $X=2.085 $Y=2.4 $X2=0 $Y2=0
cc_132 A2 N_A_77_368#_c_424_n 0.0478981f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_133 N_A2_c_118_n N_A_77_368#_c_424_n 4.90062e-19 $X=2.09 $Y=1.515 $X2=0 $Y2=0
cc_134 N_A2_M1016_g N_A_77_368#_c_408_n 2.33577e-19 $X=2.085 $Y=2.4 $X2=0 $Y2=0
cc_135 N_A2_M1009_g N_A_77_368#_c_429_n 8.84614e-19 $X=1.185 $Y=2.4 $X2=0 $Y2=0
cc_136 A2 N_A_77_368#_c_429_n 0.0189743f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_137 N_A2_c_118_n N_A_77_368#_c_429_n 5.52655e-19 $X=2.09 $Y=1.515 $X2=0 $Y2=0
cc_138 A2 N_A_77_368#_c_432_n 0.0041057f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_139 N_A2_M1006_g N_VPWR_c_499_n 0.0027763f $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_140 N_A2_M1009_g N_VPWR_c_499_n 0.00156821f $X=1.185 $Y=2.4 $X2=0 $Y2=0
cc_141 N_A2_M1009_g N_VPWR_c_500_n 5.60169e-19 $X=1.185 $Y=2.4 $X2=0 $Y2=0
cc_142 N_A2_M1011_g N_VPWR_c_500_n 0.0130872f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_143 N_A2_M1016_g N_VPWR_c_500_n 0.0129584f $X=2.085 $Y=2.4 $X2=0 $Y2=0
cc_144 N_A2_M1016_g N_VPWR_c_501_n 0.00460063f $X=2.085 $Y=2.4 $X2=0 $Y2=0
cc_145 N_A2_M1016_g N_VPWR_c_502_n 5.41206e-19 $X=2.085 $Y=2.4 $X2=0 $Y2=0
cc_146 N_A2_M1006_g N_VPWR_c_504_n 0.005209f $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_147 N_A2_M1009_g N_VPWR_c_506_n 0.005209f $X=1.185 $Y=2.4 $X2=0 $Y2=0
cc_148 N_A2_M1011_g N_VPWR_c_506_n 0.00460063f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_149 N_A2_M1006_g N_VPWR_c_498_n 0.00986584f $X=0.735 $Y=2.4 $X2=0 $Y2=0
cc_150 N_A2_M1009_g N_VPWR_c_498_n 0.00982266f $X=1.185 $Y=2.4 $X2=0 $Y2=0
cc_151 N_A2_M1011_g N_VPWR_c_498_n 0.00908554f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_152 N_A2_M1016_g N_VPWR_c_498_n 0.00908665f $X=2.085 $Y=2.4 $X2=0 $Y2=0
cc_153 N_A2_M1003_g N_A_92_74#_c_749_n 0.00159319f $X=0.8 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A2_M1003_g N_A_92_74#_c_750_n 0.0136535f $X=0.8 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A2_M1005_g N_A_92_74#_c_750_n 0.0130918f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_156 A2 N_A_92_74#_c_750_n 0.0517333f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_157 N_A2_c_118_n N_A_92_74#_c_750_n 0.00392608f $X=2.09 $Y=1.515 $X2=0 $Y2=0
cc_158 A2 N_A_92_74#_c_751_n 0.0224351f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_159 N_A2_c_118_n N_A_92_74#_c_751_n 6.80996e-19 $X=2.09 $Y=1.515 $X2=0 $Y2=0
cc_160 N_A2_M1005_g N_A_92_74#_c_752_n 3.92313e-19 $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_161 N_A2_M1010_g N_A_92_74#_c_752_n 3.92313e-19 $X=1.66 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A2_M1010_g N_A_92_74#_c_753_n 0.0130453f $X=1.66 $Y=0.74 $X2=0 $Y2=0
cc_163 N_A2_M1012_g N_A_92_74#_c_753_n 0.0128967f $X=2.09 $Y=0.74 $X2=0 $Y2=0
cc_164 A2 N_A_92_74#_c_753_n 0.0568851f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_165 N_A2_c_118_n N_A_92_74#_c_753_n 0.00258446f $X=2.09 $Y=1.515 $X2=0 $Y2=0
cc_166 A2 N_A_92_74#_c_756_n 0.0146029f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_167 N_A2_c_118_n N_A_92_74#_c_756_n 0.00248733f $X=2.09 $Y=1.515 $X2=0 $Y2=0
cc_168 N_A2_M1003_g N_VGND_c_800_n 0.0137191f $X=0.8 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A2_M1005_g N_VGND_c_800_n 0.0106755f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_170 N_A2_M1010_g N_VGND_c_800_n 4.71636e-19 $X=1.66 $Y=0.74 $X2=0 $Y2=0
cc_171 N_A2_M1005_g N_VGND_c_801_n 4.71636e-19 $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_172 N_A2_M1010_g N_VGND_c_801_n 0.0106755f $X=1.66 $Y=0.74 $X2=0 $Y2=0
cc_173 N_A2_M1012_g N_VGND_c_801_n 0.0107817f $X=2.09 $Y=0.74 $X2=0 $Y2=0
cc_174 N_A2_M1003_g N_VGND_c_804_n 0.00383152f $X=0.8 $Y=0.74 $X2=0 $Y2=0
cc_175 N_A2_M1005_g N_VGND_c_806_n 0.00383152f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_176 N_A2_M1010_g N_VGND_c_806_n 0.00383152f $X=1.66 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A2_M1012_g N_VGND_c_808_n 0.00383152f $X=2.09 $Y=0.74 $X2=0 $Y2=0
cc_178 N_A2_M1003_g N_VGND_c_811_n 0.00762539f $X=0.8 $Y=0.74 $X2=0 $Y2=0
cc_179 N_A2_M1005_g N_VGND_c_811_n 0.0075754f $X=1.23 $Y=0.74 $X2=0 $Y2=0
cc_180 N_A2_M1010_g N_VGND_c_811_n 0.0075754f $X=1.66 $Y=0.74 $X2=0 $Y2=0
cc_181 N_A2_M1012_g N_VGND_c_811_n 0.00757637f $X=2.09 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A1_M1027_g B1 0.00133012f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_183 N_A1_c_203_n B1 0.0148045f $X=3.69 $Y=1.515 $X2=0 $Y2=0
cc_184 N_A1_c_198_n B1 0.00937978f $X=3.885 $Y=1.515 $X2=0 $Y2=0
cc_185 N_A1_M1020_g N_A_77_368#_c_408_n 2.33577e-19 $X=2.535 $Y=2.4 $X2=0 $Y2=0
cc_186 N_A1_M1020_g N_A_77_368#_c_434_n 0.0160581f $X=2.535 $Y=2.4 $X2=0 $Y2=0
cc_187 N_A1_M1022_g N_A_77_368#_c_434_n 0.0142562f $X=2.985 $Y=2.4 $X2=0 $Y2=0
cc_188 N_A1_c_203_n N_A_77_368#_c_434_n 0.0413875f $X=3.69 $Y=1.515 $X2=0 $Y2=0
cc_189 N_A1_c_198_n N_A_77_368#_c_434_n 4.89356e-19 $X=3.885 $Y=1.515 $X2=0
+ $Y2=0
cc_190 N_A1_M1022_g N_A_77_368#_c_409_n 2.33577e-19 $X=2.985 $Y=2.4 $X2=0 $Y2=0
cc_191 N_A1_M1024_g N_A_77_368#_c_409_n 2.33577e-19 $X=3.435 $Y=2.4 $X2=0 $Y2=0
cc_192 N_A1_M1024_g N_A_77_368#_c_440_n 0.0142562f $X=3.435 $Y=2.4 $X2=0 $Y2=0
cc_193 N_A1_M1026_g N_A_77_368#_c_440_n 0.0177335f $X=3.885 $Y=2.4 $X2=0 $Y2=0
cc_194 N_A1_c_203_n N_A_77_368#_c_440_n 0.0370097f $X=3.69 $Y=1.515 $X2=0 $Y2=0
cc_195 N_A1_c_198_n N_A_77_368#_c_440_n 4.86535e-19 $X=3.885 $Y=1.515 $X2=0
+ $Y2=0
cc_196 N_A1_M1026_g N_A_77_368#_c_410_n 0.00147311f $X=3.885 $Y=2.4 $X2=0 $Y2=0
cc_197 N_A1_c_203_n N_A_77_368#_c_445_n 0.0143992f $X=3.69 $Y=1.515 $X2=0 $Y2=0
cc_198 N_A1_c_198_n N_A_77_368#_c_445_n 5.51948e-19 $X=3.885 $Y=1.515 $X2=0
+ $Y2=0
cc_199 N_A1_M1026_g N_A_77_368#_c_412_n 8.13654e-19 $X=3.885 $Y=2.4 $X2=0 $Y2=0
cc_200 N_A1_M1020_g N_VPWR_c_500_n 5.41206e-19 $X=2.535 $Y=2.4 $X2=0 $Y2=0
cc_201 N_A1_M1020_g N_VPWR_c_501_n 0.00460063f $X=2.535 $Y=2.4 $X2=0 $Y2=0
cc_202 N_A1_M1020_g N_VPWR_c_502_n 0.0129584f $X=2.535 $Y=2.4 $X2=0 $Y2=0
cc_203 N_A1_M1022_g N_VPWR_c_502_n 0.0129584f $X=2.985 $Y=2.4 $X2=0 $Y2=0
cc_204 N_A1_M1024_g N_VPWR_c_502_n 5.41206e-19 $X=3.435 $Y=2.4 $X2=0 $Y2=0
cc_205 N_A1_M1022_g N_VPWR_c_503_n 5.41206e-19 $X=2.985 $Y=2.4 $X2=0 $Y2=0
cc_206 N_A1_M1024_g N_VPWR_c_503_n 0.0129584f $X=3.435 $Y=2.4 $X2=0 $Y2=0
cc_207 N_A1_M1026_g N_VPWR_c_503_n 0.0140386f $X=3.885 $Y=2.4 $X2=0 $Y2=0
cc_208 N_A1_M1022_g N_VPWR_c_508_n 0.00460063f $X=2.985 $Y=2.4 $X2=0 $Y2=0
cc_209 N_A1_M1024_g N_VPWR_c_508_n 0.00460063f $X=3.435 $Y=2.4 $X2=0 $Y2=0
cc_210 N_A1_M1026_g N_VPWR_c_509_n 0.00460063f $X=3.885 $Y=2.4 $X2=0 $Y2=0
cc_211 N_A1_M1020_g N_VPWR_c_498_n 0.00908665f $X=2.535 $Y=2.4 $X2=0 $Y2=0
cc_212 N_A1_M1022_g N_VPWR_c_498_n 0.00908554f $X=2.985 $Y=2.4 $X2=0 $Y2=0
cc_213 N_A1_M1024_g N_VPWR_c_498_n 0.00908554f $X=3.435 $Y=2.4 $X2=0 $Y2=0
cc_214 N_A1_M1026_g N_VPWR_c_498_n 0.00913687f $X=3.885 $Y=2.4 $X2=0 $Y2=0
cc_215 N_A1_M1026_g N_A_901_368#_c_603_n 0.00186165f $X=3.885 $Y=2.4 $X2=0 $Y2=0
cc_216 N_A1_M1000_g N_Y_c_676_n 0.00450806f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_217 N_A1_M1008_g N_Y_c_676_n 0.0136469f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_218 N_A1_M1019_g N_Y_c_676_n 0.0136469f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_219 N_A1_c_203_n N_Y_c_676_n 0.0835653f $X=3.69 $Y=1.515 $X2=0 $Y2=0
cc_220 N_A1_c_198_n N_Y_c_676_n 0.00719684f $X=3.885 $Y=1.515 $X2=0 $Y2=0
cc_221 N_A1_M1027_g N_Y_c_677_n 0.0113071f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A1_c_198_n N_Y_c_677_n 0.00353991f $X=3.885 $Y=1.515 $X2=0 $Y2=0
cc_223 N_A1_M1027_g N_Y_c_683_n 0.00953159f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A1_M1000_g N_A_92_74#_c_753_n 0.0017668f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_225 N_A1_M1000_g N_A_92_74#_c_755_n 0.0146042f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_226 N_A1_M1008_g N_A_92_74#_c_755_n 0.0105399f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_227 N_A1_M1019_g N_A_92_74#_c_755_n 0.0106128f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_228 N_A1_M1027_g N_A_92_74#_c_755_n 0.0115786f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_229 N_A1_M1000_g N_VGND_c_801_n 6.39729e-19 $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_230 N_A1_M1000_g N_VGND_c_808_n 0.00291649f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_231 N_A1_M1008_g N_VGND_c_808_n 0.00291649f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_232 N_A1_M1019_g N_VGND_c_808_n 0.00291649f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A1_M1027_g N_VGND_c_808_n 0.00291649f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_234 N_A1_M1000_g N_VGND_c_811_n 0.00359219f $X=2.52 $Y=0.74 $X2=0 $Y2=0
cc_235 N_A1_M1008_g N_VGND_c_811_n 0.00359121f $X=2.95 $Y=0.74 $X2=0 $Y2=0
cc_236 N_A1_M1019_g N_VGND_c_811_n 0.00359121f $X=3.38 $Y=0.74 $X2=0 $Y2=0
cc_237 N_A1_M1027_g N_VGND_c_811_n 0.0036412f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_238 N_B1_M1018_g N_C1_M1014_g 0.0173064f $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_239 B1 N_C1_M1014_g 2.47186e-19 $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_240 N_B1_M1021_g N_C1_M1002_g 0.0180372f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_241 B1 C1 0.0284982f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_242 N_B1_c_274_n C1 0.00433573f $X=6.19 $Y=1.465 $X2=0 $Y2=0
cc_243 B1 N_C1_c_346_n 2.42588e-19 $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_244 N_B1_c_274_n N_C1_c_346_n 0.0190118f $X=6.19 $Y=1.465 $X2=0 $Y2=0
cc_245 N_B1_M1007_g N_A_77_368#_c_410_n 0.00442888f $X=4.855 $Y=2.4 $X2=0 $Y2=0
cc_246 N_B1_M1007_g N_A_77_368#_c_411_n 0.0163793f $X=4.855 $Y=2.4 $X2=0 $Y2=0
cc_247 B1 N_A_77_368#_c_411_n 0.0391524f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_248 N_B1_M1013_g N_A_77_368#_c_451_n 0.0142562f $X=5.305 $Y=2.4 $X2=0 $Y2=0
cc_249 N_B1_M1017_g N_A_77_368#_c_451_n 0.0142562f $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_250 B1 N_A_77_368#_c_451_n 0.0484052f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_251 N_B1_c_274_n N_A_77_368#_c_451_n 4.39737e-19 $X=6.19 $Y=1.465 $X2=0 $Y2=0
cc_252 N_B1_M1021_g N_A_77_368#_c_455_n 0.00341458f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_253 B1 N_A_77_368#_c_455_n 0.0167354f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_254 N_B1_c_274_n N_A_77_368#_c_455_n 4.97911e-19 $X=6.19 $Y=1.465 $X2=0 $Y2=0
cc_255 N_B1_M1021_g N_A_77_368#_c_458_n 0.00854351f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_256 N_B1_M1007_g N_A_77_368#_c_412_n 0.0034041f $X=4.855 $Y=2.4 $X2=0 $Y2=0
cc_257 B1 N_A_77_368#_c_460_n 0.0145231f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_258 N_B1_c_274_n N_A_77_368#_c_460_n 4.97911e-19 $X=6.19 $Y=1.465 $X2=0 $Y2=0
cc_259 N_B1_M1007_g N_VPWR_c_509_n 0.00333896f $X=4.855 $Y=2.4 $X2=0 $Y2=0
cc_260 N_B1_M1013_g N_VPWR_c_509_n 0.00333896f $X=5.305 $Y=2.4 $X2=0 $Y2=0
cc_261 N_B1_M1017_g N_VPWR_c_509_n 0.00333896f $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_262 N_B1_M1021_g N_VPWR_c_509_n 0.00333926f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_263 N_B1_M1007_g N_VPWR_c_498_n 0.00427818f $X=4.855 $Y=2.4 $X2=0 $Y2=0
cc_264 N_B1_M1013_g N_VPWR_c_498_n 0.00422685f $X=5.305 $Y=2.4 $X2=0 $Y2=0
cc_265 N_B1_M1017_g N_VPWR_c_498_n 0.00422685f $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_266 N_B1_M1021_g N_VPWR_c_498_n 0.00422798f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_267 N_B1_M1007_g N_A_901_368#_c_601_n 0.00953345f $X=4.855 $Y=2.4 $X2=0 $Y2=0
cc_268 N_B1_M1013_g N_A_901_368#_c_601_n 5.73047e-19 $X=5.305 $Y=2.4 $X2=0 $Y2=0
cc_269 N_B1_M1007_g N_A_901_368#_c_602_n 0.0116345f $X=4.855 $Y=2.4 $X2=0 $Y2=0
cc_270 N_B1_M1013_g N_A_901_368#_c_602_n 0.0116345f $X=5.305 $Y=2.4 $X2=0 $Y2=0
cc_271 N_B1_M1007_g N_A_901_368#_c_603_n 0.00291744f $X=4.855 $Y=2.4 $X2=0 $Y2=0
cc_272 N_B1_M1007_g N_A_901_368#_c_617_n 5.73047e-19 $X=4.855 $Y=2.4 $X2=0 $Y2=0
cc_273 N_B1_M1013_g N_A_901_368#_c_617_n 0.00951061f $X=5.305 $Y=2.4 $X2=0 $Y2=0
cc_274 N_B1_M1017_g N_A_901_368#_c_617_n 0.00963732f $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_275 N_B1_M1021_g N_A_901_368#_c_617_n 6.18421e-19 $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_276 N_B1_M1017_g N_A_901_368#_c_604_n 0.0116345f $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_277 N_B1_M1021_g N_A_901_368#_c_604_n 0.0139961f $X=6.205 $Y=2.4 $X2=0 $Y2=0
cc_278 N_B1_M1013_g N_A_901_368#_c_608_n 0.00194226f $X=5.305 $Y=2.4 $X2=0 $Y2=0
cc_279 N_B1_M1017_g N_A_901_368#_c_608_n 0.00194226f $X=5.755 $Y=2.4 $X2=0 $Y2=0
cc_280 B1 N_Y_c_677_n 0.0736923f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_281 N_B1_c_274_n N_Y_c_677_n 0.0158549f $X=6.19 $Y=1.465 $X2=0 $Y2=0
cc_282 N_B1_M1001_g N_Y_c_678_n 0.00159319f $X=5.76 $Y=0.74 $X2=0 $Y2=0
cc_283 N_B1_M1001_g N_Y_c_679_n 0.012695f $X=5.76 $Y=0.74 $X2=0 $Y2=0
cc_284 N_B1_M1018_g N_Y_c_679_n 0.0170661f $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_285 B1 N_Y_c_679_n 0.036928f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_286 N_B1_c_274_n N_Y_c_679_n 0.0049477f $X=6.19 $Y=1.465 $X2=0 $Y2=0
cc_287 N_B1_M1018_g N_Y_c_680_n 3.92313e-19 $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_288 B1 N_Y_c_684_n 0.0216392f $X=5.915 $Y=1.58 $X2=0 $Y2=0
cc_289 N_B1_c_274_n N_Y_c_684_n 0.00645498f $X=6.19 $Y=1.465 $X2=0 $Y2=0
cc_290 N_B1_M1018_g N_Y_c_685_n 0.00158218f $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_291 N_B1_M1001_g N_VGND_c_802_n 0.0125716f $X=5.76 $Y=0.74 $X2=0 $Y2=0
cc_292 N_B1_M1018_g N_VGND_c_802_n 0.00955691f $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_293 N_B1_M1018_g N_VGND_c_803_n 4.71636e-19 $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_294 N_B1_M1001_g N_VGND_c_808_n 0.00383152f $X=5.76 $Y=0.74 $X2=0 $Y2=0
cc_295 N_B1_M1018_g N_VGND_c_809_n 0.00383152f $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_296 N_B1_M1001_g N_VGND_c_811_n 0.00762539f $X=5.76 $Y=0.74 $X2=0 $Y2=0
cc_297 N_B1_M1018_g N_VGND_c_811_n 0.00757637f $X=6.19 $Y=0.74 $X2=0 $Y2=0
cc_298 N_C1_M1002_g N_VPWR_c_509_n 0.00333896f $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_299 N_C1_M1004_g N_VPWR_c_509_n 0.00333896f $X=7.105 $Y=2.4 $X2=0 $Y2=0
cc_300 N_C1_M1023_g N_VPWR_c_509_n 0.00333896f $X=7.555 $Y=2.4 $X2=0 $Y2=0
cc_301 N_C1_M1025_g N_VPWR_c_509_n 0.00333896f $X=8.005 $Y=2.4 $X2=0 $Y2=0
cc_302 N_C1_M1002_g N_VPWR_c_498_n 0.00422796f $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_303 N_C1_M1004_g N_VPWR_c_498_n 0.00422685f $X=7.105 $Y=2.4 $X2=0 $Y2=0
cc_304 N_C1_M1023_g N_VPWR_c_498_n 0.00422685f $X=7.555 $Y=2.4 $X2=0 $Y2=0
cc_305 N_C1_M1025_g N_VPWR_c_498_n 0.00426801f $X=8.005 $Y=2.4 $X2=0 $Y2=0
cc_306 N_C1_M1002_g N_A_901_368#_c_625_n 0.0129423f $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_307 N_C1_M1004_g N_A_901_368#_c_625_n 6.28485e-19 $X=7.105 $Y=2.4 $X2=0 $Y2=0
cc_308 C1 N_A_901_368#_c_625_n 0.0174392f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_309 N_C1_M1002_g N_A_901_368#_c_605_n 0.0116345f $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_310 N_C1_M1004_g N_A_901_368#_c_605_n 0.0116345f $X=7.105 $Y=2.4 $X2=0 $Y2=0
cc_311 N_C1_M1002_g N_A_901_368#_c_630_n 5.73047e-19 $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_312 N_C1_M1004_g N_A_901_368#_c_630_n 0.00892729f $X=7.105 $Y=2.4 $X2=0 $Y2=0
cc_313 N_C1_M1023_g N_A_901_368#_c_630_n 0.00892729f $X=7.555 $Y=2.4 $X2=0 $Y2=0
cc_314 N_C1_M1025_g N_A_901_368#_c_630_n 5.73047e-19 $X=8.005 $Y=2.4 $X2=0 $Y2=0
cc_315 N_C1_M1023_g N_A_901_368#_c_606_n 0.0116345f $X=7.555 $Y=2.4 $X2=0 $Y2=0
cc_316 N_C1_M1025_g N_A_901_368#_c_606_n 0.014552f $X=8.005 $Y=2.4 $X2=0 $Y2=0
cc_317 N_C1_M1023_g N_A_901_368#_c_607_n 5.99467e-19 $X=7.555 $Y=2.4 $X2=0 $Y2=0
cc_318 N_C1_M1025_g N_A_901_368#_c_607_n 0.013348f $X=8.005 $Y=2.4 $X2=0 $Y2=0
cc_319 N_C1_M1002_g N_A_901_368#_c_609_n 0.001916f $X=6.655 $Y=2.4 $X2=0 $Y2=0
cc_320 N_C1_M1004_g N_A_901_368#_c_610_n 0.00194226f $X=7.105 $Y=2.4 $X2=0 $Y2=0
cc_321 N_C1_M1023_g N_A_901_368#_c_610_n 0.00194226f $X=7.555 $Y=2.4 $X2=0 $Y2=0
cc_322 N_C1_M1014_g N_Y_c_680_n 3.92313e-19 $X=6.62 $Y=0.74 $X2=0 $Y2=0
cc_323 N_C1_M1014_g N_Y_c_681_n 0.0129459f $X=6.62 $Y=0.74 $X2=0 $Y2=0
cc_324 N_C1_M1015_g N_Y_c_681_n 0.0139042f $X=7.05 $Y=0.74 $X2=0 $Y2=0
cc_325 C1 N_Y_c_681_n 0.0519673f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_326 N_C1_c_346_n N_Y_c_681_n 0.00404583f $X=8.005 $Y=1.5 $X2=0 $Y2=0
cc_327 N_C1_M1015_g N_Y_c_682_n 0.00528327f $X=7.05 $Y=0.74 $X2=0 $Y2=0
cc_328 N_C1_M1004_g N_Y_c_682_n 0.0142175f $X=7.105 $Y=2.4 $X2=0 $Y2=0
cc_329 N_C1_M1023_g N_Y_c_682_n 0.0226851f $X=7.555 $Y=2.4 $X2=0 $Y2=0
cc_330 N_C1_M1025_g N_Y_c_682_n 0.0205449f $X=8.005 $Y=2.4 $X2=0 $Y2=0
cc_331 C1 N_Y_c_682_n 0.10804f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_332 N_C1_c_346_n N_Y_c_682_n 0.05745f $X=8.005 $Y=1.5 $X2=0 $Y2=0
cc_333 C1 N_Y_c_685_n 0.011271f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_334 C1 N_Y_c_718_n 0.0143992f $X=7.355 $Y=1.58 $X2=0 $Y2=0
cc_335 N_C1_c_346_n N_Y_c_718_n 5.51551e-19 $X=8.005 $Y=1.5 $X2=0 $Y2=0
cc_336 N_C1_M1014_g N_VGND_c_802_n 4.56715e-19 $X=6.62 $Y=0.74 $X2=0 $Y2=0
cc_337 N_C1_M1014_g N_VGND_c_803_n 0.0106755f $X=6.62 $Y=0.74 $X2=0 $Y2=0
cc_338 N_C1_M1015_g N_VGND_c_803_n 0.0137064f $X=7.05 $Y=0.74 $X2=0 $Y2=0
cc_339 N_C1_M1014_g N_VGND_c_809_n 0.00383152f $X=6.62 $Y=0.74 $X2=0 $Y2=0
cc_340 N_C1_M1015_g N_VGND_c_810_n 0.00383152f $X=7.05 $Y=0.74 $X2=0 $Y2=0
cc_341 N_C1_M1014_g N_VGND_c_811_n 0.00757637f $X=6.62 $Y=0.74 $X2=0 $Y2=0
cc_342 N_C1_M1015_g N_VGND_c_811_n 0.00762539f $X=7.05 $Y=0.74 $X2=0 $Y2=0
cc_343 N_A_77_368#_c_417_n N_VPWR_M1006_d 0.00314376f $X=1.245 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_344 N_A_77_368#_c_424_n N_VPWR_M1011_d 0.00314376f $X=2.225 $Y=2.035 $X2=0
+ $Y2=0
cc_345 N_A_77_368#_c_434_n N_VPWR_M1020_d 0.00314376f $X=3.125 $Y=2.035 $X2=0
+ $Y2=0
cc_346 N_A_77_368#_c_440_n N_VPWR_M1024_d 0.00314376f $X=4.025 $Y=2.035 $X2=0
+ $Y2=0
cc_347 N_A_77_368#_c_406_n N_VPWR_c_499_n 0.0233699f $X=0.51 $Y=2.815 $X2=0
+ $Y2=0
cc_348 N_A_77_368#_c_417_n N_VPWR_c_499_n 0.0126919f $X=1.245 $Y=2.035 $X2=0
+ $Y2=0
cc_349 N_A_77_368#_c_407_n N_VPWR_c_499_n 0.022423f $X=1.41 $Y=2.445 $X2=0 $Y2=0
cc_350 N_A_77_368#_c_407_n N_VPWR_c_500_n 0.0234083f $X=1.41 $Y=2.445 $X2=0
+ $Y2=0
cc_351 N_A_77_368#_c_424_n N_VPWR_c_500_n 0.0170259f $X=2.225 $Y=2.035 $X2=0
+ $Y2=0
cc_352 N_A_77_368#_c_408_n N_VPWR_c_500_n 0.0233699f $X=2.31 $Y=2.445 $X2=0
+ $Y2=0
cc_353 N_A_77_368#_c_408_n N_VPWR_c_501_n 0.00749631f $X=2.31 $Y=2.445 $X2=0
+ $Y2=0
cc_354 N_A_77_368#_c_408_n N_VPWR_c_502_n 0.0233699f $X=2.31 $Y=2.445 $X2=0
+ $Y2=0
cc_355 N_A_77_368#_c_434_n N_VPWR_c_502_n 0.0170259f $X=3.125 $Y=2.035 $X2=0
+ $Y2=0
cc_356 N_A_77_368#_c_409_n N_VPWR_c_502_n 0.0233699f $X=3.21 $Y=2.445 $X2=0
+ $Y2=0
cc_357 N_A_77_368#_c_409_n N_VPWR_c_503_n 0.0233699f $X=3.21 $Y=2.445 $X2=0
+ $Y2=0
cc_358 N_A_77_368#_c_440_n N_VPWR_c_503_n 0.0170259f $X=4.025 $Y=2.035 $X2=0
+ $Y2=0
cc_359 N_A_77_368#_c_410_n N_VPWR_c_503_n 0.0234083f $X=4.11 $Y=2.4 $X2=0 $Y2=0
cc_360 N_A_77_368#_c_406_n N_VPWR_c_504_n 0.014549f $X=0.51 $Y=2.815 $X2=0 $Y2=0
cc_361 N_A_77_368#_c_407_n N_VPWR_c_506_n 0.0109793f $X=1.41 $Y=2.445 $X2=0
+ $Y2=0
cc_362 N_A_77_368#_c_409_n N_VPWR_c_508_n 0.00749631f $X=3.21 $Y=2.445 $X2=0
+ $Y2=0
cc_363 N_A_77_368#_c_410_n N_VPWR_c_509_n 0.011066f $X=4.11 $Y=2.4 $X2=0 $Y2=0
cc_364 N_A_77_368#_c_406_n N_VPWR_c_498_n 0.0119743f $X=0.51 $Y=2.815 $X2=0
+ $Y2=0
cc_365 N_A_77_368#_c_407_n N_VPWR_c_498_n 0.00901959f $X=1.41 $Y=2.445 $X2=0
+ $Y2=0
cc_366 N_A_77_368#_c_408_n N_VPWR_c_498_n 0.0062048f $X=2.31 $Y=2.445 $X2=0
+ $Y2=0
cc_367 N_A_77_368#_c_409_n N_VPWR_c_498_n 0.0062048f $X=3.21 $Y=2.445 $X2=0
+ $Y2=0
cc_368 N_A_77_368#_c_410_n N_VPWR_c_498_n 0.00915947f $X=4.11 $Y=2.4 $X2=0 $Y2=0
cc_369 N_A_77_368#_c_411_n N_A_901_368#_M1007_s 0.00506503f $X=4.995 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_370 N_A_77_368#_c_451_n N_A_901_368#_M1013_s 0.00315967f $X=5.895 $Y=2.035
+ $X2=0 $Y2=0
cc_371 N_A_77_368#_c_410_n N_A_901_368#_c_601_n 0.0463432f $X=4.11 $Y=2.4 $X2=0
+ $Y2=0
cc_372 N_A_77_368#_c_411_n N_A_901_368#_c_601_n 0.0219767f $X=4.995 $Y=2.035
+ $X2=0 $Y2=0
cc_373 N_A_77_368#_M1007_d N_A_901_368#_c_602_n 0.00165831f $X=4.945 $Y=1.84
+ $X2=0 $Y2=0
cc_374 N_A_77_368#_c_493_p N_A_901_368#_c_602_n 0.0118736f $X=5.08 $Y=2.57 $X2=0
+ $Y2=0
cc_375 N_A_77_368#_c_410_n N_A_901_368#_c_603_n 0.00601303f $X=4.11 $Y=2.4 $X2=0
+ $Y2=0
cc_376 N_A_77_368#_c_451_n N_A_901_368#_c_617_n 0.0170259f $X=5.895 $Y=2.035
+ $X2=0 $Y2=0
cc_377 N_A_77_368#_M1017_d N_A_901_368#_c_604_n 0.00165831f $X=5.845 $Y=1.84
+ $X2=0 $Y2=0
cc_378 N_A_77_368#_c_458_n N_A_901_368#_c_604_n 0.0139027f $X=5.98 $Y=2.57 $X2=0
+ $Y2=0
cc_379 N_VPWR_c_509_n N_A_901_368#_c_602_n 0.0357927f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_380 N_VPWR_c_498_n N_A_901_368#_c_602_n 0.0200586f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_381 N_VPWR_c_503_n N_A_901_368#_c_603_n 0.00293392f $X=3.66 $Y=2.41 $X2=0
+ $Y2=0
cc_382 N_VPWR_c_509_n N_A_901_368#_c_603_n 0.0235512f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_383 N_VPWR_c_498_n N_A_901_368#_c_603_n 0.0126924f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_384 N_VPWR_c_509_n N_A_901_368#_c_604_n 0.0389233f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_385 N_VPWR_c_498_n N_A_901_368#_c_604_n 0.0218015f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_386 N_VPWR_c_509_n N_A_901_368#_c_605_n 0.0357927f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_387 N_VPWR_c_498_n N_A_901_368#_c_605_n 0.0200586f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_388 N_VPWR_c_509_n N_A_901_368#_c_606_n 0.0593439f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_389 N_VPWR_c_498_n N_A_901_368#_c_606_n 0.032751f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_390 N_VPWR_c_509_n N_A_901_368#_c_608_n 0.0234458f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_391 N_VPWR_c_498_n N_A_901_368#_c_608_n 0.0125551f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_392 N_VPWR_c_509_n N_A_901_368#_c_609_n 0.0199669f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_393 N_VPWR_c_498_n N_A_901_368#_c_609_n 0.0107485f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_394 N_VPWR_c_509_n N_A_901_368#_c_610_n 0.0234458f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_395 N_VPWR_c_498_n N_A_901_368#_c_610_n 0.0125551f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_396 N_A_901_368#_c_605_n N_Y_M1002_d 0.00165831f $X=7.165 $Y=2.99 $X2=0 $Y2=0
cc_397 N_A_901_368#_c_606_n N_Y_M1023_d 0.00165831f $X=8.065 $Y=2.99 $X2=0 $Y2=0
cc_398 N_A_901_368#_M1004_s N_Y_c_682_n 0.00314376f $X=7.195 $Y=1.84 $X2=0 $Y2=0
cc_399 N_A_901_368#_M1025_s N_Y_c_682_n 0.00273353f $X=8.095 $Y=1.84 $X2=0 $Y2=0
cc_400 N_A_901_368#_c_630_n N_Y_c_682_n 0.0170259f $X=7.33 $Y=2.455 $X2=0 $Y2=0
cc_401 N_A_901_368#_c_606_n N_Y_c_682_n 0.0118736f $X=8.065 $Y=2.99 $X2=0 $Y2=0
cc_402 N_A_901_368#_c_607_n N_Y_c_682_n 0.0243696f $X=8.23 $Y=2.285 $X2=0 $Y2=0
cc_403 N_A_901_368#_c_605_n N_Y_c_718_n 0.0118736f $X=7.165 $Y=2.99 $X2=0 $Y2=0
cc_404 N_Y_c_676_n N_A_92_74#_M1008_d 0.00177483f $X=3.588 $Y=0.957 $X2=0 $Y2=0
cc_405 N_Y_c_677_n N_A_92_74#_M1027_d 0.00425265f $X=5.38 $Y=1.045 $X2=0 $Y2=0
cc_406 N_Y_c_676_n N_A_92_74#_c_753_n 0.00561736f $X=3.588 $Y=0.957 $X2=0 $Y2=0
cc_407 N_Y_M1000_s N_A_92_74#_c_755_n 0.00179328f $X=2.595 $Y=0.37 $X2=0 $Y2=0
cc_408 N_Y_M1019_s N_A_92_74#_c_755_n 0.00179328f $X=3.455 $Y=0.37 $X2=0 $Y2=0
cc_409 N_Y_c_676_n N_A_92_74#_c_755_n 0.0630655f $X=3.588 $Y=0.957 $X2=0 $Y2=0
cc_410 N_Y_c_677_n N_A_92_74#_c_755_n 0.0160707f $X=5.38 $Y=1.045 $X2=0 $Y2=0
cc_411 N_Y_c_679_n N_VGND_M1001_s 0.00176461f $X=6.32 $Y=1.045 $X2=0 $Y2=0
cc_412 N_Y_c_681_n N_VGND_M1014_d 0.00176461f $X=7.18 $Y=1.095 $X2=0 $Y2=0
cc_413 N_Y_c_678_n N_VGND_c_802_n 0.0164982f $X=5.545 $Y=0.515 $X2=0 $Y2=0
cc_414 N_Y_c_679_n N_VGND_c_802_n 0.0170777f $X=6.32 $Y=1.045 $X2=0 $Y2=0
cc_415 N_Y_c_680_n N_VGND_c_802_n 0.0164567f $X=6.405 $Y=0.515 $X2=0 $Y2=0
cc_416 N_Y_c_680_n N_VGND_c_803_n 0.0182488f $X=6.405 $Y=0.515 $X2=0 $Y2=0
cc_417 N_Y_c_681_n N_VGND_c_803_n 0.0170777f $X=7.18 $Y=1.095 $X2=0 $Y2=0
cc_418 N_Y_c_682_n N_VGND_c_803_n 0.0184913f $X=7.695 $Y=2.035 $X2=0 $Y2=0
cc_419 N_Y_c_678_n N_VGND_c_808_n 0.011066f $X=5.545 $Y=0.515 $X2=0 $Y2=0
cc_420 N_Y_c_680_n N_VGND_c_809_n 0.00749631f $X=6.405 $Y=0.515 $X2=0 $Y2=0
cc_421 N_Y_c_682_n N_VGND_c_810_n 0.0595689f $X=7.695 $Y=2.035 $X2=0 $Y2=0
cc_422 N_Y_c_678_n N_VGND_c_811_n 0.00915947f $X=5.545 $Y=0.515 $X2=0 $Y2=0
cc_423 N_Y_c_680_n N_VGND_c_811_n 0.0062048f $X=6.405 $Y=0.515 $X2=0 $Y2=0
cc_424 N_Y_c_682_n N_VGND_c_811_n 0.049306f $X=7.695 $Y=2.035 $X2=0 $Y2=0
cc_425 N_A_92_74#_c_750_n N_VGND_M1003_d 0.00176461f $X=1.36 $Y=1.095 $X2=-0.19
+ $Y2=-0.245
cc_426 N_A_92_74#_c_753_n N_VGND_M1010_d 0.00176461f $X=2.22 $Y=1.095 $X2=0
+ $Y2=0
cc_427 N_A_92_74#_c_749_n N_VGND_c_800_n 0.0182902f $X=0.585 $Y=0.515 $X2=0
+ $Y2=0
cc_428 N_A_92_74#_c_750_n N_VGND_c_800_n 0.0170777f $X=1.36 $Y=1.095 $X2=0 $Y2=0
cc_429 N_A_92_74#_c_752_n N_VGND_c_800_n 0.0182488f $X=1.445 $Y=0.515 $X2=0
+ $Y2=0
cc_430 N_A_92_74#_c_752_n N_VGND_c_801_n 0.0182488f $X=1.445 $Y=0.515 $X2=0
+ $Y2=0
cc_431 N_A_92_74#_c_753_n N_VGND_c_801_n 0.0170777f $X=2.22 $Y=1.095 $X2=0 $Y2=0
cc_432 N_A_92_74#_c_754_n N_VGND_c_801_n 0.0103909f $X=2.305 $Y=0.615 $X2=0
+ $Y2=0
cc_433 N_A_92_74#_c_749_n N_VGND_c_804_n 0.011066f $X=0.585 $Y=0.515 $X2=0 $Y2=0
cc_434 N_A_92_74#_c_752_n N_VGND_c_806_n 0.00749631f $X=1.445 $Y=0.515 $X2=0
+ $Y2=0
cc_435 N_A_92_74#_c_754_n N_VGND_c_808_n 0.00758556f $X=2.305 $Y=0.615 $X2=0
+ $Y2=0
cc_436 N_A_92_74#_c_755_n N_VGND_c_808_n 0.0732318f $X=4.025 $Y=0.515 $X2=0
+ $Y2=0
cc_437 N_A_92_74#_c_749_n N_VGND_c_811_n 0.00915947f $X=0.585 $Y=0.515 $X2=0
+ $Y2=0
cc_438 N_A_92_74#_c_752_n N_VGND_c_811_n 0.0062048f $X=1.445 $Y=0.515 $X2=0
+ $Y2=0
cc_439 N_A_92_74#_c_754_n N_VGND_c_811_n 0.00627867f $X=2.305 $Y=0.615 $X2=0
+ $Y2=0
cc_440 N_A_92_74#_c_755_n N_VGND_c_811_n 0.0615843f $X=4.025 $Y=0.515 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__xor2_1.pex.spice
* Created: Fri Aug 28 18:18:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__XOR2_1%B 1 3 6 10 14 19 21 27 28 32
c69 32 0 6.81261e-20 $X=2.515 $Y=1.565
c70 28 0 1.31541e-19 $X=2.68 $Y=1.515
c71 14 0 1.72297e-19 $X=2.755 $Y=2.4
r72 27 30 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.515
+ $X2=2.68 $Y2=1.68
r73 27 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.515
+ $X2=2.68 $Y2=1.35
r74 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.515 $X2=2.68 $Y2=1.515
r75 21 28 1.07204 $w=4.28e-07 $l=4e-08 $layer=LI1_cond $X=2.64 $Y=1.565 $X2=2.68
+ $Y2=1.565
r76 21 32 4.00257 $w=4.28e-07 $l=1.25e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.515 $Y2=1.565
r77 19 25 38.4319 $w=3.01e-07 $l=2.4e-07 $layer=POLY_cond $X=1.45 $Y=1.605
+ $X2=1.69 $Y2=1.605
r78 18 32 37.1925 $w=3.28e-07 $l=1.065e-06 $layer=LI1_cond $X=1.45 $Y=1.53
+ $X2=2.515 $Y2=1.53
r79 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.45
+ $Y=1.53 $X2=1.45 $Y2=1.53
r80 14 30 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.755 $Y=2.4
+ $X2=2.755 $Y2=1.68
r81 10 29 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.59 $Y=0.805
+ $X2=2.59 $Y2=1.35
r82 4 25 19.0468 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.69 $Y=1.365
+ $X2=1.69 $Y2=1.605
r83 4 6 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.69 $Y=1.365
+ $X2=1.69 $Y2=0.9
r84 1 19 50.4419 $w=3.01e-07 $l=4.18121e-07 $layer=POLY_cond $X=1.135 $Y=1.845
+ $X2=1.45 $Y2=1.605
r85 1 3 164.683 $w=1.8e-07 $l=6.15e-07 $layer=POLY_cond $X=1.135 $Y=1.845
+ $X2=1.135 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__XOR2_1%A 1 3 8 9 10 11 13 18 20 22 26
c56 18 0 1.05828e-19 $X=2.2 $Y=0.805
c57 1 0 6.81261e-20 $X=0.715 $Y=1.765
r58 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.45 $X2=0.61 $Y2=1.45
r59 22 26 9.80239 $w=4.33e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.397
+ $X2=0.61 $Y2=1.397
r60 20 25 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.625 $Y=1.45
+ $X2=0.61 $Y2=1.45
r61 18 21 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.2 $Y=0.805
+ $X2=2.2 $Y2=1.25
r62 15 18 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.2 $Y=0.255 $X2=2.2
+ $Y2=0.805
r63 11 21 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.185 $Y=1.34
+ $X2=2.185 $Y2=1.25
r64 11 13 412.032 $w=1.8e-07 $l=1.06e-06 $layer=POLY_cond $X=2.185 $Y=1.34
+ $X2=2.185 $Y2=2.4
r65 9 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.125 $Y=0.18
+ $X2=2.2 $Y2=0.255
r66 9 10 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=2.125 $Y=0.18
+ $X2=0.97 $Y2=0.18
r67 6 20 41.3672 $w=2.16e-07 $l=2.16852e-07 $layer=POLY_cond $X=0.895 $Y=1.285
+ $X2=0.775 $Y2=1.45
r68 6 8 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.895 $Y=1.285
+ $X2=0.895 $Y2=0.9
r69 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.895 $Y=0.255
+ $X2=0.97 $Y2=0.18
r70 5 8 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=0.895 $Y=0.255
+ $X2=0.895 $Y2=0.9
r71 1 20 71.7726 $w=2.16e-07 $l=3.43693e-07 $layer=POLY_cond $X=0.715 $Y=1.765
+ $X2=0.775 $Y2=1.45
r72 1 3 270.153 $w=1.8e-07 $l=6.95e-07 $layer=POLY_cond $X=0.715 $Y=1.765
+ $X2=0.715 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__XOR2_1%A_194_125# 1 2 9 13 16 19 21 23 25 28 30 34
+ 35
c87 35 0 1.71893e-19 $X=3.25 $Y=1.485
c88 23 0 1.05828e-19 $X=1.475 $Y=0.875
c89 13 0 1.31541e-19 $X=3.255 $Y=2.4
r90 35 39 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=1.485
+ $X2=3.25 $Y2=1.65
r91 35 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.25 $Y=1.485
+ $X2=3.25 $Y2=1.32
r92 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.25
+ $Y=1.485 $X2=3.25 $Y2=1.485
r93 31 34 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=3.11 $Y=1.485
+ $X2=3.25 $Y2=1.485
r94 27 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.11 $Y=1.65
+ $X2=3.11 $Y2=1.485
r95 27 28 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.11 $Y=1.65 $X2=3.11
+ $Y2=1.95
r96 26 30 4.29663 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=1.525 $Y=2.035
+ $X2=1.235 $Y2=2.035
r97 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.025 $Y=2.035
+ $X2=3.11 $Y2=1.95
r98 25 26 97.861 $w=1.68e-07 $l=1.5e-06 $layer=LI1_cond $X=3.025 $Y=2.035
+ $X2=1.525 $Y2=2.035
r99 21 23 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.115 $Y=0.875
+ $X2=1.475 $Y2=0.875
r100 17 30 2.56749 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=2.12
+ $X2=1.235 $Y2=2.035
r101 17 19 14.3323 $w=5.78e-07 $l=6.95e-07 $layer=LI1_cond $X=1.235 $Y=2.12
+ $X2=1.235 $Y2=2.815
r102 16 30 2.56749 $w=3.75e-07 $l=2.43824e-07 $layer=LI1_cond $X=1.03 $Y=1.95
+ $X2=1.235 $Y2=2.035
r103 15 21 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.03 $Y=1.04
+ $X2=1.115 $Y2=0.875
r104 15 16 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=1.03 $Y=1.04
+ $X2=1.03 $Y2=1.95
r105 13 39 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=3.255 $Y=2.4
+ $X2=3.255 $Y2=1.65
r106 9 38 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=3.16 $Y=0.805
+ $X2=3.16 $Y2=1.32
r107 2 30 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=1.225
+ $Y=1.96 $X2=1.36 $Y2=2.115
r108 2 19 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.225
+ $Y=1.96 $X2=1.36 $Y2=2.815
r109 1 23 91 $w=1.7e-07 $l=6.17475e-07 $layer=licon1_NDIFF $count=2 $X=0.97
+ $Y=0.625 $X2=1.475 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_MS__XOR2_1%VPWR 1 2 9 15 18 19 20 26 35 36 39
r42 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 36 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r45 33 39 10.4332 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=2.695 $Y=3.33
+ $X2=2.475 $Y2=3.33
r46 33 35 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=2.695 $Y=3.33
+ $X2=3.6 $Y2=3.33
r47 32 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 28 31 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 26 39 10.4332 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=2.255 $Y=3.33
+ $X2=2.475 $Y2=3.33
r52 26 31 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.255 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 24 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r55 20 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r56 20 29 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 18 23 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.325 $Y=3.33
+ $X2=0.24 $Y2=3.33
r58 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.325 $Y=3.33
+ $X2=0.49 $Y2=3.33
r59 17 28 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=0.655 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.655 $Y=3.33
+ $X2=0.49 $Y2=3.33
r61 13 39 1.73497 $w=4.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=3.245
+ $X2=2.475 $Y2=3.33
r62 13 15 11.2625 $w=4.38e-07 $l=4.3e-07 $layer=LI1_cond $X=2.475 $Y=3.245
+ $X2=2.475 $Y2=2.815
r63 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.49 $Y=2.105 $X2=0.49
+ $Y2=2.815
r64 7 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.49 $Y=3.245 $X2=0.49
+ $Y2=3.33
r65 7 12 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.49 $Y=3.245
+ $X2=0.49 $Y2=2.815
r66 2 15 600 $w=1.7e-07 $l=1.07034e-06 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=1.84 $X2=2.475 $Y2=2.815
r67 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.345
+ $Y=1.96 $X2=0.49 $Y2=2.815
r68 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.345
+ $Y=1.96 $X2=0.49 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_MS__XOR2_1%A_355_368# 1 2 9 14 16
c23 16 0 3.44191e-19 $X=3.03 $Y=2.455
r24 10 14 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.085 $Y=2.375
+ $X2=1.92 $Y2=2.375
r25 9 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.865 $Y=2.375
+ $X2=3.03 $Y2=2.375
r26 9 10 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=2.865 $Y=2.375
+ $X2=2.085 $Y2=2.375
r27 2 16 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=2.845
+ $Y=1.84 $X2=3.03 $Y2=2.455
r28 1 14 300 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_PDIFF $count=2 $X=1.775
+ $Y=1.84 $X2=1.92 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_MS__XOR2_1%X 1 2 7 11 16 17 18 19 23 31
r36 23 31 1.42437 $w=4.43e-07 $l=5.5e-08 $layer=LI1_cond $X=2.747 $Y=0.98
+ $X2=2.747 $Y2=0.925
r37 19 23 2.41799 $w=4.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.747 $Y=1.065
+ $X2=2.747 $Y2=0.98
r38 19 31 0.388464 $w=4.43e-07 $l=1.5e-08 $layer=LI1_cond $X=2.747 $Y=0.91
+ $X2=2.747 $Y2=0.925
r39 19 28 8.54621 $w=4.43e-07 $l=3.3e-07 $layer=LI1_cond $X=2.747 $Y=0.91
+ $X2=2.747 $Y2=0.58
r40 18 28 0.64744 $w=4.43e-07 $l=2.5e-08 $layer=LI1_cond $X=2.747 $Y=0.555
+ $X2=2.747 $Y2=0.58
r41 16 17 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=3.56 $Y=1.985
+ $X2=3.56 $Y2=1.82
r42 13 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.67 $Y=1.15
+ $X2=3.67 $Y2=1.82
r43 9 16 0.886495 $w=3.88e-07 $l=3e-08 $layer=LI1_cond $X=3.56 $Y=2.015 $X2=3.56
+ $Y2=1.985
r44 9 11 23.6399 $w=3.88e-07 $l=8e-07 $layer=LI1_cond $X=3.56 $Y=2.015 $X2=3.56
+ $Y2=2.815
r45 8 19 6.34366 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=2.97 $Y=1.065
+ $X2=2.747 $Y2=1.065
r46 7 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.585 $Y=1.065
+ $X2=3.67 $Y2=1.15
r47 7 8 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=3.585 $Y=1.065
+ $X2=2.97 $Y2=1.065
r48 2 16 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=3.345
+ $Y=1.84 $X2=3.53 $Y2=1.985
r49 2 11 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=3.345
+ $Y=1.84 $X2=3.53 $Y2=2.815
r50 1 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.665
+ $Y=0.435 $X2=2.805 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__XOR2_1%VGND 1 2 3 10 12 16 22 25 26 27 28 29 30 44
r42 47 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r43 46 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r44 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r45 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r46 41 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r47 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r48 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r49 37 40 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r50 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r51 35 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r52 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r53 32 46 6.94742 $w=1.7e-07 $l=3.88e-07 $layer=LI1_cond $X=0.775 $Y=0 $X2=0.387
+ $Y2=0
r54 32 34 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=0.775 $Y=0 $X2=1.68
+ $Y2=0
r55 30 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r56 30 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r57 28 40 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.21 $Y=0 $X2=3.12
+ $Y2=0
r58 28 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.21 $Y=0 $X2=3.375
+ $Y2=0
r59 27 43 4.30588 $w=1.7e-07 $l=6e-08 $layer=LI1_cond $X=3.54 $Y=0 $X2=3.6 $Y2=0
r60 27 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.54 $Y=0 $X2=3.375
+ $Y2=0
r61 25 34 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.82 $Y=0 $X2=1.68
+ $Y2=0
r62 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.82 $Y=0 $X2=1.985
+ $Y2=0
r63 24 37 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=2.15 $Y=0 $X2=2.16
+ $Y2=0
r64 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.15 $Y=0 $X2=1.985
+ $Y2=0
r65 20 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.375 $Y=0.085
+ $X2=3.375 $Y2=0
r66 20 22 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=3.375 $Y=0.085
+ $X2=3.375 $Y2=0.58
r67 16 18 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.985 $Y=0.58
+ $X2=1.985 $Y2=1.03
r68 14 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.985 $Y=0.085
+ $X2=1.985 $Y2=0
r69 14 16 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=1.985 $Y=0.085
+ $X2=1.985 $Y2=0.58
r70 10 46 3.09769 $w=6e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.475 $Y=0.085
+ $X2=0.387 $Y2=0
r71 10 12 14.7516 $w=5.98e-07 $l=7.4e-07 $layer=LI1_cond $X=0.475 $Y=0.085
+ $X2=0.475 $Y2=0.825
r72 3 22 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.235
+ $Y=0.435 $X2=3.375 $Y2=0.58
r73 2 18 182 $w=1.7e-07 $l=5.03115e-07 $layer=licon1_NDIFF $count=1 $X=1.765
+ $Y=0.625 $X2=1.985 $Y2=1.03
r74 2 16 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=1.765
+ $Y=0.625 $X2=1.985 $Y2=0.58
r75 1 12 91 $w=1.7e-07 $l=5.5608e-07 $layer=licon1_NDIFF $count=2 $X=0.215
+ $Y=0.625 $X2=0.68 $Y2=0.825
.ends


# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__nor4_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__nor4_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.640000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.028400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.045000 1.300000 8.515000 1.630000 ;
        RECT 7.805000 1.180000 8.515000 1.300000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.028400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.350000 6.595000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.028400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.435000 1.350000 3.785000 1.780000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  1.028400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.350000 1.875000 1.780000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  3.147200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.010000 7.570000 1.130000 ;
        RECT 0.125000 1.130000 4.590000 1.180000 ;
        RECT 0.125000 1.180000 0.355000 1.950000 ;
        RECT 0.125000 1.950000 1.895000 2.120000 ;
        RECT 0.615000 0.350000 1.740000 1.010000 ;
        RECT 0.615000 2.120000 0.945000 2.735000 ;
        RECT 1.565000 2.120000 1.895000 2.735000 ;
        RECT 2.410000 0.350000 3.590000 1.010000 ;
        RECT 4.260000 0.350000 4.590000 0.960000 ;
        RECT 4.260000 0.960000 7.860000 1.010000 ;
        RECT 7.240000 0.340000 7.860000 0.960000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.640000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.640000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.640000 0.085000 ;
      RECT 0.000000  3.245000 8.640000 3.415000 ;
      RECT 0.115000  0.085000 0.445000 0.840000 ;
      RECT 0.115000  2.290000 0.445000 2.905000 ;
      RECT 0.115000  2.905000 2.265000 3.075000 ;
      RECT 1.145000  2.290000 1.395000 2.905000 ;
      RECT 1.910000  0.085000 2.240000 0.840000 ;
      RECT 2.095000  1.820000 2.265000 1.950000 ;
      RECT 2.095000  1.950000 4.145000 2.120000 ;
      RECT 2.095000  2.120000 2.265000 2.905000 ;
      RECT 2.465000  2.290000 2.795000 2.905000 ;
      RECT 2.465000  2.905000 6.075000 3.075000 ;
      RECT 2.970000  2.120000 3.190000 2.735000 ;
      RECT 3.365000  2.290000 3.695000 2.905000 ;
      RECT 3.760000  0.085000 4.090000 0.840000 ;
      RECT 3.895000  2.120000 4.145000 2.735000 ;
      RECT 4.375000  1.950000 8.525000 2.120000 ;
      RECT 4.375000  2.120000 4.625000 2.735000 ;
      RECT 4.760000  0.085000 7.070000 0.790000 ;
      RECT 4.825000  2.300000 5.155000 2.905000 ;
      RECT 5.340000  2.120000 5.560000 2.735000 ;
      RECT 5.745000  2.300000 6.075000 2.905000 ;
      RECT 6.255000  2.120000 6.525000 2.980000 ;
      RECT 6.695000  2.290000 7.025000 3.245000 ;
      RECT 7.195000  2.120000 7.525000 2.980000 ;
      RECT 7.695000  2.290000 8.025000 3.245000 ;
      RECT 8.030000  0.085000 8.360000 1.010000 ;
      RECT 8.195000  1.820000 8.525000 1.950000 ;
      RECT 8.195000  2.120000 8.525000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
  END
END sky130_fd_sc_ms__nor4_4

* File: sky130_fd_sc_ms__o21bai_2.spice
* Created: Fri Aug 28 17:56:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o21bai_2.pex.spice"
.subckt sky130_fd_sc_ms__o21bai_2  VNB VPB B1_N A1 A2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2	A2
* A1	A1
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_B1_N_M1011_g N_A_27_74#_M1011_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.1824 PD=1.85 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_A_225_74#_M1007_d N_A_27_74#_M1007_g N_Y_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.5 A=0.111 P=1.78 MULT=1
MM1013 N_A_225_74#_M1013_d N_A_27_74#_M1013_g N_Y_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1004 N_A_225_74#_M1013_d N_A1_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1406 PD=1.09 PS=1.12 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1005 N_A_225_74#_M1005_d N_A2_M1005_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1406 PD=1.02 PS=1.12 NRD=0 NRS=4.86 M=1 R=4.93333 SA=75001.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1010 N_A_225_74#_M1005_d N_A2_M1010_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1006 N_A_225_74#_M1006_d N_A1_M1006_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1000 N_VPWR_M1000_d N_B1_N_M1000_g N_A_27_74#_M1000_s VPB PSHORT L=0.18 W=1
+ AD=0.302358 AS=0.29 PD=1.61321 PS=2.58 NRD=47.5952 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90003.3 A=0.18 P=2.36 MULT=1
MM1008 N_Y_M1008_d N_A_27_74#_M1008_g N_VPWR_M1000_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.338642 PD=1.39 PS=1.80679 NRD=0 NRS=12.2928 M=1 R=6.22222
+ SA=90000.9 SB=90002.5 A=0.2016 P=2.6 MULT=1
MM1009 N_Y_M1008_d N_A_27_74#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2016 PD=1.39 PS=1.48 NRD=0 NRS=2.6201 M=1 R=6.22222 SA=90001.4
+ SB=90002.1 A=0.2016 P=2.6 MULT=1
MM1001 N_A_510_368#_M1001_d N_A1_M1001_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2016 PD=1.39 PS=1.48 NRD=0 NRS=11.426 M=1 R=6.22222 SA=90001.9
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1002 N_Y_M1002_d N_A2_M1002_g N_A_510_368#_M1001_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.3
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1003 N_Y_M1002_d N_A2_M1003_g N_A_510_368#_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.154 PD=1.39 PS=1.395 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.8
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1012 N_A_510_368#_M1003_s N_A1_M1012_g N_VPWR_M1012_s VPB PSHORT L=0.18 W=1.12
+ AD=0.154 AS=0.3136 PD=1.395 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.742 P=13.12
*
.include "sky130_fd_sc_ms__o21bai_2.pxi.spice"
*
.ends
*
*

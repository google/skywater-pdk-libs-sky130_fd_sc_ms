* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__fa_2 A B CIN VGND VNB VPB VPWR COUT SUM
X0 a_487_347# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X1 a_27_79# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 VGND CIN a_701_79# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 a_1097_347# B a_1205_368# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X4 VGND A a_701_79# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 a_686_347# B VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X6 SUM a_995_347# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X7 VGND a_339_347# COUT VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X8 a_27_378# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X9 a_701_79# a_339_347# a_995_347# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X10 a_995_347# CIN a_1097_347# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X11 VPWR B a_27_378# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X12 VGND B a_27_79# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X13 a_686_347# a_339_347# a_995_347# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X14 VPWR CIN a_686_347# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X15 COUT a_339_347# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X16 VGND a_995_347# SUM VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X17 a_995_347# CIN a_1119_79# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 a_487_79# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X19 a_339_347# B a_487_79# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X20 VPWR a_995_347# SUM VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X21 a_1205_79# A VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 a_1205_368# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X23 a_1119_79# B a_1205_79# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X24 SUM a_995_347# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X25 VPWR a_339_347# COUT VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X26 a_27_79# CIN a_339_347# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X27 a_339_347# B a_487_347# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X28 VPWR A a_686_347# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X29 a_27_378# CIN a_339_347# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X30 COUT a_339_347# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X31 a_701_79# B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

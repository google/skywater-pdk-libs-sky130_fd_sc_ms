* NGSPICE file created from sky130_fd_sc_ms__a2bb2oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 Y B2 a_615_74# VNB nlowvt w=740000u l=150000u
+  ad=4.144e+11p pd=4.08e+06u as=5.994e+11p ps=6.06e+06u
M1001 a_212_392# A1_N VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.1e+11p pd=2.42e+06u as=8.648e+11p ps=8.08e+06u
M1002 Y a_212_102# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=8.17e+11p ps=8.02e+06u
M1003 Y a_212_102# a_424_368# VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=1.1872e+12p ps=1.108e+07u
M1004 a_424_368# a_212_102# Y VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_615_74# B1 VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_615_74# B2 Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2_N a_212_102# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.93e+06u
M1008 VPWR B2 a_424_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_424_368# B2 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR B1 a_424_368# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_212_102# A1_N VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_212_102# Y VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_424_368# B1 VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND B1 a_615_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_212_102# A2_N a_212_392# VPB pshort w=1e+06u l=180000u
+  ad=2.6e+11p pd=2.52e+06u as=0p ps=0u
.ends


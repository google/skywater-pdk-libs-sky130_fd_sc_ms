* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfrtp_4 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 a_834_93# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_225_81# a_27_74# a_312_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X2 a_225_81# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X3 a_1367_112# a_1037_387# a_1745_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 Q a_2339_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 VPWR a_1745_74# a_2339_74# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X6 a_1955_74# a_2003_48# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X7 Q a_2339_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X8 a_343_464# D a_415_81# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X9 a_517_464# SCD VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X10 a_2003_48# a_1745_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X11 VGND RESET_B a_2141_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X12 a_834_93# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X13 a_2141_74# a_1745_74# a_2003_48# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X14 VPWR RESET_B a_2003_48# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X15 VPWR a_834_93# a_1037_387# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X16 a_27_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X17 a_1745_74# a_1037_387# a_1985_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X18 a_1233_138# a_1037_387# a_1319_138# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X19 VPWR a_1233_138# a_1367_112# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X20 a_312_81# D a_415_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X21 a_2339_74# a_1745_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X22 VGND a_2339_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X23 a_1345_463# a_1367_112# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X24 VPWR a_2339_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X25 a_415_81# a_1037_387# a_1233_138# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X26 a_1397_138# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X27 VPWR RESET_B a_1233_138# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X28 VPWR a_2339_74# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X29 Q a_2339_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X30 a_2339_74# a_1745_74# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X31 a_1745_74# a_834_93# a_1955_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X32 a_415_81# a_27_74# a_517_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X33 Q a_2339_74# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X34 a_415_81# SCE a_555_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X35 VGND a_2339_74# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X36 a_1233_138# a_834_93# a_1345_463# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X37 VGND a_834_93# a_1037_387# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X38 a_555_81# SCD a_225_81# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X39 VPWR RESET_B a_415_81# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X40 a_1985_508# a_2003_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X41 a_415_81# a_834_93# a_1233_138# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X42 a_1367_112# a_834_93# a_1745_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X43 VPWR SCE a_343_464# VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X44 a_27_74# SCE VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X45 a_1319_138# a_1367_112# a_1397_138# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X46 VGND a_1233_138# a_1367_112# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
.ends

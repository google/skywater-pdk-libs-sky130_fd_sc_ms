* File: sky130_fd_sc_ms__a222o_2.spice
* Created: Wed Sep  2 11:52:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a222o_2.pex.spice"
.subckt sky130_fd_sc_ms__a222o_2  VNB VPB C1 C2 A1 B1 B2 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* B2	B2
* B1	B1
* A1	A1
* C2	C2
* C1	C1
* VPB	VPB
* VNB	VNB
MM1004 A_114_82# N_C1_M1004_g N_A_27_82#_M1004_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1824 PD=0.88 PS=1.85 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.8 A=0.096 P=1.58 MULT=1
MM1015 N_VGND_M1015_d N_C2_M1015_g A_114_82# VNB NLOWVT L=0.15 W=0.64
+ AD=0.192649 AS=0.0768 PD=1.25217 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667
+ SA=75000.6 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1005 N_X_M1005_d N_A_27_82#_M1005_g N_VGND_M1015_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.222751 PD=1.02 PS=1.44783 NRD=0 NRS=53.508 M=1 R=4.93333
+ SA=75001.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1010 N_X_M1005_d N_A_27_82#_M1010_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2586 PD=1.02 PS=2.67 NRD=0 NRS=47.748 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_A_27_82#_M1007_d N_A1_M1007_g N_A_557_74#_M1007_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1504 AS=0.1971 PD=1.11 PS=1.92 NRD=20.616 NRS=6.552 M=1 R=4.26667
+ SA=75000.2 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1011 A_775_74# N_B1_M1011_g N_A_27_82#_M1007_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1504 PD=0.88 PS=1.11 NRD=12.18 NRS=14.988 M=1 R=4.26667
+ SA=75000.9 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1012 N_VGND_M1012_d N_B2_M1012_g A_775_74# VNB NLOWVT L=0.15 W=0.64 AD=0.1344
+ AS=0.0768 PD=1.06 PS=0.88 NRD=3.744 NRS=12.18 M=1 R=4.26667 SA=75001.2
+ SB=75000.8 A=0.096 P=1.58 MULT=1
MM1000 N_A_557_74#_M1000_d N_A2_M1000_g N_VGND_M1012_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.1344 PD=1.85 PS=1.06 NRD=0 NRS=22.488 M=1 R=4.26667 SA=75001.8
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_A_119_392#_M1001_d N_C1_M1001_g N_A_27_82#_M1001_s VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.28 PD=1.27 PS=2.56 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1002 N_A_27_82#_M1002_d N_C2_M1002_g N_A_119_392#_M1001_d VPB PSHORT L=0.18
+ W=1 AD=0.28 AS=0.135 PD=2.56 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90000.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1006 N_X_M1006_d N_A_27_82#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.32385 PD=1.39 PS=3.09 NRD=0 NRS=14.9326 M=1 R=6.22222
+ SA=90000.2 SB=90002.7 A=0.2016 P=2.6 MULT=1
MM1008 N_X_M1006_d N_A_27_82#_M1008_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.264785 PD=1.39 PS=1.7117 NRD=0 NRS=14.9326 M=1 R=6.22222
+ SA=90000.6 SB=90002.2 A=0.2016 P=2.6 MULT=1
MM1003 N_A_642_368#_M1003_d N_A1_M1003_g N_VPWR_M1008_s VPB PSHORT L=0.18 W=1
+ AD=0.26675 AS=0.236415 PD=1.655 PS=1.5283 NRD=19.6803 NRS=16.7253 M=1
+ R=5.55556 SA=90001.2 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1013 N_A_119_392#_M1013_d N_B1_M1013_g N_A_642_368#_M1003_d VPB PSHORT L=0.18
+ W=1 AD=0.135 AS=0.26675 PD=1.27 PS=1.655 NRD=0 NRS=41.7049 M=1 R=5.55556
+ SA=90001.9 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1014 N_A_642_368#_M1014_d N_B2_M1014_g N_A_119_392#_M1013_d VPB PSHORT L=0.18
+ W=1 AD=0.185 AS=0.135 PD=1.37 PS=1.27 NRD=8.8453 NRS=0 M=1 R=5.55556
+ SA=90002.3 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_A2_M1009_g N_A_642_368#_M1014_d VPB PSHORT L=0.18 W=1
+ AD=0.28 AS=0.185 PD=2.56 PS=1.37 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90002.9
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX16_noxref VNB VPB NWDIODE A=10.5276 P=15.04
c_675 A_775_74# 0 2.49076e-20 $X=3.875 $Y=0.37
*
.include "sky130_fd_sc_ms__a222o_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__dfbbp_1.spice
* Created: Wed Sep  2 12:02:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dfbbp_1.pex.spice"
.subckt sky130_fd_sc_ms__dfbbp_1  VNB VPB CLK D SET_B RESET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1029 N_VGND_M1029_d N_CLK_M1029_g N_A_27_74#_M1029_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.2109 PD=1.09 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1017 N_A_214_74#_M1017_d N_A_27_74#_M1017_g N_VGND_M1029_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1032 N_A_422_125#_M1032_d N_D_M1032_g N_VGND_M1032_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.088025 AS=0.1197 PD=0.95 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1004 N_A_520_87#_M1004_d N_A_27_74#_M1004_g N_A_422_125#_M1032_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.088025 PD=0.7 PS=0.95 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75000.5 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1025 A_606_87# N_A_214_74#_M1025_g N_A_520_87#_M1004_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.08225 AS=0.0588 PD=0.905 PS=0.7 NRD=40.236 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1036 N_VGND_M1036_d N_A_671_93#_M1036_g A_606_87# VNB NLOWVT L=0.15 W=0.42
+ AD=0.205962 AS=0.08225 PD=1.31629 PS=0.905 NRD=124.392 NRS=40.236 M=1 R=2.8
+ SA=75001 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1033 N_A_872_119#_M1033_d N_SET_B_M1033_g N_VGND_M1036_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.192025 AS=0.269713 PD=1.335 PS=1.72371 NRD=64.164 NRS=94.992 M=1
+ R=3.66667 SA=75001.5 SB=75001.4 A=0.0825 P=1.4 MULT=1
MM1022 N_A_671_93#_M1022_d N_A_520_87#_M1022_g N_A_872_119#_M1033_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.192025 PD=0.83 PS=1.335 NRD=0 NRS=64.164 M=1
+ R=3.66667 SA=75002.1 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1030 N_A_872_119#_M1030_d N_A_1062_93#_M1030_g N_A_671_93#_M1022_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.26245 AS=0.077 PD=2.29 PS=0.83 NRD=92.112 NRS=0 M=1
+ R=3.66667 SA=75002.6 SB=75000.3 A=0.0825 P=1.4 MULT=1
MM1006 A_1318_119# N_A_671_93#_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.05775 AS=0.26105 PD=0.76 PS=2.28 NRD=10.908 NRS=0 M=1 R=3.66667
+ SA=75000.3 SB=75001.5 A=0.0825 P=1.4 MULT=1
MM1012 N_A_1314_424#_M1012_d N_A_214_74#_M1012_g A_1318_119# VNB NLOWVT L=0.15
+ W=0.55 AD=0.131376 AS=0.05775 PD=1.32113 PS=0.76 NRD=0 NRS=10.908 M=1
+ R=3.66667 SA=75000.6 SB=75001.1 A=0.0825 P=1.4 MULT=1
MM1014 A_1498_74# N_A_27_74#_M1014_g N_A_1314_424#_M1012_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0819 AS=0.100324 PD=0.81 PS=1.00887 NRD=39.996 NRS=32.856 M=1
+ R=2.8 SA=75000.6 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_A_1474_446#_M1021_g A_1498_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0877655 AS=0.0819 PD=0.796552 PS=0.81 NRD=22.848 NRS=39.996 M=1 R=2.8
+ SA=75001.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1034 N_A_1708_74#_M1034_d N_SET_B_M1034_g N_VGND_M1021_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1295 AS=0.154634 PD=1.09 PS=1.40345 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1027 N_A_1474_446#_M1027_d N_A_1314_424#_M1027_g N_A_1708_74#_M1034_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.10545 AS=0.1295 PD=1.025 PS=1.09 NRD=0.804 NRS=0 M=1
+ R=4.93333 SA=75001.6 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1031 N_A_1708_74#_M1031_d N_A_1062_93#_M1031_g N_A_1474_446#_M1027_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.2294 AS=0.10545 PD=2.1 PS=1.025 NRD=4.044 NRS=0 M=1
+ R=4.93333 SA=75002 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1007_d N_RESET_B_M1007_g N_A_1062_93#_M1007_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.0943552 AS=0.1197 PD=0.847241 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1002 N_Q_N_M1002_d N_A_1474_446#_M1002_g N_VGND_M1007_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.166245 PD=2.05 PS=1.49276 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1019 N_VGND_M1019_d N_A_1474_446#_M1019_g N_A_2320_410#_M1019_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0783879 AS=0.1197 PD=0.771207 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1038 N_Q_M1038_d N_A_2320_410#_M1038_g N_VGND_M1019_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1998 AS=0.138112 PD=2.02 PS=1.35879 NRD=0 NRS=7.296 M=1 R=4.93333
+ SA=75000.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1018 N_VPWR_M1018_d N_CLK_M1018_g N_A_27_74#_M1018_s VPB PSHORT L=0.18 W=1.12
+ AD=0.224 AS=0.3136 PD=1.52 PS=2.8 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.8 A=0.2016 P=2.6 MULT=1
MM1028 N_A_214_74#_M1028_d N_A_27_74#_M1028_g N_VPWR_M1018_d VPB PSHORT L=0.18
+ W=1.12 AD=0.2912 AS=0.224 PD=2.76 PS=1.52 NRD=0 NRS=13.1793 M=1 R=6.22222
+ SA=90000.8 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1013 N_A_422_125#_M1013_d N_D_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.18 W=0.42
+ AD=0.0567 AS=0.2541 PD=0.69 PS=2.05 NRD=0 NRS=0 M=1 R=2.33333 SA=90000.5
+ SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1016 N_A_520_87#_M1016_d N_A_214_74#_M1016_g N_A_422_125#_M1013_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.10815 AS=0.0567 PD=1.18 PS=0.69 NRD=94.9737 NRS=0 M=1
+ R=2.33333 SA=90001 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1039 A_716_379# N_A_27_74#_M1039_g N_A_520_87#_M1016_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0441 AS=0.10815 PD=0.63 PS=1.18 NRD=23.443 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90002.9 A=0.0756 P=1.2 MULT=1
MM1009 N_VPWR_M1009_d N_A_671_93#_M1009_g A_716_379# VPB PSHORT L=0.18 W=0.42
+ AD=0.0924 AS=0.0441 PD=0.833333 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.33333
+ SA=90000.6 SB=90002.5 A=0.0756 P=1.2 MULT=1
MM1020 N_A_671_93#_M1020_d N_SET_B_M1020_g N_VPWR_M1009_d VPB PSHORT L=0.18
+ W=0.84 AD=0.1512 AS=0.1848 PD=1.2 PS=1.66667 NRD=19.9167 NRS=31.6579 M=1
+ R=4.66667 SA=90000.7 SB=90002.7 A=0.1512 P=2.04 MULT=1
MM1035 A_1020_379# N_A_520_87#_M1035_g N_A_671_93#_M1020_d VPB PSHORT L=0.18
+ W=0.84 AD=0.1008 AS=0.1512 PD=1.08 PS=1.2 NRD=15.2281 NRS=0 M=1 R=4.66667
+ SA=90001.2 SB=90002.2 A=0.1512 P=2.04 MULT=1
MM1011 N_VPWR_M1011_d N_A_1062_93#_M1011_g A_1020_379# VPB PSHORT L=0.18 W=0.84
+ AD=0.1386 AS=0.1008 PD=1.17 PS=1.08 NRD=5.8509 NRS=15.2281 M=1 R=4.66667
+ SA=90001.6 SB=90001.8 A=0.1512 P=2.04 MULT=1
MM1003 A_1206_379# N_A_671_93#_M1003_g N_VPWR_M1011_d VPB PSHORT L=0.18 W=0.84
+ AD=0.16695 AS=0.1386 PD=1.425 PS=1.17 NRD=33.7067 NRS=5.8509 M=1 R=4.66667
+ SA=90002.1 SB=90001.3 A=0.1512 P=2.04 MULT=1
MM1005 N_A_1314_424#_M1005_d N_A_27_74#_M1005_g A_1206_379# VPB PSHORT L=0.18
+ W=0.84 AD=0.1778 AS=0.16695 PD=1.59333 PS=1.425 NRD=0 NRS=33.7067 M=1
+ R=4.66667 SA=90001.9 SB=90001.7 A=0.1512 P=2.04 MULT=1
MM1001 A_1421_508# N_A_214_74#_M1001_g N_A_1314_424#_M1005_d VPB PSHORT L=0.18
+ W=0.42 AD=0.05565 AS=0.0889 PD=0.685 PS=0.796667 NRD=36.3465 NRS=37.5088 M=1
+ R=2.33333 SA=90001.6 SB=90002.6 A=0.0756 P=1.2 MULT=1
MM1015 N_VPWR_M1015_d N_A_1474_446#_M1015_g A_1421_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.147237 AS=0.05565 PD=1.08845 PS=0.685 NRD=16.4101 NRS=36.3465 M=1
+ R=2.33333 SA=90002.1 SB=90002.1 A=0.0756 P=1.2 MULT=1
MM1023 N_A_1474_446#_M1023_d N_SET_B_M1023_g N_VPWR_M1015_d VPB PSHORT L=0.18
+ W=1 AD=0.1675 AS=0.350563 PD=1.335 PS=2.59155 NRD=11.8003 NRS=0 M=1 R=5.55556
+ SA=90001.4 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1010 A_1817_392# N_A_1314_424#_M1010_g N_A_1474_446#_M1023_d VPB PSHORT L=0.18
+ W=1 AD=0.1175 AS=0.1675 PD=1.235 PS=1.335 NRD=12.2928 NRS=0 M=1 R=5.55556
+ SA=90001.9 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1024 N_VPWR_M1024_d N_A_1062_93#_M1024_g A_1817_392# VPB PSHORT L=0.18 W=1
+ AD=0.28 AS=0.1175 PD=2.56 PS=1.235 NRD=0 NRS=12.2928 M=1 R=5.55556 SA=90002.3
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_RESET_B_M1000_g N_A_1062_93#_M1000_s VPB PSHORT L=0.18
+ W=0.64 AD=0.123345 AS=0.1664 PD=1.05818 PS=1.8 NRD=42.3747 NRS=0 M=1 R=3.55556
+ SA=90000.2 SB=90000.7 A=0.1152 P=1.64 MULT=1
MM1008 N_Q_N_M1008_d N_A_1474_446#_M1008_g N_VPWR_M1000_d VPB PSHORT L=0.18
+ W=1.12 AD=0.2912 AS=0.215855 PD=2.76 PS=1.85182 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.5 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1026 N_VPWR_M1026_d N_A_1474_446#_M1026_g N_A_2320_410#_M1026_s VPB PSHORT
+ L=0.18 W=0.84 AD=0.1518 AS=0.2184 PD=1.24714 PS=2.2 NRD=28.7226 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1037 N_Q_M1037_d N_A_2320_410#_M1037_g N_VPWR_M1026_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3024 AS=0.2024 PD=2.78 PS=1.66286 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX40_noxref VNB VPB NWDIODE A=24.8124 P=30.4
c_157 VNB 0 1.25678e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__dfbbp_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__o41ai_4.pex.spice
* Created: Fri Aug 28 18:05:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O41AI_4%B1 3 5 7 8 10 13 15 17 18 19 20 22 23 24 35
c68 15 0 6.95413e-20 $X=1.355 $Y=1.185
c69 8 0 6.95413e-20 $X=0.925 $Y=1.185
r70 34 36 11.4038 $w=3.17e-07 $l=7.5e-08 $layer=POLY_cond $X=0.98 $Y=1.367
+ $X2=1.055 $Y2=1.367
r71 34 35 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.98
+ $Y=1.385 $X2=0.98 $Y2=1.385
r72 32 34 8.36278 $w=3.17e-07 $l=5.5e-08 $layer=POLY_cond $X=0.925 $Y=1.367
+ $X2=0.98 $Y2=1.367
r73 31 32 63.8612 $w=3.17e-07 $l=4.2e-07 $layer=POLY_cond $X=0.505 $Y=1.367
+ $X2=0.925 $Y2=1.367
r74 30 31 1.5205 $w=3.17e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.367
+ $X2=0.505 $Y2=1.367
r75 28 30 29.6498 $w=3.17e-07 $l=1.95e-07 $layer=POLY_cond $X=0.3 $Y=1.367
+ $X2=0.495 $Y2=1.367
r76 28 29 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.3
+ $Y=1.385 $X2=0.3 $Y2=1.385
r77 24 35 8.09825 $w=3.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=0.98 $Y2=1.365
r78 24 29 13.0818 $w=3.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.72 $Y=1.365
+ $X2=0.3 $Y2=1.365
r79 23 29 1.86883 $w=3.68e-07 $l=6e-08 $layer=LI1_cond $X=0.24 $Y=1.365 $X2=0.3
+ $Y2=1.365
r80 20 22 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.855 $Y=1.185
+ $X2=1.855 $Y2=0.74
r81 18 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.78 $Y=1.26
+ $X2=1.855 $Y2=1.185
r82 18 19 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.78 $Y=1.26
+ $X2=1.43 $Y2=1.26
r83 15 19 24.856 $w=3.17e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.355 $Y=1.185
+ $X2=1.43 $Y2=1.26
r84 15 36 45.6151 $w=3.17e-07 $l=3.80263e-07 $layer=POLY_cond $X=1.355 $Y=1.185
+ $X2=1.055 $Y2=1.367
r85 15 17 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.355 $Y=1.185
+ $X2=1.355 $Y2=0.74
r86 11 36 15.9969 $w=1.8e-07 $l=1.83e-07 $layer=POLY_cond $X=1.055 $Y=1.55
+ $X2=1.055 $Y2=1.367
r87 11 13 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=1.055 $Y=1.55
+ $X2=1.055 $Y2=2.4
r88 8 32 20.269 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=0.925 $Y=1.185
+ $X2=0.925 $Y2=1.367
r89 8 10 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.925 $Y=1.185
+ $X2=0.925 $Y2=0.74
r90 5 30 20.269 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=0.495 $Y=1.185
+ $X2=0.495 $Y2=1.367
r91 5 7 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=0.495 $Y=1.185
+ $X2=0.495 $Y2=0.74
r92 1 31 15.9969 $w=1.8e-07 $l=1.83e-07 $layer=POLY_cond $X=0.505 $Y=1.55
+ $X2=0.505 $Y2=1.367
r93 1 3 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=0.505 $Y=1.55
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O41AI_4%A4 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 23
+ 24 26 27 28 40
c104 24 0 3.37137e-19 $X=3.97 $Y=1.185
c105 23 0 1.72039e-20 $X=3.615 $Y=1.26
c106 22 0 8.21537e-20 $X=3.895 $Y=1.26
c107 19 0 1.95112e-19 $X=3.54 $Y=1.185
c108 4 0 1.05859e-19 $X=2.355 $Y=1.185
r109 41 42 33.6992 $w=4.72e-07 $l=3.3e-07 $layer=POLY_cond $X=3.085 $Y=1.455
+ $X2=3.415 $Y2=1.455
r110 39 41 9.19068 $w=4.72e-07 $l=9e-08 $layer=POLY_cond $X=2.995 $Y=1.455
+ $X2=3.085 $Y2=1.455
r111 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.995
+ $Y=1.385 $X2=2.995 $Y2=1.385
r112 37 39 3.06356 $w=4.72e-07 $l=3e-08 $layer=POLY_cond $X=2.965 $Y=1.455
+ $X2=2.995 $Y2=1.455
r113 36 37 45.9534 $w=4.72e-07 $l=4.5e-07 $layer=POLY_cond $X=2.515 $Y=1.455
+ $X2=2.965 $Y2=1.455
r114 35 36 16.339 $w=4.72e-07 $l=1.6e-07 $layer=POLY_cond $X=2.355 $Y=1.455
+ $X2=2.515 $Y2=1.455
r115 33 35 4.08475 $w=4.72e-07 $l=4e-08 $layer=POLY_cond $X=2.315 $Y=1.455
+ $X2=2.355 $Y2=1.455
r116 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.315
+ $Y=1.385 $X2=2.315 $Y2=1.385
r117 28 40 11.0572 $w=3.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.64 $Y=1.365
+ $X2=2.995 $Y2=1.365
r118 28 34 10.1228 $w=3.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.64 $Y=1.365
+ $X2=2.315 $Y2=1.365
r119 27 34 4.8278 $w=3.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.16 $Y=1.365
+ $X2=2.315 $Y2=1.365
r120 24 26 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.97 $Y=1.185
+ $X2=3.97 $Y2=0.74
r121 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.895 $Y=1.26
+ $X2=3.97 $Y2=1.185
r122 22 23 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.895 $Y=1.26
+ $X2=3.615 $Y2=1.26
r123 19 23 32.0248 $w=4.72e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.54 $Y=1.185
+ $X2=3.615 $Y2=1.26
r124 19 42 12.7648 $w=4.72e-07 $l=3.26573e-07 $layer=POLY_cond $X=3.54 $Y=1.185
+ $X2=3.415 $Y2=1.455
r125 19 21 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.54 $Y=1.185
+ $X2=3.54 $Y2=0.74
r126 16 42 25.4515 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=3.415 $Y=1.725
+ $X2=3.415 $Y2=1.455
r127 16 18 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.415 $Y=1.725
+ $X2=3.415 $Y2=2.4
r128 13 41 29.9582 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.085 $Y=1.185
+ $X2=3.085 $Y2=1.455
r129 13 15 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.085 $Y=1.185
+ $X2=3.085 $Y2=0.74
r130 10 37 25.4515 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=2.965 $Y=1.725
+ $X2=2.965 $Y2=1.455
r131 10 12 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=2.965 $Y=1.725
+ $X2=2.965 $Y2=2.4
r132 7 36 25.4515 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=2.515 $Y=1.725
+ $X2=2.515 $Y2=1.455
r133 7 9 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=2.515 $Y=1.725
+ $X2=2.515 $Y2=2.4
r134 4 35 29.9582 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.355 $Y=1.185
+ $X2=2.355 $Y2=1.455
r135 4 6 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.355 $Y=1.185
+ $X2=2.355 $Y2=0.74
r136 1 33 25.5297 $w=4.72e-07 $l=3.747e-07 $layer=POLY_cond $X=2.065 $Y=1.725
+ $X2=2.315 $Y2=1.455
r137 1 3 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=2.065 $Y=1.725
+ $X2=2.065 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O41AI_4%A3 1 3 4 5 6 8 9 11 12 14 15 17 18 20 21 23
+ 24 26 27 28 29 30 44
c103 30 0 1.39749e-19 $X=6 $Y=1.295
c104 1 0 2.87561e-19 $X=3.865 $Y=1.725
r105 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.58
+ $Y=1.385 $X2=5.58 $Y2=1.385
r106 42 44 27.8935 $w=4.32e-07 $l=2.5e-07 $layer=POLY_cond $X=5.33 $Y=1.472
+ $X2=5.58 $Y2=1.472
r107 41 42 1.67361 $w=4.32e-07 $l=1.5e-08 $layer=POLY_cond $X=5.315 $Y=1.472
+ $X2=5.33 $Y2=1.472
r108 39 41 46.3032 $w=4.32e-07 $l=4.15e-07 $layer=POLY_cond $X=4.9 $Y=1.472
+ $X2=5.315 $Y2=1.472
r109 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.9
+ $Y=1.385 $X2=4.9 $Y2=1.385
r110 37 39 3.90509 $w=4.32e-07 $l=3.5e-08 $layer=POLY_cond $X=4.865 $Y=1.472
+ $X2=4.9 $Y2=1.472
r111 36 37 50.2083 $w=4.32e-07 $l=4.5e-07 $layer=POLY_cond $X=4.415 $Y=1.472
+ $X2=4.865 $Y2=1.472
r112 35 36 1.67361 $w=4.32e-07 $l=1.5e-08 $layer=POLY_cond $X=4.4 $Y=1.472
+ $X2=4.415 $Y2=1.472
r113 30 45 13.0818 $w=3.68e-07 $l=4.2e-07 $layer=LI1_cond $X=6 $Y=1.365 $X2=5.58
+ $Y2=1.365
r114 29 45 1.86883 $w=3.68e-07 $l=6e-08 $layer=LI1_cond $X=5.52 $Y=1.365
+ $X2=5.58 $Y2=1.365
r115 28 29 14.9506 $w=3.68e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.365
+ $X2=5.52 $Y2=1.365
r116 28 40 4.3606 $w=3.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.04 $Y=1.365
+ $X2=4.9 $Y2=1.365
r117 27 40 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.56 $Y=1.365 $X2=4.9
+ $Y2=1.365
r118 24 44 27.8935 $w=4.32e-07 $l=3.55674e-07 $layer=POLY_cond $X=5.83 $Y=1.22
+ $X2=5.58 $Y2=1.472
r119 24 26 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.83 $Y=1.22
+ $X2=5.83 $Y2=0.74
r120 21 42 27.7542 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=5.33 $Y=1.22
+ $X2=5.33 $Y2=1.472
r121 21 23 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.33 $Y=1.22
+ $X2=5.33 $Y2=0.74
r122 18 41 23.3057 $w=1.8e-07 $l=2.53e-07 $layer=POLY_cond $X=5.315 $Y=1.725
+ $X2=5.315 $Y2=1.472
r123 18 20 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=5.315 $Y=1.725
+ $X2=5.315 $Y2=2.4
r124 15 39 27.7542 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=4.9 $Y=1.22
+ $X2=4.9 $Y2=1.472
r125 15 17 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.9 $Y=1.22 $X2=4.9
+ $Y2=0.74
r126 12 37 23.3057 $w=1.8e-07 $l=2.53e-07 $layer=POLY_cond $X=4.865 $Y=1.725
+ $X2=4.865 $Y2=1.472
r127 12 14 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=4.865 $Y=1.725
+ $X2=4.865 $Y2=2.4
r128 9 36 23.3057 $w=1.8e-07 $l=2.53e-07 $layer=POLY_cond $X=4.415 $Y=1.725
+ $X2=4.415 $Y2=1.472
r129 9 11 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=4.415 $Y=1.725
+ $X2=4.415 $Y2=2.4
r130 6 35 27.7542 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=4.4 $Y=1.22 $X2=4.4
+ $Y2=1.472
r131 6 8 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.4 $Y=1.22 $X2=4.4
+ $Y2=0.74
r132 4 35 30.2215 $w=4.32e-07 $l=2.12212e-07 $layer=POLY_cond $X=4.325 $Y=1.65
+ $X2=4.4 $Y2=1.472
r133 4 5 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.325 $Y=1.65
+ $X2=3.955 $Y2=1.65
r134 1 5 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.865 $Y=1.725
+ $X2=3.955 $Y2=1.65
r135 1 3 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.865 $Y=1.725
+ $X2=3.865 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O41AI_4%A2 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 51
c97 27 0 4.367e-20 $X=7.675 $Y=2.4
c98 20 0 9.87313e-20 $X=7.225 $Y=2.4
r99 50 51 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=7.655 $Y=1.385
+ $X2=7.675 $Y2=1.385
r100 48 50 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=7.55 $Y=1.385
+ $X2=7.655 $Y2=1.385
r101 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.55
+ $Y=1.385 $X2=7.55 $Y2=1.385
r102 46 48 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=7.225 $Y=1.385
+ $X2=7.55 $Y2=1.385
r103 45 46 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=7.19 $Y=1.385
+ $X2=7.225 $Y2=1.385
r104 44 45 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=6.775 $Y=1.385
+ $X2=7.19 $Y2=1.385
r105 43 44 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.76 $Y=1.385
+ $X2=6.775 $Y2=1.385
r106 41 43 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=6.53 $Y=1.385
+ $X2=6.76 $Y2=1.385
r107 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.53
+ $Y=1.385 $X2=6.53 $Y2=1.385
r108 39 41 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=6.325 $Y=1.385
+ $X2=6.53 $Y2=1.385
r109 37 39 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=6.26 $Y=1.385
+ $X2=6.325 $Y2=1.385
r110 32 49 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.92 $Y=1.365
+ $X2=7.55 $Y2=1.365
r111 31 49 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=7.44 $Y=1.365
+ $X2=7.55 $Y2=1.365
r112 30 31 14.9506 $w=3.68e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.365
+ $X2=7.44 $Y2=1.365
r113 30 42 13.3933 $w=3.68e-07 $l=4.3e-07 $layer=LI1_cond $X=6.96 $Y=1.365
+ $X2=6.53 $Y2=1.365
r114 29 42 1.55736 $w=3.68e-07 $l=5e-08 $layer=LI1_cond $X=6.48 $Y=1.365
+ $X2=6.53 $Y2=1.365
r115 25 51 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.675 $Y=1.55
+ $X2=7.675 $Y2=1.385
r116 25 27 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=7.675 $Y=1.55
+ $X2=7.675 $Y2=2.4
r117 22 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.22
+ $X2=7.655 $Y2=1.385
r118 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.655 $Y=1.22
+ $X2=7.655 $Y2=0.74
r119 18 46 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.225 $Y=1.55
+ $X2=7.225 $Y2=1.385
r120 18 20 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=7.225 $Y=1.55
+ $X2=7.225 $Y2=2.4
r121 15 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.19 $Y=1.22
+ $X2=7.19 $Y2=1.385
r122 15 17 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.19 $Y=1.22
+ $X2=7.19 $Y2=0.74
r123 11 44 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.775 $Y=1.55
+ $X2=6.775 $Y2=1.385
r124 11 13 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=6.775 $Y=1.55
+ $X2=6.775 $Y2=2.4
r125 8 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.76 $Y=1.22
+ $X2=6.76 $Y2=1.385
r126 8 10 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.76 $Y=1.22 $X2=6.76
+ $Y2=0.74
r127 4 39 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.325 $Y=1.55
+ $X2=6.325 $Y2=1.385
r128 4 6 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=6.325 $Y=1.55
+ $X2=6.325 $Y2=2.4
r129 1 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.26 $Y=1.22
+ $X2=6.26 $Y2=1.385
r130 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.26 $Y=1.22 $X2=6.26
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O41AI_4%A1 3 5 7 10 12 14 17 19 21 22 24 26 28 29 30
+ 31 32
r81 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.47
+ $Y=1.385 $X2=9.47 $Y2=1.385
r82 45 47 55.7267 $w=3.33e-07 $l=3.85e-07 $layer=POLY_cond $X=9.085 $Y=1.43
+ $X2=9.47 $Y2=1.43
r83 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.79
+ $Y=1.385 $X2=8.79 $Y2=1.385
r84 40 42 19.5405 $w=3.33e-07 $l=1.35e-07 $layer=POLY_cond $X=8.655 $Y=1.43
+ $X2=8.79 $Y2=1.43
r85 37 38 2.17117 $w=3.33e-07 $l=1.5e-08 $layer=POLY_cond $X=8.125 $Y=1.43
+ $X2=8.14 $Y2=1.43
r86 32 48 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.84 $Y=1.365
+ $X2=9.47 $Y2=1.365
r87 31 48 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=9.36 $Y=1.365
+ $X2=9.47 $Y2=1.365
r88 30 31 14.9506 $w=3.68e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.365
+ $X2=9.36 $Y2=1.365
r89 30 43 2.80324 $w=3.68e-07 $l=9e-08 $layer=LI1_cond $X=8.88 $Y=1.365 $X2=8.79
+ $Y2=1.365
r90 29 43 12.1474 $w=3.68e-07 $l=3.9e-07 $layer=LI1_cond $X=8.4 $Y=1.365
+ $X2=8.79 $Y2=1.365
r91 26 50 21.4384 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=9.585 $Y=1.22
+ $X2=9.585 $Y2=1.43
r92 26 28 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.585 $Y=1.22
+ $X2=9.585 $Y2=0.74
r93 22 50 1.44745 $w=3.33e-07 $l=1e-08 $layer=POLY_cond $X=9.575 $Y=1.43
+ $X2=9.585 $Y2=1.43
r94 22 47 15.1982 $w=3.33e-07 $l=1.05e-07 $layer=POLY_cond $X=9.575 $Y=1.43
+ $X2=9.47 $Y2=1.43
r95 22 24 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=9.575 $Y=1.55
+ $X2=9.575 $Y2=2.4
r96 19 45 21.4384 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=9.085 $Y=1.22
+ $X2=9.085 $Y2=1.43
r97 19 21 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.085 $Y=1.22
+ $X2=9.085 $Y2=0.74
r98 15 45 1.44745 $w=3.33e-07 $l=1e-08 $layer=POLY_cond $X=9.075 $Y=1.43
+ $X2=9.085 $Y2=1.43
r99 15 42 41.2523 $w=3.33e-07 $l=2.85e-07 $layer=POLY_cond $X=9.075 $Y=1.43
+ $X2=8.79 $Y2=1.43
r100 15 17 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=9.075 $Y=1.55
+ $X2=9.075 $Y2=2.4
r101 12 40 21.4384 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=8.655 $Y=1.22
+ $X2=8.655 $Y2=1.43
r102 12 14 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.655 $Y=1.22
+ $X2=8.655 $Y2=0.74
r103 8 40 4.34234 $w=3.33e-07 $l=3e-08 $layer=POLY_cond $X=8.625 $Y=1.43
+ $X2=8.655 $Y2=1.43
r104 8 38 70.2012 $w=3.33e-07 $l=4.85e-07 $layer=POLY_cond $X=8.625 $Y=1.43
+ $X2=8.14 $Y2=1.43
r105 8 10 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=8.625 $Y=1.55
+ $X2=8.625 $Y2=2.4
r106 5 38 21.4384 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=8.14 $Y=1.22
+ $X2=8.14 $Y2=1.43
r107 5 7 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.14 $Y=1.22 $X2=8.14
+ $Y2=0.74
r108 1 37 17.1428 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=8.125 $Y=1.64
+ $X2=8.125 $Y2=1.43
r109 1 3 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=8.125 $Y=1.64
+ $X2=8.125 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O41AI_4%VPWR 1 2 3 4 13 15 21 25 29 31 33 38 46 53
+ 54 60 63 66
r107 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r108 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r109 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r110 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r111 54 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r112 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r113 51 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.515 $Y=3.33
+ $X2=9.35 $Y2=3.33
r114 51 53 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.515 $Y=3.33
+ $X2=9.84 $Y2=3.33
r115 50 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r116 50 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r117 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r118 47 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.515 $Y=3.33
+ $X2=8.35 $Y2=3.33
r119 47 49 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.515 $Y=3.33
+ $X2=8.88 $Y2=3.33
r120 46 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.185 $Y=3.33
+ $X2=9.35 $Y2=3.33
r121 46 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.185 $Y=3.33
+ $X2=8.88 $Y2=3.33
r122 45 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r123 44 45 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r124 42 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r125 41 44 407.102 $w=1.68e-07 $l=6.24e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=7.92 $Y2=3.33
r126 41 42 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r127 39 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=3.33
+ $X2=1.28 $Y2=3.33
r128 39 41 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.445 $Y=3.33
+ $X2=1.68 $Y2=3.33
r129 38 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.185 $Y=3.33
+ $X2=8.35 $Y2=3.33
r130 38 44 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.185 $Y=3.33
+ $X2=7.92 $Y2=3.33
r131 37 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r132 37 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r133 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r134 34 57 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r135 34 36 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r136 33 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=1.28 $Y2=3.33
r137 33 36 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=0.72 $Y2=3.33
r138 31 45 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=7.92 $Y2=3.33
r139 31 42 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=1.68 $Y2=3.33
r140 27 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.35 $Y=3.245
+ $X2=9.35 $Y2=3.33
r141 27 29 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=9.35 $Y=3.245
+ $X2=9.35 $Y2=2.225
r142 23 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.35 $Y=3.245
+ $X2=8.35 $Y2=3.33
r143 23 25 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=8.35 $Y=3.245
+ $X2=8.35 $Y2=2.225
r144 19 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=3.245
+ $X2=1.28 $Y2=3.33
r145 19 21 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=1.28 $Y=3.245
+ $X2=1.28 $Y2=2.225
r146 15 18 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r147 13 57 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r148 13 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.815
r149 4 29 300 $w=1.7e-07 $l=4.68455e-07 $layer=licon1_PDIFF $count=2 $X=9.165
+ $Y=1.84 $X2=9.35 $Y2=2.225
r150 3 25 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=8.215
+ $Y=1.84 $X2=8.35 $Y2=2.225
r151 2 21 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=1.145
+ $Y=1.84 $X2=1.28 $Y2=2.225
r152 1 18 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r153 1 15 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__O41AI_4%Y 1 2 3 4 5 18 22 24 25 26 27 28 35 41 44 45
+ 46 50
c80 46 0 2.87561e-19 $X=3.12 $Y=2.035
c81 26 0 1.05859e-19 $X=1.64 $Y=1.01
r82 46 50 2.84726 $w=4.3e-07 $l=1.4e-07 $layer=LI1_cond $X=3.19 $Y=1.935
+ $X2=3.05 $Y2=1.935
r83 46 50 0.214408 $w=4.28e-07 $l=8e-09 $layer=LI1_cond $X=3.042 $Y=1.935
+ $X2=3.05 $Y2=1.935
r84 45 46 10.774 $w=4.28e-07 $l=4.02e-07 $layer=LI1_cond $X=2.64 $Y=1.935
+ $X2=3.042 $Y2=1.935
r85 42 45 5.62821 $w=4.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.43 $Y=1.935
+ $X2=2.64 $Y2=1.935
r86 42 44 4.87592 $w=3e-07 $l=1.4e-07 $layer=LI1_cond $X=2.43 $Y=1.935 $X2=2.29
+ $Y2=1.935
r87 35 37 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.71 $Y=0.8
+ $X2=0.71 $Y2=0.925
r88 29 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=1.805
+ $X2=1.64 $Y2=1.805
r89 28 44 4.87592 $w=3e-07 $l=1.94422e-07 $layer=LI1_cond $X=2.15 $Y=1.805
+ $X2=2.29 $Y2=1.935
r90 28 29 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.15 $Y=1.805
+ $X2=1.805 $Y2=1.805
r91 27 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=1.72 $X2=1.64
+ $Y2=1.805
r92 26 40 3.25678 $w=3.3e-07 $l=2.08e-07 $layer=LI1_cond $X=1.64 $Y=1.01
+ $X2=1.64 $Y2=0.802
r93 26 27 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.64 $Y=1.01 $X2=1.64
+ $Y2=1.72
r94 24 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.475 $Y=1.805
+ $X2=1.64 $Y2=1.805
r95 24 25 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.475 $Y=1.805
+ $X2=0.945 $Y2=1.805
r96 23 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=0.925
+ $X2=0.71 $Y2=0.925
r97 22 40 4.50939 $w=1.7e-07 $l=2.17991e-07 $layer=LI1_cond $X=1.475 $Y=0.925
+ $X2=1.64 $Y2=0.802
r98 22 23 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.475 $Y=0.925
+ $X2=0.795 $Y2=0.925
r99 18 20 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.78 $Y=1.985
+ $X2=0.78 $Y2=2.815
r100 16 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.78 $Y=1.89
+ $X2=0.945 $Y2=1.805
r101 16 18 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.78 $Y=1.89
+ $X2=0.78 $Y2=1.985
r102 5 46 300 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=2 $X=3.055
+ $Y=1.84 $X2=3.19 $Y2=1.965
r103 4 44 300 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=2 $X=2.155
+ $Y=1.84 $X2=2.29 $Y2=1.965
r104 3 20 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.78 $Y2=2.815
r105 3 18 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.84 $X2=0.78 $Y2=1.985
r106 2 40 182 $w=1.7e-07 $l=5.85662e-07 $layer=licon1_NDIFF $count=1 $X=1.43
+ $Y=0.37 $X2=1.64 $Y2=0.86
r107 1 35 182 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_MS__O41AI_4%A_339_368# 1 2 3 4 5 18 20 21 24 26 30 34 38
+ 40 44 46 47 48
c94 30 0 2.24545e-20 $X=3.64 $Y=1.965
r95 42 44 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=5.54 $Y=2.905
+ $X2=5.54 $Y2=2.145
r96 41 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.805 $Y=2.99
+ $X2=4.64 $Y2=2.99
r97 40 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.375 $Y=2.99
+ $X2=5.54 $Y2=2.905
r98 40 41 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.375 $Y=2.99
+ $X2=4.805 $Y2=2.99
r99 36 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.64 $Y=2.905
+ $X2=4.64 $Y2=2.99
r100 36 38 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=4.64 $Y=2.905
+ $X2=4.64 $Y2=2.145
r101 35 47 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=3.805 $Y=2.99
+ $X2=3.652 $Y2=2.99
r102 34 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.475 $Y=2.99
+ $X2=4.64 $Y2=2.99
r103 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.475 $Y=2.99
+ $X2=3.805 $Y2=2.99
r104 30 33 32.873 $w=3.03e-07 $l=8.7e-07 $layer=LI1_cond $X=3.652 $Y=1.965
+ $X2=3.652 $Y2=2.835
r105 28 47 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.652 $Y=2.905
+ $X2=3.652 $Y2=2.99
r106 28 33 2.64495 $w=3.03e-07 $l=7e-08 $layer=LI1_cond $X=3.652 $Y=2.905
+ $X2=3.652 $Y2=2.835
r107 27 46 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.88 $Y=2.99 $X2=2.74
+ $Y2=2.99
r108 26 47 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.5 $Y=2.99
+ $X2=3.652 $Y2=2.99
r109 26 27 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.5 $Y=2.99
+ $X2=2.88 $Y2=2.99
r110 22 46 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.74 $Y=2.905
+ $X2=2.74 $Y2=2.99
r111 22 24 17.2866 $w=2.78e-07 $l=4.2e-07 $layer=LI1_cond $X=2.74 $Y=2.905
+ $X2=2.74 $Y2=2.485
r112 20 46 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.6 $Y=2.99 $X2=2.74
+ $Y2=2.99
r113 20 21 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.6 $Y=2.99
+ $X2=1.98 $Y2=2.99
r114 16 21 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=1.827 $Y=2.905
+ $X2=1.98 $Y2=2.99
r115 16 18 25.6938 $w=3.03e-07 $l=6.8e-07 $layer=LI1_cond $X=1.827 $Y=2.905
+ $X2=1.827 $Y2=2.225
r116 5 44 300 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_PDIFF $count=2 $X=5.405
+ $Y=1.84 $X2=5.54 $Y2=2.145
r117 4 38 300 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_PDIFF $count=2 $X=4.505
+ $Y=1.84 $X2=4.64 $Y2=2.145
r118 3 33 400 $w=1.7e-07 $l=1.06035e-06 $layer=licon1_PDIFF $count=1 $X=3.505
+ $Y=1.84 $X2=3.64 $Y2=2.835
r119 3 30 400 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=3.505
+ $Y=1.84 $X2=3.64 $Y2=1.965
r120 2 24 300 $w=1.7e-07 $l=7.09295e-07 $layer=licon1_PDIFF $count=2 $X=2.605
+ $Y=1.84 $X2=2.74 $Y2=2.485
r121 1 18 300 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_PDIFF $count=2 $X=1.695
+ $Y=1.84 $X2=1.84 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_MS__O41AI_4%A_791_368# 1 2 3 4 15 17 18 21 23 27 29 33
+ 35 36
c46 18 0 7.69031e-20 $X=4.305 $Y=1.805
r47 31 33 7.76646 $w=2.28e-07 $l=1.55e-07 $layer=LI1_cond $X=7.45 $Y=1.89
+ $X2=7.45 $Y2=2.045
r48 30 36 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=6.665 $Y=1.805
+ $X2=6.55 $Y2=1.805
r49 29 31 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=7.335 $Y=1.805
+ $X2=7.45 $Y2=1.89
r50 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.335 $Y=1.805
+ $X2=6.665 $Y2=1.805
r51 25 36 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.55 $Y=1.89
+ $X2=6.55 $Y2=1.805
r52 25 27 3.75797 $w=2.28e-07 $l=7.5e-08 $layer=LI1_cond $X=6.55 $Y=1.89
+ $X2=6.55 $Y2=1.965
r53 24 35 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.205 $Y=1.805
+ $X2=5.09 $Y2=1.805
r54 23 36 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=6.435 $Y=1.805
+ $X2=6.55 $Y2=1.805
r55 23 24 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=6.435 $Y=1.805
+ $X2=5.205 $Y2=1.805
r56 19 35 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.09 $Y=1.89
+ $X2=5.09 $Y2=1.805
r57 19 21 3.75797 $w=2.28e-07 $l=7.5e-08 $layer=LI1_cond $X=5.09 $Y=1.89
+ $X2=5.09 $Y2=1.965
r58 17 35 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.975 $Y=1.805
+ $X2=5.09 $Y2=1.805
r59 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.975 $Y=1.805
+ $X2=4.305 $Y2=1.805
r60 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.14 $Y=1.89
+ $X2=4.305 $Y2=1.805
r61 13 15 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=4.14 $Y=1.89
+ $X2=4.14 $Y2=2.045
r62 4 33 300 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_PDIFF $count=2 $X=7.315
+ $Y=1.84 $X2=7.45 $Y2=2.045
r63 3 27 300 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=2 $X=6.415
+ $Y=1.84 $X2=6.55 $Y2=1.965
r64 2 21 300 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=2 $X=4.955
+ $Y=1.84 $X2=5.09 $Y2=1.965
r65 1 15 300 $w=1.7e-07 $l=2.82754e-07 $layer=licon1_PDIFF $count=2 $X=3.955
+ $Y=1.84 $X2=4.14 $Y2=2.045
.ends

.subckt PM_SKY130_FD_SC_MS__O41AI_4%A_1191_368# 1 2 3 4 5 18 20 21 24 26 31 34
+ 35 38 42 46 50 51
c81 50 0 4.367e-20 $X=7 $Y=2.982
c82 35 0 9.87313e-20 $X=8.015 $Y=1.805
r83 46 48 35.8081 $w=2.78e-07 $l=8.7e-07 $layer=LI1_cond $X=9.825 $Y=1.965
+ $X2=9.825 $Y2=2.835
r84 44 46 3.0869 $w=2.78e-07 $l=7.5e-08 $layer=LI1_cond $X=9.825 $Y=1.89
+ $X2=9.825 $Y2=1.965
r85 43 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.015 $Y=1.805
+ $X2=8.85 $Y2=1.805
r86 42 44 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=9.685 $Y=1.805
+ $X2=9.825 $Y2=1.89
r87 42 43 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.685 $Y=1.805
+ $X2=9.015 $Y2=1.805
r88 38 40 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=8.85 $Y=1.965
+ $X2=8.85 $Y2=2.835
r89 36 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.85 $Y=1.89 $X2=8.85
+ $Y2=1.805
r90 36 38 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=8.85 $Y=1.89
+ $X2=8.85 $Y2=1.965
r91 34 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.685 $Y=1.805
+ $X2=8.85 $Y2=1.805
r92 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.685 $Y=1.805
+ $X2=8.015 $Y2=1.805
r93 31 33 35.8081 $w=2.78e-07 $l=8.7e-07 $layer=LI1_cond $X=7.875 $Y=1.965
+ $X2=7.875 $Y2=2.835
r94 29 33 2.88111 $w=2.78e-07 $l=7e-08 $layer=LI1_cond $X=7.875 $Y=2.905
+ $X2=7.875 $Y2=2.835
r95 28 35 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=7.875 $Y=1.89
+ $X2=8.015 $Y2=1.805
r96 28 31 3.0869 $w=2.78e-07 $l=7.5e-08 $layer=LI1_cond $X=7.875 $Y=1.89
+ $X2=7.875 $Y2=1.965
r97 27 50 8.35232 $w=1.77e-07 $l=1.68953e-07 $layer=LI1_cond $X=7.165 $Y=2.99
+ $X2=7 $Y2=2.982
r98 26 29 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=7.735 $Y=2.99
+ $X2=7.875 $Y2=2.905
r99 26 27 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=7.735 $Y=2.99
+ $X2=7.165 $Y2=2.99
r100 22 50 0.762005 $w=3.3e-07 $l=9.2e-08 $layer=LI1_cond $X=7 $Y=2.89 $X2=7
+ $Y2=2.982
r101 22 24 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=7 $Y=2.89 $X2=7
+ $Y2=2.145
r102 20 50 8.35232 $w=1.77e-07 $l=1.65e-07 $layer=LI1_cond $X=6.835 $Y=2.982
+ $X2=7 $Y2=2.982
r103 20 21 34.172 $w=1.83e-07 $l=5.7e-07 $layer=LI1_cond $X=6.835 $Y=2.982
+ $X2=6.265 $Y2=2.982
r104 16 21 7.54394 $w=1.85e-07 $l=2.05925e-07 $layer=LI1_cond $X=6.1 $Y=2.89
+ $X2=6.265 $Y2=2.982
r105 16 18 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=6.1 $Y=2.89
+ $X2=6.1 $Y2=2.145
r106 5 48 400 $w=1.7e-07 $l=1.06035e-06 $layer=licon1_PDIFF $count=1 $X=9.665
+ $Y=1.84 $X2=9.8 $Y2=2.835
r107 5 46 400 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=9.665
+ $Y=1.84 $X2=9.8 $Y2=1.965
r108 4 40 400 $w=1.7e-07 $l=1.06035e-06 $layer=licon1_PDIFF $count=1 $X=8.715
+ $Y=1.84 $X2=8.85 $Y2=2.835
r109 4 38 400 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=8.715
+ $Y=1.84 $X2=8.85 $Y2=1.965
r110 3 33 400 $w=1.7e-07 $l=1.06035e-06 $layer=licon1_PDIFF $count=1 $X=7.765
+ $Y=1.84 $X2=7.9 $Y2=2.835
r111 3 31 400 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_PDIFF $count=1 $X=7.765
+ $Y=1.84 $X2=7.9 $Y2=1.965
r112 2 24 300 $w=1.7e-07 $l=3.66333e-07 $layer=licon1_PDIFF $count=2 $X=6.865
+ $Y=1.84 $X2=7 $Y2=2.145
r113 1 18 300 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_PDIFF $count=2 $X=5.955
+ $Y=1.84 $X2=6.1 $Y2=2.145
.ends

.subckt PM_SKY130_FD_SC_MS__O41AI_4%A_27_74# 1 2 3 4 5 6 7 8 9 10 11 36 38 39 40
+ 45 46 47 50 53 54 55 58 61 62 66 68 72 74 78 80 84 86 90 92 94 96 98 103 104
+ 106 108 110 112 113
c190 61 0 1.95112e-19 $X=4.105 $Y=1.3
c191 53 0 1.97387e-19 $X=3.415 $Y=1.3
c192 40 0 6.95413e-20 $X=1.975 $Y=0.34
c193 38 0 6.95413e-20 $X=0.975 $Y=0.34
r194 98 101 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=1.14 $Y=0.34
+ $X2=1.14 $Y2=0.55
r195 94 115 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.84 $Y=0.84
+ $X2=9.84 $Y2=0.925
r196 94 96 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=9.84 $Y=0.84
+ $X2=9.84 $Y2=0.515
r197 93 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.035 $Y=0.925
+ $X2=8.87 $Y2=0.925
r198 92 115 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.715 $Y=0.925
+ $X2=9.84 $Y2=0.925
r199 92 93 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.715 $Y=0.925
+ $X2=9.035 $Y2=0.925
r200 88 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.87 $Y=0.84
+ $X2=8.87 $Y2=0.925
r201 88 90 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=8.87 $Y=0.84
+ $X2=8.87 $Y2=0.515
r202 87 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.035 $Y=0.925
+ $X2=7.91 $Y2=0.925
r203 86 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.705 $Y=0.925
+ $X2=8.87 $Y2=0.925
r204 86 87 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.705 $Y=0.925
+ $X2=8.035 $Y2=0.925
r205 82 112 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.91 $Y=0.84
+ $X2=7.91 $Y2=0.925
r206 82 84 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=7.91 $Y=0.84
+ $X2=7.91 $Y2=0.515
r207 81 110 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.06 $Y=0.925
+ $X2=6.975 $Y2=0.925
r208 80 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.785 $Y=0.925
+ $X2=7.91 $Y2=0.925
r209 80 81 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=7.785 $Y=0.925
+ $X2=7.06 $Y2=0.925
r210 76 110 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.975 $Y=0.84
+ $X2=6.975 $Y2=0.925
r211 76 78 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=6.975 $Y=0.84
+ $X2=6.975 $Y2=0.515
r212 75 108 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.21 $Y=0.925
+ $X2=6.085 $Y2=0.925
r213 74 110 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=0.925
+ $X2=6.975 $Y2=0.925
r214 74 75 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.89 $Y=0.925
+ $X2=6.21 $Y2=0.925
r215 70 108 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.085 $Y=0.84
+ $X2=6.085 $Y2=0.925
r216 70 72 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=6.085 $Y=0.84
+ $X2=6.085 $Y2=0.515
r217 69 106 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.28 $Y=0.925
+ $X2=5.155 $Y2=0.925
r218 68 108 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.96 $Y=0.925
+ $X2=6.085 $Y2=0.925
r219 68 69 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.96 $Y=0.925
+ $X2=5.28 $Y2=0.925
r220 64 106 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.155 $Y=0.84
+ $X2=5.155 $Y2=0.925
r221 64 66 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=5.155 $Y=0.84
+ $X2=5.155 $Y2=0.515
r222 63 104 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.35 $Y=0.925
+ $X2=4.185 $Y2=0.925
r223 62 106 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.03 $Y=0.925
+ $X2=5.155 $Y2=0.925
r224 62 63 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.03 $Y=0.925
+ $X2=4.35 $Y2=0.925
r225 60 104 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.105 $Y=1.01
+ $X2=4.185 $Y2=0.925
r226 60 61 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.105 $Y=1.01
+ $X2=4.105 $Y2=1.3
r227 56 104 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.185 $Y=0.84
+ $X2=4.185 $Y2=0.925
r228 56 58 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.185 $Y=0.84
+ $X2=4.185 $Y2=0.515
r229 54 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.02 $Y=1.385
+ $X2=4.105 $Y2=1.3
r230 54 55 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.02 $Y=1.385
+ $X2=3.5 $Y2=1.385
r231 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.415 $Y=1.3
+ $X2=3.5 $Y2=1.385
r232 52 103 3.64284 $w=2.55e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.415 $Y=1.01
+ $X2=3.33 $Y2=0.925
r233 52 53 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.415 $Y=1.01
+ $X2=3.415 $Y2=1.3
r234 48 103 3.64284 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=0.84
+ $X2=3.33 $Y2=0.925
r235 48 50 11.016 $w=3.38e-07 $l=3.25e-07 $layer=LI1_cond $X=3.33 $Y=0.84
+ $X2=3.33 $Y2=0.515
r236 46 103 2.83584 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.16 $Y=0.925
+ $X2=3.33 $Y2=0.925
r237 46 47 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=3.16 $Y=0.925
+ $X2=2.305 $Y2=0.925
r238 43 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.14 $Y=0.84
+ $X2=2.305 $Y2=0.925
r239 43 45 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.14 $Y=0.84
+ $X2=2.14 $Y2=0.515
r240 42 45 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.14 $Y=0.425
+ $X2=2.14 $Y2=0.515
r241 41 98 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=0.34
+ $X2=1.14 $Y2=0.34
r242 40 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.975 $Y=0.34
+ $X2=2.14 $Y2=0.425
r243 40 41 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.975 $Y=0.34
+ $X2=1.305 $Y2=0.34
r244 38 98 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0.34
+ $X2=1.14 $Y2=0.34
r245 38 39 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=0.975 $Y=0.34
+ $X2=0.445 $Y2=0.34
r246 34 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.425
+ $X2=0.445 $Y2=0.34
r247 34 36 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=0.425
+ $X2=0.28 $Y2=0.515
r248 11 115 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=9.66
+ $Y=0.37 $X2=9.8 $Y2=0.925
r249 11 96 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=9.66
+ $Y=0.37 $X2=9.8 $Y2=0.515
r250 10 90 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.73
+ $Y=0.37 $X2=8.87 $Y2=0.515
r251 9 112 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=7.73
+ $Y=0.37 $X2=7.87 $Y2=0.925
r252 9 84 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.73
+ $Y=0.37 $X2=7.87 $Y2=0.515
r253 8 110 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=6.835
+ $Y=0.37 $X2=6.975 $Y2=0.925
r254 8 78 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.835
+ $Y=0.37 $X2=6.975 $Y2=0.515
r255 7 108 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=5.905
+ $Y=0.37 $X2=6.045 $Y2=0.925
r256 7 72 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.905
+ $Y=0.37 $X2=6.045 $Y2=0.515
r257 6 106 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=4.975
+ $Y=0.37 $X2=5.115 $Y2=0.925
r258 6 66 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.975
+ $Y=0.37 $X2=5.115 $Y2=0.515
r259 5 58 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.045
+ $Y=0.37 $X2=4.185 $Y2=0.515
r260 4 50 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=3.16
+ $Y=0.37 $X2=3.325 $Y2=0.515
r261 3 45 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=1.93
+ $Y=0.37 $X2=2.14 $Y2=0.515
r262 2 101 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=1 $Y=0.37
+ $X2=1.14 $Y2=0.55
r263 1 36 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O41AI_4%VGND 1 2 3 4 5 6 7 8 27 29 33 35 39 43 47 51
+ 55 57 58 59 61 73 78 83 88 95 96 106 109 112 115 118 121
r149 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r150 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r151 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r152 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r153 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r154 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r155 96 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=9.36 $Y2=0
r156 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r157 93 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.535 $Y=0
+ $X2=9.37 $Y2=0
r158 93 95 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.535 $Y=0
+ $X2=9.84 $Y2=0
r159 92 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r160 92 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r161 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r162 89 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.535 $Y=0
+ $X2=8.37 $Y2=0
r163 89 91 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.535 $Y=0 $X2=8.88
+ $Y2=0
r164 88 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.205 $Y=0
+ $X2=9.37 $Y2=0
r165 88 91 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.205 $Y=0
+ $X2=8.88 $Y2=0
r166 87 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r167 87 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r168 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r169 84 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.57 $Y=0
+ $X2=7.405 $Y2=0
r170 84 86 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=7.57 $Y=0 $X2=7.92
+ $Y2=0
r171 83 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.205 $Y=0
+ $X2=8.37 $Y2=0
r172 83 86 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=8.205 $Y=0
+ $X2=7.92 $Y2=0
r173 82 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r174 82 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=6.48 $Y2=0
r175 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r176 79 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.71 $Y=0
+ $X2=6.545 $Y2=0
r177 79 81 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.71 $Y=0 $X2=6.96
+ $Y2=0
r178 78 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.24 $Y=0
+ $X2=7.405 $Y2=0
r179 78 81 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.24 $Y=0 $X2=6.96
+ $Y2=0
r180 77 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r181 77 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r182 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r183 74 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.78 $Y=0
+ $X2=5.615 $Y2=0
r184 74 76 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.78 $Y=0 $X2=6
+ $Y2=0
r185 73 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.38 $Y=0
+ $X2=6.545 $Y2=0
r186 73 76 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.38 $Y=0 $X2=6
+ $Y2=0
r187 72 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r188 72 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r189 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r190 69 71 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.99 $Y=0 $X2=3.6
+ $Y2=0
r191 68 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=2.64 $Y2=0
r192 67 68 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r193 64 68 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=2.16 $Y2=0
r194 63 67 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r195 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r196 61 103 11.9608 $w=5.13e-07 $l=5.15e-07 $layer=LI1_cond $X=2.732 $Y=0
+ $X2=2.732 $Y2=0.515
r197 61 69 7.34265 $w=1.7e-07 $l=2.58e-07 $layer=LI1_cond $X=2.732 $Y=0 $X2=2.99
+ $Y2=0
r198 61 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r199 61 67 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.475 $Y=0
+ $X2=2.16 $Y2=0
r200 59 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r201 59 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=4.56 $Y2=0
r202 57 71 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.67 $Y=0 $X2=3.6
+ $Y2=0
r203 57 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=0 $X2=3.755
+ $Y2=0
r204 53 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.37 $Y=0.085
+ $X2=9.37 $Y2=0
r205 53 55 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=9.37 $Y=0.085
+ $X2=9.37 $Y2=0.55
r206 49 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.37 $Y=0.085
+ $X2=8.37 $Y2=0
r207 49 51 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=8.37 $Y=0.085
+ $X2=8.37 $Y2=0.55
r208 45 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.405 $Y=0.085
+ $X2=7.405 $Y2=0
r209 45 47 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=7.405 $Y=0.085
+ $X2=7.405 $Y2=0.55
r210 41 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.545 $Y=0.085
+ $X2=6.545 $Y2=0
r211 41 43 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=6.545 $Y=0.085
+ $X2=6.545 $Y2=0.55
r212 37 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.615 $Y=0.085
+ $X2=5.615 $Y2=0
r213 37 39 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=5.615 $Y=0.085
+ $X2=5.615 $Y2=0.55
r214 36 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.85 $Y=0
+ $X2=4.685 $Y2=0
r215 35 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.45 $Y=0
+ $X2=5.615 $Y2=0
r216 35 36 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.45 $Y=0 $X2=4.85
+ $Y2=0
r217 31 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.685 $Y=0.085
+ $X2=4.685 $Y2=0
r218 31 33 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.685 $Y=0.085
+ $X2=4.685 $Y2=0.55
r219 30 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.84 $Y=0 $X2=3.755
+ $Y2=0
r220 29 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.52 $Y=0
+ $X2=4.685 $Y2=0
r221 29 30 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.52 $Y=0 $X2=3.84
+ $Y2=0
r222 25 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.755 $Y=0.085
+ $X2=3.755 $Y2=0
r223 25 27 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.755 $Y=0.085
+ $X2=3.755 $Y2=0.515
r224 8 55 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=9.16
+ $Y=0.37 $X2=9.37 $Y2=0.55
r225 7 51 182 $w=1.7e-07 $l=2.45561e-07 $layer=licon1_NDIFF $count=1 $X=8.215
+ $Y=0.37 $X2=8.37 $Y2=0.55
r226 6 47 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=7.265
+ $Y=0.37 $X2=7.405 $Y2=0.55
r227 5 43 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=6.335
+ $Y=0.37 $X2=6.545 $Y2=0.55
r228 4 39 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=5.405
+ $Y=0.37 $X2=5.615 $Y2=0.55
r229 3 33 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=4.475
+ $Y=0.37 $X2=4.685 $Y2=0.55
r230 2 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.615
+ $Y=0.37 $X2=3.755 $Y2=0.515
r231 1 103 182 $w=1.7e-07 $l=3.65377e-07 $layer=licon1_NDIFF $count=1 $X=2.43
+ $Y=0.37 $X2=2.73 $Y2=0.515
.ends


* File: sky130_fd_sc_ms__nor2_8.pex.spice
* Created: Wed Sep  2 12:15:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NOR2_8%A 1 3 4 5 6 8 9 11 13 14 18 20 22 25 27 29 30
+ 32 35 37 39 42 44 46 47 48 49 50 51 52 53 72
c129 30 0 1.96393e-19 $X=2.855 $Y=1.725
c130 20 0 1.96393e-19 $X=1.905 $Y=1.725
c131 11 0 1.90646e-19 $X=1.455 $Y=1.725
c132 6 0 3.09093e-19 $X=1.005 $Y=1.725
r133 70 72 39.0447 $w=3.58e-07 $l=2.9e-07 $layer=POLY_cond $X=3.42 $Y=1.537
+ $X2=3.71 $Y2=1.537
r134 70 71 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.42
+ $Y=1.515 $X2=3.42 $Y2=1.515
r135 68 70 15.4832 $w=3.58e-07 $l=1.15e-07 $layer=POLY_cond $X=3.305 $Y=1.537
+ $X2=3.42 $Y2=1.537
r136 67 68 12.7905 $w=3.58e-07 $l=9.5e-08 $layer=POLY_cond $X=3.21 $Y=1.537
+ $X2=3.305 $Y2=1.537
r137 66 67 47.7961 $w=3.58e-07 $l=3.55e-07 $layer=POLY_cond $X=2.855 $Y=1.537
+ $X2=3.21 $Y2=1.537
r138 65 66 67.3184 $w=3.58e-07 $l=5e-07 $layer=POLY_cond $X=2.355 $Y=1.537
+ $X2=2.855 $Y2=1.537
r139 64 65 6.05866 $w=3.58e-07 $l=4.5e-08 $layer=POLY_cond $X=2.31 $Y=1.537
+ $X2=2.355 $Y2=1.537
r140 62 64 33.6592 $w=3.58e-07 $l=2.5e-07 $layer=POLY_cond $X=2.06 $Y=1.537
+ $X2=2.31 $Y2=1.537
r141 62 63 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.06
+ $Y=1.515 $X2=2.06 $Y2=1.515
r142 60 62 20.8687 $w=3.58e-07 $l=1.55e-07 $layer=POLY_cond $X=1.905 $Y=1.537
+ $X2=2.06 $Y2=1.537
r143 59 60 12.7905 $w=3.58e-07 $l=9.5e-08 $layer=POLY_cond $X=1.81 $Y=1.537
+ $X2=1.905 $Y2=1.537
r144 53 71 4.82418 $w=4.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.6 $Y=1.565
+ $X2=3.42 $Y2=1.565
r145 52 71 8.0403 $w=4.28e-07 $l=3e-07 $layer=LI1_cond $X=3.12 $Y=1.565 $X2=3.42
+ $Y2=1.565
r146 51 52 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.12 $Y2=1.565
r147 50 51 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.565
+ $X2=2.64 $Y2=1.565
r148 50 63 2.6801 $w=4.28e-07 $l=1e-07 $layer=LI1_cond $X=2.16 $Y=1.565 $X2=2.06
+ $Y2=1.565
r149 49 63 10.1844 $w=4.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.68 $Y=1.565
+ $X2=2.06 $Y2=1.565
r150 44 72 19.5223 $w=3.58e-07 $l=2.50208e-07 $layer=POLY_cond $X=3.855 $Y=1.725
+ $X2=3.71 $Y2=1.537
r151 44 46 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.855 $Y=1.725
+ $X2=3.855 $Y2=2.4
r152 40 72 23.1716 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=3.71 $Y=1.35
+ $X2=3.71 $Y2=1.537
r153 40 42 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.71 $Y=1.35
+ $X2=3.71 $Y2=0.74
r154 37 68 18.8375 $w=1.8e-07 $l=1.88e-07 $layer=POLY_cond $X=3.305 $Y=1.725
+ $X2=3.305 $Y2=1.537
r155 37 39 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.305 $Y=1.725
+ $X2=3.305 $Y2=2.4
r156 33 67 23.1716 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=3.21 $Y=1.35
+ $X2=3.21 $Y2=1.537
r157 33 35 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.21 $Y=1.35
+ $X2=3.21 $Y2=0.74
r158 30 66 18.8375 $w=1.8e-07 $l=1.88e-07 $layer=POLY_cond $X=2.855 $Y=1.725
+ $X2=2.855 $Y2=1.537
r159 30 32 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=2.855 $Y=1.725
+ $X2=2.855 $Y2=2.4
r160 27 65 18.8375 $w=1.8e-07 $l=1.88e-07 $layer=POLY_cond $X=2.355 $Y=1.725
+ $X2=2.355 $Y2=1.537
r161 27 29 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=2.355 $Y=1.725
+ $X2=2.355 $Y2=2.4
r162 23 64 23.1716 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=2.31 $Y=1.35
+ $X2=2.31 $Y2=1.537
r163 23 25 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.31 $Y=1.35
+ $X2=2.31 $Y2=0.74
r164 20 60 18.8375 $w=1.8e-07 $l=1.88e-07 $layer=POLY_cond $X=1.905 $Y=1.725
+ $X2=1.905 $Y2=1.537
r165 20 22 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=1.905 $Y=1.725
+ $X2=1.905 $Y2=2.4
r166 16 59 23.1716 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=1.81 $Y=1.35
+ $X2=1.81 $Y2=1.537
r167 16 18 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.81 $Y=1.35
+ $X2=1.81 $Y2=0.74
r168 15 48 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.545 $Y=1.65
+ $X2=1.455 $Y2=1.65
r169 14 59 26.7661 $w=3.58e-07 $l=1.45753e-07 $layer=POLY_cond $X=1.735 $Y=1.65
+ $X2=1.81 $Y2=1.537
r170 14 15 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.735 $Y=1.65
+ $X2=1.545 $Y2=1.65
r171 11 48 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=1.455 $Y=1.725
+ $X2=1.455 $Y2=1.65
r172 11 13 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=1.455 $Y=1.725
+ $X2=1.455 $Y2=2.4
r173 10 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.095 $Y=1.65
+ $X2=1.005 $Y2=1.65
r174 9 48 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.365 $Y=1.65
+ $X2=1.455 $Y2=1.65
r175 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.365 $Y=1.65
+ $X2=1.095 $Y2=1.65
r176 6 47 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=1.005 $Y=1.725
+ $X2=1.005 $Y2=1.65
r177 6 8 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=1.005 $Y=1.725
+ $X2=1.005 $Y2=2.4
r178 4 47 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.915 $Y=1.65
+ $X2=1.005 $Y2=1.65
r179 4 5 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.915 $Y=1.65
+ $X2=0.595 $Y2=1.65
r180 1 5 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=0.505 $Y=1.725
+ $X2=0.595 $Y2=1.65
r181 1 3 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=0.505 $Y=1.725
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__NOR2_8%B 1 3 6 8 12 14 18 20 22 23 27 29 31 34 36 38
+ 39 40 43 45 49 53 55 56 57 62 64 66 67 71 72
r134 75 76 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.39
+ $Y=1.145 $X2=7.39 $Y2=1.145
r135 71 75 57.7492 $w=6.3e-07 $l=6.8e-07 $layer=POLY_cond $X=7.38 $Y=0.465
+ $X2=7.38 $Y2=1.145
r136 71 72 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.39
+ $Y=0.465 $X2=7.39 $Y2=0.465
r137 67 76 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=7.39 $Y=0.925
+ $X2=7.39 $Y2=1.145
r138 66 67 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=7.39 $Y=0.555
+ $X2=7.39 $Y2=0.925
r139 66 72 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=7.39 $Y=0.555
+ $X2=7.39 $Y2=0.465
r140 63 75 3.39701 $w=6.3e-07 $l=4e-08 $layer=POLY_cond $X=7.38 $Y=1.185
+ $X2=7.38 $Y2=1.145
r141 63 64 6.3694 $w=6.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.38 $Y=1.185
+ $X2=7.38 $Y2=1.26
r142 47 64 36.8168 $w=6.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.38 $Y=1.335
+ $X2=7.38 $Y2=1.26
r143 47 53 413.976 $w=1.8e-07 $l=1.065e-06 $layer=POLY_cond $X=7.605 $Y=1.335
+ $X2=7.605 $Y2=2.4
r144 47 49 413.976 $w=1.8e-07 $l=1.065e-06 $layer=POLY_cond $X=7.155 $Y=1.335
+ $X2=7.155 $Y2=2.4
r145 46 62 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.745 $Y=1.26
+ $X2=6.655 $Y2=1.26
r146 45 64 37.3437 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=7.065 $Y=1.26
+ $X2=7.38 $Y2=1.26
r147 45 46 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.065 $Y=1.26
+ $X2=6.745 $Y2=1.26
r148 41 62 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=6.655 $Y=1.335
+ $X2=6.655 $Y2=1.26
r149 41 43 413.976 $w=1.8e-07 $l=1.065e-06 $layer=POLY_cond $X=6.655 $Y=1.335
+ $X2=6.655 $Y2=2.4
r150 40 61 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.4 $Y=1.26
+ $X2=6.325 $Y2=1.26
r151 39 62 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.565 $Y=1.26
+ $X2=6.655 $Y2=1.26
r152 39 40 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.565 $Y=1.26
+ $X2=6.4 $Y2=1.26
r153 36 61 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.325 $Y=1.185
+ $X2=6.325 $Y2=1.26
r154 36 38 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=6.325 $Y=1.185
+ $X2=6.325 $Y2=0.74
r155 32 61 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=6.205 $Y=1.26
+ $X2=6.325 $Y2=1.26
r156 32 59 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=6.205 $Y=1.26
+ $X2=5.895 $Y2=1.26
r157 32 34 413.976 $w=1.8e-07 $l=1.065e-06 $layer=POLY_cond $X=6.205 $Y=1.335
+ $X2=6.205 $Y2=2.4
r158 29 59 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.895 $Y=1.185
+ $X2=5.895 $Y2=1.26
r159 29 31 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.895 $Y=1.185
+ $X2=5.895 $Y2=0.74
r160 25 59 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=5.755 $Y=1.26
+ $X2=5.895 $Y2=1.26
r161 25 27 413.976 $w=1.8e-07 $l=1.065e-06 $layer=POLY_cond $X=5.755 $Y=1.335
+ $X2=5.755 $Y2=2.4
r162 24 57 13.2179 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=5.4 $Y=1.26
+ $X2=5.307 $Y2=1.26
r163 23 25 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.665 $Y=1.26
+ $X2=5.755 $Y2=1.26
r164 23 24 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=5.665 $Y=1.26
+ $X2=5.4 $Y2=1.26
r165 20 57 10.9219 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=5.325 $Y=1.185
+ $X2=5.307 $Y2=1.26
r166 20 22 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.325 $Y=1.185
+ $X2=5.325 $Y2=0.74
r167 16 57 10.9219 $w=1.8e-07 $l=7.59934e-08 $layer=POLY_cond $X=5.305 $Y=1.335
+ $X2=5.307 $Y2=1.26
r168 16 18 413.976 $w=1.8e-07 $l=1.065e-06 $layer=POLY_cond $X=5.305 $Y=1.335
+ $X2=5.305 $Y2=2.4
r169 15 56 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.895 $Y=1.26
+ $X2=4.805 $Y2=1.26
r170 14 57 13.2179 $w=1.5e-07 $l=9.2e-08 $layer=POLY_cond $X=5.215 $Y=1.26
+ $X2=5.307 $Y2=1.26
r171 14 15 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.215 $Y=1.26
+ $X2=4.895 $Y2=1.26
r172 10 56 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.805 $Y=1.335
+ $X2=4.805 $Y2=1.26
r173 10 12 413.976 $w=1.8e-07 $l=1.065e-06 $layer=POLY_cond $X=4.805 $Y=1.335
+ $X2=4.805 $Y2=2.4
r174 9 55 6.66866 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=4.395 $Y=1.26
+ $X2=4.265 $Y2=1.26
r175 8 56 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.715 $Y=1.26
+ $X2=4.805 $Y2=1.26
r176 8 9 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.715 $Y=1.26
+ $X2=4.395 $Y2=1.26
r177 4 55 18.8402 $w=1.65e-07 $l=9.28709e-08 $layer=POLY_cond $X=4.305 $Y=1.335
+ $X2=4.265 $Y2=1.26
r178 4 6 413.976 $w=1.8e-07 $l=1.065e-06 $layer=POLY_cond $X=4.305 $Y=1.335
+ $X2=4.305 $Y2=2.4
r179 1 55 18.8402 $w=1.65e-07 $l=9.87421e-08 $layer=POLY_cond $X=4.21 $Y=1.185
+ $X2=4.265 $Y2=1.26
r180 1 3 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=4.21 $Y=1.185
+ $X2=4.21 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__NOR2_8%A_27_368# 1 2 3 4 5 6 7 8 9 30 34 35 38 40 44
+ 46 50 52 54 57 58 59 62 66 70 74 78 82 86 90 95 97 100 101 102
c130 90 0 1.18447e-19 $X=1.23 $Y=1.865
c131 50 0 1.96393e-19 $X=3.08 $Y=2.435
c132 44 0 1.96393e-19 $X=2.13 $Y=2.435
c133 38 0 3.81292e-19 $X=1.23 $Y=2.435
r134 90 93 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.23 $Y=1.865
+ $X2=1.23 $Y2=2.035
r135 86 89 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=7.88 $Y=1.985
+ $X2=7.88 $Y2=2.815
r136 84 89 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=7.88 $Y=2.905
+ $X2=7.88 $Y2=2.815
r137 83 102 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.035 $Y=2.99
+ $X2=6.905 $Y2=2.99
r138 82 84 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.715 $Y=2.99
+ $X2=7.88 $Y2=2.905
r139 82 83 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.715 $Y=2.99
+ $X2=7.035 $Y2=2.99
r140 78 81 36.7895 $w=2.58e-07 $l=8.3e-07 $layer=LI1_cond $X=6.905 $Y=1.985
+ $X2=6.905 $Y2=2.815
r141 76 102 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.905 $Y=2.905
+ $X2=6.905 $Y2=2.99
r142 76 81 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=6.905 $Y=2.905
+ $X2=6.905 $Y2=2.815
r143 75 101 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=6.08 $Y=2.99
+ $X2=5.977 $Y2=2.99
r144 74 102 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.775 $Y=2.99
+ $X2=6.905 $Y2=2.99
r145 74 75 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.775 $Y=2.99
+ $X2=6.08 $Y2=2.99
r146 70 73 44.9047 $w=2.03e-07 $l=8.3e-07 $layer=LI1_cond $X=5.977 $Y=1.985
+ $X2=5.977 $Y2=2.815
r147 68 101 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.977 $Y=2.905
+ $X2=5.977 $Y2=2.99
r148 68 73 4.86918 $w=2.03e-07 $l=9e-08 $layer=LI1_cond $X=5.977 $Y=2.905
+ $X2=5.977 $Y2=2.815
r149 67 100 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.185 $Y=2.99
+ $X2=5.055 $Y2=2.99
r150 66 101 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=5.875 $Y=2.99
+ $X2=5.977 $Y2=2.99
r151 66 67 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.875 $Y=2.99
+ $X2=5.185 $Y2=2.99
r152 62 65 31.0273 $w=2.58e-07 $l=7e-07 $layer=LI1_cond $X=5.055 $Y=2.115
+ $X2=5.055 $Y2=2.815
r153 60 100 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.055 $Y=2.905
+ $X2=5.055 $Y2=2.99
r154 60 65 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=5.055 $Y=2.905
+ $X2=5.055 $Y2=2.815
r155 58 100 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.925 $Y=2.99
+ $X2=5.055 $Y2=2.99
r156 58 59 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.925 $Y=2.99
+ $X2=4.245 $Y2=2.99
r157 55 59 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.08 $Y=2.905
+ $X2=4.245 $Y2=2.99
r158 55 57 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.08 $Y=2.905
+ $X2=4.08 $Y2=2.815
r159 54 99 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.08 $Y=2.12 $X2=4.08
+ $Y2=2.035
r160 54 57 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.08 $Y=2.12
+ $X2=4.08 $Y2=2.815
r161 53 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.245 $Y=2.035
+ $X2=3.12 $Y2=2.035
r162 52 99 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.915 $Y=2.035
+ $X2=4.08 $Y2=2.035
r163 52 53 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.915 $Y=2.035
+ $X2=3.245 $Y2=2.035
r164 48 97 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=2.12
+ $X2=3.12 $Y2=2.035
r165 48 50 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=3.12 $Y=2.12
+ $X2=3.12 $Y2=2.435
r166 47 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.295 $Y=2.035
+ $X2=2.17 $Y2=2.035
r167 46 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.995 $Y=2.035
+ $X2=3.12 $Y2=2.035
r168 46 47 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.995 $Y=2.035
+ $X2=2.295 $Y2=2.035
r169 42 95 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=2.12
+ $X2=2.17 $Y2=2.035
r170 42 44 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=2.17 $Y=2.12
+ $X2=2.17 $Y2=2.435
r171 41 93 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.315 $Y=2.035
+ $X2=1.23 $Y2=2.035
r172 40 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.045 $Y=2.035
+ $X2=2.17 $Y2=2.035
r173 40 41 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.045 $Y=2.035
+ $X2=1.315 $Y2=2.035
r174 36 93 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=2.12
+ $X2=1.23 $Y2=2.035
r175 36 38 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.23 $Y=2.12
+ $X2=1.23 $Y2=2.435
r176 34 90 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=1.865
+ $X2=1.23 $Y2=1.865
r177 34 35 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.145 $Y=1.865
+ $X2=0.445 $Y2=1.865
r178 30 32 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.28 $Y=1.985
+ $X2=0.28 $Y2=2.815
r179 28 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=1.95
+ $X2=0.445 $Y2=1.865
r180 28 30 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.28 $Y=1.95
+ $X2=0.28 $Y2=1.985
r181 9 89 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=7.695
+ $Y=1.84 $X2=7.88 $Y2=2.815
r182 9 86 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=7.695
+ $Y=1.84 $X2=7.88 $Y2=1.985
r183 8 81 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.84 $X2=6.93 $Y2=2.815
r184 8 78 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.84 $X2=6.93 $Y2=1.985
r185 7 73 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.845
+ $Y=1.84 $X2=5.98 $Y2=2.815
r186 7 70 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.845
+ $Y=1.84 $X2=5.98 $Y2=1.985
r187 6 65 400 $w=1.7e-07 $l=1.06348e-06 $layer=licon1_PDIFF $count=1 $X=4.895
+ $Y=1.84 $X2=5.08 $Y2=2.815
r188 6 62 400 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_PDIFF $count=1 $X=4.895
+ $Y=1.84 $X2=5.08 $Y2=2.115
r189 5 99 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=3.945
+ $Y=1.84 $X2=4.08 $Y2=2.035
r190 5 57 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.945
+ $Y=1.84 $X2=4.08 $Y2=2.815
r191 4 97 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=2.945
+ $Y=1.84 $X2=3.08 $Y2=2.035
r192 4 50 300 $w=1.7e-07 $l=6.59052e-07 $layer=licon1_PDIFF $count=2 $X=2.945
+ $Y=1.84 $X2=3.08 $Y2=2.435
r193 3 95 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.84 $X2=2.13 $Y2=2.035
r194 3 44 300 $w=1.7e-07 $l=6.59052e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.84 $X2=2.13 $Y2=2.435
r195 2 93 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=1.84 $X2=1.23 $Y2=2.035
r196 2 38 300 $w=1.7e-07 $l=6.59052e-07 $layer=licon1_PDIFF $count=2 $X=1.095
+ $Y=1.84 $X2=1.23 $Y2=2.435
r197 1 32 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r198 1 30 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__NOR2_8%VPWR 1 2 3 4 15 19 23 27 29 31 36 41 46 56 57
+ 60 63 66 69
r99 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r100 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r101 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r102 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r103 56 57 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r104 53 56 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=7.92 $Y2=3.33
r105 51 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.745 $Y=3.33
+ $X2=3.58 $Y2=3.33
r106 51 53 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.745 $Y=3.33
+ $X2=4.08 $Y2=3.33
r107 50 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r108 50 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r109 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r110 47 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.795 $Y=3.33
+ $X2=2.63 $Y2=3.33
r111 47 49 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.795 $Y=3.33
+ $X2=3.12 $Y2=3.33
r112 46 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.415 $Y=3.33
+ $X2=3.58 $Y2=3.33
r113 46 49 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.415 $Y=3.33
+ $X2=3.12 $Y2=3.33
r114 45 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r115 45 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r116 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r117 42 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=1.68 $Y2=3.33
r118 42 44 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=2.16 $Y2=3.33
r119 41 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=3.33
+ $X2=2.63 $Y2=3.33
r120 41 44 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.465 $Y=3.33
+ $X2=2.16 $Y2=3.33
r121 40 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r122 40 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r123 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r124 37 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r125 37 39 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r126 36 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.515 $Y=3.33
+ $X2=1.68 $Y2=3.33
r127 36 39 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.515 $Y=3.33
+ $X2=1.2 $Y2=3.33
r128 34 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r129 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r130 31 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r131 31 33 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r132 29 57 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=7.92 $Y2=3.33
r133 29 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r134 29 53 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r135 25 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.58 $Y=3.245
+ $X2=3.58 $Y2=3.33
r136 25 27 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=3.58 $Y=3.245
+ $X2=3.58 $Y2=2.455
r137 21 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=3.245
+ $X2=2.63 $Y2=3.33
r138 21 23 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.63 $Y=3.245
+ $X2=2.63 $Y2=2.455
r139 17 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=3.245
+ $X2=1.68 $Y2=3.33
r140 17 19 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=1.68 $Y=3.245
+ $X2=1.68 $Y2=2.455
r141 13 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r142 13 15 33.5256 $w=3.28e-07 $l=9.6e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.285
r143 4 27 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=3.395
+ $Y=1.84 $X2=3.58 $Y2=2.455
r144 3 23 300 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_PDIFF $count=2 $X=2.445
+ $Y=1.84 $X2=2.63 $Y2=2.455
r145 2 19 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.84 $X2=1.68 $Y2=2.455
r146 1 15 300 $w=1.7e-07 $l=5.29481e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.84 $X2=0.78 $Y2=2.285
.ends

.subckt PM_SKY130_FD_SC_MS__NOR2_8%Y 1 2 3 4 5 6 7 8 27 29 30 33 35 39 45 51 55
+ 59 60 63 67 68 73
r109 76 77 5.99298 $w=8.55e-07 $l=4.2e-07 $layer=LI1_cond $X=5.11 $Y=1.14
+ $X2=5.53 $Y2=1.14
r110 74 76 7.56257 $w=8.55e-07 $l=5.3e-07 $layer=LI1_cond $X=4.58 $Y=1.14
+ $X2=5.11 $Y2=1.14
r111 73 74 0.28538 $w=8.55e-07 $l=2e-08 $layer=LI1_cond $X=4.56 $Y=1.14 $X2=4.58
+ $Y2=1.14
r112 71 73 1.92632 $w=8.55e-07 $l=1.35e-07 $layer=LI1_cond $X=4.425 $Y=1.14
+ $X2=4.56 $Y2=1.14
r113 68 73 10.6563 $w=1.7e-07 $l=5.25e-07 $layer=LI1_cond $X=4.56 $Y=1.665
+ $X2=4.56 $Y2=1.14
r114 63 65 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.38 $Y=1.97
+ $X2=7.38 $Y2=2.65
r115 61 63 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=7.38 $Y=1.65
+ $X2=7.38 $Y2=1.97
r116 59 61 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.215 $Y=1.565
+ $X2=7.38 $Y2=1.65
r117 59 60 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=7.215 $Y=1.565
+ $X2=6.595 $Y2=1.565
r118 55 57 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.43 $Y=1.97
+ $X2=6.43 $Y2=2.65
r119 53 60 12.0026 $w=8.55e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.43 $Y=1.65
+ $X2=6.595 $Y2=1.565
r120 53 55 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=6.43 $Y=1.65
+ $X2=6.43 $Y2=1.97
r121 49 53 4.56608 $w=8.55e-07 $l=6.50615e-07 $layer=LI1_cond $X=6.11 $Y=1.14
+ $X2=6.43 $Y2=1.65
r122 49 77 8.27602 $w=8.55e-07 $l=5.8e-07 $layer=LI1_cond $X=6.11 $Y=1.14
+ $X2=5.53 $Y2=1.14
r123 49 51 21.8266 $w=3.28e-07 $l=6.25e-07 $layer=LI1_cond $X=6.11 $Y=1.14
+ $X2=6.11 $Y2=0.515
r124 45 47 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.53 $Y=1.97
+ $X2=5.53 $Y2=2.65
r125 43 77 6.368 $w=3.3e-07 $l=6.4e-07 $layer=LI1_cond $X=5.53 $Y=1.78 $X2=5.53
+ $Y2=1.14
r126 43 45 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=5.53 $Y=1.78
+ $X2=5.53 $Y2=1.97
r127 39 41 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.58 $Y=1.97
+ $X2=4.58 $Y2=2.65
r128 37 74 6.368 $w=3.3e-07 $l=6.4e-07 $layer=LI1_cond $X=4.58 $Y=1.78 $X2=4.58
+ $Y2=1.14
r129 37 39 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.58 $Y=1.78
+ $X2=4.58 $Y2=1.97
r130 36 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.59 $Y=1.095
+ $X2=3.425 $Y2=1.095
r131 35 71 12.0026 $w=8.55e-07 $l=1.86145e-07 $layer=LI1_cond $X=4.26 $Y=1.095
+ $X2=4.425 $Y2=1.14
r132 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.26 $Y=1.095
+ $X2=3.59 $Y2=1.095
r133 31 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.425 $Y=1.01
+ $X2=3.425 $Y2=1.095
r134 31 33 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=3.425 $Y=1.01
+ $X2=3.425 $Y2=0.515
r135 29 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.26 $Y=1.095
+ $X2=3.425 $Y2=1.095
r136 29 30 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=3.26 $Y=1.095
+ $X2=2.19 $Y2=1.095
r137 25 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.025 $Y=1.01
+ $X2=2.19 $Y2=1.095
r138 25 27 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.025 $Y=1.01
+ $X2=2.025 $Y2=0.515
r139 8 65 400 $w=1.7e-07 $l=8.749e-07 $layer=licon1_PDIFF $count=1 $X=7.245
+ $Y=1.84 $X2=7.38 $Y2=2.65
r140 8 63 400 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_PDIFF $count=1 $X=7.245
+ $Y=1.84 $X2=7.38 $Y2=1.97
r141 7 57 400 $w=1.7e-07 $l=8.749e-07 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=1.84 $X2=6.43 $Y2=2.65
r142 7 55 400 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=1.84 $X2=6.43 $Y2=1.97
r143 6 47 400 $w=1.7e-07 $l=8.749e-07 $layer=licon1_PDIFF $count=1 $X=5.395
+ $Y=1.84 $X2=5.53 $Y2=2.65
r144 6 45 400 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_PDIFF $count=1 $X=5.395
+ $Y=1.84 $X2=5.53 $Y2=1.97
r145 5 41 400 $w=1.7e-07 $l=8.97747e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.84 $X2=4.58 $Y2=2.65
r146 5 39 400 $w=1.7e-07 $l=2.41402e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.84 $X2=4.58 $Y2=1.97
r147 4 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.97
+ $Y=0.37 $X2=6.11 $Y2=0.515
r148 3 76 60.6667 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_NDIFF $count=3
+ $X=4.285 $Y=0.37 $X2=5.11 $Y2=0.515
r149 3 71 60.6667 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=3
+ $X=4.285 $Y=0.37 $X2=4.425 $Y2=0.515
r150 2 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.285
+ $Y=0.37 $X2=3.425 $Y2=0.515
r151 1 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.885
+ $Y=0.37 $X2=2.025 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__NOR2_8%VGND 1 2 3 4 5 20 25 29 31 35 37 41 43 45 50
+ 60 61 64 69 72 75 78
r78 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r79 76 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r80 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r81 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r82 65 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r83 64 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r84 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r85 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r86 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r87 58 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r88 57 60 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r89 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r90 55 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.775 $Y=0 $X2=6.61
+ $Y2=0
r91 55 57 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=6.775 $Y=0 $X2=6.96
+ $Y2=0
r92 54 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r93 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r94 51 69 13.9655 $w=1.7e-07 $l=3.65e-07 $layer=LI1_cond $X=3.09 $Y=0 $X2=2.725
+ $Y2=0
r95 51 53 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.09 $Y=0 $X2=3.6
+ $Y2=0
r96 50 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.925
+ $Y2=0
r97 50 53 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.6
+ $Y2=0
r98 49 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r99 49 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r100 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r101 46 64 16.5844 $w=1.7e-07 $l=5.2e-07 $layer=LI1_cond $X=1.69 $Y=0 $X2=1.17
+ $Y2=0
r102 46 48 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=1.69 $Y=0 $X2=2.16
+ $Y2=0
r103 45 69 13.9655 $w=1.7e-07 $l=3.65e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.725
+ $Y2=0
r104 45 48 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.16
+ $Y2=0
r105 43 76 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=5.52 $Y2=0
r106 43 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r107 43 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r108 39 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.61 $Y=0.085
+ $X2=6.61 $Y2=0
r109 39 41 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=6.61 $Y=0.085
+ $X2=6.61 $Y2=0.515
r110 38 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.775 $Y=0 $X2=5.61
+ $Y2=0
r111 37 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.445 $Y=0 $X2=6.61
+ $Y2=0
r112 37 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.445 $Y=0
+ $X2=5.775 $Y2=0
r113 33 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.61 $Y=0.085
+ $X2=5.61 $Y2=0
r114 33 35 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.61 $Y=0.085
+ $X2=5.61 $Y2=0.515
r115 32 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.09 $Y=0 $X2=3.925
+ $Y2=0
r116 31 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.445 $Y=0 $X2=5.61
+ $Y2=0
r117 31 32 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=5.445 $Y=0
+ $X2=4.09 $Y2=0
r118 27 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.925 $Y=0.085
+ $X2=3.925 $Y2=0
r119 27 29 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=3.925 $Y=0.085
+ $X2=3.925 $Y2=0.675
r120 23 69 2.94957 $w=7.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=0.085
+ $X2=2.725 $Y2=0
r121 23 25 9.66693 $w=7.28e-07 $l=5.9e-07 $layer=LI1_cond $X=2.725 $Y=0.085
+ $X2=2.725 $Y2=0.675
r122 18 64 3.59326 $w=1.04e-06 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=0.085
+ $X2=1.17 $Y2=0
r123 18 20 5.04423 $w=1.038e-06 $l=4.3e-07 $layer=LI1_cond $X=1.17 $Y=0.085
+ $X2=1.17 $Y2=0.515
r124 5 41 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=6.4
+ $Y=0.37 $X2=6.61 $Y2=0.515
r125 4 35 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=5.4
+ $Y=0.37 $X2=5.61 $Y2=0.515
r126 3 29 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=3.785
+ $Y=0.37 $X2=3.925 $Y2=0.675
r127 2 25 91 $w=1.7e-07 $l=7.47094e-07 $layer=licon1_NDIFF $count=2 $X=2.385
+ $Y=0.37 $X2=2.995 $Y2=0.675
r128 1 20 60.6667 $w=1.7e-07 $l=9.94862e-07 $layer=licon1_NDIFF $count=3 $X=0.67
+ $Y=0.37 $X2=1.595 $Y2=0.515
r129 1 20 60.6667 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=3 $X=0.67
+ $Y=0.37 $X2=0.885 $Y2=0.515
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__a222o_1 A1 A2 B1 B2 C1 C2 VGND VNB VPB VPWR X
X0 a_340_390# B1 a_27_390# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X1 VPWR a_32_74# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X2 a_651_74# A2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X3 a_27_390# B2 a_340_390# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X4 a_119_74# C2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X5 a_32_74# C1 a_119_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 VPWR A1 a_340_390# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X7 a_32_74# A1 a_651_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 VGND a_32_74# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 a_386_74# B1 a_32_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X10 a_32_74# C2 a_27_390# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X11 VGND B2 a_386_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X12 a_27_390# C1 a_32_74# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X13 a_340_390# A2 VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
.ends

* File: sky130_fd_sc_ms__a31o_1.spice
* Created: Wed Sep  2 11:55:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a31o_1.pex.spice"
.subckt sky130_fd_sc_ms__a31o_1  VNB VPB A3 A2 A1 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_81_270#_M1006_g N_X_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.221517 AS=0.1961 PD=1.42638 PS=2.01 NRD=25.128 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75002.1 A=0.111 P=1.78 MULT=1
MM1008 A_265_120# N_A3_M1008_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.64 AD=0.0672
+ AS=0.191583 PD=0.85 PS=1.23362 NRD=9.372 NRS=29.52 M=1 R=4.26667 SA=75000.9
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1005 A_337_120# N_A2_M1005_g A_265_120# VNB NLOWVT L=0.15 W=0.64 AD=0.125625
+ AS=0.0672 PD=1.045 PS=0.85 NRD=26.484 NRS=9.372 M=1 R=4.26667 SA=75001.3
+ SB=75001.3 A=0.096 P=1.58 MULT=1
MM1009 N_A_81_270#_M1009_d N_A1_M1009_g A_337_120# VNB NLOWVT L=0.15 W=0.64
+ AD=0.1408 AS=0.125625 PD=1.08 PS=1.045 NRD=14.988 NRS=26.484 M=1 R=4.26667
+ SA=75001.8 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1000_d N_B1_M1000_g N_A_81_270#_M1009_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1696 AS=0.1408 PD=1.81 PS=1.08 NRD=0 NRS=14.988 M=1 R=4.26667 SA=75002.4
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_VPWR_M1007_d N_A_81_270#_M1007_g N_X_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.28 AS=0.2912 PD=1.7117 PS=2.76 NRD=19.3454 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90002.1 A=0.2016 P=2.6 MULT=1
MM1003 N_A_253_392#_M1003_d N_A3_M1003_g N_VPWR_M1007_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.25 PD=1.27 PS=1.5283 NRD=0 NRS=21.67 M=1 R=5.55556 SA=90000.8
+ SB=90001.7 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_A2_M1004_g N_A_253_392#_M1003_d VPB PSHORT L=0.18 W=1
+ AD=0.225 AS=0.135 PD=1.45 PS=1.27 NRD=16.7253 NRS=0 M=1 R=5.55556 SA=90001.3
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1001 N_A_253_392#_M1001_d N_A1_M1001_g N_VPWR_M1004_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.225 PD=1.27 PS=1.45 NRD=0 NRS=16.7253 M=1 R=5.55556 SA=90001.9
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1002 N_A_81_270#_M1002_d N_B1_M1002_g N_A_253_392#_M1001_d VPB PSHORT L=0.18
+ W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556 SA=90002.4
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__a31o_1.pxi.spice"
*
.ends
*
*

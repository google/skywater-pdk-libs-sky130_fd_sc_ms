* File: sky130_fd_sc_ms__nand4bb_2.spice
* Created: Fri Aug 28 17:46:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__nand4bb_2.pex.spice"
.subckt sky130_fd_sc_ms__nand4bb_2  VNB VPB A_N B_N C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B_N	B_N
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1018 N_VGND_M1018_d N_A_N_M1018_g N_A_27_368#_M1018_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1344 AS=0.1824 PD=1.06 PS=1.85 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.8 A=0.096 P=1.58 MULT=1
MM1005 N_A_231_74#_M1005_d N_B_N_M1005_g N_VGND_M1018_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.1344 PD=1.85 PS=1.06 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75000.8
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1012 N_A_373_74#_M1012_d N_A_27_368#_M1012_g N_Y_M1012_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2442 AS=0.11285 PD=2.14 PS=1.045 NRD=7.296 NRS=4.044 M=1 R=4.93333
+ SA=75000.3 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1016 N_A_373_74#_M1016_d N_A_27_368#_M1016_g N_Y_M1012_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1773 AS=0.11285 PD=1.28 PS=1.045 NRD=13.776 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1002 N_A_373_74#_M1016_d N_A_231_74#_M1002_g N_A_678_74#_M1002_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.1773 AS=0.1036 PD=1.28 PS=1.02 NRD=13.776 NRS=0 M=1
+ R=4.93333 SA=75001.3 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1015 N_A_373_74#_M1015_d N_A_231_74#_M1015_g N_A_678_74#_M1002_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2516 AS=0.1036 PD=2.16 PS=1.02 NRD=4.044 NRS=0 M=1
+ R=4.93333 SA=75001.7 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1013 N_A_886_74#_M1013_d N_C_M1013_g N_A_678_74#_M1013_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.2 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1019 N_A_886_74#_M1019_d N_C_M1019_g N_A_678_74#_M1013_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.7 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1006 N_A_886_74#_M1019_d N_D_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.1
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1009 N_A_886_74#_M1009_d N_D_M1009_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1295 PD=2.05 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 N_VPWR_M1010_d N_A_N_M1010_g N_A_27_368#_M1010_s VPB PSHORT L=0.18 W=1
+ AD=0.22725 AS=0.28 PD=1.49 PS=2.56 NRD=15.7403 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90000.9 A=0.18 P=2.36 MULT=1
MM1017 N_A_231_74#_M1017_d N_B_N_M1017_g N_VPWR_M1010_d VPB PSHORT L=0.18 W=1
+ AD=0.38 AS=0.22725 PD=2.76 PS=1.49 NRD=8.8453 NRS=15.7403 M=1 R=5.55556
+ SA=90000.8 SB=90000.3 A=0.18 P=2.36 MULT=1
MM1003 N_Y_M1003_d N_A_27_368#_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.2
+ SB=90004.1 A=0.2016 P=2.6 MULT=1
MM1007 N_Y_M1003_d N_A_27_368#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.7
+ SB=90003.7 A=0.2016 P=2.6 MULT=1
MM1000 N_Y_M1000_d N_A_231_74#_M1000_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90001.2
+ SB=90003.1 A=0.2016 P=2.6 MULT=1
MM1004 N_Y_M1000_d N_A_231_74#_M1004_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.448 PD=1.39 PS=1.92 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.7
+ SB=90002.7 A=0.2016 P=2.6 MULT=1
MM1001 N_Y_M1001_d N_C_M1001_g N_VPWR_M1004_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.448 PD=1.39 PS=1.92 NRD=0 NRS=0 M=1 R=6.22222 SA=90002.7 SB=90001.7
+ A=0.2016 P=2.6 MULT=1
MM1011 N_Y_M1001_d N_C_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12 AD=0.1512
+ AS=0.2072 PD=1.39 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003.1 SB=90001.2
+ A=0.2016 P=2.6 MULT=1
MM1008 N_Y_M1008_d N_D_M1008_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12 AD=0.1736
+ AS=0.2072 PD=1.43 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90003.7 SB=90000.7
+ A=0.2016 P=2.6 MULT=1
MM1014 N_Y_M1008_d N_D_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1.12 AD=0.1736
+ AS=0.3248 PD=1.43 PS=2.82 NRD=6.1464 NRS=0.8668 M=1 R=6.22222 SA=90004.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX20_noxref VNB VPB NWDIODE A=13.206 P=17.92
*
.include "sky130_fd_sc_ms__nand4bb_2.pxi.spice"
*
.ends
*
*

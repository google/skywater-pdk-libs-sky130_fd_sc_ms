* File: sky130_fd_sc_ms__ebufn_8.pxi.spice
* Created: Fri Aug 28 17:32:13 2020
* 
x_PM_SKY130_FD_SC_MS__EBUFN_8%A_84_48# N_A_84_48#_M1011_d N_A_84_48#_M1026_d
+ N_A_84_48#_M1007_g N_A_84_48#_M1001_g N_A_84_48#_M1013_g N_A_84_48#_M1002_g
+ N_A_84_48#_M1019_g N_A_84_48#_M1005_g N_A_84_48#_M1027_g N_A_84_48#_M1006_g
+ N_A_84_48#_M1030_g N_A_84_48#_M1008_g N_A_84_48#_M1012_g N_A_84_48#_M1031_g
+ N_A_84_48#_M1014_g N_A_84_48#_M1033_g N_A_84_48#_M1035_g N_A_84_48#_M1036_g
+ N_A_84_48#_c_342_p N_A_84_48#_c_230_n N_A_84_48#_c_242_n N_A_84_48#_c_256_p
+ N_A_84_48#_c_305_p N_A_84_48#_c_243_n N_A_84_48#_c_253_p N_A_84_48#_c_244_n
+ N_A_84_48#_c_288_p N_A_84_48#_c_231_n N_A_84_48#_c_293_p N_A_84_48#_c_245_n
+ N_A_84_48#_c_246_n N_A_84_48#_c_232_n N_A_84_48#_c_272_p N_A_84_48#_c_287_p
+ N_A_84_48#_c_233_n PM_SKY130_FD_SC_MS__EBUFN_8%A_84_48#
x_PM_SKY130_FD_SC_MS__EBUFN_8%A_833_48# N_A_833_48#_M1029_s N_A_833_48#_M1028_s
+ N_A_833_48#_c_490_n N_A_833_48#_M1000_g N_A_833_48#_c_491_n
+ N_A_833_48#_c_492_n N_A_833_48#_c_493_n N_A_833_48#_M1003_g
+ N_A_833_48#_c_494_n N_A_833_48#_c_495_n N_A_833_48#_M1004_g
+ N_A_833_48#_c_496_n N_A_833_48#_c_497_n N_A_833_48#_M1020_g
+ N_A_833_48#_c_498_n N_A_833_48#_c_499_n N_A_833_48#_M1024_g
+ N_A_833_48#_c_500_n N_A_833_48#_c_501_n N_A_833_48#_M1025_g
+ N_A_833_48#_c_502_n N_A_833_48#_c_503_n N_A_833_48#_M1034_g
+ N_A_833_48#_c_504_n N_A_833_48#_c_505_n N_A_833_48#_M1037_g
+ N_A_833_48#_c_506_n N_A_833_48#_c_507_n N_A_833_48#_c_508_n
+ N_A_833_48#_c_509_n N_A_833_48#_c_510_n N_A_833_48#_c_511_n
+ N_A_833_48#_c_512_n N_A_833_48#_c_513_n N_A_833_48#_c_514_n
+ N_A_833_48#_c_515_n N_A_833_48#_c_516_n N_A_833_48#_c_517_n
+ N_A_833_48#_c_518_n N_A_833_48#_c_519_n N_A_833_48#_c_525_n
+ N_A_833_48#_c_521_n PM_SKY130_FD_SC_MS__EBUFN_8%A_833_48#
x_PM_SKY130_FD_SC_MS__EBUFN_8%TE_B N_TE_B_c_676_n N_TE_B_M1009_g N_TE_B_c_655_n
+ N_TE_B_c_656_n N_TE_B_c_679_n N_TE_B_M1010_g N_TE_B_c_657_n N_TE_B_c_681_n
+ N_TE_B_M1015_g N_TE_B_c_658_n N_TE_B_c_683_n N_TE_B_M1016_g N_TE_B_c_659_n
+ N_TE_B_c_685_n N_TE_B_M1017_g N_TE_B_c_660_n N_TE_B_c_687_n N_TE_B_M1018_g
+ N_TE_B_c_661_n N_TE_B_c_689_n N_TE_B_M1021_g N_TE_B_c_662_n N_TE_B_c_691_n
+ N_TE_B_M1022_g N_TE_B_c_663_n N_TE_B_c_664_n N_TE_B_c_694_n N_TE_B_M1028_g
+ N_TE_B_c_665_n N_TE_B_M1029_g N_TE_B_c_666_n N_TE_B_c_667_n N_TE_B_c_668_n
+ N_TE_B_c_669_n N_TE_B_c_670_n N_TE_B_c_671_n N_TE_B_c_672_n TE_B TE_B TE_B
+ N_TE_B_c_674_n N_TE_B_c_675_n PM_SKY130_FD_SC_MS__EBUFN_8%TE_B
x_PM_SKY130_FD_SC_MS__EBUFN_8%A N_A_M1026_g N_A_c_838_n N_A_M1011_g N_A_M1032_g
+ N_A_c_840_n N_A_M1023_g A N_A_c_842_n PM_SKY130_FD_SC_MS__EBUFN_8%A
x_PM_SKY130_FD_SC_MS__EBUFN_8%A_28_368# N_A_28_368#_M1001_s N_A_28_368#_M1002_s
+ N_A_28_368#_M1006_s N_A_28_368#_M1012_s N_A_28_368#_M1035_s
+ N_A_28_368#_M1010_d N_A_28_368#_M1016_d N_A_28_368#_M1018_d
+ N_A_28_368#_M1022_d N_A_28_368#_c_887_n N_A_28_368#_c_888_n
+ N_A_28_368#_c_889_n N_A_28_368#_c_910_n N_A_28_368#_c_890_n
+ N_A_28_368#_c_971_p N_A_28_368#_c_891_n N_A_28_368#_c_974_p
+ N_A_28_368#_c_892_n N_A_28_368#_c_918_n N_A_28_368#_c_921_n
+ N_A_28_368#_c_923_n N_A_28_368#_c_924_n N_A_28_368#_c_925_n
+ N_A_28_368#_c_926_n N_A_28_368#_c_893_n N_A_28_368#_c_894_n
+ N_A_28_368#_c_895_n N_A_28_368#_c_896_n N_A_28_368#_c_897_n
+ N_A_28_368#_c_898_n N_A_28_368#_c_899_n PM_SKY130_FD_SC_MS__EBUFN_8%A_28_368#
x_PM_SKY130_FD_SC_MS__EBUFN_8%Z N_Z_M1007_s N_Z_M1019_s N_Z_M1030_s N_Z_M1033_s
+ N_Z_M1001_d N_Z_M1005_d N_Z_M1008_d N_Z_M1014_d N_Z_c_1038_n N_Z_c_1023_n
+ N_Z_c_1030_n N_Z_c_1049_n N_Z_c_1053_n N_Z_c_1024_n N_Z_c_1031_n N_Z_c_1063_n
+ N_Z_c_1067_n N_Z_c_1032_n N_Z_c_1025_n N_Z_c_1033_n N_Z_c_1083_n N_Z_c_1085_n
+ N_Z_c_1034_n N_Z_c_1026_n N_Z_c_1035_n N_Z_c_1036_n N_Z_c_1027_n Z Z Z
+ N_Z_c_1110_n Z PM_SKY130_FD_SC_MS__EBUFN_8%Z
x_PM_SKY130_FD_SC_MS__EBUFN_8%VPWR N_VPWR_M1009_s N_VPWR_M1015_s N_VPWR_M1017_s
+ N_VPWR_M1021_s N_VPWR_M1028_d N_VPWR_M1032_s N_VPWR_c_1153_n N_VPWR_c_1154_n
+ N_VPWR_c_1155_n N_VPWR_c_1156_n N_VPWR_c_1157_n N_VPWR_c_1158_n
+ N_VPWR_c_1159_n N_VPWR_c_1160_n VPWR N_VPWR_c_1161_n N_VPWR_c_1162_n
+ N_VPWR_c_1163_n N_VPWR_c_1164_n N_VPWR_c_1165_n N_VPWR_c_1166_n
+ N_VPWR_c_1167_n N_VPWR_c_1168_n N_VPWR_c_1169_n N_VPWR_c_1170_n
+ N_VPWR_c_1152_n PM_SKY130_FD_SC_MS__EBUFN_8%VPWR
x_PM_SKY130_FD_SC_MS__EBUFN_8%A_27_74# N_A_27_74#_M1007_d N_A_27_74#_M1013_d
+ N_A_27_74#_M1027_d N_A_27_74#_M1031_d N_A_27_74#_M1036_d N_A_27_74#_M1003_d
+ N_A_27_74#_M1020_d N_A_27_74#_M1025_d N_A_27_74#_M1037_d N_A_27_74#_c_1281_n
+ N_A_27_74#_c_1282_n N_A_27_74#_c_1283_n N_A_27_74#_c_1306_n
+ N_A_27_74#_c_1284_n N_A_27_74#_c_1309_n N_A_27_74#_c_1285_n
+ N_A_27_74#_c_1313_n N_A_27_74#_c_1286_n N_A_27_74#_c_1287_n
+ N_A_27_74#_c_1288_n N_A_27_74#_c_1289_n N_A_27_74#_c_1290_n
+ N_A_27_74#_c_1291_n N_A_27_74#_c_1292_n N_A_27_74#_c_1293_n
+ N_A_27_74#_c_1294_n N_A_27_74#_c_1295_n N_A_27_74#_c_1296_n
+ N_A_27_74#_c_1297_n N_A_27_74#_c_1298_n N_A_27_74#_c_1299_n
+ N_A_27_74#_c_1300_n N_A_27_74#_c_1301_n N_A_27_74#_c_1302_n
+ PM_SKY130_FD_SC_MS__EBUFN_8%A_27_74#
x_PM_SKY130_FD_SC_MS__EBUFN_8%VGND N_VGND_M1000_s N_VGND_M1004_s N_VGND_M1024_s
+ N_VGND_M1034_s N_VGND_M1029_d N_VGND_M1023_s N_VGND_c_1446_n N_VGND_c_1447_n
+ N_VGND_c_1448_n N_VGND_c_1449_n N_VGND_c_1450_n N_VGND_c_1451_n
+ N_VGND_c_1452_n N_VGND_c_1453_n N_VGND_c_1454_n N_VGND_c_1455_n
+ N_VGND_c_1456_n N_VGND_c_1457_n N_VGND_c_1458_n VGND N_VGND_c_1459_n
+ N_VGND_c_1460_n N_VGND_c_1461_n N_VGND_c_1462_n N_VGND_c_1463_n
+ N_VGND_c_1464_n PM_SKY130_FD_SC_MS__EBUFN_8%VGND
cc_1 VNB N_A_84_48#_M1007_g 0.02824f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_2 VNB N_A_84_48#_M1001_g 7.19436e-19 $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_3 VNB N_A_84_48#_M1013_g 0.0212213f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_4 VNB N_A_84_48#_M1002_g 4.76169e-19 $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_5 VNB N_A_84_48#_M1019_g 0.0212477f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=0.74
cc_6 VNB N_A_84_48#_M1005_g 4.96766e-19 $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=2.4
cc_7 VNB N_A_84_48#_M1027_g 0.0218518f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=0.74
cc_8 VNB N_A_84_48#_M1006_g 4.97118e-19 $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=2.4
cc_9 VNB N_A_84_48#_M1030_g 0.0227695f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=0.74
cc_10 VNB N_A_84_48#_M1008_g 4.78866e-19 $X=-0.19 $Y=-0.245 $X2=2.36 $Y2=2.4
cc_11 VNB N_A_84_48#_M1012_g 4.97118e-19 $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=2.4
cc_12 VNB N_A_84_48#_M1031_g 0.0229504f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=0.74
cc_13 VNB N_A_84_48#_M1014_g 5.09481e-19 $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=2.4
cc_14 VNB N_A_84_48#_M1033_g 0.0227562f $X=-0.19 $Y=-0.245 $X2=3.325 $Y2=0.74
cc_15 VNB N_A_84_48#_M1035_g 4.60318e-19 $X=-0.19 $Y=-0.245 $X2=3.795 $Y2=2.4
cc_16 VNB N_A_84_48#_M1036_g 0.022169f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=0.74
cc_17 VNB N_A_84_48#_c_230_n 0.00906377f $X=-0.19 $Y=-0.245 $X2=3.87 $Y2=1.565
cc_18 VNB N_A_84_48#_c_231_n 0.00210925f $X=-0.19 $Y=-0.245 $X2=9.845 $Y2=0.505
cc_19 VNB N_A_84_48#_c_232_n 0.0247114f $X=-0.19 $Y=-0.245 $X2=10.23 $Y2=1.72
cc_20 VNB N_A_84_48#_c_233_n 0.196838f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=1.485
cc_21 VNB N_A_833_48#_c_490_n 0.0145547f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.32
cc_22 VNB N_A_833_48#_c_491_n 0.0127756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_833_48#_c_492_n 0.00774194f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.65
cc_24 VNB N_A_833_48#_c_493_n 0.0143293f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_25 VNB N_A_833_48#_c_494_n 0.0109932f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.32
cc_26 VNB N_A_833_48#_c_495_n 0.0149279f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.74
cc_27 VNB N_A_833_48#_c_496_n 0.0102563f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_28 VNB N_A_833_48#_c_497_n 0.0149544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_833_48#_c_498_n 0.0109799f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=0.74
cc_30 VNB N_A_833_48#_c_499_n 0.0145943f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.65
cc_31 VNB N_A_833_48#_c_500_n 0.0102563f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_833_48#_c_501_n 0.0149561f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=0.74
cc_33 VNB N_A_833_48#_c_502_n 0.0109799f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=1.65
cc_34 VNB N_A_833_48#_c_503_n 0.0145943f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=2.4
cc_35 VNB N_A_833_48#_c_504_n 0.0102563f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=0.74
cc_36 VNB N_A_833_48#_c_505_n 0.0183025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_833_48#_c_506_n 0.0292022f $X=-0.19 $Y=-0.245 $X2=2.36 $Y2=2.4
cc_38 VNB N_A_833_48#_c_507_n 0.0299788f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=2.4
cc_39 VNB N_A_833_48#_c_508_n 0.00523367f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=2.4
cc_40 VNB N_A_833_48#_c_509_n 0.00436985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_833_48#_c_510_n 0.00436985f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=1.32
cc_42 VNB N_A_833_48#_c_511_n 0.00438315f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=0.74
cc_43 VNB N_A_833_48#_c_512_n 0.00436985f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=0.74
cc_44 VNB N_A_833_48#_c_513_n 0.00438315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_833_48#_c_514_n 0.00436985f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=1.65
cc_46 VNB N_A_833_48#_c_515_n 0.0152858f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=2.4
cc_47 VNB N_A_833_48#_c_516_n 0.020453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_833_48#_c_517_n 0.0111351f $X=-0.19 $Y=-0.245 $X2=3.325 $Y2=1.32
cc_49 VNB N_A_833_48#_c_518_n 0.0795427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_833_48#_c_519_n 0.0141642f $X=-0.19 $Y=-0.245 $X2=3.795 $Y2=2.4
cc_51 VNB N_TE_B_c_655_n 0.00891422f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_TE_B_c_656_n 0.0053384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_TE_B_c_657_n 0.00647609f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.74
cc_54 VNB N_TE_B_c_658_n 0.00886076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_TE_B_c_659_n 0.00649511f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.65
cc_56 VNB N_TE_B_c_660_n 0.00886067f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=0.74
cc_57 VNB N_TE_B_c_661_n 0.00649511f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=2.4
cc_58 VNB N_TE_B_c_662_n 0.0105865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_TE_B_c_663_n 0.0344152f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=0.74
cc_60 VNB N_TE_B_c_664_n 0.0283125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_TE_B_c_665_n 0.0227572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_TE_B_c_666_n 0.00439505f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=2.4
cc_63 VNB N_TE_B_c_667_n 0.00441496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_TE_B_c_668_n 0.00441486f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=1.32
cc_65 VNB N_TE_B_c_669_n 0.00441496f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=0.74
cc_66 VNB N_TE_B_c_670_n 0.00441496f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=0.74
cc_67 VNB N_TE_B_c_671_n 0.00441491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_TE_B_c_672_n 0.00681471f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=1.65
cc_69 VNB TE_B 0.0193491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_TE_B_c_674_n 0.0100304f $X=-0.19 $Y=-0.245 $X2=3.795 $Y2=2.4
cc_71 VNB N_TE_B_c_675_n 0.0234895f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=1.32
cc_72 VNB N_A_M1026_g 0.00619936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_c_838_n 0.0172452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_M1032_g 0.00628897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_c_840_n 0.0188503f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=2.4
cc_76 VNB A 0.0035636f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.32
cc_77 VNB N_A_c_842_n 0.0439932f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=0.74
cc_78 VNB N_Z_c_1023_n 0.00261517f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=2.4
cc_79 VNB N_Z_c_1024_n 0.00307912f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=0.74
cc_80 VNB N_Z_c_1025_n 0.00559895f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=1.65
cc_81 VNB N_Z_c_1026_n 0.00229628f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=0.74
cc_82 VNB N_Z_c_1027_n 0.00229411f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.485
cc_83 VNB Z 2.27624e-19 $X=-0.19 $Y=-0.245 $X2=3.87 $Y2=1.565
cc_84 VNB Z 0.00172469f $X=-0.19 $Y=-0.245 $X2=3.655 $Y2=1.565
cc_85 VNB N_VPWR_c_1152_n 0.442315f $X=-0.19 $Y=-0.245 $X2=9.93 $Y2=0.925
cc_86 VNB N_A_27_74#_c_1281_n 0.0362361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_27_74#_c_1282_n 0.0027626f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=0.74
cc_88 VNB N_A_27_74#_c_1283_n 0.00931596f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=0.74
cc_89 VNB N_A_27_74#_c_1284_n 0.0028694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_27_74#_c_1285_n 0.00280532f $X=-0.19 $Y=-0.245 $X2=2.36 $Y2=2.4
cc_91 VNB N_A_27_74#_c_1286_n 0.00488489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_27_74#_c_1287_n 4.66026e-19 $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=1.65
cc_93 VNB N_A_27_74#_c_1288_n 0.00627739f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=2.4
cc_94 VNB N_A_27_74#_c_1289_n 0.00583076f $X=-0.19 $Y=-0.245 $X2=3.31 $Y2=2.4
cc_95 VNB N_A_27_74#_c_1290_n 0.0023333f $X=-0.19 $Y=-0.245 $X2=3.325 $Y2=0.74
cc_96 VNB N_A_27_74#_c_1291_n 0.00528215f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_27_74#_c_1292_n 0.00263046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_27_74#_c_1293_n 0.00563126f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=0.74
cc_99 VNB N_A_27_74#_c_1294_n 0.00263046f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.485
cc_100 VNB N_A_27_74#_c_1295_n 0.00976772f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.485
cc_101 VNB N_A_27_74#_c_1296_n 0.00266546f $X=-0.19 $Y=-0.245 $X2=3.955 $Y2=1.65
cc_102 VNB N_A_27_74#_c_1297_n 0.00121874f $X=-0.19 $Y=-0.245 $X2=7.585
+ $Y2=2.135
cc_103 VNB N_A_27_74#_c_1298_n 0.00220535f $X=-0.19 $Y=-0.245 $X2=4.04 $Y2=2.135
cc_104 VNB N_A_27_74#_c_1299_n 0.00233543f $X=-0.19 $Y=-0.245 $X2=9.665
+ $Y2=2.305
cc_105 VNB N_A_27_74#_c_1300_n 0.0105845f $X=-0.19 $Y=-0.245 $X2=7.755 $Y2=2.305
cc_106 VNB N_A_27_74#_c_1301_n 0.00238685f $X=-0.19 $Y=-0.245 $X2=9.83 $Y2=1.985
cc_107 VNB N_A_27_74#_c_1302_n 0.00238685f $X=-0.19 $Y=-0.245 $X2=9.805 $Y2=2.39
cc_108 VNB N_VGND_c_1446_n 0.00334323f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=2.4
cc_109 VNB N_VGND_c_1447_n 0.00789915f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=0.74
cc_110 VNB N_VGND_c_1448_n 0.00582552f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=2.4
cc_111 VNB N_VGND_c_1449_n 0.00659784f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=0.74
cc_112 VNB N_VGND_c_1450_n 0.00719205f $X=-0.19 $Y=-0.245 $X2=1.91 $Y2=2.4
cc_113 VNB N_VGND_c_1451_n 0.0120978f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=1.32
cc_114 VNB N_VGND_c_1452_n 0.0189538f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=0.74
cc_115 VNB N_VGND_c_1453_n 0.0998102f $X=-0.19 $Y=-0.245 $X2=2.36 $Y2=2.4
cc_116 VNB N_VGND_c_1454_n 0.00604233f $X=-0.19 $Y=-0.245 $X2=2.36 $Y2=2.4
cc_117 VNB N_VGND_c_1455_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=1.65
cc_118 VNB N_VGND_c_1456_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=2.4
cc_119 VNB N_VGND_c_1457_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1458_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=2.81 $Y2=1.32
cc_121 VNB N_VGND_c_1459_n 0.0172524f $X=-0.19 $Y=-0.245 $X2=3.81 $Y2=1.32
cc_122 VNB N_VGND_c_1460_n 0.0569499f $X=-0.19 $Y=-0.245 $X2=3.49 $Y2=1.485
cc_123 VNB N_VGND_c_1461_n 0.0172141f $X=-0.19 $Y=-0.245 $X2=3.87 $Y2=1.565
cc_124 VNB N_VGND_c_1462_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=9.665 $Y2=2.305
cc_125 VNB N_VGND_c_1463_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=9.805 $Y2=2.22
cc_126 VNB N_VGND_c_1464_n 0.558924f $X=-0.19 $Y=-0.245 $X2=9.805 $Y2=2.815
cc_127 VPB N_A_84_48#_M1001_g 0.028056f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=2.4
cc_128 VPB N_A_84_48#_M1002_g 0.0213209f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_129 VPB N_A_84_48#_M1005_g 0.0219683f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=2.4
cc_130 VPB N_A_84_48#_M1006_g 0.0219916f $X=-0.19 $Y=1.66 $X2=1.91 $Y2=2.4
cc_131 VPB N_A_84_48#_M1008_g 0.0213688f $X=-0.19 $Y=1.66 $X2=2.36 $Y2=2.4
cc_132 VPB N_A_84_48#_M1012_g 0.0219916f $X=-0.19 $Y=1.66 $X2=2.81 $Y2=2.4
cc_133 VPB N_A_84_48#_M1014_g 0.0224243f $X=-0.19 $Y=1.66 $X2=3.31 $Y2=2.4
cc_134 VPB N_A_84_48#_M1035_g 0.0214723f $X=-0.19 $Y=1.66 $X2=3.795 $Y2=2.4
cc_135 VPB N_A_84_48#_c_242_n 0.00168561f $X=-0.19 $Y=1.66 $X2=3.955 $Y2=2.05
cc_136 VPB N_A_84_48#_c_243_n 0.0123659f $X=-0.19 $Y=1.66 $X2=9.665 $Y2=2.305
cc_137 VPB N_A_84_48#_c_244_n 0.00229053f $X=-0.19 $Y=1.66 $X2=9.83 $Y2=2.815
cc_138 VPB N_A_84_48#_c_245_n 0.00503473f $X=-0.19 $Y=1.66 $X2=10.145 $Y2=1.805
cc_139 VPB N_A_84_48#_c_246_n 0.00205111f $X=-0.19 $Y=1.66 $X2=9.945 $Y2=1.805
cc_140 VPB N_A_84_48#_c_232_n 0.00255885f $X=-0.19 $Y=1.66 $X2=10.23 $Y2=1.72
cc_141 VPB N_A_833_48#_c_516_n 0.00116802f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_833_48#_c_521_n 0.0122037f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=0.74
cc_143 VPB N_TE_B_c_676_n 0.0174312f $X=-0.19 $Y=1.66 $X2=9.705 $Y2=0.37
cc_144 VPB N_TE_B_c_655_n 0.00867498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_145 VPB N_TE_B_c_656_n 0.00409831f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_146 VPB N_TE_B_c_679_n 0.0175592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_147 VPB N_TE_B_c_657_n 0.00515318f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.74
cc_148 VPB N_TE_B_c_681_n 0.017561f $X=-0.19 $Y=1.66 $X2=0.51 $Y2=1.65
cc_149 VPB N_TE_B_c_658_n 0.00867498f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_TE_B_c_683_n 0.017561f $X=-0.19 $Y=1.66 $X2=0.925 $Y2=0.74
cc_151 VPB N_TE_B_c_659_n 0.00515318f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=1.65
cc_152 VPB N_TE_B_c_685_n 0.017561f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_153 VPB N_TE_B_c_660_n 0.00867498f $X=-0.19 $Y=1.66 $X2=1.38 $Y2=0.74
cc_154 VPB N_TE_B_c_687_n 0.017562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_TE_B_c_661_n 0.00515318f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=2.4
cc_156 VPB N_TE_B_c_689_n 0.0180248f $X=-0.19 $Y=1.66 $X2=1.81 $Y2=1.32
cc_157 VPB N_TE_B_c_662_n 0.0111142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_158 VPB N_TE_B_c_691_n 0.0224806f $X=-0.19 $Y=1.66 $X2=1.91 $Y2=2.4
cc_159 VPB N_TE_B_c_663_n 0.014664f $X=-0.19 $Y=1.66 $X2=2.31 $Y2=0.74
cc_160 VPB N_TE_B_c_664_n 0.00960941f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_TE_B_c_694_n 0.0222086f $X=-0.19 $Y=1.66 $X2=2.36 $Y2=1.65
cc_162 VPB N_TE_B_c_666_n 0.00200584f $X=-0.19 $Y=1.66 $X2=2.81 $Y2=2.4
cc_163 VPB N_TE_B_c_667_n 0.00200584f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_164 VPB N_TE_B_c_668_n 0.00200584f $X=-0.19 $Y=1.66 $X2=2.81 $Y2=1.32
cc_165 VPB N_TE_B_c_669_n 0.00200584f $X=-0.19 $Y=1.66 $X2=2.81 $Y2=0.74
cc_166 VPB N_TE_B_c_670_n 0.00200584f $X=-0.19 $Y=1.66 $X2=2.81 $Y2=0.74
cc_167 VPB N_TE_B_c_671_n 0.00200584f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_TE_B_c_672_n 0.00200584f $X=-0.19 $Y=1.66 $X2=3.31 $Y2=1.65
cc_169 VPB N_TE_B_c_674_n 0.00782129f $X=-0.19 $Y=1.66 $X2=3.795 $Y2=2.4
cc_170 VPB N_TE_B_c_675_n 0.00427266f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=1.32
cc_171 VPB N_A_M1026_g 0.0230335f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_172 VPB N_A_M1032_g 0.0249374f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_173 VPB N_A_28_368#_c_887_n 0.0501872f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_174 VPB N_A_28_368#_c_888_n 0.0025134f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_28_368#_c_889_n 0.00929469f $X=-0.19 $Y=1.66 $X2=1.91 $Y2=1.65
cc_176 VPB N_A_28_368#_c_890_n 0.00262732f $X=-0.19 $Y=1.66 $X2=2.31 $Y2=0.74
cc_177 VPB N_A_28_368#_c_891_n 0.00240659f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_28_368#_c_892_n 0.00445308f $X=-0.19 $Y=1.66 $X2=2.81 $Y2=0.74
cc_179 VPB N_A_28_368#_c_893_n 0.00171072f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=0.74
cc_180 VPB N_A_28_368#_c_894_n 0.00123754f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=0.74
cc_181 VPB N_A_28_368#_c_895_n 0.00196551f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_28_368#_c_896_n 0.0023101f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=1.485
cc_183 VPB N_A_28_368#_c_897_n 0.0023101f $X=-0.19 $Y=1.66 $X2=3.87 $Y2=1.565
cc_184 VPB N_A_28_368#_c_898_n 0.0023101f $X=-0.19 $Y=1.66 $X2=3.955 $Y2=2.05
cc_185 VPB N_A_28_368#_c_899_n 0.0187412f $X=-0.19 $Y=1.66 $X2=9.665 $Y2=2.305
cc_186 VPB N_Z_c_1030_n 0.00236883f $X=-0.19 $Y=1.66 $X2=1.81 $Y2=1.32
cc_187 VPB N_Z_c_1031_n 0.00219429f $X=-0.19 $Y=1.66 $X2=2.36 $Y2=1.65
cc_188 VPB N_Z_c_1032_n 0.00249468f $X=-0.19 $Y=1.66 $X2=2.81 $Y2=0.74
cc_189 VPB N_Z_c_1033_n 0.00256624f $X=-0.19 $Y=1.66 $X2=3.31 $Y2=2.4
cc_190 VPB N_Z_c_1034_n 5.31124e-19 $X=-0.19 $Y=1.66 $X2=3.81 $Y2=1.32
cc_191 VPB N_Z_c_1035_n 0.00236205f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_Z_c_1036_n 0.00224287f $X=-0.19 $Y=1.66 $X2=1.14 $Y2=1.485
cc_193 VPB Z 0.00153546f $X=-0.19 $Y=1.66 $X2=3.655 $Y2=1.565
cc_194 VPB N_VPWR_c_1153_n 0.00858545f $X=-0.19 $Y=1.66 $X2=0.96 $Y2=2.4
cc_195 VPB N_VPWR_c_1154_n 0.0083004f $X=-0.19 $Y=1.66 $X2=1.38 $Y2=0.74
cc_196 VPB N_VPWR_c_1155_n 0.00899828f $X=-0.19 $Y=1.66 $X2=1.41 $Y2=2.4
cc_197 VPB N_VPWR_c_1156_n 0.0188241f $X=-0.19 $Y=1.66 $X2=1.81 $Y2=1.32
cc_198 VPB N_VPWR_c_1157_n 0.00802001f $X=-0.19 $Y=1.66 $X2=1.91 $Y2=1.65
cc_199 VPB N_VPWR_c_1158_n 0.00556529f $X=-0.19 $Y=1.66 $X2=2.31 $Y2=1.32
cc_200 VPB N_VPWR_c_1159_n 0.0119967f $X=-0.19 $Y=1.66 $X2=2.31 $Y2=0.74
cc_201 VPB N_VPWR_c_1160_n 0.0442765f $X=-0.19 $Y=1.66 $X2=2.36 $Y2=1.65
cc_202 VPB N_VPWR_c_1161_n 0.101612f $X=-0.19 $Y=1.66 $X2=2.81 $Y2=2.4
cc_203 VPB N_VPWR_c_1162_n 0.0186948f $X=-0.19 $Y=1.66 $X2=3.31 $Y2=2.4
cc_204 VPB N_VPWR_c_1163_n 0.0186948f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1164_n 0.0417371f $X=-0.19 $Y=1.66 $X2=3.81 $Y2=1.32
cc_206 VPB N_VPWR_c_1165_n 0.0173363f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1166_n 0.00631813f $X=-0.19 $Y=1.66 $X2=4.04 $Y2=2.135
cc_208 VPB N_VPWR_c_1167_n 0.00632182f $X=-0.19 $Y=1.66 $X2=9.805 $Y2=1.89
cc_209 VPB N_VPWR_c_1168_n 0.00632182f $X=-0.19 $Y=1.66 $X2=9.83 $Y2=1.985
cc_210 VPB N_VPWR_c_1169_n 0.00631222f $X=-0.19 $Y=1.66 $X2=9.83 $Y2=2.815
cc_211 VPB N_VPWR_c_1170_n 0.0061274f $X=-0.19 $Y=1.66 $X2=9.805 $Y2=0.505
cc_212 VPB N_VPWR_c_1152_n 0.110087f $X=-0.19 $Y=1.66 $X2=9.93 $Y2=0.925
cc_213 N_A_84_48#_c_243_n N_A_833_48#_M1028_s 0.0237719f $X=9.665 $Y=2.305 $X2=0
+ $Y2=0
cc_214 N_A_84_48#_M1036_g N_A_833_48#_c_490_n 0.00835898f $X=3.81 $Y=0.74 $X2=0
+ $Y2=0
cc_215 N_A_84_48#_c_233_n N_A_833_48#_c_492_n 0.00835898f $X=3.81 $Y=1.485 $X2=0
+ $Y2=0
cc_216 N_A_84_48#_c_243_n N_A_833_48#_c_525_n 0.00891814f $X=9.665 $Y=2.305
+ $X2=0 $Y2=0
cc_217 N_A_84_48#_c_243_n N_A_833_48#_c_521_n 0.0673532f $X=9.665 $Y=2.305 $X2=0
+ $Y2=0
cc_218 N_A_84_48#_c_253_p N_A_833_48#_c_521_n 0.00425919f $X=9.83 $Y=1.985 $X2=0
+ $Y2=0
cc_219 N_A_84_48#_c_246_n N_A_833_48#_c_521_n 0.00254866f $X=9.945 $Y=1.805
+ $X2=0 $Y2=0
cc_220 N_A_84_48#_M1035_g N_TE_B_c_676_n 0.0170175f $X=3.795 $Y=2.4 $X2=-0.19
+ $Y2=-0.245
cc_221 N_A_84_48#_c_256_p N_TE_B_c_676_n 0.0172321f $X=7.585 $Y=2.135 $X2=-0.19
+ $Y2=-0.245
cc_222 N_A_84_48#_c_256_p N_TE_B_c_655_n 0.00575192f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_223 N_A_84_48#_c_230_n N_TE_B_c_656_n 0.00106842f $X=3.87 $Y=1.565 $X2=0
+ $Y2=0
cc_224 N_A_84_48#_c_242_n N_TE_B_c_656_n 0.00889779f $X=3.955 $Y=2.05 $X2=0
+ $Y2=0
cc_225 N_A_84_48#_c_233_n N_TE_B_c_656_n 0.0170175f $X=3.81 $Y=1.485 $X2=0 $Y2=0
cc_226 N_A_84_48#_c_256_p N_TE_B_c_679_n 0.0139722f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_227 N_A_84_48#_c_256_p N_TE_B_c_657_n 0.00181991f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_228 N_A_84_48#_c_256_p N_TE_B_c_681_n 0.0139992f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_229 N_A_84_48#_c_256_p N_TE_B_c_658_n 0.00382113f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_230 N_A_84_48#_c_256_p N_TE_B_c_683_n 0.0139971f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_231 N_A_84_48#_c_256_p N_TE_B_c_659_n 0.00181018f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_232 N_A_84_48#_c_256_p N_TE_B_c_685_n 0.0139992f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_233 N_A_84_48#_c_256_p N_TE_B_c_660_n 0.00382012f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_234 N_A_84_48#_c_256_p N_TE_B_c_687_n 0.0139469f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_235 N_A_84_48#_c_256_p N_TE_B_c_661_n 0.00181018f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_236 N_A_84_48#_c_256_p N_TE_B_c_689_n 0.0145205f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_237 N_A_84_48#_c_272_p N_TE_B_c_689_n 0.00373646f $X=7.67 $Y=2.135 $X2=0
+ $Y2=0
cc_238 N_A_84_48#_c_256_p N_TE_B_c_662_n 0.00327121f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_239 N_A_84_48#_c_272_p N_TE_B_c_662_n 0.00376009f $X=7.67 $Y=2.135 $X2=0
+ $Y2=0
cc_240 N_A_84_48#_c_243_n N_TE_B_c_691_n 0.0169228f $X=9.665 $Y=2.305 $X2=0
+ $Y2=0
cc_241 N_A_84_48#_c_243_n N_TE_B_c_694_n 0.020923f $X=9.665 $Y=2.305 $X2=0 $Y2=0
cc_242 N_A_84_48#_c_253_p N_TE_B_c_694_n 0.00128021f $X=9.83 $Y=1.985 $X2=0
+ $Y2=0
cc_243 N_A_84_48#_c_244_n N_TE_B_c_694_n 8.43479e-19 $X=9.83 $Y=2.815 $X2=0
+ $Y2=0
cc_244 N_A_84_48#_c_243_n TE_B 0.0103192f $X=9.665 $Y=2.305 $X2=0 $Y2=0
cc_245 N_A_84_48#_c_243_n N_TE_B_c_674_n 0.00121335f $X=9.665 $Y=2.305 $X2=0
+ $Y2=0
cc_246 N_A_84_48#_c_243_n N_TE_B_c_675_n 0.0012261f $X=9.665 $Y=2.305 $X2=0
+ $Y2=0
cc_247 N_A_84_48#_c_246_n N_TE_B_c_675_n 6.8077e-19 $X=9.945 $Y=1.805 $X2=0
+ $Y2=0
cc_248 N_A_84_48#_c_243_n N_A_M1026_g 0.0174522f $X=9.665 $Y=2.305 $X2=0 $Y2=0
cc_249 N_A_84_48#_c_253_p N_A_M1026_g 0.00673876f $X=9.83 $Y=1.985 $X2=0 $Y2=0
cc_250 N_A_84_48#_c_244_n N_A_M1026_g 0.00872778f $X=9.83 $Y=2.815 $X2=0 $Y2=0
cc_251 N_A_84_48#_c_246_n N_A_M1026_g 0.00532279f $X=9.945 $Y=1.805 $X2=0 $Y2=0
cc_252 N_A_84_48#_c_287_p N_A_M1026_g 4.64231e-19 $X=9.805 $Y=2.305 $X2=0 $Y2=0
cc_253 N_A_84_48#_c_288_p N_A_c_838_n 0.00208866f $X=9.805 $Y=0.84 $X2=0 $Y2=0
cc_254 N_A_84_48#_c_231_n N_A_c_838_n 0.00591333f $X=9.845 $Y=0.505 $X2=0 $Y2=0
cc_255 N_A_84_48#_c_244_n N_A_M1032_g 2.69566e-19 $X=9.83 $Y=2.815 $X2=0 $Y2=0
cc_256 N_A_84_48#_c_245_n N_A_M1032_g 0.0218164f $X=10.145 $Y=1.805 $X2=0 $Y2=0
cc_257 N_A_84_48#_c_231_n N_A_c_840_n 3.45303e-19 $X=9.845 $Y=0.505 $X2=0 $Y2=0
cc_258 N_A_84_48#_c_293_p N_A_c_840_n 0.0152487f $X=10.145 $Y=0.925 $X2=0 $Y2=0
cc_259 N_A_84_48#_c_232_n N_A_c_840_n 0.0057552f $X=10.23 $Y=1.72 $X2=0 $Y2=0
cc_260 N_A_84_48#_c_243_n A 4.25182e-19 $X=9.665 $Y=2.305 $X2=0 $Y2=0
cc_261 N_A_84_48#_c_288_p A 0.0190643f $X=9.805 $Y=0.84 $X2=0 $Y2=0
cc_262 N_A_84_48#_c_245_n A 0.00213835f $X=10.145 $Y=1.805 $X2=0 $Y2=0
cc_263 N_A_84_48#_c_246_n A 0.023783f $X=9.945 $Y=1.805 $X2=0 $Y2=0
cc_264 N_A_84_48#_c_232_n A 0.0279669f $X=10.23 $Y=1.72 $X2=0 $Y2=0
cc_265 N_A_84_48#_c_288_p N_A_c_842_n 7.03839e-19 $X=9.805 $Y=0.84 $X2=0 $Y2=0
cc_266 N_A_84_48#_c_246_n N_A_c_842_n 7.11382e-19 $X=9.945 $Y=1.805 $X2=0 $Y2=0
cc_267 N_A_84_48#_c_232_n N_A_c_842_n 0.0174675f $X=10.23 $Y=1.72 $X2=0 $Y2=0
cc_268 N_A_84_48#_c_242_n N_A_28_368#_M1035_s 0.00236618f $X=3.955 $Y=2.05 $X2=0
+ $Y2=0
cc_269 N_A_84_48#_c_256_p N_A_28_368#_M1035_s 0.00351257f $X=7.585 $Y=2.135
+ $X2=0 $Y2=0
cc_270 N_A_84_48#_c_305_p N_A_28_368#_M1035_s 0.00107343f $X=4.04 $Y=2.135 $X2=0
+ $Y2=0
cc_271 N_A_84_48#_c_256_p N_A_28_368#_M1010_d 0.00425773f $X=7.585 $Y=2.135
+ $X2=0 $Y2=0
cc_272 N_A_84_48#_c_256_p N_A_28_368#_M1016_d 0.00427366f $X=7.585 $Y=2.135
+ $X2=0 $Y2=0
cc_273 N_A_84_48#_c_256_p N_A_28_368#_M1018_d 0.00427366f $X=7.585 $Y=2.135
+ $X2=0 $Y2=0
cc_274 N_A_84_48#_c_243_n N_A_28_368#_M1022_d 0.00541402f $X=9.665 $Y=2.305
+ $X2=0 $Y2=0
cc_275 N_A_84_48#_M1001_g N_A_28_368#_c_887_n 0.00146508f $X=0.51 $Y=2.4 $X2=0
+ $Y2=0
cc_276 N_A_84_48#_M1001_g N_A_28_368#_c_888_n 0.0142242f $X=0.51 $Y=2.4 $X2=0
+ $Y2=0
cc_277 N_A_84_48#_M1002_g N_A_28_368#_c_888_n 0.0140221f $X=0.96 $Y=2.4 $X2=0
+ $Y2=0
cc_278 N_A_84_48#_M1005_g N_A_28_368#_c_910_n 0.0110737f $X=1.41 $Y=2.4 $X2=0
+ $Y2=0
cc_279 N_A_84_48#_M1006_g N_A_28_368#_c_910_n 5.44871e-19 $X=1.91 $Y=2.4 $X2=0
+ $Y2=0
cc_280 N_A_84_48#_M1005_g N_A_28_368#_c_890_n 0.0119307f $X=1.41 $Y=2.4 $X2=0
+ $Y2=0
cc_281 N_A_84_48#_M1006_g N_A_28_368#_c_890_n 0.0143183f $X=1.91 $Y=2.4 $X2=0
+ $Y2=0
cc_282 N_A_84_48#_M1008_g N_A_28_368#_c_891_n 0.0140221f $X=2.36 $Y=2.4 $X2=0
+ $Y2=0
cc_283 N_A_84_48#_M1012_g N_A_28_368#_c_891_n 0.0142213f $X=2.81 $Y=2.4 $X2=0
+ $Y2=0
cc_284 N_A_84_48#_M1014_g N_A_28_368#_c_892_n 0.0144328f $X=3.31 $Y=2.4 $X2=0
+ $Y2=0
cc_285 N_A_84_48#_M1035_g N_A_28_368#_c_892_n 0.0144843f $X=3.795 $Y=2.4 $X2=0
+ $Y2=0
cc_286 N_A_84_48#_M1035_g N_A_28_368#_c_918_n 0.00194303f $X=3.795 $Y=2.4 $X2=0
+ $Y2=0
cc_287 N_A_84_48#_c_256_p N_A_28_368#_c_918_n 0.00815076f $X=7.585 $Y=2.135
+ $X2=0 $Y2=0
cc_288 N_A_84_48#_c_305_p N_A_28_368#_c_918_n 0.0100237f $X=4.04 $Y=2.135 $X2=0
+ $Y2=0
cc_289 N_A_84_48#_M1014_g N_A_28_368#_c_921_n 5.36803e-19 $X=3.31 $Y=2.4 $X2=0
+ $Y2=0
cc_290 N_A_84_48#_M1035_g N_A_28_368#_c_921_n 0.00489895f $X=3.795 $Y=2.4 $X2=0
+ $Y2=0
cc_291 N_A_84_48#_c_256_p N_A_28_368#_c_923_n 0.0388605f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_292 N_A_84_48#_c_256_p N_A_28_368#_c_924_n 0.0388605f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_293 N_A_84_48#_c_256_p N_A_28_368#_c_925_n 0.0388943f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_294 N_A_84_48#_c_256_p N_A_28_368#_c_926_n 0.0136015f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_295 N_A_84_48#_c_243_n N_A_28_368#_c_926_n 0.0101671f $X=9.665 $Y=2.305 $X2=0
+ $Y2=0
cc_296 N_A_84_48#_c_272_p N_A_28_368#_c_926_n 0.0113151f $X=7.67 $Y=2.135 $X2=0
+ $Y2=0
cc_297 N_A_84_48#_M1005_g N_A_28_368#_c_893_n 0.00194226f $X=1.41 $Y=2.4 $X2=0
+ $Y2=0
cc_298 N_A_84_48#_c_256_p N_A_28_368#_c_896_n 0.0169819f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_299 N_A_84_48#_c_256_p N_A_28_368#_c_897_n 0.0169819f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_300 N_A_84_48#_c_256_p N_A_28_368#_c_898_n 0.0168295f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_301 N_A_84_48#_c_243_n N_A_28_368#_c_899_n 0.0211182f $X=9.665 $Y=2.305 $X2=0
+ $Y2=0
cc_302 N_A_84_48#_M1001_g N_Z_c_1038_n 0.0108799f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_303 N_A_84_48#_M1002_g N_Z_c_1038_n 0.0103925f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_304 N_A_84_48#_M1005_g N_Z_c_1038_n 6.52534e-19 $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_305 N_A_84_48#_M1013_g N_Z_c_1023_n 0.0108901f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_306 N_A_84_48#_M1019_g N_Z_c_1023_n 0.00906272f $X=1.38 $Y=0.74 $X2=0 $Y2=0
cc_307 N_A_84_48#_c_342_p N_Z_c_1023_n 0.0291873f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_308 N_A_84_48#_c_233_n N_Z_c_1023_n 0.00299956f $X=3.81 $Y=1.485 $X2=0 $Y2=0
cc_309 N_A_84_48#_M1002_g N_Z_c_1030_n 0.0149064f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_310 N_A_84_48#_M1005_g N_Z_c_1030_n 0.0145117f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_311 N_A_84_48#_c_342_p N_Z_c_1030_n 0.0356865f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_312 N_A_84_48#_c_233_n N_Z_c_1030_n 0.00207695f $X=3.81 $Y=1.485 $X2=0 $Y2=0
cc_313 N_A_84_48#_M1013_g N_Z_c_1049_n 5.43234e-19 $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_314 N_A_84_48#_M1019_g N_Z_c_1049_n 0.00600998f $X=1.38 $Y=0.74 $X2=0 $Y2=0
cc_315 N_A_84_48#_M1027_g N_Z_c_1049_n 0.00618702f $X=1.81 $Y=0.74 $X2=0 $Y2=0
cc_316 N_A_84_48#_M1030_g N_Z_c_1049_n 4.62714e-19 $X=2.31 $Y=0.74 $X2=0 $Y2=0
cc_317 N_A_84_48#_M1006_g N_Z_c_1053_n 0.0104648f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_318 N_A_84_48#_M1008_g N_Z_c_1053_n 6.14153e-19 $X=2.36 $Y=2.4 $X2=0 $Y2=0
cc_319 N_A_84_48#_M1027_g N_Z_c_1024_n 0.00930697f $X=1.81 $Y=0.74 $X2=0 $Y2=0
cc_320 N_A_84_48#_M1030_g N_Z_c_1024_n 0.0128277f $X=2.31 $Y=0.74 $X2=0 $Y2=0
cc_321 N_A_84_48#_c_342_p N_Z_c_1024_n 0.0492574f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_322 N_A_84_48#_c_233_n N_Z_c_1024_n 0.00426458f $X=3.81 $Y=1.485 $X2=0 $Y2=0
cc_323 N_A_84_48#_M1006_g N_Z_c_1031_n 0.012931f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_324 N_A_84_48#_M1008_g N_Z_c_1031_n 0.012931f $X=2.36 $Y=2.4 $X2=0 $Y2=0
cc_325 N_A_84_48#_c_342_p N_Z_c_1031_n 0.0416512f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_326 N_A_84_48#_c_233_n N_Z_c_1031_n 0.00215575f $X=3.81 $Y=1.485 $X2=0 $Y2=0
cc_327 N_A_84_48#_M1006_g N_Z_c_1063_n 6.14153e-19 $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_328 N_A_84_48#_M1008_g N_Z_c_1063_n 0.0104648f $X=2.36 $Y=2.4 $X2=0 $Y2=0
cc_329 N_A_84_48#_M1012_g N_Z_c_1063_n 0.0102924f $X=2.81 $Y=2.4 $X2=0 $Y2=0
cc_330 N_A_84_48#_M1014_g N_Z_c_1063_n 5.83379e-19 $X=3.31 $Y=2.4 $X2=0 $Y2=0
cc_331 N_A_84_48#_M1031_g N_Z_c_1067_n 0.00620791f $X=2.81 $Y=0.74 $X2=0 $Y2=0
cc_332 N_A_84_48#_M1033_g N_Z_c_1067_n 4.62024e-19 $X=3.325 $Y=0.74 $X2=0 $Y2=0
cc_333 N_A_84_48#_M1012_g N_Z_c_1032_n 0.0132272f $X=2.81 $Y=2.4 $X2=0 $Y2=0
cc_334 N_A_84_48#_M1014_g N_Z_c_1032_n 0.0132272f $X=3.31 $Y=2.4 $X2=0 $Y2=0
cc_335 N_A_84_48#_c_342_p N_Z_c_1032_n 0.045409f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_336 N_A_84_48#_c_233_n N_Z_c_1032_n 0.00313888f $X=3.81 $Y=1.485 $X2=0 $Y2=0
cc_337 N_A_84_48#_M1031_g N_Z_c_1025_n 0.00938204f $X=2.81 $Y=0.74 $X2=0 $Y2=0
cc_338 N_A_84_48#_M1033_g N_Z_c_1025_n 0.0130129f $X=3.325 $Y=0.74 $X2=0 $Y2=0
cc_339 N_A_84_48#_M1036_g N_Z_c_1025_n 0.00461775f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_340 N_A_84_48#_c_342_p N_Z_c_1025_n 0.0678816f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_341 N_A_84_48#_c_230_n N_Z_c_1025_n 0.0049593f $X=3.87 $Y=1.565 $X2=0 $Y2=0
cc_342 N_A_84_48#_c_233_n N_Z_c_1025_n 0.00802702f $X=3.81 $Y=1.485 $X2=0 $Y2=0
cc_343 N_A_84_48#_M1014_g N_Z_c_1033_n 0.00110956f $X=3.31 $Y=2.4 $X2=0 $Y2=0
cc_344 N_A_84_48#_c_342_p N_Z_c_1033_n 0.0274622f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_345 N_A_84_48#_c_242_n N_Z_c_1033_n 0.00667444f $X=3.955 $Y=2.05 $X2=0 $Y2=0
cc_346 N_A_84_48#_c_233_n N_Z_c_1033_n 0.00291196f $X=3.81 $Y=1.485 $X2=0 $Y2=0
cc_347 N_A_84_48#_M1012_g N_Z_c_1083_n 5.90928e-19 $X=2.81 $Y=2.4 $X2=0 $Y2=0
cc_348 N_A_84_48#_M1014_g N_Z_c_1083_n 0.010427f $X=3.31 $Y=2.4 $X2=0 $Y2=0
cc_349 N_A_84_48#_M1036_g N_Z_c_1085_n 0.00457683f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_350 N_A_84_48#_M1001_g N_Z_c_1034_n 0.00254215f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_351 N_A_84_48#_M1002_g N_Z_c_1034_n 0.00153805f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_352 N_A_84_48#_M1019_g N_Z_c_1026_n 0.00277555f $X=1.38 $Y=0.74 $X2=0 $Y2=0
cc_353 N_A_84_48#_M1027_g N_Z_c_1026_n 0.00277555f $X=1.81 $Y=0.74 $X2=0 $Y2=0
cc_354 N_A_84_48#_c_342_p N_Z_c_1026_n 0.0271537f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_355 N_A_84_48#_c_233_n N_Z_c_1026_n 0.00248949f $X=3.81 $Y=1.485 $X2=0 $Y2=0
cc_356 N_A_84_48#_M1006_g N_Z_c_1035_n 0.00115436f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_357 N_A_84_48#_c_342_p N_Z_c_1035_n 0.0276979f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_358 N_A_84_48#_c_233_n N_Z_c_1035_n 0.00359665f $X=3.81 $Y=1.485 $X2=0 $Y2=0
cc_359 N_A_84_48#_M1008_g N_Z_c_1036_n 0.00112087f $X=2.36 $Y=2.4 $X2=0 $Y2=0
cc_360 N_A_84_48#_M1012_g N_Z_c_1036_n 0.00112087f $X=2.81 $Y=2.4 $X2=0 $Y2=0
cc_361 N_A_84_48#_c_342_p N_Z_c_1036_n 0.0275631f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_362 N_A_84_48#_c_233_n N_Z_c_1036_n 0.00209661f $X=3.81 $Y=1.485 $X2=0 $Y2=0
cc_363 N_A_84_48#_M1031_g N_Z_c_1027_n 0.00317348f $X=2.81 $Y=0.74 $X2=0 $Y2=0
cc_364 N_A_84_48#_c_342_p N_Z_c_1027_n 0.0272627f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_365 N_A_84_48#_c_233_n N_Z_c_1027_n 0.00424593f $X=3.81 $Y=1.485 $X2=0 $Y2=0
cc_366 N_A_84_48#_M1007_g Z 0.00463107f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_367 N_A_84_48#_M1013_g Z 0.00311186f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_368 N_A_84_48#_M1007_g Z 0.00883951f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_369 N_A_84_48#_M1001_g Z 0.00918156f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_370 N_A_84_48#_M1013_g Z 0.00469957f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_371 N_A_84_48#_M1002_g Z 0.00458897f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_372 N_A_84_48#_c_342_p Z 0.0227592f $X=3.49 $Y=1.485 $X2=0 $Y2=0
cc_373 N_A_84_48#_c_233_n Z 0.0320249f $X=3.81 $Y=1.485 $X2=0 $Y2=0
cc_374 N_A_84_48#_M1007_g N_Z_c_1110_n 0.00480711f $X=0.495 $Y=0.74 $X2=0 $Y2=0
cc_375 N_A_84_48#_M1013_g N_Z_c_1110_n 0.00588517f $X=0.925 $Y=0.74 $X2=0 $Y2=0
cc_376 N_A_84_48#_M1019_g N_Z_c_1110_n 5.35511e-19 $X=1.38 $Y=0.74 $X2=0 $Y2=0
cc_377 N_A_84_48#_c_256_p N_VPWR_M1009_s 0.00775066f $X=7.585 $Y=2.135 $X2=-0.19
+ $Y2=-0.245
cc_378 N_A_84_48#_c_256_p N_VPWR_M1015_s 0.00690732f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_379 N_A_84_48#_c_256_p N_VPWR_M1017_s 0.00690586f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_380 N_A_84_48#_c_256_p N_VPWR_M1021_s 0.00625322f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_381 N_A_84_48#_c_272_p N_VPWR_M1021_s 0.00748716f $X=7.67 $Y=2.135 $X2=0
+ $Y2=0
cc_382 N_A_84_48#_c_243_n N_VPWR_M1028_d 0.00647629f $X=9.665 $Y=2.305 $X2=0
+ $Y2=0
cc_383 N_A_84_48#_c_245_n N_VPWR_M1032_s 0.00349386f $X=10.145 $Y=1.805 $X2=0
+ $Y2=0
cc_384 N_A_84_48#_c_243_n N_VPWR_c_1158_n 0.0189268f $X=9.665 $Y=2.305 $X2=0
+ $Y2=0
cc_385 N_A_84_48#_c_244_n N_VPWR_c_1158_n 0.0161582f $X=9.83 $Y=2.815 $X2=0
+ $Y2=0
cc_386 N_A_84_48#_c_244_n N_VPWR_c_1160_n 0.0229093f $X=9.83 $Y=2.815 $X2=0
+ $Y2=0
cc_387 N_A_84_48#_c_245_n N_VPWR_c_1160_n 0.0123212f $X=10.145 $Y=1.805 $X2=0
+ $Y2=0
cc_388 N_A_84_48#_M1001_g N_VPWR_c_1161_n 0.00333926f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_389 N_A_84_48#_M1002_g N_VPWR_c_1161_n 0.00333926f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_390 N_A_84_48#_M1005_g N_VPWR_c_1161_n 0.00333896f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_391 N_A_84_48#_M1006_g N_VPWR_c_1161_n 0.00333926f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_392 N_A_84_48#_M1008_g N_VPWR_c_1161_n 0.00333926f $X=2.36 $Y=2.4 $X2=0 $Y2=0
cc_393 N_A_84_48#_M1012_g N_VPWR_c_1161_n 0.00333926f $X=2.81 $Y=2.4 $X2=0 $Y2=0
cc_394 N_A_84_48#_M1014_g N_VPWR_c_1161_n 0.00333926f $X=3.31 $Y=2.4 $X2=0 $Y2=0
cc_395 N_A_84_48#_M1035_g N_VPWR_c_1161_n 0.00333911f $X=3.795 $Y=2.4 $X2=0
+ $Y2=0
cc_396 N_A_84_48#_c_244_n N_VPWR_c_1165_n 0.0123179f $X=9.83 $Y=2.815 $X2=0
+ $Y2=0
cc_397 N_A_84_48#_M1001_g N_VPWR_c_1152_n 0.00426447f $X=0.51 $Y=2.4 $X2=0 $Y2=0
cc_398 N_A_84_48#_M1002_g N_VPWR_c_1152_n 0.00422687f $X=0.96 $Y=2.4 $X2=0 $Y2=0
cc_399 N_A_84_48#_M1005_g N_VPWR_c_1152_n 0.00423173f $X=1.41 $Y=2.4 $X2=0 $Y2=0
cc_400 N_A_84_48#_M1006_g N_VPWR_c_1152_n 0.00423176f $X=1.91 $Y=2.4 $X2=0 $Y2=0
cc_401 N_A_84_48#_M1008_g N_VPWR_c_1152_n 0.00422687f $X=2.36 $Y=2.4 $X2=0 $Y2=0
cc_402 N_A_84_48#_M1012_g N_VPWR_c_1152_n 0.00423176f $X=2.81 $Y=2.4 $X2=0 $Y2=0
cc_403 N_A_84_48#_M1014_g N_VPWR_c_1152_n 0.00423522f $X=3.31 $Y=2.4 $X2=0 $Y2=0
cc_404 N_A_84_48#_M1035_g N_VPWR_c_1152_n 0.00423285f $X=3.795 $Y=2.4 $X2=0
+ $Y2=0
cc_405 N_A_84_48#_c_244_n N_VPWR_c_1152_n 0.0101276f $X=9.83 $Y=2.815 $X2=0
+ $Y2=0
cc_406 N_A_84_48#_M1007_g N_A_27_74#_c_1281_n 0.00159289f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_407 N_A_84_48#_M1007_g N_A_27_74#_c_1282_n 0.0132617f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_408 N_A_84_48#_M1013_g N_A_27_74#_c_1282_n 0.0108851f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_409 N_A_84_48#_M1019_g N_A_27_74#_c_1306_n 0.00394726f $X=1.38 $Y=0.74 $X2=0
+ $Y2=0
cc_410 N_A_84_48#_M1019_g N_A_27_74#_c_1284_n 0.0108851f $X=1.38 $Y=0.74 $X2=0
+ $Y2=0
cc_411 N_A_84_48#_M1027_g N_A_27_74#_c_1284_n 0.0111293f $X=1.81 $Y=0.74 $X2=0
+ $Y2=0
cc_412 N_A_84_48#_M1030_g N_A_27_74#_c_1309_n 0.0061935f $X=2.31 $Y=0.74 $X2=0
+ $Y2=0
cc_413 N_A_84_48#_M1031_g N_A_27_74#_c_1309_n 4.62714e-19 $X=2.81 $Y=0.74 $X2=0
+ $Y2=0
cc_414 N_A_84_48#_M1030_g N_A_27_74#_c_1285_n 0.00822804f $X=2.31 $Y=0.74 $X2=0
+ $Y2=0
cc_415 N_A_84_48#_M1031_g N_A_27_74#_c_1285_n 0.0115976f $X=2.81 $Y=0.74 $X2=0
+ $Y2=0
cc_416 N_A_84_48#_M1033_g N_A_27_74#_c_1313_n 0.00542481f $X=3.325 $Y=0.74 $X2=0
+ $Y2=0
cc_417 N_A_84_48#_M1036_g N_A_27_74#_c_1313_n 7.18008e-19 $X=3.81 $Y=0.74 $X2=0
+ $Y2=0
cc_418 N_A_84_48#_M1033_g N_A_27_74#_c_1286_n 0.00879688f $X=3.325 $Y=0.74 $X2=0
+ $Y2=0
cc_419 N_A_84_48#_M1036_g N_A_27_74#_c_1286_n 0.0123192f $X=3.81 $Y=0.74 $X2=0
+ $Y2=0
cc_420 N_A_84_48#_M1036_g N_A_27_74#_c_1287_n 4.60332e-19 $X=3.81 $Y=0.74 $X2=0
+ $Y2=0
cc_421 N_A_84_48#_M1036_g N_A_27_74#_c_1289_n 0.00514561f $X=3.81 $Y=0.74 $X2=0
+ $Y2=0
cc_422 N_A_84_48#_c_230_n N_A_27_74#_c_1289_n 0.00936976f $X=3.87 $Y=1.565 $X2=0
+ $Y2=0
cc_423 N_A_84_48#_c_256_p N_A_27_74#_c_1291_n 0.0140299f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_424 N_A_84_48#_c_256_p N_A_27_74#_c_1293_n 0.0154654f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_425 N_A_84_48#_c_256_p N_A_27_74#_c_1295_n 0.0233169f $X=7.585 $Y=2.135 $X2=0
+ $Y2=0
cc_426 N_A_84_48#_M1030_g N_A_27_74#_c_1298_n 0.00294698f $X=2.31 $Y=0.74 $X2=0
+ $Y2=0
cc_427 N_A_84_48#_M1033_g N_A_27_74#_c_1299_n 0.00270885f $X=3.325 $Y=0.74 $X2=0
+ $Y2=0
cc_428 N_A_84_48#_c_256_p N_A_27_74#_c_1300_n 0.00981245f $X=7.585 $Y=2.135
+ $X2=0 $Y2=0
cc_429 N_A_84_48#_c_256_p N_A_27_74#_c_1301_n 0.00746164f $X=7.585 $Y=2.135
+ $X2=0 $Y2=0
cc_430 N_A_84_48#_c_256_p N_A_27_74#_c_1302_n 0.00813622f $X=7.585 $Y=2.135
+ $X2=0 $Y2=0
cc_431 N_A_84_48#_c_293_p N_VGND_M1023_s 0.00916777f $X=10.145 $Y=0.925 $X2=0
+ $Y2=0
cc_432 N_A_84_48#_c_232_n N_VGND_M1023_s 0.0037774f $X=10.23 $Y=1.72 $X2=0 $Y2=0
cc_433 N_A_84_48#_c_231_n N_VGND_c_1450_n 0.0181878f $X=9.845 $Y=0.505 $X2=0
+ $Y2=0
cc_434 N_A_84_48#_c_231_n N_VGND_c_1452_n 0.0104513f $X=9.845 $Y=0.505 $X2=0
+ $Y2=0
cc_435 N_A_84_48#_c_293_p N_VGND_c_1452_n 0.00936242f $X=10.145 $Y=0.925 $X2=0
+ $Y2=0
cc_436 N_A_84_48#_M1007_g N_VGND_c_1453_n 0.00278271f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_437 N_A_84_48#_M1013_g N_VGND_c_1453_n 0.00278271f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_438 N_A_84_48#_M1019_g N_VGND_c_1453_n 0.00278271f $X=1.38 $Y=0.74 $X2=0
+ $Y2=0
cc_439 N_A_84_48#_M1027_g N_VGND_c_1453_n 0.00278271f $X=1.81 $Y=0.74 $X2=0
+ $Y2=0
cc_440 N_A_84_48#_M1030_g N_VGND_c_1453_n 0.00278247f $X=2.31 $Y=0.74 $X2=0
+ $Y2=0
cc_441 N_A_84_48#_M1031_g N_VGND_c_1453_n 0.00278271f $X=2.81 $Y=0.74 $X2=0
+ $Y2=0
cc_442 N_A_84_48#_M1033_g N_VGND_c_1453_n 0.00278262f $X=3.325 $Y=0.74 $X2=0
+ $Y2=0
cc_443 N_A_84_48#_M1036_g N_VGND_c_1453_n 0.00278271f $X=3.81 $Y=0.74 $X2=0
+ $Y2=0
cc_444 N_A_84_48#_c_231_n N_VGND_c_1461_n 0.0114427f $X=9.845 $Y=0.505 $X2=0
+ $Y2=0
cc_445 N_A_84_48#_M1007_g N_VGND_c_1464_n 0.00357086f $X=0.495 $Y=0.74 $X2=0
+ $Y2=0
cc_446 N_A_84_48#_M1013_g N_VGND_c_1464_n 0.00353674f $X=0.925 $Y=0.74 $X2=0
+ $Y2=0
cc_447 N_A_84_48#_M1019_g N_VGND_c_1464_n 0.00353674f $X=1.38 $Y=0.74 $X2=0
+ $Y2=0
cc_448 N_A_84_48#_M1027_g N_VGND_c_1464_n 0.00354087f $X=1.81 $Y=0.74 $X2=0
+ $Y2=0
cc_449 N_A_84_48#_M1030_g N_VGND_c_1464_n 0.00354743f $X=2.31 $Y=0.74 $X2=0
+ $Y2=0
cc_450 N_A_84_48#_M1031_g N_VGND_c_1464_n 0.00354875f $X=2.81 $Y=0.74 $X2=0
+ $Y2=0
cc_451 N_A_84_48#_M1033_g N_VGND_c_1464_n 0.0035474f $X=3.325 $Y=0.74 $X2=0
+ $Y2=0
cc_452 N_A_84_48#_M1036_g N_VGND_c_1464_n 0.0035405f $X=3.81 $Y=0.74 $X2=0 $Y2=0
cc_453 N_A_84_48#_c_231_n N_VGND_c_1464_n 0.00909435f $X=9.845 $Y=0.505 $X2=0
+ $Y2=0
cc_454 N_A_84_48#_c_293_p N_VGND_c_1464_n 0.00616274f $X=10.145 $Y=0.925 $X2=0
+ $Y2=0
cc_455 N_A_833_48#_c_491_n N_TE_B_c_655_n 0.0115273f $X=4.595 $Y=1.26 $X2=0
+ $Y2=0
cc_456 N_A_833_48#_c_492_n N_TE_B_c_656_n 0.0115273f $X=4.315 $Y=1.26 $X2=0
+ $Y2=0
cc_457 N_A_833_48#_c_494_n N_TE_B_c_657_n 0.0115273f $X=5.025 $Y=1.26 $X2=0
+ $Y2=0
cc_458 N_A_833_48#_c_496_n N_TE_B_c_658_n 0.0115273f $X=5.455 $Y=1.26 $X2=0
+ $Y2=0
cc_459 N_A_833_48#_c_498_n N_TE_B_c_659_n 0.0115273f $X=5.885 $Y=1.26 $X2=0
+ $Y2=0
cc_460 N_A_833_48#_c_500_n N_TE_B_c_660_n 0.0115273f $X=6.315 $Y=1.26 $X2=0
+ $Y2=0
cc_461 N_A_833_48#_c_502_n N_TE_B_c_661_n 0.0115273f $X=6.745 $Y=1.26 $X2=0
+ $Y2=0
cc_462 N_A_833_48#_c_525_n N_TE_B_c_689_n 0.00112842f $X=8.095 $Y=1.925 $X2=0
+ $Y2=0
cc_463 N_A_833_48#_c_504_n N_TE_B_c_662_n 0.0115273f $X=7.175 $Y=1.26 $X2=0
+ $Y2=0
cc_464 N_A_833_48#_c_516_n N_TE_B_c_691_n 0.00126213f $X=8.01 $Y=1.8 $X2=0 $Y2=0
cc_465 N_A_833_48#_c_525_n N_TE_B_c_691_n 0.01282f $X=8.095 $Y=1.925 $X2=0 $Y2=0
cc_466 N_A_833_48#_c_506_n N_TE_B_c_664_n 0.00317119f $X=7.72 $Y=1.26 $X2=0
+ $Y2=0
cc_467 N_A_833_48#_c_516_n N_TE_B_c_664_n 0.00462536f $X=8.01 $Y=1.8 $X2=0 $Y2=0
cc_468 N_A_833_48#_c_518_n N_TE_B_c_664_n 0.00756727f $X=8.565 $Y=0.505 $X2=0
+ $Y2=0
cc_469 N_A_833_48#_c_519_n N_TE_B_c_664_n 0.00456187f $X=8.985 $Y=0.515 $X2=0
+ $Y2=0
cc_470 N_A_833_48#_c_521_n N_TE_B_c_694_n 0.0119787f $X=8.77 $Y=1.965 $X2=0
+ $Y2=0
cc_471 N_A_833_48#_c_518_n N_TE_B_c_665_n 0.00516259f $X=8.565 $Y=0.505 $X2=0
+ $Y2=0
cc_472 N_A_833_48#_c_519_n N_TE_B_c_665_n 0.00794536f $X=8.985 $Y=0.515 $X2=0
+ $Y2=0
cc_473 N_A_833_48#_c_508_n N_TE_B_c_666_n 0.0115273f $X=4.67 $Y=1.26 $X2=0 $Y2=0
cc_474 N_A_833_48#_c_509_n N_TE_B_c_667_n 0.0115273f $X=5.1 $Y=1.26 $X2=0 $Y2=0
cc_475 N_A_833_48#_c_510_n N_TE_B_c_668_n 0.0115273f $X=5.53 $Y=1.26 $X2=0 $Y2=0
cc_476 N_A_833_48#_c_511_n N_TE_B_c_669_n 0.0115273f $X=5.96 $Y=1.26 $X2=0 $Y2=0
cc_477 N_A_833_48#_c_512_n N_TE_B_c_670_n 0.0115273f $X=6.39 $Y=1.26 $X2=0 $Y2=0
cc_478 N_A_833_48#_c_513_n N_TE_B_c_671_n 0.0115273f $X=6.82 $Y=1.26 $X2=0 $Y2=0
cc_479 N_A_833_48#_c_514_n N_TE_B_c_672_n 0.0115273f $X=7.25 $Y=1.26 $X2=0 $Y2=0
cc_480 N_A_833_48#_c_516_n N_TE_B_c_672_n 0.00836196f $X=8.01 $Y=1.8 $X2=0 $Y2=0
cc_481 N_A_833_48#_c_516_n TE_B 0.0295862f $X=8.01 $Y=1.8 $X2=0 $Y2=0
cc_482 N_A_833_48#_c_518_n TE_B 9.40747e-19 $X=8.565 $Y=0.505 $X2=0 $Y2=0
cc_483 N_A_833_48#_c_519_n TE_B 0.0751834f $X=8.985 $Y=0.515 $X2=0 $Y2=0
cc_484 N_A_833_48#_c_521_n TE_B 0.0454738f $X=8.77 $Y=1.965 $X2=0 $Y2=0
cc_485 N_A_833_48#_c_516_n N_TE_B_c_674_n 0.0121043f $X=8.01 $Y=1.8 $X2=0 $Y2=0
cc_486 N_A_833_48#_c_519_n N_TE_B_c_674_n 0.00437509f $X=8.985 $Y=0.515 $X2=0
+ $Y2=0
cc_487 N_A_833_48#_c_521_n N_TE_B_c_674_n 0.0273001f $X=8.77 $Y=1.965 $X2=0
+ $Y2=0
cc_488 N_A_833_48#_c_521_n N_A_M1026_g 7.4873e-19 $X=8.77 $Y=1.965 $X2=0 $Y2=0
cc_489 N_A_833_48#_c_525_n N_A_28_368#_M1022_d 7.54356e-19 $X=8.095 $Y=1.925
+ $X2=0 $Y2=0
cc_490 N_A_833_48#_c_521_n N_A_28_368#_M1022_d 0.00223631f $X=8.77 $Y=1.965
+ $X2=0 $Y2=0
cc_491 N_A_833_48#_c_490_n N_A_27_74#_c_1286_n 9.48753e-19 $X=4.24 $Y=1.185
+ $X2=0 $Y2=0
cc_492 N_A_833_48#_c_490_n N_A_27_74#_c_1287_n 9.29165e-19 $X=4.24 $Y=1.185
+ $X2=0 $Y2=0
cc_493 N_A_833_48#_c_490_n N_A_27_74#_c_1288_n 0.00741157f $X=4.24 $Y=1.185
+ $X2=0 $Y2=0
cc_494 N_A_833_48#_c_491_n N_A_27_74#_c_1288_n 0.00839174f $X=4.595 $Y=1.26
+ $X2=0 $Y2=0
cc_495 N_A_833_48#_c_492_n N_A_27_74#_c_1288_n 0.0049686f $X=4.315 $Y=1.26 $X2=0
+ $Y2=0
cc_496 N_A_833_48#_c_493_n N_A_27_74#_c_1288_n 0.00605219f $X=4.67 $Y=1.185
+ $X2=0 $Y2=0
cc_497 N_A_833_48#_c_508_n N_A_27_74#_c_1288_n 0.00349533f $X=4.67 $Y=1.26 $X2=0
+ $Y2=0
cc_498 N_A_833_48#_c_493_n N_A_27_74#_c_1290_n 0.00112526f $X=4.67 $Y=1.185
+ $X2=0 $Y2=0
cc_499 N_A_833_48#_c_495_n N_A_27_74#_c_1290_n 0.00943354f $X=5.1 $Y=1.185 $X2=0
+ $Y2=0
cc_500 N_A_833_48#_c_497_n N_A_27_74#_c_1290_n 3.92634e-19 $X=5.53 $Y=1.185
+ $X2=0 $Y2=0
cc_501 N_A_833_48#_c_496_n N_A_27_74#_c_1291_n 0.00945505f $X=5.455 $Y=1.26
+ $X2=0 $Y2=0
cc_502 N_A_833_48#_c_509_n N_A_27_74#_c_1291_n 0.00691356f $X=5.1 $Y=1.26 $X2=0
+ $Y2=0
cc_503 N_A_833_48#_c_510_n N_A_27_74#_c_1291_n 0.00675192f $X=5.53 $Y=1.26 $X2=0
+ $Y2=0
cc_504 N_A_833_48#_c_495_n N_A_27_74#_c_1292_n 3.93664e-19 $X=5.1 $Y=1.185 $X2=0
+ $Y2=0
cc_505 N_A_833_48#_c_497_n N_A_27_74#_c_1292_n 0.0106304f $X=5.53 $Y=1.185 $X2=0
+ $Y2=0
cc_506 N_A_833_48#_c_498_n N_A_27_74#_c_1292_n 0.00787652f $X=5.885 $Y=1.26
+ $X2=0 $Y2=0
cc_507 N_A_833_48#_c_499_n N_A_27_74#_c_1292_n 0.00126428f $X=5.96 $Y=1.185
+ $X2=0 $Y2=0
cc_508 N_A_833_48#_c_510_n N_A_27_74#_c_1292_n 0.00308673f $X=5.53 $Y=1.26 $X2=0
+ $Y2=0
cc_509 N_A_833_48#_c_498_n N_A_27_74#_c_1293_n 0.0028859f $X=5.885 $Y=1.26 $X2=0
+ $Y2=0
cc_510 N_A_833_48#_c_500_n N_A_27_74#_c_1293_n 0.00777301f $X=6.315 $Y=1.26
+ $X2=0 $Y2=0
cc_511 N_A_833_48#_c_511_n N_A_27_74#_c_1293_n 0.00743366f $X=5.96 $Y=1.26 $X2=0
+ $Y2=0
cc_512 N_A_833_48#_c_512_n N_A_27_74#_c_1293_n 0.00675192f $X=6.39 $Y=1.26 $X2=0
+ $Y2=0
cc_513 N_A_833_48#_c_499_n N_A_27_74#_c_1294_n 4.44315e-19 $X=5.96 $Y=1.185
+ $X2=0 $Y2=0
cc_514 N_A_833_48#_c_501_n N_A_27_74#_c_1294_n 0.0106978f $X=6.39 $Y=1.185 $X2=0
+ $Y2=0
cc_515 N_A_833_48#_c_502_n N_A_27_74#_c_1294_n 0.00787652f $X=6.745 $Y=1.26
+ $X2=0 $Y2=0
cc_516 N_A_833_48#_c_503_n N_A_27_74#_c_1294_n 0.00126428f $X=6.82 $Y=1.185
+ $X2=0 $Y2=0
cc_517 N_A_833_48#_c_512_n N_A_27_74#_c_1294_n 0.00333129f $X=6.39 $Y=1.26 $X2=0
+ $Y2=0
cc_518 N_A_833_48#_c_502_n N_A_27_74#_c_1295_n 0.0028859f $X=6.745 $Y=1.26 $X2=0
+ $Y2=0
cc_519 N_A_833_48#_c_504_n N_A_27_74#_c_1295_n 0.00777301f $X=7.175 $Y=1.26
+ $X2=0 $Y2=0
cc_520 N_A_833_48#_c_506_n N_A_27_74#_c_1295_n 0.00293227f $X=7.72 $Y=1.26 $X2=0
+ $Y2=0
cc_521 N_A_833_48#_c_513_n N_A_27_74#_c_1295_n 0.00743366f $X=6.82 $Y=1.26 $X2=0
+ $Y2=0
cc_522 N_A_833_48#_c_514_n N_A_27_74#_c_1295_n 0.00701045f $X=7.25 $Y=1.26 $X2=0
+ $Y2=0
cc_523 N_A_833_48#_c_516_n N_A_27_74#_c_1295_n 0.00812414f $X=8.01 $Y=1.8 $X2=0
+ $Y2=0
cc_524 N_A_833_48#_c_503_n N_A_27_74#_c_1296_n 4.44315e-19 $X=6.82 $Y=1.185
+ $X2=0 $Y2=0
cc_525 N_A_833_48#_c_505_n N_A_27_74#_c_1296_n 0.011062f $X=7.25 $Y=1.185 $X2=0
+ $Y2=0
cc_526 N_A_833_48#_c_506_n N_A_27_74#_c_1296_n 0.00763221f $X=7.72 $Y=1.26 $X2=0
+ $Y2=0
cc_527 N_A_833_48#_c_507_n N_A_27_74#_c_1296_n 0.00481512f $X=7.795 $Y=1.185
+ $X2=0 $Y2=0
cc_528 N_A_833_48#_c_514_n N_A_27_74#_c_1296_n 0.00333129f $X=7.25 $Y=1.26 $X2=0
+ $Y2=0
cc_529 N_A_833_48#_c_515_n N_A_27_74#_c_1296_n 0.00117099f $X=7.87 $Y=0.505
+ $X2=0 $Y2=0
cc_530 N_A_833_48#_c_516_n N_A_27_74#_c_1296_n 0.0123137f $X=8.01 $Y=1.8 $X2=0
+ $Y2=0
cc_531 N_A_833_48#_c_517_n N_A_27_74#_c_1296_n 0.0423085f $X=8.095 $Y=0.675
+ $X2=0 $Y2=0
cc_532 N_A_833_48#_c_493_n N_A_27_74#_c_1300_n 0.00190168f $X=4.67 $Y=1.185
+ $X2=0 $Y2=0
cc_533 N_A_833_48#_c_494_n N_A_27_74#_c_1300_n 0.00829432f $X=5.025 $Y=1.26
+ $X2=0 $Y2=0
cc_534 N_A_833_48#_c_495_n N_A_27_74#_c_1300_n 0.00128545f $X=5.1 $Y=1.185 $X2=0
+ $Y2=0
cc_535 N_A_833_48#_c_508_n N_A_27_74#_c_1300_n 0.00207909f $X=4.67 $Y=1.26 $X2=0
+ $Y2=0
cc_536 N_A_833_48#_c_509_n N_A_27_74#_c_1300_n 0.00346919f $X=5.1 $Y=1.26 $X2=0
+ $Y2=0
cc_537 N_A_833_48#_c_498_n N_A_27_74#_c_1301_n 0.00231645f $X=5.885 $Y=1.26
+ $X2=0 $Y2=0
cc_538 N_A_833_48#_c_510_n N_A_27_74#_c_1301_n 2.58532e-19 $X=5.53 $Y=1.26 $X2=0
+ $Y2=0
cc_539 N_A_833_48#_c_502_n N_A_27_74#_c_1302_n 0.00231645f $X=6.745 $Y=1.26
+ $X2=0 $Y2=0
cc_540 N_A_833_48#_c_512_n N_A_27_74#_c_1302_n 2.58532e-19 $X=6.39 $Y=1.26 $X2=0
+ $Y2=0
cc_541 N_A_833_48#_c_490_n N_VGND_c_1446_n 0.0100283f $X=4.24 $Y=1.185 $X2=0
+ $Y2=0
cc_542 N_A_833_48#_c_491_n N_VGND_c_1446_n 7.11061e-19 $X=4.595 $Y=1.26 $X2=0
+ $Y2=0
cc_543 N_A_833_48#_c_493_n N_VGND_c_1446_n 0.0108109f $X=4.67 $Y=1.185 $X2=0
+ $Y2=0
cc_544 N_A_833_48#_c_495_n N_VGND_c_1446_n 5.57989e-19 $X=5.1 $Y=1.185 $X2=0
+ $Y2=0
cc_545 N_A_833_48#_c_495_n N_VGND_c_1447_n 0.001891f $X=5.1 $Y=1.185 $X2=0 $Y2=0
cc_546 N_A_833_48#_c_496_n N_VGND_c_1447_n 0.00230361f $X=5.455 $Y=1.26 $X2=0
+ $Y2=0
cc_547 N_A_833_48#_c_497_n N_VGND_c_1447_n 0.001891f $X=5.53 $Y=1.185 $X2=0
+ $Y2=0
cc_548 N_A_833_48#_c_497_n N_VGND_c_1448_n 6.16849e-19 $X=5.53 $Y=1.185 $X2=0
+ $Y2=0
cc_549 N_A_833_48#_c_499_n N_VGND_c_1448_n 0.0128208f $X=5.96 $Y=1.185 $X2=0
+ $Y2=0
cc_550 N_A_833_48#_c_500_n N_VGND_c_1448_n 0.00230361f $X=6.315 $Y=1.26 $X2=0
+ $Y2=0
cc_551 N_A_833_48#_c_501_n N_VGND_c_1448_n 0.00198331f $X=6.39 $Y=1.185 $X2=0
+ $Y2=0
cc_552 N_A_833_48#_c_501_n N_VGND_c_1449_n 6.16849e-19 $X=6.39 $Y=1.185 $X2=0
+ $Y2=0
cc_553 N_A_833_48#_c_503_n N_VGND_c_1449_n 0.0128208f $X=6.82 $Y=1.185 $X2=0
+ $Y2=0
cc_554 N_A_833_48#_c_504_n N_VGND_c_1449_n 0.00230361f $X=7.175 $Y=1.26 $X2=0
+ $Y2=0
cc_555 N_A_833_48#_c_505_n N_VGND_c_1449_n 0.00321968f $X=7.25 $Y=1.185 $X2=0
+ $Y2=0
cc_556 N_A_833_48#_c_517_n N_VGND_c_1449_n 3.11442e-19 $X=8.095 $Y=0.675 $X2=0
+ $Y2=0
cc_557 N_A_833_48#_c_519_n N_VGND_c_1450_n 0.0278867f $X=8.985 $Y=0.515 $X2=0
+ $Y2=0
cc_558 N_A_833_48#_c_490_n N_VGND_c_1453_n 0.00383152f $X=4.24 $Y=1.185 $X2=0
+ $Y2=0
cc_559 N_A_833_48#_c_493_n N_VGND_c_1455_n 0.00383152f $X=4.67 $Y=1.185 $X2=0
+ $Y2=0
cc_560 N_A_833_48#_c_495_n N_VGND_c_1455_n 0.00434272f $X=5.1 $Y=1.185 $X2=0
+ $Y2=0
cc_561 N_A_833_48#_c_497_n N_VGND_c_1457_n 0.00434272f $X=5.53 $Y=1.185 $X2=0
+ $Y2=0
cc_562 N_A_833_48#_c_499_n N_VGND_c_1457_n 0.00383152f $X=5.96 $Y=1.185 $X2=0
+ $Y2=0
cc_563 N_A_833_48#_c_501_n N_VGND_c_1459_n 0.00434272f $X=6.39 $Y=1.185 $X2=0
+ $Y2=0
cc_564 N_A_833_48#_c_503_n N_VGND_c_1459_n 0.00383152f $X=6.82 $Y=1.185 $X2=0
+ $Y2=0
cc_565 N_A_833_48#_c_505_n N_VGND_c_1460_n 0.00434272f $X=7.25 $Y=1.185 $X2=0
+ $Y2=0
cc_566 N_A_833_48#_c_515_n N_VGND_c_1460_n 0.00215305f $X=7.87 $Y=0.505 $X2=0
+ $Y2=0
cc_567 N_A_833_48#_c_517_n N_VGND_c_1460_n 0.0158548f $X=8.095 $Y=0.675 $X2=0
+ $Y2=0
cc_568 N_A_833_48#_c_518_n N_VGND_c_1460_n 0.0129945f $X=8.565 $Y=0.505 $X2=0
+ $Y2=0
cc_569 N_A_833_48#_c_519_n N_VGND_c_1460_n 0.0467562f $X=8.985 $Y=0.515 $X2=0
+ $Y2=0
cc_570 N_A_833_48#_c_490_n N_VGND_c_1464_n 0.00757637f $X=4.24 $Y=1.185 $X2=0
+ $Y2=0
cc_571 N_A_833_48#_c_493_n N_VGND_c_1464_n 0.0075754f $X=4.67 $Y=1.185 $X2=0
+ $Y2=0
cc_572 N_A_833_48#_c_495_n N_VGND_c_1464_n 0.00820284f $X=5.1 $Y=1.185 $X2=0
+ $Y2=0
cc_573 N_A_833_48#_c_497_n N_VGND_c_1464_n 0.00820284f $X=5.53 $Y=1.185 $X2=0
+ $Y2=0
cc_574 N_A_833_48#_c_499_n N_VGND_c_1464_n 0.0075754f $X=5.96 $Y=1.185 $X2=0
+ $Y2=0
cc_575 N_A_833_48#_c_501_n N_VGND_c_1464_n 0.00820284f $X=6.39 $Y=1.185 $X2=0
+ $Y2=0
cc_576 N_A_833_48#_c_503_n N_VGND_c_1464_n 0.0075754f $X=6.82 $Y=1.185 $X2=0
+ $Y2=0
cc_577 N_A_833_48#_c_505_n N_VGND_c_1464_n 0.00825283f $X=7.25 $Y=1.185 $X2=0
+ $Y2=0
cc_578 N_A_833_48#_c_517_n N_VGND_c_1464_n 0.0134631f $X=8.095 $Y=0.675 $X2=0
+ $Y2=0
cc_579 N_A_833_48#_c_518_n N_VGND_c_1464_n 0.0193081f $X=8.565 $Y=0.505 $X2=0
+ $Y2=0
cc_580 N_A_833_48#_c_519_n N_VGND_c_1464_n 0.0385205f $X=8.985 $Y=0.515 $X2=0
+ $Y2=0
cc_581 N_TE_B_c_675_n N_A_M1026_g 0.0461591f $X=9.11 $Y=1.385 $X2=0 $Y2=0
cc_582 N_TE_B_c_665_n N_A_c_838_n 0.0133063f $X=9.2 $Y=1.22 $X2=0 $Y2=0
cc_583 TE_B N_A_c_838_n 2.95037e-19 $X=9.275 $Y=1.21 $X2=0 $Y2=0
cc_584 N_TE_B_c_665_n A 2.69981e-19 $X=9.2 $Y=1.22 $X2=0 $Y2=0
cc_585 TE_B A 0.0309922f $X=9.275 $Y=1.21 $X2=0 $Y2=0
cc_586 TE_B N_A_c_842_n 0.00304313f $X=9.275 $Y=1.21 $X2=0 $Y2=0
cc_587 N_TE_B_c_675_n N_A_c_842_n 0.0180472f $X=9.11 $Y=1.385 $X2=0 $Y2=0
cc_588 N_TE_B_c_676_n N_A_28_368#_c_892_n 0.00344915f $X=4.26 $Y=1.765 $X2=0
+ $Y2=0
cc_589 N_TE_B_c_676_n N_A_28_368#_c_918_n 8.84747e-19 $X=4.26 $Y=1.765 $X2=0
+ $Y2=0
cc_590 N_TE_B_c_676_n N_A_28_368#_c_921_n 0.00555833f $X=4.26 $Y=1.765 $X2=0
+ $Y2=0
cc_591 N_TE_B_c_679_n N_A_28_368#_c_921_n 3.0069e-19 $X=4.81 $Y=1.765 $X2=0
+ $Y2=0
cc_592 N_TE_B_c_676_n N_A_28_368#_c_923_n 0.0100971f $X=4.26 $Y=1.765 $X2=0
+ $Y2=0
cc_593 N_TE_B_c_679_n N_A_28_368#_c_923_n 0.0100971f $X=4.81 $Y=1.765 $X2=0
+ $Y2=0
cc_594 N_TE_B_c_681_n N_A_28_368#_c_924_n 0.0100971f $X=5.26 $Y=1.765 $X2=0
+ $Y2=0
cc_595 N_TE_B_c_683_n N_A_28_368#_c_924_n 0.0100971f $X=5.81 $Y=1.765 $X2=0
+ $Y2=0
cc_596 N_TE_B_c_685_n N_A_28_368#_c_925_n 0.0100971f $X=6.26 $Y=1.765 $X2=0
+ $Y2=0
cc_597 N_TE_B_c_687_n N_A_28_368#_c_925_n 0.0111227f $X=6.81 $Y=1.765 $X2=0
+ $Y2=0
cc_598 N_TE_B_c_689_n N_A_28_368#_c_926_n 0.0122021f $X=7.26 $Y=1.765 $X2=0
+ $Y2=0
cc_599 N_TE_B_c_691_n N_A_28_368#_c_926_n 0.0108004f $X=7.88 $Y=1.765 $X2=0
+ $Y2=0
cc_600 N_TE_B_c_676_n N_A_28_368#_c_896_n 3.16734e-19 $X=4.26 $Y=1.765 $X2=0
+ $Y2=0
cc_601 N_TE_B_c_679_n N_A_28_368#_c_896_n 0.0077957f $X=4.81 $Y=1.765 $X2=0
+ $Y2=0
cc_602 N_TE_B_c_681_n N_A_28_368#_c_896_n 0.0077957f $X=5.26 $Y=1.765 $X2=0
+ $Y2=0
cc_603 N_TE_B_c_683_n N_A_28_368#_c_896_n 3.16734e-19 $X=5.81 $Y=1.765 $X2=0
+ $Y2=0
cc_604 N_TE_B_c_681_n N_A_28_368#_c_897_n 3.16734e-19 $X=5.26 $Y=1.765 $X2=0
+ $Y2=0
cc_605 N_TE_B_c_683_n N_A_28_368#_c_897_n 0.0077957f $X=5.81 $Y=1.765 $X2=0
+ $Y2=0
cc_606 N_TE_B_c_685_n N_A_28_368#_c_897_n 0.0077957f $X=6.26 $Y=1.765 $X2=0
+ $Y2=0
cc_607 N_TE_B_c_687_n N_A_28_368#_c_897_n 3.16734e-19 $X=6.81 $Y=1.765 $X2=0
+ $Y2=0
cc_608 N_TE_B_c_685_n N_A_28_368#_c_898_n 3.95442e-19 $X=6.26 $Y=1.765 $X2=0
+ $Y2=0
cc_609 N_TE_B_c_687_n N_A_28_368#_c_898_n 0.0083162f $X=6.81 $Y=1.765 $X2=0
+ $Y2=0
cc_610 N_TE_B_c_689_n N_A_28_368#_c_898_n 0.0102618f $X=7.26 $Y=1.765 $X2=0
+ $Y2=0
cc_611 N_TE_B_c_691_n N_A_28_368#_c_898_n 0.00160728f $X=7.88 $Y=1.765 $X2=0
+ $Y2=0
cc_612 N_TE_B_c_689_n N_A_28_368#_c_899_n 8.48629e-19 $X=7.26 $Y=1.765 $X2=0
+ $Y2=0
cc_613 N_TE_B_c_691_n N_A_28_368#_c_899_n 0.00703488f $X=7.88 $Y=1.765 $X2=0
+ $Y2=0
cc_614 N_TE_B_c_676_n N_VPWR_c_1153_n 0.00150551f $X=4.26 $Y=1.765 $X2=0 $Y2=0
cc_615 N_TE_B_c_679_n N_VPWR_c_1153_n 0.00203999f $X=4.81 $Y=1.765 $X2=0 $Y2=0
cc_616 N_TE_B_c_681_n N_VPWR_c_1154_n 0.00203999f $X=5.26 $Y=1.765 $X2=0 $Y2=0
cc_617 N_TE_B_c_683_n N_VPWR_c_1154_n 0.00203999f $X=5.81 $Y=1.765 $X2=0 $Y2=0
cc_618 N_TE_B_c_685_n N_VPWR_c_1155_n 0.00203999f $X=6.26 $Y=1.765 $X2=0 $Y2=0
cc_619 N_TE_B_c_687_n N_VPWR_c_1155_n 0.00343717f $X=6.81 $Y=1.765 $X2=0 $Y2=0
cc_620 N_TE_B_c_687_n N_VPWR_c_1156_n 0.005209f $X=6.81 $Y=1.765 $X2=0 $Y2=0
cc_621 N_TE_B_c_689_n N_VPWR_c_1156_n 0.00381803f $X=7.26 $Y=1.765 $X2=0 $Y2=0
cc_622 N_TE_B_c_689_n N_VPWR_c_1157_n 0.00378775f $X=7.26 $Y=1.765 $X2=0 $Y2=0
cc_623 N_TE_B_c_691_n N_VPWR_c_1157_n 0.00378775f $X=7.88 $Y=1.765 $X2=0 $Y2=0
cc_624 N_TE_B_c_694_n N_VPWR_c_1158_n 0.0262737f $X=9.105 $Y=1.765 $X2=0 $Y2=0
cc_625 N_TE_B_c_676_n N_VPWR_c_1161_n 0.00517089f $X=4.26 $Y=1.765 $X2=0 $Y2=0
cc_626 N_TE_B_c_679_n N_VPWR_c_1162_n 0.005209f $X=4.81 $Y=1.765 $X2=0 $Y2=0
cc_627 N_TE_B_c_681_n N_VPWR_c_1162_n 0.005209f $X=5.26 $Y=1.765 $X2=0 $Y2=0
cc_628 N_TE_B_c_683_n N_VPWR_c_1163_n 0.005209f $X=5.81 $Y=1.765 $X2=0 $Y2=0
cc_629 N_TE_B_c_685_n N_VPWR_c_1163_n 0.005209f $X=6.26 $Y=1.765 $X2=0 $Y2=0
cc_630 N_TE_B_c_691_n N_VPWR_c_1164_n 0.00381803f $X=7.88 $Y=1.765 $X2=0 $Y2=0
cc_631 N_TE_B_c_694_n N_VPWR_c_1164_n 0.00460063f $X=9.105 $Y=1.765 $X2=0 $Y2=0
cc_632 N_TE_B_c_676_n N_VPWR_c_1152_n 0.00515763f $X=4.26 $Y=1.765 $X2=0 $Y2=0
cc_633 N_TE_B_c_679_n N_VPWR_c_1152_n 0.00515684f $X=4.81 $Y=1.765 $X2=0 $Y2=0
cc_634 N_TE_B_c_681_n N_VPWR_c_1152_n 0.00515684f $X=5.26 $Y=1.765 $X2=0 $Y2=0
cc_635 N_TE_B_c_683_n N_VPWR_c_1152_n 0.00515684f $X=5.81 $Y=1.765 $X2=0 $Y2=0
cc_636 N_TE_B_c_685_n N_VPWR_c_1152_n 0.00515684f $X=6.26 $Y=1.765 $X2=0 $Y2=0
cc_637 N_TE_B_c_687_n N_VPWR_c_1152_n 0.00515684f $X=6.81 $Y=1.765 $X2=0 $Y2=0
cc_638 N_TE_B_c_689_n N_VPWR_c_1152_n 0.00475291f $X=7.26 $Y=1.765 $X2=0 $Y2=0
cc_639 N_TE_B_c_691_n N_VPWR_c_1152_n 0.00480425f $X=7.88 $Y=1.765 $X2=0 $Y2=0
cc_640 N_TE_B_c_694_n N_VPWR_c_1152_n 0.00913687f $X=9.105 $Y=1.765 $X2=0 $Y2=0
cc_641 N_TE_B_c_656_n N_A_27_74#_c_1288_n 0.00368482f $X=4.35 $Y=1.69 $X2=0
+ $Y2=0
cc_642 N_TE_B_c_657_n N_A_27_74#_c_1291_n 0.00592187f $X=5.17 $Y=1.69 $X2=0
+ $Y2=0
cc_643 N_TE_B_c_668_n N_A_27_74#_c_1293_n 0.00696604f $X=5.81 $Y=1.69 $X2=0
+ $Y2=0
cc_644 N_TE_B_c_660_n N_A_27_74#_c_1295_n 0.00696604f $X=6.72 $Y=1.69 $X2=0
+ $Y2=0
cc_645 N_TE_B_c_671_n N_A_27_74#_c_1295_n 0.00341127f $X=7.26 $Y=1.69 $X2=0
+ $Y2=0
cc_646 N_TE_B_c_666_n N_A_27_74#_c_1300_n 0.00448635f $X=4.81 $Y=1.69 $X2=0
+ $Y2=0
cc_647 N_TE_B_c_658_n N_A_27_74#_c_1301_n 0.003502f $X=5.72 $Y=1.69 $X2=0 $Y2=0
cc_648 N_TE_B_c_660_n N_A_27_74#_c_1302_n 0.00329532f $X=6.72 $Y=1.69 $X2=0
+ $Y2=0
cc_649 N_TE_B_c_665_n N_VGND_c_1450_n 0.00259633f $X=9.2 $Y=1.22 $X2=0 $Y2=0
cc_650 TE_B N_VGND_c_1450_n 0.0125437f $X=9.275 $Y=1.21 $X2=0 $Y2=0
cc_651 N_TE_B_c_665_n N_VGND_c_1460_n 0.00432935f $X=9.2 $Y=1.22 $X2=0 $Y2=0
cc_652 N_TE_B_c_665_n N_VGND_c_1464_n 0.00821561f $X=9.2 $Y=1.22 $X2=0 $Y2=0
cc_653 N_A_M1026_g N_VPWR_c_1158_n 0.00212264f $X=9.605 $Y=2.4 $X2=0 $Y2=0
cc_654 N_A_M1026_g N_VPWR_c_1160_n 6.0886e-19 $X=9.605 $Y=2.4 $X2=0 $Y2=0
cc_655 N_A_M1032_g N_VPWR_c_1160_n 0.0160409f $X=10.055 $Y=2.4 $X2=0 $Y2=0
cc_656 N_A_M1026_g N_VPWR_c_1165_n 0.005209f $X=9.605 $Y=2.4 $X2=0 $Y2=0
cc_657 N_A_M1032_g N_VPWR_c_1165_n 0.00460063f $X=10.055 $Y=2.4 $X2=0 $Y2=0
cc_658 N_A_M1026_g N_VPWR_c_1152_n 0.0098216f $X=9.605 $Y=2.4 $X2=0 $Y2=0
cc_659 N_A_M1032_g N_VPWR_c_1152_n 0.00908554f $X=10.055 $Y=2.4 $X2=0 $Y2=0
cc_660 N_A_c_838_n N_VGND_c_1450_n 0.00144568f $X=9.63 $Y=1.22 $X2=0 $Y2=0
cc_661 N_A_c_838_n N_VGND_c_1452_n 3.97405e-19 $X=9.63 $Y=1.22 $X2=0 $Y2=0
cc_662 N_A_c_840_n N_VGND_c_1452_n 0.00805371f $X=10.06 $Y=1.22 $X2=0 $Y2=0
cc_663 N_A_c_838_n N_VGND_c_1461_n 0.00434054f $X=9.63 $Y=1.22 $X2=0 $Y2=0
cc_664 N_A_c_840_n N_VGND_c_1461_n 0.00383152f $X=10.06 $Y=1.22 $X2=0 $Y2=0
cc_665 N_A_c_838_n N_VGND_c_1464_n 0.00820221f $X=9.63 $Y=1.22 $X2=0 $Y2=0
cc_666 N_A_c_840_n N_VGND_c_1464_n 0.00383967f $X=10.06 $Y=1.22 $X2=0 $Y2=0
cc_667 N_A_28_368#_c_888_n N_Z_M1001_d 0.00165831f $X=1.085 $Y=2.99 $X2=0 $Y2=0
cc_668 N_A_28_368#_c_890_n N_Z_M1005_d 0.00218982f $X=2.05 $Y=2.99 $X2=0 $Y2=0
cc_669 N_A_28_368#_c_891_n N_Z_M1008_d 0.00165831f $X=2.92 $Y=2.99 $X2=0 $Y2=0
cc_670 N_A_28_368#_c_892_n N_Z_M1014_d 0.00203037f $X=3.87 $Y=2.99 $X2=0 $Y2=0
cc_671 N_A_28_368#_c_888_n N_Z_c_1038_n 0.0177131f $X=1.085 $Y=2.99 $X2=0 $Y2=0
cc_672 N_A_28_368#_M1002_s N_Z_c_1030_n 0.00165831f $X=1.05 $Y=1.84 $X2=0 $Y2=0
cc_673 N_A_28_368#_c_910_n N_Z_c_1030_n 0.0148589f $X=1.185 $Y=2.325 $X2=0 $Y2=0
cc_674 N_A_28_368#_c_890_n N_Z_c_1053_n 0.0177084f $X=2.05 $Y=2.99 $X2=0 $Y2=0
cc_675 N_A_28_368#_M1006_s N_Z_c_1031_n 0.00165831f $X=2 $Y=1.84 $X2=0 $Y2=0
cc_676 N_A_28_368#_c_971_p N_Z_c_1031_n 0.0126919f $X=2.135 $Y=2.325 $X2=0 $Y2=0
cc_677 N_A_28_368#_c_891_n N_Z_c_1063_n 0.0159318f $X=2.92 $Y=2.99 $X2=0 $Y2=0
cc_678 N_A_28_368#_M1012_s N_Z_c_1032_n 0.00218982f $X=2.9 $Y=1.84 $X2=0 $Y2=0
cc_679 N_A_28_368#_c_974_p N_Z_c_1032_n 0.0167599f $X=3.085 $Y=2.325 $X2=0 $Y2=0
cc_680 N_A_28_368#_c_892_n N_Z_c_1083_n 0.0165667f $X=3.87 $Y=2.99 $X2=0 $Y2=0
cc_681 N_A_28_368#_c_887_n N_Z_c_1034_n 0.00774108f $X=0.285 $Y=1.985 $X2=0
+ $Y2=0
cc_682 N_A_28_368#_c_923_n N_VPWR_M1009_s 0.00532667f $X=4.87 $Y=2.475 $X2=-0.19
+ $Y2=1.66
cc_683 N_A_28_368#_c_924_n N_VPWR_M1015_s 0.00532667f $X=5.87 $Y=2.475 $X2=0
+ $Y2=0
cc_684 N_A_28_368#_c_925_n N_VPWR_M1017_s 0.00532667f $X=6.87 $Y=2.475 $X2=0
+ $Y2=0
cc_685 N_A_28_368#_c_926_n N_VPWR_M1021_s 0.00823786f $X=7.94 $Y=2.645 $X2=0
+ $Y2=0
cc_686 N_A_28_368#_c_892_n N_VPWR_c_1153_n 0.0119238f $X=3.87 $Y=2.99 $X2=0
+ $Y2=0
cc_687 N_A_28_368#_c_923_n N_VPWR_c_1153_n 0.0202465f $X=4.87 $Y=2.475 $X2=0
+ $Y2=0
cc_688 N_A_28_368#_c_896_n N_VPWR_c_1153_n 0.0101711f $X=5.035 $Y=2.475 $X2=0
+ $Y2=0
cc_689 N_A_28_368#_c_924_n N_VPWR_c_1154_n 0.0202465f $X=5.87 $Y=2.475 $X2=0
+ $Y2=0
cc_690 N_A_28_368#_c_896_n N_VPWR_c_1154_n 0.0101711f $X=5.035 $Y=2.475 $X2=0
+ $Y2=0
cc_691 N_A_28_368#_c_897_n N_VPWR_c_1154_n 0.0101711f $X=6.035 $Y=2.475 $X2=0
+ $Y2=0
cc_692 N_A_28_368#_c_925_n N_VPWR_c_1155_n 0.0202465f $X=6.87 $Y=2.475 $X2=0
+ $Y2=0
cc_693 N_A_28_368#_c_897_n N_VPWR_c_1155_n 0.0101711f $X=6.035 $Y=2.475 $X2=0
+ $Y2=0
cc_694 N_A_28_368#_c_898_n N_VPWR_c_1155_n 0.0101711f $X=7.035 $Y=2.475 $X2=0
+ $Y2=0
cc_695 N_A_28_368#_c_926_n N_VPWR_c_1156_n 0.00324117f $X=7.94 $Y=2.645 $X2=0
+ $Y2=0
cc_696 N_A_28_368#_c_898_n N_VPWR_c_1156_n 0.0143153f $X=7.035 $Y=2.475 $X2=0
+ $Y2=0
cc_697 N_A_28_368#_c_926_n N_VPWR_c_1157_n 0.0245684f $X=7.94 $Y=2.645 $X2=0
+ $Y2=0
cc_698 N_A_28_368#_c_898_n N_VPWR_c_1157_n 0.00327717f $X=7.035 $Y=2.475 $X2=0
+ $Y2=0
cc_699 N_A_28_368#_c_899_n N_VPWR_c_1157_n 0.00327717f $X=8.105 $Y=2.645 $X2=0
+ $Y2=0
cc_700 N_A_28_368#_c_888_n N_VPWR_c_1161_n 0.0449528f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_701 N_A_28_368#_c_889_n N_VPWR_c_1161_n 0.0179217f $X=0.37 $Y=2.99 $X2=0
+ $Y2=0
cc_702 N_A_28_368#_c_890_n N_VPWR_c_1161_n 0.0440768f $X=2.05 $Y=2.99 $X2=0
+ $Y2=0
cc_703 N_A_28_368#_c_891_n N_VPWR_c_1161_n 0.0439866f $X=2.92 $Y=2.99 $X2=0
+ $Y2=0
cc_704 N_A_28_368#_c_892_n N_VPWR_c_1161_n 0.0662563f $X=3.87 $Y=2.99 $X2=0
+ $Y2=0
cc_705 N_A_28_368#_c_893_n N_VPWR_c_1161_n 0.0188916f $X=1.217 $Y=2.99 $X2=0
+ $Y2=0
cc_706 N_A_28_368#_c_894_n N_VPWR_c_1161_n 0.0121867f $X=2.135 $Y=2.99 $X2=0
+ $Y2=0
cc_707 N_A_28_368#_c_895_n N_VPWR_c_1161_n 0.0193554f $X=3.055 $Y=2.99 $X2=0
+ $Y2=0
cc_708 N_A_28_368#_c_896_n N_VPWR_c_1162_n 0.0143153f $X=5.035 $Y=2.475 $X2=0
+ $Y2=0
cc_709 N_A_28_368#_c_897_n N_VPWR_c_1163_n 0.0143153f $X=6.035 $Y=2.475 $X2=0
+ $Y2=0
cc_710 N_A_28_368#_c_926_n N_VPWR_c_1164_n 0.00324117f $X=7.94 $Y=2.645 $X2=0
+ $Y2=0
cc_711 N_A_28_368#_c_899_n N_VPWR_c_1164_n 0.0140571f $X=8.105 $Y=2.645 $X2=0
+ $Y2=0
cc_712 N_A_28_368#_c_888_n N_VPWR_c_1152_n 0.0252362f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_713 N_A_28_368#_c_889_n N_VPWR_c_1152_n 0.00971942f $X=0.37 $Y=2.99 $X2=0
+ $Y2=0
cc_714 N_A_28_368#_c_890_n N_VPWR_c_1152_n 0.0248093f $X=2.05 $Y=2.99 $X2=0
+ $Y2=0
cc_715 N_A_28_368#_c_891_n N_VPWR_c_1152_n 0.0246722f $X=2.92 $Y=2.99 $X2=0
+ $Y2=0
cc_716 N_A_28_368#_c_892_n N_VPWR_c_1152_n 0.0366153f $X=3.87 $Y=2.99 $X2=0
+ $Y2=0
cc_717 N_A_28_368#_c_923_n N_VPWR_c_1152_n 0.0115311f $X=4.87 $Y=2.475 $X2=0
+ $Y2=0
cc_718 N_A_28_368#_c_924_n N_VPWR_c_1152_n 0.0115311f $X=5.87 $Y=2.475 $X2=0
+ $Y2=0
cc_719 N_A_28_368#_c_925_n N_VPWR_c_1152_n 0.0115442f $X=6.87 $Y=2.475 $X2=0
+ $Y2=0
cc_720 N_A_28_368#_c_926_n N_VPWR_c_1152_n 0.0121916f $X=7.94 $Y=2.645 $X2=0
+ $Y2=0
cc_721 N_A_28_368#_c_893_n N_VPWR_c_1152_n 0.0101653f $X=1.217 $Y=2.99 $X2=0
+ $Y2=0
cc_722 N_A_28_368#_c_894_n N_VPWR_c_1152_n 0.00660921f $X=2.135 $Y=2.99 $X2=0
+ $Y2=0
cc_723 N_A_28_368#_c_895_n N_VPWR_c_1152_n 0.010497f $X=3.055 $Y=2.99 $X2=0
+ $Y2=0
cc_724 N_A_28_368#_c_896_n N_VPWR_c_1152_n 0.0117766f $X=5.035 $Y=2.475 $X2=0
+ $Y2=0
cc_725 N_A_28_368#_c_897_n N_VPWR_c_1152_n 0.0117766f $X=6.035 $Y=2.475 $X2=0
+ $Y2=0
cc_726 N_A_28_368#_c_898_n N_VPWR_c_1152_n 0.0117766f $X=7.035 $Y=2.475 $X2=0
+ $Y2=0
cc_727 N_A_28_368#_c_899_n N_VPWR_c_1152_n 0.011784f $X=8.105 $Y=2.645 $X2=0
+ $Y2=0
cc_728 N_Z_c_1023_n N_A_27_74#_M1013_d 0.00221449f $X=1.43 $Y=1.065 $X2=0 $Y2=0
cc_729 N_Z_c_1024_n N_A_27_74#_M1027_d 0.00250873f $X=2.43 $Y=1.065 $X2=0 $Y2=0
cc_730 N_Z_c_1025_n N_A_27_74#_M1031_d 0.00270388f $X=3.43 $Y=1.065 $X2=0 $Y2=0
cc_731 Z N_A_27_74#_c_1281_n 0.00676472f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_732 N_Z_M1007_s N_A_27_74#_c_1282_n 0.00176461f $X=0.57 $Y=0.37 $X2=0 $Y2=0
cc_733 N_Z_c_1023_n N_A_27_74#_c_1282_n 0.00319222f $X=1.43 $Y=1.065 $X2=0 $Y2=0
cc_734 N_Z_c_1110_n N_A_27_74#_c_1282_n 0.0159544f $X=0.71 $Y=0.76 $X2=0 $Y2=0
cc_735 N_Z_c_1023_n N_A_27_74#_c_1306_n 0.0133644f $X=1.43 $Y=1.065 $X2=0 $Y2=0
cc_736 N_Z_c_1049_n N_A_27_74#_c_1306_n 0.0137413f $X=1.595 $Y=0.76 $X2=0 $Y2=0
cc_737 N_Z_M1019_s N_A_27_74#_c_1284_n 0.00176461f $X=1.455 $Y=0.37 $X2=0 $Y2=0
cc_738 N_Z_c_1023_n N_A_27_74#_c_1284_n 0.00386975f $X=1.43 $Y=1.065 $X2=0 $Y2=0
cc_739 N_Z_c_1049_n N_A_27_74#_c_1284_n 0.0157331f $X=1.595 $Y=0.76 $X2=0 $Y2=0
cc_740 N_Z_c_1024_n N_A_27_74#_c_1284_n 0.00319222f $X=2.43 $Y=1.065 $X2=0 $Y2=0
cc_741 N_Z_c_1024_n N_A_27_74#_c_1309_n 0.0206429f $X=2.43 $Y=1.065 $X2=0 $Y2=0
cc_742 N_Z_M1030_s N_A_27_74#_c_1285_n 0.00250873f $X=2.385 $Y=0.37 $X2=0 $Y2=0
cc_743 N_Z_c_1024_n N_A_27_74#_c_1285_n 0.00319222f $X=2.43 $Y=1.065 $X2=0 $Y2=0
cc_744 N_Z_c_1067_n N_A_27_74#_c_1285_n 0.0193319f $X=2.595 $Y=0.76 $X2=0 $Y2=0
cc_745 N_Z_c_1025_n N_A_27_74#_c_1285_n 0.00319222f $X=3.43 $Y=1.065 $X2=0 $Y2=0
cc_746 N_Z_c_1025_n N_A_27_74#_c_1313_n 0.0207199f $X=3.43 $Y=1.065 $X2=0 $Y2=0
cc_747 N_Z_M1033_s N_A_27_74#_c_1286_n 0.00234927f $X=3.4 $Y=0.37 $X2=0 $Y2=0
cc_748 N_Z_c_1025_n N_A_27_74#_c_1286_n 0.00357683f $X=3.43 $Y=1.065 $X2=0 $Y2=0
cc_749 N_Z_c_1085_n N_A_27_74#_c_1286_n 0.0182078f $X=3.595 $Y=0.76 $X2=0 $Y2=0
cc_750 N_Z_c_1025_n N_A_27_74#_c_1287_n 0.00745191f $X=3.43 $Y=1.065 $X2=0 $Y2=0
cc_751 N_Z_c_1025_n N_A_27_74#_c_1289_n 8.53482e-19 $X=3.43 $Y=1.065 $X2=0 $Y2=0
cc_752 N_A_27_74#_c_1286_n N_VGND_c_1446_n 0.0112234f $X=3.94 $Y=0.34 $X2=0
+ $Y2=0
cc_753 N_A_27_74#_c_1288_n N_VGND_c_1446_n 0.0216086f $X=4.72 $Y=1.225 $X2=0
+ $Y2=0
cc_754 N_A_27_74#_c_1290_n N_VGND_c_1446_n 0.0229496f $X=4.885 $Y=0.515 $X2=0
+ $Y2=0
cc_755 N_A_27_74#_c_1290_n N_VGND_c_1447_n 0.0281649f $X=4.885 $Y=0.515 $X2=0
+ $Y2=0
cc_756 N_A_27_74#_c_1291_n N_VGND_c_1447_n 0.0135549f $X=5.58 $Y=1.385 $X2=0
+ $Y2=0
cc_757 N_A_27_74#_c_1292_n N_VGND_c_1447_n 0.0281649f $X=5.745 $Y=0.515 $X2=0
+ $Y2=0
cc_758 N_A_27_74#_c_1292_n N_VGND_c_1448_n 0.0282477f $X=5.745 $Y=0.515 $X2=0
+ $Y2=0
cc_759 N_A_27_74#_c_1293_n N_VGND_c_1448_n 0.0198685f $X=6.44 $Y=1.385 $X2=0
+ $Y2=0
cc_760 N_A_27_74#_c_1294_n N_VGND_c_1448_n 0.0282477f $X=6.605 $Y=0.515 $X2=0
+ $Y2=0
cc_761 N_A_27_74#_c_1294_n N_VGND_c_1449_n 0.0282477f $X=6.605 $Y=0.515 $X2=0
+ $Y2=0
cc_762 N_A_27_74#_c_1295_n N_VGND_c_1449_n 0.0198685f $X=7.3 $Y=1.385 $X2=0
+ $Y2=0
cc_763 N_A_27_74#_c_1296_n N_VGND_c_1449_n 0.0282477f $X=7.465 $Y=0.515 $X2=0
+ $Y2=0
cc_764 N_A_27_74#_c_1282_n N_VGND_c_1453_n 0.043517f $X=1.055 $Y=0.34 $X2=0
+ $Y2=0
cc_765 N_A_27_74#_c_1283_n N_VGND_c_1453_n 0.0179217f $X=0.365 $Y=0.34 $X2=0
+ $Y2=0
cc_766 N_A_27_74#_c_1284_n N_VGND_c_1453_n 0.0444833f $X=1.93 $Y=0.34 $X2=0
+ $Y2=0
cc_767 N_A_27_74#_c_1285_n N_VGND_c_1453_n 0.0423044f $X=2.93 $Y=0.34 $X2=0
+ $Y2=0
cc_768 N_A_27_74#_c_1286_n N_VGND_c_1453_n 0.0550916f $X=3.94 $Y=0.34 $X2=0
+ $Y2=0
cc_769 N_A_27_74#_c_1297_n N_VGND_c_1453_n 0.0120038f $X=1.14 $Y=0.34 $X2=0
+ $Y2=0
cc_770 N_A_27_74#_c_1298_n N_VGND_c_1453_n 0.0232138f $X=2.095 $Y=0.34 $X2=0
+ $Y2=0
cc_771 N_A_27_74#_c_1299_n N_VGND_c_1453_n 0.0232651f $X=3.095 $Y=0.34 $X2=0
+ $Y2=0
cc_772 N_A_27_74#_c_1290_n N_VGND_c_1455_n 0.0109942f $X=4.885 $Y=0.515 $X2=0
+ $Y2=0
cc_773 N_A_27_74#_c_1292_n N_VGND_c_1457_n 0.0109942f $X=5.745 $Y=0.515 $X2=0
+ $Y2=0
cc_774 N_A_27_74#_c_1294_n N_VGND_c_1459_n 0.0109942f $X=6.605 $Y=0.515 $X2=0
+ $Y2=0
cc_775 N_A_27_74#_c_1296_n N_VGND_c_1460_n 0.0109942f $X=7.465 $Y=0.515 $X2=0
+ $Y2=0
cc_776 N_A_27_74#_c_1282_n N_VGND_c_1464_n 0.0245693f $X=1.055 $Y=0.34 $X2=0
+ $Y2=0
cc_777 N_A_27_74#_c_1283_n N_VGND_c_1464_n 0.00971942f $X=0.365 $Y=0.34 $X2=0
+ $Y2=0
cc_778 N_A_27_74#_c_1284_n N_VGND_c_1464_n 0.0251332f $X=1.93 $Y=0.34 $X2=0
+ $Y2=0
cc_779 N_A_27_74#_c_1285_n N_VGND_c_1464_n 0.0239316f $X=2.93 $Y=0.34 $X2=0
+ $Y2=0
cc_780 N_A_27_74#_c_1286_n N_VGND_c_1464_n 0.0308486f $X=3.94 $Y=0.34 $X2=0
+ $Y2=0
cc_781 N_A_27_74#_c_1290_n N_VGND_c_1464_n 0.00904371f $X=4.885 $Y=0.515 $X2=0
+ $Y2=0
cc_782 N_A_27_74#_c_1292_n N_VGND_c_1464_n 0.00904371f $X=5.745 $Y=0.515 $X2=0
+ $Y2=0
cc_783 N_A_27_74#_c_1294_n N_VGND_c_1464_n 0.00904371f $X=6.605 $Y=0.515 $X2=0
+ $Y2=0
cc_784 N_A_27_74#_c_1296_n N_VGND_c_1464_n 0.00904371f $X=7.465 $Y=0.515 $X2=0
+ $Y2=0
cc_785 N_A_27_74#_c_1297_n N_VGND_c_1464_n 0.00657483f $X=1.14 $Y=0.34 $X2=0
+ $Y2=0
cc_786 N_A_27_74#_c_1298_n N_VGND_c_1464_n 0.0126482f $X=2.095 $Y=0.34 $X2=0
+ $Y2=0
cc_787 N_A_27_74#_c_1299_n N_VGND_c_1464_n 0.0127168f $X=3.095 $Y=0.34 $X2=0
+ $Y2=0

* File: sky130_fd_sc_ms__a22oi_1.pxi.spice
* Created: Fri Aug 28 17:03:18 2020
* 
x_PM_SKY130_FD_SC_MS__A22OI_1%B2 N_B2_M1004_g N_B2_c_51_n N_B2_M1001_g
+ N_B2_c_52_n N_B2_c_53_n B2 B2 PM_SKY130_FD_SC_MS__A22OI_1%B2
x_PM_SKY130_FD_SC_MS__A22OI_1%B1 N_B1_M1000_g N_B1_M1005_g B1 N_B1_c_83_n
+ N_B1_c_84_n PM_SKY130_FD_SC_MS__A22OI_1%B1
x_PM_SKY130_FD_SC_MS__A22OI_1%A1 N_A1_M1003_g N_A1_M1002_g A1 N_A1_c_121_n
+ N_A1_c_122_n PM_SKY130_FD_SC_MS__A22OI_1%A1
x_PM_SKY130_FD_SC_MS__A22OI_1%A2 N_A2_M1007_g N_A2_M1006_g A2 A2 N_A2_c_157_n
+ PM_SKY130_FD_SC_MS__A22OI_1%A2
x_PM_SKY130_FD_SC_MS__A22OI_1%A_71_368# N_A_71_368#_M1004_s N_A_71_368#_M1005_d
+ N_A_71_368#_M1006_d N_A_71_368#_c_185_n N_A_71_368#_c_186_n
+ N_A_71_368#_c_187_n N_A_71_368#_c_197_n N_A_71_368#_c_194_n
+ N_A_71_368#_c_202_n N_A_71_368#_c_188_n N_A_71_368#_c_189_n
+ PM_SKY130_FD_SC_MS__A22OI_1%A_71_368#
x_PM_SKY130_FD_SC_MS__A22OI_1%Y N_Y_M1000_d N_Y_M1004_d N_Y_c_226_n N_Y_c_227_n
+ N_Y_c_228_n N_Y_c_233_n Y Y PM_SKY130_FD_SC_MS__A22OI_1%Y
x_PM_SKY130_FD_SC_MS__A22OI_1%VPWR N_VPWR_M1002_d N_VPWR_c_263_n N_VPWR_c_264_n
+ N_VPWR_c_265_n VPWR N_VPWR_c_266_n N_VPWR_c_262_n
+ PM_SKY130_FD_SC_MS__A22OI_1%VPWR
x_PM_SKY130_FD_SC_MS__A22OI_1%VGND N_VGND_M1001_s N_VGND_M1007_d N_VGND_c_290_n
+ N_VGND_c_291_n N_VGND_c_292_n N_VGND_c_293_n N_VGND_c_294_n N_VGND_c_295_n
+ VGND N_VGND_c_296_n N_VGND_c_297_n PM_SKY130_FD_SC_MS__A22OI_1%VGND
cc_1 VNB N_B2_M1004_g 0.00631372f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.4
cc_2 VNB N_B2_c_51_n 0.018672f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.22
cc_3 VNB N_B2_c_52_n 0.0687936f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.385
cc_4 VNB N_B2_c_53_n 0.0105106f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.385
cc_5 VNB B2 0.0170831f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_B1_M1000_g 0.0244201f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.4
cc_7 VNB N_B1_c_83_n 0.026255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B1_c_84_n 0.00166449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A1_M1003_g 0.0273876f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.4
cc_10 VNB N_A1_c_121_n 0.0262412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A1_c_122_n 0.00689463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_M1007_g 0.0338413f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.4
cc_13 VNB A2 0.0275005f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_14 VNB N_A2_c_157_n 0.027381f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_15 VNB N_Y_c_226_n 0.0155629f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.74
cc_16 VNB N_Y_c_227_n 0.0028102f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.385
cc_17 VNB N_Y_c_228_n 0.00336771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB Y 0.00493162f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_19 VNB N_VPWR_c_262_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_20 VNB N_VGND_c_290_n 0.0285265f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.385
cc_21 VNB N_VGND_c_291_n 0.0419806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_292_n 0.0129628f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.385
cc_23 VNB N_VGND_c_293_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_294_n 0.0452046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_295_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_296_n 0.0129628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_297_n 0.214622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VPB N_B2_M1004_g 0.0250413f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=2.4
cc_29 VPB B2 0.0160066f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_30 VPB N_B1_M1005_g 0.020253f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_31 VPB N_B1_c_83_n 0.00556367f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_32 VPB N_B1_c_84_n 0.00410931f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_33 VPB N_A1_M1002_g 0.0216409f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_34 VPB N_A1_c_121_n 0.00562372f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_A1_c_122_n 0.00200044f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_A2_M1006_g 0.0288606f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_37 VPB A2 0.0168401f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_38 VPB N_A2_c_157_n 0.00576404f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_39 VPB N_A_71_368#_c_185_n 0.0243557f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A_71_368#_c_186_n 0.00457669f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_41 VPB N_A_71_368#_c_187_n 0.00969936f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_42 VPB N_A_71_368#_c_188_n 0.0075508f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.665
cc_43 VPB N_A_71_368#_c_189_n 0.0358769f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_44 VPB Y 0.00456928f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.665
cc_45 VPB N_VPWR_c_263_n 0.00678734f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=0.74
cc_46 VPB N_VPWR_c_264_n 0.0446773f $X=-0.19 $Y=1.66 $X2=0.705 $Y2=1.385
cc_47 VPB N_VPWR_c_265_n 0.00653059f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_48 VPB N_VPWR_c_266_n 0.0255159f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.385
cc_49 VPB N_VPWR_c_262_n 0.0714703f $X=-0.19 $Y=1.66 $X2=0.27 $Y2=1.665
cc_50 N_B2_c_51_n N_B1_M1000_g 0.0432601f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_51 N_B2_M1004_g N_B1_M1005_g 0.0282551f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_52 N_B2_c_53_n N_B1_c_83_n 0.0432601f $X=0.705 $Y=1.385 $X2=0 $Y2=0
cc_53 N_B2_M1004_g N_B1_c_84_n 3.16626e-19 $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_54 N_B2_c_53_n N_B1_c_84_n 3.78988e-19 $X=0.705 $Y=1.385 $X2=0 $Y2=0
cc_55 N_B2_M1004_g N_A_71_368#_c_185_n 0.00892729f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_56 B2 N_A_71_368#_c_185_n 0.00493998f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_57 N_B2_M1004_g N_A_71_368#_c_186_n 0.0115958f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_58 N_B2_M1004_g N_A_71_368#_c_187_n 0.00291744f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_59 N_B2_M1004_g N_A_71_368#_c_194_n 6.26485e-19 $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_60 N_B2_c_51_n N_Y_c_227_n 0.0133235f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_61 N_B2_c_51_n N_Y_c_228_n 0.00217641f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_62 N_B2_M1004_g N_Y_c_233_n 0.0127764f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_63 N_B2_M1004_g Y 0.0141652f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_64 N_B2_c_51_n Y 0.00119049f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_65 N_B2_c_52_n Y 0.00514616f $X=0.615 $Y=1.385 $X2=0 $Y2=0
cc_66 N_B2_c_53_n Y 0.00696127f $X=0.705 $Y=1.385 $X2=0 $Y2=0
cc_67 B2 Y 0.045939f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_68 N_B2_M1004_g N_VPWR_c_264_n 0.00333896f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_69 N_B2_M1004_g N_VPWR_c_262_n 0.0042706f $X=0.705 $Y=2.4 $X2=0 $Y2=0
cc_70 N_B2_c_51_n N_VGND_c_290_n 0.0154153f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_71 N_B2_c_52_n N_VGND_c_290_n 0.00639332f $X=0.615 $Y=1.385 $X2=0 $Y2=0
cc_72 B2 N_VGND_c_290_n 0.00521723f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_73 N_B2_c_51_n N_VGND_c_294_n 0.00383152f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_74 N_B2_c_51_n N_VGND_c_297_n 0.0075694f $X=0.72 $Y=1.22 $X2=0 $Y2=0
cc_75 N_B1_M1000_g N_A1_M1003_g 0.014794f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_76 N_B1_M1005_g N_A1_M1002_g 0.0160353f $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_77 N_B1_c_84_n N_A1_M1002_g 6.26118e-19 $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_78 N_B1_c_83_n N_A1_c_121_n 0.0201104f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_79 N_B1_c_84_n N_A1_c_121_n 0.00114936f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_80 N_B1_c_83_n N_A1_c_122_n 0.00114936f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_81 N_B1_c_84_n N_A1_c_122_n 0.0276388f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_82 N_B1_M1005_g N_A_71_368#_c_185_n 5.73047e-19 $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_83 N_B1_M1005_g N_A_71_368#_c_186_n 0.0136313f $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_84 N_B1_M1005_g N_A_71_368#_c_197_n 0.00242345f $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_85 N_B1_c_83_n N_A_71_368#_c_197_n 4.052e-19 $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_86 N_B1_c_84_n N_A_71_368#_c_197_n 0.00774613f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_87 N_B1_M1005_g N_A_71_368#_c_194_n 0.0105282f $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_88 N_B1_M1000_g N_Y_c_226_n 0.0124193f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_89 N_B1_c_83_n N_Y_c_226_n 0.00140824f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_90 N_B1_c_84_n N_Y_c_226_n 0.0265531f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_91 N_B1_M1000_g N_Y_c_228_n 0.012242f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_92 N_B1_c_84_n N_Y_c_233_n 4.64867e-19 $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_93 N_B1_M1000_g Y 0.00536895f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_94 N_B1_M1005_g Y 0.0017316f $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_95 N_B1_c_84_n Y 0.0334882f $X=1.17 $Y=1.515 $X2=0 $Y2=0
cc_96 N_B1_M1005_g N_VPWR_c_263_n 3.13927e-19 $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_97 N_B1_M1005_g N_VPWR_c_264_n 0.00333896f $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_98 N_B1_M1005_g N_VPWR_c_262_n 0.00423185f $X=1.155 $Y=2.4 $X2=0 $Y2=0
cc_99 N_B1_M1000_g N_VGND_c_290_n 0.00190254f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_100 N_B1_M1000_g N_VGND_c_294_n 0.00434272f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_101 N_B1_M1000_g N_VGND_c_297_n 0.00821699f $X=1.08 $Y=0.74 $X2=0 $Y2=0
cc_102 N_A1_M1003_g N_A2_M1007_g 0.0328884f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_103 N_A1_M1002_g N_A2_M1006_g 0.0239398f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_104 N_A1_c_122_n N_A2_M1006_g 3.34283e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_105 N_A1_M1002_g A2 2.9613e-19 $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_106 N_A1_c_121_n A2 0.00201442f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_107 N_A1_c_122_n A2 0.0366314f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_108 N_A1_c_121_n N_A2_c_157_n 0.0206382f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_109 N_A1_c_122_n N_A2_c_157_n 3.7859e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_110 N_A1_M1002_g N_A_71_368#_c_186_n 0.00110243f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_111 N_A1_M1002_g N_A_71_368#_c_202_n 0.0153112f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_112 N_A1_c_121_n N_A_71_368#_c_202_n 7.08634e-19 $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_113 N_A1_c_122_n N_A_71_368#_c_202_n 0.0229716f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_114 N_A1_M1002_g N_A_71_368#_c_189_n 8.67149e-19 $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_115 N_A1_M1003_g N_Y_c_226_n 0.00484582f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A1_c_122_n N_Y_c_226_n 0.00196319f $X=1.71 $Y=1.515 $X2=0 $Y2=0
cc_117 N_A1_M1003_g N_Y_c_228_n 0.0144523f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_118 N_A1_M1002_g N_VPWR_c_263_n 0.0106839f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A1_M1002_g N_VPWR_c_264_n 0.00521592f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A1_M1002_g N_VPWR_c_262_n 0.0102937f $X=1.635 $Y=2.4 $X2=0 $Y2=0
cc_121 N_A1_M1003_g N_VGND_c_291_n 0.00294701f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_122 N_A1_M1003_g N_VGND_c_294_n 0.00434272f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_123 N_A1_M1003_g N_VGND_c_297_n 0.00823328f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_124 N_A2_M1006_g N_A_71_368#_c_202_n 0.0133817f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_125 A2 N_A_71_368#_c_202_n 0.012644f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_126 N_A2_M1006_g N_A_71_368#_c_188_n 8.84614e-19 $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_127 A2 N_A_71_368#_c_188_n 0.0264311f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_128 N_A2_c_157_n N_A_71_368#_c_188_n 7.81657e-19 $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_129 N_A2_M1006_g N_A_71_368#_c_189_n 0.0119414f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_130 N_A2_M1007_g N_Y_c_226_n 6.02297e-19 $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_131 N_A2_M1007_g N_Y_c_228_n 0.00204985f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_132 N_A2_M1006_g N_VPWR_c_263_n 0.00345508f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_133 N_A2_M1006_g N_VPWR_c_266_n 0.005209f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_134 N_A2_M1006_g N_VPWR_c_262_n 0.0098676f $X=2.175 $Y=2.4 $X2=0 $Y2=0
cc_135 N_A2_M1007_g N_VGND_c_291_n 0.022716f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_136 A2 N_VGND_c_291_n 0.0236581f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_137 N_A2_c_157_n N_VGND_c_291_n 0.00419666f $X=2.25 $Y=1.515 $X2=0 $Y2=0
cc_138 N_A2_M1007_g N_VGND_c_294_n 0.00383152f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A2_M1007_g N_VGND_c_297_n 0.00758569f $X=2.16 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A_71_368#_c_186_n N_Y_M1004_d 0.00165831f $X=1.215 $Y=2.99 $X2=0 $Y2=0
cc_141 N_A_71_368#_c_185_n N_Y_c_233_n 0.00216696f $X=0.48 $Y=2.455 $X2=0 $Y2=0
cc_142 N_A_71_368#_c_186_n N_Y_c_233_n 0.0117822f $X=1.215 $Y=2.99 $X2=0 $Y2=0
cc_143 N_A_71_368#_c_202_n N_VPWR_M1002_d 0.00928873f $X=2.235 $Y=2.035
+ $X2=-0.19 $Y2=1.66
cc_144 N_A_71_368#_c_186_n N_VPWR_c_263_n 0.0138772f $X=1.215 $Y=2.99 $X2=0
+ $Y2=0
cc_145 N_A_71_368#_c_194_n N_VPWR_c_263_n 0.0488299f $X=1.38 $Y=2.815 $X2=0
+ $Y2=0
cc_146 N_A_71_368#_c_202_n N_VPWR_c_263_n 0.0206577f $X=2.235 $Y=2.035 $X2=0
+ $Y2=0
cc_147 N_A_71_368#_c_189_n N_VPWR_c_263_n 0.026688f $X=2.4 $Y=2.815 $X2=0 $Y2=0
cc_148 N_A_71_368#_c_186_n N_VPWR_c_264_n 0.0593439f $X=1.215 $Y=2.99 $X2=0
+ $Y2=0
cc_149 N_A_71_368#_c_187_n N_VPWR_c_264_n 0.0235512f $X=0.645 $Y=2.99 $X2=0
+ $Y2=0
cc_150 N_A_71_368#_c_189_n N_VPWR_c_266_n 0.014549f $X=2.4 $Y=2.815 $X2=0 $Y2=0
cc_151 N_A_71_368#_c_186_n N_VPWR_c_262_n 0.032751f $X=1.215 $Y=2.99 $X2=0 $Y2=0
cc_152 N_A_71_368#_c_187_n N_VPWR_c_262_n 0.0126924f $X=0.645 $Y=2.99 $X2=0
+ $Y2=0
cc_153 N_A_71_368#_c_189_n N_VPWR_c_262_n 0.0119743f $X=2.4 $Y=2.815 $X2=0 $Y2=0
cc_154 N_Y_c_227_n N_VGND_c_290_n 0.0019893f $X=0.835 $Y=1.095 $X2=0 $Y2=0
cc_155 N_Y_c_228_n N_VGND_c_290_n 0.0167629f $X=1.35 $Y=0.515 $X2=0 $Y2=0
cc_156 N_Y_c_226_n N_VGND_c_291_n 0.00316703f $X=1.13 $Y=1.095 $X2=0 $Y2=0
cc_157 N_Y_c_228_n N_VGND_c_291_n 0.0167858f $X=1.35 $Y=0.515 $X2=0 $Y2=0
cc_158 N_Y_c_228_n N_VGND_c_294_n 0.0194005f $X=1.35 $Y=0.515 $X2=0 $Y2=0
cc_159 N_Y_c_228_n N_VGND_c_297_n 0.0159453f $X=1.35 $Y=0.515 $X2=0 $Y2=0
cc_160 N_Y_c_226_n A_159_74# 0.00366293f $X=1.13 $Y=1.095 $X2=-0.19 $Y2=-0.245

* File: sky130_fd_sc_ms__o221a_1.spice
* Created: Wed Sep  2 12:22:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o221a_1.pex.spice"
.subckt sky130_fd_sc_ms__o221a_1  VNB VPB A1 A2 B2 B1 C1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* C1	C1
* B1	B1
* B2	B2
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_83_264#_M1004_g N_X_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.166607 AS=0.2109 PD=1.25478 PS=2.05 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1003 N_A_245_94#_M1003_d N_A1_M1003_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.112 AS=0.144093 PD=0.99 PS=1.08522 NRD=0 NRS=15.468 M=1 R=4.26667
+ SA=75000.8 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_245_94#_M1003_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.112 PD=1.85 PS=0.99 NRD=0 NRS=13.116 M=1 R=4.26667 SA=75001.3
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_A_245_94#_M1001_d N_B2_M1001_g N_A_456_74#_M1001_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.2336 PD=0.92 PS=2.01 NRD=0 NRS=7.488 M=1 R=4.26667
+ SA=75000.3 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1008 N_A_456_74#_M1008_d N_B1_M1008_g N_A_245_94#_M1001_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.112 AS=0.0896 PD=0.99 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1006 N_A_83_264#_M1006_d N_C1_M1006_g N_A_456_74#_M1008_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.2944 AS=0.112 PD=2.2 PS=0.99 NRD=13.116 NRS=0 M=1 R=4.26667
+ SA=75001.2 SB=75000.4 A=0.096 P=1.58 MULT=1
MM1007 N_VPWR_M1007_d N_A_83_264#_M1007_g N_X_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.311698 AS=0.3136 PD=1.77509 PS=2.8 NRD=23.7385 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90003.1 A=0.2016 P=2.6 MULT=1
MM1010 A_267_392# N_A1_M1010_g N_VPWR_M1007_d VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.278302 PD=1.24 PS=1.58491 NRD=12.7853 NRS=28.565 M=1 R=5.55556 SA=90000.9
+ SB=90002.8 A=0.18 P=2.36 MULT=1
MM1002 N_A_83_264#_M1002_d N_A2_M1002_g A_267_392# VPB PSHORT L=0.18 W=1
+ AD=0.195 AS=0.12 PD=1.39 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556 SA=90001.3
+ SB=90002.3 A=0.18 P=2.36 MULT=1
MM1011 A_465_392# N_B2_M1011_g N_A_83_264#_M1002_d VPB PSHORT L=0.18 W=1
+ AD=0.195 AS=0.195 PD=1.39 PS=1.39 NRD=27.5603 NRS=22.6353 M=1 R=5.55556
+ SA=90001.9 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_B1_M1005_g A_465_392# VPB PSHORT L=0.18 W=1 AD=0.415
+ AS=0.195 PD=1.83 PS=1.39 NRD=0 NRS=27.5603 M=1 R=5.55556 SA=90002.5 SB=90001.2
+ A=0.18 P=2.36 MULT=1
MM1009 N_A_83_264#_M1009_d N_C1_M1009_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=1
+ AD=0.28 AS=0.415 PD=2.56 PS=1.83 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90003.5
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.742 P=13.12
c_44 VNB 0 1.2498e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__o221a_1.pxi.spice"
*
.ends
*
*

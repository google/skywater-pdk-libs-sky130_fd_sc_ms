* File: sky130_fd_sc_ms__or2_1.pxi.spice
* Created: Wed Sep  2 12:27:30 2020
* 
x_PM_SKY130_FD_SC_MS__OR2_1%B N_B_M1001_g N_B_c_44_n N_B_M1003_g B N_B_c_45_n
+ N_B_c_46_n PM_SKY130_FD_SC_MS__OR2_1%B
x_PM_SKY130_FD_SC_MS__OR2_1%A N_A_M1005_g N_A_M1002_g A N_A_c_71_n N_A_c_72_n
+ PM_SKY130_FD_SC_MS__OR2_1%A
x_PM_SKY130_FD_SC_MS__OR2_1%A_63_368# N_A_63_368#_M1003_d N_A_63_368#_M1001_s
+ N_A_63_368#_M1004_g N_A_63_368#_M1000_g N_A_63_368#_c_121_n
+ N_A_63_368#_c_112_n N_A_63_368#_c_113_n N_A_63_368#_c_114_n
+ N_A_63_368#_c_115_n N_A_63_368#_c_116_n N_A_63_368#_c_120_n
+ N_A_63_368#_c_117_n PM_SKY130_FD_SC_MS__OR2_1%A_63_368#
x_PM_SKY130_FD_SC_MS__OR2_1%VPWR N_VPWR_M1005_d N_VPWR_c_184_n VPWR
+ N_VPWR_c_185_n N_VPWR_c_186_n N_VPWR_c_183_n N_VPWR_c_188_n
+ PM_SKY130_FD_SC_MS__OR2_1%VPWR
x_PM_SKY130_FD_SC_MS__OR2_1%X N_X_M1000_d N_X_M1004_d N_X_c_208_n N_X_c_209_n X
+ X X X N_X_c_210_n PM_SKY130_FD_SC_MS__OR2_1%X
x_PM_SKY130_FD_SC_MS__OR2_1%VGND N_VGND_M1003_s N_VGND_M1002_d N_VGND_c_233_n
+ N_VGND_c_234_n N_VGND_c_235_n N_VGND_c_236_n VGND N_VGND_c_237_n
+ N_VGND_c_238_n N_VGND_c_239_n N_VGND_c_240_n PM_SKY130_FD_SC_MS__OR2_1%VGND
cc_1 VNB N_B_M1001_g 0.00922557f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=2.26
cc_2 VNB N_B_c_44_n 0.0221254f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.22
cc_3 VNB N_B_c_45_n 0.0701489f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_4 VNB N_B_c_46_n 0.0293162f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_5 VNB N_A_M1002_g 0.027266f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.22
cc_6 VNB N_A_c_71_n 0.030309f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_7 VNB N_A_c_72_n 0.00189714f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_8 VNB N_A_63_368#_M1004_g 0.00187335f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.835
cc_9 VNB N_A_63_368#_M1000_g 0.0286452f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_10 VNB N_A_63_368#_c_112_n 0.0038832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_63_368#_c_113_n 0.00741821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_63_368#_c_114_n 0.00541617f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_63_368#_c_115_n 0.00770034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_63_368#_c_116_n 4.1382e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_63_368#_c_117_n 0.0340765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_183_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.365
cc_17 VNB N_X_c_208_n 0.0265168f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.835
cc_18 VNB N_X_c_209_n 0.0133911f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_19 VNB N_X_c_210_n 0.0246392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_233_n 0.0267471f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.835
cc_21 VNB N_VGND_c_234_n 0.0168543f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.385
cc_22 VNB N_VGND_c_235_n 0.0115308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_236_n 0.00682834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_237_n 0.0239783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_238_n 0.0189562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_239_n 0.177517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_240_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VPB N_B_M1001_g 0.0311086f $X=-0.19 $Y=1.66 $X2=0.685 $Y2=2.26
cc_29 VPB N_A_M1005_g 0.0230515f $X=-0.19 $Y=1.66 $X2=0.685 $Y2=1.55
cc_30 VPB N_A_c_71_n 0.0074916f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_31 VPB N_A_c_72_n 0.0024512f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_32 VPB N_A_63_368#_M1004_g 0.0309948f $X=-0.19 $Y=1.66 $X2=0.7 $Y2=0.835
cc_33 VPB N_A_63_368#_c_116_n 0.00317467f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_34 VPB N_A_63_368#_c_120_n 0.0403242f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_184_n 0.0226065f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_185_n 0.0377411f $X=-0.19 $Y=1.66 $X2=0.155 $Y2=1.21
cc_37 VPB N_VPWR_c_186_n 0.0189562f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_183_n 0.0741763f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.365
cc_39 VPB N_VPWR_c_188_n 0.0118997f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB X 0.0133306f $X=-0.19 $Y=1.66 $X2=0.61 $Y2=1.385
cc_41 VPB X 0.0413779f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_X_c_210_n 0.0074668f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_43 N_B_M1001_g N_A_M1005_g 0.0344424f $X=0.685 $Y=2.26 $X2=0 $Y2=0
cc_44 N_B_c_44_n N_A_M1002_g 0.0135545f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_45 N_B_c_46_n N_A_M1002_g 9.09937e-19 $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_46 N_B_c_45_n N_A_c_71_n 0.042824f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_47 N_B_c_46_n N_A_c_71_n 7.73509e-19 $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_48 N_B_c_45_n N_A_c_72_n 0.00166706f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_49 N_B_c_46_n N_A_c_72_n 0.0109438f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_50 N_B_M1001_g N_A_63_368#_c_121_n 0.0139236f $X=0.685 $Y=2.26 $X2=0 $Y2=0
cc_51 N_B_c_46_n N_A_63_368#_c_121_n 0.00540887f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_52 N_B_c_44_n N_A_63_368#_c_112_n 0.00461704f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_53 N_B_c_44_n N_A_63_368#_c_114_n 0.00500991f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_54 N_B_M1001_g N_A_63_368#_c_120_n 0.0186809f $X=0.685 $Y=2.26 $X2=0 $Y2=0
cc_55 N_B_c_45_n N_A_63_368#_c_120_n 0.00659078f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_56 N_B_c_46_n N_A_63_368#_c_120_n 0.0197016f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_57 N_B_M1001_g N_VPWR_c_184_n 0.00168079f $X=0.685 $Y=2.26 $X2=0 $Y2=0
cc_58 N_B_M1001_g N_VPWR_c_185_n 0.00465228f $X=0.685 $Y=2.26 $X2=0 $Y2=0
cc_59 N_B_M1001_g N_VPWR_c_183_n 0.00555093f $X=0.685 $Y=2.26 $X2=0 $Y2=0
cc_60 N_B_c_44_n N_VGND_c_233_n 0.0135644f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_61 N_B_c_45_n N_VGND_c_233_n 0.00215303f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_62 N_B_c_46_n N_VGND_c_233_n 0.0264066f $X=0.61 $Y=1.385 $X2=0 $Y2=0
cc_63 N_B_c_44_n N_VGND_c_237_n 0.00375057f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_64 N_B_c_44_n N_VGND_c_239_n 0.00409726f $X=0.7 $Y=1.22 $X2=0 $Y2=0
cc_65 N_A_M1005_g N_A_63_368#_M1004_g 0.00934911f $X=1.105 $Y=2.26 $X2=0 $Y2=0
cc_66 N_A_c_71_n N_A_63_368#_M1004_g 0.00112359f $X=1.21 $Y=1.515 $X2=0 $Y2=0
cc_67 N_A_M1002_g N_A_63_368#_M1000_g 0.0176009f $X=1.325 $Y=0.835 $X2=0 $Y2=0
cc_68 N_A_M1005_g N_A_63_368#_c_121_n 0.0181138f $X=1.105 $Y=2.26 $X2=0 $Y2=0
cc_69 N_A_c_71_n N_A_63_368#_c_121_n 0.00183271f $X=1.21 $Y=1.515 $X2=0 $Y2=0
cc_70 N_A_c_72_n N_A_63_368#_c_121_n 0.0231721f $X=1.21 $Y=1.515 $X2=0 $Y2=0
cc_71 N_A_M1002_g N_A_63_368#_c_112_n 6.93808e-19 $X=1.325 $Y=0.835 $X2=0 $Y2=0
cc_72 N_A_M1002_g N_A_63_368#_c_113_n 0.0162525f $X=1.325 $Y=0.835 $X2=0 $Y2=0
cc_73 N_A_c_72_n N_A_63_368#_c_113_n 0.00982684f $X=1.21 $Y=1.515 $X2=0 $Y2=0
cc_74 N_A_c_71_n N_A_63_368#_c_114_n 0.00268859f $X=1.21 $Y=1.515 $X2=0 $Y2=0
cc_75 N_A_c_72_n N_A_63_368#_c_114_n 0.0166608f $X=1.21 $Y=1.515 $X2=0 $Y2=0
cc_76 N_A_M1002_g N_A_63_368#_c_115_n 0.00546476f $X=1.325 $Y=0.835 $X2=0 $Y2=0
cc_77 N_A_c_72_n N_A_63_368#_c_115_n 0.0172973f $X=1.21 $Y=1.515 $X2=0 $Y2=0
cc_78 N_A_M1005_g N_A_63_368#_c_116_n 0.00325935f $X=1.105 $Y=2.26 $X2=0 $Y2=0
cc_79 N_A_c_71_n N_A_63_368#_c_116_n 3.97332e-19 $X=1.21 $Y=1.515 $X2=0 $Y2=0
cc_80 N_A_c_72_n N_A_63_368#_c_116_n 0.00910636f $X=1.21 $Y=1.515 $X2=0 $Y2=0
cc_81 N_A_M1005_g N_A_63_368#_c_120_n 0.00260222f $X=1.105 $Y=2.26 $X2=0 $Y2=0
cc_82 N_A_M1002_g N_A_63_368#_c_117_n 0.0174761f $X=1.325 $Y=0.835 $X2=0 $Y2=0
cc_83 N_A_c_72_n N_A_63_368#_c_117_n 3.285e-19 $X=1.21 $Y=1.515 $X2=0 $Y2=0
cc_84 N_A_M1005_g N_VPWR_c_184_n 0.0154658f $X=1.105 $Y=2.26 $X2=0 $Y2=0
cc_85 N_A_M1005_g N_VPWR_c_185_n 0.00401533f $X=1.105 $Y=2.26 $X2=0 $Y2=0
cc_86 N_A_M1005_g N_VPWR_c_183_n 0.00465661f $X=1.105 $Y=2.26 $X2=0 $Y2=0
cc_87 N_A_M1002_g N_X_c_208_n 8.51118e-19 $X=1.325 $Y=0.835 $X2=0 $Y2=0
cc_88 N_A_M1002_g N_VGND_c_233_n 6.19635e-19 $X=1.325 $Y=0.835 $X2=0 $Y2=0
cc_89 N_A_M1002_g N_VGND_c_234_n 0.00508306f $X=1.325 $Y=0.835 $X2=0 $Y2=0
cc_90 N_A_M1002_g N_VGND_c_237_n 0.00451272f $X=1.325 $Y=0.835 $X2=0 $Y2=0
cc_91 N_A_M1002_g N_VGND_c_239_n 0.00487769f $X=1.325 $Y=0.835 $X2=0 $Y2=0
cc_92 N_A_63_368#_c_121_n A_155_368# 0.0096152f $X=1.615 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_93 N_A_63_368#_c_121_n N_VPWR_M1005_d 0.0183317f $X=1.615 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_94 N_A_63_368#_c_116_n N_VPWR_M1005_d 0.0023593f $X=1.7 $Y=1.95 $X2=-0.19
+ $Y2=-0.245
cc_95 N_A_63_368#_M1004_g N_VPWR_c_184_n 0.0057523f $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_96 N_A_63_368#_c_121_n N_VPWR_c_184_n 0.0436101f $X=1.615 $Y=2.035 $X2=0
+ $Y2=0
cc_97 N_A_63_368#_c_120_n N_VPWR_c_184_n 0.0125255f $X=0.46 $Y=1.985 $X2=0 $Y2=0
cc_98 N_A_63_368#_c_117_n N_VPWR_c_184_n 3.89356e-19 $X=1.805 $Y=1.465 $X2=0
+ $Y2=0
cc_99 N_A_63_368#_c_120_n N_VPWR_c_185_n 0.0066444f $X=0.46 $Y=1.985 $X2=0 $Y2=0
cc_100 N_A_63_368#_M1004_g N_VPWR_c_186_n 0.005209f $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_101 N_A_63_368#_M1004_g N_VPWR_c_183_n 0.00990469f $X=1.895 $Y=2.4 $X2=0
+ $Y2=0
cc_102 N_A_63_368#_c_120_n N_VPWR_c_183_n 0.00995531f $X=0.46 $Y=1.985 $X2=0
+ $Y2=0
cc_103 N_A_63_368#_M1000_g N_X_c_208_n 0.00926861f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_104 N_A_63_368#_M1000_g N_X_c_209_n 0.00352004f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A_63_368#_c_115_n N_X_c_209_n 0.00658407f $X=1.7 $Y=1.63 $X2=0 $Y2=0
cc_106 N_A_63_368#_c_117_n N_X_c_209_n 2.41927e-19 $X=1.805 $Y=1.465 $X2=0 $Y2=0
cc_107 N_A_63_368#_M1004_g X 0.00344691f $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_108 N_A_63_368#_c_115_n X 0.00102654f $X=1.7 $Y=1.63 $X2=0 $Y2=0
cc_109 N_A_63_368#_c_116_n X 0.00564757f $X=1.7 $Y=1.95 $X2=0 $Y2=0
cc_110 N_A_63_368#_M1004_g X 0.0188008f $X=1.895 $Y=2.4 $X2=0 $Y2=0
cc_111 N_A_63_368#_M1000_g N_X_c_210_n 0.00255066f $X=1.905 $Y=0.74 $X2=0 $Y2=0
cc_112 N_A_63_368#_c_115_n N_X_c_210_n 0.0304892f $X=1.7 $Y=1.63 $X2=0 $Y2=0
cc_113 N_A_63_368#_c_116_n N_X_c_210_n 0.00628992f $X=1.7 $Y=1.95 $X2=0 $Y2=0
cc_114 N_A_63_368#_c_117_n N_X_c_210_n 0.0106954f $X=1.805 $Y=1.465 $X2=0 $Y2=0
cc_115 N_A_63_368#_c_113_n N_VGND_M1002_d 0.00185525f $X=1.615 $Y=1.095 $X2=0
+ $Y2=0
cc_116 N_A_63_368#_c_115_n N_VGND_M1002_d 0.002623f $X=1.7 $Y=1.63 $X2=0 $Y2=0
cc_117 N_A_63_368#_c_112_n N_VGND_c_233_n 0.0231039f $X=1.075 $Y=0.82 $X2=0
+ $Y2=0
cc_118 N_A_63_368#_M1000_g N_VGND_c_234_n 0.00879154f $X=1.905 $Y=0.74 $X2=0
+ $Y2=0
cc_119 N_A_63_368#_c_112_n N_VGND_c_234_n 0.00132933f $X=1.075 $Y=0.82 $X2=0
+ $Y2=0
cc_120 N_A_63_368#_c_113_n N_VGND_c_234_n 0.0128182f $X=1.615 $Y=1.095 $X2=0
+ $Y2=0
cc_121 N_A_63_368#_c_115_n N_VGND_c_234_n 0.0142456f $X=1.7 $Y=1.63 $X2=0 $Y2=0
cc_122 N_A_63_368#_c_117_n N_VGND_c_234_n 5.87857e-19 $X=1.805 $Y=1.465 $X2=0
+ $Y2=0
cc_123 N_A_63_368#_c_112_n N_VGND_c_237_n 0.00729875f $X=1.075 $Y=0.82 $X2=0
+ $Y2=0
cc_124 N_A_63_368#_M1000_g N_VGND_c_238_n 0.00434272f $X=1.905 $Y=0.74 $X2=0
+ $Y2=0
cc_125 N_A_63_368#_M1000_g N_VGND_c_239_n 0.00828717f $X=1.905 $Y=0.74 $X2=0
+ $Y2=0
cc_126 N_A_63_368#_c_112_n N_VGND_c_239_n 0.00950289f $X=1.075 $Y=0.82 $X2=0
+ $Y2=0
cc_127 N_VPWR_c_184_n X 0.0270509f $X=1.67 $Y=2.455 $X2=0 $Y2=0
cc_128 N_VPWR_c_186_n X 0.0156645f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_129 N_VPWR_c_183_n X 0.0128976f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_130 N_X_c_208_n N_VGND_c_234_n 0.0193831f $X=2.12 $Y=0.515 $X2=0 $Y2=0
cc_131 N_X_c_208_n N_VGND_c_238_n 0.0156794f $X=2.12 $Y=0.515 $X2=0 $Y2=0
cc_132 N_X_c_208_n N_VGND_c_239_n 0.0129217f $X=2.12 $Y=0.515 $X2=0 $Y2=0

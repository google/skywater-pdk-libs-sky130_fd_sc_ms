* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__o2bb2ai_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 VPWR A1_N a_136_387# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X1 a_136_387# A2_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X2 a_518_74# B2 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X3 VGND B2 a_518_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 a_799_368# B2 Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X5 a_134_74# A2_N a_136_387# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X6 VGND B1 a_518_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 VGND A1_N a_134_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X8 a_518_74# B1 VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X9 VPWR A2_N a_136_387# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X10 a_136_387# A1_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X11 Y a_136_387# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X12 VPWR a_136_387# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X13 a_518_74# a_136_387# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X14 VPWR B1 a_799_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X15 Y B2 a_799_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X16 a_134_74# A1_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X17 Y a_136_387# a_518_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X18 a_799_368# B1 VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X19 a_136_387# A2_N a_134_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
.ends

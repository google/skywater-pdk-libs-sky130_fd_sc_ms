* File: sky130_fd_sc_ms__sdfbbn_2.spice
* Created: Wed Sep  2 12:29:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdfbbn_2.pex.spice"
.subckt sky130_fd_sc_ms__sdfbbn_2  VNB VPB SCD D SCE CLK_N SET_B RESET_B VPWR
+ Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* CLK_N	CLK_N
* SCE	SCE
* D	D
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1008 A_119_119# N_SCD_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1037 N_A_197_119#_M1037_d N_SCE_M1037_g A_119_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1428 AS=0.0504 PD=1.1 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1044 A_363_119# N_D_M1044_g N_A_197_119#_M1037_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1428 PD=0.66 PS=1.1 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1028 N_VGND_M1028_d N_A_341_410#_M1028_g A_363_119# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0504 PD=0.95 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.8
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1039 N_A_341_410#_M1039_d N_SCE_M1039_g N_VGND_M1028_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.1113 PD=1.41 PS=0.95 NRD=0 NRS=71.424 M=1 R=2.8
+ SA=75002.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1038 N_VGND_M1038_d N_CLK_N_M1038_g N_A_688_98#_M1038_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.30025 AS=0.2109 PD=1.74 PS=2.05 NRD=56.868 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1046 N_A_871_368#_M1046_d N_A_688_98#_M1046_g N_VGND_M1038_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.30025 PD=2.05 PS=1.74 NRD=0 NRS=56.868 M=1 R=4.93333
+ SA=75001.1 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1031 A_1185_125# N_A_1007_366#_M1031_g N_VGND_M1031_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.24385 PD=0.63 PS=2.14 NRD=14.28 NRS=150.168 M=1 R=2.8
+ SA=75000.3 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1016 N_A_1157_464#_M1016_d N_A_688_98#_M1016_g A_1185_125# VNB NLOWVT L=0.15
+ W=0.42 AD=0.06405 AS=0.0441 PD=0.725 PS=0.63 NRD=7.14 NRS=14.28 M=1 R=2.8
+ SA=75000.7 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1009 N_A_197_119#_M1009_d N_A_871_368#_M1009_g N_A_1157_464#_M1016_d VNB
+ NLOWVT L=0.15 W=0.42 AD=0.1491 AS=0.06405 PD=1.55 PS=0.725 NRD=19.992 NRS=0
+ M=1 R=2.8 SA=75001.1 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1019 N_A_1007_366#_M1019_d N_A_1157_464#_M1019_g N_A_1473_73#_M1019_s VNB
+ NLOWVT L=0.15 W=0.55 AD=0.077 AS=0.3531 PD=0.83 PS=2.54 NRD=0 NRS=128.064 M=1
+ R=3.66667 SA=75000.4 SB=75003.2 A=0.0825 P=1.4 MULT=1
MM1020 N_A_1473_73#_M1020_d N_A_1643_257#_M1020_g N_A_1007_366#_M1019_d VNB
+ NLOWVT L=0.15 W=0.55 AD=0.125125 AS=0.077 PD=1.005 PS=0.83 NRD=26.172 NRS=0
+ M=1 R=3.66667 SA=75000.8 SB=75002.8 A=0.0825 P=1.4 MULT=1
MM1051 N_VGND_M1051_d N_SET_B_M1051_g N_A_1473_73#_M1020_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.09625 AS=0.125125 PD=0.9 PS=1.005 NRD=15.264 NRS=11.988 M=1
+ R=3.66667 SA=75001.4 SB=75002.2 A=0.0825 P=1.4 MULT=1
MM1049 A_1902_125# N_A_1007_366#_M1049_g N_VGND_M1051_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.108187 AS=0.09625 PD=1.09 PS=0.9 NRD=30.912 NRS=0 M=1 R=3.66667
+ SA=75001.9 SB=75001.7 A=0.0825 P=1.4 MULT=1
MM1023 N_A_1997_82#_M1023_d N_A_688_98#_M1023_g A_1902_125# VNB NLOWVT L=0.15
+ W=0.55 AD=0.280387 AS=0.108187 PD=1.87113 PS=1.09 NRD=0 NRS=30.912 M=1
+ R=3.66667 SA=75001.5 SB=75002.7 A=0.0825 P=1.4 MULT=1
MM1015 A_2247_82# N_A_871_368#_M1015_g N_A_1997_82#_M1023_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.214113 PD=0.66 PS=1.42887 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75002.5 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1047 N_VGND_M1047_d N_A_2216_410#_M1047_g A_2247_82# VNB NLOWVT L=0.15 W=0.42
+ AD=0.125656 AS=0.0504 PD=1.01017 PS=0.66 NRD=30 NRS=18.564 M=1 R=2.8
+ SA=75002.9 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1006 N_A_2452_74#_M1006_d N_SET_B_M1006_g N_VGND_M1047_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1369 AS=0.221394 PD=1.11 PS=1.77983 NRD=0 NRS=39.588 M=1 R=4.93333
+ SA=75002.1 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1041 N_A_2216_410#_M1041_d N_A_1643_257#_M1041_g N_A_2452_74#_M1006_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.1036 AS=0.1369 PD=1.02 PS=1.11 NRD=0 NRS=7.296 M=1
+ R=4.93333 SA=75002.6 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1011 N_A_2452_74#_M1011_d N_A_1997_82#_M1011_g N_A_2216_410#_M1041_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.30055 AS=0.1036 PD=2.42 PS=1.02 NRD=13.776 NRS=0 M=1
+ R=4.93333 SA=75003 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1010 N_VGND_M1010_d N_RESET_B_M1010_g N_A_1643_257#_M1010_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.136772 AS=0.1176 PD=1.32517 PS=1.4 NRD=172.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1010_d N_A_2216_410#_M1007_g N_Q_N_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.240978 AS=0.1036 PD=2.33483 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.5 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1024 N_VGND_M1024_d N_A_2216_410#_M1024_g N_Q_N_M1007_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2294 AS=0.1036 PD=2.1 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.9
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1021_d N_A_2216_410#_M1021_g N_A_3272_94#_M1021_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.150029 AS=0.1824 PD=1.10377 PS=1.85 NRD=19.212 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1025 N_Q_M1025_d N_A_3272_94#_M1025_g N_VGND_M1021_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.173471 PD=1.02 PS=1.27623 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1043 N_Q_M1025_d N_A_3272_94#_M1043_g N_VGND_M1043_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2072 PD=1.02 PS=2.04 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.2
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1012 N_VPWR_M1012_d N_SCD_M1012_g N_A_27_464#_M1012_s VPB PSHORT L=0.18 W=0.64
+ AD=0.0864 AS=0.1792 PD=0.91 PS=1.84 NRD=0 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90001.5 A=0.1152 P=1.64 MULT=1
MM1013 A_209_464# N_SCE_M1013_g N_VPWR_M1012_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0672 AS=0.0864 PD=0.85 PS=0.91 NRD=15.3857 NRS=0 M=1 R=3.55556 SA=90000.6
+ SB=90001 A=0.1152 P=1.64 MULT=1
MM1042 N_A_197_119#_M1042_d N_D_M1042_g A_209_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.0864 AS=0.0672 PD=0.91 PS=0.85 NRD=0 NRS=15.3857 M=1 R=3.55556 SA=90001
+ SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1045 N_A_27_464#_M1045_d N_A_341_410#_M1045_g N_A_197_119#_M1042_d VPB PSHORT
+ L=0.18 W=0.64 AD=0.1792 AS=0.0864 PD=1.84 PS=0.91 NRD=0 NRS=0 M=1 R=3.55556
+ SA=90001.5 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1017 N_A_341_410#_M1017_d N_SCE_M1017_g N_VPWR_M1017_s VPB PSHORT L=0.18
+ W=0.64 AD=0.1792 AS=0.1792 PD=1.84 PS=1.84 NRD=0 NRS=0 M=1 R=3.55556
+ SA=90000.2 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1048 N_VPWR_M1048_d N_CLK_N_M1048_g N_A_688_98#_M1048_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1001 N_A_871_368#_M1001_d N_A_688_98#_M1001_g N_VPWR_M1048_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.1512 PD=2.8 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1030 A_1073_464# N_A_1007_366#_M1030_g N_VPWR_M1030_s VPB PSHORT L=0.18 W=0.42
+ AD=0.0504 AS=0.1176 PD=0.66 PS=1.4 NRD=30.4759 NRS=0 M=1 R=2.33333 SA=90000.2
+ SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1003 N_A_1157_464#_M1003_d N_A_871_368#_M1003_g A_1073_464# VPB PSHORT L=0.18
+ W=0.42 AD=0.0834849 AS=0.0504 PD=0.788491 PS=0.66 NRD=37.5088 NRS=30.4759 M=1
+ R=2.33333 SA=90000.6 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1018 N_A_197_119#_M1018_d N_A_688_98#_M1018_g N_A_1157_464#_M1003_d VPB PSHORT
+ L=0.18 W=0.64 AD=0.2112 AS=0.127215 PD=1.94 PS=1.20151 NRD=13.8491 NRS=0 M=1
+ R=3.55556 SA=90000.8 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1004 A_1595_424# N_A_1157_464#_M1004_g N_A_1007_366#_M1004_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1008 AS=0.735 PD=1.08 PS=3.43 NRD=15.2281 NRS=0 M=1 R=4.66667
+ SA=90000.8 SB=90001.1 A=0.1512 P=2.04 MULT=1
MM1033 N_VPWR_M1033_d N_A_1643_257#_M1033_g A_1595_424# VPB PSHORT L=0.18 W=0.84
+ AD=0.1512 AS=0.1008 PD=1.2 PS=1.08 NRD=0 NRS=15.2281 M=1 R=4.66667 SA=90001.2
+ SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1050 N_A_1007_366#_M1050_d N_SET_B_M1050_g N_VPWR_M1033_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.1512 PD=2.24 PS=1.2 NRD=0 NRS=19.9167 M=1 R=4.66667
+ SA=90001.7 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1022 A_1989_424# N_A_1007_366#_M1022_g N_VPWR_M1022_s VPB PSHORT L=0.18 W=0.84
+ AD=0.0882 AS=0.2352 PD=1.05 PS=2.24 NRD=11.7215 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90001 A=0.1512 P=2.04 MULT=1
MM1027 N_A_1997_82#_M1027_d N_A_871_368#_M1027_g A_1989_424# VPB PSHORT L=0.18
+ W=0.84 AD=0.1778 AS=0.0882 PD=1.59333 PS=1.05 NRD=0 NRS=11.7215 M=1 R=4.66667
+ SA=90000.6 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1002 A_2174_508# N_A_688_98#_M1002_g N_A_1997_82#_M1027_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0441 AS=0.0889 PD=0.63 PS=0.796667 NRD=23.443 NRS=37.5088 M=1
+ R=2.33333 SA=90001.1 SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1036 N_VPWR_M1036_d N_A_2216_410#_M1036_g A_2174_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.1176 AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.33333 SA=90001.5
+ SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1005 N_VPWR_M1005_d N_SET_B_M1005_g N_A_2216_410#_M1005_s VPB PSHORT L=0.18
+ W=1 AD=0.165 AS=0.28 PD=1.33 PS=2.56 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1034 A_2559_392# N_A_1643_257#_M1034_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.165 PD=1.24 PS=1.33 NRD=12.7853 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1040 N_A_2216_410#_M1040_d N_A_1997_82#_M1040_g A_2559_392# VPB PSHORT L=0.18
+ W=1 AD=0.28 AS=0.12 PD=2.56 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556 SA=90001.1
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_RESET_B_M1000_g N_A_1643_257#_M1000_s VPB PSHORT L=0.18
+ W=0.64 AD=0.416409 AS=0.1792 PD=1.68364 PS=1.84 NRD=197.768 NRS=0 M=1
+ R=3.55556 SA=90000.2 SB=90001.8 A=0.1152 P=1.64 MULT=1
MM1026 N_Q_N_M1026_d N_A_2216_410#_M1026_g N_VPWR_M1000_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.728716 PD=1.39 PS=2.94636 NRD=0 NRS=14.3613 M=1
+ R=6.22222 SA=90001 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1032 N_Q_N_M1026_d N_A_2216_410#_M1032_g N_VPWR_M1032_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3024 PD=1.39 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.5 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1014 N_VPWR_M1014_d N_A_2216_410#_M1014_g N_A_3272_94#_M1014_s VPB PSHORT
+ L=0.18 W=1 AD=0.177264 AS=0.275 PD=1.38208 PS=2.55 NRD=13.7703 NRS=0 M=1
+ R=5.55556 SA=90000.2 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1029 N_Q_M1029_d N_A_3272_94#_M1029_g N_VPWR_M1014_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.198536 PD=1.39 PS=1.54792 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.7
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1035 N_Q_M1029_d N_A_3272_94#_M1035_g N_VPWR_M1035_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX52_noxref VNB VPB NWDIODE A=34.6332 P=40.96
c_199 VNB 0 3.69273e-19 $X=0 $Y=0
c_378 VPB 0 5.99464e-20 $X=0 $Y=3.085
c_2893 A_1185_125# 0 1.91291e-19 $X=5.925 $Y=0.625
c_2937 A_1902_125# 0 7.74904e-20 $X=9.51 $Y=0.625
*
.include "sky130_fd_sc_ms__sdfbbn_2.pxi.spice"
*
.ends
*
*

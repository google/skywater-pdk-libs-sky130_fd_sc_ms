* File: sky130_fd_sc_ms__a21bo_1.spice
* Created: Wed Sep  2 11:50:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__a21bo_1.pex.spice"
.subckt sky130_fd_sc_ms__a21bo_1  VNB VPB A2 A1 B1_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1_N	B1_N
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1002 A_122_136# N_A2_M1002_g N_VGND_M1002_s VNB NLOWVT L=0.15 W=0.64 AD=0.0672
+ AS=0.1696 PD=0.85 PS=1.81 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2 SB=75001.1
+ A=0.096 P=1.58 MULT=1
MM1009 N_A_194_136#_M1009_d N_A1_M1009_g A_122_136# VNB NLOWVT L=0.15 W=0.64
+ AD=0.1248 AS=0.0672 PD=1.03 PS=0.85 NRD=3.744 NRS=9.372 M=1 R=4.26667
+ SA=75000.6 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1004 N_VGND_M1004_d N_A_272_110#_M1004_g N_A_194_136#_M1009_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.1248 PD=1.81 PS=1.03 NRD=0 NRS=16.872 M=1
+ R=4.26667 SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 N_VGND_M1008_d N_B1_N_M1008_g N_A_272_110#_M1008_s VNB NLOWVT L=0.15
+ W=0.55 AD=0.0964632 AS=0.15675 PD=0.90814 PS=1.67 NRD=4.356 NRS=0 M=1
+ R=3.66667 SA=75000.2 SB=75000.7 A=0.0825 P=1.4 MULT=1
MM1003 N_X_M1003_d N_A_194_136#_M1003_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.129787 PD=2.01 PS=1.22186 NRD=0 NRS=4.044 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_VPWR_M1006_d N_A2_M1006_g N_A_34_392#_M1006_s VPB PSHORT L=0.18 W=1
+ AD=0.15 AS=0.26 PD=1.3 PS=2.52 NRD=1.9503 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1000 N_A_34_392#_M1000_d N_A1_M1000_g N_VPWR_M1006_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.15 PD=1.27 PS=1.3 NRD=0 NRS=1.9503 M=1 R=5.55556 SA=90000.6
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1005 N_A_194_136#_M1005_d N_A_272_110#_M1005_g N_A_34_392#_M1000_d VPB PSHORT
+ L=0.18 W=1 AD=0.26 AS=0.135 PD=2.52 PS=1.27 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90001.1 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_B1_N_M1007_g N_A_272_110#_M1007_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1614 AS=0.2184 PD=1.26429 PS=2.2 NRD=32.1504 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1001 N_X_M1001_d N_A_194_136#_M1001_g N_VPWR_M1007_d VPB PSHORT L=0.18 W=1.12
+ AD=0.2912 AS=0.2152 PD=2.76 PS=1.68571 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8492 P=12.16
c_44 VNB 0 9.10919e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__a21bo_1.pxi.spice"
*
.ends
*
*

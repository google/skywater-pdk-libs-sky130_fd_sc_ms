* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfxtp_4 CLK D SCD SCE VGND VNB VPB VPWR Q
M1000 VPWR SCD a_415_464# VPB pshort w=640000u l=180000u
+  ad=2.83978e+12p pd=2.238e+07u as=2.304e+11p ps=2e+06u
M1001 a_630_74# CLK VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1002 a_1026_100# a_828_74# a_301_74# VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=2.904e+11p ps=3.22e+06u
M1003 a_630_74# CLK VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=1.77695e+12p ps=1.604e+07u
M1004 VGND a_1814_48# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=4.773e+11p ps=4.25e+06u
M1005 Q a_1814_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1006 a_1217_506# a_630_74# a_1026_100# VPB pshort w=420000u l=180000u
+  ad=1.512e+11p pd=1.56e+06u as=0p ps=0u
M1007 VPWR a_1814_48# a_1767_476# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1008 VPWR a_1587_74# a_1814_48# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.268e+11p ps=2.22e+06u
M1009 VPWR a_1257_74# a_1217_506# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND SCD a_452_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1011 a_452_74# SCE a_301_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=3.738e+11p ps=3.46e+06u
M1012 a_1162_100# a_828_74# a_1026_100# VNB nlowvt w=420000u l=150000u
+  ad=1.995e+11p pd=1.79e+06u as=2.226e+11p ps=1.9e+06u
M1013 a_241_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1014 VPWR a_1814_48# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR SCE a_36_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1016 Q a_1814_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Q a_1814_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_1814_48# a_1766_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1019 Q a_1814_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1766_74# a_630_74# a_1587_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=4e+11p ps=2.59e+06u
M1021 a_828_74# a_630_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1022 a_223_74# a_36_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1023 a_301_74# D a_223_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_1814_48# Q VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_828_74# a_630_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1026 a_301_74# D a_241_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1026_100# a_630_74# a_301_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1814_48# a_1587_74# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_415_464# a_36_74# a_301_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VGND a_1587_74# a_1814_48# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1031 VGND a_1814_48# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1587_74# a_828_74# a_1257_74# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=2.365e+11p ps=1.96e+06u
M1033 a_1587_74# a_630_74# a_1257_74# VPB pshort w=840000u l=180000u
+  ad=2.709e+11p pd=2.4e+06u as=7.308e+11p ps=3.42e+06u
M1034 VGND a_1257_74# a_1162_100# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1257_74# a_1026_100# VGND VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND SCE a_36_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1037 a_1257_74# a_1026_100# VPWR VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1767_476# a_828_74# a_1587_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* File: sky130_fd_sc_ms__sedfxbp_1.spice
* Created: Wed Sep  2 12:32:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sedfxbp_1.pex.spice"
.subckt sky130_fd_sc_ms__sedfxbp_1  VNB VPB D DE SCD SCE CLK VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCE	SCE
* SCD	SCD
* DE	DE
* D	D
* VPB	VPB
* VNB	VNB
MM1021 A_157_90# N_D_M1021_g N_A_27_90#_M1021_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.21 PD=0.66 PS=1.84 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_DE_M1022_g A_157_90# VNB NLOWVT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.8 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_DE_M1019_g N_A_161_394#_M1019_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1017 A_533_113# N_A_161_394#_M1017_g N_VGND_M1019_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_A_27_90#_M1006_d N_A_575_305#_M1006_g A_533_113# VNB NLOWVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75001.1 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1033 N_A_697_113#_M1033_d N_A_667_87#_M1033_g N_A_27_90#_M1006_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.1491 AS=0.0588 PD=1.55 PS=0.7 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1042 N_VGND_M1042_d N_SCE_M1042_g N_A_667_87#_M1042_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0756 AS=0.1197 PD=0.78 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1028 A_1075_125# N_SCD_M1028_g N_VGND_M1042_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0756 PD=0.66 PS=0.78 NRD=18.564 NRS=2.856 M=1 R=2.8 SA=75000.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1018 N_A_697_113#_M1018_d N_SCE_M1018_g A_1075_125# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 N_A_1351_74#_M1023_d N_CLK_M1023_g N_VGND_M1023_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1011 N_A_1549_74#_M1011_d N_A_1351_74#_M1011_g N_VGND_M1011_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.2109 PD=2.05 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_A_1747_118#_M1001_d N_A_1351_74#_M1001_g N_A_697_113#_M1001_s VNB
+ NLOWVT L=0.15 W=0.42 AD=0.1239 AS=0.1197 PD=1.01 PS=1.41 NRD=79.992 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1002 A_1895_118# N_A_1549_74#_M1002_g N_A_1747_118#_M1001_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.08085 AS=0.1239 PD=0.805 PS=1.01 NRD=39.276 NRS=8.568 M=1 R=2.8
+ SA=75000.9 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1027 N_VGND_M1027_d N_A_1972_92#_M1027_g A_1895_118# VNB NLOWVT L=0.15 W=0.42
+ AD=0.163364 AS=0.08085 PD=1.03811 PS=0.805 NRD=34.284 NRS=39.276 M=1 R=2.8
+ SA=75001.5 SB=75001 A=0.063 P=1.14 MULT=1
MM1040 N_A_1972_92#_M1040_d N_A_1747_118#_M1040_g N_VGND_M1027_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.192 AS=0.248936 PD=1.88 PS=1.58189 NRD=2.808 NRS=51.552 M=1
+ R=4.26667 SA=75001.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1024 A_2391_74# N_A_1972_92#_M1024_g N_VGND_M1024_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1824 PD=0.85 PS=1.85 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.8 A=0.096 P=1.58 MULT=1
MM1025 N_A_2463_74#_M1025_d N_A_1549_74#_M1025_g A_2391_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.129147 AS=0.0672 PD=1.20755 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667
+ SA=75000.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1036 A_2565_74# N_A_1351_74#_M1036_g N_A_2463_74#_M1025_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0847528 PD=0.66 PS=0.792453 NRD=18.564 NRS=23.568 M=1
+ R=2.8 SA=75001.1 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1037 N_VGND_M1037_d N_A_575_305#_M1037_g A_2565_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.165742 AS=0.0504 PD=1.19264 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.5
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1031 N_A_575_305#_M1031_d N_A_2463_74#_M1031_g N_VGND_M1037_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.252558 PD=1.85 PS=1.81736 NRD=0 NRS=13.116 M=1
+ R=4.26667 SA=75001.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1041 N_VGND_M1041_d N_A_2463_74#_M1041_g N_Q_M1041_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1961 AS=0.2109 PD=1.27 PS=2.05 NRD=40.536 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.9 A=0.111 P=1.78 MULT=1
MM1004 N_Q_N_M1004_d N_A_575_305#_M1004_g N_VGND_M1041_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1961 PD=2.05 PS=1.27 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1012 A_119_464# N_D_M1012_g N_A_27_90#_M1012_s VPB PSHORT L=0.18 W=0.64
+ AD=0.0672 AS=0.1792 PD=0.85 PS=1.84 NRD=15.3857 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1029 N_VPWR_M1029_d N_A_161_394#_M1029_g A_119_464# VPB PSHORT L=0.18 W=0.64
+ AD=0.1792 AS=0.0672 PD=1.84 PS=0.85 NRD=0 NRS=15.3857 M=1 R=3.55556 SA=90000.6
+ SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1005 N_VPWR_M1005_d N_DE_M1005_g N_A_161_394#_M1005_s VPB PSHORT L=0.18 W=0.64
+ AD=0.16 AS=0.1792 PD=1.14 PS=1.84 NRD=69.2455 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90001.7 A=0.1152 P=1.64 MULT=1
MM1026 A_559_464# N_DE_M1026_g N_VPWR_M1005_d VPB PSHORT L=0.18 W=0.64 AD=0.0768
+ AS=0.16 PD=0.88 PS=1.14 NRD=19.9955 NRS=0 M=1 R=3.55556 SA=90000.9 SB=90001.1
+ A=0.1152 P=1.64 MULT=1
MM1030 N_A_27_90#_M1030_d N_A_575_305#_M1030_g A_559_464# VPB PSHORT L=0.18
+ W=0.64 AD=0.0864 AS=0.0768 PD=0.91 PS=0.88 NRD=0 NRS=19.9955 M=1 R=3.55556
+ SA=90001.3 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1039 N_A_697_113#_M1039_d N_SCE_M1039_g N_A_27_90#_M1030_d VPB PSHORT L=0.18
+ W=0.64 AD=0.1792 AS=0.0864 PD=1.84 PS=0.91 NRD=0 NRS=0 M=1 R=3.55556
+ SA=90001.7 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1038 N_VPWR_M1038_d N_SCE_M1038_g N_A_667_87#_M1038_s VPB PSHORT L=0.18 W=0.64
+ AD=0.1392 AS=0.2208 PD=1.075 PS=1.97 NRD=49.2303 NRS=18.4589 M=1 R=3.55556
+ SA=90000.3 SB=90001.2 A=0.1152 P=1.64 MULT=1
MM1008 A_1071_462# N_SCD_M1008_g N_VPWR_M1038_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0672 AS=0.1392 PD=0.85 PS=1.075 NRD=15.3857 NRS=0 M=1 R=3.55556
+ SA=90000.9 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1032 N_A_697_113#_M1032_d N_A_667_87#_M1032_g A_1071_462# VPB PSHORT L=0.18
+ W=0.64 AD=0.1792 AS=0.0672 PD=1.84 PS=0.85 NRD=0 NRS=15.3857 M=1 R=3.55556
+ SA=90001.3 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1016 N_A_1351_74#_M1016_d N_CLK_M1016_g N_VPWR_M1016_s VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.3136 PD=2.8 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1000 N_A_1549_74#_M1000_d N_A_1351_74#_M1000_g N_VPWR_M1000_s VPB PSHORT
+ L=0.18 W=1.12 AD=0.3136 AS=0.3136 PD=2.8 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1010 N_A_1747_118#_M1010_d N_A_1549_74#_M1010_g N_A_697_113#_M1010_s VPB
+ PSHORT L=0.18 W=0.42 AD=0.0672 AS=0.1239 PD=0.74 PS=1.43 NRD=21.0987
+ NRS=2.3443 M=1 R=2.33333 SA=90000.2 SB=90001.5 A=0.0756 P=1.2 MULT=1
MM1009 A_1934_508# N_A_1351_74#_M1009_g N_A_1747_118#_M1010_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0525 AS=0.0672 PD=0.67 PS=0.74 NRD=32.8202 NRS=0 M=1 R=2.33333
+ SA=90000.7 SB=90001 A=0.0756 P=1.2 MULT=1
MM1013 N_VPWR_M1013_d N_A_1972_92#_M1013_g A_1934_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.0936833 AS=0.0525 PD=0.89 PS=0.67 NRD=2.3443 NRS=32.8202 M=1 R=2.33333
+ SA=90001.1 SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1035 N_A_1972_92#_M1035_d N_A_1747_118#_M1035_g N_VPWR_M1013_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.2352 AS=0.187367 PD=2.24 PS=1.78 NRD=0 NRS=19.9167 M=1
+ R=4.66667 SA=90000.7 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1043 A_2348_392# N_A_1972_92#_M1043_g N_VPWR_M1043_s VPB PSHORT L=0.18 W=1
+ AD=0.3975 AS=0.3882 PD=1.795 PS=2.89 NRD=67.4528 NRS=16.7253 M=1 R=5.55556
+ SA=90000.3 SB=90001.9 A=0.18 P=2.36 MULT=1
MM1034 N_A_2463_74#_M1034_d N_A_1351_74#_M1034_g A_2348_392# VPB PSHORT L=0.18
+ W=1 AD=0.219366 AS=0.3975 PD=1.90845 PS=1.795 NRD=0 NRS=67.4528 M=1 R=5.55556
+ SA=90001.2 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1007 A_2650_508# N_A_1549_74#_M1007_g N_A_2463_74#_M1034_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0921338 PD=0.66 PS=0.801549 NRD=30.4759 NRS=37.5088 M=1
+ R=2.33333 SA=90001.8 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1020 N_VPWR_M1020_d N_A_575_305#_M1020_g A_2650_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.108727 AS=0.0504 PD=0.90507 PS=0.66 NRD=58.6272 NRS=30.4759 M=1 R=2.33333
+ SA=90002.2 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1003 N_A_575_305#_M1003_d N_A_2463_74#_M1003_g N_VPWR_M1020_d VPB PSHORT
+ L=0.18 W=1 AD=0.28 AS=0.258873 PD=2.56 PS=2.15493 NRD=0 NRS=24.6053 M=1
+ R=5.55556 SA=90001.3 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1015 N_VPWR_M1015_d N_A_2463_74#_M1015_g N_Q_M1015_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.3136 PD=1.44 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1014 N_Q_N_M1014_d N_A_575_305#_M1014_g N_VPWR_M1015_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.1792 PD=2.8 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90000.7 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX44_noxref VNB VPB NWDIODE A=31.062 P=37.12
c_175 VNB 0 1.45871e-19 $X=0 $Y=0
c_333 VPB 0 1.97671e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__sedfxbp_1.pxi.spice"
*
.ends
*
*

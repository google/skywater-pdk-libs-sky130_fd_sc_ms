# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__sdfxbp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_ms__sdfxbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.44000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.470000 1.655000 1.800000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.590000 1.800000 10.950000 1.970000 ;
        RECT 10.590000 1.970000 10.840000 2.980000 ;
        RECT 10.620000 0.350000 10.950000 1.130000 ;
        RECT 10.780000 1.130000 10.950000 1.800000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.520700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.550000 0.900000 13.315000 1.150000 ;
        RECT 12.555000 1.820000 13.315000 2.150000 ;
        RECT 12.555000 2.150000 12.835000 2.980000 ;
        RECT 13.075000 1.150000 13.315000 1.820000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.405000 1.775000 2.755000 2.150000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.900000 2.075000 1.230000 ;
        RECT 1.565000 0.810000 2.075000 0.900000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.312600 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.265000 1.350000 3.685000 1.780000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 13.440000 0.085000 ;
        RECT  0.660000  0.085000  0.990000 0.730000 ;
        RECT  2.695000  0.085000  2.945000 1.130000 ;
        RECT  3.685000  0.085000  4.015000 0.840000 ;
        RECT  6.340000  0.085000  6.670000 0.600000 ;
        RECT  8.680000  0.085000  9.390000 0.715000 ;
        RECT 10.120000  0.085000 10.450000 1.130000 ;
        RECT 11.130000  0.085000 11.380000 1.130000 ;
        RECT 12.120000  0.085000 12.450000 0.730000 ;
        RECT 12.120000  0.730000 12.380000 1.150000 ;
        RECT 12.995000  0.085000 13.325000 0.730000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 13.440000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 13.440000 3.415000 ;
        RECT  0.725000 2.310000  1.055000 3.245000 ;
        RECT  2.670000 2.710000  3.090000 3.245000 ;
        RECT  4.075000 2.710000  4.405000 3.245000 ;
        RECT  6.575000 2.955000  6.905000 3.245000 ;
        RECT  8.860000 2.650000  9.430000 3.245000 ;
        RECT 10.140000 1.820000 10.390000 3.245000 ;
        RECT 11.040000 2.140000 11.370000 3.245000 ;
        RECT 11.120000 1.820000 11.370000 2.140000 ;
        RECT 12.105000 1.820000 12.355000 3.245000 ;
        RECT 13.005000 2.320000 13.335000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 13.440000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.085000 0.350000  0.490000 0.730000 ;
      RECT  0.085000 0.730000  0.255000 1.470000 ;
      RECT  0.085000 1.470000  0.915000 1.800000 ;
      RECT  0.085000 1.800000  0.520000 2.925000 ;
      RECT  0.745000 1.800000  0.915000 1.970000 ;
      RECT  0.745000 1.970000  2.195000 2.140000 ;
      RECT  1.480000 0.390000  2.415000 0.640000 ;
      RECT  1.650000 2.310000  1.980000 2.370000 ;
      RECT  1.650000 2.370000  4.745000 2.495000 ;
      RECT  1.650000 2.495000  5.335000 2.540000 ;
      RECT  1.650000 2.540000  1.980000 2.925000 ;
      RECT  1.865000 1.725000  2.195000 1.970000 ;
      RECT  2.245000 0.640000  2.415000 1.350000 ;
      RECT  2.245000 1.350000  3.095000 1.520000 ;
      RECT  2.925000 1.520000  3.095000 2.370000 ;
      RECT  3.125000 0.350000  3.455000 1.010000 ;
      RECT  3.125000 1.010000  4.025000 1.180000 ;
      RECT  3.295000 1.950000  4.095000 2.200000 ;
      RECT  3.855000 1.180000  4.025000 1.350000 ;
      RECT  3.855000 1.350000  4.095000 1.950000 ;
      RECT  4.195000 0.255000  6.080000 0.425000 ;
      RECT  4.195000 0.425000  4.445000 1.130000 ;
      RECT  4.265000 1.480000  4.900000 1.650000 ;
      RECT  4.265000 1.650000  4.435000 2.370000 ;
      RECT  4.575000 2.540000  5.335000 2.665000 ;
      RECT  4.605000 1.820000  4.855000 2.005000 ;
      RECT  4.605000 2.005000  5.335000 2.200000 ;
      RECT  4.650000 0.595000  4.900000 1.480000 ;
      RECT  5.005000 2.200000  5.335000 2.325000 ;
      RECT  5.070000 0.425000  5.240000 2.005000 ;
      RECT  5.085000 2.665000  5.335000 2.935000 ;
      RECT  5.410000 0.595000  5.740000 0.875000 ;
      RECT  5.410000 0.875000  5.580000 1.575000 ;
      RECT  5.410000 1.575000  7.010000 1.745000 ;
      RECT  5.505000 1.745000  5.675000 2.475000 ;
      RECT  5.505000 2.475000  5.865000 2.935000 ;
      RECT  5.750000 1.045000  6.080000 1.375000 ;
      RECT  5.845000 1.915000  6.205000 2.245000 ;
      RECT  5.910000 0.425000  6.080000 0.770000 ;
      RECT  5.910000 0.770000  7.010000 0.940000 ;
      RECT  5.910000 0.940000  6.080000 1.045000 ;
      RECT  6.035000 2.245000  6.205000 2.615000 ;
      RECT  6.035000 2.615000  7.735000 2.785000 ;
      RECT  6.250000 1.110000  7.350000 1.405000 ;
      RECT  6.730000 1.745000  7.010000 1.945000 ;
      RECT  6.840000 0.255000  7.690000 0.425000 ;
      RECT  6.840000 0.425000  7.010000 0.770000 ;
      RECT  7.110000 2.115000  7.395000 2.445000 ;
      RECT  7.180000 0.595000  7.350000 1.110000 ;
      RECT  7.180000 1.405000  7.350000 2.115000 ;
      RECT  7.520000 0.425000  7.690000 1.030000 ;
      RECT  7.520000 1.030000  7.780000 1.225000 ;
      RECT  7.520000 1.225000  8.680000 1.395000 ;
      RECT  7.565000 1.600000  7.895000 1.930000 ;
      RECT  7.565000 1.930000  7.735000 2.615000 ;
      RECT  7.860000 0.350000  8.190000 0.810000 ;
      RECT  7.905000 2.100000  8.235000 2.980000 ;
      RECT  8.020000 0.810000  8.190000 0.885000 ;
      RECT  8.020000 0.885000  9.020000 1.055000 ;
      RECT  8.065000 1.720000  9.020000 1.890000 ;
      RECT  8.065000 1.890000  8.235000 2.100000 ;
      RECT  8.350000 1.395000  8.680000 1.550000 ;
      RECT  8.710000 2.060000  9.950000 2.380000 ;
      RECT  8.850000 1.055000  9.610000 1.225000 ;
      RECT  8.850000 1.225000  9.020000 1.720000 ;
      RECT  9.280000 1.225000  9.610000 1.550000 ;
      RECT  9.560000 0.350000  9.950000 0.885000 ;
      RECT  9.600000 1.940000  9.950000 2.060000 ;
      RECT  9.600000 2.380000  9.950000 2.980000 ;
      RECT  9.780000 0.885000  9.950000 1.300000 ;
      RECT  9.780000 1.300000 10.610000 1.630000 ;
      RECT  9.780000 1.630000  9.950000 1.940000 ;
      RECT 11.580000 0.560000 11.940000 1.320000 ;
      RECT 11.580000 1.320000 12.735000 1.650000 ;
      RECT 11.580000 1.650000 11.910000 2.860000 ;
  END
END sky130_fd_sc_ms__sdfxbp_2

* File: sky130_fd_sc_ms__sdfstp_2.pex.spice
* Created: Fri Aug 28 18:13:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SDFSTP_2%SCE 2 5 9 11 13 17 24 25 27 28 32 36
r78 36 38 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.635
+ $X2=0.61 $Y2=1.47
r79 32 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.64
+ $Y=1.635 $X2=0.64 $Y2=1.635
r80 28 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.96 $Y=1.415
+ $X2=1.96 $Y2=1.25
r81 27 30 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=1.92 $Y=1.415 $X2=1.92
+ $Y2=1.495
r82 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.96
+ $Y=1.415 $X2=1.96 $Y2=1.415
r83 25 32 9.23067 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.805 $Y=1.495
+ $X2=0.72 $Y2=1.58
r84 24 30 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.795 $Y=1.495
+ $X2=1.92 $Y2=1.495
r85 24 25 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=1.795 $Y=1.495
+ $X2=0.805 $Y2=1.495
r86 17 40 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.94 $Y=0.58
+ $X2=1.94 $Y2=1.25
r87 11 13 194.355 $w=1.8e-07 $l=5e-07 $layer=POLY_cond $X=0.955 $Y=2.14
+ $X2=0.955 $Y2=2.64
r88 9 38 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=0.495 $Y=0.58
+ $X2=0.495 $Y2=1.47
r89 3 5 194.355 $w=1.8e-07 $l=5e-07 $layer=POLY_cond $X=0.505 $Y=2.14 $X2=0.505
+ $Y2=2.64
r90 2 11 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=0.61 $Y=2.065
+ $X2=0.955 $Y2=2.065
r91 2 3 53.8404 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=0.61 $Y=2.065
+ $X2=0.505 $Y2=2.065
r92 1 36 4.27811 $w=3.9e-07 $l=3e-08 $layer=POLY_cond $X=0.61 $Y=1.665 $X2=0.61
+ $Y2=1.635
r93 1 2 46.3462 $w=3.9e-07 $l=3.25e-07 $layer=POLY_cond $X=0.61 $Y=1.665
+ $X2=0.61 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_2%A_27_74# 1 2 9 12 16 19 22 26 27 31 32 34
+ 36 38
c79 27 0 1.86174e-19 $X=1.06 $Y=1.065
c80 22 0 1.61244e-19 $X=1.795 $Y=2.405
r81 32 42 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.96 $Y=1.995
+ $X2=1.96 $Y2=2.16
r82 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.96
+ $Y=1.995 $X2=1.96 $Y2=1.995
r83 29 31 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=1.92 $Y=2.32
+ $X2=1.92 $Y2=1.995
r84 27 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=1.065
+ $X2=1.06 $Y2=0.9
r85 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.06
+ $Y=1.065 $X2=1.06 $Y2=1.065
r86 24 34 0.364692 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=1.065
+ $X2=0.28 $Y2=1.065
r87 24 26 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=0.445 $Y=1.065
+ $X2=1.06 $Y2=1.065
r88 23 36 2.11342 $w=1.7e-07 $l=1.27475e-07 $layer=LI1_cond $X=0.365 $Y=2.405
+ $X2=0.24 $Y2=2.4
r89 22 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.795 $Y=2.405
+ $X2=1.92 $Y2=2.32
r90 22 23 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=1.795 $Y=2.405
+ $X2=0.365 $Y2=2.405
r91 19 36 4.3182 $w=2.1e-07 $l=1.08167e-07 $layer=LI1_cond $X=0.2 $Y=2.31
+ $X2=0.24 $Y2=2.4
r92 18 34 6.46576 $w=2.5e-07 $l=2.0106e-07 $layer=LI1_cond $X=0.2 $Y=1.23
+ $X2=0.28 $Y2=1.065
r93 18 19 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=0.2 $Y=1.23 $X2=0.2
+ $Y2=2.31
r94 14 34 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=0.9 $X2=0.28
+ $Y2=1.065
r95 14 16 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.28 $Y=0.9 $X2=0.28
+ $Y2=0.58
r96 12 42 186.581 $w=1.8e-07 $l=4.8e-07 $layer=POLY_cond $X=2.005 $Y=2.64
+ $X2=2.005 $Y2=2.16
r97 9 38 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.12 $Y=0.58 $X2=1.12
+ $Y2=0.9
r98 2 36 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.475
r99 1 16 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_2%D 3 7 9 12 13
c44 12 0 4.46515e-20 $X=1.42 $Y=1.985
r45 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=1.985
+ $X2=1.42 $Y2=2.15
r46 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=1.985
+ $X2=1.42 $Y2=1.82
r47 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.42
+ $Y=1.985 $X2=1.42 $Y2=1.985
r48 9 13 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.2 $Y=1.985 $X2=1.42
+ $Y2=1.985
r49 7 14 635.83 $w=1.5e-07 $l=1.24e-06 $layer=POLY_cond $X=1.51 $Y=0.58 $X2=1.51
+ $Y2=1.82
r50 3 15 190.468 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=1.375 $Y=2.64
+ $X2=1.375 $Y2=2.15
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_2%SCD 3 6 9 11 12 13 18 22
c44 11 0 1.0588e-19 $X=2.64 $Y=1.295
c45 9 0 1.61244e-19 $X=2.425 $Y=2.64
r46 22 24 40.6549 $w=4.95e-07 $l=1.65e-07 $layer=POLY_cond $X=2.582 $Y=1.985
+ $X2=2.582 $Y2=2.15
r47 18 20 46.3954 $w=4.95e-07 $l=1.65e-07 $layer=POLY_cond $X=2.582 $Y=1.305
+ $X2=2.582 $Y2=1.14
r48 13 22 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.665
+ $Y=1.985 $X2=2.665 $Y2=1.985
r49 12 13 16.3903 $w=2.23e-07 $l=3.2e-07 $layer=LI1_cond $X=2.667 $Y=1.665
+ $X2=2.667 $Y2=1.985
r50 11 12 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=2.667 $Y=1.295
+ $X2=2.667 $Y2=1.665
r51 11 18 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.665
+ $Y=1.305 $X2=2.665 $Y2=1.305
r52 9 24 190.468 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=2.425 $Y=2.64
+ $X2=2.425 $Y2=2.15
r53 6 22 8.86311 $w=4.95e-07 $l=8.2e-08 $layer=POLY_cond $X=2.582 $Y=1.903
+ $X2=2.582 $Y2=1.985
r54 5 18 8.86311 $w=4.95e-07 $l=8.2e-08 $layer=POLY_cond $X=2.582 $Y=1.387
+ $X2=2.582 $Y2=1.305
r55 5 6 55.7728 $w=4.95e-07 $l=5.16e-07 $layer=POLY_cond $X=2.582 $Y=1.387
+ $X2=2.582 $Y2=1.903
r56 3 20 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.41 $Y=0.58 $X2=2.41
+ $Y2=1.14
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_2%CLK 3 6 8 11 13
c38 11 0 1.80078e-19 $X=3.42 $Y=1.385
c39 6 0 1.0588e-19 $X=3.485 $Y=2.4
r40 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.42 $Y=1.385
+ $X2=3.42 $Y2=1.55
r41 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.42 $Y=1.385
+ $X2=3.42 $Y2=1.22
r42 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.42
+ $Y=1.385 $X2=3.42 $Y2=1.385
r43 8 12 5.60648 $w=3.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.6 $Y=1.365 $X2=3.42
+ $Y2=1.365
r44 6 14 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.485 $Y=2.4
+ $X2=3.485 $Y2=1.55
r45 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.4 $Y=0.74 $X2=3.4
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_2%A_795_74# 1 2 9 11 13 17 21 22 23 25 26 28
+ 30 33 36 39 43 45 46 47 48 51 55 56 57 58 61 62 63 65 67 68 72 75 76 80 86 87
+ 95 96 97 101
c278 75 0 3.7885e-19 $X=10.555 $Y=1.97
c279 68 0 3.47781e-20 $X=10 $Y=1.64
c280 28 0 3.01101e-20 $X=10.13 $Y=1.085
c281 11 0 1.3233e-19 $X=5.4 $Y=1.655
c282 9 0 4.72054e-20 $X=4.975 $Y=2.495
r283 96 97 24.9528 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.565 $Y=1.655
+ $X2=5.565 $Y2=1.58
r284 94 95 33.0969 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.975 $Y=1.565
+ $X2=5.065 $Y2=1.565
r285 86 87 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=8.255 $Y=1.685
+ $X2=8.425 $Y2=1.685
r286 84 96 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=5.565 $Y=1.88
+ $X2=5.565 $Y2=1.655
r287 83 85 16.0091 $w=2.21e-07 $l=2.9e-07 $layer=LI1_cond $X=5.602 $Y=1.88
+ $X2=5.602 $Y2=2.17
r288 83 84 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.565
+ $Y=1.88 $X2=5.565 $Y2=1.88
r289 76 105 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.555 $Y=1.97
+ $X2=10.555 $Y2=2.135
r290 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.555
+ $Y=1.97 $X2=10.555 $Y2=1.97
r291 73 75 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=10.17 $Y=1.97
+ $X2=10.555 $Y2=1.97
r292 72 101 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.975 $Y=1.64
+ $X2=8.975 $Y2=1.475
r293 71 87 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=8.975 $Y=1.64
+ $X2=8.425 $Y2=1.64
r294 71 72 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.975
+ $Y=1.64 $X2=8.975 $Y2=1.64
r295 68 73 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=10.085 $Y=1.64
+ $X2=10.085 $Y2=1.97
r296 68 71 35.7956 $w=3.28e-07 $l=1.025e-06 $layer=LI1_cond $X=10 $Y=1.64
+ $X2=8.975 $Y2=1.64
r297 67 86 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=7.365 $Y=1.81
+ $X2=8.255 $Y2=1.81
r298 64 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.28 $Y=1.895
+ $X2=7.365 $Y2=1.81
r299 64 65 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=7.28 $Y=1.895
+ $X2=7.28 $Y2=2.905
r300 62 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.195 $Y=2.99
+ $X2=7.28 $Y2=2.905
r301 62 63 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.195 $Y=2.99
+ $X2=6.685 $Y2=2.99
r302 61 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.6 $Y=2.905
+ $X2=6.685 $Y2=2.99
r303 60 61 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.6 $Y=2.255
+ $X2=6.6 $Y2=2.905
r304 59 85 2.27611 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=5.73 $Y=2.17
+ $X2=5.602 $Y2=2.17
r305 58 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.515 $Y=2.17
+ $X2=6.6 $Y2=2.255
r306 58 59 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=6.515 $Y=2.17
+ $X2=5.73 $Y2=2.17
r307 56 85 5.3732 $w=2.21e-07 $l=1.04307e-07 $layer=LI1_cond $X=5.645 $Y=2.255
+ $X2=5.602 $Y2=2.17
r308 56 57 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.645 $Y=2.255
+ $X2=5.645 $Y2=2.895
r309 55 80 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.085 $Y=1.015
+ $X2=5.085 $Y2=1.1
r310 54 55 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.085 $Y=0.425
+ $X2=5.085 $Y2=1.015
r311 52 94 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=4.875 $Y=1.565
+ $X2=4.975 $Y2=1.565
r312 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.875
+ $Y=1.565 $X2=4.875 $Y2=1.565
r313 49 80 14.5487 $w=1.68e-07 $l=2.23e-07 $layer=LI1_cond $X=4.862 $Y=1.1
+ $X2=5.085 $Y2=1.1
r314 49 51 20.5588 $w=2.03e-07 $l=3.8e-07 $layer=LI1_cond $X=4.862 $Y=1.185
+ $X2=4.862 $Y2=1.565
r315 47 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.56 $Y=2.98
+ $X2=5.645 $Y2=2.895
r316 47 48 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=5.56 $Y=2.98
+ $X2=4.325 $Y2=2.98
r317 45 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5 $Y=0.34
+ $X2=5.085 $Y2=0.425
r318 45 46 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=5 $Y=0.34 $X2=4.2
+ $Y2=0.34
r319 41 48 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.2 $Y=2.895
+ $X2=4.325 $Y2=2.98
r320 41 43 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=4.2 $Y=2.895
+ $X2=4.2 $Y2=2.78
r321 37 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.115 $Y=0.425
+ $X2=4.2 $Y2=0.34
r322 37 39 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.115 $Y=0.425
+ $X2=4.115 $Y2=0.515
r323 33 105 239.056 $w=1.8e-07 $l=6.15e-07 $layer=POLY_cond $X=10.63 $Y=2.75
+ $X2=10.63 $Y2=2.135
r324 28 30 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=10.13 $Y=1.085
+ $X2=10.13 $Y2=0.69
r325 27 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.775 $Y=1.16
+ $X2=9.7 $Y2=1.16
r326 26 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.055 $Y=1.16
+ $X2=10.13 $Y2=1.085
r327 26 27 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=10.055 $Y=1.16
+ $X2=9.775 $Y2=1.16
r328 23 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.7 $Y=1.085
+ $X2=9.7 $Y2=1.16
r329 23 25 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=9.7 $Y=1.085
+ $X2=9.7 $Y2=0.69
r330 21 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.625 $Y=1.16
+ $X2=9.7 $Y2=1.16
r331 21 22 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=9.625 $Y=1.16
+ $X2=9.14 $Y2=1.16
r332 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.065 $Y=1.235
+ $X2=9.14 $Y2=1.16
r333 19 101 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=9.065 $Y=1.235
+ $X2=9.065 $Y2=1.475
r334 17 35 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=5.64 $Y=0.615
+ $X2=5.64 $Y2=1.26
r335 13 35 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.625 $Y=1.35
+ $X2=5.625 $Y2=1.26
r336 13 97 89.4032 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=5.625 $Y=1.35
+ $X2=5.625 $Y2=1.58
r337 11 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.4 $Y=1.655
+ $X2=5.565 $Y2=1.655
r338 11 95 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.4 $Y=1.655
+ $X2=5.065 $Y2=1.655
r339 7 94 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.975 $Y=1.73
+ $X2=4.975 $Y2=1.565
r340 7 9 297.363 $w=1.8e-07 $l=7.65e-07 $layer=POLY_cond $X=4.975 $Y=1.73
+ $X2=4.975 $Y2=2.495
r341 2 43 600 $w=1.7e-07 $l=1.00524e-06 $layer=licon1_PDIFF $count=1 $X=4.025
+ $Y=1.84 $X2=4.16 $Y2=2.78
r342 1 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.975
+ $Y=0.37 $X2=4.115 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_2%A_1185_55# 1 2 7 9 12 14 18 21 23 24 27 31
+ 33 35 40
c96 33 0 1.75838e-19 $X=6.27 $Y=1.815
c97 7 0 5.96633e-20 $X=6 $Y=0.935
r98 35 37 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=6.855 $Y=0.525
+ $X2=6.855 $Y2=0.615
r99 31 41 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.105 $Y=1.815
+ $X2=6.105 $Y2=1.98
r100 31 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.105 $Y=1.815
+ $X2=6.105 $Y2=1.65
r101 30 33 9.43135 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=6.105 $Y=1.815
+ $X2=6.27 $Y2=1.815
r102 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.105
+ $Y=1.815 $X2=6.105 $Y2=1.815
r103 25 27 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=6.94 $Y=1.915
+ $X2=6.94 $Y2=2.515
r104 23 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.69 $Y=0.615
+ $X2=6.855 $Y2=0.615
r105 23 24 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.69 $Y=0.615
+ $X2=6.31 $Y2=0.615
r106 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.855 $Y=1.83
+ $X2=6.94 $Y2=1.915
r107 21 33 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=6.855 $Y=1.83
+ $X2=6.27 $Y2=1.83
r108 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.145
+ $Y=1.1 $X2=6.145 $Y2=1.1
r109 16 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.145 $Y=0.7
+ $X2=6.31 $Y2=0.615
r110 16 18 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=6.145 $Y=0.7 $X2=6.145
+ $Y2=1.1
r111 14 19 38.8445 $w=3.55e-07 $l=1.93533e-07 $layer=POLY_cond $X=6.055 $Y=1.265
+ $X2=6.117 $Y2=1.1
r112 14 40 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=6.055 $Y=1.265
+ $X2=6.055 $Y2=1.65
r113 12 41 211.847 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=6.03 $Y=2.525
+ $X2=6.03 $Y2=1.98
r114 7 19 38.8445 $w=3.55e-07 $l=2.15708e-07 $layer=POLY_cond $X=6 $Y=0.935
+ $X2=6.117 $Y2=1.1
r115 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6 $Y=0.935 $X2=6
+ $Y2=0.615
r116 2 27 600 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_PDIFF $count=1 $X=6.805
+ $Y=2.315 $X2=6.94 $Y2=2.515
r117 1 35 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=6.71
+ $Y=0.37 $X2=6.855 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_2%A_991_81# 1 2 7 9 11 13 16 18 20 23 25 27
+ 31 34 36 42 44 45 49 50 51 52 55 60 62 68
c182 52 0 5.96633e-20 $X=6.88 $Y=0.955
c183 42 0 2.09475e-20 $X=5.425 $Y=0.615
c184 34 0 1.3233e-19 $X=5.24 $Y=2.39
c185 31 0 2.52187e-20 $X=7.07 $Y=0.94
c186 9 0 1.75838e-19 $X=6.715 $Y=2.525
r187 67 68 24.0272 $w=3.31e-07 $l=1.65e-07 $layer=POLY_cond $X=8.13 $Y=1.32
+ $X2=8.295 $Y2=1.32
r188 61 67 30.5801 $w=3.31e-07 $l=2.1e-07 $layer=POLY_cond $X=7.92 $Y=1.32
+ $X2=8.13 $Y2=1.32
r189 61 65 10.9215 $w=3.31e-07 $l=7.5e-08 $layer=POLY_cond $X=7.92 $Y=1.32
+ $X2=7.845 $Y2=1.32
r190 60 62 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.92 $Y=1.39
+ $X2=7.92 $Y2=1.225
r191 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.92
+ $Y=1.39 $X2=7.92 $Y2=1.39
r192 53 62 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=7.84 $Y=1.04
+ $X2=7.84 $Y2=1.225
r193 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.755 $Y=0.955
+ $X2=7.84 $Y2=1.04
r194 51 52 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=7.755 $Y=0.955
+ $X2=6.88 $Y2=0.955
r195 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.715
+ $Y=1.065 $X2=6.715 $Y2=1.065
r196 47 49 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=6.715 $Y=1.375
+ $X2=6.715 $Y2=1.065
r197 46 52 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.715 $Y=1.04
+ $X2=6.88 $Y2=0.955
r198 46 49 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=6.715 $Y=1.04
+ $X2=6.715 $Y2=1.065
r199 44 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.55 $Y=1.46
+ $X2=6.715 $Y2=1.375
r200 44 45 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.55 $Y=1.46
+ $X2=5.59 $Y2=1.46
r201 40 45 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.465 $Y=1.46
+ $X2=5.59 $Y2=1.46
r202 40 56 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.465 $Y=1.46
+ $X2=5.22 $Y2=1.46
r203 40 42 35.0343 $w=2.48e-07 $l=7.6e-07 $layer=LI1_cond $X=5.465 $Y=1.375
+ $X2=5.465 $Y2=0.615
r204 38 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.22 $Y=1.545
+ $X2=5.22 $Y2=1.46
r205 38 55 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=5.22 $Y=1.545
+ $X2=5.22 $Y2=2.265
r206 34 55 6.55365 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=5.24 $Y=2.39
+ $X2=5.24 $Y2=2.265
r207 34 36 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=5.24 $Y=2.39
+ $X2=5.24 $Y2=2.495
r208 33 50 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.715 $Y=1.405
+ $X2=6.715 $Y2=1.065
r209 29 50 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=6.715 $Y=1.015
+ $X2=6.715 $Y2=1.065
r210 29 31 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=6.715 $Y=0.94
+ $X2=7.07 $Y2=0.94
r211 25 68 38.5891 $w=3.31e-07 $l=3.64005e-07 $layer=POLY_cond $X=8.56 $Y=1.085
+ $X2=8.295 $Y2=1.32
r212 25 27 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.56 $Y=1.085
+ $X2=8.56 $Y2=0.69
r213 21 68 17.0024 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=8.295 $Y=1.555
+ $X2=8.295 $Y2=1.32
r214 21 23 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=8.295 $Y=1.555
+ $X2=8.295 $Y2=2.315
r215 18 67 21.295 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=8.13 $Y=1.085
+ $X2=8.13 $Y2=1.32
r216 18 20 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.13 $Y=1.085
+ $X2=8.13 $Y2=0.69
r217 14 65 17.0024 $w=1.8e-07 $l=2.35e-07 $layer=POLY_cond $X=7.845 $Y=1.555
+ $X2=7.845 $Y2=1.32
r218 14 16 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=7.845 $Y=1.555
+ $X2=7.845 $Y2=2.315
r219 11 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.07 $Y=0.865
+ $X2=7.07 $Y2=0.94
r220 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.07 $Y=0.865
+ $X2=7.07 $Y2=0.58
r221 7 33 34.7712 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.715 $Y=1.57
+ $X2=6.715 $Y2=1.405
r222 7 9 371.218 $w=1.8e-07 $l=9.55e-07 $layer=POLY_cond $X=6.715 $Y=1.57
+ $X2=6.715 $Y2=2.525
r223 2 36 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=5.065
+ $Y=2.285 $X2=5.2 $Y2=2.495
r224 1 42 182 $w=1.7e-07 $l=5.65332e-07 $layer=licon1_NDIFF $count=1 $X=4.955
+ $Y=0.405 $X2=5.425 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_2%SET_B 3 7 11 15 17 18 21 23 30 33 41
c132 23 0 5.34496e-20 $X=11.76 $Y=1.295
c133 15 0 7.44554e-20 $X=11.59 $Y=0.58
c134 11 0 3.15842e-21 $X=11.47 $Y=2.75
c135 7 0 1.09822e-19 $X=7.46 $Y=0.58
r136 34 41 9.11234 $w=4.28e-07 $l=3.4e-07 $layer=LI1_cond $X=11.66 $Y=1.635
+ $X2=11.66 $Y2=1.295
r137 33 36 39.8861 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=11.577 $Y=1.635
+ $X2=11.577 $Y2=1.8
r138 33 35 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=11.577 $Y=1.635
+ $X2=11.577 $Y2=1.47
r139 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.61
+ $Y=1.635 $X2=11.61 $Y2=1.635
r140 28 30 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.37 $Y=1.39 $X2=7.46
+ $Y2=1.39
r141 25 28 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=7.21 $Y=1.39
+ $X2=7.37 $Y2=1.39
r142 23 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=1.295
+ $X2=11.76 $Y2=1.295
r143 21 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.37
+ $Y=1.39 $X2=7.37 $Y2=1.39
r144 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=1.295
+ $X2=7.44 $Y2=1.295
r145 18 20 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.585 $Y=1.295
+ $X2=7.44 $Y2=1.295
r146 17 23 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.615 $Y=1.295
+ $X2=11.76 $Y2=1.295
r147 17 18 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=11.615 $Y=1.295
+ $X2=7.585 $Y2=1.295
r148 15 35 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=11.59 $Y=0.58
+ $X2=11.59 $Y2=1.47
r149 11 36 369.274 $w=1.8e-07 $l=9.5e-07 $layer=POLY_cond $X=11.47 $Y=2.75
+ $X2=11.47 $Y2=1.8
r150 5 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.46 $Y=1.225
+ $X2=7.46 $Y2=1.39
r151 5 7 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=7.46 $Y=1.225
+ $X2=7.46 $Y2=0.58
r152 1 25 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.21 $Y=1.555
+ $X2=7.21 $Y2=1.39
r153 1 3 377.048 $w=1.8e-07 $l=9.7e-07 $layer=POLY_cond $X=7.21 $Y=1.555
+ $X2=7.21 $Y2=2.525
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_2%A_608_74# 1 2 9 13 16 20 21 22 23 24 27 31
+ 33 38 39 40 41 43 45 48 50 51 52 53 56 59 60 61 66 69 74
c198 66 0 1.80078e-19 $X=4.05 $Y=1.515
c199 21 0 2.09475e-20 $X=4.805 $Y=1.115
r200 70 72 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=3.9 $Y=1.515
+ $X2=3.935 $Y2=1.515
r201 67 74 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=4.05 $Y=1.515
+ $X2=4.425 $Y2=1.515
r202 67 72 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=4.05 $Y=1.515
+ $X2=3.935 $Y2=1.515
r203 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.05
+ $Y=1.515 $X2=4.05 $Y2=1.515
r204 64 66 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.05 $Y=1.82
+ $X2=4.05 $Y2=1.515
r205 61 63 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=3.13 $Y=1.945
+ $X2=3.26 $Y2=1.945
r206 60 64 6.98653 $w=2.5e-07 $l=2.18746e-07 $layer=LI1_cond $X=3.885 $Y=1.945
+ $X2=4.05 $Y2=1.82
r207 60 63 28.8111 $w=2.48e-07 $l=6.25e-07 $layer=LI1_cond $X=3.885 $Y=1.945
+ $X2=3.26 $Y2=1.945
r208 59 61 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.045 $Y=1.82
+ $X2=3.13 $Y2=1.945
r209 59 69 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=3.045 $Y=1.82
+ $X2=3.045 $Y2=1.01
r210 54 69 9.49412 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=3.155 $Y=0.815
+ $X2=3.155 $Y2=1.01
r211 54 56 8.86495 $w=3.88e-07 $l=3e-07 $layer=LI1_cond $X=3.155 $Y=0.815
+ $X2=3.155 $Y2=0.515
r212 50 51 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=4.44 $Y=1.97
+ $X2=4.44 $Y2=2.12
r213 46 48 443.543 $w=1.5e-07 $l=8.65e-07 $layer=POLY_cond $X=10.63 $Y=1.445
+ $X2=10.63 $Y2=0.58
r214 43 45 143.261 $w=1.8e-07 $l=5.35e-07 $layer=POLY_cond $X=9.89 $Y=3.075
+ $X2=9.89 $Y2=2.54
r215 42 53 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.53 $Y=3.15 $X2=9.44
+ $Y2=3.15
r216 41 43 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=9.8 $Y=3.15
+ $X2=9.89 $Y2=3.075
r217 41 42 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.8 $Y=3.15
+ $X2=9.53 $Y2=3.15
r218 39 46 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.555 $Y=1.52
+ $X2=10.63 $Y2=1.445
r219 39 40 525.585 $w=1.5e-07 $l=1.025e-06 $layer=POLY_cond $X=10.555 $Y=1.52
+ $X2=9.53 $Y2=1.52
r220 36 53 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.44 $Y=3.075
+ $X2=9.44 $Y2=3.15
r221 36 38 207.96 $w=1.8e-07 $l=5.35e-07 $layer=POLY_cond $X=9.44 $Y=3.075
+ $X2=9.44 $Y2=2.54
r222 35 40 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=9.44 $Y=1.595
+ $X2=9.53 $Y2=1.52
r223 35 38 367.331 $w=1.8e-07 $l=9.45e-07 $layer=POLY_cond $X=9.44 $Y=1.595
+ $X2=9.44 $Y2=2.54
r224 34 52 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.6 $Y=3.15 $X2=5.51
+ $Y2=3.15
r225 33 53 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.35 $Y=3.15 $X2=9.44
+ $Y2=3.15
r226 33 34 1922.87 $w=1.5e-07 $l=3.75e-06 $layer=POLY_cond $X=9.35 $Y=3.15
+ $X2=5.6 $Y2=3.15
r227 29 52 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=5.51 $Y=3.075
+ $X2=5.51 $Y2=3.15
r228 29 31 174.919 $w=1.8e-07 $l=4.5e-07 $layer=POLY_cond $X=5.51 $Y=3.075
+ $X2=5.51 $Y2=2.625
r229 25 27 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=4.88 $Y=1.04
+ $X2=4.88 $Y2=0.615
r230 23 52 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.42 $Y=3.15 $X2=5.51
+ $Y2=3.15
r231 23 24 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=5.42 $Y=3.15
+ $X2=4.53 $Y2=3.15
r232 21 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.805 $Y=1.115
+ $X2=4.88 $Y2=1.04
r233 21 22 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=4.805 $Y=1.115
+ $X2=4.5 $Y2=1.115
r234 20 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.455 $Y=3.075
+ $X2=4.53 $Y2=3.15
r235 20 51 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=4.455 $Y=3.075
+ $X2=4.455 $Y2=2.12
r236 17 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.425 $Y=1.68
+ $X2=4.425 $Y2=1.515
r237 17 50 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.425 $Y=1.68
+ $X2=4.425 $Y2=1.97
r238 16 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.425 $Y=1.35
+ $X2=4.425 $Y2=1.515
r239 15 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.425 $Y=1.19
+ $X2=4.5 $Y2=1.115
r240 15 16 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=4.425 $Y=1.19
+ $X2=4.425 $Y2=1.35
r241 11 72 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.935 $Y=1.68
+ $X2=3.935 $Y2=1.515
r242 11 13 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=3.935 $Y=1.68
+ $X2=3.935 $Y2=2.4
r243 7 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.9 $Y=1.35 $X2=3.9
+ $Y2=1.515
r244 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.9 $Y=1.35 $X2=3.9
+ $Y2=0.74
r245 2 63 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.125
+ $Y=1.84 $X2=3.26 $Y2=1.985
r246 1 56 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=3.04
+ $Y=0.37 $X2=3.185 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_2%A_2186_367# 1 2 7 9 13 16 17 21 23 24 27 30
+ 31 35 37 39
c104 35 0 6.56335e-20 $X=11.11 $Y=1.065
c105 16 0 3.1683e-20 $X=11.02 $Y=1.835
c106 9 0 1.88308e-19 $X=11.02 $Y=2.75
c107 7 0 1.557e-19 $X=11.02 $Y=1.925
r108 35 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.11 $Y=1.065
+ $X2=11.11 $Y2=1.23
r109 35 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.11 $Y=1.065
+ $X2=11.11 $Y2=0.9
r110 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.11
+ $Y=1.065 $X2=11.11 $Y2=1.065
r111 31 34 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=11.11 $Y=0.875
+ $X2=11.11 $Y2=1.065
r112 29 37 3.87901 $w=2.37e-07 $l=1.14039e-07 $layer=LI1_cond $X=12.72 $Y=0.96
+ $X2=12.652 $Y2=0.875
r113 29 30 88.0749 $w=1.68e-07 $l=1.35e-06 $layer=LI1_cond $X=12.72 $Y=0.96
+ $X2=12.72 $Y2=2.31
r114 25 37 3.87901 $w=2.37e-07 $l=8.5e-08 $layer=LI1_cond $X=12.652 $Y=0.79
+ $X2=12.652 $Y2=0.875
r115 25 27 7.93485 $w=3.03e-07 $l=2.1e-07 $layer=LI1_cond $X=12.652 $Y=0.79
+ $X2=12.652 $Y2=0.58
r116 23 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.635 $Y=2.395
+ $X2=12.72 $Y2=2.31
r117 23 24 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=12.635 $Y=2.395
+ $X2=12.31 $Y2=2.395
r118 19 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=12.185 $Y=2.48
+ $X2=12.31 $Y2=2.395
r119 19 21 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=12.185 $Y=2.48
+ $X2=12.185 $Y2=2.75
r120 18 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.275 $Y=0.875
+ $X2=11.11 $Y2=0.875
r121 17 37 2.57001 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=12.5 $Y=0.875
+ $X2=12.652 $Y2=0.875
r122 17 18 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=12.5 $Y=0.875
+ $X2=11.275 $Y2=0.875
r123 16 40 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=11.035 $Y=1.835
+ $X2=11.035 $Y2=1.23
r124 13 39 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.02 $Y=0.58
+ $X2=11.02 $Y2=0.9
r125 7 16 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=11.02 $Y=1.925
+ $X2=11.02 $Y2=1.835
r126 7 9 320.685 $w=1.8e-07 $l=8.25e-07 $layer=POLY_cond $X=11.02 $Y=1.925
+ $X2=11.02 $Y2=2.75
r127 2 21 600 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_PDIFF $count=1 $X=12.095
+ $Y=2.54 $X2=12.225 $Y2=2.75
r128 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.5
+ $Y=0.37 $X2=12.64 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_2%A_1804_424# 1 2 3 4 5 18 22 24 26 28 31 35
+ 36 39 41 42 43 48 52 54 56 57 58 60 63 65 67 69 70 72 77 79 81 84
c192 57 0 1.93538e-19 $X=10.89 $Y=1.485
c193 36 0 5.67555e-20 $X=13.43 $Y=1.365
r194 84 85 66.7385 $w=3.75e-07 $l=4.5e-07 $layer=POLY_cond $X=12.322 $Y=1.975
+ $X2=12.322 $Y2=1.525
r195 83 84 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=12.3
+ $Y=1.975 $X2=12.3 $Y2=1.975
r196 80 81 9.54788 $w=5.03e-07 $l=1.65e-07 $layer=LI1_cond $X=11.695 $Y=2.222
+ $X2=11.86 $Y2=2.222
r197 72 75 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=9.415 $Y=0.34
+ $X2=9.415 $Y2=0.53
r198 70 85 23.988 $w=2.62e-07 $l=1.98e-07 $layer=POLY_cond $X=12.322 $Y=1.327
+ $X2=12.322 $Y2=1.525
r199 69 70 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=12.3
+ $Y=1.295 $X2=12.3 $Y2=1.295
r200 67 83 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.3 $Y=1.97 $X2=12.3
+ $Y2=2.055
r201 67 69 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=12.3 $Y=1.97
+ $X2=12.3 $Y2=1.295
r202 65 83 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.135 $Y=2.055
+ $X2=12.3 $Y2=2.055
r203 65 81 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=12.135 $Y=2.055
+ $X2=11.86 $Y2=2.055
r204 61 80 3.22715 $w=3.3e-07 $l=2.53e-07 $layer=LI1_cond $X=11.695 $Y=2.475
+ $X2=11.695 $Y2=2.222
r205 61 63 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=11.695 $Y=2.475
+ $X2=11.695 $Y2=2.75
r206 60 80 17.053 $w=5.03e-07 $l=7.2e-07 $layer=LI1_cond $X=10.975 $Y=2.222
+ $X2=11.695 $Y2=2.222
r207 60 79 7.65311 $w=5.03e-07 $l=8.5e-08 $layer=LI1_cond $X=10.975 $Y=2.222
+ $X2=10.89 $Y2=2.222
r208 59 60 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=10.975 $Y=1.57
+ $X2=10.975 $Y2=1.97
r209 57 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.89 $Y=1.485
+ $X2=10.975 $Y2=1.57
r210 57 58 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.89 $Y=1.485
+ $X2=10.58 $Y2=1.485
r211 56 79 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=10.435 $Y=2.39
+ $X2=10.89 $Y2=2.39
r212 54 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.495 $Y=1.4
+ $X2=10.58 $Y2=1.485
r213 54 77 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=10.495 $Y=1.4
+ $X2=10.495 $Y2=0.81
r214 50 77 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=10.415 $Y=0.645
+ $X2=10.415 $Y2=0.81
r215 50 52 2.26996 $w=3.28e-07 $l=6.5e-08 $layer=LI1_cond $X=10.415 $Y=0.645
+ $X2=10.415 $Y2=0.58
r216 49 52 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=10.415 $Y=0.425
+ $X2=10.415 $Y2=0.58
r217 46 48 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=10.27 $Y=2.905
+ $X2=10.27 $Y2=2.745
r218 45 56 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.27 $Y=2.475
+ $X2=10.435 $Y2=2.39
r219 45 48 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=10.27 $Y=2.475
+ $X2=10.27 $Y2=2.745
r220 44 72 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.58 $Y=0.34
+ $X2=9.415 $Y2=0.34
r221 43 49 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.25 $Y=0.34
+ $X2=10.415 $Y2=0.425
r222 43 44 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.25 $Y=0.34
+ $X2=9.58 $Y2=0.34
r223 41 46 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.105 $Y=2.99
+ $X2=10.27 $Y2=2.905
r224 41 42 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=10.105 $Y=2.99
+ $X2=9.33 $Y2=2.99
r225 37 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.165 $Y=2.905
+ $X2=9.33 $Y2=2.99
r226 37 39 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=9.165 $Y=2.905
+ $X2=9.165 $Y2=2.4
r227 34 84 2.22462 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=12.322 $Y=1.99
+ $X2=12.322 $Y2=1.975
r228 34 35 37.3423 $w=3.75e-07 $l=1.5e-07 $layer=POLY_cond $X=12.337 $Y=1.99
+ $X2=12.337 $Y2=2.14
r229 29 36 33.9972 $w=1.65e-07 $l=1.6e-07 $layer=POLY_cond $X=13.43 $Y=1.525
+ $X2=13.43 $Y2=1.365
r230 29 31 363.444 $w=1.8e-07 $l=9.35e-07 $layer=POLY_cond $X=13.43 $Y=1.525
+ $X2=13.43 $Y2=2.46
r231 26 36 33.9972 $w=1.65e-07 $l=1.67332e-07 $layer=POLY_cond $X=13.415
+ $Y=1.205 $X2=13.43 $Y2=1.365
r232 26 28 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=13.415 $Y=1.205
+ $X2=13.415 $Y2=0.81
r233 25 70 2.52859 $w=3.2e-07 $l=2.06126e-07 $layer=POLY_cond $X=12.51 $Y=1.365
+ $X2=12.322 $Y2=1.327
r234 24 36 3.5291 $w=3.2e-07 $l=9e-08 $layer=POLY_cond $X=13.34 $Y=1.365
+ $X2=13.43 $Y2=1.365
r235 24 25 149.67 $w=3.2e-07 $l=8.3e-07 $layer=POLY_cond $X=13.34 $Y=1.365
+ $X2=12.51 $Y2=1.365
r236 22 35 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=12.45 $Y=2.75
+ $X2=12.45 $Y2=2.14
r237 16 70 23.988 $w=2.62e-07 $l=2.43105e-07 $layer=POLY_cond $X=12.425 $Y=1.13
+ $X2=12.322 $Y2=1.327
r238 16 18 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=12.425 $Y=1.13
+ $X2=12.425 $Y2=0.58
r239 5 63 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=11.56
+ $Y=2.54 $X2=11.695 $Y2=2.75
r240 4 48 600 $w=1.7e-07 $l=7.56224e-07 $layer=licon1_PDIFF $count=1 $X=9.98
+ $Y=2.12 $X2=10.27 $Y2=2.745
r241 3 39 300 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_PDIFF $count=2 $X=9.02
+ $Y=2.12 $X2=9.165 $Y2=2.4
r242 2 52 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=10.205
+ $Y=0.37 $X2=10.415 $Y2=0.58
r243 1 75 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=9.27
+ $Y=0.37 $X2=9.415 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_2%A_2611_98# 1 2 9 13 15 17 20 24 28 34 37 41
c77 28 0 7.29682e-20 $X=13.205 $Y=2.105
r78 41 42 2.02521 $w=3.57e-07 $l=1.5e-08 $layer=POLY_cond $X=14.37 $Y=1.427
+ $X2=14.385 $Y2=1.427
r79 35 39 5.40056 $w=3.57e-07 $l=4e-08 $layer=POLY_cond $X=13.895 $Y=1.427
+ $X2=13.935 $Y2=1.427
r80 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.895
+ $Y=1.485 $X2=13.895 $Y2=1.485
r81 32 37 1.36975 $w=3.3e-07 $l=1.68e-07 $layer=LI1_cond $X=13.37 $Y=1.485
+ $X2=13.202 $Y2=1.485
r82 32 34 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=13.37 $Y=1.485
+ $X2=13.895 $Y2=1.485
r83 28 30 24.4249 $w=3.33e-07 $l=7.1e-07 $layer=LI1_cond $X=13.202 $Y=2.105
+ $X2=13.202 $Y2=2.815
r84 26 37 5.13366 $w=3.32e-07 $l=1.65e-07 $layer=LI1_cond $X=13.202 $Y=1.65
+ $X2=13.202 $Y2=1.485
r85 26 28 15.6526 $w=3.33e-07 $l=4.55e-07 $layer=LI1_cond $X=13.202 $Y=1.65
+ $X2=13.202 $Y2=2.105
r86 22 37 5.13366 $w=3.32e-07 $l=1.65997e-07 $layer=LI1_cond $X=13.2 $Y=1.32
+ $X2=13.202 $Y2=1.485
r87 22 24 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=13.2 $Y=1.32
+ $X2=13.2 $Y2=0.635
r88 18 42 18.7718 $w=1.8e-07 $l=2.23e-07 $layer=POLY_cond $X=14.385 $Y=1.65
+ $X2=14.385 $Y2=1.427
r89 18 20 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=14.385 $Y=1.65
+ $X2=14.385 $Y2=2.4
r90 15 41 23.1043 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=14.37 $Y=1.205
+ $X2=14.37 $Y2=1.427
r91 15 17 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=14.37 $Y=1.205
+ $X2=14.37 $Y2=0.76
r92 11 41 58.056 $w=3.57e-07 $l=4.3e-07 $layer=POLY_cond $X=13.94 $Y=1.427
+ $X2=14.37 $Y2=1.427
r93 11 39 0.67507 $w=3.57e-07 $l=5e-09 $layer=POLY_cond $X=13.94 $Y=1.427
+ $X2=13.935 $Y2=1.427
r94 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=13.94 $Y=1.32
+ $X2=13.94 $Y2=0.76
r95 7 39 18.7718 $w=1.8e-07 $l=2.23e-07 $layer=POLY_cond $X=13.935 $Y=1.65
+ $X2=13.935 $Y2=1.427
r96 7 9 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=13.935 $Y=1.65
+ $X2=13.935 $Y2=2.4
r97 2 30 400 $w=1.7e-07 $l=9.17701e-07 $layer=licon1_PDIFF $count=1 $X=13.075
+ $Y=1.96 $X2=13.205 $Y2=2.815
r98 2 28 400 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_PDIFF $count=1 $X=13.075
+ $Y=1.96 $X2=13.205 $Y2=2.105
r99 1 24 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=13.055
+ $Y=0.49 $X2=13.2 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_2%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 39 43 47 51
+ 55 59 63 67 71 73 76 77 79 80 82 83 84 86 91 112 119 124 129 135 138 141 144
+ 147 150 154
c182 55 0 3.47781e-20 $X=8.52 $Y=2.58
r183 153 154 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r184 150 151 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r185 147 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r186 144 145 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r187 141 142 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r188 139 142 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r189 138 139 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r190 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r191 133 154 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=14.64 $Y2=3.33
r192 133 151 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.68 $Y2=3.33
r193 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r194 130 150 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=13.825 $Y=3.33
+ $X2=13.682 $Y2=3.33
r195 130 132 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=13.825 $Y=3.33
+ $X2=14.16 $Y2=3.33
r196 129 153 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=14.445 $Y=3.33
+ $X2=14.662 $Y2=3.33
r197 129 132 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=14.445 $Y=3.33
+ $X2=14.16 $Y2=3.33
r198 128 151 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r199 128 148 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.72 $Y2=3.33
r200 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r201 125 147 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.84 $Y=3.33
+ $X2=12.675 $Y2=3.33
r202 125 127 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=12.84 $Y=3.33
+ $X2=13.2 $Y2=3.33
r203 124 150 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=13.54 $Y=3.33
+ $X2=13.682 $Y2=3.33
r204 124 127 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=13.54 $Y=3.33
+ $X2=13.2 $Y2=3.33
r205 123 148 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r206 123 145 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.28 $Y2=3.33
r207 122 123 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r208 120 144 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.33 $Y=3.33
+ $X2=11.205 $Y2=3.33
r209 120 122 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=11.33 $Y=3.33
+ $X2=12.24 $Y2=3.33
r210 119 147 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.51 $Y=3.33
+ $X2=12.675 $Y2=3.33
r211 119 122 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=12.51 $Y=3.33
+ $X2=12.24 $Y2=3.33
r212 118 145 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r213 117 118 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r214 115 118 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=10.8 $Y2=3.33
r215 114 117 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=10.8 $Y2=3.33
r216 114 115 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r217 112 144 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.08 $Y=3.33
+ $X2=11.205 $Y2=3.33
r218 112 117 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=11.08 $Y=3.33
+ $X2=10.8 $Y2=3.33
r219 111 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r220 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r221 104 107 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r222 104 105 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r223 102 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r224 101 102 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r225 99 102 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=6 $Y2=3.33
r226 99 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r227 98 101 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=6 $Y2=3.33
r228 98 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r229 96 141 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=3.71 $Y2=3.33
r230 96 98 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=4.08 $Y2=3.33
r231 95 139 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r232 95 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r233 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r234 92 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r235 92 94 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r236 91 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=3.33
+ $X2=2.725 $Y2=3.33
r237 91 94 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.56 $Y=3.33
+ $X2=1.2 $Y2=3.33
r238 89 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r239 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r240 86 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r241 86 88 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r242 84 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r243 84 105 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r244 84 107 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r245 82 110 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=8.435 $Y=3.33
+ $X2=8.4 $Y2=3.33
r246 82 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.435 $Y=3.33
+ $X2=8.56 $Y2=3.33
r247 81 114 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=8.685 $Y=3.33
+ $X2=8.88 $Y2=3.33
r248 81 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.685 $Y=3.33
+ $X2=8.56 $Y2=3.33
r249 79 107 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=7.535 $Y=3.33
+ $X2=7.44 $Y2=3.33
r250 79 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.535 $Y=3.33
+ $X2=7.62 $Y2=3.33
r251 78 110 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=7.705 $Y=3.33
+ $X2=8.4 $Y2=3.33
r252 78 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.705 $Y=3.33
+ $X2=7.62 $Y2=3.33
r253 76 101 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=6.095 $Y=3.33
+ $X2=6 $Y2=3.33
r254 76 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.095 $Y=3.33
+ $X2=6.22 $Y2=3.33
r255 75 104 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.345 $Y=3.33
+ $X2=6.48 $Y2=3.33
r256 75 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.345 $Y=3.33
+ $X2=6.22 $Y2=3.33
r257 71 153 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=14.61 $Y=3.245
+ $X2=14.662 $Y2=3.33
r258 71 73 29.3349 $w=3.28e-07 $l=8.4e-07 $layer=LI1_cond $X=14.61 $Y=3.245
+ $X2=14.61 $Y2=2.405
r259 67 70 29.5187 $w=2.83e-07 $l=7.3e-07 $layer=LI1_cond $X=13.682 $Y=2.085
+ $X2=13.682 $Y2=2.815
r260 65 150 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=13.682 $Y=3.245
+ $X2=13.682 $Y2=3.33
r261 65 70 17.3877 $w=2.83e-07 $l=4.3e-07 $layer=LI1_cond $X=13.682 $Y=3.245
+ $X2=13.682 $Y2=2.815
r262 61 147 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.675 $Y=3.245
+ $X2=12.675 $Y2=3.33
r263 61 63 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=12.675 $Y=3.245
+ $X2=12.675 $Y2=2.815
r264 57 144 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.205 $Y=3.245
+ $X2=11.205 $Y2=3.33
r265 57 59 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=11.205 $Y=3.245
+ $X2=11.205 $Y2=2.81
r266 53 83 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.56 $Y=3.245
+ $X2=8.56 $Y2=3.33
r267 53 55 30.655 $w=2.48e-07 $l=6.65e-07 $layer=LI1_cond $X=8.56 $Y=3.245
+ $X2=8.56 $Y2=2.58
r268 49 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.62 $Y=3.245
+ $X2=7.62 $Y2=3.33
r269 49 51 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=7.62 $Y=3.245
+ $X2=7.62 $Y2=2.23
r270 45 77 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.22 $Y=3.245
+ $X2=6.22 $Y2=3.33
r271 45 47 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=6.22 $Y=3.245
+ $X2=6.22 $Y2=2.59
r272 41 141 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.71 $Y=3.245
+ $X2=3.71 $Y2=3.33
r273 41 43 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.71 $Y=3.245
+ $X2=3.71 $Y2=2.78
r274 40 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.89 $Y=3.33
+ $X2=2.725 $Y2=3.33
r275 39 141 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.545 $Y=3.33
+ $X2=3.71 $Y2=3.33
r276 39 40 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.545 $Y=3.33
+ $X2=2.89 $Y2=3.33
r277 35 138 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=3.245
+ $X2=2.725 $Y2=3.33
r278 35 37 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.725 $Y=3.245
+ $X2=2.725 $Y2=2.995
r279 31 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r280 31 33 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.78
r281 10 73 300 $w=1.7e-07 $l=6.28888e-07 $layer=licon1_PDIFF $count=2 $X=14.475
+ $Y=1.84 $X2=14.61 $Y2=2.405
r282 9 70 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=13.52
+ $Y=1.96 $X2=13.705 $Y2=2.815
r283 9 67 400 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_PDIFF $count=1 $X=13.52
+ $Y=1.96 $X2=13.705 $Y2=2.085
r284 8 63 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=12.54
+ $Y=2.54 $X2=12.675 $Y2=2.815
r285 7 59 600 $w=1.7e-07 $l=3.30681e-07 $layer=licon1_PDIFF $count=1 $X=11.11
+ $Y=2.54 $X2=11.245 $Y2=2.81
r286 6 55 600 $w=1.7e-07 $l=7.49466e-07 $layer=licon1_PDIFF $count=1 $X=8.385
+ $Y=1.895 $X2=8.52 $Y2=2.58
r287 5 51 300 $w=1.7e-07 $l=3.6e-07 $layer=licon1_PDIFF $count=2 $X=7.3 $Y=2.315
+ $X2=7.62 $Y2=2.23
r288 4 47 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=6.12
+ $Y=2.315 $X2=6.26 $Y2=2.59
r289 3 43 600 $w=1.7e-07 $l=1.00524e-06 $layer=licon1_PDIFF $count=1 $X=3.575
+ $Y=1.84 $X2=3.71 $Y2=2.78
r290 2 37 600 $w=1.7e-07 $l=7.729e-07 $layer=licon1_PDIFF $count=1 $X=2.515
+ $Y=2.32 $X2=2.725 $Y2=2.995
r291 1 33 600 $w=1.7e-07 $l=5.23163e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=2.32 $X2=0.73 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_2%A_293_464# 1 2 3 4 13 19 21 22 24 25 27 32
+ 33 36 43 45 46 47
c132 27 0 4.72054e-20 $X=4.585 $Y=2.325
c133 24 0 4.46515e-20 $X=2.3 $Y=2.49
c134 22 0 1.77325e-19 $X=1.89 $Y=0.995
c135 19 0 8.84878e-21 $X=1.725 $Y=0.58
r136 47 49 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.75 $Y=2.325
+ $X2=4.75 $Y2=2.495
r137 45 46 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.667 $Y=1.9
+ $X2=4.667 $Y2=2.07
r138 40 43 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=4.505 $Y=0.72
+ $X2=4.665 $Y2=0.72
r139 36 38 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.035 $Y=2.325
+ $X2=3.035 $Y2=2.575
r140 32 47 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.75 $Y=2.24
+ $X2=4.75 $Y2=2.325
r141 32 46 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.75 $Y=2.24
+ $X2=4.75 $Y2=2.07
r142 29 40 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.505 $Y=0.845
+ $X2=4.505 $Y2=0.72
r143 29 45 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=4.505 $Y=0.845
+ $X2=4.505 $Y2=1.9
r144 28 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=2.325
+ $X2=3.035 $Y2=2.325
r145 27 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.585 $Y=2.325
+ $X2=4.75 $Y2=2.325
r146 27 28 95.5775 $w=1.68e-07 $l=1.465e-06 $layer=LI1_cond $X=4.585 $Y=2.325
+ $X2=3.12 $Y2=2.325
r147 26 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=2.575
+ $X2=2.3 $Y2=2.575
r148 25 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.95 $Y=2.575
+ $X2=3.035 $Y2=2.575
r149 25 26 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.95 $Y=2.575
+ $X2=2.385 $Y2=2.575
r150 24 33 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=2.49 $X2=2.3
+ $Y2=2.575
r151 23 24 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=2.3 $Y=1.08
+ $X2=2.3 $Y2=2.49
r152 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.215 $Y=0.995
+ $X2=2.3 $Y2=1.08
r153 21 22 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.215 $Y=0.995
+ $X2=1.89 $Y2=0.995
r154 17 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.725 $Y=0.91
+ $X2=1.89 $Y2=0.995
r155 17 19 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.725 $Y=0.91
+ $X2=1.725 $Y2=0.58
r156 13 33 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.3 $Y=2.785
+ $X2=2.3 $Y2=2.575
r157 13 15 24.2013 $w=2.48e-07 $l=5.25e-07 $layer=LI1_cond $X=2.215 $Y=2.785
+ $X2=1.69 $Y2=2.785
r158 4 49 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=4.605
+ $Y=2.285 $X2=4.75 $Y2=2.495
r159 3 15 600 $w=1.7e-07 $l=5.25595e-07 $layer=licon1_PDIFF $count=1 $X=1.465
+ $Y=2.32 $X2=1.69 $Y2=2.745
r160 2 43 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=4.525
+ $Y=0.405 $X2=4.665 $Y2=0.68
r161 1 19 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.37 $X2=1.725 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_2%A_1587_379# 1 2 9 11 15 18 19
r34 19 21 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=8.68 $Y=2.06 $X2=8.68
+ $Y2=2.15
r35 13 15 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=9.665 $Y=2.145
+ $X2=9.665 $Y2=2.265
r36 12 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.765 $Y=2.06
+ $X2=8.68 $Y2=2.06
r37 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.5 $Y=2.06
+ $X2=9.665 $Y2=2.145
r38 11 12 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=9.5 $Y=2.06
+ $X2=8.765 $Y2=2.06
r39 10 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.235 $Y=2.15
+ $X2=8.07 $Y2=2.15
r40 9 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.595 $Y=2.15
+ $X2=8.68 $Y2=2.15
r41 9 10 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.595 $Y=2.15
+ $X2=8.235 $Y2=2.15
r42 2 15 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=9.53
+ $Y=2.12 $X2=9.665 $Y2=2.265
r43 1 18 300 $w=1.7e-07 $l=3.968e-07 $layer=licon1_PDIFF $count=2 $X=7.935
+ $Y=1.895 $X2=8.07 $Y2=2.23
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_2%Q 1 2 9 13 17 19 20 21 22
c41 20 0 5.67555e-20 $X=14.465 $Y=1.49
r42 28 31 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=14.135 $Y=1.985
+ $X2=14.16 $Y2=1.985
r43 25 31 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=14.54 $Y=1.985
+ $X2=14.16 $Y2=1.985
r44 22 25 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=14.64 $Y=1.985
+ $X2=14.54 $Y2=1.985
r45 21 25 4.15415 $w=4.28e-07 $l=1.55e-07 $layer=LI1_cond $X=14.54 $Y=1.665
+ $X2=14.54 $Y2=1.82
r46 20 21 4.69018 $w=4.28e-07 $l=1.75e-07 $layer=LI1_cond $X=14.54 $Y=1.49
+ $X2=14.54 $Y2=1.665
r47 19 20 8.9189 $w=4.28e-07 $l=1.7e-07 $layer=LI1_cond $X=14.465 $Y=1.32
+ $X2=14.465 $Y2=1.49
r48 17 19 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=14.26 $Y=1.15
+ $X2=14.26 $Y2=1.32
r49 11 28 1.70047 $w=2.8e-07 $l=1.65e-07 $layer=LI1_cond $X=14.135 $Y=2.15
+ $X2=14.135 $Y2=1.985
r50 11 13 10.7013 $w=2.78e-07 $l=2.6e-07 $layer=LI1_cond $X=14.135 $Y=2.15
+ $X2=14.135 $Y2=2.41
r51 7 17 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=14.167 $Y=0.973
+ $X2=14.167 $Y2=1.15
r52 7 9 14.2189 $w=3.53e-07 $l=4.38e-07 $layer=LI1_cond $X=14.167 $Y=0.973
+ $X2=14.167 $Y2=0.535
r53 2 31 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=14.025
+ $Y=1.84 $X2=14.16 $Y2=1.985
r54 2 13 300 $w=1.7e-07 $l=6.33916e-07 $layer=licon1_PDIFF $count=2 $X=14.025
+ $Y=1.84 $X2=14.16 $Y2=2.41
r55 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.015
+ $Y=0.39 $X2=14.155 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_2%VGND 1 2 3 4 5 6 7 8 9 30 34 36 40 44 48 52
+ 54 56 58 59 65 67 72 87 94 107 112 118 121 124 127 130 135 141 143 147
c162 147 0 2.52187e-20 $X=14.64 $Y=0
r163 146 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r164 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r165 139 141 9.39905 $w=6.83e-07 $l=9e-08 $layer=LI1_cond $X=12.24 $Y=0.257
+ $X2=12.33 $Y2=0.257
r166 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r167 137 139 1.30957 $w=6.83e-07 $l=7.5e-08 $layer=LI1_cond $X=12.165 $Y=0.257
+ $X2=12.24 $Y2=0.257
r168 134 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r169 133 137 7.0717 $w=6.83e-07 $l=4.05e-07 $layer=LI1_cond $X=11.76 $Y=0.257
+ $X2=12.165 $Y2=0.257
r170 133 135 9.92288 $w=6.83e-07 $l=1.2e-07 $layer=LI1_cond $X=11.76 $Y=0.257
+ $X2=11.64 $Y2=0.257
r171 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r172 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r173 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r174 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r175 122 125 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.6 $Y2=0
r176 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r177 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r178 116 147 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=14.64 $Y2=0
r179 116 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=13.68 $Y2=0
r180 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r181 113 143 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.805 $Y=0
+ $X2=13.68 $Y2=0
r182 113 115 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=13.805 $Y=0
+ $X2=14.16 $Y2=0
r183 112 146 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=14.515 $Y=0
+ $X2=14.697 $Y2=0
r184 112 115 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=14.515 $Y=0
+ $X2=14.16 $Y2=0
r185 111 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=13.68 $Y2=0
r186 111 140 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=12.24 $Y2=0
r187 110 141 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=13.2 $Y=0
+ $X2=12.33 $Y2=0
r188 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r189 107 143 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.555 $Y=0
+ $X2=13.68 $Y2=0
r190 107 110 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=13.555 $Y=0
+ $X2=13.2 $Y2=0
r191 106 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r192 105 135 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=11.28 $Y=0
+ $X2=11.64 $Y2=0
r193 105 106 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r194 103 106 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=11.28 $Y2=0
r195 103 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r196 102 105 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=9.36 $Y=0
+ $X2=11.28 $Y2=0
r197 102 103 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r198 100 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.02 $Y=0
+ $X2=8.855 $Y2=0
r199 100 102 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=9.02 $Y=0
+ $X2=9.36 $Y2=0
r200 98 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r201 98 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r202 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r203 95 127 11.2921 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=8.01 $Y=0 $X2=7.76
+ $Y2=0
r204 95 97 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=8.01 $Y=0 $X2=8.4
+ $Y2=0
r205 94 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.69 $Y=0
+ $X2=8.855 $Y2=0
r206 94 97 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=8.69 $Y=0 $X2=8.4
+ $Y2=0
r207 89 92 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r208 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r209 87 127 11.2921 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=7.51 $Y=0 $X2=7.76
+ $Y2=0
r210 87 92 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=7.51 $Y=0 $X2=7.44
+ $Y2=0
r211 86 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r212 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r213 83 86 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r214 83 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r215 82 85 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r216 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r217 80 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.85 $Y=0
+ $X2=3.685 $Y2=0
r218 80 82 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.85 $Y=0 $X2=4.08
+ $Y2=0
r219 79 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=2.64 $Y2=0
r220 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r221 76 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r222 76 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r223 75 78 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r224 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r225 73 118 10.6558 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=1.07 $Y=0
+ $X2=0.842 $Y2=0
r226 73 75 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.07 $Y=0 $X2=1.2
+ $Y2=0
r227 72 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.46 $Y=0
+ $X2=2.625 $Y2=0
r228 72 78 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.46 $Y=0 $X2=2.16
+ $Y2=0
r229 70 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r230 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r231 67 118 10.6558 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.842 $Y2=0
r232 67 69 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r233 65 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r234 65 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.48
+ $Y2=0
r235 65 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r236 61 89 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=6.46 $Y=0 $X2=6.48
+ $Y2=0
r237 59 85 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=6.13 $Y=0 $X2=6
+ $Y2=0
r238 58 63 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.295 $Y=0
+ $X2=6.295 $Y2=0.275
r239 58 61 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.295 $Y=0 $X2=6.46
+ $Y2=0
r240 58 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.295 $Y=0 $X2=6.13
+ $Y2=0
r241 54 146 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=14.64 $Y=0.085
+ $X2=14.697 $Y2=0
r242 54 56 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=14.64 $Y=0.085
+ $X2=14.64 $Y2=0.525
r243 50 143 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.68 $Y=0.085
+ $X2=13.68 $Y2=0
r244 50 52 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=13.68 $Y=0.085
+ $X2=13.68 $Y2=0.535
r245 46 130 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.855 $Y=0.085
+ $X2=8.855 $Y2=0
r246 46 48 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=8.855 $Y=0.085
+ $X2=8.855 $Y2=0.53
r247 42 127 2.07448 $w=5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.76 $Y=0.085
+ $X2=7.76 $Y2=0
r248 42 44 10.2863 $w=4.98e-07 $l=4.3e-07 $layer=LI1_cond $X=7.76 $Y=0.085
+ $X2=7.76 $Y2=0.515
r249 38 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=0.085
+ $X2=3.685 $Y2=0
r250 38 40 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.685 $Y=0.085
+ $X2=3.685 $Y2=0.515
r251 37 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.79 $Y=0
+ $X2=2.625 $Y2=0
r252 36 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.52 $Y=0
+ $X2=3.685 $Y2=0
r253 36 37 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.52 $Y=0 $X2=2.79
+ $Y2=0
r254 32 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.625 $Y=0.085
+ $X2=2.625 $Y2=0
r255 32 34 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=2.625 $Y=0.085
+ $X2=2.625 $Y2=0.545
r256 28 118 1.82608 $w=4.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.842 $Y=0.085
+ $X2=0.842 $Y2=0
r257 28 30 11.3036 $w=4.53e-07 $l=4.3e-07 $layer=LI1_cond $X=0.842 $Y=0.085
+ $X2=0.842 $Y2=0.515
r258 9 56 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=14.445
+ $Y=0.39 $X2=14.6 $Y2=0.525
r259 8 52 91 $w=1.7e-07 $l=2.51496e-07 $layer=licon1_NDIFF $count=2 $X=13.49
+ $Y=0.49 $X2=13.72 $Y2=0.535
r260 7 137 91 $w=1.7e-07 $l=5.67891e-07 $layer=licon1_NDIFF $count=2 $X=11.665
+ $Y=0.37 $X2=12.165 $Y2=0.515
r261 6 48 182 $w=1.7e-07 $l=2.89137e-07 $layer=licon1_NDIFF $count=1 $X=8.635
+ $Y=0.37 $X2=8.855 $Y2=0.53
r262 5 44 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=7.535
+ $Y=0.37 $X2=7.76 $Y2=0.515
r263 4 63 182 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_NDIFF $count=1 $X=6.075
+ $Y=0.405 $X2=6.295 $Y2=0.275
r264 3 40 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=3.475
+ $Y=0.37 $X2=3.685 $Y2=0.515
r265 2 34 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=0.37 $X2=2.625 $Y2=0.545
r266 1 30 182 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.84 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSTP_2%A_1641_74# 1 2 9 11 12 14
c42 12 0 1.09822e-19 $X=8.51 $Y=0.97
c43 11 0 3.01101e-20 $X=9.75 $Y=0.97
r44 14 16 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=9.915 $Y=0.81
+ $X2=9.915 $Y2=0.97
r45 11 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.75 $Y=0.97
+ $X2=9.915 $Y2=0.97
r46 11 12 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=9.75 $Y=0.97
+ $X2=8.51 $Y2=0.97
r47 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.345 $Y=0.885
+ $X2=8.51 $Y2=0.97
r48 7 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.345 $Y=0.885
+ $X2=8.345 $Y2=0.515
r49 2 14 182 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_NDIFF $count=1 $X=9.775
+ $Y=0.37 $X2=9.915 $Y2=0.81
r50 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.205
+ $Y=0.37 $X2=8.345 $Y2=0.515
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
X0 VGND a_179_48# X VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X1 a_179_48# D VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X2 VPWR a_179_48# X VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X3 a_647_74# D VGND VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X4 VGND B_N a_503_48# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X5 VPWR a_27_74# a_179_48# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X6 a_27_74# A_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X7 VPWR C a_179_48# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X8 a_455_74# a_503_48# a_533_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X9 a_179_48# a_27_74# a_455_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X10 a_179_48# a_503_48# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X11 VPWR B_N a_503_48# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X12 a_533_74# C a_647_74# VNB sky130_fd_pr__nfet_01v8_lvt w=640000u l=150000u
X13 a_27_74# A_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
.ends

* File: sky130_fd_sc_ms__xnor2_1.spice
* Created: Wed Sep  2 12:33:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__xnor2_1.pex.spice"
.subckt sky130_fd_sc_ms__xnor2_1  VNB VPB B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1006 A_112_119# N_A_M1006_g N_VGND_M1006_s VNB NLOWVT L=0.15 W=0.64 AD=0.0672
+ AS=0.176 PD=0.85 PS=1.83 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75000.2 SB=75000.6
+ A=0.096 P=1.58 MULT=1
MM1002 N_A_141_385#_M1002_d N_B_M1002_g A_112_119# VNB NLOWVT L=0.15 W=0.64
+ AD=0.176 AS=0.0672 PD=1.83 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_VGND_M1000_d N_A_M1000_g N_A_293_74#_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.182 AS=0.2035 PD=1.345 PS=2.03 NRD=12.156 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1008 N_A_293_74#_M1008_d N_B_M1008_g N_VGND_M1000_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.182 PD=1.02 PS=1.345 NRD=0 NRS=12.972 M=1 R=4.93333 SA=75000.8
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1004 N_Y_M1004_d N_A_141_385#_M1004_g N_A_293_74#_M1008_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2294 AS=0.1036 PD=2.1 PS=1.02 NRD=4.044 NRS=0 M=1 R=4.93333
+ SA=75001.2 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1007 N_A_141_385#_M1007_d N_A_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.2772 PD=1.11 PS=2.34 NRD=0 NRS=10.5395 M=1 R=4.66667 SA=90000.2
+ SB=90002.4 A=0.1512 P=2.04 MULT=1
MM1001 N_VPWR_M1001_d N_B_M1001_g N_A_141_385#_M1007_d VPB PSHORT L=0.18 W=0.84
+ AD=0.234107 AS=0.1134 PD=1.44 PS=1.11 NRD=147.75 NRS=0 M=1 R=4.66667
+ SA=90000.7 SB=90001.9 A=0.1512 P=2.04 MULT=1
MM1003 A_379_368# N_A_M1003_g N_VPWR_M1001_d VPB PSHORT L=0.18 W=1.12 AD=0.1344
+ AS=0.312143 PD=1.36 PS=1.92 NRD=11.426 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1005 N_Y_M1005_d N_B_M1005_g A_379_368# VPB PSHORT L=0.18 W=1.12 AD=0.2184
+ AS=0.1344 PD=1.51 PS=1.36 NRD=11.426 NRS=11.426 M=1 R=6.22222 SA=90001.5
+ SB=90000.8 A=0.2016 P=2.6 MULT=1
MM1009 N_VPWR_M1009_d N_A_141_385#_M1009_g N_Y_M1005_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.2184 PD=2.8 PS=1.51 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9564 P=11.2
*
.include "sky130_fd_sc_ms__xnor2_1.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__nor3b_2.pxi.spice
* Created: Wed Sep  2 12:16:24 2020
* 
x_PM_SKY130_FD_SC_MS__NOR3B_2%C_N N_C_N_M1003_g N_C_N_M1008_g C_N N_C_N_c_82_n
+ PM_SKY130_FD_SC_MS__NOR3B_2%C_N
x_PM_SKY130_FD_SC_MS__NOR3B_2%A_27_392# N_A_27_392#_M1008_s N_A_27_392#_M1003_s
+ N_A_27_392#_c_114_n N_A_27_392#_M1000_g N_A_27_392#_M1005_g
+ N_A_27_392#_c_116_n N_A_27_392#_M1012_g N_A_27_392#_M1006_g
+ N_A_27_392#_c_118_n N_A_27_392#_c_126_n N_A_27_392#_c_127_n
+ N_A_27_392#_c_119_n N_A_27_392#_c_120_n N_A_27_392#_c_121_n
+ N_A_27_392#_c_122_n N_A_27_392#_c_123_n PM_SKY130_FD_SC_MS__NOR3B_2%A_27_392#
x_PM_SKY130_FD_SC_MS__NOR3B_2%B N_B_M1001_g N_B_M1007_g N_B_M1013_g N_B_M1010_g
+ B N_B_c_196_n N_B_c_197_n PM_SKY130_FD_SC_MS__NOR3B_2%B
x_PM_SKY130_FD_SC_MS__NOR3B_2%A N_A_M1002_g N_A_M1009_g N_A_M1004_g N_A_M1011_g
+ A A A N_A_c_248_n PM_SKY130_FD_SC_MS__NOR3B_2%A
x_PM_SKY130_FD_SC_MS__NOR3B_2%VPWR N_VPWR_M1003_d N_VPWR_M1009_s N_VPWR_M1011_s
+ N_VPWR_c_293_n N_VPWR_c_294_n N_VPWR_c_295_n N_VPWR_c_296_n VPWR
+ N_VPWR_c_297_n N_VPWR_c_298_n N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_301_n
+ N_VPWR_c_292_n PM_SKY130_FD_SC_MS__NOR3B_2%VPWR
x_PM_SKY130_FD_SC_MS__NOR3B_2%A_227_368# N_A_227_368#_M1005_s
+ N_A_227_368#_M1006_s N_A_227_368#_M1010_s N_A_227_368#_c_348_n
+ N_A_227_368#_c_349_n N_A_227_368#_c_350_n N_A_227_368#_c_351_n
+ N_A_227_368#_c_352_n N_A_227_368#_c_353_n N_A_227_368#_c_354_n
+ PM_SKY130_FD_SC_MS__NOR3B_2%A_227_368#
x_PM_SKY130_FD_SC_MS__NOR3B_2%Y N_Y_M1000_s N_Y_M1001_d N_Y_M1002_d N_Y_M1005_d
+ N_Y_c_392_n N_Y_c_393_n N_Y_c_394_n N_Y_c_395_n N_Y_c_396_n N_Y_c_397_n
+ N_Y_c_398_n Y Y N_Y_c_399_n PM_SKY130_FD_SC_MS__NOR3B_2%Y
x_PM_SKY130_FD_SC_MS__NOR3B_2%A_498_368# N_A_498_368#_M1007_d
+ N_A_498_368#_M1009_d N_A_498_368#_c_451_n N_A_498_368#_c_463_n
+ N_A_498_368#_c_452_n N_A_498_368#_c_456_n
+ PM_SKY130_FD_SC_MS__NOR3B_2%A_498_368#
x_PM_SKY130_FD_SC_MS__NOR3B_2%VGND N_VGND_M1008_d N_VGND_M1012_d N_VGND_M1013_s
+ N_VGND_M1004_s N_VGND_c_478_n N_VGND_c_479_n N_VGND_c_480_n VGND
+ N_VGND_c_481_n N_VGND_c_482_n N_VGND_c_483_n N_VGND_c_484_n N_VGND_c_485_n
+ N_VGND_c_486_n N_VGND_c_487_n N_VGND_c_488_n PM_SKY130_FD_SC_MS__NOR3B_2%VGND
cc_1 VNB N_C_N_M1008_g 0.045041f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.69
cc_2 VNB C_N 0.00302227f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_3 VNB N_C_N_c_82_n 0.0212084f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_4 VNB N_A_27_392#_c_114_n 0.0176119f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.69
cc_5 VNB N_A_27_392#_M1005_g 0.00721961f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.615
cc_6 VNB N_A_27_392#_c_116_n 0.0192011f $X=-0.19 $Y=-0.245 $X2=0.582 $Y2=1.45
cc_7 VNB N_A_27_392#_M1006_g 0.00705856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_392#_c_118_n 0.0335242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_392#_c_119_n 0.012887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_392#_c_120_n 0.0117556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_392#_c_121_n 0.0179582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_392#_c_122_n 0.00730665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_392#_c_123_n 0.0789656f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B_M1001_g 0.0259199f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.46
cc_15 VNB N_B_M1013_g 0.0317091f $X=-0.19 $Y=-0.245 $X2=0.582 $Y2=1.615
cc_16 VNB B 0.00231327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B_c_196_n 0.0307078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B_c_197_n 0.0248648f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_M1002_g 0.0324424f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.46
cc_20 VNB N_A_M1004_g 0.0324934f $X=-0.19 $Y=-0.245 $X2=0.582 $Y2=1.615
cc_21 VNB A 0.0211459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_c_248_n 0.043067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_292_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_392_n 0.00228526f $X=-0.19 $Y=-0.245 $X2=0.582 $Y2=1.78
cc_25 VNB N_Y_c_393_n 0.00408474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_394_n 0.00195796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_395_n 0.0156942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_396_n 0.00261132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_397_n 0.0142336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_398_n 0.00325261f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_399_n 5.03809e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_478_n 0.00890068f $X=-0.19 $Y=-0.245 $X2=0.582 $Y2=1.78
cc_33 VNB N_VGND_c_479_n 0.0120457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_480_n 0.0420237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_481_n 0.0190372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_482_n 0.0166972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_483_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_484_n 0.0172153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_485_n 0.020831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_486_n 0.0137748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_487_n 0.0243803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_488_n 0.265014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_C_N_M1003_g 0.0323753f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=2.46
cc_44 VPB C_N 0.00255821f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_45 VPB N_C_N_c_82_n 0.0140189f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_46 VPB N_A_27_392#_M1005_g 0.0265469f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_47 VPB N_A_27_392#_M1006_g 0.0217399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_27_392#_c_126_n 0.00691932f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_A_27_392#_c_127_n 0.0367495f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_50 VPB N_A_27_392#_c_121_n 0.0137991f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_51 VPB N_B_M1007_g 0.0207433f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=0.69
cc_52 VPB N_B_M1010_g 0.0250876f $X=-0.19 $Y=1.66 $X2=0.582 $Y2=1.78
cc_53 VPB B 0.00657804f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_B_c_196_n 0.00423142f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_B_c_197_n 0.0106168f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_A_M1009_g 0.0253599f $X=-0.19 $Y=1.66 $X2=0.5 $Y2=0.69
cc_57 VPB N_A_M1011_g 0.0246355f $X=-0.19 $Y=1.66 $X2=0.582 $Y2=1.78
cc_58 VPB A 0.0151336f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_A_c_248_n 0.0069886f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_293_n 0.0179682f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_61 VPB N_VPWR_c_294_n 0.0118814f $X=-0.19 $Y=1.66 $X2=0.72 $Y2=1.615
cc_62 VPB N_VPWR_c_295_n 0.0107811f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_296_n 0.0499696f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_297_n 0.0176729f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_298_n 0.0611154f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_299_n 0.018048f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_300_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_301_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_292_n 0.0817021f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_70 VPB N_A_227_368#_c_348_n 0.0130846f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_71 VPB N_A_227_368#_c_349_n 0.00192243f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_72 VPB N_A_227_368#_c_350_n 0.00411341f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_73 VPB N_A_227_368#_c_351_n 0.0103669f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_74 VPB N_A_227_368#_c_352_n 0.00615921f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_75 VPB N_A_227_368#_c_353_n 0.00560044f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_76 VPB N_A_227_368#_c_354_n 0.00181992f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_77 VPB N_Y_c_393_n 0.00394095f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_78 VPB N_A_498_368#_c_451_n 0.0173379f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_79 VPB N_A_498_368#_c_452_n 0.00202354f $X=-0.19 $Y=1.66 $X2=0.59 $Y2=1.615
cc_80 N_C_N_M1008_g N_A_27_392#_c_114_n 0.0286f $X=0.5 $Y=0.69 $X2=0 $Y2=0
cc_81 C_N N_A_27_392#_M1005_g 0.0040108f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_82 N_C_N_c_82_n N_A_27_392#_M1005_g 0.00284553f $X=0.59 $Y=1.615 $X2=0 $Y2=0
cc_83 N_C_N_M1008_g N_A_27_392#_c_118_n 0.0122317f $X=0.5 $Y=0.69 $X2=0 $Y2=0
cc_84 N_C_N_M1003_g N_A_27_392#_c_126_n 7.04192e-19 $X=0.5 $Y=2.46 $X2=0 $Y2=0
cc_85 N_C_N_M1008_g N_A_27_392#_c_119_n 0.0117984f $X=0.5 $Y=0.69 $X2=0 $Y2=0
cc_86 C_N N_A_27_392#_c_119_n 0.0287637f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_87 N_C_N_c_82_n N_A_27_392#_c_119_n 0.0040948f $X=0.59 $Y=1.615 $X2=0 $Y2=0
cc_88 N_C_N_M1008_g N_A_27_392#_c_120_n 0.0042843f $X=0.5 $Y=0.69 $X2=0 $Y2=0
cc_89 C_N N_A_27_392#_c_120_n 0.00199562f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_90 N_C_N_c_82_n N_A_27_392#_c_120_n 7.25782e-19 $X=0.59 $Y=1.615 $X2=0 $Y2=0
cc_91 N_C_N_M1008_g N_A_27_392#_c_121_n 0.0040915f $X=0.5 $Y=0.69 $X2=0 $Y2=0
cc_92 C_N N_A_27_392#_c_121_n 0.0251881f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_93 N_C_N_c_82_n N_A_27_392#_c_121_n 0.0118711f $X=0.59 $Y=1.615 $X2=0 $Y2=0
cc_94 N_C_N_M1008_g N_A_27_392#_c_122_n 0.00105106f $X=0.5 $Y=0.69 $X2=0 $Y2=0
cc_95 C_N N_A_27_392#_c_122_n 0.00801071f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_96 C_N N_A_27_392#_c_123_n 6.87608e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_97 N_C_N_c_82_n N_A_27_392#_c_123_n 0.00557301f $X=0.59 $Y=1.615 $X2=0 $Y2=0
cc_98 N_C_N_M1003_g N_VPWR_c_293_n 0.0214472f $X=0.5 $Y=2.46 $X2=0 $Y2=0
cc_99 C_N N_VPWR_c_293_n 0.0233068f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_100 N_C_N_c_82_n N_VPWR_c_293_n 0.00384378f $X=0.59 $Y=1.615 $X2=0 $Y2=0
cc_101 N_C_N_M1003_g N_VPWR_c_297_n 0.00460063f $X=0.5 $Y=2.46 $X2=0 $Y2=0
cc_102 N_C_N_M1003_g N_VPWR_c_292_n 0.00912278f $X=0.5 $Y=2.46 $X2=0 $Y2=0
cc_103 N_C_N_M1003_g N_A_227_368#_c_348_n 0.00506032f $X=0.5 $Y=2.46 $X2=0 $Y2=0
cc_104 N_C_N_M1003_g N_A_227_368#_c_350_n 6.0406e-19 $X=0.5 $Y=2.46 $X2=0 $Y2=0
cc_105 N_C_N_M1008_g N_VGND_c_478_n 0.00683336f $X=0.5 $Y=0.69 $X2=0 $Y2=0
cc_106 N_C_N_M1008_g N_VGND_c_481_n 0.00434272f $X=0.5 $Y=0.69 $X2=0 $Y2=0
cc_107 N_C_N_M1008_g N_VGND_c_488_n 0.00824987f $X=0.5 $Y=0.69 $X2=0 $Y2=0
cc_108 N_A_27_392#_c_116_n N_B_M1001_g 0.00650474f $X=1.515 $Y=1.22 $X2=0 $Y2=0
cc_109 N_A_27_392#_c_123_n N_B_M1001_g 0.0204061f $X=1.515 $Y=1.385 $X2=0 $Y2=0
cc_110 N_A_27_392#_c_123_n B 0.00131605f $X=1.515 $Y=1.385 $X2=0 $Y2=0
cc_111 N_A_27_392#_M1006_g N_B_c_196_n 0.0204061f $X=1.95 $Y=2.4 $X2=0 $Y2=0
cc_112 N_A_27_392#_M1005_g N_VPWR_c_293_n 0.00262876f $X=1.5 $Y=2.4 $X2=0 $Y2=0
cc_113 N_A_27_392#_c_126_n N_VPWR_c_293_n 0.0349444f $X=0.222 $Y=2.087 $X2=0
+ $Y2=0
cc_114 N_A_27_392#_c_119_n N_VPWR_c_293_n 0.00174444f $X=1.005 $Y=1.195 $X2=0
+ $Y2=0
cc_115 N_A_27_392#_c_127_n N_VPWR_c_297_n 0.0121815f $X=0.275 $Y=2.115 $X2=0
+ $Y2=0
cc_116 N_A_27_392#_M1005_g N_VPWR_c_298_n 0.00333896f $X=1.5 $Y=2.4 $X2=0 $Y2=0
cc_117 N_A_27_392#_M1006_g N_VPWR_c_298_n 0.00333896f $X=1.95 $Y=2.4 $X2=0 $Y2=0
cc_118 N_A_27_392#_M1005_g N_VPWR_c_292_n 0.00427818f $X=1.5 $Y=2.4 $X2=0 $Y2=0
cc_119 N_A_27_392#_M1006_g N_VPWR_c_292_n 0.00422796f $X=1.95 $Y=2.4 $X2=0 $Y2=0
cc_120 N_A_27_392#_c_127_n N_VPWR_c_292_n 0.0100828f $X=0.275 $Y=2.115 $X2=0
+ $Y2=0
cc_121 N_A_27_392#_M1005_g N_A_227_368#_c_348_n 0.0170023f $X=1.5 $Y=2.4 $X2=0
+ $Y2=0
cc_122 N_A_27_392#_M1006_g N_A_227_368#_c_348_n 7.21661e-19 $X=1.95 $Y=2.4 $X2=0
+ $Y2=0
cc_123 N_A_27_392#_c_122_n N_A_227_368#_c_348_n 0.0136266f $X=1.17 $Y=1.195
+ $X2=0 $Y2=0
cc_124 N_A_27_392#_c_123_n N_A_227_368#_c_348_n 0.00490664f $X=1.515 $Y=1.385
+ $X2=0 $Y2=0
cc_125 N_A_27_392#_M1005_g N_A_227_368#_c_349_n 0.0116345f $X=1.5 $Y=2.4 $X2=0
+ $Y2=0
cc_126 N_A_27_392#_M1006_g N_A_227_368#_c_349_n 0.0116345f $X=1.95 $Y=2.4 $X2=0
+ $Y2=0
cc_127 N_A_27_392#_M1005_g N_A_227_368#_c_350_n 0.00291744f $X=1.5 $Y=2.4 $X2=0
+ $Y2=0
cc_128 N_A_27_392#_M1005_g N_A_227_368#_c_351_n 7.23423e-19 $X=1.5 $Y=2.4 $X2=0
+ $Y2=0
cc_129 N_A_27_392#_M1006_g N_A_227_368#_c_351_n 0.0161868f $X=1.95 $Y=2.4 $X2=0
+ $Y2=0
cc_130 N_A_27_392#_M1006_g N_A_227_368#_c_354_n 0.001916f $X=1.95 $Y=2.4 $X2=0
+ $Y2=0
cc_131 N_A_27_392#_c_122_n N_Y_M1000_s 0.00206393f $X=1.17 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_132 N_A_27_392#_c_114_n N_Y_c_392_n 0.00474752f $X=1.07 $Y=1.22 $X2=0 $Y2=0
cc_133 N_A_27_392#_c_116_n N_Y_c_393_n 0.00123263f $X=1.515 $Y=1.22 $X2=0 $Y2=0
cc_134 N_A_27_392#_M1006_g N_Y_c_393_n 0.00795747f $X=1.95 $Y=2.4 $X2=0 $Y2=0
cc_135 N_A_27_392#_c_122_n N_Y_c_393_n 0.0195623f $X=1.17 $Y=1.195 $X2=0 $Y2=0
cc_136 N_A_27_392#_c_123_n N_Y_c_393_n 0.0295116f $X=1.515 $Y=1.385 $X2=0 $Y2=0
cc_137 N_A_27_392#_c_123_n N_Y_c_397_n 0.0112113f $X=1.515 $Y=1.385 $X2=0 $Y2=0
cc_138 N_A_27_392#_c_114_n N_Y_c_399_n 0.00268071f $X=1.07 $Y=1.22 $X2=0 $Y2=0
cc_139 N_A_27_392#_c_116_n N_Y_c_399_n 0.0232602f $X=1.515 $Y=1.22 $X2=0 $Y2=0
cc_140 N_A_27_392#_c_122_n N_Y_c_399_n 0.0171358f $X=1.17 $Y=1.195 $X2=0 $Y2=0
cc_141 N_A_27_392#_c_123_n N_Y_c_399_n 0.00364771f $X=1.515 $Y=1.385 $X2=0 $Y2=0
cc_142 N_A_27_392#_c_114_n N_VGND_c_478_n 0.00538033f $X=1.07 $Y=1.22 $X2=0
+ $Y2=0
cc_143 N_A_27_392#_c_118_n N_VGND_c_478_n 0.0232729f $X=0.285 $Y=0.515 $X2=0
+ $Y2=0
cc_144 N_A_27_392#_c_119_n N_VGND_c_478_n 0.0261348f $X=1.005 $Y=1.195 $X2=0
+ $Y2=0
cc_145 N_A_27_392#_c_118_n N_VGND_c_481_n 0.0161257f $X=0.285 $Y=0.515 $X2=0
+ $Y2=0
cc_146 N_A_27_392#_c_114_n N_VGND_c_484_n 0.00434272f $X=1.07 $Y=1.22 $X2=0
+ $Y2=0
cc_147 N_A_27_392#_c_116_n N_VGND_c_484_n 0.00383152f $X=1.515 $Y=1.22 $X2=0
+ $Y2=0
cc_148 N_A_27_392#_c_114_n N_VGND_c_485_n 4.13256e-19 $X=1.07 $Y=1.22 $X2=0
+ $Y2=0
cc_149 N_A_27_392#_c_116_n N_VGND_c_485_n 0.00815797f $X=1.515 $Y=1.22 $X2=0
+ $Y2=0
cc_150 N_A_27_392#_c_123_n N_VGND_c_485_n 8.53107e-19 $X=1.515 $Y=1.385 $X2=0
+ $Y2=0
cc_151 N_A_27_392#_c_114_n N_VGND_c_488_n 0.00821461f $X=1.07 $Y=1.22 $X2=0
+ $Y2=0
cc_152 N_A_27_392#_c_116_n N_VGND_c_488_n 0.00367677f $X=1.515 $Y=1.22 $X2=0
+ $Y2=0
cc_153 N_A_27_392#_c_118_n N_VGND_c_488_n 0.013291f $X=0.285 $Y=0.515 $X2=0
+ $Y2=0
cc_154 B N_A_M1009_g 4.34161e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_155 N_B_M1010_g A 3.94742e-19 $X=2.85 $Y=2.4 $X2=0 $Y2=0
cc_156 B A 0.0329499f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_157 N_B_c_197_n A 0.00149566f $X=3.11 $Y=1.515 $X2=0 $Y2=0
cc_158 B N_A_c_248_n 3.07261e-19 $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_159 N_B_c_197_n N_A_c_248_n 0.00878683f $X=3.11 $Y=1.515 $X2=0 $Y2=0
cc_160 N_B_M1010_g N_VPWR_c_294_n 8.93777e-19 $X=2.85 $Y=2.4 $X2=0 $Y2=0
cc_161 N_B_M1007_g N_VPWR_c_298_n 0.00333926f $X=2.4 $Y=2.4 $X2=0 $Y2=0
cc_162 N_B_M1010_g N_VPWR_c_298_n 0.00333926f $X=2.85 $Y=2.4 $X2=0 $Y2=0
cc_163 N_B_M1007_g N_VPWR_c_292_n 0.00422798f $X=2.4 $Y=2.4 $X2=0 $Y2=0
cc_164 N_B_M1010_g N_VPWR_c_292_n 0.0042782f $X=2.85 $Y=2.4 $X2=0 $Y2=0
cc_165 N_B_M1007_g N_A_227_368#_c_351_n 7.5548e-19 $X=2.4 $Y=2.4 $X2=0 $Y2=0
cc_166 N_B_M1007_g N_A_227_368#_c_352_n 0.0139518f $X=2.4 $Y=2.4 $X2=0 $Y2=0
cc_167 N_B_M1010_g N_A_227_368#_c_352_n 0.0149887f $X=2.85 $Y=2.4 $X2=0 $Y2=0
cc_168 N_B_M1001_g N_Y_c_393_n 0.00287038f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_169 N_B_M1001_g N_Y_c_394_n 3.94489e-19 $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_170 N_B_M1013_g N_Y_c_394_n 3.98786e-19 $X=2.815 $Y=0.74 $X2=0 $Y2=0
cc_171 N_B_M1013_g N_Y_c_395_n 0.0148202f $X=2.815 $Y=0.74 $X2=0 $Y2=0
cc_172 B N_Y_c_395_n 0.036025f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_173 N_B_c_196_n N_Y_c_395_n 0.00851701f $X=2.94 $Y=1.515 $X2=0 $Y2=0
cc_174 N_B_M1001_g N_Y_c_397_n 0.0232011f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_175 B N_Y_c_398_n 0.00637318f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_176 N_B_c_196_n N_Y_c_398_n 0.00344949f $X=2.94 $Y=1.515 $X2=0 $Y2=0
cc_177 N_B_M1010_g N_A_498_368#_c_451_n 0.0150541f $X=2.85 $Y=2.4 $X2=0 $Y2=0
cc_178 B N_A_498_368#_c_451_n 0.0356032f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_179 N_B_c_197_n N_A_498_368#_c_451_n 0.00172015f $X=3.11 $Y=1.515 $X2=0 $Y2=0
cc_180 N_B_M1007_g N_A_498_368#_c_456_n 0.0133055f $X=2.4 $Y=2.4 $X2=0 $Y2=0
cc_181 N_B_M1010_g N_A_498_368#_c_456_n 0.0167082f $X=2.85 $Y=2.4 $X2=0 $Y2=0
cc_182 B N_A_498_368#_c_456_n 0.0135427f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_183 N_B_c_196_n N_A_498_368#_c_456_n 0.0013974f $X=2.94 $Y=1.515 $X2=0 $Y2=0
cc_184 N_B_M1001_g N_VGND_c_485_n 0.00799625f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_185 N_B_M1013_g N_VGND_c_485_n 3.93732e-19 $X=2.815 $Y=0.74 $X2=0 $Y2=0
cc_186 N_B_M1001_g N_VGND_c_486_n 0.00230732f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_187 N_B_M1013_g N_VGND_c_486_n 0.00230732f $X=2.815 $Y=0.74 $X2=0 $Y2=0
cc_188 N_B_M1001_g N_VGND_c_487_n 4.40756e-19 $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_189 N_B_M1013_g N_VGND_c_487_n 0.0111471f $X=2.815 $Y=0.74 $X2=0 $Y2=0
cc_190 N_B_M1001_g N_VGND_c_488_n 0.00367737f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_191 N_B_M1013_g N_VGND_c_488_n 0.00752925f $X=2.815 $Y=0.74 $X2=0 $Y2=0
cc_192 N_A_M1009_g N_VPWR_c_294_n 0.0145968f $X=3.85 $Y=2.4 $X2=0 $Y2=0
cc_193 N_A_M1011_g N_VPWR_c_294_n 5.58229e-19 $X=4.3 $Y=2.4 $X2=0 $Y2=0
cc_194 N_A_M1011_g N_VPWR_c_296_n 0.00376978f $X=4.3 $Y=2.4 $X2=0 $Y2=0
cc_195 A N_VPWR_c_296_n 0.0210862f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_196 N_A_M1009_g N_VPWR_c_299_n 0.00460063f $X=3.85 $Y=2.4 $X2=0 $Y2=0
cc_197 N_A_M1011_g N_VPWR_c_299_n 0.005209f $X=4.3 $Y=2.4 $X2=0 $Y2=0
cc_198 N_A_M1009_g N_VPWR_c_292_n 0.00908554f $X=3.85 $Y=2.4 $X2=0 $Y2=0
cc_199 N_A_M1011_g N_VPWR_c_292_n 0.00985654f $X=4.3 $Y=2.4 $X2=0 $Y2=0
cc_200 N_A_M1009_g N_A_227_368#_c_352_n 6.0406e-19 $X=3.85 $Y=2.4 $X2=0 $Y2=0
cc_201 N_A_M1009_g N_A_227_368#_c_353_n 0.00106876f $X=3.85 $Y=2.4 $X2=0 $Y2=0
cc_202 N_A_M1002_g N_Y_c_395_n 0.0148141f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_203 A N_Y_c_395_n 0.0465213f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_204 N_A_c_248_n N_Y_c_395_n 0.00449551f $X=4.3 $Y=1.515 $X2=0 $Y2=0
cc_205 N_A_M1002_g N_Y_c_396_n 4.55721e-19 $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_206 N_A_M1004_g N_Y_c_396_n 4.75407e-19 $X=4.285 $Y=0.74 $X2=0 $Y2=0
cc_207 N_A_M1009_g N_A_498_368#_c_451_n 0.0163793f $X=3.85 $Y=2.4 $X2=0 $Y2=0
cc_208 A N_A_498_368#_c_451_n 0.0351003f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_209 N_A_c_248_n N_A_498_368#_c_451_n 2.76642e-19 $X=4.3 $Y=1.515 $X2=0 $Y2=0
cc_210 N_A_M1011_g N_A_498_368#_c_463_n 0.00249027f $X=4.3 $Y=2.4 $X2=0 $Y2=0
cc_211 A N_A_498_368#_c_463_n 0.0189743f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_212 N_A_c_248_n N_A_498_368#_c_463_n 5.54777e-19 $X=4.3 $Y=1.515 $X2=0 $Y2=0
cc_213 N_A_M1009_g N_A_498_368#_c_452_n 2.17858e-19 $X=3.85 $Y=2.4 $X2=0 $Y2=0
cc_214 N_A_M1011_g N_A_498_368#_c_452_n 0.0110065f $X=4.3 $Y=2.4 $X2=0 $Y2=0
cc_215 N_A_M1002_g N_VGND_c_480_n 5.17057e-19 $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_216 N_A_M1004_g N_VGND_c_480_n 0.0130256f $X=4.285 $Y=0.74 $X2=0 $Y2=0
cc_217 A N_VGND_c_480_n 0.023824f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_218 N_A_c_248_n N_VGND_c_480_n 7.92882e-19 $X=4.3 $Y=1.515 $X2=0 $Y2=0
cc_219 N_A_M1002_g N_VGND_c_482_n 0.00383152f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_220 N_A_M1004_g N_VGND_c_482_n 0.00444681f $X=4.285 $Y=0.74 $X2=0 $Y2=0
cc_221 N_A_M1002_g N_VGND_c_487_n 0.0113336f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_222 N_A_M1004_g N_VGND_c_487_n 4.39287e-19 $X=4.285 $Y=0.74 $X2=0 $Y2=0
cc_223 N_A_M1002_g N_VGND_c_488_n 0.00753404f $X=3.805 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A_M1004_g N_VGND_c_488_n 0.00877997f $X=4.285 $Y=0.74 $X2=0 $Y2=0
cc_225 N_VPWR_c_293_n N_A_227_368#_c_348_n 0.0663622f $X=0.725 $Y=2.115 $X2=0
+ $Y2=0
cc_226 N_VPWR_c_298_n N_A_227_368#_c_349_n 0.0357927f $X=3.46 $Y=3.33 $X2=0
+ $Y2=0
cc_227 N_VPWR_c_292_n N_A_227_368#_c_349_n 0.0200586f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_228 N_VPWR_c_293_n N_A_227_368#_c_350_n 0.0125436f $X=0.725 $Y=2.115 $X2=0
+ $Y2=0
cc_229 N_VPWR_c_298_n N_A_227_368#_c_350_n 0.0235512f $X=3.46 $Y=3.33 $X2=0
+ $Y2=0
cc_230 N_VPWR_c_292_n N_A_227_368#_c_350_n 0.0126924f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_231 N_VPWR_c_294_n N_A_227_368#_c_352_n 0.0125436f $X=3.625 $Y=2.395 $X2=0
+ $Y2=0
cc_232 N_VPWR_c_298_n N_A_227_368#_c_352_n 0.0620536f $X=3.46 $Y=3.33 $X2=0
+ $Y2=0
cc_233 N_VPWR_c_292_n N_A_227_368#_c_352_n 0.0344172f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_234 N_VPWR_c_294_n N_A_227_368#_c_353_n 0.0420849f $X=3.625 $Y=2.395 $X2=0
+ $Y2=0
cc_235 N_VPWR_c_298_n N_A_227_368#_c_354_n 0.0199669f $X=3.46 $Y=3.33 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_292_n N_A_227_368#_c_354_n 0.0107485f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_237 N_VPWR_M1009_s N_A_498_368#_c_451_n 0.00549825f $X=3.485 $Y=1.84 $X2=0
+ $Y2=0
cc_238 N_VPWR_c_294_n N_A_498_368#_c_451_n 0.0219302f $X=3.625 $Y=2.395 $X2=0
+ $Y2=0
cc_239 N_VPWR_c_294_n N_A_498_368#_c_452_n 0.0234083f $X=3.625 $Y=2.395 $X2=0
+ $Y2=0
cc_240 N_VPWR_c_296_n N_A_498_368#_c_452_n 0.0295855f $X=4.525 $Y=2.115 $X2=0
+ $Y2=0
cc_241 N_VPWR_c_299_n N_A_498_368#_c_452_n 0.0109793f $X=4.425 $Y=3.33 $X2=0
+ $Y2=0
cc_242 N_VPWR_c_292_n N_A_498_368#_c_452_n 0.00901959f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_243 N_A_227_368#_c_349_n N_Y_M1005_d 0.00165831f $X=2.01 $Y=2.99 $X2=0 $Y2=0
cc_244 N_A_227_368#_c_348_n N_Y_c_393_n 0.0307826f $X=1.275 $Y=1.985 $X2=0 $Y2=0
cc_245 N_A_227_368#_c_349_n N_Y_c_393_n 0.0118736f $X=2.01 $Y=2.99 $X2=0 $Y2=0
cc_246 N_A_227_368#_c_351_n N_Y_c_393_n 0.0300333f $X=2.175 $Y=1.985 $X2=0 $Y2=0
cc_247 N_A_227_368#_c_352_n N_A_498_368#_M1007_d 0.00165831f $X=2.97 $Y=2.99
+ $X2=-0.19 $Y2=1.66
cc_248 N_A_227_368#_M1010_s N_A_498_368#_c_451_n 0.0050953f $X=2.94 $Y=1.84
+ $X2=0 $Y2=0
cc_249 N_A_227_368#_c_353_n N_A_498_368#_c_451_n 0.0197632f $X=3.075 $Y=2.455
+ $X2=0 $Y2=0
cc_250 N_A_227_368#_c_352_n N_A_498_368#_c_456_n 0.0159318f $X=2.97 $Y=2.99
+ $X2=0 $Y2=0
cc_251 N_Y_c_397_n N_VGND_M1012_d 0.0100206f $X=2.505 $Y=0.95 $X2=0 $Y2=0
cc_252 N_Y_c_399_n N_VGND_M1012_d 0.00237017f $X=1.81 $Y=0.95 $X2=0 $Y2=0
cc_253 N_Y_c_395_n N_VGND_M1013_s 0.0120678f $X=3.925 $Y=1.045 $X2=0 $Y2=0
cc_254 N_Y_c_392_n N_VGND_c_478_n 0.0160793f $X=1.285 $Y=0.515 $X2=0 $Y2=0
cc_255 N_Y_c_395_n N_VGND_c_480_n 0.00729485f $X=3.925 $Y=1.045 $X2=0 $Y2=0
cc_256 N_Y_c_396_n N_VGND_c_480_n 0.0236511f $X=4.02 $Y=0.515 $X2=0 $Y2=0
cc_257 N_Y_c_396_n N_VGND_c_482_n 0.0115122f $X=4.02 $Y=0.515 $X2=0 $Y2=0
cc_258 N_Y_c_392_n N_VGND_c_484_n 0.011986f $X=1.285 $Y=0.515 $X2=0 $Y2=0
cc_259 N_Y_c_392_n N_VGND_c_485_n 0.0112611f $X=1.285 $Y=0.515 $X2=0 $Y2=0
cc_260 N_Y_c_394_n N_VGND_c_485_n 0.011219f $X=2.6 $Y=0.515 $X2=0 $Y2=0
cc_261 N_Y_c_397_n N_VGND_c_485_n 0.0385023f $X=2.505 $Y=0.95 $X2=0 $Y2=0
cc_262 N_Y_c_399_n N_VGND_c_485_n 0.016076f $X=1.81 $Y=0.95 $X2=0 $Y2=0
cc_263 N_Y_c_394_n N_VGND_c_486_n 0.00838873f $X=2.6 $Y=0.515 $X2=0 $Y2=0
cc_264 N_Y_c_394_n N_VGND_c_487_n 0.0183801f $X=2.6 $Y=0.515 $X2=0 $Y2=0
cc_265 N_Y_c_395_n N_VGND_c_487_n 0.0575387f $X=3.925 $Y=1.045 $X2=0 $Y2=0
cc_266 N_Y_c_396_n N_VGND_c_487_n 0.0184157f $X=4.02 $Y=0.515 $X2=0 $Y2=0
cc_267 N_Y_c_392_n N_VGND_c_488_n 0.00991881f $X=1.285 $Y=0.515 $X2=0 $Y2=0
cc_268 N_Y_c_394_n N_VGND_c_488_n 0.00694347f $X=2.6 $Y=0.515 $X2=0 $Y2=0
cc_269 N_Y_c_396_n N_VGND_c_488_n 0.0095288f $X=4.02 $Y=0.515 $X2=0 $Y2=0
cc_270 N_Y_c_397_n N_VGND_c_488_n 0.00769121f $X=2.505 $Y=0.95 $X2=0 $Y2=0
cc_271 N_Y_c_399_n N_VGND_c_488_n 0.00627259f $X=1.81 $Y=0.95 $X2=0 $Y2=0

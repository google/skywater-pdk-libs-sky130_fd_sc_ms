* File: sky130_fd_sc_ms__xor3_2.spice
* Created: Wed Sep  2 12:34:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__xor3_2.pex.spice"
.subckt sky130_fd_sc_ms__xor3_2  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1018 N_VGND_M1018_d N_A_83_289#_M1018_g N_A_27_134#_M1018_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.34745 AS=0.1824 PD=1.81 PS=1.85 NRD=91.476 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1000 N_A_83_289#_M1000_d N_A_M1000_g N_VGND_M1018_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.169862 AS=0.34745 PD=1.275 PS=1.81 NRD=0 NRS=91.476 M=1 R=4.26667
+ SA=75001 SB=75002 A=0.096 P=1.58 MULT=1
MM1020 N_A_416_113#_M1020_d N_B_M1020_g N_A_83_289#_M1000_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.125283 AS=0.169862 PD=1.19547 PS=1.275 NRD=0 NRS=47.808 M=1
+ R=4.26667 SA=75001.5 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1010 N_A_27_134#_M1010_d N_A_440_315#_M1010_g N_A_416_113#_M1020_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.125326 AS=0.082217 PD=0.919245 PS=0.784528 NRD=19.992
+ NRS=20.712 M=1 R=2.8 SA=75002.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1017 N_A_375_419#_M1017_d N_B_M1017_g N_A_27_134#_M1010_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.1495 AS=0.190974 PD=1.14 PS=1.40075 NRD=15.468 NRS=31.872 M=1
+ R=4.26667 SA=75002 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1021 N_A_83_289#_M1021_d N_A_440_315#_M1021_g N_A_375_419#_M1017_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.2848 AS=0.1495 PD=2.17 PS=1.14 NRD=31.872 NRS=15.468 M=1
+ R=4.26667 SA=75002.6 SB=75000.4 A=0.096 P=1.58 MULT=1
MM1011 N_VGND_M1011_d N_B_M1011_g N_A_440_315#_M1011_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.46725 AS=0.2035 PD=2.88 PS=2.03 NRD=93.468 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.4 A=0.111 P=1.78 MULT=1
MM1005 N_A_1198_424#_M1005_d N_A_1162_379#_M1005_g N_A_375_419#_M1005_s VNB
+ NLOWVT L=0.15 W=0.64 AD=0.169775 AS=0.176 PD=1.24 PS=1.83 NRD=47.808 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1009 N_A_416_113#_M1009_d N_C_M1009_g N_A_1198_424#_M1005_d VNB NLOWVT L=0.15
+ W=0.64 AD=0.2144 AS=0.169775 PD=1.95 PS=1.24 NRD=4.68 NRS=0 M=1 R=4.26667
+ SA=75000.8 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1019 N_VGND_M1019_d N_C_M1019_g N_A_1162_379#_M1019_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.106521 AS=0.1197 PD=0.847241 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1019_d N_A_1198_424#_M1002_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.187679 AS=0.1036 PD=1.49276 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1014 N_VGND_M1014_d N_A_1198_424#_M1014_g N_X_M1002_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1006 N_VPWR_M1006_d N_A_83_289#_M1006_g N_A_27_134#_M1006_s VPB PSHORT L=0.18
+ W=1 AD=0.2075 AS=0.28 PD=1.415 PS=2.56 NRD=8.8453 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90002.4 A=0.18 P=2.36 MULT=1
MM1008 N_A_83_289#_M1008_d N_A_M1008_g N_VPWR_M1006_d VPB PSHORT L=0.18 W=1
+ AD=0.186413 AS=0.2075 PD=1.47283 PS=1.415 NRD=0 NRS=17.73 M=1 R=5.55556
+ SA=90000.8 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1023 N_A_375_419#_M1023_d N_B_M1023_g N_A_83_289#_M1008_d VPB PSHORT L=0.18
+ W=0.84 AD=0.146432 AS=0.156587 PD=1.32243 PS=1.23717 NRD=0 NRS=18.7544 M=1
+ R=4.66667 SA=90001.3 SB=90001.6 A=0.1512 P=2.04 MULT=1
MM1001 N_A_27_134#_M1001_d N_A_440_315#_M1001_g N_A_375_419#_M1023_d VPB PSHORT
+ L=0.18 W=0.64 AD=0.0864 AS=0.111568 PD=0.91 PS=1.00757 NRD=0 NRS=13.8491 M=1
+ R=3.55556 SA=90001.8 SB=90001.5 A=0.1152 P=1.64 MULT=1
MM1003 N_A_416_113#_M1003_d N_B_M1003_g N_A_27_134#_M1001_d VPB PSHORT L=0.18
+ W=0.64 AD=0.122465 AS=0.0864 PD=1.03351 PS=0.91 NRD=26.1616 NRS=0 M=1
+ R=3.55556 SA=90002.3 SB=90001.1 A=0.1152 P=1.64 MULT=1
MM1013 N_A_83_289#_M1013_d N_A_440_315#_M1013_g N_A_416_113#_M1003_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.5418 AS=0.160735 PD=2.97 PS=1.35649 NRD=71.511 NRS=0 M=1
+ R=4.66667 SA=90002.2 SB=90000.6 A=0.1512 P=2.04 MULT=1
MM1022 N_VPWR_M1022_d N_B_M1022_g N_A_440_315#_M1022_s VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.3136 PD=2.8 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1015 N_A_1198_424#_M1015_d N_A_1162_379#_M1015_g N_A_416_113#_M1015_s VPB
+ PSHORT L=0.18 W=0.84 AD=0.2436 AS=0.2352 PD=1.42 PS=2.24 NRD=71.511 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90000.9 A=0.1512 P=2.04 MULT=1
MM1012 N_A_375_419#_M1012_d N_C_M1012_g N_A_1198_424#_M1015_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.2436 PD=2.24 PS=1.42 NRD=0 NRS=0 M=1 R=4.66667
+ SA=90000.9 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1016 N_VPWR_M1016_d N_C_M1016_g N_A_1162_379#_M1016_s VPB PSHORT L=0.18 W=0.64
+ AD=0.278109 AS=0.2304 PD=1.33455 PS=2 NRD=25.3933 NRS=23.0687 M=1 R=3.55556
+ SA=90000.3 SB=90001.5 A=0.1152 P=1.64 MULT=1
MM1004 N_X_M1004_d N_A_1198_424#_M1004_g N_VPWR_M1016_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.486691 PD=1.39 PS=2.33545 NRD=0 NRS=62.4293 M=1 R=6.22222
+ SA=90000.9 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1007 N_X_M1004_d N_A_1198_424#_M1007_g N_VPWR_M1007_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.4
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX24_noxref VNB VPB NWDIODE A=18.5628 P=23.68
c_109 VNB 0 1.49322e-19 $X=0 $Y=0
c_194 VPB 0 2.47561e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__xor3_2.pxi.spice"
*
.ends
*
*

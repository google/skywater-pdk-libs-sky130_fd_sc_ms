* File: sky130_fd_sc_ms__a41oi_4.pex.spice
* Created: Wed Sep  2 11:56:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__A41OI_4%B1 3 5 7 8 10 13 15 17 18 20 22 23 24 25 39
+ 41
c75 41 0 1.97368e-19 $X=1.595 $Y=1.532
c76 20 0 1.19863e-19 $X=1.955 $Y=1.715
r77 40 41 34.8101 $w=3.65e-07 $l=9e-08 $layer=POLY_cond $X=1.505 $Y=1.532
+ $X2=1.595 $Y2=1.532
r78 38 40 37.9425 $w=3.65e-07 $l=2.4e-07 $layer=POLY_cond $X=1.265 $Y=1.532
+ $X2=1.505 $Y2=1.532
r79 38 39 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.265
+ $Y=1.515 $X2=1.265 $Y2=1.515
r80 36 38 41.1044 $w=3.65e-07 $l=2.6e-07 $layer=POLY_cond $X=1.005 $Y=1.532
+ $X2=1.265 $Y2=1.532
r81 33 34 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.585
+ $Y=1.515 $X2=0.585 $Y2=1.515
r82 31 33 11.857 $w=3.65e-07 $l=7.5e-08 $layer=POLY_cond $X=0.51 $Y=1.532
+ $X2=0.585 $Y2=1.532
r83 25 39 1.74206 $w=4.28e-07 $l=6.5e-08 $layer=LI1_cond $X=1.2 $Y=1.565
+ $X2=1.265 $Y2=1.565
r84 24 25 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=1.2 $Y2=1.565
r85 24 34 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=1.565
+ $X2=0.585 $Y2=1.565
r86 23 34 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.24 $Y=1.565
+ $X2=0.585 $Y2=1.565
r87 20 22 183.428 $w=1.8e-07 $l=6.85e-07 $layer=POLY_cond $X=1.955 $Y=1.715
+ $X2=1.955 $Y2=2.4
r88 18 20 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.865 $Y=1.64
+ $X2=1.955 $Y2=1.715
r89 18 41 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.865 $Y=1.64
+ $X2=1.595 $Y2=1.64
r90 15 40 19.2931 $w=1.8e-07 $l=1.83e-07 $layer=POLY_cond $X=1.505 $Y=1.715
+ $X2=1.505 $Y2=1.532
r91 15 17 183.428 $w=1.8e-07 $l=6.85e-07 $layer=POLY_cond $X=1.505 $Y=1.715
+ $X2=1.505 $Y2=2.4
r92 11 36 1.58094 $w=3.65e-07 $l=1e-08 $layer=POLY_cond $X=0.995 $Y=1.532
+ $X2=1.005 $Y2=1.532
r93 11 33 64.8184 $w=3.65e-07 $l=4.1e-07 $layer=POLY_cond $X=0.995 $Y=1.532
+ $X2=0.585 $Y2=1.532
r94 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.995 $Y=1.35
+ $X2=0.995 $Y2=0.74
r95 8 36 19.2931 $w=1.8e-07 $l=1.83e-07 $layer=POLY_cond $X=1.005 $Y=1.715
+ $X2=1.005 $Y2=1.532
r96 8 10 183.428 $w=1.8e-07 $l=6.85e-07 $layer=POLY_cond $X=1.005 $Y=1.715
+ $X2=1.005 $Y2=2.4
r97 5 31 19.2931 $w=1.8e-07 $l=1.83e-07 $layer=POLY_cond $X=0.51 $Y=1.715
+ $X2=0.51 $Y2=1.532
r98 5 7 183.428 $w=1.8e-07 $l=6.85e-07 $layer=POLY_cond $X=0.51 $Y=1.715
+ $X2=0.51 $Y2=2.4
r99 1 31 2.37141 $w=3.65e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.532
+ $X2=0.51 $Y2=1.532
r100 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A41OI_4%A1 1 3 4 5 6 8 9 11 12 14 15 17 18 20 21 23
+ 24 26 27 28 39 42
c108 39 0 1.19863e-19 $X=3.13 $Y=1.515
c109 18 0 1.56189e-19 $X=3.405 $Y=1.745
c110 5 0 3.74685e-19 $X=2.06 $Y=1.28
r111 41 42 27.8268 $w=4.85e-07 $l=2.8e-07 $layer=POLY_cond $X=3.405 $Y=1.475
+ $X2=3.685 $Y2=1.475
r112 40 41 14.9072 $w=4.85e-07 $l=1.5e-07 $layer=POLY_cond $X=3.255 $Y=1.475
+ $X2=3.405 $Y2=1.475
r113 38 40 12.4227 $w=4.85e-07 $l=1.25e-07 $layer=POLY_cond $X=3.13 $Y=1.475
+ $X2=3.255 $Y2=1.475
r114 38 39 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.13
+ $Y=1.515 $X2=3.13 $Y2=1.515
r115 36 38 17.3918 $w=4.85e-07 $l=1.75e-07 $layer=POLY_cond $X=2.955 $Y=1.475
+ $X2=3.13 $Y2=1.475
r116 35 36 46.7093 $w=4.85e-07 $l=4.7e-07 $layer=POLY_cond $X=2.485 $Y=1.475
+ $X2=2.955 $Y2=1.475
r117 33 35 3.47835 $w=4.85e-07 $l=3.5e-08 $layer=POLY_cond $X=2.45 $Y=1.475
+ $X2=2.485 $Y2=1.475
r118 33 34 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.45
+ $Y=1.515 $X2=2.45 $Y2=1.515
r119 31 33 4.47217 $w=4.85e-07 $l=4.5e-08 $layer=POLY_cond $X=2.405 $Y=1.475
+ $X2=2.45 $Y2=1.475
r120 28 39 0.26801 $w=4.28e-07 $l=1e-08 $layer=LI1_cond $X=3.12 $Y=1.565
+ $X2=3.13 $Y2=1.565
r121 27 28 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=3.12 $Y2=1.565
r122 27 34 5.09219 $w=4.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.64 $Y=1.565
+ $X2=2.45 $Y2=1.565
r123 24 42 22.3608 $w=4.85e-07 $l=3.65582e-07 $layer=POLY_cond $X=3.91 $Y=1.745
+ $X2=3.685 $Y2=1.475
r124 24 26 175.394 $w=1.8e-07 $l=6.55e-07 $layer=POLY_cond $X=3.91 $Y=1.745
+ $X2=3.91 $Y2=2.4
r125 21 42 30.6402 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.685 $Y=1.205
+ $X2=3.685 $Y2=1.475
r126 21 23 149.42 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.685 $Y=1.205
+ $X2=3.685 $Y2=0.74
r127 18 41 26.1155 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=3.405 $Y=1.745
+ $X2=3.405 $Y2=1.475
r128 18 20 175.394 $w=1.8e-07 $l=6.55e-07 $layer=POLY_cond $X=3.405 $Y=1.745
+ $X2=3.405 $Y2=2.4
r129 15 40 30.6402 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.255 $Y=1.205
+ $X2=3.255 $Y2=1.475
r130 15 17 149.42 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.255 $Y=1.205
+ $X2=3.255 $Y2=0.74
r131 12 36 26.1155 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=2.955 $Y=1.745
+ $X2=2.955 $Y2=1.475
r132 12 14 175.394 $w=1.8e-07 $l=6.55e-07 $layer=POLY_cond $X=2.955 $Y=1.745
+ $X2=2.955 $Y2=2.4
r133 9 35 30.6402 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.485 $Y=1.205
+ $X2=2.485 $Y2=1.475
r134 9 11 149.42 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.485 $Y=1.205
+ $X2=2.485 $Y2=0.74
r135 6 31 26.1155 $w=1.8e-07 $l=2.7e-07 $layer=POLY_cond $X=2.405 $Y=1.745
+ $X2=2.405 $Y2=1.475
r136 6 8 175.394 $w=1.8e-07 $l=6.55e-07 $layer=POLY_cond $X=2.405 $Y=1.745
+ $X2=2.405 $Y2=2.4
r137 4 31 37.0697 $w=4.85e-07 $l=2.47841e-07 $layer=POLY_cond $X=2.285 $Y=1.28
+ $X2=2.405 $Y2=1.475
r138 4 5 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.285 $Y=1.28
+ $X2=2.06 $Y2=1.28
r139 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.985 $Y=1.205
+ $X2=2.06 $Y2=1.28
r140 1 3 149.42 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.985 $Y=1.205
+ $X2=1.985 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A41OI_4%A2 1 3 6 8 10 13 15 17 20 22 24 27 31 34 35
+ 48 50 57
c95 57 0 1.1015e-19 $X=4.675 $Y=1.55
c96 50 0 1.61301e-19 $X=4.445 $Y=1.55
c97 48 0 2.34008e-19 $X=5.545 $Y=1.427
c98 6 0 6.08204e-20 $X=4.36 $Y=2.4
c99 1 0 1.63532e-19 $X=4.185 $Y=1.205
r100 45 46 26.6334 $w=3.71e-07 $l=2.05e-07 $layer=POLY_cond $X=5.115 $Y=1.427
+ $X2=5.32 $Y2=1.427
r101 44 45 31.8302 $w=3.71e-07 $l=2.45e-07 $layer=POLY_cond $X=4.87 $Y=1.427
+ $X2=5.115 $Y2=1.427
r102 43 44 24.035 $w=3.71e-07 $l=1.85e-07 $layer=POLY_cond $X=4.685 $Y=1.427
+ $X2=4.87 $Y2=1.427
r103 42 50 0.260017 $w=4.58e-07 $l=1e-08 $layer=LI1_cond $X=4.435 $Y=1.55
+ $X2=4.445 $Y2=1.55
r104 41 43 32.4798 $w=3.71e-07 $l=2.5e-07 $layer=POLY_cond $X=4.435 $Y=1.427
+ $X2=4.685 $Y2=1.427
r105 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.435
+ $Y=1.485 $X2=4.435 $Y2=1.485
r106 39 41 9.74394 $w=3.71e-07 $l=7.5e-08 $layer=POLY_cond $X=4.36 $Y=1.427
+ $X2=4.435 $Y2=1.427
r107 35 57 3.96409 $w=4.58e-07 $l=1.15e-07 $layer=LI1_cond $X=4.56 $Y=1.55
+ $X2=4.675 $Y2=1.55
r108 35 50 2.9902 $w=4.58e-07 $l=1.15e-07 $layer=LI1_cond $X=4.56 $Y=1.55
+ $X2=4.445 $Y2=1.55
r109 34 42 9.23061 $w=4.58e-07 $l=3.55e-07 $layer=LI1_cond $X=4.08 $Y=1.55
+ $X2=4.435 $Y2=1.55
r110 32 48 11.6927 $w=3.71e-07 $l=9e-08 $layer=POLY_cond $X=5.455 $Y=1.427
+ $X2=5.545 $Y2=1.427
r111 32 46 17.5391 $w=3.71e-07 $l=1.35e-07 $layer=POLY_cond $X=5.455 $Y=1.427
+ $X2=5.32 $Y2=1.427
r112 31 57 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=5.455 $Y=1.485
+ $X2=4.675 $Y2=1.485
r113 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.455
+ $Y=1.485 $X2=5.455 $Y2=1.485
r114 25 48 35.7278 $w=3.71e-07 $l=3.70068e-07 $layer=POLY_cond $X=5.82 $Y=1.65
+ $X2=5.545 $Y2=1.427
r115 25 27 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=5.82 $Y=1.65
+ $X2=5.82 $Y2=2.4
r116 22 48 24.032 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.545 $Y=1.205
+ $X2=5.545 $Y2=1.427
r117 22 24 149.42 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.545 $Y=1.205
+ $X2=5.545 $Y2=0.74
r118 18 46 19.6776 $w=1.8e-07 $l=2.23e-07 $layer=POLY_cond $X=5.32 $Y=1.65
+ $X2=5.32 $Y2=1.427
r119 18 20 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=5.32 $Y=1.65
+ $X2=5.32 $Y2=2.4
r120 15 45 24.032 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=5.115 $Y=1.205
+ $X2=5.115 $Y2=1.427
r121 15 17 149.42 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.115 $Y=1.205
+ $X2=5.115 $Y2=0.74
r122 11 44 19.6776 $w=1.8e-07 $l=2.23e-07 $layer=POLY_cond $X=4.87 $Y=1.65
+ $X2=4.87 $Y2=1.427
r123 11 13 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=4.87 $Y=1.65
+ $X2=4.87 $Y2=2.4
r124 8 43 24.032 $w=1.5e-07 $l=2.22e-07 $layer=POLY_cond $X=4.685 $Y=1.205
+ $X2=4.685 $Y2=1.427
r125 8 10 149.42 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.685 $Y=1.205
+ $X2=4.685 $Y2=0.74
r126 4 39 19.6776 $w=1.8e-07 $l=2.23e-07 $layer=POLY_cond $X=4.36 $Y=1.65
+ $X2=4.36 $Y2=1.427
r127 4 6 291.532 $w=1.8e-07 $l=7.5e-07 $layer=POLY_cond $X=4.36 $Y=1.65 $X2=4.36
+ $Y2=2.4
r128 1 39 22.7358 $w=3.71e-07 $l=2.96874e-07 $layer=POLY_cond $X=4.185 $Y=1.205
+ $X2=4.36 $Y2=1.427
r129 1 3 149.42 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.185 $Y=1.205
+ $X2=4.185 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__A41OI_4%A3 3 7 11 15 19 23 27 31 33 34 35 36 37 57
c88 27 0 7.4136e-20 $X=7.72 $Y=2.4
c89 15 0 1.85629e-19 $X=6.965 $Y=0.74
r90 56 57 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=7.72 $Y=1.515
+ $X2=7.825 $Y2=1.515
r91 54 56 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.705 $Y=1.515
+ $X2=7.72 $Y2=1.515
r92 54 55 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=7.705
+ $Y=1.515 $X2=7.705 $Y2=1.515
r93 52 54 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=7.395 $Y=1.515
+ $X2=7.705 $Y2=1.515
r94 51 52 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=7.22 $Y=1.515
+ $X2=7.395 $Y2=1.515
r95 50 51 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=6.965 $Y=1.515
+ $X2=7.22 $Y2=1.515
r96 49 50 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=6.77 $Y=1.515
+ $X2=6.965 $Y2=1.515
r97 48 49 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=6.535 $Y=1.515
+ $X2=6.77 $Y2=1.515
r98 46 48 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=6.345 $Y=1.515
+ $X2=6.535 $Y2=1.515
r99 46 47 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=6.345
+ $Y=1.515 $X2=6.345 $Y2=1.515
r100 43 46 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.27 $Y=1.515
+ $X2=6.345 $Y2=1.515
r101 37 55 5.76222 $w=4.28e-07 $l=2.15e-07 $layer=LI1_cond $X=7.92 $Y=1.565
+ $X2=7.705 $Y2=1.565
r102 36 55 7.10226 $w=4.28e-07 $l=2.65e-07 $layer=LI1_cond $X=7.44 $Y=1.565
+ $X2=7.705 $Y2=1.565
r103 35 36 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.565
+ $X2=7.44 $Y2=1.565
r104 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.96 $Y2=1.565
r105 34 47 3.61813 $w=4.28e-07 $l=1.35e-07 $layer=LI1_cond $X=6.48 $Y=1.565
+ $X2=6.345 $Y2=1.565
r106 33 47 9.24634 $w=4.28e-07 $l=3.45e-07 $layer=LI1_cond $X=6 $Y=1.565
+ $X2=6.345 $Y2=1.565
r107 29 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.825 $Y=1.35
+ $X2=7.825 $Y2=1.515
r108 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.825 $Y=1.35
+ $X2=7.825 $Y2=0.74
r109 25 56 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.72 $Y=1.68
+ $X2=7.72 $Y2=1.515
r110 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.72 $Y=1.68
+ $X2=7.72 $Y2=2.4
r111 21 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.395 $Y=1.35
+ $X2=7.395 $Y2=1.515
r112 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.395 $Y=1.35
+ $X2=7.395 $Y2=0.74
r113 17 51 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.22 $Y=1.68
+ $X2=7.22 $Y2=1.515
r114 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=7.22 $Y=1.68
+ $X2=7.22 $Y2=2.4
r115 13 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.965 $Y=1.35
+ $X2=6.965 $Y2=1.515
r116 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.965 $Y=1.35
+ $X2=6.965 $Y2=0.74
r117 9 49 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.77 $Y=1.68
+ $X2=6.77 $Y2=1.515
r118 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.77 $Y=1.68
+ $X2=6.77 $Y2=2.4
r119 5 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.535 $Y=1.35
+ $X2=6.535 $Y2=1.515
r120 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.535 $Y=1.35
+ $X2=6.535 $Y2=0.74
r121 1 43 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.27 $Y=1.68
+ $X2=6.27 $Y2=1.515
r122 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.27 $Y=1.68 $X2=6.27
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A41OI_4%A4 3 7 11 15 19 23 27 31 33 34 35 36 55
c77 36 0 7.4136e-20 $X=9.84 $Y=1.665
c78 7 0 2.04552e-19 $X=8.255 $Y=0.74
c79 3 0 1.72297e-19 $X=8.22 $Y=2.4
r80 54 55 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=9.57 $Y=1.515
+ $X2=9.585 $Y2=1.515
r81 52 54 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=9.47 $Y=1.515 $X2=9.57
+ $Y2=1.515
r82 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.47
+ $Y=1.515 $X2=9.47 $Y2=1.515
r83 50 52 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=9.12 $Y=1.515
+ $X2=9.47 $Y2=1.515
r84 49 50 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=9.115 $Y=1.515
+ $X2=9.12 $Y2=1.515
r85 48 49 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=8.685 $Y=1.515
+ $X2=9.115 $Y2=1.515
r86 47 48 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=8.67 $Y=1.515
+ $X2=8.685 $Y2=1.515
r87 45 47 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=8.45 $Y=1.515
+ $X2=8.67 $Y2=1.515
r88 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.45
+ $Y=1.515 $X2=8.45 $Y2=1.515
r89 43 45 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=8.255 $Y=1.515
+ $X2=8.45 $Y2=1.515
r90 41 43 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=8.22 $Y=1.515
+ $X2=8.255 $Y2=1.515
r91 36 53 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=9.84 $Y=1.565
+ $X2=9.47 $Y2=1.565
r92 35 53 2.94811 $w=4.28e-07 $l=1.1e-07 $layer=LI1_cond $X=9.36 $Y=1.565
+ $X2=9.47 $Y2=1.565
r93 34 35 12.8645 $w=4.28e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.565
+ $X2=9.36 $Y2=1.565
r94 34 46 11.5244 $w=4.28e-07 $l=4.3e-07 $layer=LI1_cond $X=8.88 $Y=1.565
+ $X2=8.45 $Y2=1.565
r95 33 46 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=8.4 $Y=1.565 $X2=8.45
+ $Y2=1.565
r96 29 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.585 $Y=1.35
+ $X2=9.585 $Y2=1.515
r97 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.585 $Y=1.35
+ $X2=9.585 $Y2=0.74
r98 25 54 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.57 $Y=1.68
+ $X2=9.57 $Y2=1.515
r99 25 27 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=9.57 $Y=1.68
+ $X2=9.57 $Y2=2.4
r100 21 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.115 $Y=1.35
+ $X2=9.115 $Y2=1.515
r101 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.115 $Y=1.35
+ $X2=9.115 $Y2=0.74
r102 17 50 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.12 $Y=1.68
+ $X2=9.12 $Y2=1.515
r103 17 19 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=9.12 $Y=1.68
+ $X2=9.12 $Y2=2.4
r104 13 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.685 $Y=1.35
+ $X2=8.685 $Y2=1.515
r105 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.685 $Y=1.35
+ $X2=8.685 $Y2=0.74
r106 9 47 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.67 $Y=1.68
+ $X2=8.67 $Y2=1.515
r107 9 11 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.67 $Y=1.68
+ $X2=8.67 $Y2=2.4
r108 5 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.255 $Y=1.35
+ $X2=8.255 $Y2=1.515
r109 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.255 $Y=1.35
+ $X2=8.255 $Y2=0.74
r110 1 41 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.22 $Y=1.68
+ $X2=8.22 $Y2=1.515
r111 1 3 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=8.22 $Y=1.68 $X2=8.22
+ $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__A41OI_4%A_27_368# 1 2 3 4 5 6 7 8 9 10 11 36 40 41
+ 44 46 48 49 50 54 56 57 60 62 66 68 72 74 78 80 84 86 90 92 94 96 98 102 105
+ 107 109 111 113 115
c192 84 0 1.72297e-19 $X=7.945 $Y=2.425
c193 56 0 1.30665e-19 $X=4.135 $Y=2.12
c194 54 0 1.35778e-19 $X=3.97 $Y=2.375
r195 94 117 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.795 $Y=2.12
+ $X2=9.795 $Y2=2.035
r196 94 96 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=9.795 $Y=2.12
+ $X2=9.795 $Y2=2.815
r197 93 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.06 $Y=2.035
+ $X2=8.895 $Y2=2.035
r198 92 117 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.63 $Y=2.035
+ $X2=9.795 $Y2=2.035
r199 92 93 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=9.63 $Y=2.035
+ $X2=9.06 $Y2=2.035
r200 88 115 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.895 $Y=2.12
+ $X2=8.895 $Y2=2.035
r201 88 90 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=8.895 $Y=2.12
+ $X2=8.895 $Y2=2.815
r202 87 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.11 $Y=2.035
+ $X2=7.945 $Y2=2.035
r203 86 115 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.73 $Y=2.035
+ $X2=8.895 $Y2=2.035
r204 86 87 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=8.73 $Y=2.035
+ $X2=8.11 $Y2=2.035
r205 82 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.945 $Y=2.12
+ $X2=7.945 $Y2=2.035
r206 82 84 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=7.945 $Y=2.12
+ $X2=7.945 $Y2=2.425
r207 81 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.16 $Y=2.035
+ $X2=6.995 $Y2=2.035
r208 80 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.78 $Y=2.035
+ $X2=7.945 $Y2=2.035
r209 80 81 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=7.78 $Y=2.035
+ $X2=7.16 $Y2=2.035
r210 76 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.995 $Y=2.12
+ $X2=6.995 $Y2=2.035
r211 76 78 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=6.995 $Y=2.12
+ $X2=6.995 $Y2=2.815
r212 75 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.21 $Y=2.035
+ $X2=6.045 $Y2=2.035
r213 74 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.83 $Y=2.035
+ $X2=6.995 $Y2=2.035
r214 74 75 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=6.83 $Y=2.035
+ $X2=6.21 $Y2=2.035
r215 70 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.045 $Y=2.12
+ $X2=6.045 $Y2=2.035
r216 70 72 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=6.045 $Y=2.12
+ $X2=6.045 $Y2=2.815
r217 69 107 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=5.26 $Y=2.035
+ $X2=5.095 $Y2=1.97
r218 68 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.88 $Y=2.035
+ $X2=6.045 $Y2=2.035
r219 68 69 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=5.88 $Y=2.035
+ $X2=5.26 $Y2=2.035
r220 64 107 0.89609 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=5.095 $Y=2.12
+ $X2=5.095 $Y2=1.97
r221 64 66 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=5.095 $Y=2.12
+ $X2=5.095 $Y2=2.815
r222 63 104 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.3 $Y=2.035
+ $X2=4.135 $Y2=2.035
r223 62 107 8.61065 $w=1.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=4.93 $Y=2.035
+ $X2=5.095 $Y2=1.97
r224 62 63 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=4.93 $Y=2.035
+ $X2=4.3 $Y2=2.035
r225 58 105 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.135 $Y=2.46
+ $X2=4.135 $Y2=2.375
r226 58 60 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=4.135 $Y=2.46
+ $X2=4.135 $Y2=2.815
r227 57 105 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.135 $Y=2.29
+ $X2=4.135 $Y2=2.375
r228 56 104 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.135 $Y=2.12
+ $X2=4.135 $Y2=2.035
r229 56 57 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=4.135 $Y=2.12
+ $X2=4.135 $Y2=2.29
r230 55 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.345 $Y=2.375
+ $X2=3.18 $Y2=2.375
r231 54 105 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.97 $Y=2.375
+ $X2=4.135 $Y2=2.375
r232 54 55 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=3.97 $Y=2.375
+ $X2=3.345 $Y2=2.375
r233 51 100 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=2.375
+ $X2=2.18 $Y2=2.375
r234 50 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.015 $Y=2.375
+ $X2=3.18 $Y2=2.375
r235 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.015 $Y=2.375
+ $X2=2.345 $Y2=2.375
r236 48 100 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=2.46
+ $X2=2.18 $Y2=2.375
r237 48 49 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=2.18 $Y=2.46
+ $X2=2.18 $Y2=2.905
r238 47 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.445 $Y=2.99
+ $X2=1.28 $Y2=2.99
r239 46 49 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.015 $Y=2.99
+ $X2=2.18 $Y2=2.905
r240 46 47 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.015 $Y=2.99
+ $X2=1.445 $Y2=2.99
r241 42 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=2.905
+ $X2=1.28 $Y2=2.99
r242 42 44 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=1.28 $Y=2.905
+ $X2=1.28 $Y2=2.405
r243 40 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=2.99
+ $X2=1.28 $Y2=2.99
r244 40 41 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=2.99
+ $X2=0.445 $Y2=2.99
r245 36 39 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=0.28 $Y=2.035
+ $X2=0.28 $Y2=2.815
r246 34 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.445 $Y2=2.99
r247 34 39 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.28 $Y2=2.815
r248 11 117 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=9.66
+ $Y=1.84 $X2=9.795 $Y2=2.035
r249 11 96 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.66
+ $Y=1.84 $X2=9.795 $Y2=2.815
r250 10 115 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=8.76
+ $Y=1.84 $X2=8.895 $Y2=2.035
r251 10 90 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.76
+ $Y=1.84 $X2=8.895 $Y2=2.815
r252 9 113 600 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=7.81
+ $Y=1.84 $X2=7.945 $Y2=2.035
r253 9 84 300 $w=1.7e-07 $l=6.48999e-07 $layer=licon1_PDIFF $count=2 $X=7.81
+ $Y=1.84 $X2=7.945 $Y2=2.425
r254 8 111 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=6.86
+ $Y=1.84 $X2=6.995 $Y2=2.035
r255 8 78 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=6.86
+ $Y=1.84 $X2=6.995 $Y2=2.815
r256 7 109 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=5.91
+ $Y=1.84 $X2=6.045 $Y2=2.035
r257 7 72 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.91
+ $Y=1.84 $X2=6.045 $Y2=2.815
r258 6 107 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.96
+ $Y=1.84 $X2=5.095 $Y2=1.985
r259 6 66 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.96
+ $Y=1.84 $X2=5.095 $Y2=2.815
r260 5 104 400 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_PDIFF $count=1 $X=4
+ $Y=1.84 $X2=4.135 $Y2=2.035
r261 5 60 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4
+ $Y=1.84 $X2=4.135 $Y2=2.815
r262 4 102 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=3.045
+ $Y=1.84 $X2=3.18 $Y2=2.375
r263 3 100 300 $w=1.7e-07 $l=5.98707e-07 $layer=licon1_PDIFF $count=2 $X=2.045
+ $Y=1.84 $X2=2.18 $Y2=2.375
r264 2 44 300 $w=1.7e-07 $l=6.50961e-07 $layer=licon1_PDIFF $count=2 $X=1.095
+ $Y=1.84 $X2=1.28 $Y2=2.405
r265 1 39 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r266 1 36 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.035
.ends

.subckt PM_SKY130_FD_SC_MS__A41OI_4%Y 1 2 3 4 5 18 22 23 28 31 32 34 36 41 44 46
+ 51 55 61 63
c104 61 0 1.73187e-19 $X=3.59 $Y=1.55
c105 55 0 1.21641e-19 $X=3.515 $Y=1.58
c106 51 0 1.63532e-19 $X=3.47 $Y=0.785
c107 46 0 1.77318e-19 $X=2.105 $Y=1.97
r108 58 63 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=3.59 $Y=1.675
+ $X2=3.59 $Y2=1.665
r109 55 63 1.75171 $w=2.48e-07 $l=3.8e-08 $layer=LI1_cond $X=3.59 $Y=1.627
+ $X2=3.59 $Y2=1.665
r110 55 61 4.73668 $w=2.48e-07 $l=7.7e-08 $layer=LI1_cond $X=3.59 $Y=1.627
+ $X2=3.59 $Y2=1.55
r111 55 58 1.70562 $w=2.48e-07 $l=3.7e-08 $layer=LI1_cond $X=3.59 $Y=1.712
+ $X2=3.59 $Y2=1.675
r112 54 55 10.9713 $w=2.48e-07 $l=2.38e-07 $layer=LI1_cond $X=3.59 $Y=1.95
+ $X2=3.59 $Y2=1.712
r113 53 61 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.55 $Y=1 $X2=3.55
+ $Y2=1.55
r114 51 53 10.2083 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=3.47 $Y=0.785
+ $X2=3.47 $Y2=1
r115 45 46 7.71634 $w=2.98e-07 $l=1.45e-07 $layer=LI1_cond $X=1.96 $Y=1.97
+ $X2=2.105 $Y2=1.97
r116 43 45 8.8354 $w=2.98e-07 $l=2.3e-07 $layer=LI1_cond $X=1.73 $Y=1.97
+ $X2=1.96 $Y2=1.97
r117 43 44 5.41145 $w=2.98e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=1.97
+ $X2=1.645 $Y2=1.97
r118 36 54 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.465 $Y=2.035
+ $X2=3.59 $Y2=1.95
r119 36 46 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.465 $Y=2.035
+ $X2=2.105 $Y2=2.035
r120 32 34 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.27 $Y=1.01
+ $X2=2.27 $Y2=0.76
r121 31 45 0.922372 $w=2.9e-07 $l=1.5e-07 $layer=LI1_cond $X=1.96 $Y=1.82
+ $X2=1.96 $Y2=1.97
r122 30 32 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.96 $Y=1.095
+ $X2=2.27 $Y2=1.095
r123 30 31 25.4332 $w=2.88e-07 $l=6.4e-07 $layer=LI1_cond $X=1.96 $Y=1.18
+ $X2=1.96 $Y2=1.82
r124 26 43 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.73 $Y=2.12 $X2=1.73
+ $Y2=1.97
r125 26 28 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=1.73 $Y=2.12
+ $X2=1.73 $Y2=2.57
r126 25 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=2.035
+ $X2=0.78 $Y2=2.035
r127 25 44 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=0.945 $Y=2.035
+ $X2=1.645 $Y2=2.035
r128 22 30 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.815 $Y=1.095
+ $X2=1.96 $Y2=1.095
r129 22 23 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.815 $Y=1.095
+ $X2=0.875 $Y2=1.095
r130 16 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.71 $Y=1.01
+ $X2=0.875 $Y2=1.095
r131 16 18 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.71 $Y=1.01
+ $X2=0.71 $Y2=0.515
r132 5 43 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.84 $X2=1.73 $Y2=1.985
r133 5 28 600 $w=1.7e-07 $l=7.94638e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.84 $X2=1.73 $Y2=2.57
r134 4 41 300 $w=1.7e-07 $l=3.1229e-07 $layer=licon1_PDIFF $count=2 $X=0.6
+ $Y=1.84 $X2=0.78 $Y2=2.075
r135 3 51 182 $w=1.7e-07 $l=4.79922e-07 $layer=licon1_NDIFF $count=1 $X=3.33
+ $Y=0.37 $X2=3.47 $Y2=0.785
r136 2 34 182 $w=1.7e-07 $l=4.83735e-07 $layer=licon1_NDIFF $count=1 $X=2.06
+ $Y=0.37 $X2=2.27 $Y2=0.76
r137 1 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A41OI_4%VPWR 1 2 3 4 5 6 7 8 27 29 33 35 39 41 45 47
+ 51 53 57 61 65 68 69 70 72 80 90 91 94 97 100 103 106 109 112
r143 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r144 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r145 107 110 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r146 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r147 104 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r148 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r149 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r150 98 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r151 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r152 95 98 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r153 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r154 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r155 88 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.84 $Y2=3.33
r156 88 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r157 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r158 85 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.53 $Y=3.33
+ $X2=8.405 $Y2=3.33
r159 85 87 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=8.53 $Y=3.33
+ $X2=8.88 $Y2=3.33
r160 84 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r161 84 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r162 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r163 81 109 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.61 $Y=3.33
+ $X2=7.485 $Y2=3.33
r164 81 83 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=7.61 $Y=3.33
+ $X2=7.92 $Y2=3.33
r165 80 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.28 $Y=3.33
+ $X2=8.405 $Y2=3.33
r166 80 83 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.28 $Y=3.33
+ $X2=7.92 $Y2=3.33
r167 79 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r168 78 79 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r169 75 79 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r170 74 78 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r171 74 75 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r172 72 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.515 $Y=3.33
+ $X2=2.68 $Y2=3.33
r173 72 78 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.515 $Y=3.33
+ $X2=2.16 $Y2=3.33
r174 70 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r175 70 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r176 68 87 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.26 $Y=3.33
+ $X2=8.88 $Y2=3.33
r177 68 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.26 $Y=3.33
+ $X2=9.345 $Y2=3.33
r178 67 90 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=9.43 $Y=3.33
+ $X2=9.84 $Y2=3.33
r179 67 69 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.43 $Y=3.33
+ $X2=9.345 $Y2=3.33
r180 63 69 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.345 $Y=3.245
+ $X2=9.345 $Y2=3.33
r181 63 65 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=9.345 $Y=3.245
+ $X2=9.345 $Y2=2.455
r182 59 112 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.405 $Y=3.245
+ $X2=8.405 $Y2=3.33
r183 59 61 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=8.405 $Y=3.245
+ $X2=8.405 $Y2=2.455
r184 55 109 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.485 $Y=3.245
+ $X2=7.485 $Y2=3.33
r185 55 57 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=7.485 $Y=3.245
+ $X2=7.485 $Y2=2.455
r186 54 106 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.66 $Y=3.33
+ $X2=6.535 $Y2=3.33
r187 53 109 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.36 $Y=3.33
+ $X2=7.485 $Y2=3.33
r188 53 54 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=7.36 $Y=3.33 $X2=6.66
+ $Y2=3.33
r189 49 106 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.535 $Y=3.245
+ $X2=6.535 $Y2=3.33
r190 49 51 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=6.535 $Y=3.245
+ $X2=6.535 $Y2=2.455
r191 48 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.71 $Y=3.33
+ $X2=5.585 $Y2=3.33
r192 47 106 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.41 $Y=3.33
+ $X2=6.535 $Y2=3.33
r193 47 48 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=6.41 $Y=3.33 $X2=5.71
+ $Y2=3.33
r194 43 103 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.585 $Y=3.245
+ $X2=5.585 $Y2=3.33
r195 43 45 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=5.585 $Y=3.245
+ $X2=5.585 $Y2=2.455
r196 42 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.75 $Y=3.33
+ $X2=4.625 $Y2=3.33
r197 41 103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.46 $Y=3.33
+ $X2=5.585 $Y2=3.33
r198 41 42 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=5.46 $Y=3.33
+ $X2=4.75 $Y2=3.33
r199 37 100 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=3.245
+ $X2=4.625 $Y2=3.33
r200 37 39 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=4.625 $Y=3.245
+ $X2=4.625 $Y2=2.455
r201 36 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.795 $Y=3.33
+ $X2=3.67 $Y2=3.33
r202 35 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.5 $Y=3.33
+ $X2=4.625 $Y2=3.33
r203 35 36 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=4.5 $Y=3.33
+ $X2=3.795 $Y2=3.33
r204 31 97 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=3.245
+ $X2=3.67 $Y2=3.33
r205 31 33 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=3.67 $Y=3.245
+ $X2=3.67 $Y2=2.795
r206 30 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.845 $Y=3.33
+ $X2=2.68 $Y2=3.33
r207 29 97 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.545 $Y=3.33
+ $X2=3.67 $Y2=3.33
r208 29 30 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.545 $Y=3.33
+ $X2=2.845 $Y2=3.33
r209 25 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=3.245
+ $X2=2.68 $Y2=3.33
r210 25 27 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=2.68 $Y=3.245
+ $X2=2.68 $Y2=2.735
r211 8 65 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=9.21
+ $Y=1.84 $X2=9.345 $Y2=2.455
r212 7 61 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=8.31
+ $Y=1.84 $X2=8.445 $Y2=2.455
r213 6 57 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=7.31
+ $Y=1.84 $X2=7.445 $Y2=2.455
r214 5 51 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=6.36
+ $Y=1.84 $X2=6.495 $Y2=2.455
r215 4 45 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=5.41
+ $Y=1.84 $X2=5.545 $Y2=2.455
r216 3 39 300 $w=1.7e-07 $l=6.79154e-07 $layer=licon1_PDIFF $count=2 $X=4.45
+ $Y=1.84 $X2=4.585 $Y2=2.455
r217 2 33 600 $w=1.7e-07 $l=1.02027e-06 $layer=licon1_PDIFF $count=1 $X=3.495
+ $Y=1.84 $X2=3.63 $Y2=2.795
r218 1 27 600 $w=1.7e-07 $l=9.83158e-07 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=1.84 $X2=2.68 $Y2=2.735
.ends

.subckt PM_SKY130_FD_SC_MS__A41OI_4%VGND 1 2 3 4 13 15 19 23 27 29 31 36 44 51
+ 52 58 61 64
r99 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r100 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r101 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r102 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r103 52 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=9.36
+ $Y2=0
r104 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r105 49 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.495 $Y=0 $X2=9.33
+ $Y2=0
r106 49 51 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.495 $Y=0 $X2=9.84
+ $Y2=0
r107 48 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r108 48 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r109 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r110 45 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.635 $Y=0 $X2=8.47
+ $Y2=0
r111 45 47 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=8.635 $Y=0 $X2=8.88
+ $Y2=0
r112 44 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.165 $Y=0 $X2=9.33
+ $Y2=0
r113 44 47 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.165 $Y=0
+ $X2=8.88 $Y2=0
r114 43 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r115 42 43 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r116 40 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r117 39 42 407.102 $w=1.68e-07 $l=6.24e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=7.92
+ $Y2=0
r118 39 40 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r119 37 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.21
+ $Y2=0
r120 37 39 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.375 $Y=0
+ $X2=1.68 $Y2=0
r121 36 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.305 $Y=0 $X2=8.47
+ $Y2=0
r122 36 42 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=8.305 $Y=0
+ $X2=7.92 $Y2=0
r123 35 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r124 35 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r125 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r126 32 55 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r127 32 34 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.72 $Y2=0
r128 31 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.21
+ $Y2=0
r129 31 34 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=0
+ $X2=0.72 $Y2=0
r130 29 43 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=7.92 $Y2=0
r131 29 40 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=1.68 $Y2=0
r132 25 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.33 $Y=0.085
+ $X2=9.33 $Y2=0
r133 25 27 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=9.33 $Y=0.085
+ $X2=9.33 $Y2=0.675
r134 21 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.47 $Y=0.085
+ $X2=8.47 $Y2=0
r135 21 23 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=8.47 $Y=0.085
+ $X2=8.47 $Y2=0.675
r136 17 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0
r137 17 19 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0.675
r138 13 55 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r139 13 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.515
r140 4 27 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=9.19
+ $Y=0.37 $X2=9.33 $Y2=0.675
r141 3 23 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=8.33
+ $Y=0.37 $X2=8.47 $Y2=0.675
r142 2 19 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.37 $X2=1.21 $Y2=0.675
r143 1 15 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__A41OI_4%A_325_74# 1 2 3 4 5 18 20 21 24 26 34 36 38
r63 32 34 27.1535 $w=3.63e-07 $l=8.6e-07 $layer=LI1_cond $X=4.9 $Y=0.437
+ $X2=5.76 $Y2=0.437
r64 30 38 6.12952 $w=2.67e-07 $l=1.65e-07 $layer=LI1_cond $X=4.135 $Y=0.437
+ $X2=3.97 $Y2=0.437
r65 30 32 24.1539 $w=3.63e-07 $l=7.65e-07 $layer=LI1_cond $X=4.135 $Y=0.437
+ $X2=4.9 $Y2=0.437
r66 27 36 11.6921 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=3.135 $Y=0.34
+ $X2=2.87 $Y2=0.34
r67 26 38 6.12952 $w=2.67e-07 $l=2.07918e-07 $layer=LI1_cond $X=3.805 $Y=0.34
+ $X2=3.97 $Y2=0.437
r68 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.805 $Y=0.34
+ $X2=3.135 $Y2=0.34
r69 22 36 2.222 $w=5.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=0.425 $X2=2.87
+ $Y2=0.34
r70 22 24 2.03108 $w=5.28e-07 $l=9e-08 $layer=LI1_cond $X=2.87 $Y=0.425 $X2=2.87
+ $Y2=0.515
r71 20 36 11.6921 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=2.605 $Y=0.34
+ $X2=2.87 $Y2=0.34
r72 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.605 $Y=0.34
+ $X2=1.935 $Y2=0.34
r73 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.77 $Y=0.425
+ $X2=1.935 $Y2=0.34
r74 16 18 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.77 $Y=0.425
+ $X2=1.77 $Y2=0.655
r75 5 34 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.62
+ $Y=0.37 $X2=5.76 $Y2=0.515
r76 4 32 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.76
+ $Y=0.37 $X2=4.9 $Y2=0.515
r77 3 38 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=3.76
+ $Y=0.37 $X2=3.97 $Y2=0.515
r78 2 24 45.5 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_NDIFF $count=4 $X=2.56
+ $Y=0.37 $X2=3.04 $Y2=0.515
r79 1 18 182 $w=1.7e-07 $l=3.50071e-07 $layer=licon1_NDIFF $count=1 $X=1.625
+ $Y=0.37 $X2=1.77 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_MS__A41OI_4%A_852_74# 1 2 3 4 22 23
c31 22 0 1.35727e-19 $X=7.61 $Y=0.95
r32 22 23 5.33064 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=7.61 $Y=0.95
+ $X2=7.445 $Y2=0.95
r33 20 23 23.5573 $w=3.38e-07 $l=6.95e-07 $layer=LI1_cond $X=6.75 $Y=0.96
+ $X2=7.445 $Y2=0.96
r34 18 20 48.1314 $w=3.38e-07 $l=1.42e-06 $layer=LI1_cond $X=5.33 $Y=0.96
+ $X2=6.75 $Y2=0.96
r35 15 18 29.15 $w=3.38e-07 $l=8.6e-07 $layer=LI1_cond $X=4.47 $Y=0.96 $X2=5.33
+ $Y2=0.96
r36 4 22 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=7.47
+ $Y=0.37 $X2=7.61 $Y2=0.95
r37 3 20 182 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_NDIFF $count=1 $X=6.61
+ $Y=0.37 $X2=6.75 $Y2=0.96
r38 2 18 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=5.19
+ $Y=0.37 $X2=5.33 $Y2=0.95
r39 1 15 182 $w=1.7e-07 $l=6.76905e-07 $layer=licon1_NDIFF $count=1 $X=4.26
+ $Y=0.37 $X2=4.47 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_MS__A41OI_4%A_1235_74# 1 2 3 4 5 16 20 24 25 28 30 34 39
+ 42
c55 39 0 9.28144e-20 $X=6.485 $Y=0.485
c56 20 0 1.6164e-19 $X=8.04 $Y=0.6
r57 37 39 7.12439 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.32 $Y=0.485
+ $X2=6.485 $Y2=0.485
r58 32 34 22.8184 $w=2.48e-07 $l=4.95e-07 $layer=LI1_cond $X=9.84 $Y=1.01
+ $X2=9.84 $Y2=0.515
r59 31 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.985 $Y=1.095
+ $X2=8.9 $Y2=1.095
r60 30 32 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.715 $Y=1.095
+ $X2=9.84 $Y2=1.01
r61 30 31 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=9.715 $Y=1.095
+ $X2=8.985 $Y2=1.095
r62 26 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.9 $Y=1.01 $X2=8.9
+ $Y2=1.095
r63 26 28 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=8.9 $Y=1.01 $X2=8.9
+ $Y2=0.515
r64 24 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.815 $Y=1.095
+ $X2=8.9 $Y2=1.095
r65 24 25 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.815 $Y=1.095
+ $X2=8.125 $Y2=1.095
r66 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.04 $Y=1.01
+ $X2=8.125 $Y2=1.095
r67 21 23 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=8.04 $Y=1.01
+ $X2=8.04 $Y2=0.965
r68 20 41 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.04 $Y=0.6 $X2=8.04
+ $Y2=0.475
r69 20 23 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.04 $Y=0.6
+ $X2=8.04 $Y2=0.965
r70 19 39 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=7.18 $Y=0.475
+ $X2=6.485 $Y2=0.475
r71 16 41 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.955 $Y=0.475
+ $X2=8.04 $Y2=0.475
r72 16 19 35.7257 $w=2.48e-07 $l=7.75e-07 $layer=LI1_cond $X=7.955 $Y=0.475
+ $X2=7.18 $Y2=0.475
r73 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.66
+ $Y=0.37 $X2=9.8 $Y2=0.515
r74 4 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.76
+ $Y=0.37 $X2=8.9 $Y2=0.515
r75 3 41 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.9
+ $Y=0.37 $X2=8.04 $Y2=0.515
r76 3 23 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=7.9
+ $Y=0.37 $X2=8.04 $Y2=0.965
r77 2 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.04
+ $Y=0.37 $X2=7.18 $Y2=0.515
r78 1 37 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=6.175
+ $Y=0.37 $X2=6.32 $Y2=0.525
.ends


* File: sky130_fd_sc_ms__dlrtp_2.spice
* Created: Wed Sep  2 12:05:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dlrtp_2.pex.spice"
.subckt sky130_fd_sc_ms__dlrtp_2  VNB VPB D GATE RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_D_M1012_g N_A_27_392#_M1012_s VNB NLOWVT L=0.15 W=0.55
+ AD=0.129591 AS=0.15675 PD=0.997674 PS=1.67 NRD=18 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75000.8 A=0.0825 P=1.4 MULT=1
MM1021 N_A_235_74#_M1021_d N_GATE_M1021_g N_VGND_M1012_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.174359 PD=2.05 PS=1.34233 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.7 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_VGND_M1001_d N_A_235_74#_M1001_g N_A_347_98#_M1001_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.205216 AS=0.2701 PD=1.59797 PS=2.21 NRD=36.048 NRS=12.972 M=1
+ R=4.93333 SA=75000.3 SB=75001.4 A=0.111 P=1.78 MULT=1
MM1003 A_568_74# N_A_27_392#_M1003_g N_VGND_M1001_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0768 AS=0.177484 PD=0.88 PS=1.38203 NRD=12.18 NRS=15.936 M=1 R=4.26667
+ SA=75000.8 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1004 N_A_646_74#_M1004_d N_A_347_98#_M1004_g A_568_74# VNB NLOWVT L=0.15
+ W=0.64 AD=0.194158 AS=0.0768 PD=1.42491 PS=0.88 NRD=16.872 NRS=12.18 M=1
+ R=4.26667 SA=75001.2 SB=75001 A=0.096 P=1.58 MULT=1
MM1019 A_784_81# N_A_235_74#_M1019_g N_A_646_74#_M1004_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.127417 PD=0.66 PS=0.935094 NRD=18.564 NRS=48.564 M=1
+ R=2.8 SA=75001.8 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_832_55#_M1020_g A_784_81# VNB NLOWVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 A_1060_74# N_A_646_74#_M1017_g N_A_832_55#_M1017_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.0888 AS=0.2109 PD=0.98 PS=2.05 NRD=10.536 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001.7 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_RESET_B_M1005_g A_1060_74# VNB NLOWVT L=0.15 W=0.74
+ AD=0.1628 AS=0.0888 PD=1.18 PS=0.98 NRD=14.592 NRS=10.536 M=1 R=4.93333
+ SA=75000.6 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1006 N_Q_M1006_d N_A_832_55#_M1006_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1073 AS=0.1628 PD=1.03 PS=1.18 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.2
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1018 N_Q_M1006_d N_A_832_55#_M1018_g N_VGND_M1018_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1073 AS=0.2553 PD=1.03 PS=2.17 NRD=1.62 NRS=9.72 M=1 R=4.93333 SA=75001.6
+ SB=75000.3 A=0.111 P=1.78 MULT=1
MM1002 N_VPWR_M1002_d N_D_M1002_g N_A_27_392#_M1002_s VPB PSHORT L=0.18 W=0.84
+ AD=0.22685 AS=0.2352 PD=1.57 PS=2.24 NRD=50.432 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90000.8 A=0.1512 P=2.04 MULT=1
MM1015 N_A_235_74#_M1015_d N_GATE_M1015_g N_VPWR_M1002_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2352 AS=0.22685 PD=2.24 PS=1.57 NRD=0 NRS=50.432 M=1 R=4.66667
+ SA=90000.8 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1007 N_VPWR_M1007_d N_A_235_74#_M1007_g N_A_347_98#_M1007_s VPB PSHORT L=0.18
+ W=0.84 AD=0.210023 AS=0.2352 PD=1.42891 PS=2.24 NRD=45.7237 NRS=0 M=1
+ R=4.66667 SA=90000.2 SB=90002.3 A=0.1512 P=2.04 MULT=1
MM1014 A_568_392# N_A_27_392#_M1014_g N_VPWR_M1007_d VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.250027 PD=1.24 PS=1.70109 NRD=12.7853 NRS=15.7403 M=1 R=5.55556
+ SA=90000.7 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1016 N_A_646_74#_M1016_d N_A_235_74#_M1016_g A_568_392# VPB PSHORT L=0.18 W=1
+ AD=0.219366 AS=0.12 PD=1.90845 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556
+ SA=90001.1 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1000 A_759_508# N_A_347_98#_M1000_g N_A_646_74#_M1016_d VPB PSHORT L=0.18
+ W=0.42 AD=0.10605 AS=0.0921338 PD=0.925 PS=0.801549 NRD=92.6294 NRS=39.8531
+ M=1 R=2.33333 SA=90001.6 SB=90003.2 A=0.0756 P=1.2 MULT=1
MM1011 N_VPWR_M1011_d N_A_832_55#_M1011_g A_759_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.119318 AS=0.10605 PD=0.951818 PS=0.925 NRD=68.0044 NRS=92.6294 M=1
+ R=2.33333 SA=90002.2 SB=90002.5 A=0.0756 P=1.2 MULT=1
MM1009 N_A_832_55#_M1009_d N_A_646_74#_M1009_g N_VPWR_M1011_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.318182 PD=1.39 PS=2.53818 NRD=0 NRS=35.1645 M=1
+ R=6.22222 SA=90001.2 SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1010 N_VPWR_M1010_d N_RESET_B_M1010_g N_A_832_55#_M1009_d VPB PSHORT L=0.18
+ W=1.12 AD=0.2072 AS=0.1512 PD=1.49 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90001.7 SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1008 N_Q_M1008_d N_A_832_55#_M1008_g N_VPWR_M1010_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1596 AS=0.2072 PD=1.405 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.2
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1013 N_Q_M1008_d N_A_832_55#_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1596 AS=0.3528 PD=1.405 PS=2.87 NRD=1.7533 NRS=5.2599 M=1 R=6.22222
+ SA=90002.7 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX22_noxref VNB VPB NWDIODE A=14.0988 P=18.88
c_1051 A_784_81# 0 1.78997e-19 $X=3.92 $Y=0.405
*
.include "sky130_fd_sc_ms__dlrtp_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__dlrbn_1.pex.spice
* Created: Wed Sep  2 12:04:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__DLRBN_1%D 2 5 9 11 12 15
r35 15 17 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.425
+ $X2=0.59 $Y2=1.26
r36 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.6
+ $Y=1.425 $X2=0.6 $Y2=1.425
r37 12 16 2.24265 $w=6.38e-07 $l=1.2e-07 $layer=LI1_cond $X=0.72 $Y=1.58 $X2=0.6
+ $Y2=1.58
r38 9 17 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=0.5 $Y=0.835 $X2=0.5
+ $Y2=1.26
r39 5 11 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=0.505 $Y=2.54
+ $X2=0.505 $Y2=1.93
r40 2 11 42.4214 $w=3.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.59 $Y=1.755
+ $X2=0.59 $Y2=1.93
r41 1 15 1.64869 $w=3.5e-07 $l=1e-08 $layer=POLY_cond $X=0.59 $Y=1.435 $X2=0.59
+ $Y2=1.425
r42 1 2 52.7581 $w=3.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.59 $Y=1.435 $X2=0.59
+ $Y2=1.755
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_1%GATE_N 3 6 9 11 12 15 16
r36 15 17 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.425
+ $X2=1.18 $Y2=1.26
r37 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.17
+ $Y=1.425 $X2=1.17 $Y2=1.425
r38 12 16 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.17 $Y=1.665
+ $X2=1.17 $Y2=1.425
r39 9 11 237.113 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=1.265 $Y=2.54
+ $X2=1.265 $Y2=1.93
r40 6 11 42.4214 $w=3.5e-07 $l=1.75e-07 $layer=POLY_cond $X=1.18 $Y=1.755
+ $X2=1.18 $Y2=1.93
r41 5 15 1.64869 $w=3.5e-07 $l=1e-08 $layer=POLY_cond $X=1.18 $Y=1.435 $X2=1.18
+ $Y2=1.425
r42 5 6 52.7581 $w=3.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.18 $Y=1.435 $X2=1.18
+ $Y2=1.755
r43 3 17 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.08 $Y=0.74 $X2=1.08
+ $Y2=1.26
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_1%A_231_74# 1 2 9 12 16 19 23 26 27 30 32 33
+ 34 37 38 41 44 45 49 53 57 59 63 66 69
c149 53 0 9.3463e-20 $X=2.35 $Y=1.385
c150 26 0 5.58535e-20 $X=2.47 $Y=2.22
r151 63 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.445 $Y=1.285
+ $X2=3.445 $Y2=1.12
r152 62 64 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.445 $Y=1.285
+ $X2=3.445 $Y2=1.45
r153 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.445
+ $Y=1.285 $X2=3.445 $Y2=1.285
r154 59 62 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=3.445 $Y=1.215
+ $X2=3.445 $Y2=1.285
r155 55 57 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.205 $Y=2.055
+ $X2=3.365 $Y2=2.055
r156 53 67 40.9207 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.332 $Y=1.385
+ $X2=2.332 $Y2=1.55
r157 53 66 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.332 $Y=1.385
+ $X2=2.332 $Y2=1.22
r158 52 54 8.53881 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.37 $Y=1.385
+ $X2=2.37 $Y2=1.55
r159 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.35
+ $Y=1.385 $X2=2.35 $Y2=1.385
r160 49 52 5.29501 $w=3.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.37 $Y=1.215
+ $X2=2.37 $Y2=1.385
r161 44 47 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.54 $Y=2.305
+ $X2=1.54 $Y2=2.33
r162 44 45 10.3232 $w=2.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.54 $Y=2.305
+ $X2=1.54 $Y2=2.1
r163 43 45 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=1.59 $Y=1.09
+ $X2=1.59 $Y2=2.1
r164 41 43 18.7979 $w=5.43e-07 $l=5.75e-07 $layer=LI1_cond $X=1.402 $Y=0.515
+ $X2=1.402 $Y2=1.09
r165 38 71 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=4.125 $Y=2.215
+ $X2=3.935 $Y2=2.215
r166 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.125
+ $Y=2.215 $X2=4.125 $Y2=2.215
r167 35 37 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=4.125 $Y=2.905
+ $X2=4.125 $Y2=2.215
r168 33 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.96 $Y=2.99
+ $X2=4.125 $Y2=2.905
r169 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.96 $Y=2.99
+ $X2=3.29 $Y2=2.99
r170 32 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.365 $Y=1.97
+ $X2=3.365 $Y2=2.055
r171 32 64 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.365 $Y=1.97
+ $X2=3.365 $Y2=1.45
r172 30 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.205 $Y=2.905
+ $X2=3.29 $Y2=2.99
r173 29 55 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.205 $Y=2.14
+ $X2=3.205 $Y2=2.055
r174 29 30 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=3.205 $Y=2.14
+ $X2=3.205 $Y2=2.905
r175 28 49 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.555 $Y=1.215
+ $X2=2.37 $Y2=1.215
r176 27 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.28 $Y=1.215
+ $X2=3.445 $Y2=1.215
r177 27 28 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.28 $Y=1.215
+ $X2=2.555 $Y2=1.215
r178 26 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.47 $Y=2.22
+ $X2=2.47 $Y2=1.55
r179 24 44 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.675 $Y=2.305
+ $X2=1.54 $Y2=2.305
r180 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.385 $Y=2.305
+ $X2=2.47 $Y2=2.22
r181 23 24 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.385 $Y=2.305
+ $X2=1.675 $Y2=2.305
r182 17 71 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.935 $Y=2.38
+ $X2=3.935 $Y2=2.215
r183 17 19 143.823 $w=1.8e-07 $l=3.7e-07 $layer=POLY_cond $X=3.935 $Y=2.38
+ $X2=3.935 $Y2=2.75
r184 16 69 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.355 $Y=0.69
+ $X2=3.355 $Y2=1.12
r185 12 67 322.629 $w=1.8e-07 $l=8.3e-07 $layer=POLY_cond $X=2.36 $Y=2.38
+ $X2=2.36 $Y2=1.55
r186 9 66 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.225 $Y=0.74
+ $X2=2.225 $Y2=1.22
r187 2 47 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=1.355
+ $Y=2.12 $X2=1.49 $Y2=2.33
r188 1 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.155
+ $Y=0.37 $X2=1.295 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_1%A_27_424# 1 2 9 13 15 19 22 24 27 28 29 30
+ 33 34 35 36 41 42
c103 41 0 2.24964e-19 $X=2.905 $Y=1.635
c104 33 0 1.66804e-19 $X=2.825 $Y=2.56
r105 42 47 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.905 $Y=1.635
+ $X2=2.905 $Y2=1.8
r106 42 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.905 $Y=1.635
+ $X2=2.905 $Y2=1.47
r107 41 44 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.905 $Y=1.635
+ $X2=2.905 $Y2=1.8
r108 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.905
+ $Y=1.635 $X2=2.905 $Y2=1.635
r109 36 38 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.93 $Y=2.645
+ $X2=1.93 $Y2=2.815
r110 33 44 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.825 $Y=2.56
+ $X2=2.825 $Y2=1.8
r111 31 36 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.015 $Y=2.645
+ $X2=1.93 $Y2=2.645
r112 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.74 $Y=2.645
+ $X2=2.825 $Y2=2.56
r113 30 31 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=2.74 $Y=2.645
+ $X2=2.015 $Y2=2.645
r114 28 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.845 $Y=2.815
+ $X2=1.93 $Y2=2.815
r115 28 29 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.845 $Y=2.815
+ $X2=1.235 $Y2=2.815
r116 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.15 $Y=2.73
+ $X2=1.235 $Y2=2.815
r117 26 27 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.15 $Y=2.24
+ $X2=1.15 $Y2=2.73
r118 25 35 2.28545 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.365 $Y=2.155
+ $X2=0.23 $Y2=2.155
r119 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.065 $Y=2.155
+ $X2=1.15 $Y2=2.24
r120 24 25 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.065 $Y=2.155
+ $X2=0.365 $Y2=2.155
r121 20 35 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.23 $Y=2.24
+ $X2=0.23 $Y2=2.155
r122 20 22 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.23 $Y=2.24
+ $X2=0.23 $Y2=2.265
r123 19 35 4.14756 $w=2.2e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.18 $Y=2.07
+ $X2=0.23 $Y2=2.155
r124 19 34 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=0.18 $Y=2.07
+ $X2=0.18 $Y2=1.09
r125 15 34 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=0.272 $Y=0.913
+ $X2=0.272 $Y2=1.09
r126 15 17 3.36789 $w=3.55e-07 $l=9.8e-08 $layer=LI1_cond $X=0.272 $Y=0.913
+ $X2=0.272 $Y2=0.815
r127 13 47 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.98 $Y=2.46
+ $X2=2.98 $Y2=1.8
r128 9 46 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.965 $Y=0.69
+ $X2=2.965 $Y2=1.47
r129 2 22 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.12 $X2=0.28 $Y2=2.265
r130 1 17 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.56 $X2=0.285 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_1%A_373_74# 1 2 7 9 10 11 13 16 19 22 23 27 28
+ 30 34 37
c96 23 0 1.8903e-19 $X=3.875 $Y=0.865
c97 11 0 2.98305e-19 $X=3.49 $Y=1.765
r98 31 34 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.93 $Y=1.885
+ $X2=2.05 $Y2=1.885
r99 28 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.04 $Y=1.285
+ $X2=4.04 $Y2=1.45
r100 28 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.04 $Y=1.285
+ $X2=4.04 $Y2=1.12
r101 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.04
+ $Y=1.285 $X2=4.04 $Y2=1.285
r102 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.04 $Y=0.95
+ $X2=4.04 $Y2=1.285
r103 24 30 2.76166 $w=1.7e-07 $l=1.67481e-07 $layer=LI1_cond $X=2.175 $Y=0.865
+ $X2=2.01 $Y2=0.87
r104 23 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.875 $Y=0.865
+ $X2=4.04 $Y2=0.95
r105 23 24 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=3.875 $Y=0.865
+ $X2=2.175 $Y2=0.865
r106 22 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.93 $Y=1.72
+ $X2=1.93 $Y2=1.885
r107 21 30 3.70735 $w=2.5e-07 $l=1.23693e-07 $layer=LI1_cond $X=1.93 $Y=0.96
+ $X2=2.01 $Y2=0.87
r108 21 22 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=1.93 $Y=0.96
+ $X2=1.93 $Y2=1.72
r109 17 30 3.70735 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=2.01 $Y=0.78 $X2=2.01
+ $Y2=0.87
r110 17 19 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.01 $Y=0.78
+ $X2=2.01 $Y2=0.515
r111 16 37 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.13 $Y=0.8
+ $X2=4.13 $Y2=1.12
r112 13 38 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.95 $Y=1.69
+ $X2=3.95 $Y2=1.45
r113 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.875 $Y=1.765
+ $X2=3.95 $Y2=1.69
r114 10 11 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=3.875 $Y=1.765
+ $X2=3.49 $Y2=1.765
r115 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.4 $Y=1.84
+ $X2=3.49 $Y2=1.765
r116 7 9 166.022 $w=1.8e-07 $l=6.2e-07 $layer=POLY_cond $X=3.4 $Y=1.84 $X2=3.4
+ $Y2=2.46
r117 2 34 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.905
+ $Y=1.74 $X2=2.05 $Y2=1.885
r118 1 19 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.865
+ $Y=0.37 $X2=2.01 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_1%A_889_92# 1 2 9 11 13 15 17 20 24 28 30 31
+ 32 33 42 45 48 50 53 54 56 59 63
c136 53 0 1.11337e-19 $X=6.435 $Y=1.72
c137 20 0 1.44146e-19 $X=6.535 $Y=2.27
c138 9 0 1.8903e-19 $X=4.52 $Y=0.8
r139 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.645
+ $Y=1.385 $X2=6.645 $Y2=1.385
r140 60 63 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=6.435 $Y=1.385
+ $X2=6.645 $Y2=1.385
r141 58 59 9.96101 $w=5.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.78 $Y=2.005
+ $X2=5.945 $Y2=2.005
r142 55 58 8.49845 $w=5.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.375 $Y=2.005
+ $X2=5.78 $Y2=2.005
r143 55 56 3.88629 $w=5.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.375 $Y=2.005
+ $X2=5.29 $Y2=2.005
r144 52 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.435 $Y=1.55
+ $X2=6.435 $Y2=1.385
r145 52 53 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.435 $Y=1.55
+ $X2=6.435 $Y2=1.72
r146 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.35 $Y=1.805
+ $X2=6.435 $Y2=1.72
r147 50 59 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=6.35 $Y=1.805
+ $X2=5.945 $Y2=1.805
r148 46 58 3.93508 $w=3.3e-07 $l=2.85e-07 $layer=LI1_cond $X=5.78 $Y=2.29
+ $X2=5.78 $Y2=2.005
r149 46 48 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=5.78 $Y=2.29
+ $X2=5.78 $Y2=2.685
r150 45 55 7.98728 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=5.375 $Y=1.72
+ $X2=5.375 $Y2=2.005
r151 45 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.375 $Y=1.72
+ $X2=5.375 $Y2=1.05
r152 40 54 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=5.335 $Y=0.925
+ $X2=5.335 $Y2=1.05
r153 40 42 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=5.335 $Y=0.925
+ $X2=5.335 $Y2=0.515
r154 37 56 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=4.695 $Y=2.125
+ $X2=5.29 $Y2=2.125
r155 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.695
+ $Y=2.125 $X2=4.695 $Y2=2.125
r156 32 64 100.982 $w=3.6e-07 $l=6.3e-07 $layer=POLY_cond $X=7.275 $Y=1.4
+ $X2=6.645 $Y2=1.4
r157 31 34 66.6233 $w=4.1e-07 $l=3.6e-07 $layer=POLY_cond $X=7.48 $Y=1.4
+ $X2=7.48 $Y2=1.76
r158 31 33 47.9425 $w=4.1e-07 $l=1.8e-07 $layer=POLY_cond $X=7.48 $Y=1.4
+ $X2=7.48 $Y2=1.22
r159 31 32 5.91772 $w=3.6e-07 $l=2.05e-07 $layer=POLY_cond $X=7.48 $Y=1.4
+ $X2=7.275 $Y2=1.4
r160 29 64 3.20579 $w=3.6e-07 $l=2e-08 $layer=POLY_cond $X=6.625 $Y=1.4
+ $X2=6.645 $Y2=1.4
r161 29 30 4.93351 $w=3.6e-07 $l=9e-08 $layer=POLY_cond $X=6.625 $Y=1.4
+ $X2=6.535 $Y2=1.4
r162 28 33 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=7.61 $Y=0.835
+ $X2=7.61 $Y2=1.22
r163 24 34 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=7.595 $Y=2.34
+ $X2=7.595 $Y2=1.76
r164 18 30 36.864 $w=1.65e-07 $l=1.8e-07 $layer=POLY_cond $X=6.535 $Y=1.58
+ $X2=6.535 $Y2=1.4
r165 18 20 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=6.535 $Y=1.58
+ $X2=6.535 $Y2=2.27
r166 15 30 36.864 $w=1.65e-07 $l=1.8735e-07 $layer=POLY_cond $X=6.52 $Y=1.22
+ $X2=6.535 $Y2=1.4
r167 15 17 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.52 $Y=1.22
+ $X2=6.52 $Y2=0.74
r168 11 38 34.8237 $w=2.7e-07 $l=1.80291e-07 $layer=POLY_cond $X=4.62 $Y=2.29
+ $X2=4.652 $Y2=2.125
r169 11 13 178.806 $w=1.8e-07 $l=4.6e-07 $layer=POLY_cond $X=4.62 $Y=2.29
+ $X2=4.62 $Y2=2.75
r170 7 38 87.1026 $w=2.7e-07 $l=4.96634e-07 $layer=POLY_cond $X=4.52 $Y=1.69
+ $X2=4.652 $Y2=2.125
r171 7 9 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=4.52 $Y=1.69 $X2=4.52
+ $Y2=0.8
r172 2 58 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.635
+ $Y=1.71 $X2=5.78 $Y2=1.885
r173 2 48 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=5.635
+ $Y=1.71 $X2=5.78 $Y2=2.685
r174 1 42 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=5.23
+ $Y=0.37 $X2=5.375 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_1%A_686_74# 1 2 9 11 13 14 15 16 22 23 28 32
+ 33 35 36
r95 35 37 10.5366 $w=3.48e-07 $l=3.2e-07 $layer=LI1_cond $X=4.55 $Y=1.385
+ $X2=4.55 $Y2=1.705
r96 35 36 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.55 $Y=1.385
+ $X2=4.55 $Y2=1.22
r97 32 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.625 $Y=2.57
+ $X2=3.625 $Y2=2.405
r98 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.005
+ $Y=1.385 $X2=5.005 $Y2=1.385
r99 26 35 1.07274 $w=3.3e-07 $l=1.75e-07 $layer=LI1_cond $X=4.725 $Y=1.385
+ $X2=4.55 $Y2=1.385
r100 26 28 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=4.725 $Y=1.385
+ $X2=5.005 $Y2=1.385
r101 24 36 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.46 $Y=0.61
+ $X2=4.46 $Y2=1.22
r102 22 37 4.974 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=4.375 $Y=1.705
+ $X2=4.55 $Y2=1.705
r103 22 23 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=4.375 $Y=1.705
+ $X2=3.79 $Y2=1.705
r104 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.705 $Y=1.79
+ $X2=3.79 $Y2=1.705
r105 20 33 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=3.705 $Y=1.79
+ $X2=3.705 $Y2=2.405
r106 16 24 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.375 $Y=0.485
+ $X2=4.46 $Y2=0.61
r107 16 18 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=4.375 $Y=0.485
+ $X2=3.72 $Y2=0.485
r108 14 29 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=5.455 $Y=1.385
+ $X2=5.005 $Y2=1.385
r109 14 15 3.90195 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.455 $Y=1.385
+ $X2=5.455 $Y2=1.22
r110 11 15 34.7346 $w=1.65e-07 $l=1.35e-07 $layer=POLY_cond $X=5.59 $Y=1.22
+ $X2=5.455 $Y2=1.22
r111 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.59 $Y=1.22
+ $X2=5.59 $Y2=0.74
r112 7 15 34.7346 $w=1.65e-07 $l=3.7229e-07 $layer=POLY_cond $X=5.545 $Y=1.55
+ $X2=5.455 $Y2=1.22
r113 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=5.545 $Y=1.55
+ $X2=5.545 $Y2=2.27
r114 2 32 600 $w=1.7e-07 $l=6.74129e-07 $layer=licon1_PDIFF $count=1 $X=3.49
+ $Y=1.96 $X2=3.625 $Y2=2.57
r115 1 18 182 $w=1.7e-07 $l=3.59235e-07 $layer=licon1_NDIFF $count=1 $X=3.43
+ $Y=0.37 $X2=3.72 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_1%RESET_B 3 6 8 11 13
c35 13 0 1.84321e-19 $X=6.04 $Y=1.22
r36 11 14 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.04 $Y=1.385
+ $X2=6.04 $Y2=1.55
r37 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.04 $Y=1.385
+ $X2=6.04 $Y2=1.22
r38 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.04
+ $Y=1.385 $X2=6.04 $Y2=1.385
r39 8 12 3.40065 $w=3.03e-07 $l=9e-08 $layer=LI1_cond $X=6.027 $Y=1.295
+ $X2=6.027 $Y2=1.385
r40 6 14 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=6.005 $Y=2.27
+ $X2=6.005 $Y2=1.55
r41 3 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.98 $Y=0.74 $X2=5.98
+ $Y2=1.22
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_1%A_1437_112# 1 2 9 13 17 21 25 26 28
c42 21 0 1.44146e-19 $X=7.37 $Y=2.065
r43 26 31 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.06 $Y=1.465
+ $X2=8.06 $Y2=1.63
r44 26 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.06 $Y=1.465
+ $X2=8.06 $Y2=1.3
r45 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.06
+ $Y=1.465 $X2=8.06 $Y2=1.465
r46 23 28 0.533013 $w=3.3e-07 $l=1.38e-07 $layer=LI1_cond $X=7.56 $Y=1.465
+ $X2=7.422 $Y2=1.465
r47 23 25 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=7.56 $Y=1.465 $X2=8.06
+ $Y2=1.465
r48 19 28 6.22203 $w=2.62e-07 $l=1.70895e-07 $layer=LI1_cond $X=7.41 $Y=1.63
+ $X2=7.422 $Y2=1.465
r49 19 21 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=7.41 $Y=1.63
+ $X2=7.41 $Y2=2.065
r50 15 28 6.22203 $w=2.62e-07 $l=1.65e-07 $layer=LI1_cond $X=7.422 $Y=1.3
+ $X2=7.422 $Y2=1.465
r51 15 17 19.4868 $w=2.73e-07 $l=4.65e-07 $layer=LI1_cond $X=7.422 $Y=1.3
+ $X2=7.422 $Y2=0.835
r52 13 30 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=8.125 $Y=0.74
+ $X2=8.125 $Y2=1.3
r53 9 31 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=8.135 $Y=2.4
+ $X2=8.135 $Y2=1.63
r54 2 21 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=7.245
+ $Y=1.92 $X2=7.37 $Y2=2.065
r55 1 17 182 $w=1.7e-07 $l=3.65205e-07 $layer=licon1_NDIFF $count=1 $X=7.185
+ $Y=0.56 $X2=7.395 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_1%VPWR 1 2 3 4 5 18 22 26 30 35 36 37 39 44 52
+ 64 73 74 77 80 83 90
c105 4 0 1.11337e-19 $X=6.095 $Y=1.71
r106 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r107 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r108 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r109 74 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r110 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r111 71 90 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=8.01 $Y=3.33
+ $X2=7.877 $Y2=3.33
r112 71 73 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=8.01 $Y=3.33
+ $X2=8.4 $Y2=3.33
r113 70 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r114 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r115 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r116 66 69 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r117 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r118 64 90 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=7.745 $Y=3.33
+ $X2=7.877 $Y2=3.33
r119 64 69 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.745 $Y=3.33
+ $X2=7.44 $Y2=3.33
r120 63 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r121 63 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.04
+ $Y2=3.33
r122 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r123 60 62 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=5.445 $Y=3.33
+ $X2=6 $Y2=3.33
r124 59 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r125 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r126 56 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r127 55 58 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r128 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r129 53 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=2.67 $Y2=3.33
r130 53 55 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=3.12 $Y2=3.33
r131 52 60 9.90988 $w=1.7e-07 $l=3.83e-07 $layer=LI1_cond $X=5.062 $Y=3.33
+ $X2=5.445 $Y2=3.33
r132 52 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r133 52 83 10.0846 $w=7.63e-07 $l=6.45e-07 $layer=LI1_cond $X=5.062 $Y=3.33
+ $X2=5.062 $Y2=2.685
r134 52 58 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.68 $Y=3.33
+ $X2=4.56 $Y2=3.33
r135 51 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r136 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r137 48 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r138 48 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r139 47 50 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r140 47 48 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r141 45 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r142 45 47 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r143 44 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.67 $Y2=3.33
r144 44 50 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.16 $Y2=3.33
r145 42 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r146 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r147 39 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r148 39 41 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r149 37 59 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r150 37 56 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=3.12 $Y2=3.33
r151 35 62 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.115 $Y=3.33
+ $X2=6 $Y2=3.33
r152 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.115 $Y=3.33
+ $X2=6.28 $Y2=3.33
r153 34 66 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=6.445 $Y=3.33
+ $X2=6.48 $Y2=3.33
r154 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.445 $Y=3.33
+ $X2=6.28 $Y2=3.33
r155 30 33 36.0954 $w=2.63e-07 $l=8.3e-07 $layer=LI1_cond $X=7.877 $Y=1.985
+ $X2=7.877 $Y2=2.815
r156 28 90 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=7.877 $Y=3.245
+ $X2=7.877 $Y2=3.33
r157 28 33 18.7 $w=2.63e-07 $l=4.3e-07 $layer=LI1_cond $X=7.877 $Y=3.245
+ $X2=7.877 $Y2=2.815
r158 24 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.28 $Y=3.245
+ $X2=6.28 $Y2=3.33
r159 24 26 38.4148 $w=3.28e-07 $l=1.1e-06 $layer=LI1_cond $X=6.28 $Y=3.245
+ $X2=6.28 $Y2=2.145
r160 20 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.67 $Y=3.245
+ $X2=2.67 $Y2=3.33
r161 20 22 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.67 $Y=3.245
+ $X2=2.67 $Y2=2.985
r162 16 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r163 16 18 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.495
r164 5 33 600 $w=1.7e-07 $l=1.0012e-06 $layer=licon1_PDIFF $count=1 $X=7.685
+ $Y=1.92 $X2=7.91 $Y2=2.815
r165 5 30 300 $w=1.7e-07 $l=2.55441e-07 $layer=licon1_PDIFF $count=2 $X=7.685
+ $Y=1.92 $X2=7.91 $Y2=1.985
r166 4 26 300 $w=1.7e-07 $l=5.19326e-07 $layer=licon1_PDIFF $count=2 $X=6.095
+ $Y=1.71 $X2=6.28 $Y2=2.145
r167 3 83 300 $w=1.7e-07 $l=6.38396e-07 $layer=licon1_PDIFF $count=2 $X=4.71
+ $Y=2.54 $X2=5.28 $Y2=2.685
r168 2 22 600 $w=1.7e-07 $l=1.12966e-06 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.96 $X2=2.67 $Y2=2.985
r169 1 18 300 $w=1.7e-07 $l=4.37321e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=2.12 $X2=0.73 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_1%Q 1 2 11 12 13 14 15 16 29
c32 29 0 1.84321e-19 $X=6.735 $Y=0.515
r33 16 26 7.59257 $w=4.23e-07 $l=2.8e-07 $layer=LI1_cond $X=6.902 $Y=2.405
+ $X2=6.902 $Y2=2.685
r34 15 16 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=6.902 $Y=2.035
+ $X2=6.902 $Y2=2.405
r35 14 35 8.96211 $w=5.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.84 $Y=0.925
+ $X2=6.84 $Y2=1.05
r36 13 14 8.04635 $w=5.48e-07 $l=3.7e-07 $layer=LI1_cond $X=6.84 $Y=0.555
+ $X2=6.84 $Y2=0.925
r37 13 29 0.869875 $w=5.48e-07 $l=4e-08 $layer=LI1_cond $X=6.84 $Y=0.555
+ $X2=6.84 $Y2=0.515
r38 12 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.03 $Y=1.72
+ $X2=7.03 $Y2=1.05
r39 11 12 8.76046 $w=4.23e-07 $l=1.65e-07 $layer=LI1_cond $X=6.902 $Y=1.885
+ $X2=6.902 $Y2=1.72
r40 9 15 2.79298 $w=4.23e-07 $l=1.03e-07 $layer=LI1_cond $X=6.902 $Y=1.932
+ $X2=6.902 $Y2=2.035
r41 9 11 1.27447 $w=4.23e-07 $l=4.7e-08 $layer=LI1_cond $X=6.902 $Y=1.932
+ $X2=6.902 $Y2=1.885
r42 2 26 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=6.625
+ $Y=1.71 $X2=6.775 $Y2=2.685
r43 2 11 400 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=6.625
+ $Y=1.71 $X2=6.775 $Y2=1.885
r44 1 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.595
+ $Y=0.37 $X2=6.735 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_1%Q_N 1 2 9 13 14 15 16 23 32
r18 21 23 1.65126 $w=3.33e-07 $l=4.8e-08 $layer=LI1_cond $X=8.362 $Y=1.987
+ $X2=8.362 $Y2=2.035
r19 15 16 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=8.362 $Y=2.405
+ $X2=8.362 $Y2=2.775
r20 14 21 0.653624 $w=3.33e-07 $l=1.9e-08 $layer=LI1_cond $X=8.362 $Y=1.968
+ $X2=8.362 $Y2=1.987
r21 14 32 7.88131 $w=3.33e-07 $l=1.48e-07 $layer=LI1_cond $X=8.362 $Y=1.968
+ $X2=8.362 $Y2=1.82
r22 14 15 12.1093 $w=3.33e-07 $l=3.52e-07 $layer=LI1_cond $X=8.362 $Y=2.053
+ $X2=8.362 $Y2=2.405
r23 14 23 0.619223 $w=3.33e-07 $l=1.8e-08 $layer=LI1_cond $X=8.362 $Y=2.053
+ $X2=8.362 $Y2=2.035
r24 13 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.445 $Y=1.13
+ $X2=8.445 $Y2=1.82
r25 7 13 7.60349 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=8.387 $Y=0.988
+ $X2=8.387 $Y2=1.13
r26 7 9 19.1265 $w=2.83e-07 $l=4.73e-07 $layer=LI1_cond $X=8.387 $Y=0.988
+ $X2=8.387 $Y2=0.515
r27 2 14 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.225
+ $Y=1.84 $X2=8.36 $Y2=1.985
r28 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=8.225
+ $Y=1.84 $X2=8.36 $Y2=2.815
r29 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.2 $Y=0.37
+ $X2=8.34 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__DLRBN_1%VGND 1 2 3 4 5 18 24 28 32 37 38 40 41 42 44
+ 49 70 79 80 83 87 93
r91 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r92 87 90 10.8067 $w=5.68e-07 $l=5.15e-07 $layer=LI1_cond $X=2.63 $Y=0 $X2=2.63
+ $Y2=0.515
r93 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r94 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r95 80 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r96 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r97 77 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.075 $Y=0 $X2=7.91
+ $Y2=0
r98 77 79 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.075 $Y=0 $X2=8.4
+ $Y2=0
r99 76 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r100 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r101 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r102 72 75 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r103 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r104 70 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.745 $Y=0 $X2=7.91
+ $Y2=0
r105 70 75 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.745 $Y=0
+ $X2=7.44 $Y2=0
r106 69 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r107 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r108 66 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r109 65 68 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r110 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r111 63 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r112 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r113 60 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r114 59 62 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.56
+ $Y2=0
r115 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r116 57 87 7.98728 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=2.63
+ $Y2=0
r117 57 59 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.915 $Y=0
+ $X2=3.12 $Y2=0
r118 56 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r119 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r120 53 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r121 53 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r122 52 55 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r123 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r124 50 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=0.795
+ $Y2=0
r125 50 52 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r126 49 87 7.98728 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=2.345 $Y=0 $X2=2.63
+ $Y2=0
r127 49 55 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.345 $Y=0
+ $X2=2.16 $Y2=0
r128 47 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r129 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r130 44 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.795
+ $Y2=0
r131 44 46 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.24
+ $Y2=0
r132 42 63 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.56 $Y2=0
r133 42 60 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.32 $Y=0 $X2=3.12
+ $Y2=0
r134 40 68 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=6.03 $Y=0 $X2=6 $Y2=0
r135 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.03 $Y=0 $X2=6.195
+ $Y2=0
r136 39 72 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=6.36 $Y=0 $X2=6.48
+ $Y2=0
r137 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.36 $Y=0 $X2=6.195
+ $Y2=0
r138 37 62 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.73 $Y=0 $X2=4.56
+ $Y2=0
r139 37 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.73 $Y=0 $X2=4.855
+ $Y2=0
r140 36 65 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=4.98 $Y=0 $X2=5.04
+ $Y2=0
r141 36 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.98 $Y=0 $X2=4.855
+ $Y2=0
r142 32 34 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=7.91 $Y=0.495
+ $X2=7.91 $Y2=0.965
r143 30 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0
r144 30 32 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=7.91 $Y=0.085
+ $X2=7.91 $Y2=0.495
r145 26 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.195 $Y=0.085
+ $X2=6.195 $Y2=0
r146 26 28 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.195 $Y=0.085
+ $X2=6.195 $Y2=0.495
r147 22 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.855 $Y=0.085
+ $X2=4.855 $Y2=0
r148 22 24 32.9599 $w=2.48e-07 $l=7.15e-07 $layer=LI1_cond $X=4.855 $Y=0.085
+ $X2=4.855 $Y2=0.8
r149 18 20 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.795 $Y=0.515
+ $X2=0.795 $Y2=0.925
r150 16 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=0.085
+ $X2=0.795 $Y2=0
r151 16 18 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.795 $Y=0.085
+ $X2=0.795 $Y2=0.515
r152 5 34 182 $w=1.7e-07 $l=5.05124e-07 $layer=licon1_NDIFF $count=1 $X=7.685
+ $Y=0.56 $X2=7.91 $Y2=0.965
r153 5 32 182 $w=1.7e-07 $l=2.55441e-07 $layer=licon1_NDIFF $count=1 $X=7.685
+ $Y=0.56 $X2=7.91 $Y2=0.495
r154 4 28 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=6.055
+ $Y=0.37 $X2=6.195 $Y2=0.495
r155 3 24 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=4.595
+ $Y=0.59 $X2=4.815 $Y2=0.8
r156 2 90 182 $w=1.7e-07 $l=3.95917e-07 $layer=licon1_NDIFF $count=1 $X=2.3
+ $Y=0.37 $X2=2.63 $Y2=0.515
r157 1 20 182 $w=1.7e-07 $l=4.62088e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.56 $X2=0.795 $Y2=0.925
r158 1 18 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.56 $X2=0.795 $Y2=0.515
.ends


* File: sky130_fd_sc_ms__sdfxtp_2.spice
* Created: Wed Sep  2 12:31:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__sdfxtp_2.pex.spice"
.subckt sky130_fd_sc_ms__sdfxtp_2  VNB VPB SCE D SCD CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1033 N_VGND_M1033_d N_SCE_M1033_g N_A_27_74#_M1033_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0735 AS=0.1386 PD=0.77 PS=1.5 NRD=19.992 NRS=7.14 M=1 R=2.8 SA=75000.3
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1015 A_223_74# N_A_27_74#_M1015_g N_VGND_M1033_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0735 PD=0.66 PS=0.77 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.8
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1016 N_A_301_74#_M1016_d N_D_M1016_g A_223_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.11655 AS=0.0504 PD=0.975 PS=0.66 NRD=38.568 NRS=18.564 M=1 R=2.8
+ SA=75001.1 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1013 A_442_74# N_SCE_M1013_g N_A_301_74#_M1016_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.11655 PD=0.66 PS=0.975 NRD=18.564 NRS=39.996 M=1 R=2.8
+ SA=75001.8 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_SCD_M1004_g A_442_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0968897 AS=0.0504 PD=0.84 PS=0.66 NRD=32.856 NRS=18.564 M=1 R=2.8
+ SA=75002.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1031 N_A_634_74#_M1031_d N_CLK_M1031_g N_VGND_M1004_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.17071 PD=2.05 PS=1.48 NRD=0 NRS=4.044 M=1 R=4.93333 SA=75001.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1030 N_A_846_74#_M1030_d N_A_634_74#_M1030_g N_VGND_M1030_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.2627 PD=2.05 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75000.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1001 N_A_1044_100#_M1001_d N_A_634_74#_M1001_g N_A_301_74#_M1001_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.15225 AS=0.1197 PD=1.145 PS=1.41 NRD=71.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.4 A=0.063 P=1.14 MULT=1
MM1007 A_1219_100# N_A_846_74#_M1007_g N_A_1044_100#_M1001_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0882 AS=0.15225 PD=0.84 PS=1.145 NRD=44.28 NRS=55.704 M=1 R=2.8
+ SA=75001.1 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_1287_320#_M1010_g A_1219_100# VNB NLOWVT L=0.15 W=0.42
+ AD=0.195473 AS=0.0882 PD=1.25567 PS=0.84 NRD=117.252 NRS=44.28 M=1 R=2.8
+ SA=75001.7 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1008 N_A_1287_320#_M1008_d N_A_1044_100#_M1008_g N_VGND_M1010_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.18975 AS=0.255977 PD=1.24 PS=1.64433 NRD=0 NRS=90.54 M=1
+ R=3.66667 SA=75002.1 SB=75002.1 A=0.0825 P=1.4 MULT=1
MM1011 N_A_1595_424#_M1011_d N_A_846_74#_M1011_g N_A_1287_320#_M1008_d VNB
+ NLOWVT L=0.15 W=0.55 AD=0.10674 AS=0.18975 PD=1.03196 PS=1.24 NRD=0 NRS=89.448
+ M=1 R=3.66667 SA=75003 SB=75001.3 A=0.0825 P=1.4 MULT=1
MM1021 A_1787_74# N_A_634_74#_M1021_g N_A_1595_424#_M1011_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0815103 PD=0.66 PS=0.788041 NRD=18.564 NRS=22.848 M=1
+ R=2.8 SA=75003.3 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_A_1829_398#_M1022_g A_1787_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0821897 AS=0.0504 PD=0.78931 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75003.7 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1017 N_A_1829_398#_M1017_d N_A_1595_424#_M1017_g N_VGND_M1022_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.14481 PD=2.05 PS=1.39069 NRD=0 NRS=11.34 M=1
+ R=4.93333 SA=75002.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_VGND_M1005_d N_A_1829_398#_M1005_g N_Q_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2627 AS=0.12025 PD=2.19 PS=1.065 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.3
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1024 N_VGND_M1024_d N_A_1829_398#_M1024_g N_Q_M1005_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2294 AS=0.12025 PD=2.1 PS=1.065 NRD=4.044 NRS=7.296 M=1 R=4.93333
+ SA=75000.8 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1002 N_VPWR_M1002_d N_SCE_M1002_g N_A_27_74#_M1002_s VPB PSHORT L=0.18 W=0.64
+ AD=0.1024 AS=0.1792 PD=0.96 PS=1.84 NRD=13.8491 NRS=0 M=1 R=3.55556 SA=90000.2
+ SB=90003 A=0.1152 P=1.64 MULT=1
MM1032 A_219_453# N_SCE_M1032_g N_VPWR_M1002_d VPB PSHORT L=0.18 W=0.64
+ AD=0.0768 AS=0.1024 PD=0.88 PS=0.96 NRD=19.9955 NRS=0 M=1 R=3.55556 SA=90000.7
+ SB=90002.5 A=0.1152 P=1.64 MULT=1
MM1006 N_A_301_74#_M1006_d N_D_M1006_g A_219_453# VPB PSHORT L=0.18 W=0.64
+ AD=0.1648 AS=0.0768 PD=1.155 PS=0.88 NRD=35.3812 NRS=19.9955 M=1 R=3.55556
+ SA=90001.1 SB=90002 A=0.1152 P=1.64 MULT=1
MM1029 A_442_453# N_A_27_74#_M1029_g N_A_301_74#_M1006_d VPB PSHORT L=0.18
+ W=0.64 AD=0.0768 AS=0.1648 PD=0.88 PS=1.155 NRD=19.9955 NRS=36.9178 M=1
+ R=3.55556 SA=90001.8 SB=90001.3 A=0.1152 P=1.64 MULT=1
MM1018 N_VPWR_M1018_d N_SCD_M1018_g A_442_453# VPB PSHORT L=0.18 W=0.64
+ AD=0.199536 AS=0.0768 PD=1.32364 PS=0.88 NRD=44.6205 NRS=19.9955 M=1 R=3.55556
+ SA=90002.2 SB=90000.9 A=0.1152 P=1.64 MULT=1
MM1012 N_A_634_74#_M1012_d N_CLK_M1012_g N_VPWR_M1018_d VPB PSHORT L=0.18 W=1.12
+ AD=0.3136 AS=0.349189 PD=2.8 PS=2.31636 NRD=0 NRS=25.4918 M=1 R=6.22222
+ SA=90001.8 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1019 N_A_846_74#_M1019_d N_A_634_74#_M1019_g N_VPWR_M1019_s VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.6258 PD=2.8 PS=3.53 NRD=0 NRS=27.2451 M=1 R=6.22222
+ SA=90000.4 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1023 N_A_1044_100#_M1023_d N_A_846_74#_M1023_g N_A_301_74#_M1023_s VPB PSHORT
+ L=0.18 W=0.42 AD=0.0567 AS=0.1176 PD=0.69 PS=1.4 NRD=0 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90004.4 A=0.0756 P=1.2 MULT=1
MM1025 A_1213_508# N_A_634_74#_M1025_g N_A_1044_100#_M1023_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0777 AS=0.0567 PD=0.79 PS=0.69 NRD=60.9715 NRS=0 M=1 R=2.33333
+ SA=90000.6 SB=90003.9 A=0.0756 P=1.2 MULT=1
MM1020 N_VPWR_M1020_d N_A_1287_320#_M1020_g A_1213_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.105 AS=0.0777 PD=0.893333 PS=0.79 NRD=0 NRS=60.9715 M=1 R=2.33333
+ SA=90001.2 SB=90003.4 A=0.0756 P=1.2 MULT=1
MM1027 N_A_1287_320#_M1027_d N_A_1044_100#_M1027_g N_VPWR_M1020_d VPB PSHORT
+ L=0.18 W=0.84 AD=0.21 AS=0.21 PD=1.34 PS=1.78667 NRD=0 NRS=52.7566 M=1
+ R=4.66667 SA=90001 SB=90001.9 A=0.1512 P=2.04 MULT=1
MM1003 N_A_1595_424#_M1003_d N_A_634_74#_M1003_g N_A_1287_320#_M1027_d VPB
+ PSHORT L=0.18 W=0.84 AD=0.1836 AS=0.21 PD=1.62667 PS=1.34 NRD=0 NRS=52.7566
+ M=1 R=4.66667 SA=90001.7 SB=90001.3 A=0.1512 P=2.04 MULT=1
MM1000 A_1707_496# N_A_846_74#_M1000_g N_A_1595_424#_M1003_d VPB PSHORT L=0.18
+ W=0.42 AD=0.1281 AS=0.0918 PD=1.03 PS=0.813333 NRD=117.254 NRS=49.25 M=1
+ R=2.33333 SA=90002.9 SB=90001.8 A=0.0756 P=1.2 MULT=1
MM1014 N_VPWR_M1014_d N_A_1829_398#_M1014_g A_1707_496# VPB PSHORT L=0.18 W=0.42
+ AD=0.119907 AS=0.1281 PD=0.95831 PS=1.03 NRD=0 NRS=117.254 M=1 R=2.33333
+ SA=90003.7 SB=90001 A=0.0756 P=1.2 MULT=1
MM1009 N_A_1829_398#_M1009_d N_A_1595_424#_M1009_g N_VPWR_M1014_d VPB PSHORT
+ L=0.18 W=1 AD=0.28 AS=0.285493 PD=2.56 PS=2.28169 NRD=0 NRS=0 M=1 R=5.55556
+ SA=90002 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1026 N_Q_M1026_d N_A_1829_398#_M1026_g N_VPWR_M1026_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1028 N_Q_M1026_d N_A_1829_398#_M1028_g N_VPWR_M1028_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX34_noxref VNB VPB NWDIODE A=23.0268 P=28.48
c_130 VNB 0 1.87953e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__sdfxtp_2.pxi.spice"
*
.ends
*
*

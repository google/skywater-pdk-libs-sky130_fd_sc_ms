* File: sky130_fd_sc_ms__and4bb_4.spice
* Created: Wed Sep  2 11:59:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__and4bb_4.pex.spice"
.subckt sky130_fd_sc_ms__and4bb_4  VNB VPB B_N A_N C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* A_N	A_N
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1023 N_VGND_M1023_d N_B_N_M1023_g N_A_27_74#_M1023_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1024 N_A_200_74#_M1024_d N_A_N_M1024_g N_VGND_M1023_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1915 AS=0.0896 PD=1.99 PS=0.92 NRD=13.116 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1009 N_A_475_388#_M1009_d N_A_200_74#_M1009_g N_A_412_140#_M1009_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.2272 PD=0.92 PS=1.99 NRD=0 NRS=13.116 M=1
+ R=4.26667 SA=75000.3 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1027 N_A_475_388#_M1009_d N_A_200_74#_M1027_g N_A_412_140#_M1027_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1000 N_A_685_140#_M1000_d N_A_27_74#_M1000_g N_A_412_140#_M1027_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.1 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1002 N_A_685_140#_M1000_d N_A_27_74#_M1002_g N_A_412_140#_M1002_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_A_685_140#_M1001_d N_C_M1001_g N_A_882_137#_M1001_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.2272 PD=0.92 PS=1.99 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75000.3 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1025 N_A_685_140#_M1001_d N_C_M1025_g N_A_882_137#_M1025_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1010 N_VGND_M1010_d N_D_M1010_g N_A_882_137#_M1010_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.6 A=0.096 P=1.58 MULT=1
MM1026 N_VGND_M1026_d N_D_M1026_g N_A_882_137#_M1010_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.115478 AS=0.0896 PD=1.01101 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1008 N_VGND_M1026_d N_A_475_388#_M1008_g N_X_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.133522 AS=0.1036 PD=1.16899 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333
+ SA=75001 SB=75001.6 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_A_475_388#_M1012_g N_X_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1406 AS=0.1036 PD=1.12 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75001.4
+ SB=75001.2 A=0.111 P=1.78 MULT=1
MM1013 N_VGND_M1012_d N_A_475_388#_M1013_g N_X_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1406 AS=0.1184 PD=1.12 PS=1.06 NRD=4.86 NRS=6.48 M=1 R=4.93333 SA=75002
+ SB=75000.7 A=0.111 P=1.78 MULT=1
MM1021 N_VGND_M1021_d N_A_475_388#_M1021_g N_X_M1013_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2146 AS=0.1184 PD=2.06 PS=1.06 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.4
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1003 N_VPWR_M1003_d N_B_N_M1003_g N_A_27_74#_M1003_s VPB PSHORT L=0.18 W=1
+ AD=0.185 AS=0.28 PD=1.37 PS=2.56 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90000.2
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1022 N_A_200_74#_M1022_d N_A_N_M1022_g N_VPWR_M1003_d VPB PSHORT L=0.18 W=1
+ AD=0.28 AS=0.185 PD=2.56 PS=1.37 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90000.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1015 N_A_475_388#_M1015_d N_A_200_74#_M1015_g N_VPWR_M1015_s VPB PSHORT L=0.18
+ W=1 AD=0.22 AS=0.305 PD=1.44 PS=2.61 NRD=15.7403 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90006.3 A=0.18 P=2.36 MULT=1
MM1017 N_A_475_388#_M1015_d N_A_200_74#_M1017_g N_VPWR_M1017_s VPB PSHORT L=0.18
+ W=1 AD=0.22 AS=0.145 PD=1.44 PS=1.29 NRD=15.7403 NRS=0 M=1 R=5.55556
+ SA=90000.8 SB=90005.7 A=0.18 P=2.36 MULT=1
MM1019 N_VPWR_M1017_s N_A_27_74#_M1019_g N_A_475_388#_M1019_s VPB PSHORT L=0.18
+ W=1 AD=0.145 AS=0.15 PD=1.29 PS=1.3 NRD=2.9353 NRS=4.9053 M=1 R=5.55556
+ SA=90001.3 SB=90005.2 A=0.18 P=2.36 MULT=1
MM1020 N_VPWR_M1020_d N_A_27_74#_M1020_g N_A_475_388#_M1019_s VPB PSHORT L=0.18
+ W=1 AD=0.185 AS=0.15 PD=1.37 PS=1.3 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90001.8
+ SB=90004.7 A=0.18 P=2.36 MULT=1
MM1016 N_A_475_388#_M1016_d N_C_M1016_g N_VPWR_M1020_d VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.185 PD=1.27 PS=1.37 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90002.3
+ SB=90004.2 A=0.18 P=2.36 MULT=1
MM1018 N_A_475_388#_M1016_d N_C_M1018_g N_VPWR_M1018_s VPB PSHORT L=0.18 W=1
+ AD=0.135 AS=0.595 PD=1.27 PS=2.19 NRD=0 NRS=8.8453 M=1 R=5.55556 SA=90002.8
+ SB=90003.7 A=0.18 P=2.36 MULT=1
MM1004 N_A_475_388#_M1004_d N_D_M1004_g N_VPWR_M1018_s VPB PSHORT L=0.18 W=1
+ AD=0.17125 AS=0.595 PD=1.425 PS=2.19 NRD=8.8453 NRS=0 M=1 R=5.55556 SA=90004.2
+ SB=90002.3 A=0.18 P=2.36 MULT=1
MM1014 N_A_475_388#_M1004_d N_D_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1
+ AD=0.17125 AS=0.183302 PD=1.425 PS=1.39151 NRD=0 NRS=16.2525 M=1 R=5.55556
+ SA=90004.2 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1005 N_X_M1005_d N_A_475_388#_M1005_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.205298 PD=1.39 PS=1.55849 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.3
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1006 N_X_M1005_d N_A_475_388#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90004.7
+ SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1007 N_X_M1007_d N_A_475_388#_M1007_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90005.2
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1011 N_X_M1007_d N_A_475_388#_M1011_g N_VPWR_M1011_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90005.6
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX28_noxref VNB VPB NWDIODE A=17.245 P=22.92
c_87 VNB 0 5.63592e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__and4bb_4.pxi.spice"
*
.ends
*
*

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
M1000 a_1273_392# B a_1063_392# VPB pshort w=1e+06u l=180000u
+  ad=8.3e+11p pd=7.66e+06u as=5.9e+11p ps=5.18e+06u
M1001 VGND a_193_277# X VNB nlowvt w=740000u l=150000u
+  ad=2.0924e+12p pd=1.558e+07u as=6.919e+11p ps=4.83e+06u
M1002 a_1273_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=1.5228e+12p ps=1.154e+07u
M1003 X a_193_277# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=9.184e+11p pd=6.12e+06u as=0p ps=0u
M1004 VPWR A a_1273_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_193_277# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_193_277# a_27_94# a_791_392# VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=8.3e+11p ps=7.66e+06u
M1007 VGND A a_193_277# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=1.4134e+12p ps=6.78e+06u
M1008 VGND D_N a_27_94# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1009 a_681_368# C_N VGND VNB nlowvt w=640000u l=150000u
+  ad=1.719e+11p pd=1.85e+06u as=0p ps=0u
M1010 a_791_392# a_27_94# a_193_277# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR D_N a_27_94# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1012 X a_193_277# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_193_277# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_193_277# B VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_193_277# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_791_392# a_681_368# a_1063_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_193_277# a_27_94# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1063_392# a_681_368# a_791_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_193_277# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_193_277# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_681_368# a_193_277# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_681_368# C_N VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1023 a_1063_392# B a_1273_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__nor3b_1 A B C_N VGND VNB VPB VPWR Y
X0 a_347_368# a_27_112# Y VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X1 a_27_112# C_N VGND VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X2 a_27_112# C_N VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X3 VPWR A a_263_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X4 VGND a_27_112# Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X6 Y B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X7 a_263_368# B a_347_368# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
.ends

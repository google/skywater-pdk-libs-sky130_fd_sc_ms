* File: sky130_fd_sc_ms__nor2_1.pex.spice
* Created: Fri Aug 28 17:46:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__NOR2_1%A 3 7 9 13 16
r27 15 16 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.505 $Y=1.465
+ $X2=0.515 $Y2=1.465
r28 12 15 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.29 $Y=1.465
+ $X2=0.505 $Y2=1.465
r29 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.465 $X2=0.29 $Y2=1.465
r30 9 13 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.29 $Y=1.665 $X2=0.29
+ $Y2=1.465
r31 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.3
+ $X2=0.515 $Y2=1.465
r32 5 7 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.515 $Y=1.3 $X2=0.515
+ $Y2=0.74
r33 1 15 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=1.465
r34 1 3 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.505 $Y=1.63
+ $X2=0.505 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__NOR2_1%B 3 7 9 15 16
r23 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.465 $X2=1.15 $Y2=1.465
r24 13 15 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.945 $Y=1.465
+ $X2=1.15 $Y2=1.465
r25 11 13 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=0.925 $Y=1.465
+ $X2=0.945 $Y2=1.465
r26 9 16 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=1.15 $Y=1.665 $X2=1.15
+ $Y2=1.465
r27 5 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=1.3
+ $X2=0.945 $Y2=1.465
r28 5 7 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.945 $Y=1.3 $X2=0.945
+ $Y2=0.74
r29 1 11 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.63
+ $X2=0.925 $Y2=1.465
r30 1 3 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.925 $Y=1.63
+ $X2=0.925 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__NOR2_1%VPWR 1 4 6 10 14 15
r16 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r17 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r18 12 18 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r19 12 14 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=1.2 $Y2=3.33
r20 10 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r21 10 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r22 6 9 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=0.28 $Y=2.115 $X2=0.28
+ $Y2=2.815
r23 4 18 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r24 4 9 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.28 $Y=3.245 $X2=0.28
+ $Y2=2.815
r25 1 9 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.815
r26 1 6 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.84 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__NOR2_1%Y 1 2 9 12 13 14 15
c26 12 0 1.80995e-20 $X=0.73 $Y=1.95
r27 14 15 7.05312 $w=6.4e-07 $l=3.7e-07 $layer=LI1_cond $X=0.98 $Y=2.405
+ $X2=0.98 $Y2=2.775
r28 14 19 5.52812 $w=6.4e-07 $l=2.9e-07 $layer=LI1_cond $X=0.98 $Y=2.405
+ $X2=0.98 $Y2=2.115
r29 12 19 10.6252 $w=6.4e-07 $l=3.22102e-07 $layer=LI1_cond $X=0.73 $Y=1.95
+ $X2=0.98 $Y2=2.115
r30 12 13 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.73 $Y=1.95
+ $X2=0.73 $Y2=1.13
r31 7 13 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.69 $Y=1.005
+ $X2=0.69 $Y2=1.13
r32 7 9 22.5879 $w=2.48e-07 $l=4.9e-07 $layer=LI1_cond $X=0.69 $Y=1.005 $X2=0.69
+ $Y2=0.515
r33 2 15 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.015
+ $Y=1.84 $X2=1.15 $Y2=2.815
r34 2 19 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.015
+ $Y=1.84 $X2=1.15 $Y2=2.115
r35 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.59
+ $Y=0.37 $X2=0.73 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__NOR2_1%VGND 1 2 7 9 11 13 15 17 27
r21 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r22 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r23 18 23 3.98448 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=0 $X2=0.192
+ $Y2=0
r24 18 20 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.385 $Y=0 $X2=0.72
+ $Y2=0
r25 17 26 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=1.217
+ $Y2=0
r26 17 20 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.995 $Y=0 $X2=0.72
+ $Y2=0
r27 15 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r28 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r29 15 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r30 11 26 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=1.16 $Y=0.085
+ $X2=1.217 $Y2=0
r31 11 13 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.16 $Y=0.085
+ $X2=1.16 $Y2=0.515
r32 7 23 3.15868 $w=2.5e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.192 $Y2=0
r33 7 9 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.26 $Y=0.085 $X2=0.26
+ $Y2=0.515
r34 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.02
+ $Y=0.37 $X2=1.16 $Y2=0.515
r35 1 9 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.155
+ $Y=0.37 $X2=0.3 $Y2=0.515
.ends


* File: sky130_fd_sc_ms__dfrbp_2.spice
* Created: Wed Sep  2 12:02:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dfrbp_2.pex.spice"
.subckt sky130_fd_sc_ms__dfrbp_2  VNB VPB D RESET_B CLK VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* CLK	CLK
* RESET_B	RESET_B
* D	D
* VPB	VPB
* VNB	VNB
MM1012 A_156_74# N_D_M1012_g N_A_70_74#_M1012_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1176 PD=0.63 PS=1.4 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1037 N_VGND_M1037_d N_RESET_B_M1037_g A_156_74# VNB NLOWVT L=0.15 W=0.42
+ AD=0.111861 AS=0.0441 PD=0.973966 PS=0.63 NRD=8.568 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1031 N_A_334_119#_M1031_d N_A_298_294#_M1031_g N_VGND_M1037_d VNB NLOWVT
+ L=0.15 W=0.74 AD=0.2109 AS=0.197089 PD=2.05 PS=1.71603 NRD=0 NRS=12.156 M=1
+ R=4.93333 SA=75000.5 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1028 A_536_81# N_RESET_B_M1028_g N_VGND_M1028_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1281 PD=0.66 PS=1.45 NRD=18.564 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1015 N_A_614_81#_M1015_d N_A_334_119#_M1015_g A_536_81# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1281 AS=0.0504 PD=1.45 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_A_298_294#_M1006_d N_A_728_331#_M1006_g N_A_70_74#_M1006_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1456 PD=0.7 PS=1.63 NRD=0 NRS=25.704 M=1 R=2.8
+ SA=75000.3 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1032 N_A_614_81#_M1032_d N_A_818_418#_M1032_g N_A_298_294#_M1006_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.2184 AS=0.0588 PD=1.88 PS=0.7 NRD=71.424 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75000.4 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_A_728_331#_M1029_g N_A_818_418#_M1029_s VNB NLOWVT
+ L=0.15 W=0.74 AD=0.3983 AS=0.1998 PD=2.005 PS=2.02 NRD=78.36 NRS=0 M=1
+ R=4.93333 SA=75000.2 SB=75001.3 A=0.111 P=1.78 MULT=1
MM1007 N_A_728_331#_M1007_d N_CLK_M1007_g N_VGND_M1029_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.3983 PD=2.05 PS=2.005 NRD=0 NRS=78.36 M=1 R=4.93333
+ SA=75001.3 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1017 N_A_1586_149#_M1017_d N_A_728_331#_M1017_g N_A_1499_149#_M1017_s VNB
+ NLOWVT L=0.15 W=0.42 AD=0.0783879 AS=0.1197 PD=0.771207 PS=1.41 NRD=5.712
+ NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1025 N_A_334_119#_M1025_d N_A_818_418#_M1025_g N_A_1586_149#_M1017_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.31255 AS=0.138112 PD=2.62 PS=1.35879 NRD=59.568
+ NRS=4.044 M=1 R=4.93333 SA=75000.5 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1008 N_VGND_M1008_d N_A_1800_291#_M1008_g N_A_1499_149#_M1008_s VNB NLOWVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1155 PD=0.7 PS=1.39 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1021 A_1974_74# N_RESET_B_M1021_g N_VGND_M1008_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1018 N_A_1800_291#_M1018_d N_A_1586_149#_M1018_g A_1974_74# VNB NLOWVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_1586_149#_M1010_g N_Q_N_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75001 A=0.111 P=1.78 MULT=1
MM1033 N_VGND_M1033_d N_A_1586_149#_M1033_g N_Q_N_M1010_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.124942 AS=0.1036 PD=1.14217 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1022 N_A_2366_352#_M1022_d N_A_1586_149#_M1022_g N_VGND_M1033_d VNB NLOWVT
+ L=0.15 W=0.64 AD=0.1728 AS=0.108058 PD=1.82 PS=0.987826 NRD=0 NRS=7.488 M=1
+ R=4.26667 SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1001 N_Q_M1001_d N_A_2366_352#_M1001_g N_VGND_M1001_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1998 PD=1.02 PS=2.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1016 N_Q_M1001_d N_A_2366_352#_M1016_g N_VGND_M1016_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1998 PD=1.02 PS=2.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1036 N_A_70_74#_M1036_d N_D_M1036_g N_VPWR_M1036_s VPB PSHORT L=0.18 W=0.42
+ AD=0.0567 AS=0.1386 PD=0.69 PS=1.5 NRD=0 NRS=21.0987 M=1 R=2.33333 SA=90000.2
+ SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1004 N_VPWR_M1004_d N_RESET_B_M1004_g N_A_70_74#_M1036_d VPB PSHORT L=0.18
+ W=0.42 AD=0.221875 AS=0.0567 PD=1.57944 PS=0.69 NRD=221.98 NRS=0 M=1 R=2.33333
+ SA=90000.7 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1023 N_A_334_119#_M1023_d N_A_298_294#_M1023_g N_VPWR_M1004_d VPB PSHORT
+ L=0.18 W=1 AD=0.28 AS=0.528275 PD=2.56 PS=3.76056 NRD=0 NRS=93.2204 M=1
+ R=5.55556 SA=90000.8 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1011_d N_RESET_B_M1011_g N_A_298_294#_M1011_s VPB PSHORT L=0.18
+ W=0.42 AD=0.135175 AS=0.1113 PD=1.09 PS=1.37 NRD=107.877 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90002.2 A=0.0756 P=1.2 MULT=1
MM1013 A_686_485# N_A_334_119#_M1013_g N_VPWR_M1011_d VPB PSHORT L=0.18 W=0.42
+ AD=0.0441 AS=0.135175 PD=0.63 PS=1.09 NRD=23.443 NRS=39.8531 M=1 R=2.33333
+ SA=90000.9 SB=90001.4 A=0.0756 P=1.2 MULT=1
MM1024 N_A_298_294#_M1024_d N_A_728_331#_M1024_g A_686_485# VPB PSHORT L=0.18
+ W=0.42 AD=0.0567 AS=0.0441 PD=0.69 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.33333
+ SA=90001.3 SB=90001 A=0.0756 P=1.2 MULT=1
MM1026 N_A_70_74#_M1026_d N_A_818_418#_M1026_g N_A_298_294#_M1024_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.273 AS=0.0567 PD=2.14 PS=0.69 NRD=21.0987 NRS=0 M=1
+ R=2.33333 SA=90001.8 SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1034 N_VPWR_M1034_d N_A_728_331#_M1034_g N_A_818_418#_M1034_s VPB PSHORT
+ L=0.18 W=1.12 AD=0.355425 AS=0.3136 PD=1.775 PS=2.8 NRD=29.8849 NRS=0 M=1
+ R=6.22222 SA=90000.2 SB=90001 A=0.2016 P=2.6 MULT=1
MM1009 N_A_728_331#_M1009_d N_CLK_M1009_g N_VPWR_M1034_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3136 AS=0.355425 PD=2.8 PS=1.775 NRD=0 NRS=29.8849 M=1 R=6.22222
+ SA=90001 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1027 N_A_1586_149#_M1027_d N_A_728_331#_M1027_g N_A_334_119#_M1027_s VPB
+ PSHORT L=0.18 W=1 AD=0.25 AS=0.265 PD=2.11268 PS=2.53 NRD=44.3053 NRS=0 M=1
+ R=5.55556 SA=90000.2 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1005 A_1758_389# N_A_818_418#_M1005_g N_A_1586_149#_M1027_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.105 PD=0.66 PS=0.887324 NRD=30.4759 NRS=0 M=1 R=2.33333
+ SA=90000.9 SB=90003.3 A=0.0756 P=1.2 MULT=1
MM1014 N_VPWR_M1014_d N_A_1800_291#_M1014_g A_1758_389# VPB PSHORT L=0.18 W=0.42
+ AD=0.1363 AS=0.0504 PD=1.125 PS=0.66 NRD=126.415 NRS=30.4759 M=1 R=2.33333
+ SA=90001.3 SB=90002.9 A=0.0756 P=1.2 MULT=1
MM1002 N_A_1800_291#_M1002_d N_RESET_B_M1002_g N_VPWR_M1014_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0567 AS=0.1363 PD=0.69 PS=1.125 NRD=0 NRS=126.415 M=1 R=2.33333
+ SA=90001.9 SB=90002.3 A=0.0756 P=1.2 MULT=1
MM1019 N_VPWR_M1019_d N_A_1586_149#_M1019_g N_A_1800_291#_M1002_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.0926045 AS=0.0567 PD=0.804545 PS=0.69 NRD=39.8531 NRS=0 M=1
+ R=2.33333 SA=90002.4 SB=90001.8 A=0.0756 P=1.2 MULT=1
MM1030 N_Q_N_M1030_d N_A_1586_149#_M1030_g N_VPWR_M1019_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.246945 PD=1.39 PS=2.14545 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.2 SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1035 N_Q_N_M1030_d N_A_1586_149#_M1035_g N_VPWR_M1035_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.205298 PD=1.39 PS=1.55849 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.7 SB=90000.8 A=0.2016 P=2.6 MULT=1
MM1020 N_A_2366_352#_M1020_d N_A_1586_149#_M1020_g N_VPWR_M1035_s VPB PSHORT
+ L=0.18 W=1 AD=0.375 AS=0.183302 PD=2.75 PS=1.39151 NRD=17.73 NRS=16.0752 M=1
+ R=5.55556 SA=90002.3 SB=90000.3 A=0.18 P=2.36 MULT=1
MM1000 N_Q_M1000_d N_A_2366_352#_M1000_g N_VPWR_M1000_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.2
+ SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1003 N_Q_M1000_d N_A_2366_352#_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.7
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX38_noxref VNB VPB NWDIODE A=24.9576 P=33.65
c_153 VNB 0 7.64129e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_ms__dfrbp_2.pxi.spice"
*
.ends
*
*

* File: sky130_fd_sc_ms__or2b_1.pxi.spice
* Created: Wed Sep  2 12:27:51 2020
* 
x_PM_SKY130_FD_SC_MS__OR2B_1%B_N N_B_N_c_60_n N_B_N_M1005_g N_B_N_c_61_n
+ N_B_N_c_62_n N_B_N_M1003_g B_N PM_SKY130_FD_SC_MS__OR2B_1%B_N
x_PM_SKY130_FD_SC_MS__OR2B_1%A_27_112# N_A_27_112#_M1003_s N_A_27_112#_M1005_s
+ N_A_27_112#_M1000_g N_A_27_112#_M1004_g N_A_27_112#_c_94_n N_A_27_112#_c_95_n
+ N_A_27_112#_c_101_n N_A_27_112#_c_102_n N_A_27_112#_c_103_n
+ N_A_27_112#_c_115_n N_A_27_112#_c_96_n N_A_27_112#_c_97_n N_A_27_112#_c_98_n
+ N_A_27_112#_c_99_n PM_SKY130_FD_SC_MS__OR2B_1%A_27_112#
x_PM_SKY130_FD_SC_MS__OR2B_1%A N_A_M1001_g N_A_M1006_g A N_A_c_160_n N_A_c_161_n
+ PM_SKY130_FD_SC_MS__OR2B_1%A
x_PM_SKY130_FD_SC_MS__OR2B_1%A_264_368# N_A_264_368#_M1000_d
+ N_A_264_368#_M1004_s N_A_264_368#_M1002_g N_A_264_368#_M1007_g
+ N_A_264_368#_c_202_n N_A_264_368#_c_196_n N_A_264_368#_c_197_n
+ N_A_264_368#_c_198_n N_A_264_368#_c_204_n N_A_264_368#_c_199_n
+ N_A_264_368#_c_200_n PM_SKY130_FD_SC_MS__OR2B_1%A_264_368#
x_PM_SKY130_FD_SC_MS__OR2B_1%VPWR N_VPWR_M1005_d N_VPWR_M1006_d N_VPWR_c_265_n
+ N_VPWR_c_266_n N_VPWR_c_267_n N_VPWR_c_268_n VPWR N_VPWR_c_269_n
+ N_VPWR_c_270_n N_VPWR_c_264_n N_VPWR_c_272_n PM_SKY130_FD_SC_MS__OR2B_1%VPWR
x_PM_SKY130_FD_SC_MS__OR2B_1%X N_X_M1007_d N_X_M1002_d N_X_c_302_n N_X_c_303_n X
+ X X N_X_c_306_n N_X_c_304_n X PM_SKY130_FD_SC_MS__OR2B_1%X
x_PM_SKY130_FD_SC_MS__OR2B_1%VGND N_VGND_M1003_d N_VGND_M1001_d N_VGND_c_327_n
+ N_VGND_c_328_n N_VGND_c_329_n N_VGND_c_330_n VGND N_VGND_c_331_n
+ N_VGND_c_332_n N_VGND_c_333_n N_VGND_c_334_n PM_SKY130_FD_SC_MS__OR2B_1%VGND
cc_1 VNB N_B_N_c_60_n 0.0695094f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.7
cc_2 VNB N_B_N_c_61_n 0.02624f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.295
cc_3 VNB N_B_N_c_62_n 0.0243562f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=1.22
cc_4 VNB B_N 0.00771224f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_5 VNB N_A_27_112#_M1000_g 0.0236728f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=0.835
cc_6 VNB N_A_27_112#_M1004_g 0.00228213f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.385
cc_7 VNB N_A_27_112#_c_94_n 0.0441328f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.385
cc_8 VNB N_A_27_112#_c_95_n 0.0114296f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_9 VNB N_A_27_112#_c_96_n 0.00279704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_112#_c_97_n 0.00409161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_112#_c_98_n 0.0155571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_112#_c_99_n 0.0144242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_M1001_g 0.0263428f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.54
cc_14 VNB N_A_c_160_n 0.0281456f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.295
cc_15 VNB N_A_c_161_n 0.00180753f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.385
cc_16 VNB N_A_264_368#_M1002_g 0.00179278f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=0.835
cc_17 VNB N_A_264_368#_M1007_g 0.0294109f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.385
cc_18 VNB N_A_264_368#_c_196_n 0.00325419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_264_368#_c_197_n 0.00335286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_264_368#_c_198_n 0.0202157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_264_368#_c_199_n 0.00626634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_264_368#_c_200_n 0.0345886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_264_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_X_c_302_n 0.0272846f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=0.835
cc_25 VNB N_X_c_303_n 0.0154926f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.385
cc_26 VNB N_X_c_304_n 0.0248898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_327_n 0.0346814f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=0.835
cc_28 VNB N_VGND_c_328_n 0.0188865f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.385
cc_29 VNB N_VGND_c_329_n 0.0216143f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_30 VNB N_VGND_c_330_n 0.00798243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_331_n 0.0310594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_332_n 0.0206731f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_333_n 0.220663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_334_n 0.0100982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VPB N_B_N_c_60_n 0.00355203f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=1.7
cc_36 VPB N_B_N_M1005_g 0.053045f $X=-0.19 $Y=1.66 $X2=0.505 $Y2=2.54
cc_37 VPB N_A_27_112#_M1004_g 0.0275937f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.385
cc_38 VPB N_A_27_112#_c_101_n 0.0431698f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_39 VPB N_A_27_112#_c_102_n 0.00235784f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_40 VPB N_A_27_112#_c_103_n 0.00979329f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_41 VPB N_A_27_112#_c_97_n 0.0104101f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_42 VPB N_A_M1006_g 0.0217955f $X=-0.19 $Y=1.66 $X2=0.88 $Y2=1.22
cc_43 VPB N_A_c_160_n 0.00613741f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.295
cc_44 VPB N_A_c_161_n 0.00425926f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.385
cc_45 VPB N_A_264_368#_M1002_g 0.0304781f $X=-0.19 $Y=1.66 $X2=0.88 $Y2=0.835
cc_46 VPB N_A_264_368#_c_202_n 0.0174287f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_47 VPB N_A_264_368#_c_197_n 0.00133625f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_48 VPB N_A_264_368#_c_204_n 0.00674445f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_265_n 0.0268834f $X=-0.19 $Y=1.66 $X2=0.88 $Y2=0.835
cc_50 VPB N_VPWR_c_266_n 0.0142501f $X=-0.19 $Y=1.66 $X2=0.36 $Y2=1.385
cc_51 VPB N_VPWR_c_267_n 0.0395991f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_268_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.385
cc_53 VPB N_VPWR_c_269_n 0.0191515f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_270_n 0.0227588f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_264_n 0.0880701f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_272_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_57 VPB X 0.0466392f $X=-0.19 $Y=1.66 $X2=0.29 $Y2=1.385
cc_58 VPB N_X_c_306_n 0.020212f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_59 VPB N_X_c_304_n 0.00790712f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_60 N_B_N_c_62_n N_A_27_112#_M1000_g 0.00726223f $X=0.88 $Y=1.22 $X2=0 $Y2=0
cc_61 N_B_N_c_60_n N_A_27_112#_c_94_n 0.00307942f $X=0.505 $Y=1.7 $X2=0 $Y2=0
cc_62 N_B_N_c_61_n N_A_27_112#_c_94_n 0.00389289f $X=0.805 $Y=1.295 $X2=0 $Y2=0
cc_63 N_B_N_M1005_g N_A_27_112#_c_101_n 0.0254932f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_64 N_B_N_M1005_g N_A_27_112#_c_102_n 0.0167703f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_65 N_B_N_c_61_n N_A_27_112#_c_102_n 0.0019038f $X=0.805 $Y=1.295 $X2=0 $Y2=0
cc_66 B_N N_A_27_112#_c_102_n 5.214e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_67 N_B_N_c_60_n N_A_27_112#_c_103_n 0.00222782f $X=0.505 $Y=1.7 $X2=0 $Y2=0
cc_68 N_B_N_M1005_g N_A_27_112#_c_103_n 0.00438675f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_69 B_N N_A_27_112#_c_103_n 0.0230941f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_70 N_B_N_c_62_n N_A_27_112#_c_115_n 0.00400158f $X=0.88 $Y=1.22 $X2=0 $Y2=0
cc_71 N_B_N_c_61_n N_A_27_112#_c_96_n 0.00871279f $X=0.805 $Y=1.295 $X2=0 $Y2=0
cc_72 N_B_N_c_62_n N_A_27_112#_c_96_n 0.00795326f $X=0.88 $Y=1.22 $X2=0 $Y2=0
cc_73 B_N N_A_27_112#_c_96_n 0.0237254f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_74 N_B_N_c_60_n N_A_27_112#_c_97_n 0.00954145f $X=0.505 $Y=1.7 $X2=0 $Y2=0
cc_75 N_B_N_M1005_g N_A_27_112#_c_97_n 0.00138205f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_76 N_B_N_c_61_n N_A_27_112#_c_97_n 0.00620548f $X=0.805 $Y=1.295 $X2=0 $Y2=0
cc_77 N_B_N_c_61_n N_A_27_112#_c_98_n 0.0101512f $X=0.805 $Y=1.295 $X2=0 $Y2=0
cc_78 N_B_N_c_60_n N_A_27_112#_c_99_n 0.0102304f $X=0.505 $Y=1.7 $X2=0 $Y2=0
cc_79 B_N N_A_27_112#_c_99_n 0.0271897f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_80 N_B_N_M1005_g N_VPWR_c_265_n 0.00914782f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_81 N_B_N_M1005_g N_VPWR_c_269_n 0.005209f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_82 N_B_N_M1005_g N_VPWR_c_264_n 0.00990469f $X=0.505 $Y=2.54 $X2=0 $Y2=0
cc_83 N_B_N_c_62_n N_VGND_c_327_n 0.0059966f $X=0.88 $Y=1.22 $X2=0 $Y2=0
cc_84 N_B_N_c_62_n N_VGND_c_331_n 0.00434478f $X=0.88 $Y=1.22 $X2=0 $Y2=0
cc_85 N_B_N_c_62_n N_VGND_c_333_n 0.00487769f $X=0.88 $Y=1.22 $X2=0 $Y2=0
cc_86 N_A_27_112#_M1000_g N_A_M1001_g 0.014193f $X=1.665 $Y=0.835 $X2=0 $Y2=0
cc_87 N_A_27_112#_M1004_g N_A_M1006_g 0.0383809f $X=1.69 $Y=2.34 $X2=0 $Y2=0
cc_88 N_A_27_112#_c_95_n N_A_c_160_n 0.052574f $X=1.59 $Y=1.3 $X2=0 $Y2=0
cc_89 N_A_27_112#_c_95_n N_A_c_161_n 4.43468e-19 $X=1.59 $Y=1.3 $X2=0 $Y2=0
cc_90 N_A_27_112#_M1004_g N_A_264_368#_c_202_n 0.0180607f $X=1.69 $Y=2.34 $X2=0
+ $Y2=0
cc_91 N_A_27_112#_M1000_g N_A_264_368#_c_196_n 0.00744356f $X=1.665 $Y=0.835
+ $X2=0 $Y2=0
cc_92 N_A_27_112#_M1000_g N_A_264_368#_c_197_n 0.00575302f $X=1.665 $Y=0.835
+ $X2=0 $Y2=0
cc_93 N_A_27_112#_M1004_g N_A_264_368#_c_197_n 0.00977134f $X=1.69 $Y=2.34 $X2=0
+ $Y2=0
cc_94 N_A_27_112#_c_95_n N_A_264_368#_c_197_n 0.00933029f $X=1.59 $Y=1.3 $X2=0
+ $Y2=0
cc_95 N_A_27_112#_c_98_n N_A_264_368#_c_197_n 0.0250314f $X=1.36 $Y=1.465 $X2=0
+ $Y2=0
cc_96 N_A_27_112#_M1004_g N_A_264_368#_c_204_n 0.0152622f $X=1.69 $Y=2.34 $X2=0
+ $Y2=0
cc_97 N_A_27_112#_c_94_n N_A_264_368#_c_204_n 0.00775559f $X=1.59 $Y=1.465 $X2=0
+ $Y2=0
cc_98 N_A_27_112#_c_97_n N_A_264_368#_c_204_n 0.00447704f $X=0.83 $Y=1.465 $X2=0
+ $Y2=0
cc_99 N_A_27_112#_c_98_n N_A_264_368#_c_204_n 0.0155529f $X=1.36 $Y=1.465 $X2=0
+ $Y2=0
cc_100 N_A_27_112#_M1000_g N_A_264_368#_c_199_n 0.0056446f $X=1.665 $Y=0.835
+ $X2=0 $Y2=0
cc_101 N_A_27_112#_M1004_g N_VPWR_c_265_n 0.00417133f $X=1.69 $Y=2.34 $X2=0
+ $Y2=0
cc_102 N_A_27_112#_c_101_n N_VPWR_c_265_n 0.0346006f $X=0.28 $Y=2.265 $X2=0
+ $Y2=0
cc_103 N_A_27_112#_c_102_n N_VPWR_c_265_n 0.00371626f $X=0.66 $Y=1.845 $X2=0
+ $Y2=0
cc_104 N_A_27_112#_c_97_n N_VPWR_c_265_n 0.0157412f $X=0.83 $Y=1.465 $X2=0 $Y2=0
cc_105 N_A_27_112#_c_98_n N_VPWR_c_265_n 0.00497979f $X=1.36 $Y=1.465 $X2=0
+ $Y2=0
cc_106 N_A_27_112#_M1004_g N_VPWR_c_267_n 0.00567889f $X=1.69 $Y=2.34 $X2=0
+ $Y2=0
cc_107 N_A_27_112#_c_101_n N_VPWR_c_269_n 0.014549f $X=0.28 $Y=2.265 $X2=0 $Y2=0
cc_108 N_A_27_112#_M1004_g N_VPWR_c_264_n 0.00610055f $X=1.69 $Y=2.34 $X2=0
+ $Y2=0
cc_109 N_A_27_112#_c_101_n N_VPWR_c_264_n 0.0119743f $X=0.28 $Y=2.265 $X2=0
+ $Y2=0
cc_110 N_A_27_112#_M1000_g N_VGND_c_327_n 0.00735506f $X=1.665 $Y=0.835 $X2=0
+ $Y2=0
cc_111 N_A_27_112#_c_94_n N_VGND_c_327_n 0.00766427f $X=1.59 $Y=1.465 $X2=0
+ $Y2=0
cc_112 N_A_27_112#_c_96_n N_VGND_c_327_n 0.00488088f $X=0.745 $Y=1.3 $X2=0 $Y2=0
cc_113 N_A_27_112#_c_98_n N_VGND_c_327_n 0.0449072f $X=1.36 $Y=1.465 $X2=0 $Y2=0
cc_114 N_A_27_112#_M1000_g N_VGND_c_329_n 0.00418801f $X=1.665 $Y=0.835 $X2=0
+ $Y2=0
cc_115 N_A_27_112#_c_115_n N_VGND_c_331_n 0.00243801f $X=0.745 $Y=1.01 $X2=0
+ $Y2=0
cc_116 N_A_27_112#_c_99_n N_VGND_c_331_n 0.00905393f $X=0.665 $Y=0.845 $X2=0
+ $Y2=0
cc_117 N_A_27_112#_M1000_g N_VGND_c_333_n 0.00487769f $X=1.665 $Y=0.835 $X2=0
+ $Y2=0
cc_118 N_A_27_112#_c_115_n N_VGND_c_333_n 0.00494557f $X=0.745 $Y=1.01 $X2=0
+ $Y2=0
cc_119 N_A_27_112#_c_99_n N_VGND_c_333_n 0.0154532f $X=0.665 $Y=0.845 $X2=0
+ $Y2=0
cc_120 N_A_M1006_g N_A_264_368#_M1002_g 0.0182493f $X=2.11 $Y=2.34 $X2=0 $Y2=0
cc_121 N_A_c_161_n N_A_264_368#_M1002_g 0.0026215f $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_122 N_A_M1001_g N_A_264_368#_M1007_g 0.0127273f $X=2.095 $Y=0.835 $X2=0 $Y2=0
cc_123 N_A_M1006_g N_A_264_368#_c_202_n 0.00255838f $X=2.11 $Y=2.34 $X2=0 $Y2=0
cc_124 N_A_M1001_g N_A_264_368#_c_196_n 0.0124806f $X=2.095 $Y=0.835 $X2=0 $Y2=0
cc_125 N_A_M1001_g N_A_264_368#_c_197_n 0.00519192f $X=2.095 $Y=0.835 $X2=0
+ $Y2=0
cc_126 N_A_c_161_n N_A_264_368#_c_197_n 0.0322792f $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_127 N_A_M1001_g N_A_264_368#_c_198_n 0.013594f $X=2.095 $Y=0.835 $X2=0 $Y2=0
cc_128 N_A_c_160_n N_A_264_368#_c_198_n 0.00309695f $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_129 N_A_c_161_n N_A_264_368#_c_198_n 0.0466983f $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_130 N_A_M1006_g N_A_264_368#_c_204_n 0.00377011f $X=2.11 $Y=2.34 $X2=0 $Y2=0
cc_131 N_A_M1001_g N_A_264_368#_c_199_n 0.00308855f $X=2.095 $Y=0.835 $X2=0
+ $Y2=0
cc_132 N_A_c_161_n N_A_264_368#_c_199_n 7.33087e-19 $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_133 N_A_M1001_g N_A_264_368#_c_200_n 0.00113203f $X=2.095 $Y=0.835 $X2=0
+ $Y2=0
cc_134 N_A_c_160_n N_A_264_368#_c_200_n 0.0176113f $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_135 N_A_c_161_n N_A_264_368#_c_200_n 3.09225e-19 $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_136 N_A_M1006_g N_VPWR_c_266_n 0.00884557f $X=2.11 $Y=2.34 $X2=0 $Y2=0
cc_137 N_A_c_160_n N_VPWR_c_266_n 6.61748e-19 $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_138 N_A_c_161_n N_VPWR_c_266_n 0.00954634f $X=2.2 $Y=1.515 $X2=0 $Y2=0
cc_139 N_A_M1006_g N_VPWR_c_267_n 0.0059286f $X=2.11 $Y=2.34 $X2=0 $Y2=0
cc_140 N_A_M1006_g N_VPWR_c_264_n 0.00610055f $X=2.11 $Y=2.34 $X2=0 $Y2=0
cc_141 N_A_M1006_g N_X_c_306_n 7.79105e-19 $X=2.11 $Y=2.34 $X2=0 $Y2=0
cc_142 N_A_M1001_g N_VGND_c_328_n 0.00665253f $X=2.095 $Y=0.835 $X2=0 $Y2=0
cc_143 N_A_M1001_g N_VGND_c_329_n 0.0043356f $X=2.095 $Y=0.835 $X2=0 $Y2=0
cc_144 N_A_M1001_g N_VGND_c_333_n 0.00487769f $X=2.095 $Y=0.835 $X2=0 $Y2=0
cc_145 N_A_264_368#_c_202_n N_VPWR_c_265_n 0.038037f $X=1.465 $Y=2.695 $X2=0
+ $Y2=0
cc_146 N_A_264_368#_M1002_g N_VPWR_c_266_n 0.00520277f $X=2.695 $Y=2.4 $X2=0
+ $Y2=0
cc_147 N_A_264_368#_c_202_n N_VPWR_c_266_n 0.0113776f $X=1.465 $Y=2.695 $X2=0
+ $Y2=0
cc_148 N_A_264_368#_c_198_n N_VPWR_c_266_n 0.00182168f $X=2.535 $Y=1.095 $X2=0
+ $Y2=0
cc_149 N_A_264_368#_c_202_n N_VPWR_c_267_n 0.00975961f $X=1.465 $Y=2.695 $X2=0
+ $Y2=0
cc_150 N_A_264_368#_M1002_g N_VPWR_c_270_n 0.005209f $X=2.695 $Y=2.4 $X2=0 $Y2=0
cc_151 N_A_264_368#_M1002_g N_VPWR_c_264_n 0.0099091f $X=2.695 $Y=2.4 $X2=0
+ $Y2=0
cc_152 N_A_264_368#_c_202_n N_VPWR_c_264_n 0.0111753f $X=1.465 $Y=2.695 $X2=0
+ $Y2=0
cc_153 N_A_264_368#_c_204_n A_356_368# 0.00300467f $X=1.78 $Y=1.905 $X2=-0.19
+ $Y2=-0.245
cc_154 N_A_264_368#_M1007_g N_X_c_302_n 0.0113949f $X=2.825 $Y=0.74 $X2=0 $Y2=0
cc_155 N_A_264_368#_M1007_g N_X_c_303_n 0.00556841f $X=2.825 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A_264_368#_c_198_n N_X_c_303_n 0.0104368f $X=2.535 $Y=1.095 $X2=0 $Y2=0
cc_157 N_A_264_368#_c_200_n N_X_c_303_n 2.77016e-19 $X=2.77 $Y=1.465 $X2=0 $Y2=0
cc_158 N_A_264_368#_M1002_g X 0.0120848f $X=2.695 $Y=2.4 $X2=0 $Y2=0
cc_159 N_A_264_368#_M1002_g N_X_c_306_n 0.00523005f $X=2.695 $Y=2.4 $X2=0 $Y2=0
cc_160 N_A_264_368#_c_198_n N_X_c_306_n 0.0138127f $X=2.535 $Y=1.095 $X2=0 $Y2=0
cc_161 N_A_264_368#_c_200_n N_X_c_306_n 0.00116022f $X=2.77 $Y=1.465 $X2=0 $Y2=0
cc_162 N_A_264_368#_M1002_g N_X_c_304_n 0.00415514f $X=2.695 $Y=2.4 $X2=0 $Y2=0
cc_163 N_A_264_368#_M1007_g N_X_c_304_n 0.00246301f $X=2.825 $Y=0.74 $X2=0 $Y2=0
cc_164 N_A_264_368#_c_198_n N_X_c_304_n 0.0302873f $X=2.535 $Y=1.095 $X2=0 $Y2=0
cc_165 N_A_264_368#_c_200_n N_X_c_304_n 0.00232633f $X=2.77 $Y=1.465 $X2=0 $Y2=0
cc_166 N_A_264_368#_c_198_n N_VGND_M1001_d 0.00843341f $X=2.535 $Y=1.095 $X2=0
+ $Y2=0
cc_167 N_A_264_368#_c_196_n N_VGND_c_327_n 0.0379888f $X=1.88 $Y=0.835 $X2=0
+ $Y2=0
cc_168 N_A_264_368#_c_199_n N_VGND_c_327_n 0.0102677f $X=1.87 $Y=1.095 $X2=0
+ $Y2=0
cc_169 N_A_264_368#_M1007_g N_VGND_c_328_n 0.0110504f $X=2.825 $Y=0.74 $X2=0
+ $Y2=0
cc_170 N_A_264_368#_c_196_n N_VGND_c_328_n 0.0195637f $X=1.88 $Y=0.835 $X2=0
+ $Y2=0
cc_171 N_A_264_368#_c_198_n N_VGND_c_328_n 0.0347439f $X=2.535 $Y=1.095 $X2=0
+ $Y2=0
cc_172 N_A_264_368#_c_200_n N_VGND_c_328_n 3.0856e-19 $X=2.77 $Y=1.465 $X2=0
+ $Y2=0
cc_173 N_A_264_368#_c_196_n N_VGND_c_329_n 0.00852231f $X=1.88 $Y=0.835 $X2=0
+ $Y2=0
cc_174 N_A_264_368#_M1007_g N_VGND_c_332_n 0.00434272f $X=2.825 $Y=0.74 $X2=0
+ $Y2=0
cc_175 N_A_264_368#_M1007_g N_VGND_c_333_n 0.00829406f $X=2.825 $Y=0.74 $X2=0
+ $Y2=0
cc_176 N_A_264_368#_c_196_n N_VGND_c_333_n 0.0112256f $X=1.88 $Y=0.835 $X2=0
+ $Y2=0
cc_177 N_VPWR_c_270_n X 0.0230269f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_178 N_VPWR_c_264_n X 0.0189916f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_179 N_VPWR_c_266_n N_X_c_306_n 0.0421814f $X=2.42 $Y=2.115 $X2=0 $Y2=0
cc_180 N_X_c_302_n N_VGND_c_328_n 0.0353629f $X=3.04 $Y=0.515 $X2=0 $Y2=0
cc_181 N_X_c_302_n N_VGND_c_332_n 0.0176874f $X=3.04 $Y=0.515 $X2=0 $Y2=0
cc_182 N_X_c_302_n N_VGND_c_333_n 0.0145837f $X=3.04 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__dfstp_1.pxi.spice
* Created: Wed Sep  2 12:03:36 2020
* 
x_PM_SKY130_FD_SC_MS__DFSTP_1%D N_D_c_239_n N_D_M1008_g N_D_M1028_g D D
+ N_D_c_241_n N_D_c_242_n N_D_c_246_n PM_SKY130_FD_SC_MS__DFSTP_1%D
x_PM_SKY130_FD_SC_MS__DFSTP_1%CLK N_CLK_M1004_g N_CLK_M1031_g CLK N_CLK_c_275_n
+ N_CLK_c_276_n PM_SKY130_FD_SC_MS__DFSTP_1%CLK
x_PM_SKY130_FD_SC_MS__DFSTP_1%A_398_74# N_A_398_74#_M1020_d N_A_398_74#_M1010_d
+ N_A_398_74#_M1017_g N_A_398_74#_c_311_n N_A_398_74#_c_312_n
+ N_A_398_74#_M1024_g N_A_398_74#_M1007_g N_A_398_74#_M1027_g
+ N_A_398_74#_c_333_n N_A_398_74#_c_314_n N_A_398_74#_c_334_n
+ N_A_398_74#_c_315_n N_A_398_74#_c_316_n N_A_398_74#_c_335_n
+ N_A_398_74#_c_336_n N_A_398_74#_c_317_n N_A_398_74#_c_337_n
+ N_A_398_74#_c_338_n N_A_398_74#_c_318_n N_A_398_74#_c_340_n
+ N_A_398_74#_c_341_n N_A_398_74#_c_342_n N_A_398_74#_c_343_n
+ N_A_398_74#_c_344_n N_A_398_74#_c_345_n N_A_398_74#_c_377_p
+ N_A_398_74#_c_419_p N_A_398_74#_c_378_p N_A_398_74#_c_346_n
+ N_A_398_74#_c_380_p N_A_398_74#_c_319_n N_A_398_74#_c_320_n
+ N_A_398_74#_c_321_n N_A_398_74#_c_322_n N_A_398_74#_c_323_n
+ N_A_398_74#_c_349_n N_A_398_74#_c_324_n N_A_398_74#_c_325_n
+ N_A_398_74#_c_326_n N_A_398_74#_c_350_n N_A_398_74#_c_327_n
+ N_A_398_74#_c_328_n N_A_398_74#_c_352_n PM_SKY130_FD_SC_MS__DFSTP_1%A_398_74#
x_PM_SKY130_FD_SC_MS__DFSTP_1%A_760_395# N_A_760_395#_M1011_s
+ N_A_760_395#_M1000_d N_A_760_395#_M1030_g N_A_760_395#_c_590_n
+ N_A_760_395#_M1022_g N_A_760_395#_c_591_n N_A_760_395#_c_596_n
+ N_A_760_395#_c_597_n N_A_760_395#_c_598_n N_A_760_395#_c_592_n
+ N_A_760_395#_c_599_n N_A_760_395#_c_600_n N_A_760_395#_c_593_n
+ PM_SKY130_FD_SC_MS__DFSTP_1%A_760_395#
x_PM_SKY130_FD_SC_MS__DFSTP_1%A_604_74# N_A_604_74#_M1013_d N_A_604_74#_M1017_d
+ N_A_604_74#_M1000_g N_A_604_74#_M1011_g N_A_604_74#_M1001_g
+ N_A_604_74#_M1003_g N_A_604_74#_c_672_n N_A_604_74#_c_673_n
+ N_A_604_74#_c_674_n N_A_604_74#_c_675_n N_A_604_74#_c_676_n
+ N_A_604_74#_c_677_n N_A_604_74#_c_678_n N_A_604_74#_c_679_n
+ N_A_604_74#_c_688_n N_A_604_74#_c_680_n N_A_604_74#_c_681_n
+ N_A_604_74#_c_682_n PM_SKY130_FD_SC_MS__DFSTP_1%A_604_74#
x_PM_SKY130_FD_SC_MS__DFSTP_1%SET_B N_SET_B_M1012_g N_SET_B_M1009_g
+ N_SET_B_c_813_n N_SET_B_M1023_g N_SET_B_c_819_n N_SET_B_M1006_g
+ N_SET_B_c_814_n N_SET_B_c_815_n N_SET_B_c_822_n N_SET_B_c_823_n
+ N_SET_B_c_824_n SET_B N_SET_B_c_826_n N_SET_B_c_816_n
+ PM_SKY130_FD_SC_MS__DFSTP_1%SET_B
x_PM_SKY130_FD_SC_MS__DFSTP_1%A_224_350# N_A_224_350#_M1031_s
+ N_A_224_350#_M1004_s N_A_224_350#_M1020_g N_A_224_350#_M1010_g
+ N_A_224_350#_c_950_n N_A_224_350#_c_938_n N_A_224_350#_c_951_n
+ N_A_224_350#_c_952_n N_A_224_350#_M1013_g N_A_224_350#_M1015_g
+ N_A_224_350#_c_954_n N_A_224_350#_M1021_g N_A_224_350#_c_940_n
+ N_A_224_350#_c_941_n N_A_224_350#_M1018_g N_A_224_350#_c_943_n
+ N_A_224_350#_c_944_n N_A_224_350#_c_945_n N_A_224_350#_c_961_n
+ N_A_224_350#_c_946_n N_A_224_350#_c_963_n N_A_224_350#_c_947_n
+ N_A_224_350#_c_948_n N_A_224_350#_c_965_n
+ PM_SKY130_FD_SC_MS__DFSTP_1%A_224_350#
x_PM_SKY130_FD_SC_MS__DFSTP_1%A_1470_48# N_A_1470_48#_M1005_d
+ N_A_1470_48#_M1016_d N_A_1470_48#_M1019_g N_A_1470_48#_M1002_g
+ N_A_1470_48#_c_1122_n N_A_1470_48#_c_1123_n N_A_1470_48#_c_1137_n
+ N_A_1470_48#_c_1124_n N_A_1470_48#_c_1125_n N_A_1470_48#_c_1129_n
+ N_A_1470_48#_c_1126_n N_A_1470_48#_c_1127_n
+ PM_SKY130_FD_SC_MS__DFSTP_1%A_1470_48#
x_PM_SKY130_FD_SC_MS__DFSTP_1%A_1301_392# N_A_1301_392#_M1007_d
+ N_A_1301_392#_M1021_d N_A_1301_392#_M1006_d N_A_1301_392#_c_1203_n
+ N_A_1301_392#_M1005_g N_A_1301_392#_M1016_g N_A_1301_392#_c_1213_n
+ N_A_1301_392#_M1026_g N_A_1301_392#_c_1215_n N_A_1301_392#_M1029_g
+ N_A_1301_392#_c_1216_n N_A_1301_392#_c_1217_n N_A_1301_392#_c_1218_n
+ N_A_1301_392#_c_1219_n N_A_1301_392#_c_1220_n N_A_1301_392#_c_1206_n
+ N_A_1301_392#_c_1221_n N_A_1301_392#_c_1222_n N_A_1301_392#_c_1223_n
+ N_A_1301_392#_c_1224_n N_A_1301_392#_c_1225_n N_A_1301_392#_c_1207_n
+ N_A_1301_392#_c_1208_n N_A_1301_392#_c_1226_n N_A_1301_392#_c_1227_n
+ N_A_1301_392#_c_1228_n N_A_1301_392#_c_1209_n N_A_1301_392#_c_1210_n
+ N_A_1301_392#_c_1229_n PM_SKY130_FD_SC_MS__DFSTP_1%A_1301_392#
x_PM_SKY130_FD_SC_MS__DFSTP_1%A_1902_74# N_A_1902_74#_M1026_s
+ N_A_1902_74#_M1029_s N_A_1902_74#_c_1376_n N_A_1902_74#_M1014_g
+ N_A_1902_74#_M1025_g N_A_1902_74#_c_1378_n N_A_1902_74#_c_1379_n
+ N_A_1902_74#_c_1380_n N_A_1902_74#_c_1381_n N_A_1902_74#_c_1382_n
+ N_A_1902_74#_c_1383_n N_A_1902_74#_c_1384_n
+ PM_SKY130_FD_SC_MS__DFSTP_1%A_1902_74#
x_PM_SKY130_FD_SC_MS__DFSTP_1%A_27_74# N_A_27_74#_M1028_s N_A_27_74#_M1013_s
+ N_A_27_74#_M1008_s N_A_27_74#_M1017_s N_A_27_74#_c_1432_n N_A_27_74#_c_1433_n
+ N_A_27_74#_c_1438_n N_A_27_74#_c_1439_n N_A_27_74#_c_1440_n
+ N_A_27_74#_c_1434_n N_A_27_74#_c_1435_n N_A_27_74#_c_1442_n
+ N_A_27_74#_c_1482_n N_A_27_74#_c_1436_n PM_SKY130_FD_SC_MS__DFSTP_1%A_27_74#
x_PM_SKY130_FD_SC_MS__DFSTP_1%VPWR N_VPWR_M1008_d N_VPWR_M1004_d N_VPWR_M1030_d
+ N_VPWR_M1012_d N_VPWR_M1002_d N_VPWR_M1016_s N_VPWR_M1029_d N_VPWR_c_1500_n
+ N_VPWR_c_1501_n N_VPWR_c_1502_n N_VPWR_c_1503_n N_VPWR_c_1504_n
+ N_VPWR_c_1505_n N_VPWR_c_1506_n N_VPWR_c_1507_n N_VPWR_c_1508_n
+ N_VPWR_c_1509_n N_VPWR_c_1510_n VPWR N_VPWR_c_1511_n N_VPWR_c_1512_n
+ N_VPWR_c_1513_n N_VPWR_c_1514_n N_VPWR_c_1515_n N_VPWR_c_1516_n
+ N_VPWR_c_1499_n N_VPWR_c_1518_n N_VPWR_c_1519_n N_VPWR_c_1520_n
+ N_VPWR_c_1521_n N_VPWR_c_1522_n PM_SKY130_FD_SC_MS__DFSTP_1%VPWR
x_PM_SKY130_FD_SC_MS__DFSTP_1%Q N_Q_M1014_d N_Q_M1025_d Q Q Q Q Q Q Q
+ N_Q_c_1638_n PM_SKY130_FD_SC_MS__DFSTP_1%Q
x_PM_SKY130_FD_SC_MS__DFSTP_1%VGND N_VGND_M1028_d N_VGND_M1031_d N_VGND_M1022_d
+ N_VGND_M1009_d N_VGND_M1023_d N_VGND_M1026_d N_VGND_c_1654_n N_VGND_c_1655_n
+ N_VGND_c_1656_n N_VGND_c_1657_n N_VGND_c_1658_n N_VGND_c_1659_n
+ N_VGND_c_1660_n N_VGND_c_1661_n N_VGND_c_1662_n N_VGND_c_1663_n VGND
+ N_VGND_c_1664_n N_VGND_c_1665_n N_VGND_c_1666_n N_VGND_c_1667_n
+ N_VGND_c_1668_n N_VGND_c_1669_n N_VGND_c_1670_n N_VGND_c_1671_n
+ N_VGND_c_1672_n PM_SKY130_FD_SC_MS__DFSTP_1%VGND
cc_1 VNB N_D_c_239_n 0.044776f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.79
cc_2 VNB N_D_M1028_g 0.0283827f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_3 VNB N_D_c_241_n 0.0265904f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_4 VNB N_D_c_242_n 0.00250659f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_5 VNB N_CLK_M1004_g 0.0012514f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.99
cc_6 VNB CLK 0.00935738f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_7 VNB N_CLK_c_275_n 0.0321883f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_8 VNB N_CLK_c_276_n 0.019965f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_398_74#_c_311_n 0.0188524f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_10 VNB N_A_398_74#_c_312_n 0.0141105f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_11 VNB N_A_398_74#_M1024_g 0.0515076f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.145
cc_12 VNB N_A_398_74#_c_314_n 0.00681347f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_13 VNB N_A_398_74#_c_315_n 0.0128874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_398_74#_c_316_n 0.00283335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_398_74#_c_317_n 8.85608e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_398_74#_c_318_n 7.34628e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_398_74#_c_319_n 0.00119326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_398_74#_c_320_n 0.00560214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_398_74#_c_321_n 0.00222263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_398_74#_c_322_n 0.015306f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_398_74#_c_323_n 0.00662299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_398_74#_c_324_n 0.00615999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_398_74#_c_325_n 0.0308207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_398_74#_c_326_n 0.00183869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_398_74#_c_327_n 0.0131519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_398_74#_c_328_n 0.0180562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_760_395#_c_590_n 0.0194532f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_28 VNB N_A_760_395#_c_591_n 0.0193805f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.145
cc_29 VNB N_A_760_395#_c_592_n 0.0182397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_760_395#_c_593_n 0.0560041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_604_74#_M1011_g 0.0235674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_604_74#_M1003_g 0.0256973f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_33 VNB N_A_604_74#_c_672_n 6.38898e-19 $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.295
cc_34 VNB N_A_604_74#_c_673_n 0.00930435f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_35 VNB N_A_604_74#_c_674_n 0.00543267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_604_74#_c_675_n 0.00363392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_604_74#_c_676_n 0.0017874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_604_74#_c_677_n 0.0329511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_604_74#_c_678_n 0.0151919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_604_74#_c_679_n 0.0256034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_604_74#_c_680_n 0.00760734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_604_74#_c_681_n 0.00372827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_604_74#_c_682_n 0.00852463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_SET_B_M1009_g 0.035936f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.98
cc_45 VNB N_SET_B_c_813_n 0.0171269f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_46 VNB N_SET_B_c_814_n 0.0751012f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_47 VNB N_SET_B_c_815_n 0.0255015f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_48 VNB N_SET_B_c_816_n 0.00308008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_224_350#_M1020_g 0.0217848f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_50 VNB N_A_224_350#_c_938_n 0.0336873f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_51 VNB N_A_224_350#_M1013_g 0.0288323f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_52 VNB N_A_224_350#_c_940_n 0.0108167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_224_350#_c_941_n 0.00127264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_224_350#_M1018_g 0.0566135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_224_350#_c_943_n 0.0111885f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_224_350#_c_944_n 0.0174729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_224_350#_c_945_n 0.024013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_224_350#_c_946_n 0.00958684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_224_350#_c_947_n 0.00191874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_224_350#_c_948_n 0.0130637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1470_48#_M1019_g 0.0329919f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_62 VNB N_A_1470_48#_M1002_g 0.00652993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1470_48#_c_1122_n 0.00354417f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.145
cc_64 VNB N_A_1470_48#_c_1123_n 0.0217852f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_65 VNB N_A_1470_48#_c_1124_n 0.022578f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.99
cc_66 VNB N_A_1470_48#_c_1125_n 0.00656706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1470_48#_c_1126_n 0.00860457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1470_48#_c_1127_n 0.0436381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1301_392#_c_1203_n 0.00991707f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.21
cc_70 VNB N_A_1301_392#_M1005_g 0.0535121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1301_392#_M1026_g 0.0605586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1301_392#_c_1206_n 0.00572865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1301_392#_c_1207_n 0.00234709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1301_392#_c_1208_n 0.0195349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1301_392#_c_1209_n 2.14136e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1301_392#_c_1210_n 0.00696087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1902_74#_c_1376_n 0.0226655f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.98
cc_78 VNB N_A_1902_74#_M1025_g 0.00735078f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_79 VNB N_A_1902_74#_c_1378_n 0.00572238f $X=-0.19 $Y=-0.245 $X2=0.64
+ $Y2=1.145
cc_80 VNB N_A_1902_74#_c_1379_n 0.00265372f $X=-0.19 $Y=-0.245 $X2=0.605
+ $Y2=1.825
cc_81 VNB N_A_1902_74#_c_1380_n 0.00232958f $X=-0.19 $Y=-0.245 $X2=0.605
+ $Y2=1.99
cc_82 VNB N_A_1902_74#_c_1381_n 0.00656177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1902_74#_c_1382_n 0.0022061f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_84 VNB N_A_1902_74#_c_1383_n 0.00342286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1902_74#_c_1384_n 0.0432868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_27_74#_c_1432_n 0.0147509f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.145
cc_87 VNB N_A_27_74#_c_1433_n 0.0402619f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.98
cc_88 VNB N_A_27_74#_c_1434_n 0.00501934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_27_74#_c_1435_n 0.00855805f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_90 VNB N_A_27_74#_c_1436_n 0.0040388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VPWR_c_1499_n 0.462217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB Q 0.0093606f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_93 VNB Q 0.0310914f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.58
cc_94 VNB N_Q_c_1638_n 0.0243787f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_95 VNB N_VGND_c_1654_n 0.0077412f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.825
cc_96 VNB N_VGND_c_1655_n 0.0224525f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.145
cc_97 VNB N_VGND_c_1656_n 0.00766269f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.665
cc_98 VNB N_VGND_c_1657_n 0.0168995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1658_n 0.0173928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1659_n 0.0106822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1660_n 0.0350591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1661_n 0.00615791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1662_n 0.034271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1663_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1664_n 0.0173128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1665_n 0.0593495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1666_n 0.0213543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1667_n 0.611249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1668_n 0.00461913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1669_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1670_n 0.007312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1671_n 0.0501753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1672_n 0.0294264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VPB N_D_c_239_n 0.0122244f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.79
cc_115 VPB N_D_M1008_g 0.0630162f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=2.75
cc_116 VPB N_D_c_242_n 0.00233492f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_117 VPB N_D_c_246_n 0.0252464f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_118 VPB N_CLK_M1004_g 0.0242591f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.99
cc_119 VPB N_A_398_74#_M1017_g 0.0239f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_120 VPB N_A_398_74#_c_311_n 0.0139588f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_121 VPB N_A_398_74#_c_312_n 8.09759e-19 $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_122 VPB N_A_398_74#_M1027_g 0.0266463f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.99
cc_123 VPB N_A_398_74#_c_333_n 0.0178571f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_124 VPB N_A_398_74#_c_334_n 0.00417353f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_125 VPB N_A_398_74#_c_335_n 0.0195502f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_126 VPB N_A_398_74#_c_336_n 0.00392743f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_127 VPB N_A_398_74#_c_337_n 0.00104738f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_128 VPB N_A_398_74#_c_338_n 0.0267392f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_129 VPB N_A_398_74#_c_318_n 0.00520082f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_130 VPB N_A_398_74#_c_340_n 0.00363609f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_131 VPB N_A_398_74#_c_341_n 0.0149448f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_132 VPB N_A_398_74#_c_342_n 0.00517621f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_133 VPB N_A_398_74#_c_343_n 0.0154856f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_134 VPB N_A_398_74#_c_344_n 0.00260538f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_135 VPB N_A_398_74#_c_345_n 0.00190156f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_136 VPB N_A_398_74#_c_346_n 9.11874e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_137 VPB N_A_398_74#_c_319_n 0.00300526f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_138 VPB N_A_398_74#_c_322_n 0.00646805f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_139 VPB N_A_398_74#_c_349_n 0.0013133f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_140 VPB N_A_398_74#_c_350_n 0.00643404f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_141 VPB N_A_398_74#_c_327_n 0.0234914f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_142 VPB N_A_398_74#_c_352_n 0.0382357f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_143 VPB N_A_760_395#_M1030_g 0.0224413f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_144 VPB N_A_760_395#_c_591_n 0.0011019f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.145
cc_145 VPB N_A_760_395#_c_596_n 0.00787198f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_146 VPB N_A_760_395#_c_597_n 0.0662587f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.99
cc_147 VPB N_A_760_395#_c_598_n 0.0029891f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_148 VPB N_A_760_395#_c_599_n 9.19853e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_149 VPB N_A_760_395#_c_600_n 0.00284926f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_150 VPB N_A_604_74#_M1000_g 0.0466672f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_151 VPB N_A_604_74#_M1001_g 0.0220037f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_152 VPB N_A_604_74#_c_677_n 0.0207793f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_153 VPB N_A_604_74#_c_678_n 0.00292093f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_154 VPB N_A_604_74#_c_679_n 0.00638595f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_155 VPB N_A_604_74#_c_688_n 0.00687801f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_156 VPB N_A_604_74#_c_680_n 0.0102885f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_157 VPB N_SET_B_M1012_g 0.0213622f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=1.99
cc_158 VPB N_SET_B_M1009_g 0.0169973f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.98
cc_159 VPB N_SET_B_c_819_n 0.0375852f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_160 VPB N_SET_B_M1006_g 0.0338545f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_161 VPB N_SET_B_c_815_n 0.0213472f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_162 VPB N_SET_B_c_822_n 0.0227051f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=0.98
cc_163 VPB N_SET_B_c_823_n 0.00140339f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.825
cc_164 VPB N_SET_B_c_824_n 0.00109254f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.99
cc_165 VPB SET_B 0.00521469f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_166 VPB N_SET_B_c_826_n 0.0397593f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_167 VPB N_SET_B_c_816_n 0.0015276f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_168 VPB N_A_224_350#_M1010_g 0.0200311f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_169 VPB N_A_224_350#_c_950_n 0.0765719f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_170 VPB N_A_224_350#_c_951_n 0.0558158f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.825
cc_171 VPB N_A_224_350#_c_952_n 0.0125859f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_172 VPB N_A_224_350#_M1015_g 0.0354475f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.665
cc_173 VPB N_A_224_350#_c_954_n 0.219497f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_174 VPB N_A_224_350#_M1021_g 0.017531f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_175 VPB N_A_224_350#_c_940_n 0.0394429f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_176 VPB N_A_224_350#_c_941_n 0.00760553f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_177 VPB N_A_224_350#_c_943_n 7.74251e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_178 VPB N_A_224_350#_c_944_n 0.00575231f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_179 VPB N_A_224_350#_c_945_n 5.67618e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_180 VPB N_A_224_350#_c_961_n 0.00898883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_181 VPB N_A_224_350#_c_946_n 0.00374312f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_182 VPB N_A_224_350#_c_963_n 0.00458484f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_183 VPB N_A_224_350#_c_947_n 7.55963e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_184 VPB N_A_224_350#_c_965_n 0.0125877f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_185 VPB N_A_1470_48#_M1002_g 0.06165f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_186 VPB N_A_1470_48#_c_1129_n 0.00620556f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_187 VPB N_A_1470_48#_c_1126_n 0.0132095f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_188 VPB N_A_1301_392#_c_1203_n 0.0107504f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.21
cc_189 VPB N_A_1301_392#_M1016_g 0.0283578f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=0.98
cc_190 VPB N_A_1301_392#_c_1213_n 0.0504309f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_191 VPB N_A_1301_392#_M1026_g 0.0077247f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_192 VPB N_A_1301_392#_c_1215_n 0.0334962f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_193 VPB N_A_1301_392#_c_1216_n 0.00827353f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_194 VPB N_A_1301_392#_c_1217_n 0.0205348f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_195 VPB N_A_1301_392#_c_1218_n 0.00290592f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_196 VPB N_A_1301_392#_c_1219_n 0.00475263f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_197 VPB N_A_1301_392#_c_1220_n 0.00270883f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_198 VPB N_A_1301_392#_c_1221_n 4.99227e-19 $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_199 VPB N_A_1301_392#_c_1222_n 0.00632069f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_200 VPB N_A_1301_392#_c_1223_n 0.0028111f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_201 VPB N_A_1301_392#_c_1224_n 0.00564138f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_202 VPB N_A_1301_392#_c_1225_n 0.0157672f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_203 VPB N_A_1301_392#_c_1226_n 0.0237245f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_204 VPB N_A_1301_392#_c_1227_n 0.00103878f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_205 VPB N_A_1301_392#_c_1228_n 0.0033822f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_206 VPB N_A_1301_392#_c_1229_n 0.00217618f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_207 VPB N_A_1902_74#_M1025_g 0.0291718f $X=-0.19 $Y=1.66 $X2=0.635 $Y2=1.58
cc_208 VPB N_A_1902_74#_c_1380_n 0.0139952f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=1.99
cc_209 VPB N_A_27_74#_c_1433_n 0.0270482f $X=-0.19 $Y=1.66 $X2=0.605 $Y2=0.98
cc_210 VPB N_A_27_74#_c_1438_n 0.0256582f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.825
cc_211 VPB N_A_27_74#_c_1439_n 0.0251386f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.145
cc_212 VPB N_A_27_74#_c_1440_n 0.013057f $X=-0.19 $Y=1.66 $X2=0.64 $Y2=1.295
cc_213 VPB N_A_27_74#_c_1434_n 0.00288606f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_214 VPB N_A_27_74#_c_1442_n 0.0109364f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1500_n 0.0114356f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1501_n 0.0062626f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1502_n 0.00520835f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1503_n 0.00629929f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1504_n 0.00795074f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1505_n 0.0126929f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1506_n 0.0141737f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1507_n 0.0303002f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1508_n 0.00330333f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1509_n 0.0532773f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1510_n 0.00324402f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1511_n 0.0177091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1512_n 0.0207798f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1513_n 0.0489399f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1514_n 0.0206844f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1515_n 0.0347486f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1516_n 0.0177091f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1499_n 0.115457f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1518_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1519_n 0.00632158f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1520_n 0.00370284f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1521_n 0.0047828f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1522_n 0.0061274f $X=-0.19 $Y=1.66 $X2=0 $Y2=0
cc_238 VPB Q 0.0544426f $X=-0.19 $Y=1.66 $X2=0.495 $Y2=0.58
cc_239 N_D_c_239_n N_CLK_M1004_g 0.00422845f $X=0.605 $Y=1.79 $X2=0 $Y2=0
cc_240 N_D_c_239_n N_CLK_c_275_n 0.00573699f $X=0.605 $Y=1.79 $X2=0 $Y2=0
cc_241 N_D_c_241_n N_CLK_c_276_n 0.00230074f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_242 N_D_c_239_n N_A_224_350#_c_946_n 0.00356228f $X=0.605 $Y=1.79 $X2=0 $Y2=0
cc_243 N_D_M1028_g N_A_224_350#_c_948_n 0.00616966f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_244 N_D_c_241_n N_A_224_350#_c_948_n 0.00356228f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_245 N_D_c_242_n N_A_224_350#_c_948_n 0.0557245f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_246 N_D_c_239_n N_A_224_350#_c_965_n 0.00288057f $X=0.605 $Y=1.79 $X2=0 $Y2=0
cc_247 N_D_M1008_g N_A_224_350#_c_965_n 0.00213438f $X=0.495 $Y=2.75 $X2=0 $Y2=0
cc_248 N_D_c_242_n N_A_224_350#_c_965_n 0.0223599f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_249 N_D_M1028_g N_A_27_74#_c_1432_n 0.00146353f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_250 N_D_M1028_g N_A_27_74#_c_1433_n 0.00594476f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_251 N_D_c_241_n N_A_27_74#_c_1433_n 0.0337586f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_252 N_D_c_242_n N_A_27_74#_c_1433_n 0.0671094f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_253 N_D_M1008_g N_A_27_74#_c_1438_n 0.00686358f $X=0.495 $Y=2.75 $X2=0 $Y2=0
cc_254 N_D_M1008_g N_A_27_74#_c_1439_n 0.022299f $X=0.495 $Y=2.75 $X2=0 $Y2=0
cc_255 N_D_c_242_n N_A_27_74#_c_1439_n 0.0197854f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_256 N_D_c_246_n N_A_27_74#_c_1439_n 0.00141894f $X=0.64 $Y=1.825 $X2=0 $Y2=0
cc_257 N_D_M1008_g N_VPWR_c_1500_n 0.0137033f $X=0.495 $Y=2.75 $X2=0 $Y2=0
cc_258 N_D_M1008_g N_VPWR_c_1511_n 0.00460063f $X=0.495 $Y=2.75 $X2=0 $Y2=0
cc_259 N_D_M1008_g N_VPWR_c_1499_n 0.00912261f $X=0.495 $Y=2.75 $X2=0 $Y2=0
cc_260 N_D_M1028_g N_VGND_c_1654_n 0.0137856f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_261 N_D_c_241_n N_VGND_c_1654_n 0.00175174f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_262 N_D_c_242_n N_VGND_c_1654_n 0.0220022f $X=0.64 $Y=1.145 $X2=0 $Y2=0
cc_263 N_D_M1028_g N_VGND_c_1664_n 0.00383152f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_264 N_D_M1028_g N_VGND_c_1667_n 0.00761198f $X=0.495 $Y=0.58 $X2=0 $Y2=0
cc_265 N_CLK_c_276_n N_A_398_74#_c_314_n 4.9956e-19 $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_266 CLK N_A_224_350#_M1020_g 0.00480673f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_267 N_CLK_c_275_n N_A_224_350#_M1020_g 0.021211f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_268 N_CLK_c_276_n N_A_224_350#_M1020_g 0.0126626f $X=1.465 $Y=1.22 $X2=0
+ $Y2=0
cc_269 N_CLK_M1004_g N_A_224_350#_c_943_n 0.0496882f $X=1.48 $Y=2.31 $X2=0 $Y2=0
cc_270 N_CLK_M1004_g N_A_224_350#_c_946_n 0.00367721f $X=1.48 $Y=2.31 $X2=0
+ $Y2=0
cc_271 CLK N_A_224_350#_c_946_n 0.0287772f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_272 N_CLK_c_275_n N_A_224_350#_c_946_n 0.00297156f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_273 N_CLK_c_276_n N_A_224_350#_c_946_n 0.00327386f $X=1.465 $Y=1.22 $X2=0
+ $Y2=0
cc_274 N_CLK_M1004_g N_A_224_350#_c_963_n 0.00927844f $X=1.48 $Y=2.31 $X2=0
+ $Y2=0
cc_275 N_CLK_c_275_n N_A_224_350#_c_963_n 0.00134523f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_276 N_CLK_M1004_g N_A_224_350#_c_947_n 8.09239e-19 $X=1.48 $Y=2.31 $X2=0
+ $Y2=0
cc_277 CLK N_A_224_350#_c_947_n 0.0217771f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_278 N_CLK_c_275_n N_A_224_350#_c_947_n 2.17092e-19 $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_279 CLK N_A_224_350#_c_948_n 0.00762435f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_280 N_CLK_c_275_n N_A_224_350#_c_948_n 0.00114344f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_281 N_CLK_c_276_n N_A_224_350#_c_948_n 0.00780781f $X=1.465 $Y=1.22 $X2=0
+ $Y2=0
cc_282 N_CLK_M1004_g N_A_224_350#_c_965_n 0.00511654f $X=1.48 $Y=2.31 $X2=0
+ $Y2=0
cc_283 CLK N_A_224_350#_c_965_n 0.0368043f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_284 N_CLK_c_275_n N_A_224_350#_c_965_n 0.00231845f $X=1.465 $Y=1.385 $X2=0
+ $Y2=0
cc_285 N_CLK_M1004_g N_A_27_74#_c_1439_n 0.0176851f $X=1.48 $Y=2.31 $X2=0 $Y2=0
cc_286 N_CLK_M1004_g N_VPWR_c_1500_n 0.00730314f $X=1.48 $Y=2.31 $X2=0 $Y2=0
cc_287 N_CLK_M1004_g N_VPWR_c_1501_n 0.0124409f $X=1.48 $Y=2.31 $X2=0 $Y2=0
cc_288 N_CLK_M1004_g N_VPWR_c_1512_n 0.00512593f $X=1.48 $Y=2.31 $X2=0 $Y2=0
cc_289 N_CLK_M1004_g N_VPWR_c_1499_n 0.00520946f $X=1.48 $Y=2.31 $X2=0 $Y2=0
cc_290 N_CLK_c_276_n N_VGND_c_1654_n 0.00299692f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_291 N_CLK_c_276_n N_VGND_c_1655_n 0.00434272f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_292 CLK N_VGND_c_1656_n 0.0145969f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_293 N_CLK_c_276_n N_VGND_c_1656_n 0.0027473f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_294 N_CLK_c_276_n N_VGND_c_1667_n 0.00825381f $X=1.465 $Y=1.22 $X2=0 $Y2=0
cc_295 N_A_398_74#_c_340_n N_A_760_395#_M1030_g 0.00330468f $X=3.67 $Y=2.905
+ $X2=0 $Y2=0
cc_296 N_A_398_74#_c_341_n N_A_760_395#_M1030_g 0.0131249f $X=4.4 $Y=2.17 $X2=0
+ $Y2=0
cc_297 N_A_398_74#_c_342_n N_A_760_395#_M1030_g 0.00210924f $X=4.485 $Y=2.905
+ $X2=0 $Y2=0
cc_298 N_A_398_74#_M1024_g N_A_760_395#_c_590_n 0.0421262f $X=3.625 $Y=0.58
+ $X2=0 $Y2=0
cc_299 N_A_398_74#_c_318_n N_A_760_395#_c_591_n 4.36009e-19 $X=3.67 $Y=1.6 $X2=0
+ $Y2=0
cc_300 N_A_398_74#_c_327_n N_A_760_395#_c_591_n 0.00484587f $X=3.67 $Y=1.51
+ $X2=0 $Y2=0
cc_301 N_A_398_74#_c_341_n N_A_760_395#_c_596_n 0.0143583f $X=4.4 $Y=2.17 $X2=0
+ $Y2=0
cc_302 N_A_398_74#_c_333_n N_A_760_395#_c_597_n 0.00127104f $X=2.95 $Y=2.105
+ $X2=0 $Y2=0
cc_303 N_A_398_74#_c_318_n N_A_760_395#_c_597_n 0.00695043f $X=3.67 $Y=1.6 $X2=0
+ $Y2=0
cc_304 N_A_398_74#_c_341_n N_A_760_395#_c_597_n 0.0196904f $X=4.4 $Y=2.17 $X2=0
+ $Y2=0
cc_305 N_A_398_74#_c_327_n N_A_760_395#_c_597_n 0.0135352f $X=3.67 $Y=1.51 $X2=0
+ $Y2=0
cc_306 N_A_398_74#_c_318_n N_A_760_395#_c_598_n 0.0114156f $X=3.67 $Y=1.6 $X2=0
+ $Y2=0
cc_307 N_A_398_74#_c_341_n N_A_760_395#_c_598_n 0.0246268f $X=4.4 $Y=2.17 $X2=0
+ $Y2=0
cc_308 N_A_398_74#_c_327_n N_A_760_395#_c_598_n 2.97122e-19 $X=3.67 $Y=1.51
+ $X2=0 $Y2=0
cc_309 N_A_398_74#_c_343_n N_A_760_395#_c_599_n 0.0189597f $X=5.195 $Y=2.99
+ $X2=0 $Y2=0
cc_310 N_A_398_74#_c_341_n N_A_760_395#_c_600_n 0.0137141f $X=4.4 $Y=2.17 $X2=0
+ $Y2=0
cc_311 N_A_398_74#_c_342_n N_A_760_395#_c_600_n 0.0195772f $X=4.485 $Y=2.905
+ $X2=0 $Y2=0
cc_312 N_A_398_74#_M1024_g N_A_760_395#_c_593_n 0.00555436f $X=3.625 $Y=0.58
+ $X2=0 $Y2=0
cc_313 N_A_398_74#_c_341_n N_A_604_74#_M1000_g 0.00203712f $X=4.4 $Y=2.17 $X2=0
+ $Y2=0
cc_314 N_A_398_74#_c_342_n N_A_604_74#_M1000_g 0.0065446f $X=4.485 $Y=2.905
+ $X2=0 $Y2=0
cc_315 N_A_398_74#_c_343_n N_A_604_74#_M1000_g 0.00336499f $X=5.195 $Y=2.99
+ $X2=0 $Y2=0
cc_316 N_A_398_74#_c_345_n N_A_604_74#_M1000_g 4.94158e-19 $X=5.28 $Y=2.905
+ $X2=0 $Y2=0
cc_317 N_A_398_74#_c_345_n N_A_604_74#_M1001_g 0.00304743f $X=5.28 $Y=2.905
+ $X2=0 $Y2=0
cc_318 N_A_398_74#_c_377_p N_A_604_74#_M1001_g 0.00955249f $X=5.805 $Y=2.405
+ $X2=0 $Y2=0
cc_319 N_A_398_74#_c_378_p N_A_604_74#_M1001_g 0.0137625f $X=5.89 $Y=2.32 $X2=0
+ $Y2=0
cc_320 N_A_398_74#_c_346_n N_A_604_74#_M1001_g 0.00326296f $X=6.235 $Y=1.8 $X2=0
+ $Y2=0
cc_321 N_A_398_74#_c_380_p N_A_604_74#_M1001_g 0.00547009f $X=5.975 $Y=1.8 $X2=0
+ $Y2=0
cc_322 N_A_398_74#_c_319_n N_A_604_74#_M1001_g 0.00479832f $X=6.32 $Y=1.715
+ $X2=0 $Y2=0
cc_323 N_A_398_74#_c_321_n N_A_604_74#_M1003_g 0.00159494f $X=6.405 $Y=0.34
+ $X2=0 $Y2=0
cc_324 N_A_398_74#_c_325_n N_A_604_74#_M1003_g 0.0170948f $X=6.48 $Y=1.285 $X2=0
+ $Y2=0
cc_325 N_A_398_74#_c_326_n N_A_604_74#_M1003_g 0.00638611f $X=6.44 $Y=1.12 $X2=0
+ $Y2=0
cc_326 N_A_398_74#_c_328_n N_A_604_74#_M1003_g 0.0211037f $X=6.48 $Y=1.12 $X2=0
+ $Y2=0
cc_327 N_A_398_74#_M1024_g N_A_604_74#_c_672_n 0.00879961f $X=3.625 $Y=0.58
+ $X2=0 $Y2=0
cc_328 N_A_398_74#_c_323_n N_A_604_74#_c_672_n 0.0193151f $X=2.952 $Y=1.435
+ $X2=0 $Y2=0
cc_329 N_A_398_74#_M1024_g N_A_604_74#_c_673_n 0.00955017f $X=3.625 $Y=0.58
+ $X2=0 $Y2=0
cc_330 N_A_398_74#_c_318_n N_A_604_74#_c_673_n 0.006417f $X=3.67 $Y=1.6 $X2=0
+ $Y2=0
cc_331 N_A_398_74#_c_327_n N_A_604_74#_c_673_n 0.00266001f $X=3.67 $Y=1.51 $X2=0
+ $Y2=0
cc_332 N_A_398_74#_M1024_g N_A_604_74#_c_674_n 0.00330172f $X=3.625 $Y=0.58
+ $X2=0 $Y2=0
cc_333 N_A_398_74#_M1024_g N_A_604_74#_c_675_n 0.00111875f $X=3.625 $Y=0.58
+ $X2=0 $Y2=0
cc_334 N_A_398_74#_c_318_n N_A_604_74#_c_675_n 0.00645396f $X=3.67 $Y=1.6 $X2=0
+ $Y2=0
cc_335 N_A_398_74#_c_341_n N_A_604_74#_c_675_n 0.00422692f $X=4.4 $Y=2.17 $X2=0
+ $Y2=0
cc_336 N_A_398_74#_c_327_n N_A_604_74#_c_675_n 8.97923e-19 $X=3.67 $Y=1.51 $X2=0
+ $Y2=0
cc_337 N_A_398_74#_c_346_n N_A_604_74#_c_678_n 0.00416421f $X=6.235 $Y=1.8 $X2=0
+ $Y2=0
cc_338 N_A_398_74#_c_380_p N_A_604_74#_c_678_n 0.0123456f $X=5.975 $Y=1.8 $X2=0
+ $Y2=0
cc_339 N_A_398_74#_c_324_n N_A_604_74#_c_678_n 0.0274363f $X=6.48 $Y=1.285 $X2=0
+ $Y2=0
cc_340 N_A_398_74#_c_325_n N_A_604_74#_c_678_n 2.48355e-19 $X=6.48 $Y=1.285
+ $X2=0 $Y2=0
cc_341 N_A_398_74#_c_346_n N_A_604_74#_c_679_n 0.00200344f $X=6.235 $Y=1.8 $X2=0
+ $Y2=0
cc_342 N_A_398_74#_c_324_n N_A_604_74#_c_679_n 0.00638611f $X=6.48 $Y=1.285
+ $X2=0 $Y2=0
cc_343 N_A_398_74#_M1017_g N_A_604_74#_c_688_n 3.3119e-19 $X=2.97 $Y=2.525 $X2=0
+ $Y2=0
cc_344 N_A_398_74#_c_333_n N_A_604_74#_c_688_n 0.00151134f $X=2.95 $Y=2.105
+ $X2=0 $Y2=0
cc_345 N_A_398_74#_c_335_n N_A_604_74#_c_688_n 0.0215749f $X=3.585 $Y=2.99 $X2=0
+ $Y2=0
cc_346 N_A_398_74#_M1017_g N_A_604_74#_c_680_n 0.00296516f $X=2.97 $Y=2.525
+ $X2=0 $Y2=0
cc_347 N_A_398_74#_c_311_n N_A_604_74#_c_680_n 0.0144113f $X=3.505 $Y=1.51 $X2=0
+ $Y2=0
cc_348 N_A_398_74#_M1024_g N_A_604_74#_c_680_n 0.00781228f $X=3.625 $Y=0.58
+ $X2=0 $Y2=0
cc_349 N_A_398_74#_c_338_n N_A_604_74#_c_680_n 0.00786297f $X=2.95 $Y=1.6 $X2=0
+ $Y2=0
cc_350 N_A_398_74#_c_318_n N_A_604_74#_c_680_n 0.0470982f $X=3.67 $Y=1.6 $X2=0
+ $Y2=0
cc_351 N_A_398_74#_c_340_n N_A_604_74#_c_680_n 0.0200517f $X=3.67 $Y=2.905 $X2=0
+ $Y2=0
cc_352 N_A_398_74#_c_323_n N_A_604_74#_c_680_n 0.0797343f $X=2.952 $Y=1.435
+ $X2=0 $Y2=0
cc_353 N_A_398_74#_c_349_n N_A_604_74#_c_680_n 0.0140926f $X=3.67 $Y=2.17 $X2=0
+ $Y2=0
cc_354 N_A_398_74#_c_327_n N_A_604_74#_c_680_n 0.0015889f $X=3.67 $Y=1.51 $X2=0
+ $Y2=0
cc_355 N_A_398_74#_c_311_n N_A_604_74#_c_681_n 0.00428766f $X=3.505 $Y=1.51
+ $X2=0 $Y2=0
cc_356 N_A_398_74#_M1024_g N_A_604_74#_c_681_n 0.0041848f $X=3.625 $Y=0.58 $X2=0
+ $Y2=0
cc_357 N_A_398_74#_c_323_n N_A_604_74#_c_681_n 0.0143558f $X=2.952 $Y=1.435
+ $X2=0 $Y2=0
cc_358 N_A_398_74#_c_343_n N_SET_B_M1012_g 0.00295426f $X=5.195 $Y=2.99 $X2=0
+ $Y2=0
cc_359 N_A_398_74#_c_345_n N_SET_B_M1012_g 0.0110953f $X=5.28 $Y=2.905 $X2=0
+ $Y2=0
cc_360 N_A_398_74#_c_419_p N_SET_B_M1012_g 0.00634474f $X=5.365 $Y=2.405 $X2=0
+ $Y2=0
cc_361 N_A_398_74#_c_377_p N_SET_B_c_822_n 0.00601312f $X=5.805 $Y=2.405 $X2=0
+ $Y2=0
cc_362 N_A_398_74#_c_378_p N_SET_B_c_822_n 0.0176974f $X=5.89 $Y=2.32 $X2=0
+ $Y2=0
cc_363 N_A_398_74#_c_346_n N_SET_B_c_822_n 0.0218701f $X=6.235 $Y=1.8 $X2=0
+ $Y2=0
cc_364 N_A_398_74#_c_322_n N_SET_B_c_822_n 0.00905213f $X=7.24 $Y=1.97 $X2=0
+ $Y2=0
cc_365 N_A_398_74#_c_324_n N_SET_B_c_822_n 0.00391432f $X=6.48 $Y=1.285 $X2=0
+ $Y2=0
cc_366 N_A_398_74#_c_350_n N_SET_B_c_822_n 0.0200203f $X=7.095 $Y=2.185 $X2=0
+ $Y2=0
cc_367 N_A_398_74#_c_352_n N_SET_B_c_822_n 0.00134681f $X=7.21 $Y=2.185 $X2=0
+ $Y2=0
cc_368 N_A_398_74#_c_377_p N_SET_B_c_823_n 0.00811829f $X=5.805 $Y=2.405 $X2=0
+ $Y2=0
cc_369 N_A_398_74#_c_378_p N_SET_B_c_823_n 0.00268218f $X=5.89 $Y=2.32 $X2=0
+ $Y2=0
cc_370 N_A_398_74#_c_377_p N_SET_B_c_824_n 0.0172394f $X=5.805 $Y=2.405 $X2=0
+ $Y2=0
cc_371 N_A_398_74#_c_419_p N_SET_B_c_824_n 0.0113152f $X=5.365 $Y=2.405 $X2=0
+ $Y2=0
cc_372 N_A_398_74#_c_378_p N_SET_B_c_824_n 0.0121171f $X=5.89 $Y=2.32 $X2=0
+ $Y2=0
cc_373 N_A_398_74#_c_377_p N_SET_B_c_826_n 0.00248274f $X=5.805 $Y=2.405 $X2=0
+ $Y2=0
cc_374 N_A_398_74#_c_419_p N_SET_B_c_826_n 0.00246772f $X=5.365 $Y=2.405 $X2=0
+ $Y2=0
cc_375 N_A_398_74#_c_378_p N_SET_B_c_826_n 2.58465e-19 $X=5.89 $Y=2.32 $X2=0
+ $Y2=0
cc_376 N_A_398_74#_c_314_n N_A_224_350#_M1020_g 0.0084694f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_377 N_A_398_74#_c_316_n N_A_224_350#_M1020_g 0.00464501f $X=2.295 $Y=0.34
+ $X2=0 $Y2=0
cc_378 N_A_398_74#_c_334_n N_A_224_350#_M1010_g 7.43518e-19 $X=2.155 $Y=2.645
+ $X2=0 $Y2=0
cc_379 N_A_398_74#_c_336_n N_A_224_350#_M1010_g 9.48272e-19 $X=2.32 $Y=2.99
+ $X2=0 $Y2=0
cc_380 N_A_398_74#_M1017_g N_A_224_350#_c_950_n 0.0185232f $X=2.97 $Y=2.525
+ $X2=0 $Y2=0
cc_381 N_A_398_74#_c_334_n N_A_224_350#_c_950_n 0.00725312f $X=2.155 $Y=2.645
+ $X2=0 $Y2=0
cc_382 N_A_398_74#_c_335_n N_A_224_350#_c_950_n 0.0118684f $X=3.585 $Y=2.99
+ $X2=0 $Y2=0
cc_383 N_A_398_74#_c_337_n N_A_224_350#_c_950_n 3.15319e-19 $X=2.95 $Y=1.6 $X2=0
+ $Y2=0
cc_384 N_A_398_74#_c_338_n N_A_224_350#_c_950_n 0.0159248f $X=2.95 $Y=1.6 $X2=0
+ $Y2=0
cc_385 N_A_398_74#_c_312_n N_A_224_350#_c_938_n 0.0133559f $X=3.115 $Y=1.51
+ $X2=0 $Y2=0
cc_386 N_A_398_74#_c_315_n N_A_224_350#_c_938_n 0.00237401f $X=2.905 $Y=0.34
+ $X2=0 $Y2=0
cc_387 N_A_398_74#_c_317_n N_A_224_350#_c_938_n 5.11203e-19 $X=2.952 $Y=1.557
+ $X2=0 $Y2=0
cc_388 N_A_398_74#_c_323_n N_A_224_350#_c_938_n 0.0066912f $X=2.952 $Y=1.435
+ $X2=0 $Y2=0
cc_389 N_A_398_74#_M1017_g N_A_224_350#_c_951_n 0.0105864f $X=2.97 $Y=2.525
+ $X2=0 $Y2=0
cc_390 N_A_398_74#_c_335_n N_A_224_350#_c_951_n 0.0128457f $X=3.585 $Y=2.99
+ $X2=0 $Y2=0
cc_391 N_A_398_74#_M1024_g N_A_224_350#_M1013_g 0.0129251f $X=3.625 $Y=0.58
+ $X2=0 $Y2=0
cc_392 N_A_398_74#_c_314_n N_A_224_350#_M1013_g 0.00314925f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_393 N_A_398_74#_c_315_n N_A_224_350#_M1013_g 0.0102552f $X=2.905 $Y=0.34
+ $X2=0 $Y2=0
cc_394 N_A_398_74#_c_323_n N_A_224_350#_M1013_g 0.0180895f $X=2.952 $Y=1.435
+ $X2=0 $Y2=0
cc_395 N_A_398_74#_M1017_g N_A_224_350#_M1015_g 0.0108836f $X=2.97 $Y=2.525
+ $X2=0 $Y2=0
cc_396 N_A_398_74#_c_311_n N_A_224_350#_M1015_g 0.00305329f $X=3.505 $Y=1.51
+ $X2=0 $Y2=0
cc_397 N_A_398_74#_c_335_n N_A_224_350#_M1015_g 0.0184583f $X=3.585 $Y=2.99
+ $X2=0 $Y2=0
cc_398 N_A_398_74#_c_340_n N_A_224_350#_M1015_g 0.00689645f $X=3.67 $Y=2.905
+ $X2=0 $Y2=0
cc_399 N_A_398_74#_c_349_n N_A_224_350#_M1015_g 5.73944e-19 $X=3.67 $Y=2.17
+ $X2=0 $Y2=0
cc_400 N_A_398_74#_c_327_n N_A_224_350#_M1015_g 0.00234104f $X=3.67 $Y=1.51
+ $X2=0 $Y2=0
cc_401 N_A_398_74#_c_335_n N_A_224_350#_c_954_n 0.00398567f $X=3.585 $Y=2.99
+ $X2=0 $Y2=0
cc_402 N_A_398_74#_c_343_n N_A_224_350#_c_954_n 0.0128618f $X=5.195 $Y=2.99
+ $X2=0 $Y2=0
cc_403 N_A_398_74#_c_344_n N_A_224_350#_c_954_n 0.00420304f $X=4.57 $Y=2.99
+ $X2=0 $Y2=0
cc_404 N_A_398_74#_c_377_p N_A_224_350#_c_954_n 0.00503936f $X=5.805 $Y=2.405
+ $X2=0 $Y2=0
cc_405 N_A_398_74#_M1027_g N_A_224_350#_M1021_g 0.00479345f $X=7.21 $Y=2.75
+ $X2=0 $Y2=0
cc_406 N_A_398_74#_c_377_p N_A_224_350#_M1021_g 6.28501e-19 $X=5.805 $Y=2.405
+ $X2=0 $Y2=0
cc_407 N_A_398_74#_c_378_p N_A_224_350#_M1021_g 0.00166737f $X=5.89 $Y=2.32
+ $X2=0 $Y2=0
cc_408 N_A_398_74#_c_346_n N_A_224_350#_M1021_g 0.00347826f $X=6.235 $Y=1.8
+ $X2=0 $Y2=0
cc_409 N_A_398_74#_c_350_n N_A_224_350#_c_940_n 0.0024242f $X=7.095 $Y=2.185
+ $X2=0 $Y2=0
cc_410 N_A_398_74#_c_352_n N_A_224_350#_c_940_n 0.0120911f $X=7.21 $Y=2.185
+ $X2=0 $Y2=0
cc_411 N_A_398_74#_c_346_n N_A_224_350#_c_941_n 0.00334934f $X=6.235 $Y=1.8
+ $X2=0 $Y2=0
cc_412 N_A_398_74#_c_319_n N_A_224_350#_c_941_n 0.00223021f $X=6.32 $Y=1.715
+ $X2=0 $Y2=0
cc_413 N_A_398_74#_c_324_n N_A_224_350#_c_941_n 9.66107e-19 $X=6.48 $Y=1.285
+ $X2=0 $Y2=0
cc_414 N_A_398_74#_c_325_n N_A_224_350#_c_941_n 0.0205958f $X=6.48 $Y=1.285
+ $X2=0 $Y2=0
cc_415 N_A_398_74#_c_319_n N_A_224_350#_M1018_g 9.07333e-19 $X=6.32 $Y=1.715
+ $X2=0 $Y2=0
cc_416 N_A_398_74#_c_320_n N_A_224_350#_M1018_g 0.0126916f $X=7.155 $Y=0.34
+ $X2=0 $Y2=0
cc_417 N_A_398_74#_c_322_n N_A_224_350#_M1018_g 0.00917f $X=7.24 $Y=1.97 $X2=0
+ $Y2=0
cc_418 N_A_398_74#_c_324_n N_A_224_350#_M1018_g 3.35466e-19 $X=6.48 $Y=1.285
+ $X2=0 $Y2=0
cc_419 N_A_398_74#_c_325_n N_A_224_350#_M1018_g 0.0120588f $X=6.48 $Y=1.285
+ $X2=0 $Y2=0
cc_420 N_A_398_74#_c_328_n N_A_224_350#_M1018_g 0.0214931f $X=6.48 $Y=1.12 $X2=0
+ $Y2=0
cc_421 N_A_398_74#_c_314_n N_A_224_350#_c_944_n 0.00161969f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_422 N_A_398_74#_c_312_n N_A_224_350#_c_945_n 0.0159248f $X=3.115 $Y=1.51
+ $X2=0 $Y2=0
cc_423 N_A_398_74#_c_314_n N_A_224_350#_c_945_n 4.83416e-19 $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_424 N_A_398_74#_c_315_n N_A_224_350#_c_945_n 0.0033832f $X=2.905 $Y=0.34
+ $X2=0 $Y2=0
cc_425 N_A_398_74#_c_317_n N_A_224_350#_c_945_n 3.15319e-19 $X=2.952 $Y=1.557
+ $X2=0 $Y2=0
cc_426 N_A_398_74#_c_323_n N_A_224_350#_c_945_n 7.28093e-19 $X=2.952 $Y=1.435
+ $X2=0 $Y2=0
cc_427 N_A_398_74#_M1010_d N_A_224_350#_c_963_n 0.00308247f $X=2.02 $Y=1.75
+ $X2=0 $Y2=0
cc_428 N_A_398_74#_c_314_n N_A_224_350#_c_963_n 4.74438e-19 $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_429 N_A_398_74#_c_314_n N_A_224_350#_c_947_n 0.0241738f $X=2.13 $Y=0.515
+ $X2=0 $Y2=0
cc_430 N_A_398_74#_c_320_n N_A_1470_48#_M1019_g 0.00193743f $X=7.155 $Y=0.34
+ $X2=0 $Y2=0
cc_431 N_A_398_74#_c_322_n N_A_1470_48#_M1019_g 0.00702399f $X=7.24 $Y=1.97
+ $X2=0 $Y2=0
cc_432 N_A_398_74#_c_322_n N_A_1470_48#_M1002_g 0.0106677f $X=7.24 $Y=1.97 $X2=0
+ $Y2=0
cc_433 N_A_398_74#_c_350_n N_A_1470_48#_M1002_g 0.00452782f $X=7.095 $Y=2.185
+ $X2=0 $Y2=0
cc_434 N_A_398_74#_c_352_n N_A_1470_48#_M1002_g 0.0578668f $X=7.21 $Y=2.185
+ $X2=0 $Y2=0
cc_435 N_A_398_74#_c_322_n N_A_1470_48#_c_1122_n 0.043508f $X=7.24 $Y=1.97 $X2=0
+ $Y2=0
cc_436 N_A_398_74#_c_322_n N_A_1470_48#_c_1137_n 0.013546f $X=7.24 $Y=1.97 $X2=0
+ $Y2=0
cc_437 N_A_398_74#_c_320_n N_A_1301_392#_M1007_d 0.0026214f $X=7.155 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_438 N_A_398_74#_M1027_g N_A_1301_392#_c_1218_n 0.00307472f $X=7.21 $Y=2.75
+ $X2=0 $Y2=0
cc_439 N_A_398_74#_c_377_p N_A_1301_392#_c_1218_n 0.00561835f $X=5.805 $Y=2.405
+ $X2=0 $Y2=0
cc_440 N_A_398_74#_M1027_g N_A_1301_392#_c_1219_n 0.0154656f $X=7.21 $Y=2.75
+ $X2=0 $Y2=0
cc_441 N_A_398_74#_c_350_n N_A_1301_392#_c_1219_n 0.0149811f $X=7.095 $Y=2.185
+ $X2=0 $Y2=0
cc_442 N_A_398_74#_c_352_n N_A_1301_392#_c_1219_n 0.00259363f $X=7.21 $Y=2.185
+ $X2=0 $Y2=0
cc_443 N_A_398_74#_c_319_n N_A_1301_392#_c_1206_n 0.00735716f $X=6.32 $Y=1.715
+ $X2=0 $Y2=0
cc_444 N_A_398_74#_c_322_n N_A_1301_392#_c_1206_n 0.0504172f $X=7.24 $Y=1.97
+ $X2=0 $Y2=0
cc_445 N_A_398_74#_c_324_n N_A_1301_392#_c_1206_n 0.0252198f $X=6.48 $Y=1.285
+ $X2=0 $Y2=0
cc_446 N_A_398_74#_c_325_n N_A_1301_392#_c_1206_n 0.00218868f $X=6.48 $Y=1.285
+ $X2=0 $Y2=0
cc_447 N_A_398_74#_c_326_n N_A_1301_392#_c_1206_n 0.00605873f $X=6.44 $Y=1.12
+ $X2=0 $Y2=0
cc_448 N_A_398_74#_c_328_n N_A_1301_392#_c_1206_n 0.00148668f $X=6.48 $Y=1.12
+ $X2=0 $Y2=0
cc_449 N_A_398_74#_M1027_g N_A_1301_392#_c_1221_n 0.00150878f $X=7.21 $Y=2.75
+ $X2=0 $Y2=0
cc_450 N_A_398_74#_c_350_n N_A_1301_392#_c_1223_n 0.00373419f $X=7.095 $Y=2.185
+ $X2=0 $Y2=0
cc_451 N_A_398_74#_c_352_n N_A_1301_392#_c_1223_n 0.00198625f $X=7.21 $Y=2.185
+ $X2=0 $Y2=0
cc_452 N_A_398_74#_c_378_p N_A_1301_392#_c_1227_n 0.00719962f $X=5.89 $Y=2.32
+ $X2=0 $Y2=0
cc_453 N_A_398_74#_c_324_n N_A_1301_392#_c_1227_n 0.00122631f $X=6.48 $Y=1.285
+ $X2=0 $Y2=0
cc_454 N_A_398_74#_c_378_p N_A_1301_392#_c_1228_n 0.00329751f $X=5.89 $Y=2.32
+ $X2=0 $Y2=0
cc_455 N_A_398_74#_c_346_n N_A_1301_392#_c_1228_n 0.00680609f $X=6.235 $Y=1.8
+ $X2=0 $Y2=0
cc_456 N_A_398_74#_c_322_n N_A_1301_392#_c_1228_n 0.00792368f $X=7.24 $Y=1.97
+ $X2=0 $Y2=0
cc_457 N_A_398_74#_c_350_n N_A_1301_392#_c_1228_n 0.0291234f $X=7.095 $Y=2.185
+ $X2=0 $Y2=0
cc_458 N_A_398_74#_c_352_n N_A_1301_392#_c_1228_n 0.00287012f $X=7.21 $Y=2.185
+ $X2=0 $Y2=0
cc_459 N_A_398_74#_c_320_n N_A_1301_392#_c_1209_n 0.0209521f $X=7.155 $Y=0.34
+ $X2=0 $Y2=0
cc_460 N_A_398_74#_c_322_n N_A_1301_392#_c_1209_n 0.0178178f $X=7.24 $Y=1.97
+ $X2=0 $Y2=0
cc_461 N_A_398_74#_c_324_n N_A_1301_392#_c_1209_n 0.00314153f $X=6.48 $Y=1.285
+ $X2=0 $Y2=0
cc_462 N_A_398_74#_c_328_n N_A_1301_392#_c_1209_n 0.00407335f $X=6.48 $Y=1.12
+ $X2=0 $Y2=0
cc_463 N_A_398_74#_c_346_n N_A_1301_392#_c_1210_n 0.00678014f $X=6.235 $Y=1.8
+ $X2=0 $Y2=0
cc_464 N_A_398_74#_c_319_n N_A_1301_392#_c_1210_n 0.00633415f $X=6.32 $Y=1.715
+ $X2=0 $Y2=0
cc_465 N_A_398_74#_c_322_n N_A_1301_392#_c_1210_n 0.0128607f $X=7.24 $Y=1.97
+ $X2=0 $Y2=0
cc_466 N_A_398_74#_c_324_n N_A_1301_392#_c_1210_n 0.00479908f $X=6.48 $Y=1.285
+ $X2=0 $Y2=0
cc_467 N_A_398_74#_c_325_n N_A_1301_392#_c_1210_n 2.04288e-19 $X=6.48 $Y=1.285
+ $X2=0 $Y2=0
cc_468 N_A_398_74#_c_350_n N_A_1301_392#_c_1210_n 3.20086e-19 $X=7.095 $Y=2.185
+ $X2=0 $Y2=0
cc_469 N_A_398_74#_c_352_n N_A_1301_392#_c_1210_n 3.12047e-19 $X=7.21 $Y=2.185
+ $X2=0 $Y2=0
cc_470 N_A_398_74#_c_315_n N_A_27_74#_M1013_s 0.00388097f $X=2.905 $Y=0.34 $X2=0
+ $Y2=0
cc_471 N_A_398_74#_M1010_d N_A_27_74#_c_1440_n 0.00451828f $X=2.02 $Y=1.75 $X2=0
+ $Y2=0
cc_472 N_A_398_74#_M1017_g N_A_27_74#_c_1440_n 0.00851295f $X=2.97 $Y=2.525
+ $X2=0 $Y2=0
cc_473 N_A_398_74#_c_333_n N_A_27_74#_c_1440_n 0.00274088f $X=2.95 $Y=2.105
+ $X2=0 $Y2=0
cc_474 N_A_398_74#_c_334_n N_A_27_74#_c_1440_n 0.0462698f $X=2.155 $Y=2.645
+ $X2=0 $Y2=0
cc_475 N_A_398_74#_c_335_n N_A_27_74#_c_1440_n 0.0336324f $X=3.585 $Y=2.99 $X2=0
+ $Y2=0
cc_476 N_A_398_74#_c_337_n N_A_27_74#_c_1440_n 0.00983953f $X=2.95 $Y=1.6 $X2=0
+ $Y2=0
cc_477 N_A_398_74#_c_312_n N_A_27_74#_c_1434_n 0.00417645f $X=3.115 $Y=1.51
+ $X2=0 $Y2=0
cc_478 N_A_398_74#_c_317_n N_A_27_74#_c_1434_n 0.0458823f $X=2.952 $Y=1.557
+ $X2=0 $Y2=0
cc_479 N_A_398_74#_c_323_n N_A_27_74#_c_1434_n 0.0281153f $X=2.952 $Y=1.435
+ $X2=0 $Y2=0
cc_480 N_A_398_74#_c_314_n N_A_27_74#_c_1436_n 0.0368021f $X=2.13 $Y=0.515 $X2=0
+ $Y2=0
cc_481 N_A_398_74#_c_315_n N_A_27_74#_c_1436_n 0.0186907f $X=2.905 $Y=0.34 $X2=0
+ $Y2=0
cc_482 N_A_398_74#_c_323_n N_A_27_74#_c_1436_n 0.0239087f $X=2.952 $Y=1.435
+ $X2=0 $Y2=0
cc_483 N_A_398_74#_c_342_n N_VPWR_M1030_d 0.00828721f $X=4.485 $Y=2.905 $X2=0
+ $Y2=0
cc_484 N_A_398_74#_c_345_n N_VPWR_M1012_d 0.00320106f $X=5.28 $Y=2.905 $X2=0
+ $Y2=0
cc_485 N_A_398_74#_c_377_p N_VPWR_M1012_d 0.00952719f $X=5.805 $Y=2.405 $X2=0
+ $Y2=0
cc_486 N_A_398_74#_c_419_p N_VPWR_M1012_d 4.61723e-19 $X=5.365 $Y=2.405 $X2=0
+ $Y2=0
cc_487 N_A_398_74#_c_334_n N_VPWR_c_1501_n 0.0122108f $X=2.155 $Y=2.645 $X2=0
+ $Y2=0
cc_488 N_A_398_74#_c_336_n N_VPWR_c_1501_n 0.0130052f $X=2.32 $Y=2.99 $X2=0
+ $Y2=0
cc_489 N_A_398_74#_c_335_n N_VPWR_c_1502_n 0.0134896f $X=3.585 $Y=2.99 $X2=0
+ $Y2=0
cc_490 N_A_398_74#_c_340_n N_VPWR_c_1502_n 0.0216392f $X=3.67 $Y=2.905 $X2=0
+ $Y2=0
cc_491 N_A_398_74#_c_341_n N_VPWR_c_1502_n 0.0201983f $X=4.4 $Y=2.17 $X2=0 $Y2=0
cc_492 N_A_398_74#_c_342_n N_VPWR_c_1502_n 0.036656f $X=4.485 $Y=2.905 $X2=0
+ $Y2=0
cc_493 N_A_398_74#_c_344_n N_VPWR_c_1502_n 0.0148639f $X=4.57 $Y=2.99 $X2=0
+ $Y2=0
cc_494 N_A_398_74#_c_343_n N_VPWR_c_1503_n 0.0146521f $X=5.195 $Y=2.99 $X2=0
+ $Y2=0
cc_495 N_A_398_74#_c_345_n N_VPWR_c_1503_n 0.0185131f $X=5.28 $Y=2.905 $X2=0
+ $Y2=0
cc_496 N_A_398_74#_c_377_p N_VPWR_c_1503_n 0.0174222f $X=5.805 $Y=2.405 $X2=0
+ $Y2=0
cc_497 N_A_398_74#_c_343_n N_VPWR_c_1507_n 0.0517789f $X=5.195 $Y=2.99 $X2=0
+ $Y2=0
cc_498 N_A_398_74#_c_344_n N_VPWR_c_1507_n 0.0115893f $X=4.57 $Y=2.99 $X2=0
+ $Y2=0
cc_499 N_A_398_74#_M1027_g N_VPWR_c_1509_n 0.00349978f $X=7.21 $Y=2.75 $X2=0
+ $Y2=0
cc_500 N_A_398_74#_c_335_n N_VPWR_c_1513_n 0.0920449f $X=3.585 $Y=2.99 $X2=0
+ $Y2=0
cc_501 N_A_398_74#_c_336_n N_VPWR_c_1513_n 0.0179117f $X=2.32 $Y=2.99 $X2=0
+ $Y2=0
cc_502 N_A_398_74#_M1027_g N_VPWR_c_1499_n 0.0043189f $X=7.21 $Y=2.75 $X2=0
+ $Y2=0
cc_503 N_A_398_74#_c_335_n N_VPWR_c_1499_n 0.0482875f $X=3.585 $Y=2.99 $X2=0
+ $Y2=0
cc_504 N_A_398_74#_c_336_n N_VPWR_c_1499_n 0.00971754f $X=2.32 $Y=2.99 $X2=0
+ $Y2=0
cc_505 N_A_398_74#_c_343_n N_VPWR_c_1499_n 0.0268314f $X=5.195 $Y=2.99 $X2=0
+ $Y2=0
cc_506 N_A_398_74#_c_344_n N_VPWR_c_1499_n 0.00583135f $X=4.57 $Y=2.99 $X2=0
+ $Y2=0
cc_507 N_A_398_74#_c_377_p N_VPWR_c_1499_n 0.0121237f $X=5.805 $Y=2.405 $X2=0
+ $Y2=0
cc_508 N_A_398_74#_c_340_n A_712_463# 0.0020577f $X=3.67 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_509 N_A_398_74#_c_346_n A_1200_341# 0.00859065f $X=6.235 $Y=1.8 $X2=-0.19
+ $Y2=-0.245
cc_510 N_A_398_74#_c_316_n N_VGND_c_1656_n 0.010974f $X=2.295 $Y=0.34 $X2=0
+ $Y2=0
cc_511 N_A_398_74#_M1024_g N_VGND_c_1657_n 0.0016309f $X=3.625 $Y=0.58 $X2=0
+ $Y2=0
cc_512 N_A_398_74#_c_321_n N_VGND_c_1658_n 0.0096522f $X=6.405 $Y=0.34 $X2=0
+ $Y2=0
cc_513 N_A_398_74#_c_326_n N_VGND_c_1658_n 0.0300437f $X=6.44 $Y=1.12 $X2=0
+ $Y2=0
cc_514 N_A_398_74#_c_328_n N_VGND_c_1658_n 4.40417e-19 $X=6.48 $Y=1.12 $X2=0
+ $Y2=0
cc_515 N_A_398_74#_M1024_g N_VGND_c_1665_n 0.00435647f $X=3.625 $Y=0.58 $X2=0
+ $Y2=0
cc_516 N_A_398_74#_c_315_n N_VGND_c_1665_n 0.0509205f $X=2.905 $Y=0.34 $X2=0
+ $Y2=0
cc_517 N_A_398_74#_c_316_n N_VGND_c_1665_n 0.0235688f $X=2.295 $Y=0.34 $X2=0
+ $Y2=0
cc_518 N_A_398_74#_M1024_g N_VGND_c_1667_n 0.00451174f $X=3.625 $Y=0.58 $X2=0
+ $Y2=0
cc_519 N_A_398_74#_c_315_n N_VGND_c_1667_n 0.0288509f $X=2.905 $Y=0.34 $X2=0
+ $Y2=0
cc_520 N_A_398_74#_c_316_n N_VGND_c_1667_n 0.0127152f $X=2.295 $Y=0.34 $X2=0
+ $Y2=0
cc_521 N_A_398_74#_c_320_n N_VGND_c_1667_n 0.0334343f $X=7.155 $Y=0.34 $X2=0
+ $Y2=0
cc_522 N_A_398_74#_c_321_n N_VGND_c_1667_n 0.00660921f $X=6.405 $Y=0.34 $X2=0
+ $Y2=0
cc_523 N_A_398_74#_c_328_n N_VGND_c_1667_n 0.00355134f $X=6.48 $Y=1.12 $X2=0
+ $Y2=0
cc_524 N_A_398_74#_c_320_n N_VGND_c_1671_n 0.0595689f $X=7.155 $Y=0.34 $X2=0
+ $Y2=0
cc_525 N_A_398_74#_c_321_n N_VGND_c_1671_n 0.0121867f $X=6.405 $Y=0.34 $X2=0
+ $Y2=0
cc_526 N_A_398_74#_c_328_n N_VGND_c_1671_n 0.00278271f $X=6.48 $Y=1.12 $X2=0
+ $Y2=0
cc_527 N_A_398_74#_c_320_n N_VGND_c_1672_n 0.00508483f $X=7.155 $Y=0.34 $X2=0
+ $Y2=0
cc_528 N_A_398_74#_c_321_n A_1215_74# 6.96266e-19 $X=6.405 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_529 N_A_398_74#_c_326_n A_1215_74# 0.00925603f $X=6.44 $Y=1.12 $X2=-0.19
+ $Y2=-0.245
cc_530 N_A_398_74#_c_322_n A_1422_74# 0.00132675f $X=7.24 $Y=1.97 $X2=-0.19
+ $Y2=-0.245
cc_531 N_A_760_395#_M1030_g N_A_604_74#_M1000_g 0.005915f $X=3.89 $Y=2.525 $X2=0
+ $Y2=0
cc_532 N_A_760_395#_c_596_n N_A_604_74#_M1000_g 0.0137688f $X=4.74 $Y=1.83 $X2=0
+ $Y2=0
cc_533 N_A_760_395#_c_597_n N_A_604_74#_M1000_g 0.0047964f $X=4.22 $Y=1.8 $X2=0
+ $Y2=0
cc_534 N_A_760_395#_c_598_n N_A_604_74#_M1000_g 3.89547e-19 $X=4.385 $Y=1.8
+ $X2=0 $Y2=0
cc_535 N_A_760_395#_c_599_n N_A_604_74#_M1000_g 0.00659412f $X=4.94 $Y=2.525
+ $X2=0 $Y2=0
cc_536 N_A_760_395#_c_600_n N_A_604_74#_M1000_g 0.00940021f $X=4.882 $Y=2.32
+ $X2=0 $Y2=0
cc_537 N_A_760_395#_c_592_n N_A_604_74#_M1011_g 0.0133534f $X=4.43 $Y=1.065
+ $X2=0 $Y2=0
cc_538 N_A_760_395#_c_593_n N_A_604_74#_M1011_g 0.00789805f $X=4.31 $Y=1.065
+ $X2=0 $Y2=0
cc_539 N_A_760_395#_c_590_n N_A_604_74#_c_672_n 0.00158982f $X=4.015 $Y=0.9
+ $X2=0 $Y2=0
cc_540 N_A_760_395#_c_590_n N_A_604_74#_c_673_n 0.00563242f $X=4.015 $Y=0.9
+ $X2=0 $Y2=0
cc_541 N_A_760_395#_c_592_n N_A_604_74#_c_673_n 0.0143115f $X=4.43 $Y=1.065
+ $X2=0 $Y2=0
cc_542 N_A_760_395#_c_593_n N_A_604_74#_c_673_n 0.00481084f $X=4.31 $Y=1.065
+ $X2=0 $Y2=0
cc_543 N_A_760_395#_c_592_n N_A_604_74#_c_674_n 0.0116769f $X=4.43 $Y=1.065
+ $X2=0 $Y2=0
cc_544 N_A_760_395#_c_593_n N_A_604_74#_c_674_n 0.00940516f $X=4.31 $Y=1.065
+ $X2=0 $Y2=0
cc_545 N_A_760_395#_c_597_n N_A_604_74#_c_675_n 0.00310835f $X=4.22 $Y=1.8 $X2=0
+ $Y2=0
cc_546 N_A_760_395#_c_598_n N_A_604_74#_c_675_n 0.00328547f $X=4.385 $Y=1.8
+ $X2=0 $Y2=0
cc_547 N_A_760_395#_c_591_n N_A_604_74#_c_676_n 7.77761e-19 $X=4.31 $Y=1.59
+ $X2=0 $Y2=0
cc_548 N_A_760_395#_c_596_n N_A_604_74#_c_676_n 0.0078376f $X=4.74 $Y=1.83 $X2=0
+ $Y2=0
cc_549 N_A_760_395#_c_592_n N_A_604_74#_c_676_n 0.0155653f $X=4.43 $Y=1.065
+ $X2=0 $Y2=0
cc_550 N_A_760_395#_c_591_n N_A_604_74#_c_677_n 0.0129763f $X=4.31 $Y=1.59 $X2=0
+ $Y2=0
cc_551 N_A_760_395#_c_596_n N_A_604_74#_c_677_n 0.00260787f $X=4.74 $Y=1.83
+ $X2=0 $Y2=0
cc_552 N_A_760_395#_c_597_n N_A_604_74#_c_677_n 0.0212162f $X=4.22 $Y=1.8 $X2=0
+ $Y2=0
cc_553 N_A_760_395#_c_592_n N_A_604_74#_c_677_n 0.00508841f $X=4.43 $Y=1.065
+ $X2=0 $Y2=0
cc_554 N_A_760_395#_c_593_n N_A_604_74#_c_677_n 9.61087e-19 $X=4.31 $Y=1.065
+ $X2=0 $Y2=0
cc_555 N_A_760_395#_c_597_n N_A_604_74#_c_680_n 5.56508e-19 $X=4.22 $Y=1.8 $X2=0
+ $Y2=0
cc_556 N_A_760_395#_c_591_n N_A_604_74#_c_682_n 0.0115265f $X=4.31 $Y=1.59 $X2=0
+ $Y2=0
cc_557 N_A_760_395#_c_596_n N_A_604_74#_c_682_n 0.0246688f $X=4.74 $Y=1.83 $X2=0
+ $Y2=0
cc_558 N_A_760_395#_c_597_n N_A_604_74#_c_682_n 0.00165923f $X=4.22 $Y=1.8 $X2=0
+ $Y2=0
cc_559 N_A_760_395#_c_598_n N_A_604_74#_c_682_n 0.0206091f $X=4.385 $Y=1.8 $X2=0
+ $Y2=0
cc_560 N_A_760_395#_c_592_n N_A_604_74#_c_682_n 0.0363264f $X=4.43 $Y=1.065
+ $X2=0 $Y2=0
cc_561 N_A_760_395#_c_593_n N_A_604_74#_c_682_n 0.00645968f $X=4.31 $Y=1.065
+ $X2=0 $Y2=0
cc_562 N_A_760_395#_c_596_n N_SET_B_M1009_g 0.00164293f $X=4.74 $Y=1.83 $X2=0
+ $Y2=0
cc_563 N_A_760_395#_c_592_n N_SET_B_M1009_g 0.00135154f $X=4.43 $Y=1.065 $X2=0
+ $Y2=0
cc_564 N_A_760_395#_c_600_n N_SET_B_c_823_n 8.99889e-19 $X=4.882 $Y=2.32 $X2=0
+ $Y2=0
cc_565 N_A_760_395#_c_596_n N_SET_B_c_824_n 0.00825937f $X=4.74 $Y=1.83 $X2=0
+ $Y2=0
cc_566 N_A_760_395#_c_600_n N_SET_B_c_824_n 0.0176783f $X=4.882 $Y=2.32 $X2=0
+ $Y2=0
cc_567 N_A_760_395#_c_596_n N_SET_B_c_826_n 7.05056e-19 $X=4.74 $Y=1.83 $X2=0
+ $Y2=0
cc_568 N_A_760_395#_c_600_n N_SET_B_c_826_n 0.00502262f $X=4.882 $Y=2.32 $X2=0
+ $Y2=0
cc_569 N_A_760_395#_M1030_g N_A_224_350#_M1015_g 0.0306235f $X=3.89 $Y=2.525
+ $X2=0 $Y2=0
cc_570 N_A_760_395#_M1030_g N_A_224_350#_c_954_n 0.0123711f $X=3.89 $Y=2.525
+ $X2=0 $Y2=0
cc_571 N_A_760_395#_M1030_g N_VPWR_c_1502_n 0.00782972f $X=3.89 $Y=2.525 $X2=0
+ $Y2=0
cc_572 N_A_760_395#_c_597_n N_VPWR_c_1502_n 0.00116235f $X=4.22 $Y=1.8 $X2=0
+ $Y2=0
cc_573 N_A_760_395#_M1030_g N_VPWR_c_1499_n 9.455e-19 $X=3.89 $Y=2.525 $X2=0
+ $Y2=0
cc_574 N_A_760_395#_c_590_n N_VGND_c_1657_n 0.011113f $X=4.015 $Y=0.9 $X2=0
+ $Y2=0
cc_575 N_A_760_395#_c_592_n N_VGND_c_1657_n 0.024793f $X=4.43 $Y=1.065 $X2=0
+ $Y2=0
cc_576 N_A_760_395#_c_593_n N_VGND_c_1657_n 0.00532336f $X=4.31 $Y=1.065 $X2=0
+ $Y2=0
cc_577 N_A_760_395#_c_592_n N_VGND_c_1658_n 0.0134505f $X=4.43 $Y=1.065 $X2=0
+ $Y2=0
cc_578 N_A_760_395#_c_592_n N_VGND_c_1660_n 0.00866682f $X=4.43 $Y=1.065 $X2=0
+ $Y2=0
cc_579 N_A_760_395#_c_590_n N_VGND_c_1665_n 0.00383152f $X=4.015 $Y=0.9 $X2=0
+ $Y2=0
cc_580 N_A_760_395#_c_590_n N_VGND_c_1667_n 0.00385559f $X=4.015 $Y=0.9 $X2=0
+ $Y2=0
cc_581 N_A_760_395#_c_592_n N_VGND_c_1667_n 0.0188048f $X=4.43 $Y=1.065 $X2=0
+ $Y2=0
cc_582 N_A_604_74#_M1001_g N_SET_B_M1012_g 0.0103384f $X=5.91 $Y=2.205 $X2=0
+ $Y2=0
cc_583 N_A_604_74#_M1011_g N_SET_B_M1009_g 0.0703762f $X=5.06 $Y=0.8 $X2=0 $Y2=0
cc_584 N_A_604_74#_M1001_g N_SET_B_M1009_g 0.0235368f $X=5.91 $Y=2.205 $X2=0
+ $Y2=0
cc_585 N_A_604_74#_M1003_g N_SET_B_M1009_g 0.0119302f $X=6 $Y=0.69 $X2=0 $Y2=0
cc_586 N_A_604_74#_c_677_n N_SET_B_M1009_g 0.0055839f $X=4.97 $Y=1.38 $X2=0
+ $Y2=0
cc_587 N_A_604_74#_c_678_n N_SET_B_M1009_g 0.0207669f $X=5.9 $Y=1.38 $X2=0 $Y2=0
cc_588 N_A_604_74#_c_679_n N_SET_B_M1009_g 0.0180957f $X=5.9 $Y=1.38 $X2=0 $Y2=0
cc_589 N_A_604_74#_M1001_g N_SET_B_c_822_n 0.00227463f $X=5.91 $Y=2.205 $X2=0
+ $Y2=0
cc_590 N_A_604_74#_c_678_n N_SET_B_c_822_n 0.0059453f $X=5.9 $Y=1.38 $X2=0 $Y2=0
cc_591 N_A_604_74#_c_679_n N_SET_B_c_822_n 0.00144973f $X=5.9 $Y=1.38 $X2=0
+ $Y2=0
cc_592 N_A_604_74#_c_678_n N_SET_B_c_823_n 0.00281639f $X=5.9 $Y=1.38 $X2=0
+ $Y2=0
cc_593 N_A_604_74#_M1000_g N_SET_B_c_824_n 3.47076e-19 $X=4.715 $Y=2.525 $X2=0
+ $Y2=0
cc_594 N_A_604_74#_M1001_g N_SET_B_c_824_n 0.00106128f $X=5.91 $Y=2.205 $X2=0
+ $Y2=0
cc_595 N_A_604_74#_c_677_n N_SET_B_c_824_n 2.37165e-19 $X=4.97 $Y=1.38 $X2=0
+ $Y2=0
cc_596 N_A_604_74#_c_678_n N_SET_B_c_824_n 0.0285069f $X=5.9 $Y=1.38 $X2=0 $Y2=0
cc_597 N_A_604_74#_M1000_g N_SET_B_c_826_n 0.0292523f $X=4.715 $Y=2.525 $X2=0
+ $Y2=0
cc_598 N_A_604_74#_c_677_n N_SET_B_c_826_n 0.00375465f $X=4.97 $Y=1.38 $X2=0
+ $Y2=0
cc_599 N_A_604_74#_c_678_n N_SET_B_c_826_n 0.00514762f $X=5.9 $Y=1.38 $X2=0
+ $Y2=0
cc_600 N_A_604_74#_c_672_n N_A_224_350#_M1013_g 0.00159443f $X=3.41 $Y=0.58
+ $X2=0 $Y2=0
cc_601 N_A_604_74#_c_680_n N_A_224_350#_M1013_g 5.73353e-19 $X=3.247 $Y=2.295
+ $X2=0 $Y2=0
cc_602 N_A_604_74#_c_681_n N_A_224_350#_M1013_g 6.98346e-19 $X=3.41 $Y=0.935
+ $X2=0 $Y2=0
cc_603 N_A_604_74#_c_688_n N_A_224_350#_M1015_g 0.00610386f $X=3.245 $Y=2.515
+ $X2=0 $Y2=0
cc_604 N_A_604_74#_c_680_n N_A_224_350#_M1015_g 0.00278796f $X=3.247 $Y=2.295
+ $X2=0 $Y2=0
cc_605 N_A_604_74#_M1000_g N_A_224_350#_c_954_n 0.0105864f $X=4.715 $Y=2.525
+ $X2=0 $Y2=0
cc_606 N_A_604_74#_M1001_g N_A_224_350#_c_954_n 0.010423f $X=5.91 $Y=2.205 $X2=0
+ $Y2=0
cc_607 N_A_604_74#_M1001_g N_A_224_350#_c_941_n 0.0433295f $X=5.91 $Y=2.205
+ $X2=0 $Y2=0
cc_608 N_A_604_74#_M1001_g N_A_1301_392#_c_1220_n 9.72093e-19 $X=5.91 $Y=2.205
+ $X2=0 $Y2=0
cc_609 N_A_604_74#_M1001_g N_A_1301_392#_c_1227_n 0.00190568f $X=5.91 $Y=2.205
+ $X2=0 $Y2=0
cc_610 N_A_604_74#_c_688_n N_A_27_74#_c_1440_n 0.0180198f $X=3.245 $Y=2.515
+ $X2=0 $Y2=0
cc_611 N_A_604_74#_c_680_n N_A_27_74#_c_1440_n 0.00645809f $X=3.247 $Y=2.295
+ $X2=0 $Y2=0
cc_612 N_A_604_74#_M1001_g N_VPWR_c_1503_n 0.00426431f $X=5.91 $Y=2.205 $X2=0
+ $Y2=0
cc_613 N_A_604_74#_M1001_g N_VPWR_c_1499_n 0.00113998f $X=5.91 $Y=2.205 $X2=0
+ $Y2=0
cc_614 N_A_604_74#_M1011_g N_VGND_c_1657_n 0.00308759f $X=5.06 $Y=0.8 $X2=0
+ $Y2=0
cc_615 N_A_604_74#_c_672_n N_VGND_c_1657_n 0.00850407f $X=3.41 $Y=0.58 $X2=0
+ $Y2=0
cc_616 N_A_604_74#_c_673_n N_VGND_c_1657_n 0.00216154f $X=3.925 $Y=0.935 $X2=0
+ $Y2=0
cc_617 N_A_604_74#_c_682_n N_VGND_c_1657_n 0.00420453f $X=4.805 $Y=1.38 $X2=0
+ $Y2=0
cc_618 N_A_604_74#_M1003_g N_VGND_c_1658_n 0.0140469f $X=6 $Y=0.69 $X2=0 $Y2=0
cc_619 N_A_604_74#_c_678_n N_VGND_c_1658_n 0.0263236f $X=5.9 $Y=1.38 $X2=0 $Y2=0
cc_620 N_A_604_74#_c_679_n N_VGND_c_1658_n 0.00480071f $X=5.9 $Y=1.38 $X2=0
+ $Y2=0
cc_621 N_A_604_74#_M1011_g N_VGND_c_1660_n 0.00416964f $X=5.06 $Y=0.8 $X2=0
+ $Y2=0
cc_622 N_A_604_74#_c_672_n N_VGND_c_1665_n 0.0102427f $X=3.41 $Y=0.58 $X2=0
+ $Y2=0
cc_623 N_A_604_74#_M1011_g N_VGND_c_1667_n 0.00479212f $X=5.06 $Y=0.8 $X2=0
+ $Y2=0
cc_624 N_A_604_74#_M1003_g N_VGND_c_1667_n 0.00758453f $X=6 $Y=0.69 $X2=0 $Y2=0
cc_625 N_A_604_74#_c_672_n N_VGND_c_1667_n 0.0114717f $X=3.41 $Y=0.58 $X2=0
+ $Y2=0
cc_626 N_A_604_74#_c_673_n N_VGND_c_1667_n 0.0156955f $X=3.925 $Y=0.935 $X2=0
+ $Y2=0
cc_627 N_A_604_74#_M1003_g N_VGND_c_1671_n 0.00383152f $X=6 $Y=0.69 $X2=0 $Y2=0
cc_628 N_SET_B_M1012_g N_A_224_350#_c_954_n 0.0109545f $X=5.165 $Y=2.525 $X2=0
+ $Y2=0
cc_629 N_SET_B_c_822_n N_A_224_350#_M1021_g 0.00930082f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_630 N_SET_B_c_822_n N_A_224_350#_c_940_n 0.00644007f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_631 N_SET_B_c_813_n N_A_1470_48#_M1019_g 0.0401587f $X=7.815 $Y=0.865 $X2=0
+ $Y2=0
cc_632 N_SET_B_c_814_n N_A_1470_48#_M1019_g 0.00361551f $X=8.267 $Y=1.377 $X2=0
+ $Y2=0
cc_633 N_SET_B_c_819_n N_A_1470_48#_M1002_g 0.0282631f $X=8.08 $Y=2.23 $X2=0
+ $Y2=0
cc_634 N_SET_B_c_815_n N_A_1470_48#_M1002_g 0.0264005f $X=8.267 $Y=1.893 $X2=0
+ $Y2=0
cc_635 N_SET_B_c_822_n N_A_1470_48#_M1002_g 0.00724986f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_636 N_SET_B_c_816_n N_A_1470_48#_M1002_g 0.00301488f $X=8.35 $Y=1.295 $X2=0
+ $Y2=0
cc_637 N_SET_B_c_814_n N_A_1470_48#_c_1122_n 0.00621167f $X=8.267 $Y=1.377 $X2=0
+ $Y2=0
cc_638 N_SET_B_c_822_n N_A_1470_48#_c_1122_n 0.00815716f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_639 N_SET_B_c_816_n N_A_1470_48#_c_1122_n 0.0143471f $X=8.35 $Y=1.295 $X2=0
+ $Y2=0
cc_640 N_SET_B_c_813_n N_A_1470_48#_c_1123_n 0.00667501f $X=7.815 $Y=0.865 $X2=0
+ $Y2=0
cc_641 N_SET_B_c_814_n N_A_1470_48#_c_1123_n 0.0300714f $X=8.267 $Y=1.377 $X2=0
+ $Y2=0
cc_642 N_SET_B_c_816_n N_A_1470_48#_c_1123_n 0.0262124f $X=8.35 $Y=1.295 $X2=0
+ $Y2=0
cc_643 N_SET_B_c_816_n N_A_1470_48#_c_1124_n 0.00221386f $X=8.35 $Y=1.295 $X2=0
+ $Y2=0
cc_644 N_SET_B_c_814_n N_A_1470_48#_c_1127_n 0.0216942f $X=8.267 $Y=1.377 $X2=0
+ $Y2=0
cc_645 N_SET_B_c_822_n N_A_1470_48#_c_1127_n 0.00460122f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_646 N_SET_B_c_816_n N_A_1470_48#_c_1127_n 0.00101327f $X=8.35 $Y=1.295 $X2=0
+ $Y2=0
cc_647 N_SET_B_c_822_n N_A_1301_392#_M1021_d 8.36767e-19 $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_648 N_SET_B_c_815_n N_A_1301_392#_c_1203_n 0.0127996f $X=8.267 $Y=1.893 $X2=0
+ $Y2=0
cc_649 N_SET_B_c_814_n N_A_1301_392#_M1005_g 0.0164387f $X=8.267 $Y=1.377 $X2=0
+ $Y2=0
cc_650 N_SET_B_c_816_n N_A_1301_392#_M1005_g 0.00132758f $X=8.35 $Y=1.295 $X2=0
+ $Y2=0
cc_651 N_SET_B_c_819_n N_A_1301_392#_c_1216_n 0.0127996f $X=8.08 $Y=2.23 $X2=0
+ $Y2=0
cc_652 SET_B N_A_1301_392#_c_1216_n 0.00406074f $X=8.315 $Y=1.95 $X2=0 $Y2=0
cc_653 N_SET_B_M1006_g N_A_1301_392#_c_1217_n 0.00230403f $X=8.08 $Y=2.75 $X2=0
+ $Y2=0
cc_654 N_SET_B_c_822_n N_A_1301_392#_c_1219_n 0.0111844f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_655 N_SET_B_M1006_g N_A_1301_392#_c_1221_n 4.33574e-19 $X=8.08 $Y=2.75 $X2=0
+ $Y2=0
cc_656 N_SET_B_M1006_g N_A_1301_392#_c_1222_n 0.0100857f $X=8.08 $Y=2.75 $X2=0
+ $Y2=0
cc_657 N_SET_B_c_822_n N_A_1301_392#_c_1222_n 0.0217589f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_658 N_SET_B_c_822_n N_A_1301_392#_c_1223_n 0.00816942f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_659 N_SET_B_M1006_g N_A_1301_392#_c_1224_n 0.00862157f $X=8.08 $Y=2.75 $X2=0
+ $Y2=0
cc_660 N_SET_B_c_819_n N_A_1301_392#_c_1225_n 3.03852e-19 $X=8.08 $Y=2.23 $X2=0
+ $Y2=0
cc_661 SET_B N_A_1301_392#_c_1225_n 0.00271215f $X=8.315 $Y=1.95 $X2=0 $Y2=0
cc_662 N_SET_B_c_816_n N_A_1301_392#_c_1225_n 0.00276823f $X=8.35 $Y=1.295 $X2=0
+ $Y2=0
cc_663 N_SET_B_c_819_n N_A_1301_392#_c_1207_n 8.5946e-19 $X=8.08 $Y=2.23 $X2=0
+ $Y2=0
cc_664 N_SET_B_c_814_n N_A_1301_392#_c_1207_n 0.00288794f $X=8.267 $Y=1.377
+ $X2=0 $Y2=0
cc_665 SET_B N_A_1301_392#_c_1207_n 0.00719608f $X=8.315 $Y=1.95 $X2=0 $Y2=0
cc_666 N_SET_B_c_816_n N_A_1301_392#_c_1207_n 0.0377878f $X=8.35 $Y=1.295 $X2=0
+ $Y2=0
cc_667 N_SET_B_c_814_n N_A_1301_392#_c_1208_n 0.0127996f $X=8.267 $Y=1.377 $X2=0
+ $Y2=0
cc_668 N_SET_B_c_816_n N_A_1301_392#_c_1208_n 0.00318354f $X=8.35 $Y=1.295 $X2=0
+ $Y2=0
cc_669 N_SET_B_c_819_n N_A_1301_392#_c_1226_n 0.00230403f $X=8.08 $Y=2.23 $X2=0
+ $Y2=0
cc_670 N_SET_B_c_822_n N_A_1301_392#_c_1227_n 0.022804f $X=8.255 $Y=2.035 $X2=0
+ $Y2=0
cc_671 N_SET_B_c_822_n N_A_1301_392#_c_1228_n 0.00766188f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_672 N_SET_B_c_822_n N_A_1301_392#_c_1210_n 0.00844252f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_673 N_SET_B_c_819_n N_A_1301_392#_c_1229_n 0.00295338f $X=8.08 $Y=2.23 $X2=0
+ $Y2=0
cc_674 N_SET_B_M1006_g N_A_1301_392#_c_1229_n 0.00480662f $X=8.08 $Y=2.75 $X2=0
+ $Y2=0
cc_675 N_SET_B_c_822_n N_A_1301_392#_c_1229_n 0.00256403f $X=8.255 $Y=2.035
+ $X2=0 $Y2=0
cc_676 SET_B N_A_1301_392#_c_1229_n 0.00615918f $X=8.315 $Y=1.95 $X2=0 $Y2=0
cc_677 N_SET_B_c_816_n N_A_1301_392#_c_1229_n 0.0207551f $X=8.35 $Y=1.295 $X2=0
+ $Y2=0
cc_678 N_SET_B_c_822_n N_VPWR_M1012_d 0.0026243f $X=8.255 $Y=2.035 $X2=0 $Y2=0
cc_679 N_SET_B_c_823_n N_VPWR_M1012_d 0.00184407f $X=5.665 $Y=2.035 $X2=0 $Y2=0
cc_680 N_SET_B_c_824_n N_VPWR_M1012_d 0.00313128f $X=5.52 $Y=2.035 $X2=0 $Y2=0
cc_681 N_SET_B_M1012_g N_VPWR_c_1503_n 7.14396e-19 $X=5.165 $Y=2.525 $X2=0 $Y2=0
cc_682 N_SET_B_M1006_g N_VPWR_c_1504_n 0.00308998f $X=8.08 $Y=2.75 $X2=0 $Y2=0
cc_683 N_SET_B_M1006_g N_VPWR_c_1505_n 0.00373364f $X=8.08 $Y=2.75 $X2=0 $Y2=0
cc_684 N_SET_B_M1006_g N_VPWR_c_1514_n 0.00522185f $X=8.08 $Y=2.75 $X2=0 $Y2=0
cc_685 N_SET_B_M1006_g N_VPWR_c_1499_n 0.0054187f $X=8.08 $Y=2.75 $X2=0 $Y2=0
cc_686 N_SET_B_c_822_n A_1200_341# 0.0150735f $X=8.255 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_687 N_SET_B_M1009_g N_VGND_c_1658_n 0.00920042f $X=5.42 $Y=0.8 $X2=0 $Y2=0
cc_688 N_SET_B_M1009_g N_VGND_c_1660_n 0.00434252f $X=5.42 $Y=0.8 $X2=0 $Y2=0
cc_689 N_SET_B_M1009_g N_VGND_c_1667_n 0.00479212f $X=5.42 $Y=0.8 $X2=0 $Y2=0
cc_690 N_SET_B_c_813_n N_VGND_c_1667_n 0.00386373f $X=7.815 $Y=0.865 $X2=0 $Y2=0
cc_691 N_SET_B_c_813_n N_VGND_c_1671_n 0.00398535f $X=7.815 $Y=0.865 $X2=0 $Y2=0
cc_692 N_SET_B_c_813_n N_VGND_c_1672_n 0.0100278f $X=7.815 $Y=0.865 $X2=0 $Y2=0
cc_693 N_SET_B_c_814_n N_VGND_c_1672_n 0.00165348f $X=8.267 $Y=1.377 $X2=0 $Y2=0
cc_694 N_A_224_350#_M1018_g N_A_1470_48#_M1019_g 0.0593492f $X=7.035 $Y=0.58
+ $X2=0 $Y2=0
cc_695 N_A_224_350#_M1018_g N_A_1470_48#_M1002_g 0.00524446f $X=7.035 $Y=0.58
+ $X2=0 $Y2=0
cc_696 N_A_224_350#_M1021_g N_A_1301_392#_c_1218_n 0.00763701f $X=6.415 $Y=2.46
+ $X2=0 $Y2=0
cc_697 N_A_224_350#_M1021_g N_A_1301_392#_c_1220_n 0.012215f $X=6.415 $Y=2.46
+ $X2=0 $Y2=0
cc_698 N_A_224_350#_c_940_n N_A_1301_392#_c_1206_n 0.00172054f $X=6.96 $Y=1.735
+ $X2=0 $Y2=0
cc_699 N_A_224_350#_M1018_g N_A_1301_392#_c_1206_n 0.0148711f $X=7.035 $Y=0.58
+ $X2=0 $Y2=0
cc_700 N_A_224_350#_M1021_g N_A_1301_392#_c_1227_n 0.00326666f $X=6.415 $Y=2.46
+ $X2=0 $Y2=0
cc_701 N_A_224_350#_c_940_n N_A_1301_392#_c_1227_n 0.00129944f $X=6.96 $Y=1.735
+ $X2=0 $Y2=0
cc_702 N_A_224_350#_M1021_g N_A_1301_392#_c_1228_n 0.00440451f $X=6.415 $Y=2.46
+ $X2=0 $Y2=0
cc_703 N_A_224_350#_c_940_n N_A_1301_392#_c_1228_n 0.00685526f $X=6.96 $Y=1.735
+ $X2=0 $Y2=0
cc_704 N_A_224_350#_M1018_g N_A_1301_392#_c_1209_n 0.00842127f $X=7.035 $Y=0.58
+ $X2=0 $Y2=0
cc_705 N_A_224_350#_c_940_n N_A_1301_392#_c_1210_n 0.0155681f $X=6.96 $Y=1.735
+ $X2=0 $Y2=0
cc_706 N_A_224_350#_M1018_g N_A_1301_392#_c_1210_n 9.65332e-19 $X=7.035 $Y=0.58
+ $X2=0 $Y2=0
cc_707 N_A_224_350#_M1004_s N_A_27_74#_c_1439_n 0.0112096f $X=1.12 $Y=1.75 $X2=0
+ $Y2=0
cc_708 N_A_224_350#_c_963_n N_A_27_74#_c_1439_n 0.00581391f $X=1.985 $Y=1.805
+ $X2=0 $Y2=0
cc_709 N_A_224_350#_c_965_n N_A_27_74#_c_1439_n 0.0299077f $X=1.42 $Y=1.89 $X2=0
+ $Y2=0
cc_710 N_A_224_350#_M1010_g N_A_27_74#_c_1440_n 0.0167256f $X=1.93 $Y=2.31 $X2=0
+ $Y2=0
cc_711 N_A_224_350#_c_950_n N_A_27_74#_c_1440_n 0.028461f $X=2.45 $Y=3.075 $X2=0
+ $Y2=0
cc_712 N_A_224_350#_c_944_n N_A_27_74#_c_1440_n 6.39267e-19 $X=2.375 $Y=1.425
+ $X2=0 $Y2=0
cc_713 N_A_224_350#_c_963_n N_A_27_74#_c_1440_n 0.033362f $X=1.985 $Y=1.805
+ $X2=0 $Y2=0
cc_714 N_A_224_350#_M1020_g N_A_27_74#_c_1434_n 7.64769e-19 $X=1.915 $Y=0.74
+ $X2=0 $Y2=0
cc_715 N_A_224_350#_M1010_g N_A_27_74#_c_1434_n 0.00106311f $X=1.93 $Y=2.31
+ $X2=0 $Y2=0
cc_716 N_A_224_350#_c_950_n N_A_27_74#_c_1434_n 0.00970648f $X=2.45 $Y=3.075
+ $X2=0 $Y2=0
cc_717 N_A_224_350#_c_938_n N_A_27_74#_c_1434_n 0.0105124f $X=2.87 $Y=1.12 $X2=0
+ $Y2=0
cc_718 N_A_224_350#_M1013_g N_A_27_74#_c_1434_n 0.00226525f $X=2.945 $Y=0.58
+ $X2=0 $Y2=0
cc_719 N_A_224_350#_c_945_n N_A_27_74#_c_1434_n 0.0140574f $X=2.45 $Y=1.317
+ $X2=0 $Y2=0
cc_720 N_A_224_350#_c_963_n N_A_27_74#_c_1434_n 0.0137401f $X=1.985 $Y=1.805
+ $X2=0 $Y2=0
cc_721 N_A_224_350#_c_947_n N_A_27_74#_c_1434_n 0.0333747f $X=2.15 $Y=1.425
+ $X2=0 $Y2=0
cc_722 N_A_224_350#_M1010_g N_A_27_74#_c_1482_n 0.00422161f $X=1.93 $Y=2.31
+ $X2=0 $Y2=0
cc_723 N_A_224_350#_c_963_n N_A_27_74#_c_1482_n 0.0101605f $X=1.985 $Y=1.805
+ $X2=0 $Y2=0
cc_724 N_A_224_350#_M1020_g N_A_27_74#_c_1436_n 6.88372e-19 $X=1.915 $Y=0.74
+ $X2=0 $Y2=0
cc_725 N_A_224_350#_c_938_n N_A_27_74#_c_1436_n 0.00290347f $X=2.87 $Y=1.12
+ $X2=0 $Y2=0
cc_726 N_A_224_350#_M1013_g N_A_27_74#_c_1436_n 0.00664053f $X=2.945 $Y=0.58
+ $X2=0 $Y2=0
cc_727 N_A_224_350#_c_963_n N_VPWR_M1004_d 0.00164828f $X=1.985 $Y=1.805 $X2=0
+ $Y2=0
cc_728 N_A_224_350#_M1010_g N_VPWR_c_1501_n 0.00786063f $X=1.93 $Y=2.31 $X2=0
+ $Y2=0
cc_729 N_A_224_350#_c_950_n N_VPWR_c_1501_n 4.3464e-19 $X=2.45 $Y=3.075 $X2=0
+ $Y2=0
cc_730 N_A_224_350#_c_952_n N_VPWR_c_1501_n 0.00272925f $X=2.525 $Y=3.15 $X2=0
+ $Y2=0
cc_731 N_A_224_350#_M1015_g N_VPWR_c_1502_n 8.75021e-19 $X=3.47 $Y=2.525 $X2=0
+ $Y2=0
cc_732 N_A_224_350#_c_954_n N_VPWR_c_1502_n 0.0227567f $X=6.325 $Y=3.15 $X2=0
+ $Y2=0
cc_733 N_A_224_350#_c_954_n N_VPWR_c_1503_n 0.021028f $X=6.325 $Y=3.15 $X2=0
+ $Y2=0
cc_734 N_A_224_350#_M1021_g N_VPWR_c_1503_n 0.00630945f $X=6.415 $Y=2.46 $X2=0
+ $Y2=0
cc_735 N_A_224_350#_c_954_n N_VPWR_c_1507_n 0.0313883f $X=6.325 $Y=3.15 $X2=0
+ $Y2=0
cc_736 N_A_224_350#_c_954_n N_VPWR_c_1509_n 0.0259651f $X=6.325 $Y=3.15 $X2=0
+ $Y2=0
cc_737 N_A_224_350#_M1010_g N_VPWR_c_1513_n 0.00512593f $X=1.93 $Y=2.31 $X2=0
+ $Y2=0
cc_738 N_A_224_350#_c_952_n N_VPWR_c_1513_n 0.0368171f $X=2.525 $Y=3.15 $X2=0
+ $Y2=0
cc_739 N_A_224_350#_M1010_g N_VPWR_c_1499_n 0.00520946f $X=1.93 $Y=2.31 $X2=0
+ $Y2=0
cc_740 N_A_224_350#_c_951_n N_VPWR_c_1499_n 0.0201297f $X=3.38 $Y=3.15 $X2=0
+ $Y2=0
cc_741 N_A_224_350#_c_952_n N_VPWR_c_1499_n 0.00604517f $X=2.525 $Y=3.15 $X2=0
+ $Y2=0
cc_742 N_A_224_350#_c_954_n N_VPWR_c_1499_n 0.0848882f $X=6.325 $Y=3.15 $X2=0
+ $Y2=0
cc_743 N_A_224_350#_c_961_n N_VPWR_c_1499_n 0.00445015f $X=3.47 $Y=3.15 $X2=0
+ $Y2=0
cc_744 N_A_224_350#_c_948_n N_VGND_c_1654_n 0.0363632f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_745 N_A_224_350#_c_948_n N_VGND_c_1655_n 0.0203368f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_746 N_A_224_350#_M1020_g N_VGND_c_1656_n 0.00115634f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_747 N_A_224_350#_c_948_n N_VGND_c_1656_n 0.0255747f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_748 N_A_224_350#_M1020_g N_VGND_c_1665_n 0.00430908f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_749 N_A_224_350#_M1013_g N_VGND_c_1665_n 0.00278159f $X=2.945 $Y=0.58 $X2=0
+ $Y2=0
cc_750 N_A_224_350#_M1020_g N_VGND_c_1667_n 0.00820779f $X=1.915 $Y=0.74 $X2=0
+ $Y2=0
cc_751 N_A_224_350#_M1013_g N_VGND_c_1667_n 0.00360393f $X=2.945 $Y=0.58 $X2=0
+ $Y2=0
cc_752 N_A_224_350#_M1018_g N_VGND_c_1667_n 0.00353931f $X=7.035 $Y=0.58 $X2=0
+ $Y2=0
cc_753 N_A_224_350#_c_948_n N_VGND_c_1667_n 0.0167889f $X=1.27 $Y=0.515 $X2=0
+ $Y2=0
cc_754 N_A_224_350#_M1018_g N_VGND_c_1671_n 0.00278271f $X=7.035 $Y=0.58 $X2=0
+ $Y2=0
cc_755 N_A_1470_48#_c_1123_n N_A_1301_392#_M1005_g 0.0110779f $X=8.93 $Y=0.875
+ $X2=0 $Y2=0
cc_756 N_A_1470_48#_c_1124_n N_A_1301_392#_M1005_g 0.0125588f $X=9.095 $Y=0.79
+ $X2=0 $Y2=0
cc_757 N_A_1470_48#_c_1125_n N_A_1301_392#_M1005_g 0.0121111f $X=9.095 $Y=0.58
+ $X2=0 $Y2=0
cc_758 N_A_1470_48#_c_1126_n N_A_1301_392#_M1005_g 0.00348663f $X=9.28 $Y=2.65
+ $X2=0 $Y2=0
cc_759 N_A_1470_48#_c_1129_n N_A_1301_392#_M1016_g 0.00604419f $X=9.28 $Y=2.815
+ $X2=0 $Y2=0
cc_760 N_A_1470_48#_c_1124_n N_A_1301_392#_c_1213_n 0.00179394f $X=9.095 $Y=0.79
+ $X2=0 $Y2=0
cc_761 N_A_1470_48#_c_1126_n N_A_1301_392#_c_1213_n 0.0146955f $X=9.28 $Y=2.65
+ $X2=0 $Y2=0
cc_762 N_A_1470_48#_c_1124_n N_A_1301_392#_M1026_g 0.0020199f $X=9.095 $Y=0.79
+ $X2=0 $Y2=0
cc_763 N_A_1470_48#_c_1125_n N_A_1301_392#_M1026_g 8.93332e-19 $X=9.095 $Y=0.58
+ $X2=0 $Y2=0
cc_764 N_A_1470_48#_c_1126_n N_A_1301_392#_M1026_g 0.00206229f $X=9.28 $Y=2.65
+ $X2=0 $Y2=0
cc_765 N_A_1470_48#_c_1129_n N_A_1301_392#_c_1215_n 0.00283772f $X=9.28 $Y=2.815
+ $X2=0 $Y2=0
cc_766 N_A_1470_48#_c_1126_n N_A_1301_392#_c_1215_n 0.00193182f $X=9.28 $Y=2.65
+ $X2=0 $Y2=0
cc_767 N_A_1470_48#_c_1126_n N_A_1301_392#_c_1217_n 0.0100461f $X=9.28 $Y=2.65
+ $X2=0 $Y2=0
cc_768 N_A_1470_48#_M1002_g N_A_1301_392#_c_1219_n 0.00915692f $X=7.63 $Y=2.75
+ $X2=0 $Y2=0
cc_769 N_A_1470_48#_M1002_g N_A_1301_392#_c_1221_n 0.00374628f $X=7.63 $Y=2.75
+ $X2=0 $Y2=0
cc_770 N_A_1470_48#_M1002_g N_A_1301_392#_c_1222_n 0.00848754f $X=7.63 $Y=2.75
+ $X2=0 $Y2=0
cc_771 N_A_1470_48#_M1002_g N_A_1301_392#_c_1223_n 0.00301525f $X=7.63 $Y=2.75
+ $X2=0 $Y2=0
cc_772 N_A_1470_48#_M1002_g N_A_1301_392#_c_1224_n 5.14899e-19 $X=7.63 $Y=2.75
+ $X2=0 $Y2=0
cc_773 N_A_1470_48#_c_1126_n N_A_1301_392#_c_1225_n 0.0135429f $X=9.28 $Y=2.65
+ $X2=0 $Y2=0
cc_774 N_A_1470_48#_c_1123_n N_A_1301_392#_c_1207_n 0.0058457f $X=8.93 $Y=0.875
+ $X2=0 $Y2=0
cc_775 N_A_1470_48#_c_1124_n N_A_1301_392#_c_1207_n 0.00843598f $X=9.095 $Y=0.79
+ $X2=0 $Y2=0
cc_776 N_A_1470_48#_c_1126_n N_A_1301_392#_c_1207_n 0.069897f $X=9.28 $Y=2.65
+ $X2=0 $Y2=0
cc_777 N_A_1470_48#_c_1124_n N_A_1301_392#_c_1208_n 0.0015596f $X=9.095 $Y=0.79
+ $X2=0 $Y2=0
cc_778 N_A_1470_48#_c_1126_n N_A_1301_392#_c_1208_n 0.00453092f $X=9.28 $Y=2.65
+ $X2=0 $Y2=0
cc_779 N_A_1470_48#_c_1126_n N_A_1301_392#_c_1226_n 0.00657792f $X=9.28 $Y=2.65
+ $X2=0 $Y2=0
cc_780 N_A_1470_48#_c_1125_n N_A_1902_74#_c_1378_n 0.0295967f $X=9.095 $Y=0.58
+ $X2=0 $Y2=0
cc_781 N_A_1470_48#_c_1124_n N_A_1902_74#_c_1379_n 0.0205377f $X=9.095 $Y=0.79
+ $X2=0 $Y2=0
cc_782 N_A_1470_48#_c_1126_n N_A_1902_74#_c_1379_n 0.00148628f $X=9.28 $Y=2.65
+ $X2=0 $Y2=0
cc_783 N_A_1470_48#_c_1126_n N_A_1902_74#_c_1380_n 0.0971011f $X=9.28 $Y=2.65
+ $X2=0 $Y2=0
cc_784 N_A_1470_48#_c_1124_n N_A_1902_74#_c_1382_n 0.00500774f $X=9.095 $Y=0.79
+ $X2=0 $Y2=0
cc_785 N_A_1470_48#_c_1126_n N_A_1902_74#_c_1383_n 0.0260062f $X=9.28 $Y=2.65
+ $X2=0 $Y2=0
cc_786 N_A_1470_48#_M1002_g N_VPWR_c_1504_n 0.00276751f $X=7.63 $Y=2.75 $X2=0
+ $Y2=0
cc_787 N_A_1470_48#_c_1129_n N_VPWR_c_1505_n 0.011548f $X=9.28 $Y=2.815 $X2=0
+ $Y2=0
cc_788 N_A_1470_48#_M1002_g N_VPWR_c_1509_n 0.00485777f $X=7.63 $Y=2.75 $X2=0
+ $Y2=0
cc_789 N_A_1470_48#_c_1129_n N_VPWR_c_1515_n 0.0142018f $X=9.28 $Y=2.815 $X2=0
+ $Y2=0
cc_790 N_A_1470_48#_M1002_g N_VPWR_c_1499_n 0.00514672f $X=7.63 $Y=2.75 $X2=0
+ $Y2=0
cc_791 N_A_1470_48#_c_1129_n N_VPWR_c_1499_n 0.0118394f $X=9.28 $Y=2.815 $X2=0
+ $Y2=0
cc_792 N_A_1470_48#_c_1125_n N_VGND_c_1662_n 0.0145091f $X=9.095 $Y=0.58 $X2=0
+ $Y2=0
cc_793 N_A_1470_48#_M1019_g N_VGND_c_1667_n 0.00893489f $X=7.425 $Y=0.58 $X2=0
+ $Y2=0
cc_794 N_A_1470_48#_c_1123_n N_VGND_c_1667_n 0.0125427f $X=8.93 $Y=0.875 $X2=0
+ $Y2=0
cc_795 N_A_1470_48#_c_1137_n N_VGND_c_1667_n 0.00964541f $X=7.73 $Y=0.875 $X2=0
+ $Y2=0
cc_796 N_A_1470_48#_c_1125_n N_VGND_c_1667_n 0.0119768f $X=9.095 $Y=0.58 $X2=0
+ $Y2=0
cc_797 N_A_1470_48#_M1019_g N_VGND_c_1671_n 0.00461464f $X=7.425 $Y=0.58 $X2=0
+ $Y2=0
cc_798 N_A_1470_48#_M1019_g N_VGND_c_1672_n 0.00107631f $X=7.425 $Y=0.58 $X2=0
+ $Y2=0
cc_799 N_A_1470_48#_c_1123_n N_VGND_c_1672_n 0.0621318f $X=8.93 $Y=0.875 $X2=0
+ $Y2=0
cc_800 N_A_1470_48#_c_1125_n N_VGND_c_1672_n 0.0102732f $X=9.095 $Y=0.58 $X2=0
+ $Y2=0
cc_801 N_A_1470_48#_c_1137_n A_1500_74# 0.00522679f $X=7.73 $Y=0.875 $X2=-0.19
+ $Y2=-0.245
cc_802 N_A_1301_392#_M1026_g N_A_1902_74#_c_1376_n 0.0199795f $X=9.87 $Y=0.645
+ $X2=0 $Y2=0
cc_803 N_A_1301_392#_M1026_g N_A_1902_74#_M1025_g 0.0044545f $X=9.87 $Y=0.645
+ $X2=0 $Y2=0
cc_804 N_A_1301_392#_c_1215_n N_A_1902_74#_M1025_g 0.0188779f $X=10.025 $Y=1.94
+ $X2=0 $Y2=0
cc_805 N_A_1301_392#_M1005_g N_A_1902_74#_c_1378_n 0.00115501f $X=8.88 $Y=0.58
+ $X2=0 $Y2=0
cc_806 N_A_1301_392#_M1026_g N_A_1902_74#_c_1378_n 0.00508808f $X=9.87 $Y=0.645
+ $X2=0 $Y2=0
cc_807 N_A_1301_392#_M1005_g N_A_1902_74#_c_1379_n 8.78745e-19 $X=8.88 $Y=0.58
+ $X2=0 $Y2=0
cc_808 N_A_1301_392#_M1026_g N_A_1902_74#_c_1379_n 0.0117529f $X=9.87 $Y=0.645
+ $X2=0 $Y2=0
cc_809 N_A_1301_392#_M1016_g N_A_1902_74#_c_1380_n 9.10639e-19 $X=9.055 $Y=2.75
+ $X2=0 $Y2=0
cc_810 N_A_1301_392#_c_1213_n N_A_1902_74#_c_1380_n 0.0100324f $X=9.795 $Y=1.865
+ $X2=0 $Y2=0
cc_811 N_A_1301_392#_M1026_g N_A_1902_74#_c_1380_n 0.00856752f $X=9.87 $Y=0.645
+ $X2=0 $Y2=0
cc_812 N_A_1301_392#_c_1215_n N_A_1902_74#_c_1380_n 0.0221494f $X=10.025 $Y=1.94
+ $X2=0 $Y2=0
cc_813 N_A_1301_392#_c_1215_n N_A_1902_74#_c_1381_n 0.00615405f $X=10.025
+ $Y=1.94 $X2=0 $Y2=0
cc_814 N_A_1301_392#_M1026_g N_A_1902_74#_c_1382_n 0.0029603f $X=9.87 $Y=0.645
+ $X2=0 $Y2=0
cc_815 N_A_1301_392#_M1005_g N_A_1902_74#_c_1383_n 5.05055e-19 $X=8.88 $Y=0.58
+ $X2=0 $Y2=0
cc_816 N_A_1301_392#_M1026_g N_A_1902_74#_c_1383_n 0.0196766f $X=9.87 $Y=0.645
+ $X2=0 $Y2=0
cc_817 N_A_1301_392#_M1026_g N_A_1902_74#_c_1384_n 0.0181207f $X=9.87 $Y=0.645
+ $X2=0 $Y2=0
cc_818 N_A_1301_392#_c_1219_n N_VPWR_c_1504_n 0.0146188f $X=7.43 $Y=2.802 $X2=0
+ $Y2=0
cc_819 N_A_1301_392#_c_1222_n N_VPWR_c_1504_n 0.0126397f $X=8.14 $Y=2.395 $X2=0
+ $Y2=0
cc_820 N_A_1301_392#_M1016_g N_VPWR_c_1505_n 0.00501904f $X=9.055 $Y=2.75 $X2=0
+ $Y2=0
cc_821 N_A_1301_392#_c_1217_n N_VPWR_c_1505_n 8.30109e-19 $X=8.96 $Y=2.38 $X2=0
+ $Y2=0
cc_822 N_A_1301_392#_c_1224_n N_VPWR_c_1505_n 0.0207365f $X=8.305 $Y=2.765 $X2=0
+ $Y2=0
cc_823 N_A_1301_392#_c_1225_n N_VPWR_c_1505_n 0.0210492f $X=8.775 $Y=2.395 $X2=0
+ $Y2=0
cc_824 N_A_1301_392#_c_1215_n N_VPWR_c_1506_n 0.00982233f $X=10.025 $Y=1.94
+ $X2=0 $Y2=0
cc_825 N_A_1301_392#_c_1219_n N_VPWR_c_1509_n 0.0331655f $X=7.43 $Y=2.802 $X2=0
+ $Y2=0
cc_826 N_A_1301_392#_c_1220_n N_VPWR_c_1509_n 0.0148583f $X=6.81 $Y=2.802 $X2=0
+ $Y2=0
cc_827 N_A_1301_392#_c_1224_n N_VPWR_c_1514_n 0.0107747f $X=8.305 $Y=2.765 $X2=0
+ $Y2=0
cc_828 N_A_1301_392#_M1016_g N_VPWR_c_1515_n 0.005209f $X=9.055 $Y=2.75 $X2=0
+ $Y2=0
cc_829 N_A_1301_392#_c_1215_n N_VPWR_c_1515_n 0.00578748f $X=10.025 $Y=1.94
+ $X2=0 $Y2=0
cc_830 N_A_1301_392#_M1016_g N_VPWR_c_1499_n 0.00579542f $X=9.055 $Y=2.75 $X2=0
+ $Y2=0
cc_831 N_A_1301_392#_c_1215_n N_VPWR_c_1499_n 0.00615499f $X=10.025 $Y=1.94
+ $X2=0 $Y2=0
cc_832 N_A_1301_392#_c_1219_n N_VPWR_c_1499_n 0.0275119f $X=7.43 $Y=2.802 $X2=0
+ $Y2=0
cc_833 N_A_1301_392#_c_1220_n N_VPWR_c_1499_n 0.012228f $X=6.81 $Y=2.802 $X2=0
+ $Y2=0
cc_834 N_A_1301_392#_c_1222_n N_VPWR_c_1499_n 0.0113201f $X=8.14 $Y=2.395 $X2=0
+ $Y2=0
cc_835 N_A_1301_392#_c_1224_n N_VPWR_c_1499_n 0.0115466f $X=8.305 $Y=2.765 $X2=0
+ $Y2=0
cc_836 N_A_1301_392#_c_1225_n N_VPWR_c_1499_n 0.0139296f $X=8.775 $Y=2.395 $X2=0
+ $Y2=0
cc_837 N_A_1301_392#_c_1219_n A_1460_508# 0.0014794f $X=7.43 $Y=2.802 $X2=-0.19
+ $Y2=-0.245
cc_838 N_A_1301_392#_c_1221_n A_1460_508# 0.00111868f $X=7.515 $Y=2.625
+ $X2=-0.19 $Y2=-0.245
cc_839 N_A_1301_392#_M1026_g N_Q_c_1638_n 2.21498e-19 $X=9.87 $Y=0.645 $X2=0
+ $Y2=0
cc_840 N_A_1301_392#_M1026_g N_VGND_c_1659_n 0.00772158f $X=9.87 $Y=0.645 $X2=0
+ $Y2=0
cc_841 N_A_1301_392#_M1005_g N_VGND_c_1662_n 0.00434272f $X=8.88 $Y=0.58 $X2=0
+ $Y2=0
cc_842 N_A_1301_392#_M1026_g N_VGND_c_1662_n 0.00434272f $X=9.87 $Y=0.645 $X2=0
+ $Y2=0
cc_843 N_A_1301_392#_M1005_g N_VGND_c_1667_n 0.00444404f $X=8.88 $Y=0.58 $X2=0
+ $Y2=0
cc_844 N_A_1301_392#_M1026_g N_VGND_c_1667_n 0.00826607f $X=9.87 $Y=0.645 $X2=0
+ $Y2=0
cc_845 N_A_1301_392#_M1005_g N_VGND_c_1672_n 0.010036f $X=8.88 $Y=0.58 $X2=0
+ $Y2=0
cc_846 N_A_1902_74#_M1025_g N_VPWR_c_1506_n 0.0236266f $X=10.545 $Y=2.4 $X2=0
+ $Y2=0
cc_847 N_A_1902_74#_c_1380_n N_VPWR_c_1506_n 0.0443705f $X=9.8 $Y=2.16 $X2=0
+ $Y2=0
cc_848 N_A_1902_74#_c_1381_n N_VPWR_c_1506_n 0.0195859f $X=10.35 $Y=1.385 $X2=0
+ $Y2=0
cc_849 N_A_1902_74#_c_1384_n N_VPWR_c_1506_n 0.00623155f $X=10.545 $Y=1.385
+ $X2=0 $Y2=0
cc_850 N_A_1902_74#_c_1380_n N_VPWR_c_1515_n 0.0101861f $X=9.8 $Y=2.16 $X2=0
+ $Y2=0
cc_851 N_A_1902_74#_M1025_g N_VPWR_c_1516_n 0.00460063f $X=10.545 $Y=2.4 $X2=0
+ $Y2=0
cc_852 N_A_1902_74#_M1025_g N_VPWR_c_1499_n 0.00912261f $X=10.545 $Y=2.4 $X2=0
+ $Y2=0
cc_853 N_A_1902_74#_c_1380_n N_VPWR_c_1499_n 0.0112917f $X=9.8 $Y=2.16 $X2=0
+ $Y2=0
cc_854 N_A_1902_74#_c_1376_n Q 0.0031284f $X=10.45 $Y=1.22 $X2=0 $Y2=0
cc_855 N_A_1902_74#_c_1381_n Q 0.00112015f $X=10.35 $Y=1.385 $X2=0 $Y2=0
cc_856 N_A_1902_74#_c_1384_n Q 0.0039352f $X=10.545 $Y=1.385 $X2=0 $Y2=0
cc_857 N_A_1902_74#_c_1376_n Q 0.00561171f $X=10.45 $Y=1.22 $X2=0 $Y2=0
cc_858 N_A_1902_74#_c_1381_n Q 0.0269563f $X=10.35 $Y=1.385 $X2=0 $Y2=0
cc_859 N_A_1902_74#_c_1384_n Q 0.0223867f $X=10.545 $Y=1.385 $X2=0 $Y2=0
cc_860 N_A_1902_74#_c_1376_n N_Q_c_1638_n 0.00562579f $X=10.45 $Y=1.22 $X2=0
+ $Y2=0
cc_861 N_A_1902_74#_c_1376_n N_VGND_c_1659_n 0.00747356f $X=10.45 $Y=1.22 $X2=0
+ $Y2=0
cc_862 N_A_1902_74#_c_1378_n N_VGND_c_1659_n 0.0289005f $X=9.655 $Y=0.605 $X2=0
+ $Y2=0
cc_863 N_A_1902_74#_c_1381_n N_VGND_c_1659_n 0.0252022f $X=10.35 $Y=1.385 $X2=0
+ $Y2=0
cc_864 N_A_1902_74#_c_1384_n N_VGND_c_1659_n 0.00328533f $X=10.545 $Y=1.385
+ $X2=0 $Y2=0
cc_865 N_A_1902_74#_c_1378_n N_VGND_c_1662_n 0.0144316f $X=9.655 $Y=0.605 $X2=0
+ $Y2=0
cc_866 N_A_1902_74#_c_1376_n N_VGND_c_1666_n 0.00434272f $X=10.45 $Y=1.22 $X2=0
+ $Y2=0
cc_867 N_A_1902_74#_c_1376_n N_VGND_c_1667_n 0.00825325f $X=10.45 $Y=1.22 $X2=0
+ $Y2=0
cc_868 N_A_1902_74#_c_1378_n N_VGND_c_1667_n 0.0119474f $X=9.655 $Y=0.605 $X2=0
+ $Y2=0
cc_869 N_A_27_74#_c_1440_n N_VPWR_M1004_d 9.92177e-19 $X=2.485 $Y=2.145 $X2=0
+ $Y2=0
cc_870 N_A_27_74#_c_1482_n N_VPWR_M1004_d 0.0051214f $X=1.675 $Y=2.145 $X2=0
+ $Y2=0
cc_871 N_A_27_74#_c_1438_n N_VPWR_c_1500_n 0.0141836f $X=0.27 $Y=2.75 $X2=0
+ $Y2=0
cc_872 N_A_27_74#_c_1439_n N_VPWR_c_1500_n 0.0244352f $X=1.59 $Y=2.315 $X2=0
+ $Y2=0
cc_873 N_A_27_74#_c_1439_n N_VPWR_c_1501_n 0.00216696f $X=1.59 $Y=2.315 $X2=0
+ $Y2=0
cc_874 N_A_27_74#_c_1440_n N_VPWR_c_1501_n 0.00236221f $X=2.485 $Y=2.145 $X2=0
+ $Y2=0
cc_875 N_A_27_74#_c_1482_n N_VPWR_c_1501_n 0.01132f $X=1.675 $Y=2.145 $X2=0
+ $Y2=0
cc_876 N_A_27_74#_c_1438_n N_VPWR_c_1511_n 0.011066f $X=0.27 $Y=2.75 $X2=0 $Y2=0
cc_877 N_A_27_74#_c_1438_n N_VPWR_c_1499_n 0.00915947f $X=0.27 $Y=2.75 $X2=0
+ $Y2=0
cc_878 N_A_27_74#_c_1432_n N_VGND_c_1654_n 0.0172649f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_879 N_A_27_74#_c_1432_n N_VGND_c_1664_n 0.011402f $X=0.28 $Y=0.58 $X2=0 $Y2=0
cc_880 N_A_27_74#_c_1432_n N_VGND_c_1667_n 0.00948645f $X=0.28 $Y=0.58 $X2=0
+ $Y2=0
cc_881 N_VPWR_c_1506_n Q 0.0395687f $X=10.32 $Y=1.985 $X2=0 $Y2=0
cc_882 N_VPWR_c_1516_n Q 0.011066f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_883 N_VPWR_c_1499_n Q 0.00915947f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_884 N_Q_c_1638_n N_VGND_c_1659_n 0.027368f $X=10.665 $Y=0.515 $X2=0 $Y2=0
cc_885 N_Q_c_1638_n N_VGND_c_1666_n 0.0192663f $X=10.665 $Y=0.515 $X2=0 $Y2=0
cc_886 N_Q_c_1638_n N_VGND_c_1667_n 0.0158831f $X=10.665 $Y=0.515 $X2=0 $Y2=0

* File: sky130_fd_sc_ms__sdfsbp_1.pex.spice
* Created: Wed Sep  2 12:30:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__SDFSBP_1%SCE 3 7 9 11 17 19 20 23 24 28 33 39
c77 39 0 1.89796e-19 $X=0.67 $Y=1.535
c78 24 0 1.10806e-19 $X=1.96 $Y=1.425
c79 23 0 1.50331e-19 $X=1.96 $Y=1.425
r80 31 33 29.4556 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.685
+ $X2=0.67 $Y2=1.685
r81 30 31 1.78519 $w=2.7e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.685
+ $X2=0.505 $Y2=1.685
r82 28 39 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.67 $Y=1.665
+ $X2=0.67 $Y2=1.535
r83 28 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.67
+ $Y=1.685 $X2=0.67 $Y2=1.685
r84 24 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.96 $Y=1.425
+ $X2=1.96 $Y2=1.26
r85 23 26 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=1.92 $Y=1.425
+ $X2=1.92 $Y2=1.535
r86 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.96
+ $Y=1.425 $X2=1.96 $Y2=1.425
r87 21 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.835 $Y=1.535
+ $X2=0.67 $Y2=1.535
r88 20 26 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.795 $Y=1.535
+ $X2=1.92 $Y2=1.535
r89 20 21 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.795 $Y=1.535
+ $X2=0.835 $Y2=1.535
r90 17 37 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.885 $Y=0.58
+ $X2=1.885 $Y2=1.26
r91 13 33 53.5556 $w=2.7e-07 $l=3.73497e-07 $layer=POLY_cond $X=0.97 $Y=1.85
+ $X2=0.67 $Y2=1.685
r92 13 19 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.97 $Y=1.85
+ $X2=0.97 $Y2=2.09
r93 9 19 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=0.955 $Y=2.18 $X2=0.955
+ $Y2=2.09
r94 9 11 178.806 $w=1.8e-07 $l=4.6e-07 $layer=POLY_cond $X=0.955 $Y=2.18
+ $X2=0.955 $Y2=2.64
r95 5 30 16.5046 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.52
+ $X2=0.495 $Y2=1.685
r96 5 7 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=0.495 $Y=1.52 $X2=0.495
+ $Y2=0.58
r97 1 31 12.2893 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.85
+ $X2=0.505 $Y2=1.685
r98 1 3 307.081 $w=1.8e-07 $l=7.9e-07 $layer=POLY_cond $X=0.505 $Y=1.85
+ $X2=0.505 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSBP_1%A_27_74# 1 2 9 13 17 20 23 25 29 30 34 35
+ 37 38
c85 34 0 1.30624e-19 $X=1.96 $Y=1.995
c86 30 0 2.93935e-19 $X=0.975 $Y=1.115
c87 25 0 1.60946e-19 $X=1.795 $Y=2.375
c88 9 0 1.50564e-19 $X=1.065 $Y=0.58
r89 35 44 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.96 $Y=1.995
+ $X2=1.96 $Y2=2.16
r90 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.96
+ $Y=1.995 $X2=1.96 $Y2=1.995
r91 32 34 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.92 $Y=2.29
+ $X2=1.92 $Y2=1.995
r92 30 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.115
+ $X2=0.975 $Y2=0.95
r93 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.115 $X2=0.975 $Y2=1.115
r94 27 37 0.695019 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=1.115
+ $X2=0.28 $Y2=1.115
r95 27 29 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=0.445 $Y=1.115
+ $X2=0.975 $Y2=1.115
r96 26 38 2.53056 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=2.375
+ $X2=0.24 $Y2=2.375
r97 25 32 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.795 $Y=2.375
+ $X2=1.92 $Y2=2.29
r98 25 26 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=1.795 $Y=2.375
+ $X2=0.365 $Y2=2.375
r99 21 38 3.91525 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=2.46
+ $X2=0.24 $Y2=2.375
r100 21 23 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.24 $Y=2.46
+ $X2=0.24 $Y2=2.465
r101 20 38 3.91525 $w=2.35e-07 $l=9.21954e-08 $layer=LI1_cond $X=0.225 $Y=2.29
+ $X2=0.24 $Y2=2.375
r102 19 37 5.99569 $w=2.75e-07 $l=1.90526e-07 $layer=LI1_cond $X=0.225 $Y=1.28
+ $X2=0.28 $Y2=1.115
r103 19 20 52.9076 $w=2.18e-07 $l=1.01e-06 $layer=LI1_cond $X=0.225 $Y=1.28
+ $X2=0.225 $Y2=2.29
r104 15 37 5.99569 $w=2.75e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=0.95
+ $X2=0.28 $Y2=1.115
r105 15 17 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=0.95
+ $X2=0.28 $Y2=0.58
r106 13 44 186.581 $w=1.8e-07 $l=4.8e-07 $layer=POLY_cond $X=2.005 $Y=2.64
+ $X2=2.005 $Y2=2.16
r107 9 40 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.065 $Y=0.58
+ $X2=1.065 $Y2=0.95
r108 2 23 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.32 $X2=0.28 $Y2=2.465
r109 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSBP_1%D 3 7 9 12 13
c39 12 0 2.35667e-19 $X=1.42 $Y=1.955
r40 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=1.955
+ $X2=1.42 $Y2=2.12
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=1.955
+ $X2=1.42 $Y2=1.79
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.42
+ $Y=1.955 $X2=1.42 $Y2=1.955
r43 9 13 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.2 $Y=1.955 $X2=1.42
+ $Y2=1.955
r44 7 14 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=1.455 $Y=0.58
+ $X2=1.455 $Y2=1.79
r45 3 15 202.129 $w=1.8e-07 $l=5.2e-07 $layer=POLY_cond $X=1.375 $Y=2.64
+ $X2=1.375 $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSBP_1%SCD 1 3 4 6 7 8 9 10 11
c44 9 0 7.19792e-20 $X=2.64 $Y=1.295
c45 8 0 1.50331e-19 $X=2.597 $Y=1.918
c46 4 0 2.91569e-19 $X=2.425 $Y=2.24
r47 11 19 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.665
+ $Y=1.985 $X2=2.665 $Y2=1.985
r48 10 11 16.9004 $w=2.08e-07 $l=3.2e-07 $layer=LI1_cond $X=2.66 $Y=1.665
+ $X2=2.66 $Y2=1.985
r49 9 10 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.66 $Y=1.295
+ $X2=2.66 $Y2=1.665
r50 9 16 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.665
+ $Y=1.305 $X2=2.665 $Y2=1.305
r51 8 19 8.51415 $w=4.65e-07 $l=7.41215e-08 $layer=POLY_cond $X=2.597 $Y=1.918
+ $X2=2.582 $Y2=1.985
r52 7 16 10.4119 $w=4.65e-07 $l=1.10535e-07 $layer=POLY_cond $X=2.597 $Y=1.372
+ $X2=2.515 $Y2=1.305
r53 7 8 65.3032 $w=4.65e-07 $l=5.46e-07 $layer=POLY_cond $X=2.597 $Y=1.372
+ $X2=2.597 $Y2=1.918
r54 4 19 45.6887 $w=3.85e-07 $l=3.2413e-07 $layer=POLY_cond $X=2.425 $Y=2.24
+ $X2=2.582 $Y2=1.985
r55 4 6 107.111 $w=1.8e-07 $l=4e-07 $layer=POLY_cond $X=2.425 $Y=2.24 $X2=2.425
+ $Y2=2.64
r56 1 16 77.4558 $w=3.42e-07 $l=5.46992e-07 $layer=POLY_cond $X=2.275 $Y=0.865
+ $X2=2.515 $Y2=1.305
r57 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.275 $Y=0.865
+ $X2=2.275 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSBP_1%CLK 1 3 4 6 7
c33 4 0 7.19792e-20 $X=3.515 $Y=1.76
c34 1 0 9.27061e-20 $X=3.33 $Y=1.22
r35 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.38
+ $Y=1.385 $X2=3.38 $Y2=1.385
r36 7 11 6.85236 $w=3.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.6 $Y=1.365 $X2=3.38
+ $Y2=1.365
r37 4 10 71.3149 $w=2.76e-07 $l=4.24264e-07 $layer=POLY_cond $X=3.515 $Y=1.76
+ $X2=3.41 $Y2=1.385
r38 4 6 171.378 $w=1.8e-07 $l=6.4e-07 $layer=POLY_cond $X=3.515 $Y=1.76
+ $X2=3.515 $Y2=2.4
r39 1 10 38.7914 $w=2.76e-07 $l=2.0106e-07 $layer=POLY_cond $X=3.33 $Y=1.22
+ $X2=3.41 $Y2=1.385
r40 1 3 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.33 $Y=1.22 $X2=3.33
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSBP_1%A_781_74# 1 2 9 15 19 23 26 30 32 33 34 35
+ 36 38 39 43 44 45 48 49 50 52 53 54 56 57 60 63 64 72 77
c207 77 0 1.72394e-19 $X=8.825 $Y=1.795
c208 56 0 3.2492e-19 $X=8.745 $Y=1.95
c209 52 0 1.38381e-19 $X=7.36 $Y=2.905
c210 33 0 9.27061e-20 $X=4.21 $Y=0.34
r211 71 72 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.5 $Y=1.855
+ $X2=5.425 $Y2=1.855
r212 69 70 59.925 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=4.925 $Y=1.765
+ $X2=4.925 $Y2=2.04
r213 64 77 60.7993 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=8.825 $Y=1.515
+ $X2=8.825 $Y2=1.795
r214 64 76 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.825 $Y=1.515
+ $X2=8.825 $Y2=1.35
r215 63 66 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.825 $Y=1.515
+ $X2=8.825 $Y2=1.68
r216 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.825
+ $Y=1.515 $X2=8.825 $Y2=1.515
r217 60 71 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=5.645 $Y=1.855
+ $X2=5.5 $Y2=1.855
r218 59 61 16.8553 $w=2.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.675 $Y=1.855
+ $X2=5.675 $Y2=2.17
r219 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.645
+ $Y=1.855 $X2=5.645 $Y2=1.855
r220 56 66 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.745 $Y=1.95
+ $X2=8.745 $Y2=1.68
r221 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.66 $Y=2.035
+ $X2=8.745 $Y2=1.95
r222 53 54 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=8.66 $Y=2.035
+ $X2=7.445 $Y2=2.035
r223 51 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.36 $Y=2.12
+ $X2=7.445 $Y2=2.035
r224 51 52 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=7.36 $Y=2.12
+ $X2=7.36 $Y2=2.905
r225 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.275 $Y=2.99
+ $X2=7.36 $Y2=2.905
r226 49 50 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.275 $Y=2.99
+ $X2=6.765 $Y2=2.99
r227 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.68 $Y=2.905
+ $X2=6.765 $Y2=2.99
r228 47 48 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.68 $Y=2.255
+ $X2=6.68 $Y2=2.905
r229 46 61 2.45823 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.81 $Y=2.17
+ $X2=5.675 $Y2=2.17
r230 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.595 $Y=2.17
+ $X2=6.68 $Y2=2.255
r231 45 46 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=6.595 $Y=2.17
+ $X2=5.81 $Y2=2.17
r232 43 61 5.36411 $w=2.28e-07 $l=1.07121e-07 $layer=LI1_cond $X=5.725 $Y=2.255
+ $X2=5.675 $Y2=2.17
r233 43 44 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.725 $Y=2.255
+ $X2=5.725 $Y2=2.905
r234 41 57 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=4.945 $Y=0.425
+ $X2=4.945 $Y2=1.37
r235 39 69 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=4.925 $Y=1.535
+ $X2=4.925 $Y2=1.765
r236 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.925
+ $Y=1.535 $X2=4.925 $Y2=1.535
r237 36 57 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.895 $Y=1.505
+ $X2=4.895 $Y2=1.37
r238 36 38 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=4.895 $Y=1.505
+ $X2=4.895 $Y2=1.535
r239 34 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.64 $Y=2.99
+ $X2=5.725 $Y2=2.905
r240 34 35 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=5.64 $Y=2.99
+ $X2=4.355 $Y2=2.99
r241 32 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.86 $Y=0.34
+ $X2=4.945 $Y2=0.425
r242 32 33 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.86 $Y=0.34
+ $X2=4.21 $Y2=0.34
r243 28 35 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.23 $Y=2.905
+ $X2=4.355 $Y2=2.99
r244 28 30 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=4.23 $Y=2.905
+ $X2=4.23 $Y2=2.765
r245 24 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.045 $Y=0.425
+ $X2=4.21 $Y2=0.34
r246 24 26 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.045 $Y=0.425
+ $X2=4.045 $Y2=0.505
r247 23 77 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=8.9 $Y=2.08
+ $X2=8.9 $Y2=1.795
r248 19 76 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.735 $Y=0.69
+ $X2=8.735 $Y2=1.35
r249 13 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.5 $Y=1.69
+ $X2=5.5 $Y2=1.855
r250 13 15 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=5.5 $Y=1.69 $X2=5.5
+ $Y2=0.58
r251 12 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.09 $Y=1.765
+ $X2=4.925 $Y2=1.765
r252 12 72 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.09 $Y=1.765
+ $X2=5.425 $Y2=1.765
r253 9 70 188.524 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=4.985 $Y=2.525
+ $X2=4.985 $Y2=2.04
r254 2 30 600 $w=1.7e-07 $l=9.90202e-07 $layer=licon1_PDIFF $count=1 $X=4.055
+ $Y=1.84 $X2=4.19 $Y2=2.765
r255 1 26 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=3.905
+ $Y=0.37 $X2=4.045 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSBP_1%A_1163_48# 1 2 7 9 10 12 15 16 18 25 32
r70 34 36 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=5.89 $Y=1.065
+ $X2=6.125 $Y2=1.065
r71 32 36 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=6.32 $Y=1.065
+ $X2=6.125 $Y2=1.065
r72 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.32
+ $Y=1.065 $X2=6.32 $Y2=1.065
r73 23 25 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.02 $Y=1.915 $X2=7.02
+ $Y2=2.515
r74 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.215
+ $Y=1.8 $X2=6.215 $Y2=1.8
r75 18 23 6.9898 $w=2.25e-07 $l=1.49579e-07 $layer=LI1_cond $X=6.935 $Y=1.802
+ $X2=7.02 $Y2=1.915
r76 18 20 36.8782 $w=2.23e-07 $l=7.2e-07 $layer=LI1_cond $X=6.935 $Y=1.802
+ $X2=6.215 $Y2=1.802
r77 16 31 3.99273 $w=3.3e-07 $l=1.33492e-07 $layer=LI1_cond $X=6.263 $Y=0.957
+ $X2=6.32 $Y2=1.065
r78 16 28 15.4164 $w=3.3e-07 $l=6.79219e-07 $layer=LI1_cond $X=6.263 $Y=0.957
+ $X2=6.765 $Y2=0.54
r79 15 21 38.7084 $w=3.43e-07 $l=1.98997e-07 $layer=POLY_cond $X=6.125 $Y=1.635
+ $X2=6.2 $Y2=1.8
r80 14 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.125 $Y=1.23
+ $X2=6.125 $Y2=1.065
r81 14 15 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=6.125 $Y=1.23
+ $X2=6.125 $Y2=1.635
r82 10 21 34.0194 $w=3.43e-07 $l=2.05122e-07 $layer=POLY_cond $X=6.11 $Y=1.965
+ $X2=6.2 $Y2=1.8
r83 10 12 217.677 $w=1.8e-07 $l=5.6e-07 $layer=POLY_cond $X=6.11 $Y=1.965
+ $X2=6.11 $Y2=2.525
r84 7 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.89 $Y=0.9 $X2=5.89
+ $Y2=1.065
r85 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.89 $Y=0.9 $X2=5.89
+ $Y2=0.58
r86 2 25 600 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_PDIFF $count=1 $X=6.885
+ $Y=2.315 $X2=7.02 $Y2=2.515
r87 1 28 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=6.62
+ $Y=0.37 $X2=6.765 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSBP_1%A_995_74# 1 2 7 9 13 17 19 21 24 27 28 30
+ 34 38 40 43 50
c128 9 0 1.19047e-19 $X=6.795 $Y=2.525
r129 43 45 3.42456 $w=2.85e-07 $l=8e-08 $layer=LI1_cond $X=6.917 $Y=1.355
+ $X2=6.917 $Y2=1.435
r130 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.89
+ $Y=1.355 $X2=6.89 $Y2=1.355
r131 35 50 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=8 $Y=1.285
+ $X2=8.345 $Y2=1.285
r132 35 47 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8 $Y=1.285
+ $X2=7.925 $Y2=1.285
r133 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8
+ $Y=1.285 $X2=8 $Y2=1.285
r134 32 34 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=8 $Y=1.075 $X2=8
+ $Y2=1.285
r135 31 43 15.6246 $w=2.85e-07 $l=4.51298e-07 $layer=LI1_cond $X=7.11 $Y=0.99
+ $X2=6.917 $Y2=1.355
r136 30 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.835 $Y=0.99
+ $X2=8 $Y2=1.075
r137 30 31 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=7.835 $Y=0.99
+ $X2=7.11 $Y2=0.99
r138 29 40 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.45 $Y=1.435
+ $X2=5.325 $Y2=1.435
r139 28 45 3.76007 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=6.725 $Y=1.435
+ $X2=6.917 $Y2=1.435
r140 28 29 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=6.725 $Y=1.435
+ $X2=5.45 $Y2=1.435
r141 27 38 8.98601 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=5.285 $Y=2.37
+ $X2=5.285 $Y2=2.55
r142 26 40 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=5.285 $Y=1.52
+ $X2=5.325 $Y2=1.435
r143 26 27 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=5.285 $Y=1.52
+ $X2=5.285 $Y2=2.37
r144 22 40 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.325 $Y=1.35
+ $X2=5.325 $Y2=1.435
r145 22 24 35.4952 $w=2.48e-07 $l=7.7e-07 $layer=LI1_cond $X=5.325 $Y=1.35
+ $X2=5.325 $Y2=0.58
r146 19 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.345 $Y=1.12
+ $X2=8.345 $Y2=1.285
r147 19 21 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.345 $Y=1.12
+ $X2=8.345 $Y2=0.69
r148 15 47 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.925 $Y=1.45
+ $X2=7.925 $Y2=1.285
r149 15 17 305.137 $w=1.8e-07 $l=7.85e-07 $layer=POLY_cond $X=7.925 $Y=1.45
+ $X2=7.925 $Y2=2.235
r150 11 44 38.5662 $w=2.97e-07 $l=2.09105e-07 $layer=POLY_cond $X=6.98 $Y=1.19
+ $X2=6.88 $Y2=1.355
r151 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.98 $Y=1.19
+ $X2=6.98 $Y2=0.58
r152 7 44 48.8089 $w=2.97e-07 $l=2.94449e-07 $layer=POLY_cond $X=6.795 $Y=1.61
+ $X2=6.88 $Y2=1.355
r153 7 9 355.669 $w=1.8e-07 $l=9.15e-07 $layer=POLY_cond $X=6.795 $Y=1.61
+ $X2=6.795 $Y2=2.525
r154 2 38 600 $w=1.7e-07 $l=3.23381e-07 $layer=licon1_PDIFF $count=1 $X=5.075
+ $Y=2.315 $X2=5.285 $Y2=2.55
r155 1 24 182 $w=1.7e-07 $l=4.01497e-07 $layer=licon1_NDIFF $count=1 $X=4.975
+ $Y=0.37 $X2=5.285 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSBP_1%SET_B 3 7 9 11 12 13 20 22 23 25 26 29 31
+ 32 37 40 41 45
c147 41 0 1.19047e-19 $X=7.46 $Y=1.41
c148 26 0 1.8354e-19 $X=10.75 $Y=1.42
c149 13 0 7.13225e-20 $X=10.31 $Y=0.94
c150 12 0 1.94471e-19 $X=10.55 $Y=0.94
c151 7 0 3.21009e-19 $X=7.385 $Y=2.525
r152 40 43 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.46 $Y=1.41
+ $X2=7.46 $Y2=1.575
r153 40 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.46 $Y=1.41
+ $X2=7.46 $Y2=1.245
r154 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.46
+ $Y=1.41 $X2=7.46 $Y2=1.41
r155 37 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=1.665
+ $X2=9.84 $Y2=1.665
r156 35 41 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=7.46 $Y=1.665
+ $X2=7.46 $Y2=1.41
r157 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=1.665
+ $X2=7.44 $Y2=1.665
r158 32 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.585 $Y=1.665
+ $X2=7.44 $Y2=1.665
r159 31 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.695 $Y=1.665
+ $X2=9.84 $Y2=1.665
r160 31 32 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=9.695 $Y=1.665
+ $X2=7.585 $Y2=1.665
r161 29 51 37.3291 $w=2.28e-07 $l=7.45e-07 $layer=LI1_cond $X=10.585 $Y=1.665
+ $X2=9.84 $Y2=1.665
r162 28 29 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=10.75 $Y=1.665
+ $X2=10.585 $Y2=1.665
r163 26 45 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=10.75 $Y=1.42
+ $X2=10.75 $Y2=1.255
r164 25 28 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=10.75 $Y=1.42
+ $X2=10.75 $Y2=1.665
r165 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.75
+ $Y=1.42 $X2=10.75 $Y2=1.42
r166 22 23 37.8919 $w=4e-07 $l=1.5e-07 $layer=POLY_cond $X=10.765 $Y=1.775
+ $X2=10.765 $Y2=1.925
r167 20 23 320.685 $w=1.8e-07 $l=8.25e-07 $layer=POLY_cond $X=10.89 $Y=2.75
+ $X2=10.89 $Y2=1.925
r168 16 26 4.86635 $w=4e-07 $l=3.5e-08 $layer=POLY_cond $X=10.75 $Y=1.455
+ $X2=10.75 $Y2=1.42
r169 16 22 44.4923 $w=4e-07 $l=3.2e-07 $layer=POLY_cond $X=10.75 $Y=1.455
+ $X2=10.75 $Y2=1.775
r170 14 45 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=10.625 $Y=1.015
+ $X2=10.625 $Y2=1.255
r171 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.55 $Y=0.94
+ $X2=10.625 $Y2=1.015
r172 12 13 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=10.55 $Y=0.94
+ $X2=10.31 $Y2=0.94
r173 9 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.235 $Y=0.865
+ $X2=10.31 $Y2=0.94
r174 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.235 $Y=0.865
+ $X2=10.235 $Y2=0.58
r175 7 43 369.274 $w=1.8e-07 $l=9.5e-07 $layer=POLY_cond $X=7.385 $Y=2.525
+ $X2=7.385 $Y2=1.575
r176 3 42 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=7.37 $Y=0.58
+ $X2=7.37 $Y2=1.245
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSBP_1%A_594_74# 1 2 7 9 12 14 17 18 20 21 24 28
+ 30 34 36 39 40 43 50 53 55 56 60 61 63 65 66
c175 56 0 2.88662e-20 $X=3.885 $Y=1.905
c176 39 0 1.73559e-19 $X=9.44 $Y=2.37
c177 36 0 1.51361e-19 $X=9.44 $Y=1.795
c178 17 0 1.81976e-19 $X=4.475 $Y=3.075
r179 65 66 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.29 $Y=1.985
+ $X2=3.455 $Y2=1.985
r180 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.05
+ $Y=1.385 $X2=4.05 $Y2=1.385
r181 58 60 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=4.05 $Y=1.82
+ $X2=4.05 $Y2=1.385
r182 56 58 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.885 $Y=1.905
+ $X2=4.05 $Y2=1.82
r183 56 66 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.885 $Y=1.905
+ $X2=3.455 $Y2=1.905
r184 55 65 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=3.105 $Y=1.985
+ $X2=3.29 $Y2=1.985
r185 53 55 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.02 $Y=1.82
+ $X2=3.105 $Y2=1.985
r186 53 63 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=3.02 $Y=1.82
+ $X2=3.02 $Y2=1.01
r187 48 63 7.21712 $w=2.63e-07 $l=1.32e-07 $layer=LI1_cond $X=3.067 $Y=0.878
+ $X2=3.067 $Y2=1.01
r188 48 50 16.2212 $w=2.63e-07 $l=3.73e-07 $layer=LI1_cond $X=3.067 $Y=0.878
+ $X2=3.067 $Y2=0.505
r189 37 39 274.04 $w=1.8e-07 $l=7.05e-07 $layer=POLY_cond $X=9.44 $Y=3.075
+ $X2=9.44 $Y2=2.37
r190 36 44 69.2234 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.44 $Y=1.72
+ $X2=9.305 $Y2=1.72
r191 36 39 223.508 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.44 $Y=1.795
+ $X2=9.44 $Y2=2.37
r192 32 44 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.305 $Y=1.645
+ $X2=9.305 $Y2=1.72
r193 32 34 546.096 $w=1.5e-07 $l=1.065e-06 $layer=POLY_cond $X=9.305 $Y=1.645
+ $X2=9.305 $Y2=0.58
r194 31 43 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.68 $Y=3.15 $X2=5.59
+ $Y2=3.15
r195 30 37 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=9.35 $Y=3.15
+ $X2=9.44 $Y2=3.075
r196 30 31 1881.85 $w=1.5e-07 $l=3.67e-06 $layer=POLY_cond $X=9.35 $Y=3.15
+ $X2=5.68 $Y2=3.15
r197 26 43 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=5.59 $Y=3.075
+ $X2=5.59 $Y2=3.15
r198 26 28 184.637 $w=1.8e-07 $l=4.75e-07 $layer=POLY_cond $X=5.59 $Y=3.075
+ $X2=5.59 $Y2=2.6
r199 22 24 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.9 $Y=0.98 $X2=4.9
+ $Y2=0.58
r200 20 43 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=5.5 $Y=3.15 $X2=5.59
+ $Y2=3.15
r201 20 21 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.5 $Y=3.15
+ $X2=4.55 $Y2=3.15
r202 19 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.55 $Y=1.055
+ $X2=4.475 $Y2=1.055
r203 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.825 $Y=1.055
+ $X2=4.9 $Y2=0.98
r204 18 19 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=4.825 $Y=1.055
+ $X2=4.55 $Y2=1.055
r205 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.475 $Y=3.075
+ $X2=4.55 $Y2=3.15
r206 16 17 781.968 $w=1.5e-07 $l=1.525e-06 $layer=POLY_cond $X=4.475 $Y=1.55
+ $X2=4.475 $Y2=3.075
r207 15 61 3.90195 $w=3.3e-07 $l=3.73497e-07 $layer=POLY_cond $X=4.055 $Y=1.385
+ $X2=3.755 $Y2=1.22
r208 14 16 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.475 $Y=1.385
+ $X2=4.475 $Y2=1.55
r209 14 40 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.475 $Y=1.385
+ $X2=4.475 $Y2=1.055
r210 14 15 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=4.4 $Y=1.385
+ $X2=4.055 $Y2=1.385
r211 10 61 34.7346 $w=1.65e-07 $l=4.22137e-07 $layer=POLY_cond $X=3.965 $Y=1.55
+ $X2=3.755 $Y2=1.22
r212 10 12 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=3.965 $Y=1.55
+ $X2=3.965 $Y2=2.4
r213 7 61 34.7346 $w=1.65e-07 $l=7.5e-08 $layer=POLY_cond $X=3.83 $Y=1.22
+ $X2=3.755 $Y2=1.22
r214 7 9 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.83 $Y=1.22 $X2=3.83
+ $Y2=0.74
r215 2 65 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.15
+ $Y=1.84 $X2=3.29 $Y2=1.985
r216 1 50 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.97
+ $Y=0.37 $X2=3.115 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSBP_1%A_1924_48# 1 2 9 11 12 13 16 18 19 22 23 27
+ 30 31 32 35 37 38 40 41 45 47
c129 41 0 7.13225e-20 $X=9.785 $Y=0.985
c130 30 0 1.8354e-19 $X=11.31 $Y=1.3
c131 27 0 1.94471e-19 $X=11.23 $Y=0.58
r132 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.785
+ $Y=1.065 $X2=9.785 $Y2=1.065
r133 41 44 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=9.785 $Y=0.985
+ $X2=9.785 $Y2=1.065
r134 39 40 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=12.15 $Y=1.47
+ $X2=12.15 $Y2=2.18
r135 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.065 $Y=2.265
+ $X2=12.15 $Y2=2.18
r136 37 38 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.065 $Y=2.265
+ $X2=11.75 $Y2=2.265
r137 33 38 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=11.625 $Y=2.35
+ $X2=11.75 $Y2=2.265
r138 33 35 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=11.625 $Y=2.35
+ $X2=11.625 $Y2=2.75
r139 31 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.065 $Y=1.385
+ $X2=12.15 $Y2=1.47
r140 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=12.065 $Y=1.385
+ $X2=11.395 $Y2=1.385
r141 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.31 $Y=1.3
+ $X2=11.395 $Y2=1.385
r142 29 47 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=11.31 $Y=1.07
+ $X2=11.23 $Y2=0.985
r143 29 30 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=11.31 $Y=1.07
+ $X2=11.31 $Y2=1.3
r144 25 47 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.23 $Y=0.9
+ $X2=11.23 $Y2=0.985
r145 25 27 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=11.23 $Y=0.9
+ $X2=11.23 $Y2=0.58
r146 24 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.95 $Y=0.985
+ $X2=9.785 $Y2=0.985
r147 23 47 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.065 $Y=0.985
+ $X2=11.23 $Y2=0.985
r148 23 24 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=11.065 $Y=0.985
+ $X2=9.95 $Y2=0.985
r149 21 45 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=9.785 $Y=1.255
+ $X2=9.785 $Y2=1.065
r150 21 22 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=9.825 $Y=1.255
+ $X2=9.825 $Y2=1.405
r151 18 45 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=9.785 $Y=1.03
+ $X2=9.785 $Y2=1.065
r152 18 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.785 $Y=1.03
+ $X2=9.785 $Y2=0.865
r153 14 16 169.089 $w=1.8e-07 $l=4.35e-07 $layer=POLY_cond $X=10.44 $Y=2.315
+ $X2=10.44 $Y2=2.75
r154 12 14 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=10.35 $Y=2.24
+ $X2=10.44 $Y2=2.315
r155 12 13 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.35 $Y=2.24
+ $X2=10.03 $Y2=2.24
r156 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.955 $Y=2.165
+ $X2=10.03 $Y2=2.24
r157 11 22 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=9.955 $Y=2.165
+ $X2=9.955 $Y2=1.405
r158 9 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.695 $Y=0.58
+ $X2=9.695 $Y2=0.865
r159 2 35 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=11.525
+ $Y=2.54 $X2=11.665 $Y2=2.75
r160 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.09
+ $Y=0.37 $X2=11.23 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSBP_1%A_1762_74# 1 2 3 10 12 14 17 21 23 24 25 27
+ 28 32 34 36 39 41 42 45 46 50 52 56 58 62 66 67 70 75 76
c187 46 0 1.91489e-19 $X=13.14 $Y=1.79
r188 75 76 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=11.115 $Y=2.75
+ $X2=11.115 $Y2=2.52
r189 70 72 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=10.085 $Y=2.035
+ $X2=10.085 $Y2=2.18
r190 66 68 0.688026 $w=3.33e-07 $l=2e-08 $layer=LI1_cond $X=9.212 $Y=2.015
+ $X2=9.212 $Y2=2.035
r191 66 67 8.46614 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=9.212 $Y=2.015
+ $X2=9.212 $Y2=1.85
r192 64 67 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=9.295 $Y=1.05
+ $X2=9.295 $Y2=1.85
r193 62 64 17.5613 $w=5.93e-07 $l=5.35e-07 $layer=LI1_cond $X=9.082 $Y=0.515
+ $X2=9.082 $Y2=1.05
r194 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.73
+ $Y=1.805 $X2=11.73 $Y2=1.805
r195 56 80 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.195 $Y=1.805
+ $X2=11.195 $Y2=2.18
r196 56 58 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=11.28 $Y=1.805
+ $X2=11.73 $Y2=1.805
r197 54 80 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=11.195 $Y=2.265
+ $X2=11.195 $Y2=2.18
r198 54 76 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.195 $Y=2.265
+ $X2=11.195 $Y2=2.52
r199 53 72 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.17 $Y=2.18
+ $X2=10.085 $Y2=2.18
r200 52 80 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.11 $Y=2.18
+ $X2=11.195 $Y2=2.18
r201 52 53 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=11.11 $Y=2.18
+ $X2=10.17 $Y2=2.18
r202 51 68 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=9.38 $Y=2.035
+ $X2=9.212 $Y2=2.035
r203 50 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10 $Y=2.035
+ $X2=10.085 $Y2=2.035
r204 50 51 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=10 $Y=2.035
+ $X2=9.38 $Y2=2.035
r205 46 47 57.9764 $w=2.12e-07 $l=2.55e-07 $layer=POLY_cond $X=13.14 $Y=1.79
+ $X2=13.395 $Y2=1.79
r206 42 59 11.3783 $w=3.55e-07 $l=7e-08 $layer=POLY_cond $X=11.8 $Y=1.792
+ $X2=11.73 $Y2=1.792
r207 42 43 13.5596 $w=3.55e-07 $l=1.30457e-07 $layer=POLY_cond $X=11.8 $Y=1.792
+ $X2=11.89 $Y2=1.885
r208 41 59 57.7042 $w=3.55e-07 $l=3.55e-07 $layer=POLY_cond $X=11.375 $Y=1.792
+ $X2=11.73 $Y2=1.792
r209 37 39 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.015 $Y=0.94
+ $X2=11.3 $Y2=0.94
r210 34 47 6.70255 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=13.395 $Y=1.94
+ $X2=13.395 $Y2=1.79
r211 34 36 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=13.395 $Y=1.94
+ $X2=13.395 $Y2=2.435
r212 30 46 10.9192 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=13.14 $Y=1.615
+ $X2=13.14 $Y2=1.79
r213 30 32 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=13.14 $Y=1.615
+ $X2=13.14 $Y2=0.835
r214 29 45 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=12.485 $Y=1.69
+ $X2=12.395 $Y2=1.69
r215 28 46 21.2379 $w=2.12e-07 $l=1.32288e-07 $layer=POLY_cond $X=13.065 $Y=1.69
+ $X2=13.14 $Y2=1.79
r216 28 29 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=13.065 $Y=1.69
+ $X2=12.485 $Y2=1.69
r217 25 45 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=12.395 $Y=1.765
+ $X2=12.395 $Y2=1.69
r218 25 27 170.039 $w=1.8e-07 $l=6.35e-07 $layer=POLY_cond $X=12.395 $Y=1.765
+ $X2=12.395 $Y2=2.4
r219 23 45 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=12.305 $Y=1.69
+ $X2=12.395 $Y2=1.69
r220 23 24 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=12.305 $Y=1.69
+ $X2=12.15 $Y2=1.69
r221 19 24 24.0479 $w=2.99e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.075
+ $Y=1.615 $X2=12.15 $Y2=1.69
r222 19 43 29.8227 $w=2.99e-07 $l=3.505e-07 $layer=POLY_cond $X=12.075 $Y=1.615
+ $X2=11.89 $Y2=1.885
r223 19 21 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=12.075 $Y=1.615
+ $X2=12.075 $Y2=0.74
r224 15 43 14.6425 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=11.89 $Y=2.095
+ $X2=11.89 $Y2=1.885
r225 15 17 254.605 $w=1.8e-07 $l=6.55e-07 $layer=POLY_cond $X=11.89 $Y=2.095
+ $X2=11.89 $Y2=2.75
r226 14 41 33.1523 $w=3.55e-07 $l=2.11197e-07 $layer=POLY_cond $X=11.3 $Y=1.615
+ $X2=11.375 $Y2=1.792
r227 13 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.3 $Y=1.015
+ $X2=11.3 $Y2=0.94
r228 13 14 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=11.3 $Y=1.015 $X2=11.3
+ $Y2=1.615
r229 10 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.015 $Y=0.865
+ $X2=11.015 $Y2=0.94
r230 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.015 $Y=0.865
+ $X2=11.015 $Y2=0.58
r231 3 75 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=10.98
+ $Y=2.54 $X2=11.115 $Y2=2.75
r232 2 66 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=8.99
+ $Y=1.87 $X2=9.21 $Y2=2.015
r233 1 62 91 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_NDIFF $count=2 $X=8.81
+ $Y=0.37 $X2=9.09 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSBP_1%A_2556_112# 1 2 9 11 13 14 15 16 18 22
r47 26 27 19.3931 $w=3.46e-07 $l=5.5e-07 $layer=LI1_cond $X=13.047 $Y=0.835
+ $X2=13.047 $Y2=1.385
r48 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.62
+ $Y=1.385 $X2=13.62 $Y2=1.385
r49 20 27 1.00354 $w=3.3e-07 $l=2.08e-07 $layer=LI1_cond $X=13.255 $Y=1.385
+ $X2=13.047 $Y2=1.385
r50 20 22 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=13.255 $Y=1.385
+ $X2=13.62 $Y2=1.385
r51 16 27 6.77755 $w=3.46e-07 $l=2.02287e-07 $layer=LI1_cond $X=13.13 $Y=1.55
+ $X2=13.047 $Y2=1.385
r52 16 18 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=13.13 $Y=1.55
+ $X2=13.13 $Y2=2.16
r53 14 23 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=13.81 $Y=1.385
+ $X2=13.62 $Y2=1.385
r54 14 15 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=13.81 $Y=1.385
+ $X2=13.9 $Y2=1.385
r55 11 15 34.7346 $w=1.65e-07 $l=1.67481e-07 $layer=POLY_cond $X=13.905 $Y=1.22
+ $X2=13.9 $Y2=1.385
r56 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=13.905 $Y=1.22
+ $X2=13.905 $Y2=0.74
r57 7 15 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=13.9 $Y=1.55
+ $X2=13.9 $Y2=1.385
r58 7 9 330.403 $w=1.8e-07 $l=8.5e-07 $layer=POLY_cond $X=13.9 $Y=1.55 $X2=13.9
+ $Y2=2.4
r59 2 18 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=13.03
+ $Y=2.015 $X2=13.17 $Y2=2.16
r60 1 26 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=12.78
+ $Y=0.56 $X2=12.925 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSBP_1%VPWR 1 2 3 4 5 6 7 8 27 31 33 37 41 45 49
+ 53 57 60 61 63 64 66 67 68 70 75 102 109 116 117 120 123 126 129 132
c155 117 0 1.90308e-19 $X=14.16 $Y=3.33
c156 37 0 2.10842e-19 $X=3.74 $Y=2.78
r157 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r158 129 130 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r159 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r160 124 127 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r161 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r162 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r163 117 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.68 $Y2=3.33
r164 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r165 114 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.785 $Y=3.33
+ $X2=13.62 $Y2=3.33
r166 114 116 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.785 $Y=3.33
+ $X2=14.16 $Y2=3.33
r167 113 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r168 113 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.24 $Y2=3.33
r169 112 113 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r170 110 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.28 $Y=3.33
+ $X2=12.115 $Y2=3.33
r171 110 112 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=12.28 $Y=3.33
+ $X2=13.2 $Y2=3.33
r172 109 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.455 $Y=3.33
+ $X2=13.62 $Y2=3.33
r173 109 112 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=13.455 $Y=3.33
+ $X2=13.2 $Y2=3.33
r174 108 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r175 107 108 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r176 105 108 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.76 $Y2=3.33
r177 104 107 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=10.8 $Y=3.33
+ $X2=11.76 $Y2=3.33
r178 104 105 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r179 102 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.95 $Y=3.33
+ $X2=12.115 $Y2=3.33
r180 102 107 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=11.95 $Y=3.33
+ $X2=11.76 $Y2=3.33
r181 101 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r182 100 101 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r183 98 101 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=10.32 $Y2=3.33
r184 97 100 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=7.92 $Y=3.33
+ $X2=10.32 $Y2=3.33
r185 97 98 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r186 95 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r187 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r188 91 94 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r189 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r190 89 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r191 88 89 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r192 86 89 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=6 $Y2=3.33
r193 86 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r194 85 88 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=3.33 $X2=6
+ $Y2=3.33
r195 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r196 83 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=3.74 $Y2=3.33
r197 83 85 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=4.08 $Y2=3.33
r198 82 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r199 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r200 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r201 79 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r202 78 81 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r203 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r204 76 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r205 76 78 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r206 75 123 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.555 $Y=3.33
+ $X2=2.687 $Y2=3.33
r207 75 81 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.555 $Y=3.33
+ $X2=2.16 $Y2=3.33
r208 73 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r209 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r210 70 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r211 70 72 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r212 68 95 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=7.44 $Y2=3.33
r213 68 92 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=6.48 $Y2=3.33
r214 66 100 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=10.58 $Y=3.33
+ $X2=10.32 $Y2=3.33
r215 66 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.58 $Y=3.33
+ $X2=10.665 $Y2=3.33
r216 65 104 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=10.75 $Y=3.33
+ $X2=10.8 $Y2=3.33
r217 65 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.75 $Y=3.33
+ $X2=10.665 $Y2=3.33
r218 63 94 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=7.615 $Y=3.33
+ $X2=7.44 $Y2=3.33
r219 63 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.615 $Y=3.33
+ $X2=7.7 $Y2=3.33
r220 62 97 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=7.785 $Y=3.33
+ $X2=7.92 $Y2=3.33
r221 62 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.785 $Y=3.33
+ $X2=7.7 $Y2=3.33
r222 60 88 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.175 $Y=3.33
+ $X2=6 $Y2=3.33
r223 60 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.175 $Y=3.33
+ $X2=6.3 $Y2=3.33
r224 59 91 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=6.425 $Y=3.33
+ $X2=6.48 $Y2=3.33
r225 59 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.425 $Y=3.33
+ $X2=6.3 $Y2=3.33
r226 55 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.62 $Y=3.245
+ $X2=13.62 $Y2=3.33
r227 55 57 37.8909 $w=3.28e-07 $l=1.085e-06 $layer=LI1_cond $X=13.62 $Y=3.245
+ $X2=13.62 $Y2=2.16
r228 51 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.115 $Y=3.245
+ $X2=12.115 $Y2=3.33
r229 51 53 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=12.115 $Y=3.245
+ $X2=12.115 $Y2=2.75
r230 47 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.665 $Y=3.245
+ $X2=10.665 $Y2=3.33
r231 47 49 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=10.665 $Y=3.245
+ $X2=10.665 $Y2=2.75
r232 43 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.7 $Y=3.245 $X2=7.7
+ $Y2=3.33
r233 43 45 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=7.7 $Y=3.245
+ $X2=7.7 $Y2=2.525
r234 39 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.3 $Y=3.245
+ $X2=6.3 $Y2=3.33
r235 39 41 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=6.3 $Y=3.245
+ $X2=6.3 $Y2=2.59
r236 35 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.74 $Y=3.245
+ $X2=3.74 $Y2=3.33
r237 35 37 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.74 $Y=3.245
+ $X2=3.74 $Y2=2.78
r238 34 123 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=2.82 $Y=3.33
+ $X2=2.687 $Y2=3.33
r239 33 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.575 $Y=3.33
+ $X2=3.74 $Y2=3.33
r240 33 34 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=3.575 $Y=3.33
+ $X2=2.82 $Y2=3.33
r241 29 123 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.687 $Y=3.245
+ $X2=2.687 $Y2=3.33
r242 29 31 18.2651 $w=2.63e-07 $l=4.2e-07 $layer=LI1_cond $X=2.687 $Y=3.245
+ $X2=2.687 $Y2=2.825
r243 25 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r244 25 27 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.805
r245 8 57 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=13.485
+ $Y=2.015 $X2=13.62 $Y2=2.16
r246 7 53 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=11.98
+ $Y=2.54 $X2=12.115 $Y2=2.75
r247 6 49 600 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_PDIFF $count=1 $X=10.53
+ $Y=2.54 $X2=10.665 $Y2=2.75
r248 5 45 600 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_PDIFF $count=1 $X=7.475
+ $Y=2.315 $X2=7.7 $Y2=2.525
r249 4 41 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=6.2
+ $Y=2.315 $X2=6.34 $Y2=2.59
r250 3 37 600 $w=1.7e-07 $l=1.00524e-06 $layer=licon1_PDIFF $count=1 $X=3.605
+ $Y=1.84 $X2=3.74 $Y2=2.78
r251 2 31 600 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_PDIFF $count=1 $X=2.515
+ $Y=2.32 $X2=2.655 $Y2=2.825
r252 1 27 600 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=2.32 $X2=0.73 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSBP_1%A_293_464# 1 2 3 4 13 19 21 22 23 26 28 29
+ 31 34 37 39 40 41 48 50
c124 26 0 1.9349e-19 $X=2.3 $Y=2.32
c125 22 0 4.07687e-19 $X=1.835 $Y=1.005
r126 45 48 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=4.505 $Y=0.76
+ $X2=4.605 $Y2=0.76
r127 41 43 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.71 $Y=2.295
+ $X2=3.71 $Y2=2.405
r128 35 50 3.67481 $w=2.52e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.757 $Y=2.38
+ $X2=4.672 $Y2=2.295
r129 35 37 4.64417 $w=3.33e-07 $l=1.35e-07 $layer=LI1_cond $X=4.757 $Y=2.38
+ $X2=4.757 $Y2=2.515
r130 34 50 3.67481 $w=2.52e-07 $l=2.05144e-07 $layer=LI1_cond $X=4.505 $Y=2.21
+ $X2=4.672 $Y2=2.295
r131 33 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.505 $Y=0.925
+ $X2=4.505 $Y2=0.76
r132 33 34 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=4.505 $Y=0.925
+ $X2=4.505 $Y2=2.21
r133 32 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.795 $Y=2.295
+ $X2=3.71 $Y2=2.295
r134 31 50 2.79892 $w=1.7e-07 $l=2.52e-07 $layer=LI1_cond $X=4.42 $Y=2.295
+ $X2=4.672 $Y2=2.295
r135 31 32 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=4.42 $Y=2.295
+ $X2=3.795 $Y2=2.295
r136 30 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=2.405
+ $X2=2.3 $Y2=2.405
r137 29 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=2.405
+ $X2=3.71 $Y2=2.405
r138 29 30 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=3.625 $Y=2.405
+ $X2=2.385 $Y2=2.405
r139 27 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=2.49 $X2=2.3
+ $Y2=2.405
r140 27 28 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.3 $Y=2.49 $X2=2.3
+ $Y2=2.63
r141 26 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=2.32 $X2=2.3
+ $Y2=2.405
r142 25 26 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=2.3 $Y=1.09 $X2=2.3
+ $Y2=2.32
r143 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.215 $Y=2.715
+ $X2=2.3 $Y2=2.63
r144 23 39 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.215 $Y=2.715
+ $X2=1.945 $Y2=2.715
r145 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.215 $Y=1.005
+ $X2=2.3 $Y2=1.09
r146 21 22 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.215 $Y=1.005
+ $X2=1.835 $Y2=1.005
r147 17 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.67 $Y=0.92
+ $X2=1.835 $Y2=1.005
r148 17 19 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.67 $Y=0.92
+ $X2=1.67 $Y2=0.58
r149 13 39 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.78 $Y=2.795
+ $X2=1.945 $Y2=2.795
r150 13 15 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.78 $Y=2.795
+ $X2=1.69 $Y2=2.795
r151 4 37 600 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_PDIFF $count=1 $X=4.625
+ $Y=2.315 $X2=4.76 $Y2=2.515
r152 3 15 600 $w=1.7e-07 $l=5.76628e-07 $layer=licon1_PDIFF $count=1 $X=1.465
+ $Y=2.32 $X2=1.69 $Y2=2.795
r153 2 48 182 $w=1.7e-07 $l=4.56782e-07 $layer=licon1_NDIFF $count=1 $X=4.46
+ $Y=0.37 $X2=4.605 $Y2=0.76
r154 1 19 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.53
+ $Y=0.37 $X2=1.67 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSBP_1%A_1603_347# 1 2 7 9 16
c34 9 0 2.69082e-19 $X=8.15 $Y=2.435
r35 9 12 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.15 $Y=2.435
+ $X2=8.15 $Y2=2.52
r36 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.315 $Y=2.435
+ $X2=8.15 $Y2=2.435
r37 7 16 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.58 $Y=2.435
+ $X2=9.705 $Y2=2.435
r38 7 8 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=9.58 $Y=2.435
+ $X2=8.315 $Y2=2.435
r39 2 16 600 $w=1.7e-07 $l=7.04273e-07 $layer=licon1_PDIFF $count=1 $X=9.53
+ $Y=1.87 $X2=9.665 $Y2=2.51
r40 1 12 600 $w=1.7e-07 $l=8.49823e-07 $layer=licon1_PDIFF $count=1 $X=8.015
+ $Y=1.735 $X2=8.15 $Y2=2.52
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSBP_1%A_1712_374# 1 2 7 11 14
c31 14 0 1.72394e-19 $X=8.695 $Y=2.855
r32 14 16 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=8.695 $Y=2.855
+ $X2=8.695 $Y2=2.99
r33 9 11 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=10.215 $Y=2.905
+ $X2=10.215 $Y2=2.75
r34 8 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.86 $Y=2.99
+ $X2=8.695 $Y2=2.99
r35 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.05 $Y=2.99
+ $X2=10.215 $Y2=2.905
r36 7 8 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=10.05 $Y=2.99
+ $X2=8.86 $Y2=2.99
r37 2 11 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=10.075
+ $Y=2.54 $X2=10.215 $Y2=2.75
r38 1 14 600 $w=1.7e-07 $l=1.05033e-06 $layer=licon1_PDIFF $count=1 $X=8.56
+ $Y=1.87 $X2=8.695 $Y2=2.855
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSBP_1%Q_N 1 2 9 11 15 16 17 28
c34 15 0 1.91489e-19 $X=12.577 $Y=1.82
r35 21 28 1.01485 $w=4.93e-07 $l=4.2e-08 $layer=LI1_cond $X=12.372 $Y=0.883
+ $X2=12.372 $Y2=0.925
r36 17 30 9.94566 $w=4.93e-07 $l=1.84e-07 $layer=LI1_cond $X=12.372 $Y=0.946
+ $X2=12.372 $Y2=1.13
r37 17 28 0.507427 $w=4.93e-07 $l=2.1e-08 $layer=LI1_cond $X=12.372 $Y=0.946
+ $X2=12.372 $Y2=0.925
r38 17 21 0.53159 $w=4.93e-07 $l=2.2e-08 $layer=LI1_cond $X=12.372 $Y=0.861
+ $X2=12.372 $Y2=0.883
r39 16 17 8.36047 $w=4.93e-07 $l=3.46e-07 $layer=LI1_cond $X=12.372 $Y=0.515
+ $X2=12.372 $Y2=0.861
r40 15 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=12.535 $Y=1.82
+ $X2=12.535 $Y2=1.13
r41 11 13 37.5109 $w=2.53e-07 $l=8.3e-07 $layer=LI1_cond $X=12.577 $Y=1.985
+ $X2=12.577 $Y2=2.815
r42 9 15 7.02311 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=12.577 $Y=1.947
+ $X2=12.577 $Y2=1.82
r43 9 11 1.71737 $w=2.53e-07 $l=3.8e-08 $layer=LI1_cond $X=12.577 $Y=1.947
+ $X2=12.577 $Y2=1.985
r44 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=12.485
+ $Y=1.84 $X2=12.62 $Y2=2.815
r45 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=12.485
+ $Y=1.84 $X2=12.62 $Y2=1.985
r46 1 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.15
+ $Y=0.37 $X2=12.29 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSBP_1%Q 1 2 7 8 9 10 11 12 13
r14 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=14.122 $Y=2.405
+ $X2=14.122 $Y2=2.775
r15 11 12 14.4485 $w=3.33e-07 $l=4.2e-07 $layer=LI1_cond $X=14.122 $Y=1.985
+ $X2=14.122 $Y2=2.405
r16 10 11 11.0084 $w=3.33e-07 $l=3.2e-07 $layer=LI1_cond $X=14.122 $Y=1.665
+ $X2=14.122 $Y2=1.985
r17 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=14.122 $Y=1.295
+ $X2=14.122 $Y2=1.665
r18 8 9 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=14.122 $Y=0.925
+ $X2=14.122 $Y2=1.295
r19 7 8 14.1045 $w=3.33e-07 $l=4.1e-07 $layer=LI1_cond $X=14.122 $Y=0.515
+ $X2=14.122 $Y2=0.925
r20 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=13.99
+ $Y=1.84 $X2=14.125 $Y2=2.815
r21 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=13.99
+ $Y=1.84 $X2=14.125 $Y2=1.985
r22 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.98
+ $Y=0.37 $X2=14.12 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__SDFSBP_1%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 50
+ 51 53 54 55 57 69 87 92 97 107 108 111 114 119 122 125 133 136
r146 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r147 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r148 126 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r149 125 130 10.098 $w=6.08e-07 $l=5.15e-07 $layer=LI1_cond $X=10.59 $Y=0
+ $X2=10.59 $Y2=0.515
r150 125 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r151 125 126 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r152 121 122 11.5563 $w=8.18e-07 $l=1.65e-07 $layer=LI1_cond $X=8.13 $Y=0.325
+ $X2=8.295 $Y2=0.325
r153 117 121 3.06313 $w=8.18e-07 $l=2.1e-07 $layer=LI1_cond $X=7.92 $Y=0.325
+ $X2=8.13 $Y2=0.325
r154 117 119 15.2758 $w=8.18e-07 $l=4.2e-07 $layer=LI1_cond $X=7.92 $Y=0.325
+ $X2=7.5 $Y2=0.325
r155 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r156 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r157 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r158 108 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=13.68 $Y2=0
r159 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r160 105 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.785 $Y=0
+ $X2=13.62 $Y2=0
r161 105 107 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.785 $Y=0
+ $X2=14.16 $Y2=0
r162 104 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=13.68 $Y2=0
r163 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r164 101 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=13.2 $Y2=0
r165 101 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r166 100 103 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=12.24 $Y=0
+ $X2=13.2 $Y2=0
r167 100 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r168 98 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.955 $Y=0
+ $X2=11.79 $Y2=0
r169 98 100 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=11.955 $Y=0
+ $X2=12.24 $Y2=0
r170 97 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.455 $Y=0
+ $X2=13.62 $Y2=0
r171 97 103 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=13.455 $Y=0
+ $X2=13.2 $Y2=0
r172 96 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r173 96 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r174 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r175 93 125 8.42348 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=10.895 $Y=0
+ $X2=10.59 $Y2=0
r176 93 95 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.895 $Y=0
+ $X2=11.28 $Y2=0
r177 92 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.625 $Y=0
+ $X2=11.79 $Y2=0
r178 92 95 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=11.625 $Y=0
+ $X2=11.28 $Y2=0
r179 91 126 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=10.32 $Y2=0
r180 91 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r181 90 122 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=8.4 $Y=0
+ $X2=8.295 $Y2=0
r182 90 91 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r183 87 125 8.42348 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=10.285 $Y=0
+ $X2=10.59 $Y2=0
r184 87 90 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=10.285 $Y=0
+ $X2=8.4 $Y2=0
r185 86 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r186 85 119 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=7.44 $Y=0 $X2=7.5
+ $Y2=0
r187 85 86 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r188 82 85 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r189 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r190 79 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r191 78 79 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r192 76 79 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r193 76 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r194 75 78 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r195 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r196 73 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.71 $Y=0
+ $X2=3.545 $Y2=0
r197 73 75 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.71 $Y=0 $X2=4.08
+ $Y2=0
r198 72 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r199 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r200 69 114 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.38 $Y=0
+ $X2=3.545 $Y2=0
r201 69 71 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.38 $Y=0 $X2=3.12
+ $Y2=0
r202 68 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r203 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r204 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r205 65 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r206 64 67 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r207 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r208 62 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0
+ $X2=0.78 $Y2=0
r209 62 64 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.2
+ $Y2=0
r210 60 112 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r211 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r212 57 111 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.78 $Y2=0
r213 57 59 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=0
+ $X2=0.24 $Y2=0
r214 55 86 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=0 $X2=7.44
+ $Y2=0
r215 55 83 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.2 $Y=0 $X2=6.48
+ $Y2=0
r216 53 78 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=6.02 $Y=0 $X2=6 $Y2=0
r217 53 54 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=6.02 $Y=0 $X2=6.195
+ $Y2=0
r218 52 82 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.37 $Y=0 $X2=6.48
+ $Y2=0
r219 52 54 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=6.37 $Y=0 $X2=6.195
+ $Y2=0
r220 50 67 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=0
+ $X2=2.16 $Y2=0
r221 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=0 $X2=2.49
+ $Y2=0
r222 49 71 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.655 $Y=0
+ $X2=3.12 $Y2=0
r223 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=0 $X2=2.49
+ $Y2=0
r224 45 136 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.62 $Y=0.085
+ $X2=13.62 $Y2=0
r225 45 47 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=13.62 $Y=0.085
+ $X2=13.62 $Y2=0.515
r226 41 133 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.79 $Y=0.085
+ $X2=11.79 $Y2=0
r227 41 43 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=11.79 $Y=0.085
+ $X2=11.79 $Y2=0.515
r228 37 54 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.195 $Y=0.085
+ $X2=6.195 $Y2=0
r229 37 39 13.0061 $w=3.48e-07 $l=3.95e-07 $layer=LI1_cond $X=6.195 $Y=0.085
+ $X2=6.195 $Y2=0.48
r230 33 114 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.545 $Y=0.085
+ $X2=3.545 $Y2=0
r231 33 35 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=3.545 $Y=0.085
+ $X2=3.545 $Y2=0.505
r232 29 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=0.085
+ $X2=2.49 $Y2=0
r233 29 31 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.49 $Y=0.085
+ $X2=2.49 $Y2=0.55
r234 25 111 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0
r235 25 27 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.78 $Y=0.085
+ $X2=0.78 $Y2=0.565
r236 8 47 91 $w=1.7e-07 $l=4.26907e-07 $layer=licon1_NDIFF $count=2 $X=13.215
+ $Y=0.56 $X2=13.62 $Y2=0.515
r237 7 43 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=11.645
+ $Y=0.37 $X2=11.79 $Y2=0.515
r238 6 130 91 $w=1.7e-07 $l=5.57808e-07 $layer=licon1_NDIFF $count=2 $X=10.31
+ $Y=0.37 $X2=10.8 $Y2=0.515
r239 5 121 91 $w=1.7e-07 $l=7.78604e-07 $layer=licon1_NDIFF $count=2 $X=7.445
+ $Y=0.37 $X2=8.13 $Y2=0.57
r240 4 39 182 $w=1.7e-07 $l=2.79643e-07 $layer=licon1_NDIFF $count=1 $X=5.965
+ $Y=0.37 $X2=6.195 $Y2=0.48
r241 3 35 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=3.405
+ $Y=0.37 $X2=3.545 $Y2=0.505
r242 2 31 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.35 $Y=0.37
+ $X2=2.49 $Y2=0.55
r243 1 27 182 $w=1.7e-07 $l=2.91633e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.78 $Y2=0.565
.ends


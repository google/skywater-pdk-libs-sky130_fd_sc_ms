* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__sdfstp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
M1000 a_1686_74# a_998_81# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=1.66425e+12p ps=1.358e+07u
M1001 a_1764_74# a_800_74# a_1686_74# VNB nlowvt w=640000u l=150000u
+  ad=3.547e+11p pd=2.44e+06u as=0p ps=0u
M1002 a_998_81# a_800_74# a_292_464# VPB pshort w=420000u l=180000u
+  ad=1.344e+11p pd=1.48e+06u as=4.056e+11p ps=3.58e+06u
M1003 a_238_74# a_27_464# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1004 VGND SCD a_402_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1005 a_402_74# SCE a_292_464# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.373e+11p ps=2.81e+06u
M1006 VGND CLK a_599_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1007 a_1613_341# a_998_81# VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.35e+11p pd=5.07e+06u as=2.003e+12p ps=1.815e+07u
M1008 a_1988_74# a_1958_48# a_1910_74# VNB nlowvt w=420000u l=150000u
+  ad=3.192e+11p pd=2.36e+06u as=1.008e+11p ps=1.32e+06u
M1009 VGND a_1198_55# a_1150_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1010 a_1131_457# a_599_74# a_998_81# VPB pshort w=420000u l=180000u
+  ad=1.407e+11p pd=1.51e+06u as=0p ps=0u
M1011 a_1150_81# a_800_74# a_998_81# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=2.562e+11p ps=2.06e+06u
M1012 VGND SET_B a_1426_118# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1013 a_418_464# a_27_464# a_292_464# VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1014 a_998_81# a_599_74# a_292_464# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_800_74# a_599_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1016 a_1613_341# a_599_74# a_1764_74# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=4.18e+11p ps=4.14e+06u
M1017 VPWR SCE a_27_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=1.76e+11p ps=1.83e+06u
M1018 a_208_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1019 VPWR SCD a_418_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_1198_55# a_1131_457# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Q a_2395_112# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1022 VGND SET_B a_1988_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q a_2395_112# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1024 VPWR SET_B a_1198_55# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1025 VGND SCE a_27_464# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1026 VPWR a_1958_48# a_1721_374# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=3.655e+11p ps=4.42e+06u
M1027 VPWR a_1764_74# a_2395_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.268e+11p ps=2.22e+06u
M1028 a_292_464# D a_208_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR CLK a_599_74# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1030 a_1198_55# a_998_81# VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1764_74# SET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1426_118# a_998_81# a_1198_55# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1033 a_800_74# a_599_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.908e+11p pd=2.8e+06u as=0p ps=0u
M1034 a_292_464# D a_238_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VPWR a_1764_74# a_1958_48# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1036 VGND a_1764_74# a_2395_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=3.85e+11p ps=2.5e+06u
M1037 a_1910_74# a_599_74# a_1764_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_1764_74# a_800_74# a_1721_374# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_1958_48# a_1764_74# VGND VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
.ends

* File: sky130_fd_sc_ms__or4_2.spice
* Created: Fri Aug 28 18:08:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__or4_2.pex.spice"
.subckt sky130_fd_sc_ms__or4_2  VNB VPB D C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1004 N_A_85_392#_M1004_d N_D_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.284075 PD=0.92 PS=2.19 NRD=0 NRS=21.552 M=1 R=4.26667
+ SA=75000.4 SB=75002.9 A=0.096 P=1.58 MULT=1
MM1006 N_VGND_M1006_d N_C_M1006_g N_A_85_392#_M1004_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.1943 AS=0.0896 PD=1.255 PS=0.92 NRD=29.052 NRS=0 M=1 R=4.26667 SA=75000.8
+ SB=75002.5 A=0.096 P=1.58 MULT=1
MM1002 N_A_85_392#_M1002_d N_B_M1002_g N_VGND_M1006_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1943 PD=0.92 PS=1.255 NRD=0 NRS=29.052 M=1 R=4.26667 SA=75001.5
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1005 N_VGND_M1005_d N_A_M1005_g N_A_85_392#_M1002_d VNB NLOWVT L=0.15 W=0.64
+ AD=0.16742 AS=0.0896 PD=1.17333 PS=0.92 NRD=24.372 NRS=0 M=1 R=4.26667
+ SA=75002 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1003 N_X_M1003_d N_A_85_392#_M1003_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.19358 PD=1.02 PS=1.35667 NRD=0 NRS=18.648 M=1 R=4.93333
+ SA=75002.3 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1007 N_X_M1003_d N_A_85_392#_M1007_g N_VGND_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75002.7
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1010 A_177_392# N_D_M1010_g N_A_85_392#_M1010_s VPB PSHORT L=0.18 W=1 AD=0.12
+ AS=0.28 PD=1.24 PS=2.56 NRD=12.7853 NRS=0 M=1 R=5.55556 SA=90000.2 SB=90002.7
+ A=0.18 P=2.36 MULT=1
MM1000 A_261_392# N_C_M1000_g A_177_392# VPB PSHORT L=0.18 W=1 AD=0.12 AS=0.12
+ PD=1.24 PS=1.24 NRD=12.7853 NRS=12.7853 M=1 R=5.55556 SA=90000.6 SB=90002.3
+ A=0.18 P=2.36 MULT=1
MM1001 A_345_392# N_B_M1001_g A_261_392# VPB PSHORT L=0.18 W=1 AD=0.2 AS=0.12
+ PD=1.4 PS=1.24 NRD=28.5453 NRS=12.7853 M=1 R=5.55556 SA=90001 SB=90001.9
+ A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1011_d N_A_M1011_g A_345_392# VPB PSHORT L=0.18 W=1 AD=0.209717
+ AS=0.2 PD=1.43868 PS=1.4 NRD=15.7403 NRS=28.5453 M=1 R=5.55556 SA=90001.6
+ SB=90001.3 A=0.18 P=2.36 MULT=1
MM1008 N_X_M1008_d N_A_85_392#_M1008_g N_VPWR_M1011_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.234883 PD=1.39 PS=1.61132 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90002 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1009 N_X_M1008_d N_A_85_392#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3696 PD=1.39 PS=2.9 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90002.4
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8492 P=12.16
*
.include "sky130_fd_sc_ms__or4_2.pxi.spice"
*
.ends
*
*

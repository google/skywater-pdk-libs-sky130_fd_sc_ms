* File: sky130_fd_sc_ms__dfbbn_2.spice
* Created: Fri Aug 28 17:21:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__dfbbn_2.pex.spice"
.subckt sky130_fd_sc_ms__dfbbn_2  VNB VPB CLK_N D SET_B RESET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* D	D
* CLK_N	CLK_N
* VPB	VPB
* VNB	VNB
MM1037 N_VGND_M1037_d N_CLK_N_M1037_g N_A_27_74#_M1037_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1038 N_A_200_74#_M1038_d N_A_27_74#_M1038_g N_VGND_M1037_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1017_d N_D_M1017_g N_A_311_119#_M1017_s VNB NLOWVT L=0.15 W=0.42
+ AD=0.133562 AS=0.1197 PD=1.08 PS=1.41 NRD=32.856 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1036 A_529_119# N_A_473_405#_M1036_g N_VGND_M1017_d VNB NLOWVT L=0.15 W=0.42
+ AD=0.0441 AS=0.133562 PD=0.63 PS=1.08 NRD=14.28 NRS=34.284 M=1 R=2.8
+ SA=75000.9 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1042 N_A_601_119#_M1042_d N_A_27_74#_M1042_g A_529_119# VNB NLOWVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1028 N_A_311_119#_M1028_d N_A_200_74#_M1028_g N_A_601_119#_M1042_d VNB NLOWVT
+ L=0.15 W=0.42 AD=0.38115 AS=0.0588 PD=2.52 PS=0.7 NRD=243.564 NRS=0 M=1 R=2.8
+ SA=75001.7 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1040 N_A_473_405#_M1040_d N_A_601_119#_M1040_g N_A_867_125#_M1040_s VNB NLOWVT
+ L=0.15 W=0.55 AD=0.077 AS=0.15675 PD=0.83 PS=1.67 NRD=0 NRS=0 M=1 R=3.66667
+ SA=75000.2 SB=75004.7 A=0.0825 P=1.4 MULT=1
MM1007 N_A_867_125#_M1007_d N_A_975_322#_M1007_g N_A_473_405#_M1040_d VNB NLOWVT
+ L=0.15 W=0.55 AD=0.09625 AS=0.077 PD=0.9 PS=0.83 NRD=15.264 NRS=0 M=1
+ R=3.66667 SA=75000.6 SB=75004.3 A=0.0825 P=1.4 MULT=1
MM1005 N_VGND_M1005_d N_SET_B_M1005_g N_A_867_125#_M1007_d VNB NLOWVT L=0.15
+ W=0.55 AD=0.09625 AS=0.09625 PD=0.9 PS=0.9 NRD=15.264 NRS=0 M=1 R=3.66667
+ SA=75001.1 SB=75003.8 A=0.0825 P=1.4 MULT=1
MM1003 A_1240_125# N_A_473_405#_M1003_g N_VGND_M1005_d VNB NLOWVT L=0.15 W=0.55
+ AD=0.0950625 AS=0.09625 PD=0.94 PS=0.9 NRD=25.704 NRS=0 M=1 R=3.66667
+ SA=75001.6 SB=75003.3 A=0.0825 P=1.4 MULT=1
MM1039 N_A_1335_112#_M1039_d N_A_27_74#_M1039_g A_1240_125# VNB NLOWVT L=0.15
+ W=0.55 AD=0.345876 AS=0.0950625 PD=2.18299 PS=0.94 NRD=0 NRS=25.704 M=1
+ R=3.66667 SA=75001.9 SB=75002.8 A=0.0825 P=1.4 MULT=1
MM1004 A_1640_138# N_A_200_74#_M1004_g N_A_1335_112#_M1039_d VNB NLOWVT L=0.15
+ W=0.42 AD=0.0504 AS=0.264124 PD=0.66 PS=1.66701 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75003.6 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_A_1555_410#_M1023_g A_1640_138# VNB NLOWVT L=0.15 W=0.42
+ AD=0.0968897 AS=0.0504 PD=0.84 PS=0.66 NRD=50.196 NRS=18.564 M=1 R=2.8
+ SA=75004 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1010 N_A_1832_74#_M1010_d N_SET_B_M1010_g N_VGND_M1023_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.17071 PD=1.02 PS=1.48 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.7 SB=75001.2 A=0.111 P=1.78 MULT=1
MM1024 N_A_1555_410#_M1024_d N_A_975_322#_M1024_g N_A_1832_74#_M1010_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.1184 AS=0.1036 PD=1.06 PS=1.02 NRD=6.48 NRS=0 M=1
+ R=4.93333 SA=75003.1 SB=75000.8 A=0.111 P=1.78 MULT=1
MM1009 N_A_1832_74#_M1009_d N_A_1335_112#_M1009_g N_A_1555_410#_M1024_d VNB
+ NLOWVT L=0.15 W=0.74 AD=0.2907 AS=0.1184 PD=2.39 PS=1.06 NRD=12.972 NRS=0 M=1
+ R=4.93333 SA=75003.6 SB=75000.3 A=0.111 P=1.78 MULT=1
MM1026 N_VGND_M1026_d N_RESET_B_M1026_g N_A_975_322#_M1026_s VNB NLOWVT L=0.15
+ W=0.42 AD=0.171892 AS=0.1176 PD=1.45552 PS=1.4 NRD=101.208 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1035 N_VGND_M1026_d N_A_1555_410#_M1035_g N_Q_N_M1035_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.302858 AS=0.1036 PD=2.56448 PS=1.02 NRD=57.444 NRS=0 M=1 R=4.93333
+ SA=75000.5 SB=75000.7 A=0.111 P=1.78 MULT=1
MM1043 N_VGND_M1043_d N_A_1555_410#_M1043_g N_Q_N_M1035_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.222 AS=0.1036 PD=2.08 PS=1.02 NRD=2.424 NRS=0 M=1 R=4.93333
+ SA=75000.9 SB=75000.2 A=0.111 P=1.78 MULT=1
MM1031 N_VGND_M1031_d N_A_1555_410#_M1031_g N_A_2516_368#_M1031_s VNB NLOWVT
+ L=0.15 W=0.64 AD=0.108058 AS=0.1824 PD=0.987826 PS=1.85 NRD=5.616 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1008 N_Q_M1008_d N_A_2516_368#_M1008_g N_VGND_M1031_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.124942 PD=1.02 PS=1.14217 NRD=0 NRS=2.424 M=1 R=4.93333
+ SA=75000.6 SB=75000.6 A=0.111 P=1.78 MULT=1
MM1032 N_Q_M1008_d N_A_2516_368#_M1032_g N_VGND_M1032_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1998 PD=1.02 PS=2.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1033 N_VPWR_M1033_d N_CLK_N_M1033_g N_A_27_74#_M1033_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3024 PD=1.39 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.2 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1034 N_A_200_74#_M1034_d N_A_27_74#_M1034_g N_VPWR_M1033_d VPB PSHORT L=0.18
+ W=1.12 AD=0.2968 AS=0.1512 PD=2.77 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.6 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1025 N_VPWR_M1025_d N_D_M1025_g N_A_311_119#_M1025_s VPB PSHORT L=0.18 W=0.42
+ AD=0.08715 AS=0.17175 PD=0.835 PS=1.72 NRD=65.6601 NRS=39.8531 M=1 R=2.33333
+ SA=90000.3 SB=90001.8 A=0.0756 P=1.2 MULT=1
MM1018 A_539_503# N_A_473_405#_M1018_g N_VPWR_M1025_d VPB PSHORT L=0.18 W=0.42
+ AD=0.0504 AS=0.08715 PD=0.66 PS=0.835 NRD=30.4759 NRS=0 M=1 R=2.33333
+ SA=90000.9 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1030 N_A_601_119#_M1030_d N_A_200_74#_M1030_g A_539_503# VPB PSHORT L=0.18
+ W=0.42 AD=0.0693 AS=0.0504 PD=0.75 PS=0.66 NRD=11.7215 NRS=30.4759 M=1
+ R=2.33333 SA=90001.3 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1011 N_A_311_119#_M1011_d N_A_27_74#_M1011_g N_A_601_119#_M1030_d VPB PSHORT
+ L=0.18 W=0.42 AD=0.159 AS=0.0693 PD=1.67 PS=0.75 NRD=30.4759 NRS=11.7215 M=1
+ R=2.33333 SA=90001.8 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1006 A_933_424# N_A_601_119#_M1006_g N_A_473_405#_M1006_s VPB PSHORT L=0.18
+ W=0.84 AD=0.1008 AS=0.2226 PD=1.08 PS=2.21 NRD=15.2281 NRS=0 M=1 R=4.66667
+ SA=90000.2 SB=90001.1 A=0.1512 P=2.04 MULT=1
MM1029 N_VPWR_M1029_d N_A_975_322#_M1029_g A_933_424# VPB PSHORT L=0.18 W=0.84
+ AD=0.1386 AS=0.1008 PD=1.17 PS=1.08 NRD=0 NRS=15.2281 M=1 R=4.66667 SA=90000.6
+ SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1014 N_A_473_405#_M1014_d N_SET_B_M1014_g N_VPWR_M1029_d VPB PSHORT L=0.18
+ W=0.84 AD=0.2226 AS=0.1386 PD=2.21 PS=1.17 NRD=0 NRS=12.8838 M=1 R=4.66667
+ SA=90001.1 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1041 A_1315_424# N_A_473_405#_M1041_g N_VPWR_M1041_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1008 AS=0.2226 PD=1.08 PS=2.21 NRD=15.2281 NRS=0 M=1 R=4.66667 SA=90000.2
+ SB=90001.1 A=0.1512 P=2.04 MULT=1
MM1022 N_A_1335_112#_M1022_d N_A_200_74#_M1022_g A_1315_424# VPB PSHORT L=0.18
+ W=0.84 AD=0.1792 AS=0.1008 PD=1.6 PS=1.08 NRD=0 NRS=15.2281 M=1 R=4.66667
+ SA=90000.6 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1002 A_1507_508# N_A_27_74#_M1002_g N_A_1335_112#_M1022_d VPB PSHORT L=0.18
+ W=0.42 AD=0.0504 AS=0.0896 PD=0.66 PS=0.8 NRD=30.4759 NRS=39.8531 M=1
+ R=2.33333 SA=90001.1 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1013 N_VPWR_M1013_d N_A_1555_410#_M1013_g A_1507_508# VPB PSHORT L=0.18 W=0.42
+ AD=0.22145 AS=0.0504 PD=2.04 PS=0.66 NRD=221.507 NRS=30.4759 M=1 R=2.33333
+ SA=90001.6 SB=90000.3 A=0.0756 P=1.2 MULT=1
MM1027 N_VPWR_M1027_d N_SET_B_M1027_g N_A_1555_410#_M1027_s VPB PSHORT L=0.18
+ W=1 AD=0.254075 AS=0.28 PD=1.675 PS=2.56 NRD=39.203 NRS=0 M=1 R=5.55556
+ SA=90000.2 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1021 A_1934_392# N_A_975_322#_M1021_g N_VPWR_M1027_d VPB PSHORT L=0.18 W=1
+ AD=0.12 AS=0.254075 PD=1.24 PS=1.675 NRD=12.7853 NRS=39.203 M=1 R=5.55556
+ SA=90000.8 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1000 N_A_1555_410#_M1000_d N_A_1335_112#_M1000_g A_1934_392# VPB PSHORT L=0.18
+ W=1 AD=0.265 AS=0.12 PD=2.53 PS=1.24 NRD=0 NRS=12.7853 M=1 R=5.55556
+ SA=90001.2 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_RESET_B_M1012_g N_A_975_322#_M1012_s VPB PSHORT L=0.18
+ W=0.64 AD=0.127418 AS=0.1696 PD=1.06545 PS=1.81 NRD=44.3447 NRS=0 M=1
+ R=3.55556 SA=90000.2 SB=90001.1 A=0.1152 P=1.64 MULT=1
MM1015 N_Q_N_M1015_d N_A_1555_410#_M1015_g N_VPWR_M1012_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.222982 PD=1.39 PS=1.86455 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.5 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1019 N_Q_N_M1015_d N_A_1555_410#_M1019_g N_VPWR_M1019_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.2968 PD=1.39 PS=2.77 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90000.9 SB=90000.2 A=0.2016 P=2.6 MULT=1
MM1001 N_VPWR_M1001_d N_A_1555_410#_M1001_g N_A_2516_368#_M1001_s VPB PSHORT
+ L=0.18 W=1 AD=0.175377 AS=0.265 PD=1.37736 PS=2.53 NRD=12.7853 NRS=0 M=1
+ R=5.55556 SA=90000.2 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1016 N_Q_M1016_d N_A_2516_368#_M1016_g N_VPWR_M1001_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.196423 PD=1.39 PS=1.54264 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1020 N_Q_M1016_d N_A_2516_368#_M1020_g N_VPWR_M1020_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3024 PD=1.39 PS=2.78 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX44_noxref VNB VPB NWDIODE A=27.4908 P=33.28
c_297 VPB 0 4.37917e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_ms__dfbbn_2.pxi.spice"
*
.ends
*
*

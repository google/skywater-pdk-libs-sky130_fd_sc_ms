* File: sky130_fd_sc_ms__mux4_4.pex.spice
* Created: Fri Aug 28 17:41:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__MUX4_4%A1 3 7 11 15 17 18 28
c43 18 0 8.41401e-20 $X=0.72 $Y=1.665
r44 27 28 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=0.925 $Y=1.615
+ $X2=0.955 $Y2=1.615
r45 25 27 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=0.725 $Y=1.615
+ $X2=0.925 $Y2=1.615
r46 23 25 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=0.505 $Y=1.615
+ $X2=0.725 $Y2=1.615
r47 21 23 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.495 $Y=1.615
+ $X2=0.505 $Y2=1.615
r48 18 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.725
+ $Y=1.615 $X2=0.725 $Y2=1.615
r49 17 18 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.615
+ $X2=0.72 $Y2=1.615
r50 13 28 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.955 $Y=1.78
+ $X2=0.955 $Y2=1.615
r51 13 15 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=0.955 $Y=1.78
+ $X2=0.955 $Y2=2.46
r52 9 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.45
+ $X2=0.925 $Y2=1.615
r53 9 11 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=0.925 $Y=1.45 $X2=0.925
+ $Y2=0.95
r54 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.45
+ $X2=0.495 $Y2=1.615
r55 5 7 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=0.495 $Y=1.45 $X2=0.495
+ $Y2=0.95
r56 1 23 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.78
+ $X2=0.505 $Y2=1.615
r57 1 3 264.323 $w=1.8e-07 $l=6.8e-07 $layer=POLY_cond $X=0.505 $Y=1.78
+ $X2=0.505 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%A0 3 7 11 15 17 18 19 23 25
c60 25 0 1.04993e-19 $X=2.19 $Y=1.635
c61 11 0 7.75212e-20 $X=1.85 $Y=0.95
c62 7 0 8.41401e-20 $X=1.42 $Y=0.95
c63 3 0 2.67665e-19 $X=1.405 $Y=2.46
r64 34 35 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=1.85 $Y=1.635
+ $X2=1.905 $Y2=1.635
r65 32 34 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.51 $Y=1.635
+ $X2=1.85 $Y2=1.635
r66 32 33 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.51
+ $Y=1.635 $X2=1.51 $Y2=1.635
r67 30 32 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.42 $Y=1.635 $X2=1.51
+ $Y2=1.635
r68 28 30 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.405 $Y=1.635
+ $X2=1.42 $Y2=1.635
r69 23 35 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.995 $Y=1.635
+ $X2=1.905 $Y2=1.635
r70 23 25 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.995 $Y=1.635
+ $X2=2.19 $Y2=1.635
r71 19 25 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.19
+ $Y=1.635 $X2=2.19 $Y2=1.635
r72 18 19 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.635
+ $X2=2.16 $Y2=1.635
r73 18 33 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.68 $Y=1.635
+ $X2=1.51 $Y2=1.635
r74 17 33 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.2 $Y=1.635 $X2=1.51
+ $Y2=1.635
r75 13 35 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.8
+ $X2=1.905 $Y2=1.635
r76 13 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.905 $Y=1.8
+ $X2=1.905 $Y2=2.46
r77 9 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.85 $Y=1.47
+ $X2=1.85 $Y2=1.635
r78 9 11 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.85 $Y=1.47 $X2=1.85
+ $Y2=0.95
r79 5 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.42 $Y=1.47
+ $X2=1.42 $Y2=1.635
r80 5 7 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.42 $Y=1.47 $X2=1.42
+ $Y2=0.95
r81 1 28 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.8
+ $X2=1.405 $Y2=1.635
r82 1 3 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=1.405 $Y=1.8 $X2=1.405
+ $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%A_758_306# 1 2 9 13 17 21 24 25 27 30 32 34
+ 37 45 49 55 57 62 66 67 69 76
c134 57 0 1.30567e-19 $X=6.54 $Y=1.53
c135 32 0 7.8786e-20 $X=6.745 $Y=1.365
c136 21 0 1.75061e-19 $X=4.335 $Y=0.915
r137 75 76 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=6.745 $Y=1.53
+ $X2=6.8 $Y2=1.53
r138 71 73 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=6.315 $Y=1.53
+ $X2=6.35 $Y2=1.53
r139 66 67 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=5.2 $Y=1.45
+ $X2=6.035 $Y2=1.45
r140 65 66 7.06528 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=5.075 $Y=1.515
+ $X2=5.2 $Y2=1.515
r141 64 65 0.104768 $w=3.28e-07 $l=3e-09 $layer=LI1_cond $X=5.072 $Y=1.515
+ $X2=5.075 $Y2=1.515
r142 62 69 31.258 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.875 $Y=1.515
+ $X2=4.71 $Y2=1.515
r143 61 64 6.87974 $w=3.28e-07 $l=1.97e-07 $layer=LI1_cond $X=4.875 $Y=1.515
+ $X2=5.072 $Y2=1.515
r144 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.875
+ $Y=1.515 $X2=4.875 $Y2=1.515
r145 58 75 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=6.54 $Y=1.53
+ $X2=6.745 $Y2=1.53
r146 58 73 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=6.54 $Y=1.53
+ $X2=6.35 $Y2=1.53
r147 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.54
+ $Y=1.53 $X2=6.54 $Y2=1.53
r148 55 67 14.2244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=6.365 $Y=1.53
+ $X2=6.035 $Y2=1.53
r149 55 57 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=6.365 $Y=1.53
+ $X2=6.54 $Y2=1.53
r150 49 51 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=5.075 $Y=1.985
+ $X2=5.075 $Y2=2.815
r151 47 65 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=5.075 $Y=1.68
+ $X2=5.075 $Y2=1.515
r152 47 49 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=5.075 $Y=1.68
+ $X2=5.075 $Y2=1.985
r153 43 64 2.26808 $w=2.55e-07 $l=1.65e-07 $layer=LI1_cond $X=5.072 $Y=1.35
+ $X2=5.072 $Y2=1.515
r154 43 45 37.7369 $w=2.53e-07 $l=8.35e-07 $layer=LI1_cond $X=5.072 $Y=1.35
+ $X2=5.072 $Y2=0.515
r155 41 42 0.937743 $w=2.57e-07 $l=5e-09 $layer=POLY_cond $X=4.33 $Y=1.547
+ $X2=4.335 $Y2=1.547
r156 40 41 79.7082 $w=2.57e-07 $l=4.25e-07 $layer=POLY_cond $X=3.905 $Y=1.547
+ $X2=4.33 $Y2=1.547
r157 39 40 4.68872 $w=2.57e-07 $l=2.5e-08 $layer=POLY_cond $X=3.88 $Y=1.547
+ $X2=3.905 $Y2=1.547
r158 35 76 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.8 $Y=1.695
+ $X2=6.8 $Y2=1.53
r159 35 37 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=6.8 $Y=1.695 $X2=6.8
+ $Y2=2.385
r160 32 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.745 $Y=1.365
+ $X2=6.745 $Y2=1.53
r161 32 34 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=6.745 $Y=1.365
+ $X2=6.745 $Y2=0.925
r162 28 73 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.35 $Y=1.695
+ $X2=6.35 $Y2=1.53
r163 28 30 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=6.35 $Y=1.695
+ $X2=6.35 $Y2=2.385
r164 25 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.315 $Y=1.365
+ $X2=6.315 $Y2=1.53
r165 25 27 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=6.315 $Y=1.365
+ $X2=6.315 $Y2=0.925
r166 24 42 15.4604 $w=2.65e-07 $l=8.5e-08 $layer=POLY_cond $X=4.42 $Y=1.547
+ $X2=4.335 $Y2=1.547
r167 24 69 65.646 $w=2.65e-07 $l=2.9e-07 $layer=POLY_cond $X=4.42 $Y=1.547
+ $X2=4.71 $Y2=1.547
r168 19 42 15.359 $w=1.5e-07 $l=1.32e-07 $layer=POLY_cond $X=4.335 $Y=1.415
+ $X2=4.335 $Y2=1.547
r169 19 21 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=4.335 $Y=1.415
+ $X2=4.335 $Y2=0.915
r170 15 41 11.1533 $w=1.8e-07 $l=1.33e-07 $layer=POLY_cond $X=4.33 $Y=1.68
+ $X2=4.33 $Y2=1.547
r171 15 17 303.194 $w=1.8e-07 $l=7.8e-07 $layer=POLY_cond $X=4.33 $Y=1.68
+ $X2=4.33 $Y2=2.46
r172 11 40 15.359 $w=1.5e-07 $l=1.32e-07 $layer=POLY_cond $X=3.905 $Y=1.415
+ $X2=3.905 $Y2=1.547
r173 11 13 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.905 $Y=1.415
+ $X2=3.905 $Y2=0.915
r174 7 39 11.1533 $w=1.8e-07 $l=1.33e-07 $layer=POLY_cond $X=3.88 $Y=1.68
+ $X2=3.88 $Y2=1.547
r175 7 9 303.194 $w=1.8e-07 $l=7.8e-07 $layer=POLY_cond $X=3.88 $Y=1.68 $X2=3.88
+ $Y2=2.46
r176 2 51 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=4.97
+ $Y=1.84 $X2=5.115 $Y2=2.815
r177 2 49 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.97
+ $Y=1.84 $X2=5.115 $Y2=1.985
r178 1 45 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=4.965
+ $Y=0.37 $X2=5.11 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%S0 3 8 9 10 13 18 19 24 25 27 29 33 37 41 45
+ 48 50 52 53 54 56 57 58 59 63
c173 59 0 1.54503e-19 $X=8.4 $Y=1.665
c174 41 0 1.64187e-19 $X=7.605 $Y=0.925
c175 37 0 4.1337e-20 $X=7.25 $Y=2.385
c176 33 0 2.75222e-19 $X=7.175 $Y=0.925
r177 72 73 14.5828 $w=3.14e-07 $l=9.5e-08 $layer=POLY_cond $X=7.605 $Y=1.56
+ $X2=7.7 $Y2=1.56
r178 70 72 22.258 $w=3.14e-07 $l=1.45e-07 $layer=POLY_cond $X=7.46 $Y=1.56
+ $X2=7.605 $Y2=1.56
r179 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.46
+ $Y=1.56 $X2=7.46 $Y2=1.56
r180 68 70 32.2357 $w=3.14e-07 $l=2.1e-07 $layer=POLY_cond $X=7.25 $Y=1.56
+ $X2=7.46 $Y2=1.56
r181 67 68 11.5127 $w=3.14e-07 $l=7.5e-08 $layer=POLY_cond $X=7.175 $Y=1.56
+ $X2=7.25 $Y2=1.56
r182 65 66 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.14
+ $Y=1.56 $X2=8.14 $Y2=1.56
r183 63 73 13.3045 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.79 $Y=1.56 $X2=7.7
+ $Y2=1.56
r184 63 65 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=7.79 $Y=1.56
+ $X2=8.14 $Y2=1.56
r185 59 66 8.8128 $w=3.38e-07 $l=2.6e-07 $layer=LI1_cond $X=8.4 $Y=1.605
+ $X2=8.14 $Y2=1.605
r186 58 66 7.45698 $w=3.38e-07 $l=2.2e-07 $layer=LI1_cond $X=7.92 $Y=1.605
+ $X2=8.14 $Y2=1.605
r187 58 71 15.5919 $w=3.38e-07 $l=4.6e-07 $layer=LI1_cond $X=7.92 $Y=1.605
+ $X2=7.46 $Y2=1.605
r188 57 71 0.677908 $w=3.38e-07 $l=2e-08 $layer=LI1_cond $X=7.44 $Y=1.605
+ $X2=7.46 $Y2=1.605
r189 56 65 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=8.155 $Y=1.56
+ $X2=8.14 $Y2=1.56
r190 51 52 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.432 $Y=1.31
+ $X2=3.432 $Y2=1.46
r191 49 50 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.957 $Y=1.31
+ $X2=2.957 $Y2=1.46
r192 48 56 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=8.23 $Y=1.395
+ $X2=8.155 $Y2=1.56
r193 47 48 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=8.23 $Y=0.255
+ $X2=8.23 $Y2=1.395
r194 43 73 15.7762 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.7 $Y=1.725
+ $X2=7.7 $Y2=1.56
r195 43 45 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=7.7 $Y=1.725
+ $X2=7.7 $Y2=2.385
r196 39 72 20.044 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.605 $Y=1.395
+ $X2=7.605 $Y2=1.56
r197 39 41 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=7.605 $Y=1.395
+ $X2=7.605 $Y2=0.925
r198 35 68 15.7762 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.25 $Y=1.725
+ $X2=7.25 $Y2=1.56
r199 35 37 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=7.25 $Y=1.725
+ $X2=7.25 $Y2=2.385
r200 31 67 20.044 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.175 $Y=1.395
+ $X2=7.175 $Y2=1.56
r201 31 33 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=7.175 $Y=1.395
+ $X2=7.175 $Y2=0.925
r202 30 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.4 $Y=0.18
+ $X2=5.325 $Y2=0.18
r203 29 47 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.155 $Y=0.18
+ $X2=8.23 $Y2=0.255
r204 29 30 1412.67 $w=1.5e-07 $l=2.755e-06 $layer=POLY_cond $X=8.155 $Y=0.18
+ $X2=5.4 $Y2=0.18
r205 25 55 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=5.34 $Y=1.275
+ $X2=5.34 $Y2=1.185
r206 25 27 437.298 $w=1.8e-07 $l=1.125e-06 $layer=POLY_cond $X=5.34 $Y=1.275
+ $X2=5.34 $Y2=2.4
r207 24 55 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.325 $Y=0.74
+ $X2=5.325 $Y2=1.185
r208 21 54 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.325 $Y=0.255
+ $X2=5.325 $Y2=0.18
r209 21 24 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=5.325 $Y=0.255
+ $X2=5.325 $Y2=0.74
r210 20 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.55 $Y=0.18
+ $X2=3.475 $Y2=0.18
r211 19 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.25 $Y=0.18
+ $X2=5.325 $Y2=0.18
r212 19 20 871.702 $w=1.5e-07 $l=1.7e-06 $layer=POLY_cond $X=5.25 $Y=0.18
+ $X2=3.55 $Y2=0.18
r213 18 51 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.475 $Y=0.915
+ $X2=3.475 $Y2=1.31
r214 15 53 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.475 $Y=0.255
+ $X2=3.475 $Y2=0.18
r215 15 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.475 $Y=0.255
+ $X2=3.475 $Y2=0.915
r216 13 52 388.71 $w=1.8e-07 $l=1e-06 $layer=POLY_cond $X=3.405 $Y=2.46
+ $X2=3.405 $Y2=1.46
r217 9 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.4 $Y=0.18
+ $X2=3.475 $Y2=0.18
r218 9 10 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=3.4 $Y=0.18
+ $X2=3.075 $Y2=0.18
r219 8 49 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3 $Y=0.915 $X2=3
+ $Y2=1.31
r220 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3 $Y=0.255
+ $X2=3.075 $Y2=0.18
r221 5 8 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3 $Y=0.255 $X2=3
+ $Y2=0.915
r222 3 50 388.71 $w=1.8e-07 $l=1e-06 $layer=POLY_cond $X=2.93 $Y=2.46 $X2=2.93
+ $Y2=1.46
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%A2 3 7 11 15 17 18 28
c59 28 0 9.16034e-20 $X=9.385 $Y=1.425
c60 15 0 1.66006e-19 $X=9.385 $Y=0.69
r61 26 28 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=9.27 $Y=1.425
+ $X2=9.385 $Y2=1.425
r62 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.27
+ $Y=1.425 $X2=9.27 $Y2=1.425
r63 24 26 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=9.245 $Y=1.425
+ $X2=9.27 $Y2=1.425
r64 23 24 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=8.955 $Y=1.425
+ $X2=9.245 $Y2=1.425
r65 21 23 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=8.795 $Y=1.425
+ $X2=8.955 $Y2=1.425
r66 18 27 2.09023 $w=5.13e-07 $l=9e-08 $layer=LI1_cond $X=9.36 $Y=1.517 $X2=9.27
+ $Y2=1.517
r67 17 27 9.05768 $w=5.13e-07 $l=3.9e-07 $layer=LI1_cond $X=8.88 $Y=1.517
+ $X2=9.27 $Y2=1.517
r68 13 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.385 $Y=1.26
+ $X2=9.385 $Y2=1.425
r69 13 15 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=9.385 $Y=1.26
+ $X2=9.385 $Y2=0.69
r70 9 24 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.245 $Y=1.59
+ $X2=9.245 $Y2=1.425
r71 9 11 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=9.245 $Y=1.59
+ $X2=9.245 $Y2=2.46
r72 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.955 $Y=1.26
+ $X2=8.955 $Y2=1.425
r73 5 7 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=8.955 $Y=1.26
+ $X2=8.955 $Y2=0.69
r74 1 21 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=8.795 $Y=1.59
+ $X2=8.795 $Y2=1.425
r75 1 3 338.177 $w=1.8e-07 $l=8.7e-07 $layer=POLY_cond $X=8.795 $Y=1.59
+ $X2=8.795 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%A3 3 7 9 11 14 17 20 22 23 31
c55 31 0 2.68867e-20 $X=10.325 $Y=1.61
c56 9 0 1.44963e-19 $X=10.245 $Y=1.085
r57 31 32 1.46951 $w=3.28e-07 $l=1e-08 $layer=POLY_cond $X=10.325 $Y=1.61
+ $X2=10.335 $Y2=1.61
r58 29 31 11.7561 $w=3.28e-07 $l=8e-08 $layer=POLY_cond $X=10.245 $Y=1.61
+ $X2=10.325 $Y2=1.61
r59 27 29 54.372 $w=3.28e-07 $l=3.7e-07 $layer=POLY_cond $X=9.875 $Y=1.61
+ $X2=10.245 $Y2=1.61
r60 26 27 8.81707 $w=3.28e-07 $l=6e-08 $layer=POLY_cond $X=9.815 $Y=1.61
+ $X2=9.875 $Y2=1.61
r61 23 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.245
+ $Y=1.61 $X2=10.245 $Y2=1.61
r62 22 23 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=9.84 $Y=1.61
+ $X2=10.245 $Y2=1.61
r63 18 20 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=10.245 $Y=1.16
+ $X2=10.335 $Y2=1.16
r64 17 32 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.335 $Y=1.445
+ $X2=10.335 $Y2=1.61
r65 16 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.335 $Y=1.235
+ $X2=10.335 $Y2=1.16
r66 16 17 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=10.335 $Y=1.235
+ $X2=10.335 $Y2=1.445
r67 12 31 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.325 $Y=1.775
+ $X2=10.325 $Y2=1.61
r68 12 14 266.266 $w=1.8e-07 $l=6.85e-07 $layer=POLY_cond $X=10.325 $Y=1.775
+ $X2=10.325 $Y2=2.46
r69 9 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.245 $Y=1.085
+ $X2=10.245 $Y2=1.16
r70 9 11 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=10.245 $Y=1.085
+ $X2=10.245 $Y2=0.69
r71 5 27 16.7902 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=9.875 $Y=1.775
+ $X2=9.875 $Y2=1.61
r72 5 7 266.266 $w=1.8e-07 $l=6.85e-07 $layer=POLY_cond $X=9.875 $Y=1.775
+ $X2=9.875 $Y2=2.46
r73 1 26 21.0783 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.815 $Y=1.445
+ $X2=9.815 $Y2=1.61
r74 1 3 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=9.815 $Y=1.445
+ $X2=9.815 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%S1 3 7 11 15 17 19 21 24 26 31 32 40 44 49 55
+ 56 58
c116 56 0 5.98463e-20 $X=12.665 $Y=1.455
c117 44 0 2.9352e-20 $X=12.315 $Y=1.36
c118 24 0 1.03922e-19 $X=14.3 $Y=2.4
c119 17 0 1.438e-19 $X=14.21 $Y=1.37
c120 15 0 8.44579e-20 $X=12.035 $Y=2.46
r121 55 56 1.63907 $w=6.48e-07 $l=5.5e-08 $layer=LI1_cond $X=12.72 $Y=1.455
+ $X2=12.665 $Y2=1.455
r122 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.315
+ $Y=1.36 $X2=12.315 $Y2=1.36
r123 40 58 9.28585 $w=6.48e-07 $l=1e-07 $layer=LI1_cond $X=12.735 $Y=1.455
+ $X2=12.835 $Y2=1.455
r124 40 55 0.276018 $w=6.48e-07 $l=1.5e-08 $layer=LI1_cond $X=12.735 $Y=1.455
+ $X2=12.72 $Y2=1.455
r125 40 56 0.355271 $w=5.03e-07 $l=1.5e-08 $layer=LI1_cond $X=12.65 $Y=1.527
+ $X2=12.665 $Y2=1.527
r126 40 45 7.93438 $w=5.03e-07 $l=3.35e-07 $layer=LI1_cond $X=12.65 $Y=1.527
+ $X2=12.315 $Y2=1.527
r127 38 49 29.4439 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.705 $Y=1.385
+ $X2=13.87 $Y2=1.385
r128 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.705
+ $Y=1.385 $X2=13.705 $Y2=1.385
r129 32 37 6.02816 $w=3.23e-07 $l=1.7e-07 $layer=LI1_cond $X=13.702 $Y=1.215
+ $X2=13.702 $Y2=1.385
r130 32 58 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=13.54 $Y=1.215
+ $X2=12.835 $Y2=1.215
r131 29 30 14.7551 $w=2.94e-07 $l=9e-08 $layer=POLY_cond $X=11.945 $Y=1.36
+ $X2=12.035 $Y2=1.36
r132 28 29 67.2177 $w=2.94e-07 $l=4.1e-07 $layer=POLY_cond $X=11.535 $Y=1.36
+ $X2=11.945 $Y2=1.36
r133 26 44 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=12.125 $Y=1.36
+ $X2=12.315 $Y2=1.36
r134 26 30 13.8324 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=12.125 $Y=1.36
+ $X2=12.035 $Y2=1.36
r135 22 31 32.4784 $w=1.65e-07 $l=1.5e-07 $layer=POLY_cond $X=14.3 $Y=1.52
+ $X2=14.3 $Y2=1.37
r136 22 24 342.065 $w=1.8e-07 $l=8.8e-07 $layer=POLY_cond $X=14.3 $Y=1.52
+ $X2=14.3 $Y2=2.4
r137 19 31 32.4784 $w=1.65e-07 $l=1.57321e-07 $layer=POLY_cond $X=14.285 $Y=1.22
+ $X2=14.3 $Y2=1.37
r138 19 21 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=14.285 $Y=1.22
+ $X2=14.285 $Y2=0.74
r139 17 31 2.73406 $w=3e-07 $l=9e-08 $layer=POLY_cond $X=14.21 $Y=1.37 $X2=14.3
+ $Y2=1.37
r140 17 49 67.9852 $w=3e-07 $l=3.4e-07 $layer=POLY_cond $X=14.21 $Y=1.37
+ $X2=13.87 $Y2=1.37
r141 13 30 14.2527 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=12.035 $Y=1.525
+ $X2=12.035 $Y2=1.36
r142 13 15 363.444 $w=1.8e-07 $l=9.35e-07 $layer=POLY_cond $X=12.035 $Y=1.525
+ $X2=12.035 $Y2=2.46
r143 9 29 18.4939 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.945 $Y=1.195
+ $X2=11.945 $Y2=1.36
r144 9 11 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=11.945 $Y=1.195
+ $X2=11.945 $Y2=0.69
r145 5 28 14.2527 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=11.535 $Y=1.525
+ $X2=11.535 $Y2=1.36
r146 5 7 363.444 $w=1.8e-07 $l=9.35e-07 $layer=POLY_cond $X=11.535 $Y=1.525
+ $X2=11.535 $Y2=2.46
r147 1 28 29.5102 $w=2.94e-07 $l=2.49199e-07 $layer=POLY_cond $X=11.355 $Y=1.195
+ $X2=11.535 $Y2=1.36
r148 1 3 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=11.355 $Y=1.195
+ $X2=11.355 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%A_2489_347# 1 2 7 9 12 14 16 19 21 25 30 32
+ 33 37 39
c85 33 0 4.75356e-20 $X=13.165 $Y=1.635
c86 32 0 2.68058e-20 $X=13.165 $Y=1.635
c87 30 0 2.3931e-20 $X=14.12 $Y=1.72
c88 21 0 1.438e-19 $X=13.875 $Y=1.805
c89 7 0 1.46885e-19 $X=12.535 $Y=1.885
r90 43 44 34.8434 $w=3.32e-07 $l=2.4e-07 $layer=POLY_cond $X=12.795 $Y=1.677
+ $X2=13.035 $Y2=1.677
r91 39 41 9.25293 $w=2.98e-07 $l=1.85e-07 $layer=LI1_cond $X=14.055 $Y=0.775
+ $X2=14.055 $Y2=0.96
r92 33 46 8.71084 $w=3.32e-07 $l=6e-08 $layer=POLY_cond $X=13.165 $Y=1.677
+ $X2=13.225 $Y2=1.677
r93 33 44 18.8735 $w=3.32e-07 $l=1.3e-07 $layer=POLY_cond $X=13.165 $Y=1.677
+ $X2=13.035 $Y2=1.677
r94 32 35 6.02816 $w=3.23e-07 $l=1.7e-07 $layer=LI1_cond $X=13.167 $Y=1.635
+ $X2=13.167 $Y2=1.805
r95 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.165
+ $Y=1.635 $X2=13.165 $Y2=1.635
r96 30 37 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=14.12 $Y=1.72
+ $X2=14.04 $Y2=1.805
r97 30 41 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=14.12 $Y=1.72
+ $X2=14.12 $Y2=0.96
r98 25 27 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=14.04 $Y=1.985
+ $X2=14.04 $Y2=2.815
r99 23 37 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=14.04 $Y=1.89
+ $X2=14.04 $Y2=1.805
r100 23 25 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=14.04 $Y=1.89
+ $X2=14.04 $Y2=1.985
r101 22 35 4.53325 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=13.33 $Y=1.805
+ $X2=13.167 $Y2=1.805
r102 21 37 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.875 $Y=1.805
+ $X2=14.04 $Y2=1.805
r103 21 22 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=13.875 $Y=1.805
+ $X2=13.33 $Y2=1.805
r104 17 46 21.3668 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=13.225 $Y=1.47
+ $X2=13.225 $Y2=1.677
r105 17 19 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=13.225 $Y=1.47
+ $X2=13.225 $Y2=0.69
r106 14 44 17.0727 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=13.035 $Y=1.885
+ $X2=13.035 $Y2=1.677
r107 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=13.035 $Y=1.885
+ $X2=13.035 $Y2=2.46
r108 10 43 21.3668 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=12.795 $Y=1.47
+ $X2=12.795 $Y2=1.677
r109 10 12 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=12.795 $Y=1.47
+ $X2=12.795 $Y2=0.69
r110 7 43 37.747 $w=3.32e-07 $l=3.48827e-07 $layer=POLY_cond $X=12.535 $Y=1.885
+ $X2=12.795 $Y2=1.677
r111 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.535 $Y=1.885
+ $X2=12.535 $Y2=2.46
r112 2 27 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=13.895
+ $Y=1.84 $X2=14.04 $Y2=2.815
r113 2 25 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=13.895
+ $Y=1.84 $X2=14.04 $Y2=1.985
r114 1 39 182 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_NDIFF $count=1 $X=13.925
+ $Y=0.37 $X2=14.07 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%A_2199_74# 1 2 3 4 5 6 21 25 29 33 37 41 45
+ 49 54 57 58 59 60 61 63 65 67 69 73 75 78 79 84 87 92 93 98 101 110
c206 110 0 2.3931e-20 $X=16.215 $Y=1.465
c207 63 0 2.5462e-21 $X=13.145 $Y=2.145
c208 61 0 5.98463e-20 $X=12.493 $Y=0.437
c209 59 0 8.44579e-20 $X=12.31 $Y=2.23
r210 110 111 14.1765 $w=3.06e-07 $l=9e-08 $layer=POLY_cond $X=16.215 $Y=1.465
+ $X2=16.305 $Y2=1.465
r211 107 108 17.3268 $w=3.06e-07 $l=1.1e-07 $layer=POLY_cond $X=15.765 $Y=1.465
+ $X2=15.875 $Y2=1.465
r212 106 107 50.4052 $w=3.06e-07 $l=3.2e-07 $layer=POLY_cond $X=15.445 $Y=1.465
+ $X2=15.765 $Y2=1.465
r213 105 106 28.3529 $w=3.06e-07 $l=1.8e-07 $layer=POLY_cond $X=15.265 $Y=1.465
+ $X2=15.445 $Y2=1.465
r214 97 98 8.52431 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=12.51 $Y=0.437
+ $X2=12.675 $Y2=0.437
r215 92 93 8.68217 $w=3.63e-07 $l=1.7e-07 $layer=LI1_cond $X=11.985 $Y=0.51
+ $X2=12.155 $Y2=0.51
r216 90 91 6.59757 $w=4.18e-07 $l=2.2e-07 $layer=LI1_cond $X=11.265 $Y=0.81
+ $X2=11.265 $Y2=1.03
r217 87 90 3.56709 $w=4.18e-07 $l=1.3e-07 $layer=LI1_cond $X=11.265 $Y=0.68
+ $X2=11.265 $Y2=0.81
r218 85 110 14.1765 $w=3.06e-07 $l=9e-08 $layer=POLY_cond $X=16.125 $Y=1.465
+ $X2=16.215 $Y2=1.465
r219 85 108 39.3791 $w=3.06e-07 $l=2.5e-07 $layer=POLY_cond $X=16.125 $Y=1.465
+ $X2=15.875 $Y2=1.465
r220 84 85 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=16.125
+ $Y=1.465 $X2=16.125 $Y2=1.465
r221 82 105 25.2026 $w=3.06e-07 $l=1.6e-07 $layer=POLY_cond $X=15.105 $Y=1.465
+ $X2=15.265 $Y2=1.465
r222 82 103 14.1765 $w=3.06e-07 $l=9e-08 $layer=POLY_cond $X=15.105 $Y=1.465
+ $X2=15.015 $Y2=1.465
r223 81 84 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=15.105 $Y=1.465
+ $X2=16.125 $Y2=1.465
r224 81 82 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=15.105
+ $Y=1.465 $X2=15.105 $Y2=1.465
r225 79 81 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=14.545 $Y=1.465
+ $X2=15.105 $Y2=1.465
r226 78 79 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=14.46 $Y=1.3
+ $X2=14.545 $Y2=1.465
r227 77 78 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=14.46 $Y=0.425
+ $X2=14.46 $Y2=1.3
r228 76 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.675 $Y=0.34
+ $X2=13.51 $Y2=0.34
r229 75 77 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.375 $Y=0.34
+ $X2=14.46 $Y2=0.425
r230 75 76 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=14.375 $Y=0.34
+ $X2=13.675 $Y2=0.34
r231 71 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.51 $Y=0.425
+ $X2=13.51 $Y2=0.34
r232 71 73 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=13.51 $Y=0.425
+ $X2=13.51 $Y2=0.495
r233 67 100 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.31 $Y=2.23
+ $X2=13.31 $Y2=2.145
r234 67 69 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=13.31 $Y=2.23
+ $X2=13.31 $Y2=2.485
r235 65 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.345 $Y=0.34
+ $X2=13.51 $Y2=0.34
r236 65 98 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=13.345 $Y=0.34
+ $X2=12.675 $Y2=0.34
r237 64 95 4.746 $w=1.7e-07 $l=1.90526e-07 $layer=LI1_cond $X=12.475 $Y=2.145
+ $X2=12.31 $Y2=2.09
r238 63 100 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.145 $Y=2.145
+ $X2=13.31 $Y2=2.145
r239 63 64 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=13.145 $Y=2.145
+ $X2=12.475 $Y2=2.145
r240 61 97 0.536754 $w=3.63e-07 $l=1.7e-08 $layer=LI1_cond $X=12.493 $Y=0.437
+ $X2=12.51 $Y2=0.437
r241 61 93 10.6719 $w=3.63e-07 $l=3.38e-07 $layer=LI1_cond $X=12.493 $Y=0.437
+ $X2=12.155 $Y2=0.437
r242 59 95 3.02018 $w=3.3e-07 $l=1.4e-07 $layer=LI1_cond $X=12.31 $Y=2.23
+ $X2=12.31 $Y2=2.09
r243 59 60 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=12.31 $Y=2.23
+ $X2=12.31 $Y2=2.565
r244 57 60 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.145 $Y=2.65
+ $X2=12.31 $Y2=2.565
r245 57 58 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=12.145 $Y=2.65
+ $X2=11.475 $Y2=2.65
r246 56 87 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=11.475 $Y=0.68
+ $X2=11.265 $Y2=0.68
r247 56 92 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=11.475 $Y=0.68
+ $X2=11.985 $Y2=0.68
r248 54 91 37.5417 $w=3.28e-07 $l=1.075e-06 $layer=LI1_cond $X=11.31 $Y=2.105
+ $X2=11.31 $Y2=1.03
r249 52 58 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.31 $Y=2.565
+ $X2=11.475 $Y2=2.65
r250 52 54 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=11.31 $Y=2.565
+ $X2=11.31 $Y2=2.105
r251 47 111 19.4347 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=16.305 $Y=1.3
+ $X2=16.305 $Y2=1.465
r252 47 49 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=16.305 $Y=1.3
+ $X2=16.305 $Y2=0.74
r253 43 110 15.178 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=16.215 $Y=1.63
+ $X2=16.215 $Y2=1.465
r254 43 45 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=16.215 $Y=1.63
+ $X2=16.215 $Y2=2.4
r255 39 108 19.4347 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.875 $Y=1.3
+ $X2=15.875 $Y2=1.465
r256 39 41 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=15.875 $Y=1.3
+ $X2=15.875 $Y2=0.74
r257 35 107 15.178 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=15.765 $Y=1.63
+ $X2=15.765 $Y2=1.465
r258 35 37 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=15.765 $Y=1.63
+ $X2=15.765 $Y2=2.4
r259 31 106 19.4347 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.445 $Y=1.3
+ $X2=15.445 $Y2=1.465
r260 31 33 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=15.445 $Y=1.3
+ $X2=15.445 $Y2=0.74
r261 27 105 15.178 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=15.265 $Y=1.63
+ $X2=15.265 $Y2=1.465
r262 27 29 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=15.265 $Y=1.63
+ $X2=15.265 $Y2=2.4
r263 23 103 19.4347 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.015 $Y=1.3
+ $X2=15.015 $Y2=1.465
r264 23 25 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=15.015 $Y=1.3
+ $X2=15.015 $Y2=0.74
r265 19 103 31.5033 $w=3.06e-07 $l=2.70185e-07 $layer=POLY_cond $X=14.815
+ $Y=1.63 $X2=15.015 $Y2=1.465
r266 19 21 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=14.815 $Y=1.63
+ $X2=14.815 $Y2=2.4
r267 6 100 600 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_PDIFF $count=1 $X=13.125
+ $Y=1.96 $X2=13.31 $Y2=2.145
r268 6 69 300 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_PDIFF $count=2 $X=13.125
+ $Y=1.96 $X2=13.31 $Y2=2.485
r269 5 95 300 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_PDIFF $count=2 $X=12.125
+ $Y=1.96 $X2=12.31 $Y2=2.115
r270 4 54 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=11.165
+ $Y=1.96 $X2=11.31 $Y2=2.105
r271 3 73 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=13.3
+ $Y=0.37 $X2=13.44 $Y2=0.495
r272 2 97 91 $w=1.7e-07 $l=5.64358e-07 $layer=licon1_NDIFF $count=2 $X=12.02
+ $Y=0.37 $X2=12.51 $Y2=0.53
r273 1 90 182 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_NDIFF $count=1 $X=10.995
+ $Y=0.37 $X2=11.14 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%VPWR 1 2 3 4 5 6 7 8 9 10 31 33 39 43 47 53
+ 57 63 65 67 70 73 77 78 80 81 83 84 85 87 92 97 105 126 134 137 140 143 151
r180 150 151 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.56 $Y=3.33
+ $X2=16.56 $Y2=3.33
r181 143 146 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=8.485 $Y=3.05
+ $X2=8.485 $Y2=3.33
r182 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r183 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r184 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r185 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r186 129 151 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.08 $Y=3.33
+ $X2=16.56 $Y2=3.33
r187 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.08 $Y=3.33
+ $X2=16.08 $Y2=3.33
r188 126 150 4.67153 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=16.325 $Y=3.33
+ $X2=16.562 $Y2=3.33
r189 126 128 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=16.325 $Y=3.33
+ $X2=16.08 $Y2=3.33
r190 125 129 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.12 $Y=3.33
+ $X2=16.08 $Y2=3.33
r191 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r192 122 125 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=15.12 $Y2=3.33
r193 121 122 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r194 119 122 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=14.16 $Y2=3.33
r195 118 121 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=10.8 $Y=3.33
+ $X2=14.16 $Y2=3.33
r196 118 119 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r197 116 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r198 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r199 113 116 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r200 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r201 110 146 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.65 $Y=3.33
+ $X2=8.485 $Y2=3.33
r202 110 112 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=8.65 $Y=3.33
+ $X2=9.36 $Y2=3.33
r203 109 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r204 108 109 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r205 106 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.73 $Y=3.33
+ $X2=5.565 $Y2=3.33
r206 106 108 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.73 $Y=3.33 $X2=6
+ $Y2=3.33
r207 105 146 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.32 $Y=3.33
+ $X2=8.485 $Y2=3.33
r208 105 108 151.358 $w=1.68e-07 $l=2.32e-06 $layer=LI1_cond $X=8.32 $Y=3.33
+ $X2=6 $Y2=3.33
r209 104 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r210 103 104 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r211 101 104 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=5.04 $Y2=3.33
r212 101 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r213 100 103 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=5.04 $Y2=3.33
r214 100 101 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r215 98 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.17 $Y2=3.33
r216 98 100 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.64 $Y2=3.33
r217 97 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.4 $Y=3.33
+ $X2=5.565 $Y2=3.33
r218 97 103 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=5.4 $Y=3.33
+ $X2=5.04 $Y2=3.33
r219 96 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r220 96 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r221 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r222 93 134 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.22 $Y2=3.33
r223 93 95 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=3.33
+ $X2=1.68 $Y2=3.33
r224 92 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.045 $Y=3.33
+ $X2=2.17 $Y2=3.33
r225 92 95 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.045 $Y=3.33
+ $X2=1.68 $Y2=3.33
r226 91 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r227 91 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r228 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r229 88 131 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r230 88 90 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r231 87 134 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.22 $Y2=3.33
r232 87 90 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.72 $Y2=3.33
r233 85 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r234 85 109 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.4 $Y=3.33 $X2=6
+ $Y2=3.33
r235 85 146 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r236 83 124 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=15.405 $Y=3.33
+ $X2=15.12 $Y2=3.33
r237 83 84 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.405 $Y=3.33
+ $X2=15.53 $Y2=3.33
r238 82 128 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=15.655 $Y=3.33
+ $X2=16.08 $Y2=3.33
r239 82 84 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.655 $Y=3.33
+ $X2=15.53 $Y2=3.33
r240 80 121 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=14.375 $Y=3.33
+ $X2=14.16 $Y2=3.33
r241 80 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.375 $Y=3.33
+ $X2=14.54 $Y2=3.33
r242 79 124 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=14.705 $Y=3.33
+ $X2=15.12 $Y2=3.33
r243 79 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.705 $Y=3.33
+ $X2=14.54 $Y2=3.33
r244 77 115 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=10.465 $Y=3.33
+ $X2=10.32 $Y2=3.33
r245 77 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.465 $Y=3.33
+ $X2=10.55 $Y2=3.33
r246 76 118 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.635 $Y=3.33
+ $X2=10.8 $Y2=3.33
r247 76 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.635 $Y=3.33
+ $X2=10.55 $Y2=3.33
r248 74 115 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=9.73 $Y=3.33
+ $X2=10.32 $Y2=3.33
r249 73 112 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=9.39 $Y=3.33
+ $X2=9.36 $Y2=3.33
r250 72 74 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=9.56 $Y=3.33
+ $X2=9.73 $Y2=3.33
r251 72 73 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=9.56 $Y=3.33
+ $X2=9.39 $Y2=3.33
r252 70 72 9.49071 $w=3.38e-07 $l=2.8e-07 $layer=LI1_cond $X=9.56 $Y=3.05
+ $X2=9.56 $Y2=3.33
r253 65 150 3.09464 $w=3.3e-07 $l=1.15521e-07 $layer=LI1_cond $X=16.49 $Y=3.245
+ $X2=16.562 $Y2=3.33
r254 65 67 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=16.49 $Y=3.245
+ $X2=16.49 $Y2=2.305
r255 61 84 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=15.53 $Y=3.245
+ $X2=15.53 $Y2=3.33
r256 61 63 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=15.53 $Y=3.245
+ $X2=15.53 $Y2=2.305
r257 57 60 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=14.54 $Y=1.985
+ $X2=14.54 $Y2=2.815
r258 55 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.54 $Y=3.245
+ $X2=14.54 $Y2=3.33
r259 55 60 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=14.54 $Y=3.245
+ $X2=14.54 $Y2=2.815
r260 51 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.55 $Y=3.245
+ $X2=10.55 $Y2=3.33
r261 51 53 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=10.55 $Y=3.245
+ $X2=10.55 $Y2=2.45
r262 47 50 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=5.565 $Y=1.985
+ $X2=5.565 $Y2=2.815
r263 45 140 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=3.245
+ $X2=5.565 $Y2=3.33
r264 45 50 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.565 $Y=3.245
+ $X2=5.565 $Y2=2.815
r265 41 137 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=3.33
r266 41 43 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=2.815
r267 37 134 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=3.245
+ $X2=1.22 $Y2=3.33
r268 37 39 35.4952 $w=2.48e-07 $l=7.7e-07 $layer=LI1_cond $X=1.22 $Y=3.245
+ $X2=1.22 $Y2=2.475
r269 33 36 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=0.24 $Y=2.115
+ $X2=0.24 $Y2=2.815
r270 31 131 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r271 31 36 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.815
r272 10 67 300 $w=1.7e-07 $l=5.49773e-07 $layer=licon1_PDIFF $count=2 $X=16.305
+ $Y=1.84 $X2=16.49 $Y2=2.305
r273 9 63 300 $w=1.7e-07 $l=5.28205e-07 $layer=licon1_PDIFF $count=2 $X=15.355
+ $Y=1.84 $X2=15.49 $Y2=2.305
r274 8 60 400 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=14.39
+ $Y=1.84 $X2=14.54 $Y2=2.815
r275 8 57 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=14.39
+ $Y=1.84 $X2=14.54 $Y2=1.985
r276 7 53 300 $w=1.7e-07 $l=5.53399e-07 $layer=licon1_PDIFF $count=2 $X=10.415
+ $Y=1.96 $X2=10.55 $Y2=2.45
r277 6 70 600 $w=1.7e-07 $l=1.19723e-06 $layer=licon1_PDIFF $count=1 $X=9.335
+ $Y=1.96 $X2=9.56 $Y2=3.05
r278 5 143 600 $w=1.7e-07 $l=1.16024e-06 $layer=licon1_PDIFF $count=1 $X=8.34
+ $Y=1.96 $X2=8.485 $Y2=3.05
r279 4 50 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=5.43
+ $Y=1.84 $X2=5.565 $Y2=2.815
r280 4 47 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.43
+ $Y=1.84 $X2=5.565 $Y2=1.985
r281 3 43 600 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.96 $X2=2.13 $Y2=2.815
r282 2 39 300 $w=1.7e-07 $l=5.78576e-07 $layer=licon1_PDIFF $count=2 $X=1.045
+ $Y=1.96 $X2=1.18 $Y2=2.475
r283 1 36 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.815
r284 1 33 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.96 $X2=0.28 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%A_119_392# 1 2 7 9 11 14 15 16 19
c63 16 0 6.40679e-20 $X=2.695 $Y=1.685
c64 14 0 2.7261e-19 $X=2.61 $Y=1.97
c65 7 0 2.19288e-19 $X=0.73 $Y=2.14
r66 17 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.105 $Y=1.77
+ $X2=4.105 $Y2=2.105
r67 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.02 $Y=1.685
+ $X2=4.105 $Y2=1.77
r68 15 16 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=4.02 $Y=1.685
+ $X2=2.695 $Y2=1.685
r69 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.61 $Y=1.77
+ $X2=2.695 $Y2=1.685
r70 13 14 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.61 $Y=1.77 $X2=2.61
+ $Y2=1.97
r71 12 22 5.03363 $w=1.7e-07 $l=1.69926e-07 $layer=LI1_cond $X=0.895 $Y=2.055
+ $X2=0.73 $Y2=2.045
r72 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.525 $Y=2.055
+ $X2=2.61 $Y2=1.97
r73 11 12 106.342 $w=1.68e-07 $l=1.63e-06 $layer=LI1_cond $X=2.525 $Y=2.055
+ $X2=0.895 $Y2=2.055
r74 7 22 2.73254 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=0.73 $Y=2.14 $X2=0.73
+ $Y2=2.045
r75 7 9 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.73 $Y=2.14 $X2=0.73
+ $Y2=2.815
r76 2 19 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.97
+ $Y=1.96 $X2=4.105 $Y2=2.105
r77 1 22 400 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.96 $X2=0.73 $Y2=2.115
r78 1 9 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.96 $X2=0.73 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%A_299_392# 1 2 9 13 16 17
c29 16 0 1.72297e-19 $X=1.68 $Y=2.475
r30 17 19 7.70758 $w=2.77e-07 $l=1.75e-07 $layer=LI1_cond $X=3.145 $Y=2.395
+ $X2=3.145 $Y2=2.57
r31 11 17 3.51151 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.145 $Y=2.31
+ $X2=3.145 $Y2=2.395
r32 11 13 7.62099 $w=3.08e-07 $l=2.05e-07 $layer=LI1_cond $X=3.145 $Y=2.31
+ $X2=3.145 $Y2=2.105
r33 10 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=2.395
+ $X2=1.68 $Y2=2.395
r34 9 17 3.59349 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=2.99 $Y=2.395
+ $X2=3.145 $Y2=2.395
r35 9 10 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=2.99 $Y=2.395
+ $X2=1.845 $Y2=2.395
r36 2 19 600 $w=1.7e-07 $l=6.74129e-07 $layer=licon1_PDIFF $count=1 $X=3.02
+ $Y=1.96 $X2=3.155 $Y2=2.57
r37 2 13 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.02
+ $Y=1.96 $X2=3.155 $Y2=2.105
r38 1 16 300 $w=1.7e-07 $l=6.00417e-07 $layer=licon1_PDIFF $count=2 $X=1.495
+ $Y=1.96 $X2=1.68 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%A_509_392# 1 2 3 4 5 6 7 8 25 27 31 37 39 41
+ 46 52 55 56 57 60 64 69 70 71 73 78 82 83 86 89 90 97
c187 90 0 1.46885e-19 $X=11.76 $Y=2.035
c188 73 0 4.75356e-20 $X=12.41 $Y=0.875
c189 5 0 1.67617e-19 $X=2.545 $Y=1.96
r190 90 94 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=11.81 $Y=2.035
+ $X2=11.81 $Y2=2.23
r191 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=2.035
+ $X2=11.76 $Y2=2.035
r192 86 97 6.8092 $w=3.43e-07 $l=1.15e-07 $layer=LI1_cond $X=4.547 $Y=2.035
+ $X2=4.547 $Y2=1.92
r193 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=2.035
+ $X2=4.56 $Y2=2.035
r194 83 85 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.705 $Y=2.035
+ $X2=4.56 $Y2=2.035
r195 82 89 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.615 $Y=2.035
+ $X2=11.76 $Y2=2.035
r196 82 83 8.55196 $w=1.4e-07 $l=6.91e-06 $layer=MET1_cond $X=11.615 $Y=2.035
+ $X2=4.705 $Y2=2.035
r197 73 75 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=12.41 $Y=0.875
+ $X2=12.41 $Y2=1.02
r198 72 90 32.4779 $w=3.28e-07 $l=9.3e-07 $layer=LI1_cond $X=11.81 $Y=1.105
+ $X2=11.81 $Y2=2.035
r199 71 97 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=4.46 $Y=1.18
+ $X2=4.46 $Y2=1.92
r200 64 67 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.705 $Y=0.34
+ $X2=2.705 $Y2=0.455
r201 60 62 6.02022 $w=3.33e-07 $l=1.75e-07 $layer=LI1_cond $X=2.692 $Y=2.815
+ $X2=2.692 $Y2=2.99
r202 58 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.495 $Y=0.875
+ $X2=12.41 $Y2=0.875
r203 57 78 3.65855 $w=3.13e-07 $l=1e-07 $layer=LI1_cond $X=13.017 $Y=0.875
+ $X2=13.017 $Y2=0.775
r204 57 58 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=12.86 $Y=0.875
+ $X2=12.495 $Y2=0.875
r205 56 72 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.975 $Y=1.02
+ $X2=11.81 $Y2=1.105
r206 55 75 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.325 $Y=1.02
+ $X2=12.41 $Y2=1.02
r207 55 56 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=12.325 $Y=1.02
+ $X2=11.975 $Y2=1.02
r208 52 54 23.7169 $w=3.43e-07 $l=7.1e-07 $layer=LI1_cond $X=4.547 $Y=2.105
+ $X2=4.547 $Y2=2.815
r209 50 54 3.00637 $w=3.43e-07 $l=9e-08 $layer=LI1_cond $X=4.547 $Y=2.905
+ $X2=4.547 $Y2=2.815
r210 49 86 1.90404 $w=3.43e-07 $l=5.7e-08 $layer=LI1_cond $X=4.547 $Y=2.092
+ $X2=4.547 $Y2=2.035
r211 49 52 0.434254 $w=3.43e-07 $l=1.3e-08 $layer=LI1_cond $X=4.547 $Y=2.092
+ $X2=4.547 $Y2=2.105
r212 44 71 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=4.545 $Y=1.01
+ $X2=4.545 $Y2=1.18
r213 44 46 8.64332 $w=3.38e-07 $l=2.55e-07 $layer=LI1_cond $X=4.545 $Y=1.01
+ $X2=4.545 $Y2=0.755
r214 43 46 11.1855 $w=3.38e-07 $l=3.3e-07 $layer=LI1_cond $X=4.545 $Y=0.425
+ $X2=4.545 $Y2=0.755
r215 42 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.82 $Y=2.99
+ $X2=3.655 $Y2=2.99
r216 41 50 7.89393 $w=1.7e-07 $l=2.10247e-07 $layer=LI1_cond $X=4.375 $Y=2.99
+ $X2=4.547 $Y2=2.905
r217 41 42 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=4.375 $Y=2.99
+ $X2=3.82 $Y2=2.99
r218 40 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.775 $Y=0.34
+ $X2=3.69 $Y2=0.34
r219 39 43 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=4.375 $Y=0.34
+ $X2=4.545 $Y2=0.425
r220 39 40 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.375 $Y=0.34
+ $X2=3.775 $Y2=0.34
r221 35 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=0.425
+ $X2=3.69 $Y2=0.34
r222 35 37 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.69 $Y=0.425
+ $X2=3.69 $Y2=0.87
r223 31 34 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.655 $Y=2.105
+ $X2=3.655 $Y2=2.815
r224 29 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.655 $Y=2.905
+ $X2=3.655 $Y2=2.99
r225 29 34 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.655 $Y=2.905
+ $X2=3.655 $Y2=2.815
r226 28 64 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.87 $Y=0.34
+ $X2=2.705 $Y2=0.34
r227 27 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.605 $Y=0.34
+ $X2=3.69 $Y2=0.34
r228 27 28 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=3.605 $Y=0.34
+ $X2=2.87 $Y2=0.34
r229 26 62 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.86 $Y=2.99
+ $X2=2.692 $Y2=2.99
r230 25 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.49 $Y=2.99
+ $X2=3.655 $Y2=2.99
r231 25 26 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.49 $Y=2.99
+ $X2=2.86 $Y2=2.99
r232 8 94 600 $w=1.7e-07 $l=3.505e-07 $layer=licon1_PDIFF $count=1 $X=11.625
+ $Y=1.96 $X2=11.81 $Y2=2.23
r233 7 54 400 $w=1.7e-07 $l=9.20027e-07 $layer=licon1_PDIFF $count=1 $X=4.42
+ $Y=1.96 $X2=4.555 $Y2=2.815
r234 7 52 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.42
+ $Y=1.96 $X2=4.555 $Y2=2.105
r235 6 34 400 $w=1.7e-07 $l=9.31571e-07 $layer=licon1_PDIFF $count=1 $X=3.495
+ $Y=1.96 $X2=3.655 $Y2=2.815
r236 6 31 400 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=3.495
+ $Y=1.96 $X2=3.655 $Y2=2.105
r237 5 60 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.545
+ $Y=1.96 $X2=2.695 $Y2=2.815
r238 4 78 182 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_NDIFF $count=1 $X=12.87
+ $Y=0.37 $X2=13.01 $Y2=0.775
r239 3 46 91 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=2 $X=4.41
+ $Y=0.595 $X2=4.55 $Y2=0.755
r240 2 37 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.55
+ $Y=0.595 $X2=3.69 $Y2=0.87
r241 1 67 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=2.56
+ $Y=0.31 $X2=2.705 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%A_1191_121# 1 2 3 4 5 6 7 8 25 27 29 31 33 35
+ 37 38 40 43 45 47 52 54 55 57 59 60 63 71 73 74 79
c172 71 0 7.97039e-20 $X=7 $Y=1.145
c173 45 0 1.54503e-19 $X=7.735 $Y=0.68
c174 37 0 7.8786e-20 $X=7 $Y=0.765
r175 74 77 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=7.86 $Y=0.68 $X2=7.86
+ $Y2=0.76
r176 61 63 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=12.81 $Y=2.905
+ $X2=12.81 $Y2=2.485
r177 59 61 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.645 $Y=2.99
+ $X2=12.81 $Y2=2.905
r178 59 60 108.952 $w=1.68e-07 $l=1.67e-06 $layer=LI1_cond $X=12.645 $Y=2.99
+ $X2=10.975 $Y2=2.99
r179 55 57 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=10.885 $Y=0.34
+ $X2=11.65 $Y2=0.34
r180 54 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.89 $Y=2.905
+ $X2=10.975 $Y2=2.99
r181 53 79 5.16603 $w=1.7e-07 $l=1.05119e-07 $layer=LI1_cond $X=10.89 $Y=2.115
+ $X2=10.845 $Y2=2.03
r182 53 54 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=10.89 $Y=2.115
+ $X2=10.89 $Y2=2.905
r183 52 79 5.16603 $w=1.7e-07 $l=1.05119e-07 $layer=LI1_cond $X=10.8 $Y=1.945
+ $X2=10.845 $Y2=2.03
r184 51 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.8 $Y=0.425
+ $X2=10.885 $Y2=0.34
r185 51 52 99.1658 $w=1.68e-07 $l=1.52e-06 $layer=LI1_cond $X=10.8 $Y=0.425
+ $X2=10.8 $Y2=1.945
r186 48 73 3.31178 $w=1.7e-07 $l=1.11216e-07 $layer=LI1_cond $X=7.125 $Y=2.03
+ $X2=7.032 $Y2=1.99
r187 48 50 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=7.125 $Y=2.03
+ $X2=7.925 $Y2=2.03
r188 47 79 1.34256 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.715 $Y=2.03
+ $X2=10.845 $Y2=2.03
r189 47 50 182.021 $w=1.68e-07 $l=2.79e-06 $layer=LI1_cond $X=10.715 $Y=2.03
+ $X2=7.925 $Y2=2.03
r190 46 70 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.125 $Y=0.68 $X2=7
+ $Y2=0.68
r191 45 74 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.735 $Y=0.68
+ $X2=7.86 $Y2=0.68
r192 45 46 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.735 $Y=0.68
+ $X2=7.125 $Y2=0.68
r193 41 73 2.79615 $w=1.85e-07 $l=1.25e-07 $layer=LI1_cond $X=7.032 $Y=2.115
+ $X2=7.032 $Y2=1.99
r194 41 43 27.2776 $w=1.83e-07 $l=4.55e-07 $layer=LI1_cond $X=7.032 $Y=2.115
+ $X2=7.032 $Y2=2.57
r195 40 73 2.79615 $w=1.85e-07 $l=1.25e-07 $layer=LI1_cond $X=7.032 $Y=1.865
+ $X2=7.032 $Y2=1.99
r196 39 71 4.18896 $w=2.17e-07 $l=1.35056e-07 $layer=LI1_cond $X=7.032 $Y=1.265
+ $X2=7 $Y2=1.145
r197 39 40 35.9705 $w=1.83e-07 $l=6e-07 $layer=LI1_cond $X=7.032 $Y=1.265
+ $X2=7.032 $Y2=1.865
r198 38 71 4.18896 $w=2.17e-07 $l=1.2e-07 $layer=LI1_cond $X=7 $Y=1.025 $X2=7
+ $Y2=1.145
r199 37 70 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7 $Y=0.765 $X2=7
+ $Y2=0.68
r200 37 38 11.9854 $w=2.48e-07 $l=2.6e-07 $layer=LI1_cond $X=7 $Y=0.765 $X2=7
+ $Y2=1.025
r201 36 68 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.21 $Y=1.95
+ $X2=6.085 $Y2=1.95
r202 35 73 3.31178 $w=1.7e-07 $l=1.102e-07 $layer=LI1_cond $X=6.94 $Y=1.95
+ $X2=7.032 $Y2=1.99
r203 35 36 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.94 $Y=1.95
+ $X2=6.21 $Y2=1.95
r204 34 66 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.185 $Y=1.11
+ $X2=6.06 $Y2=1.11
r205 33 71 2.24312 $w=1.7e-07 $l=1.41421e-07 $layer=LI1_cond $X=6.875 $Y=1.11
+ $X2=7 $Y2=1.145
r206 33 34 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.875 $Y=1.11
+ $X2=6.185 $Y2=1.11
r207 29 68 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.085 $Y=2.035
+ $X2=6.085 $Y2=1.95
r208 29 31 32.4989 $w=2.48e-07 $l=7.05e-07 $layer=LI1_cond $X=6.085 $Y=2.035
+ $X2=6.085 $Y2=2.74
r209 25 66 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.06 $Y=1.025
+ $X2=6.06 $Y2=1.11
r210 25 27 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=6.06 $Y=1.025
+ $X2=6.06 $Y2=0.75
r211 8 63 300 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_PDIFF $count=2 $X=12.625
+ $Y=1.96 $X2=12.81 $Y2=2.485
r212 7 50 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.79
+ $Y=1.885 $X2=7.925 $Y2=2.03
r213 6 73 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.89
+ $Y=1.885 $X2=7.025 $Y2=2.03
r214 6 43 600 $w=1.7e-07 $l=7.49466e-07 $layer=licon1_PDIFF $count=1 $X=6.89
+ $Y=1.885 $X2=7.025 $Y2=2.57
r215 5 68 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.98
+ $Y=1.885 $X2=6.125 $Y2=2.03
r216 5 31 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.98
+ $Y=1.885 $X2=6.125 $Y2=2.74
r217 4 57 182 $w=1.7e-07 $l=2.34521e-07 $layer=licon1_NDIFF $count=1 $X=11.43
+ $Y=0.37 $X2=11.65 $Y2=0.34
r218 3 77 182 $w=1.7e-07 $l=2.87228e-07 $layer=licon1_NDIFF $count=1 $X=7.68
+ $Y=0.605 $X2=7.9 $Y2=0.76
r219 2 70 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=6.82
+ $Y=0.605 $X2=6.96 $Y2=0.76
r220 1 66 182 $w=1.7e-07 $l=5.72931e-07 $layer=licon1_NDIFF $count=1 $X=5.955
+ $Y=0.605 $X2=6.1 $Y2=1.11
r221 1 27 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=5.955
+ $Y=0.605 $X2=6.1 $Y2=0.75
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%A_1288_377# 1 2 9 11 12 13 17 19
r55 19 21 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=8.065 $Y=2.71
+ $X2=8.065 $Y2=2.99
r56 15 17 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=10.1 $Y=2.625
+ $X2=10.1 $Y2=2.45
r57 14 19 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.15 $Y=2.71
+ $X2=8.065 $Y2=2.71
r58 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.935 $Y=2.71
+ $X2=10.1 $Y2=2.625
r59 13 14 116.455 $w=1.68e-07 $l=1.785e-06 $layer=LI1_cond $X=9.935 $Y=2.71
+ $X2=8.15 $Y2=2.71
r60 11 21 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.98 $Y=2.99
+ $X2=8.065 $Y2=2.99
r61 11 12 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=7.98 $Y=2.99
+ $X2=6.74 $Y2=2.99
r62 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.575 $Y=2.905
+ $X2=6.74 $Y2=2.99
r63 7 9 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=6.575 $Y=2.905
+ $X2=6.575 $Y2=2.315
r64 2 17 300 $w=1.7e-07 $l=5.53399e-07 $layer=licon1_PDIFF $count=2 $X=9.965
+ $Y=1.96 $X2=10.1 $Y2=2.45
r65 1 9 300 $w=1.7e-07 $l=4.929e-07 $layer=licon1_PDIFF $count=2 $X=6.44
+ $Y=1.885 $X2=6.575 $Y2=2.315
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%A_1468_377# 1 2 9 11
c21 9 0 4.1337e-20 $X=9.02 $Y=2.37
r22 11 14 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=7.475 $Y=2.37
+ $X2=7.475 $Y2=2.55
r23 7 11 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.64 $Y=2.37
+ $X2=7.475 $Y2=2.37
r24 7 9 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=7.64 $Y=2.37 $X2=9.02
+ $Y2=2.37
r25 2 9 600 $w=1.7e-07 $l=4.72705e-07 $layer=licon1_PDIFF $count=1 $X=8.885
+ $Y=1.96 $X2=9.02 $Y2=2.37
r26 1 14 600 $w=1.7e-07 $l=7.29383e-07 $layer=licon1_PDIFF $count=1 $X=7.34
+ $Y=1.885 $X2=7.475 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%X 1 2 3 4 15 21 23 24 25 26 29 35 37 39 41 42
+ 45 46
c83 24 0 1.03922e-19 $X=15.205 $Y=1.885
r84 45 46 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=16.56 $Y=1.295
+ $X2=16.56 $Y2=1.665
r85 44 46 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=16.56 $Y=1.8
+ $X2=16.56 $Y2=1.665
r86 43 45 8.26753 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=16.56 $Y=1.13
+ $X2=16.56 $Y2=1.295
r87 40 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.175 $Y=1.045
+ $X2=16.05 $Y2=1.045
r88 39 43 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=16.445 $Y=1.045
+ $X2=16.56 $Y2=1.13
r89 39 40 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=16.445 $Y=1.045
+ $X2=16.175 $Y2=1.045
r90 38 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.155 $Y=1.885
+ $X2=15.99 $Y2=1.885
r91 37 44 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=16.445 $Y=1.885
+ $X2=16.56 $Y2=1.8
r92 37 38 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=16.445 $Y=1.885
+ $X2=16.155 $Y2=1.885
r93 33 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=16.05 $Y=0.96
+ $X2=16.05 $Y2=1.045
r94 33 35 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=16.05 $Y=0.96
+ $X2=16.05 $Y2=0.515
r95 29 31 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=15.99 $Y=1.985
+ $X2=15.99 $Y2=2.815
r96 27 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.99 $Y=1.97
+ $X2=15.99 $Y2=1.885
r97 27 29 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=15.99 $Y=1.97
+ $X2=15.99 $Y2=1.985
r98 25 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.925 $Y=1.045
+ $X2=16.05 $Y2=1.045
r99 25 26 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=15.925 $Y=1.045
+ $X2=15.315 $Y2=1.045
r100 23 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.825 $Y=1.885
+ $X2=15.99 $Y2=1.885
r101 23 24 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=15.825 $Y=1.885
+ $X2=15.205 $Y2=1.885
r102 19 26 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=15.19 $Y=0.96
+ $X2=15.315 $Y2=1.045
r103 19 21 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=15.19 $Y=0.96
+ $X2=15.19 $Y2=0.515
r104 15 17 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=15.04 $Y=1.985
+ $X2=15.04 $Y2=2.815
r105 13 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=15.04 $Y=1.97
+ $X2=15.205 $Y2=1.885
r106 13 15 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=15.04 $Y=1.97
+ $X2=15.04 $Y2=1.985
r107 4 31 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=15.855
+ $Y=1.84 $X2=15.99 $Y2=2.815
r108 4 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=15.855
+ $Y=1.84 $X2=15.99 $Y2=1.985
r109 3 17 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=14.905
+ $Y=1.84 $X2=15.04 $Y2=2.815
r110 3 15 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=14.905
+ $Y=1.84 $X2=15.04 $Y2=1.985
r111 2 35 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=15.95
+ $Y=0.37 $X2=16.09 $Y2=0.515
r112 1 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=15.09
+ $Y=0.37 $X2=15.23 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%VGND 1 2 3 4 5 6 7 8 9 10 31 32 34 35 37 39
+ 43 47 51 53 57 61 65 67 69 75 76 82 83 85 86 87 89 97 122 126 135 138 141 144
+ 148
c202 57 0 2.68867e-20 $X=10.46 $Y=0.515
c203 37 0 7.75212e-20 $X=1.207 $Y=1.03
c204 35 0 1.23921e-19 $X=1.045 $Y=1.155
r205 147 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.56 $Y=0
+ $X2=16.56 $Y2=0
r206 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=0
+ $X2=15.6 $Y2=0
r207 141 142 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r208 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r209 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r210 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r211 130 148 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.08 $Y=0
+ $X2=16.56 $Y2=0
r212 130 145 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.08 $Y=0
+ $X2=15.6 $Y2=0
r213 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.08 $Y=0
+ $X2=16.08 $Y2=0
r214 127 144 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.745 $Y=0
+ $X2=15.62 $Y2=0
r215 127 129 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=15.745 $Y=0
+ $X2=16.08 $Y2=0
r216 126 147 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=16.355 $Y=0
+ $X2=16.577 $Y2=0
r217 126 129 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=16.355 $Y=0
+ $X2=16.08 $Y2=0
r218 125 145 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=0
+ $X2=15.6 $Y2=0
r219 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r220 122 144 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.495 $Y=0
+ $X2=15.62 $Y2=0
r221 122 124 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=15.495 $Y=0
+ $X2=15.12 $Y2=0
r222 121 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=15.12 $Y2=0
r223 120 121 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r224 118 121 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=14.64 $Y2=0
r225 118 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=10.32 $Y2=0
r226 117 120 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=10.8 $Y=0
+ $X2=14.64 $Y2=0
r227 117 118 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r228 115 141 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.545 $Y=0
+ $X2=10.42 $Y2=0
r229 115 117 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=10.545 $Y=0
+ $X2=10.8 $Y2=0
r230 114 142 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=10.32 $Y2=0
r231 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r232 108 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r233 107 110 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=6 $Y=0 $X2=8.4
+ $Y2=0
r234 107 108 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=0 $X2=6
+ $Y2=0
r235 105 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.705 $Y=0
+ $X2=5.54 $Y2=0
r236 105 107 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.705 $Y=0 $X2=6
+ $Y2=0
r237 104 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r238 103 104 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r239 101 104 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=5.04 $Y2=0
r240 101 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=2.16 $Y2=0
r241 100 103 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.64 $Y=0
+ $X2=5.04 $Y2=0
r242 100 101 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r243 98 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.31 $Y=0
+ $X2=2.145 $Y2=0
r244 98 100 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.64
+ $Y2=0
r245 97 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.375 $Y=0
+ $X2=5.54 $Y2=0
r246 97 103 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.375 $Y=0
+ $X2=5.04 $Y2=0
r247 96 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r248 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r249 93 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r250 93 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r251 92 95 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r252 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r253 90 132 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r254 90 92 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.72 $Y2=0
r255 89 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.98 $Y=0
+ $X2=2.145 $Y2=0
r256 89 95 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.98 $Y=0 $X2=1.68
+ $Y2=0
r257 87 114 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r258 87 108 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.4 $Y=0 $X2=6
+ $Y2=0
r259 87 110 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r260 85 120 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=14.715 $Y=0
+ $X2=14.64 $Y2=0
r261 85 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.715 $Y=0 $X2=14.8
+ $Y2=0
r262 84 124 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=14.885 $Y=0
+ $X2=15.12 $Y2=0
r263 84 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.885 $Y=0 $X2=14.8
+ $Y2=0
r264 82 113 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=9.435 $Y=0
+ $X2=9.36 $Y2=0
r265 82 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.435 $Y=0 $X2=9.56
+ $Y2=0
r266 78 113 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=8.825 $Y=0
+ $X2=9.36 $Y2=0
r267 76 110 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=8.495 $Y=0 $X2=8.4
+ $Y2=0
r268 75 80 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=8.66 $Y=0 $X2=8.66
+ $Y2=0.325
r269 75 78 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.66 $Y=0 $X2=8.825
+ $Y2=0
r270 75 76 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.66 $Y=0 $X2=8.495
+ $Y2=0
r271 67 147 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=16.52 $Y=0.085
+ $X2=16.577 $Y2=0
r272 67 69 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=16.52 $Y=0.085
+ $X2=16.52 $Y2=0.625
r273 63 144 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=15.62 $Y=0.085
+ $X2=15.62 $Y2=0
r274 63 65 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=15.62 $Y=0.085
+ $X2=15.62 $Y2=0.625
r275 59 86 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.8 $Y=0.085
+ $X2=14.8 $Y2=0
r276 59 61 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=14.8 $Y=0.085
+ $X2=14.8 $Y2=0.515
r277 55 141 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.42 $Y=0.085
+ $X2=10.42 $Y2=0
r278 55 57 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.42 $Y=0.085
+ $X2=10.42 $Y2=0.515
r279 54 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.685 $Y=0 $X2=9.56
+ $Y2=0
r280 53 141 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.295 $Y=0
+ $X2=10.42 $Y2=0
r281 53 54 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=10.295 $Y=0
+ $X2=9.685 $Y2=0
r282 49 83 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.56 $Y=0.085
+ $X2=9.56 $Y2=0
r283 49 51 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=9.56 $Y=0.085
+ $X2=9.56 $Y2=0.55
r284 45 138 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.54 $Y=0.085
+ $X2=5.54 $Y2=0
r285 45 47 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=5.54 $Y=0.085
+ $X2=5.54 $Y2=0.515
r286 41 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=0.085
+ $X2=2.145 $Y2=0
r287 41 43 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=2.145 $Y=0.085
+ $X2=2.145 $Y2=0.365
r288 37 74 3.03503 $w=3.25e-07 $l=1.25e-07 $layer=LI1_cond $X=1.207 $Y=1.03
+ $X2=1.207 $Y2=1.155
r289 37 39 7.97845 $w=3.23e-07 $l=2.25e-07 $layer=LI1_cond $X=1.207 $Y=1.03
+ $X2=1.207 $Y2=0.805
r290 36 72 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=1.155
+ $X2=0.24 $Y2=1.155
r291 35 74 3.93339 $w=2.5e-07 $l=1.62e-07 $layer=LI1_cond $X=1.045 $Y=1.155
+ $X2=1.207 $Y2=1.155
r292 35 36 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=1.045 $Y=1.155
+ $X2=0.365 $Y2=1.155
r293 32 72 3.40825 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=1.03
+ $X2=0.24 $Y2=1.155
r294 32 34 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.24 $Y=1.03
+ $X2=0.24 $Y2=0.775
r295 31 132 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r296 31 34 31.8074 $w=2.48e-07 $l=6.9e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.775
r297 10 69 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=16.38
+ $Y=0.37 $X2=16.52 $Y2=0.625
r298 9 65 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=15.52
+ $Y=0.37 $X2=15.66 $Y2=0.625
r299 8 61 91 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_NDIFF $count=2 $X=14.36
+ $Y=0.37 $X2=14.8 $Y2=0.515
r300 7 57 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=10.32
+ $Y=0.37 $X2=10.46 $Y2=0.515
r301 6 51 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=9.46 $Y=0.37
+ $X2=9.6 $Y2=0.55
r302 5 80 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=8.515
+ $Y=0.18 $X2=8.66 $Y2=0.325
r303 4 47 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.4
+ $Y=0.37 $X2=5.54 $Y2=0.515
r304 3 43 182 $w=1.7e-07 $l=3.58504e-07 $layer=licon1_NDIFF $count=1 $X=1.925
+ $Y=0.63 $X2=2.145 $Y2=0.365
r305 2 74 182 $w=1.7e-07 $l=5.93949e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.63 $X2=1.17 $Y2=1.145
r306 2 39 182 $w=1.7e-07 $l=2.45713e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.63 $X2=1.17 $Y2=0.805
r307 1 72 182 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.63 $X2=0.28 $Y2=1.115
r308 1 34 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.63 $X2=0.28 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%A_114_126# 1 2 9 11 12 14 16 19 20
c50 20 0 6.40679e-20 $X=3.05 $Y=0.842
r51 19 20 9.48656 $w=4.93e-07 $l=1.65e-07 $layer=LI1_cond $X=3.215 $Y=0.842
+ $X2=3.05 $Y2=0.842
r52 16 17 25.4121 $w=2.21e-07 $l=4.88655e-07 $layer=LI1_cond $X=2.14 $Y=0.875
+ $X2=1.692 $Y2=0.79
r53 16 20 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=2.14 $Y=0.875
+ $X2=3.05 $Y2=0.875
r54 14 17 0.366029 $w=2.35e-07 $l=1.7e-07 $layer=LI1_cond $X=1.692 $Y=0.62
+ $X2=1.692 $Y2=0.79
r55 13 14 7.35602 $w=2.33e-07 $l=1.5e-07 $layer=LI1_cond $X=1.692 $Y=0.47
+ $X2=1.692 $Y2=0.62
r56 11 13 6.89349 $w=1.95e-07 $l=1.58603e-07 $layer=LI1_cond $X=1.575 $Y=0.372
+ $X2=1.692 $Y2=0.47
r57 11 12 39.8135 $w=1.93e-07 $l=7e-07 $layer=LI1_cond $X=1.575 $Y=0.372
+ $X2=0.875 $Y2=0.372
r58 7 12 7.4197 $w=1.95e-07 $l=2.08315e-07 $layer=LI1_cond $X=0.71 $Y=0.47
+ $X2=0.875 $Y2=0.372
r59 7 9 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.71 $Y=0.47 $X2=0.71
+ $Y2=0.775
r60 2 19 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=3.075
+ $Y=0.595 $X2=3.215 $Y2=0.84
r61 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.63 $X2=0.71 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%A_299_126# 1 2 7 9 13 16 20
c42 13 0 1.75061e-19 $X=4.12 $Y=0.76
r43 20 22 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.61 $Y=1.215
+ $X2=2.61 $Y2=1.345
r44 16 18 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.675 $Y=1.125
+ $X2=1.675 $Y2=1.215
r45 11 13 23.0489 $w=2.48e-07 $l=5e-07 $layer=LI1_cond $X=4.08 $Y=1.26 $X2=4.08
+ $Y2=0.76
r46 10 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=1.345
+ $X2=2.61 $Y2=1.345
r47 9 11 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.955 $Y=1.345
+ $X2=4.08 $Y2=1.26
r48 9 10 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=3.955 $Y=1.345
+ $X2=2.695 $Y2=1.345
r49 8 18 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.8 $Y=1.215
+ $X2=1.675 $Y2=1.215
r50 7 20 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=1.215
+ $X2=2.61 $Y2=1.215
r51 7 8 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=2.525 $Y=1.215
+ $X2=1.8 $Y2=1.215
r52 2 13 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=3.98
+ $Y=0.595 $X2=4.12 $Y2=0.76
r53 1 16 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.63 $X2=1.635 $Y2=1.125
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%A_1278_121# 1 2 9 11 12 14 15 16 18
c53 18 0 1.66006e-19 $X=9.17 $Y=0.55
c54 16 0 8.44834e-20 $X=8.325 $Y=0.665
r55 18 20 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=9.13 $Y=0.55
+ $X2=9.13 $Y2=0.665
r56 15 20 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.005 $Y=0.665
+ $X2=9.13 $Y2=0.665
r57 15 16 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.005 $Y=0.665
+ $X2=8.325 $Y2=0.665
r58 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.24 $Y=0.58
+ $X2=8.325 $Y2=0.665
r59 13 14 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=8.24 $Y=0.425
+ $X2=8.24 $Y2=0.58
r60 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.155 $Y=0.34
+ $X2=8.24 $Y2=0.425
r61 11 12 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=8.155 $Y=0.34
+ $X2=6.695 $Y2=0.34
r62 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.53 $Y=0.425
+ $X2=6.695 $Y2=0.34
r63 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.53 $Y=0.425 $X2=6.53
+ $Y2=0.76
r64 2 18 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=9.03 $Y=0.37
+ $X2=9.17 $Y2=0.55
r65 1 9 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=6.39
+ $Y=0.605 $X2=6.53 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__MUX4_4%A_1450_121# 1 2 7 9 13 16 20
c50 20 0 9.16034e-20 $X=8.24 $Y=1.005
c51 16 0 1.44655e-19 $X=7.39 $Y=1.1
c52 13 0 1.44963e-19 $X=10.03 $Y=0.515
r53 20 22 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=8.24 $Y=1.005
+ $X2=8.24 $Y2=1.18
r54 16 18 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=7.43 $Y=1.1 $X2=7.43
+ $Y2=1.18
r55 11 13 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=9.99 $Y=0.92
+ $X2=9.99 $Y2=0.515
r56 10 20 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.325 $Y=1.005
+ $X2=8.24 $Y2=1.005
r57 9 11 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.865 $Y=1.005
+ $X2=9.99 $Y2=0.92
r58 9 10 100.471 $w=1.68e-07 $l=1.54e-06 $layer=LI1_cond $X=9.865 $Y=1.005
+ $X2=8.325 $Y2=1.005
r59 8 18 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.555 $Y=1.18
+ $X2=7.43 $Y2=1.18
r60 7 22 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.155 $Y=1.18
+ $X2=8.24 $Y2=1.18
r61 7 8 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=8.155 $Y=1.18 $X2=7.555
+ $Y2=1.18
r62 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.89
+ $Y=0.37 $X2=10.03 $Y2=0.515
r63 1 16 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=7.25
+ $Y=0.605 $X2=7.39 $Y2=1.1
.ends


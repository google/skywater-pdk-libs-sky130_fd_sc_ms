* File: sky130_fd_sc_ms__fahcin_1.pex.spice
* Created: Wed Sep  2 12:09:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__FAHCIN_1%A 3 7 9 15 16
r34 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.71
+ $Y=1.515 $X2=0.71 $Y2=1.515
r35 13 15 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.515 $Y=1.515
+ $X2=0.71 $Y2=1.515
r36 11 13 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.5 $Y=1.515
+ $X2=0.515 $Y2=1.515
r37 9 16 5.96091 $w=2.88e-07 $l=1.5e-07 $layer=LI1_cond $X=0.69 $Y=1.665
+ $X2=0.69 $Y2=1.515
r38 5 13 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.68
+ $X2=0.515 $Y2=1.515
r39 5 7 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=0.515 $Y=1.68
+ $X2=0.515 $Y2=2.4
r40 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.35 $X2=0.5
+ $Y2=1.515
r41 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.5 $Y=1.35 $X2=0.5
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCIN_1%A_28_74# 1 2 3 4 15 19 23 27 31 33 34 36 37
+ 38 39 40 43 47 49 57
c106 34 0 1.71384e-19 $X=1.09 $Y=2.905
r107 53 57 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=1.28 $Y=1.465
+ $X2=1.41 $Y2=1.465
r108 53 54 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.28 $Y=1.465
+ $X2=1.205 $Y2=1.465
r109 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.28
+ $Y=1.465 $X2=1.28 $Y2=1.465
r110 50 52 12.2997 $w=3.67e-07 $l=3.7e-07 $layer=LI1_cond $X=1.225 $Y=1.095
+ $X2=1.225 $Y2=1.465
r111 45 47 21.8964 $w=2.48e-07 $l=4.75e-07 $layer=LI1_cond $X=3.81 $Y=2.905
+ $X2=3.81 $Y2=2.43
r112 41 43 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2.71 $Y=0.425
+ $X2=2.71 $Y2=0.55
r113 39 41 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.585 $Y=0.34
+ $X2=2.71 $Y2=0.425
r114 39 40 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=2.585 $Y=0.34
+ $X2=1.29 $Y2=0.34
r115 37 45 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.685 $Y=2.99
+ $X2=3.81 $Y2=2.905
r116 37 38 163.754 $w=1.68e-07 $l=2.51e-06 $layer=LI1_cond $X=3.685 $Y=2.99
+ $X2=1.175 $Y2=2.99
r117 36 50 6.3706 $w=3.67e-07 $l=9.44722e-08 $layer=LI1_cond $X=1.205 $Y=1.01
+ $X2=1.225 $Y2=1.095
r118 35 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.205 $Y=0.425
+ $X2=1.29 $Y2=0.34
r119 35 36 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.205 $Y=0.425
+ $X2=1.205 $Y2=1.01
r120 34 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.09 $Y=2.905
+ $X2=1.175 $Y2=2.99
r121 33 52 9.03 $w=3.67e-07 $l=2.22486e-07 $layer=LI1_cond $X=1.09 $Y=1.63
+ $X2=1.225 $Y2=1.465
r122 33 34 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=1.09 $Y=1.63
+ $X2=1.09 $Y2=2.905
r123 32 49 3.35233 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.45 $Y=1.095
+ $X2=0.285 $Y2=1.095
r124 31 50 5.25812 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=1.005 $Y=1.095
+ $X2=1.225 $Y2=1.095
r125 31 32 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.005 $Y=1.095
+ $X2=0.45 $Y2=1.095
r126 27 29 37.5109 $w=2.53e-07 $l=8.3e-07 $layer=LI1_cond $X=0.247 $Y=1.985
+ $X2=0.247 $Y2=2.815
r127 25 49 3.22182 $w=2.92e-07 $l=1.0225e-07 $layer=LI1_cond $X=0.247 $Y=1.18
+ $X2=0.285 $Y2=1.095
r128 25 27 36.381 $w=2.53e-07 $l=8.05e-07 $layer=LI1_cond $X=0.247 $Y=1.18
+ $X2=0.247 $Y2=1.985
r129 21 49 3.22182 $w=2.92e-07 $l=8.5e-08 $layer=LI1_cond $X=0.285 $Y=1.01
+ $X2=0.285 $Y2=1.095
r130 21 23 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.285 $Y=1.01
+ $X2=0.285 $Y2=0.515
r131 17 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.3
+ $X2=1.41 $Y2=1.465
r132 17 19 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.41 $Y=1.3
+ $X2=1.41 $Y2=0.79
r133 13 54 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.205 $Y=1.63
+ $X2=1.205 $Y2=1.465
r134 13 15 275.984 $w=1.8e-07 $l=7.1e-07 $layer=POLY_cond $X=1.205 $Y=1.63
+ $X2=1.205 $Y2=2.34
r135 4 47 600 $w=1.7e-07 $l=6.20645e-07 $layer=licon1_PDIFF $count=1 $X=3.665
+ $Y=1.895 $X2=3.85 $Y2=2.43
r136 3 29 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.29 $Y2=2.815
r137 3 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.84 $X2=0.29 $Y2=1.985
r138 2 43 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=2.61 $Y=0.37
+ $X2=2.75 $Y2=0.55
r139 1 23 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.37 $X2=0.285 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCIN_1%A_492_48# 1 2 9 13 19 23 27 31 33 35 36 37
+ 41 42 44 45 49 51 52 54 60 62 65 72
c173 72 0 6.47663e-20 $X=6.09 $Y=1.42
c174 31 0 1.21008e-19 $X=6.09 $Y=0.725
c175 27 0 1.532e-19 $X=5.91 $Y=2.34
c176 9 0 1.01566e-19 $X=2.535 $Y=0.69
r177 71 72 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=5.91 $Y=1.42
+ $X2=6.09 $Y2=1.42
r178 64 66 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.575 $Y=1.545
+ $X2=3.645 $Y2=1.545
r179 64 65 16.9689 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.575 $Y=1.545
+ $X2=3.485 $Y2=1.545
r180 61 71 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=5.84 $Y=1.42 $X2=5.91
+ $Y2=1.42
r181 60 63 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=5.8 $Y=1.42
+ $X2=5.8 $Y2=1.585
r182 60 62 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=5.8 $Y=1.42
+ $X2=5.8 $Y2=1.255
r183 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.84
+ $Y=1.42 $X2=5.84 $Y2=1.42
r184 54 57 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=5.12 $Y=1.905
+ $X2=5.12 $Y2=2.055
r185 52 66 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=3.825 $Y=1.545
+ $X2=3.645 $Y2=1.545
r186 51 53 18.2271 $w=2.51e-07 $l=3.75e-07 $layer=LI1_cond $X=3.825 $Y=1.545
+ $X2=4.2 $Y2=1.545
r187 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.825
+ $Y=1.545 $X2=3.825 $Y2=1.545
r188 49 63 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.715 $Y=1.82
+ $X2=5.715 $Y2=1.585
r189 46 62 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.715 $Y=1.01
+ $X2=5.715 $Y2=1.255
r190 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.63 $Y=0.925
+ $X2=5.715 $Y2=1.01
r191 44 45 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.63 $Y=0.925
+ $X2=5.295 $Y2=0.925
r192 43 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.285 $Y=1.905
+ $X2=5.12 $Y2=1.905
r193 42 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.63 $Y=1.905
+ $X2=5.715 $Y2=1.82
r194 42 43 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.63 $Y=1.905
+ $X2=5.285 $Y2=1.905
r195 39 45 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.13 $Y=0.84
+ $X2=5.295 $Y2=0.925
r196 39 41 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.13 $Y=0.84
+ $X2=5.13 $Y2=0.585
r197 38 41 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=5.13 $Y=0.425
+ $X2=5.13 $Y2=0.585
r198 36 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.965 $Y=0.34
+ $X2=5.13 $Y2=0.425
r199 36 37 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.965 $Y=0.34
+ $X2=4.285 $Y2=0.34
r200 35 53 3.01842 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.2 $Y=1.38 $X2=4.2
+ $Y2=1.545
r201 34 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.2 $Y=0.425
+ $X2=4.285 $Y2=0.34
r202 34 35 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=4.2 $Y=0.425
+ $X2=4.2 $Y2=1.38
r203 29 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.09 $Y=1.255
+ $X2=6.09 $Y2=1.42
r204 29 31 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.09 $Y=1.255
+ $X2=6.09 $Y2=0.725
r205 25 71 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=5.91 $Y=1.585
+ $X2=5.91 $Y2=1.42
r206 25 27 293.476 $w=1.8e-07 $l=7.55e-07 $layer=POLY_cond $X=5.91 $Y=1.585
+ $X2=5.91 $Y2=2.34
r207 21 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.645 $Y=1.38
+ $X2=3.645 $Y2=1.545
r208 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.645 $Y=1.38
+ $X2=3.645 $Y2=0.915
r209 17 64 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.575 $Y=1.71
+ $X2=3.575 $Y2=1.545
r210 17 19 235.169 $w=1.8e-07 $l=6.05e-07 $layer=POLY_cond $X=3.575 $Y=1.71
+ $X2=3.575 $Y2=2.315
r211 16 33 2.09011 $w=2.85e-07 $l=9e-08 $layer=POLY_cond $X=2.64 $Y=1.522
+ $X2=2.55 $Y2=1.522
r212 16 65 177.856 $w=2.85e-07 $l=8.45e-07 $layer=POLY_cond $X=2.64 $Y=1.522
+ $X2=3.485 $Y2=1.522
r213 11 33 31.2989 $w=1.65e-07 $l=1.43e-07 $layer=POLY_cond $X=2.55 $Y=1.665
+ $X2=2.55 $Y2=1.522
r214 11 13 328.46 $w=1.8e-07 $l=8.45e-07 $layer=POLY_cond $X=2.55 $Y=1.665
+ $X2=2.55 $Y2=2.51
r215 7 33 31.2989 $w=1.65e-07 $l=1.49312e-07 $layer=POLY_cond $X=2.535 $Y=1.38
+ $X2=2.55 $Y2=1.522
r216 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.535 $Y=1.38
+ $X2=2.535 $Y2=0.69
r217 2 57 600 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=1 $X=4.975
+ $Y=1.84 $X2=5.12 $Y2=2.055
r218 1 41 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=4.985
+ $Y=0.405 $X2=5.13 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCIN_1%B 1 3 6 8 9 10 11 14 18 20 22 25 27 30 32
+ 34 35 36 38 39 40 41
c136 27 0 1.27399e-19 $X=4.835 $Y=1.255
c137 18 0 3.79173e-20 $X=4.305 $Y=0.915
c138 14 0 2.11348e-20 $X=4.29 $Y=2.315
c139 8 0 9.05624e-20 $X=4.23 $Y=0.18
c140 6 0 9.79869e-20 $X=3.04 $Y=2.51
r141 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.04
+ $Y=1.42 $X2=5.04 $Y2=1.42
r142 41 45 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=5.04 $Y=1.295
+ $X2=5.04 $Y2=1.42
r143 39 44 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=5.255 $Y=1.42
+ $X2=5.04 $Y2=1.42
r144 39 40 3.90195 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.255 $Y=1.42
+ $X2=5.345 $Y2=1.42
r145 37 44 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=4.91 $Y=1.42
+ $X2=5.04 $Y2=1.42
r146 37 38 5.03009 $w=3.3e-07 $l=1.67332e-07 $layer=POLY_cond $X=4.91 $Y=1.42
+ $X2=4.75 $Y2=1.435
r147 32 40 34.7346 $w=1.65e-07 $l=1.72337e-07 $layer=POLY_cond $X=5.36 $Y=1.255
+ $X2=5.345 $Y2=1.42
r148 32 34 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.36 $Y=1.255
+ $X2=5.36 $Y2=0.775
r149 28 40 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=5.345 $Y=1.585
+ $X2=5.345 $Y2=1.42
r150 28 30 316.798 $w=1.8e-07 $l=8.15e-07 $layer=POLY_cond $X=5.345 $Y=1.585
+ $X2=5.345 $Y2=2.4
r151 27 38 37.0704 $w=1.5e-07 $l=2.18403e-07 $layer=POLY_cond $X=4.835 $Y=1.255
+ $X2=4.75 $Y2=1.435
r152 26 27 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=4.835 $Y=0.255
+ $X2=4.835 $Y2=1.255
r153 24 38 37.0704 $w=1.5e-07 $l=1.83712e-07 $layer=POLY_cond $X=4.825 $Y=1.585
+ $X2=4.75 $Y2=1.435
r154 24 25 764.021 $w=1.5e-07 $l=1.49e-06 $layer=POLY_cond $X=4.825 $Y=1.585
+ $X2=4.825 $Y2=3.075
r155 23 35 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.38 $Y=3.15 $X2=4.29
+ $Y2=3.15
r156 22 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.75 $Y=3.15
+ $X2=4.825 $Y2=3.075
r157 22 23 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.75 $Y=3.15
+ $X2=4.38 $Y2=3.15
r158 21 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.38 $Y=0.18
+ $X2=4.305 $Y2=0.18
r159 20 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.76 $Y=0.18
+ $X2=4.835 $Y2=0.255
r160 20 21 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=4.76 $Y=0.18
+ $X2=4.38 $Y2=0.18
r161 16 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.305 $Y=0.255
+ $X2=4.305 $Y2=0.18
r162 16 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.305 $Y=0.255
+ $X2=4.305 $Y2=0.915
r163 12 35 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.29 $Y=3.075
+ $X2=4.29 $Y2=3.15
r164 12 14 295.419 $w=1.8e-07 $l=7.6e-07 $layer=POLY_cond $X=4.29 $Y=3.075
+ $X2=4.29 $Y2=2.315
r165 10 35 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.2 $Y=3.15 $X2=4.29
+ $Y2=3.15
r166 10 11 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=4.2 $Y=3.15
+ $X2=3.13 $Y2=3.15
r167 8 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.23 $Y=0.18
+ $X2=4.305 $Y2=0.18
r168 8 9 610.191 $w=1.5e-07 $l=1.19e-06 $layer=POLY_cond $X=4.23 $Y=0.18
+ $X2=3.04 $Y2=0.18
r169 4 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.04 $Y=3.075
+ $X2=3.13 $Y2=3.15
r170 4 6 219.621 $w=1.8e-07 $l=5.65e-07 $layer=POLY_cond $X=3.04 $Y=3.075
+ $X2=3.04 $Y2=2.51
r171 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.965 $Y=0.255
+ $X2=3.04 $Y2=0.18
r172 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.965 $Y=0.255
+ $X2=2.965 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCIN_1%A_608_74# 1 2 9 11 13 17 18 20 22 29 33 35
+ 38 39 40 42 43 44 46 48 49 50 52 53 56 57 58 60 61 63 64 67 68 70 71 75 79 88
c267 88 0 4.231e-20 $X=8.085 $Y=1.32
c268 70 0 3.23e-19 $X=6.605 $Y=1.675
c269 67 0 2.11348e-20 $X=3.35 $Y=2.04
c270 63 0 2.11268e-20 $X=10.41 $Y=0.405
c271 35 0 3.79173e-20 $X=4.105 $Y=1.965
r272 76 88 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=7.91 $Y=1.32
+ $X2=8.085 $Y2=1.32
r273 75 78 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=7.89 $Y=1.32
+ $X2=7.89 $Y2=1.485
r274 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.91
+ $Y=1.32 $X2=7.91 $Y2=1.32
r275 71 82 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=6.605 $Y=1.675
+ $X2=6.495 $Y2=1.675
r276 70 73 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=6.605 $Y=1.675
+ $X2=6.605 $Y2=1.84
r277 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.605
+ $Y=1.675 $X2=6.605 $Y2=1.675
r278 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.41
+ $Y=0.405 $X2=10.41 $Y2=0.405
r279 61 63 37.5001 $w=3.13e-07 $l=1.025e-06 $layer=LI1_cond $X=9.385 $Y=0.412
+ $X2=10.41 $Y2=0.412
r280 59 61 7.64049 $w=3.15e-07 $l=1.95944e-07 $layer=LI1_cond $X=9.3 $Y=0.57
+ $X2=9.385 $Y2=0.412
r281 59 60 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=9.3 $Y=0.57
+ $X2=9.3 $Y2=1.655
r282 57 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.215 $Y=1.74
+ $X2=9.3 $Y2=1.655
r283 57 58 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=9.215 $Y=1.74
+ $X2=8.715 $Y2=1.74
r284 55 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.63 $Y=1.825
+ $X2=8.715 $Y2=1.74
r285 55 56 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=8.63 $Y=1.825
+ $X2=8.63 $Y2=2.905
r286 54 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.955 $Y=2.99
+ $X2=7.87 $Y2=2.99
r287 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.545 $Y=2.99
+ $X2=8.63 $Y2=2.905
r288 53 54 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.545 $Y=2.99
+ $X2=7.955 $Y2=2.99
r289 52 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.87 $Y=2.905
+ $X2=7.87 $Y2=2.99
r290 52 78 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=7.87 $Y=2.905
+ $X2=7.87 $Y2=1.485
r291 49 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.785 $Y=2.99
+ $X2=7.87 $Y2=2.99
r292 49 50 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=7.785 $Y=2.99
+ $X2=6.65 $Y2=2.99
r293 48 68 2.84813 $w=3.35e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.565 $Y=2.39
+ $X2=6.4 $Y2=2.475
r294 48 73 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=6.565 $Y=2.39
+ $X2=6.565 $Y2=1.84
r295 46 50 9.23067 $w=1.7e-07 $l=2.89396e-07 $layer=LI1_cond $X=6.4 $Y=2.905
+ $X2=6.65 $Y2=2.99
r296 45 68 2.84813 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=6.4 $Y=2.56 $X2=6.4
+ $Y2=2.475
r297 45 46 8.25294 $w=4.98e-07 $l=3.45e-07 $layer=LI1_cond $X=6.4 $Y=2.56
+ $X2=6.4 $Y2=2.905
r298 43 68 3.86674 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=6.15 $Y=2.475
+ $X2=6.4 $Y2=2.475
r299 43 44 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=6.15 $Y=2.475
+ $X2=5.045 $Y2=2.475
r300 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.96 $Y=2.56
+ $X2=5.045 $Y2=2.475
r301 41 42 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.96 $Y=2.56
+ $X2=4.96 $Y2=2.905
r302 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.875 $Y=2.99
+ $X2=4.96 $Y2=2.905
r303 39 40 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.875 $Y=2.99
+ $X2=4.275 $Y2=2.99
r304 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.19 $Y=2.905
+ $X2=4.275 $Y2=2.99
r305 37 38 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=4.19 $Y=2.05
+ $X2=4.19 $Y2=2.905
r306 36 67 2.76166 $w=1.7e-07 $l=1.66493e-07 $layer=LI1_cond $X=3.515 $Y=1.965
+ $X2=3.35 $Y2=1.962
r307 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.105 $Y=1.965
+ $X2=4.19 $Y2=2.05
r308 35 36 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.105 $Y=1.965
+ $X2=3.515 $Y2=1.965
r309 31 67 3.70735 $w=2.5e-07 $l=1.20536e-07 $layer=LI1_cond $X=3.43 $Y=1.875
+ $X2=3.35 $Y2=1.962
r310 31 33 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=3.43 $Y=1.875
+ $X2=3.43 $Y2=0.76
r311 27 67 3.70735 $w=2.5e-07 $l=8.8e-08 $layer=LI1_cond $X=3.35 $Y=2.05
+ $X2=3.35 $Y2=1.962
r312 27 29 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=3.35 $Y=2.05
+ $X2=3.35 $Y2=2.57
r313 22 64 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=10.02 $Y=0.405
+ $X2=10.41 $Y2=0.405
r314 18 23 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=10.205 $Y=1.47
+ $X2=9.945 $Y2=1.47
r315 18 20 309.024 $w=1.8e-07 $l=7.95e-07 $layer=POLY_cond $X=10.205 $Y=1.545
+ $X2=10.205 $Y2=2.34
r316 15 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.945 $Y=1.395
+ $X2=9.945 $Y2=1.47
r317 15 17 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=9.945 $Y=1.395
+ $X2=9.945 $Y2=1
r318 14 22 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=9.945 $Y=0.57
+ $X2=10.02 $Y2=0.405
r319 14 17 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.945 $Y=0.57
+ $X2=9.945 $Y2=1
r320 11 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.085 $Y=1.155
+ $X2=8.085 $Y2=1.32
r321 11 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.085 $Y=1.155
+ $X2=8.085 $Y2=0.725
r322 7 82 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=6.495 $Y=1.84
+ $X2=6.495 $Y2=1.675
r323 7 9 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=6.495 $Y=1.84
+ $X2=6.495 $Y2=2.42
r324 2 67 600 $w=1.7e-07 $l=2.43721e-07 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=2.09 $X2=3.35 $Y2=2.04
r325 2 29 600 $w=1.7e-07 $l=5.79655e-07 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=2.09 $X2=3.35 $Y2=2.57
r326 1 33 91 $w=1.7e-07 $l=5.51543e-07 $layer=licon1_NDIFF $count=2 $X=3.04
+ $Y=0.37 $X2=3.43 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCIN_1%A_430_418# 1 2 3 4 13 15 16 17 18 19 20 22
+ 25 27 29 34 38 40 42 43 44 45 46 47 50 54 59 63 64 69 70
c213 50 0 9.79869e-20 $X=2.16 $Y=2.035
c214 42 0 1.46093e-19 $X=4.415 $Y=2.035
c215 27 0 2.11268e-20 $X=10.89 $Y=1.43
c216 16 0 1.05034e-19 $X=7.205 $Y=1.195
r217 68 70 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=10.85 $Y=1.595
+ $X2=10.89 $Y2=1.595
r218 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.85
+ $Y=1.595 $X2=10.85 $Y2=1.595
r219 65 68 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=10.655 $Y=1.595
+ $X2=10.85 $Y2=1.595
r220 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.37
+ $Y=1.335 $X2=7.37 $Y2=1.335
r221 60 69 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=10.85 $Y=2.035
+ $X2=10.85 $Y2=1.595
r222 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=2.035
+ $X2=10.8 $Y2=2.035
r223 57 64 25.6098 $w=3.13e-07 $l=7e-07 $layer=LI1_cond $X=7.397 $Y=2.035
+ $X2=7.397 $Y2=1.335
r224 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=2.035
+ $X2=7.44 $Y2=2.035
r225 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=2.035
+ $X2=4.56 $Y2=2.035
r226 50 85 7.20241 $w=4.15e-07 $l=2.45e-07 $layer=LI1_cond $X=2.265 $Y=2.035
+ $X2=2.265 $Y2=2.28
r227 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=2.035
+ $X2=2.16 $Y2=2.035
r228 47 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.585 $Y=2.035
+ $X2=7.44 $Y2=2.035
r229 46 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=10.8 $Y2=2.035
r230 46 47 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=7.585 $Y2=2.035
r231 45 53 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.705 $Y=2.035
+ $X2=4.56 $Y2=2.035
r232 44 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.295 $Y=2.035
+ $X2=7.44 $Y2=2.035
r233 44 45 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=7.295 $Y=2.035
+ $X2=4.705 $Y2=2.035
r234 43 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=2.035
+ $X2=2.16 $Y2=2.035
r235 42 53 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.415 $Y=2.035
+ $X2=4.56 $Y2=2.035
r236 42 43 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=4.415 $Y=2.035
+ $X2=2.305 $Y2=2.035
r237 40 54 1.32974 $w=2.58e-07 $l=3e-08 $layer=LI1_cond $X=4.575 $Y=2.005
+ $X2=4.575 $Y2=2.035
r238 40 41 5.76222 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=4.575 $Y=2.005
+ $X2=4.575 $Y2=1.875
r239 38 41 44.0233 $w=2.48e-07 $l=9.55e-07 $layer=LI1_cond $X=4.58 $Y=0.92
+ $X2=4.58 $Y2=1.875
r240 32 50 6.17653 $w=4.15e-07 $l=1.57003e-07 $layer=LI1_cond $X=2.29 $Y=1.89
+ $X2=2.265 $Y2=2.035
r241 32 34 51.1685 $w=2.48e-07 $l=1.11e-06 $layer=LI1_cond $X=2.29 $Y=1.89
+ $X2=2.29 $Y2=0.78
r242 31 63 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=7.37 $Y=1.725
+ $X2=7.37 $Y2=1.335
r243 30 63 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=7.37 $Y=1.27
+ $X2=7.37 $Y2=1.335
r244 27 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.89 $Y=1.43
+ $X2=10.89 $Y2=1.595
r245 27 29 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=10.89 $Y=1.43
+ $X2=10.89 $Y2=1
r246 23 65 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.655 $Y=1.76
+ $X2=10.655 $Y2=1.595
r247 23 25 225.452 $w=1.8e-07 $l=5.8e-07 $layer=POLY_cond $X=10.655 $Y=1.76
+ $X2=10.655 $Y2=2.34
r248 20 22 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=7.9 $Y=1.875
+ $X2=7.9 $Y2=2.42
r249 19 31 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=7.535 $Y=1.8
+ $X2=7.37 $Y2=1.725
r250 18 20 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=7.81 $Y=1.8
+ $X2=7.9 $Y2=1.875
r251 18 19 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=7.81 $Y=1.8
+ $X2=7.535 $Y2=1.8
r252 16 30 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=7.205 $Y=1.195
+ $X2=7.37 $Y2=1.27
r253 16 17 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.205 $Y=1.195
+ $X2=6.595 $Y2=1.195
r254 13 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.52 $Y=1.12
+ $X2=6.595 $Y2=1.195
r255 13 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.52 $Y=1.12
+ $X2=6.52 $Y2=0.725
r256 4 54 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=4.38
+ $Y=1.895 $X2=4.53 $Y2=2.04
r257 3 85 600 $w=1.7e-07 $l=2.61534e-07 $layer=licon1_PDIFF $count=1 $X=2.15
+ $Y=2.09 $X2=2.32 $Y2=2.28
r258 2 38 182 $w=1.7e-07 $l=3.9702e-07 $layer=licon1_NDIFF $count=1 $X=4.38
+ $Y=0.595 $X2=4.54 $Y2=0.92
r259 1 34 182 $w=1.7e-07 $l=4.68348e-07 $layer=licon1_NDIFF $count=1 $X=2.195
+ $Y=0.37 $X2=2.32 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCIN_1%CIN 3 5 7 8 10 12 14 15
r60 18 20 48.5406 $w=2.83e-07 $l=2.85e-07 $layer=POLY_cond $X=8.585 $Y=1.35
+ $X2=8.87 $Y2=1.35
r61 17 18 16.1802 $w=2.83e-07 $l=9.5e-08 $layer=POLY_cond $X=8.49 $Y=1.35
+ $X2=8.585 $Y2=1.35
r62 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.87
+ $Y=1.32 $X2=8.87 $Y2=1.32
r63 12 14 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=9.47 $Y=1.395
+ $X2=9.47 $Y2=0.95
r64 8 12 46.8375 $w=2.83e-07 $l=3.4187e-07 $layer=POLY_cond $X=9.195 $Y=1.545
+ $X2=9.47 $Y2=1.395
r65 8 20 55.3534 $w=2.83e-07 $l=4.11096e-07 $layer=POLY_cond $X=9.195 $Y=1.545
+ $X2=8.87 $Y2=1.35
r66 8 10 332.347 $w=1.8e-07 $l=8.55e-07 $layer=POLY_cond $X=9.195 $Y=1.545
+ $X2=9.195 $Y2=2.4
r67 5 18 17.601 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=8.585 $Y=1.155
+ $X2=8.585 $Y2=1.35
r68 5 7 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.585 $Y=1.155
+ $X2=8.585 $Y2=0.725
r69 1 17 13.3727 $w=1.8e-07 $l=1.95e-07 $layer=POLY_cond $X=8.49 $Y=1.545
+ $X2=8.49 $Y2=1.35
r70 1 3 309.024 $w=1.8e-07 $l=7.95e-07 $layer=POLY_cond $X=8.49 $Y=1.545
+ $X2=8.49 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCIN_1%A_1857_368# 1 2 3 10 12 15 20 23 28 29 32
+ 34 35 36 39 40 45 50
r91 43 50 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=11.7 $Y=1.515
+ $X2=11.775 $Y2=1.515
r92 43 47 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=11.7 $Y=1.515
+ $X2=11.465 $Y2=1.515
r93 42 45 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=11.7 $Y=1.515
+ $X2=11.89 $Y2=1.515
r94 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.7
+ $Y=1.515 $X2=11.7 $Y2=1.515
r95 38 40 8.98215 $w=3.33e-07 $l=1.8e-07 $layer=LI1_cond $X=10.975 $Y=2.907
+ $X2=11.155 $Y2=2.907
r96 38 39 8.81015 $w=3.33e-07 $l=1.75e-07 $layer=LI1_cond $X=10.975 $Y=2.907
+ $X2=10.8 $Y2=2.907
r97 35 36 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=9.64 $Y=1.995
+ $X2=9.64 $Y2=1.34
r98 34 35 7.30169 $w=4.68e-07 $l=8.5e-08 $layer=LI1_cond $X=9.49 $Y=2.08
+ $X2=9.49 $Y2=1.995
r99 31 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.89 $Y=1.68
+ $X2=11.89 $Y2=1.515
r100 31 32 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=11.89 $Y=1.68
+ $X2=11.89 $Y2=2.905
r101 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.805 $Y=2.99
+ $X2=11.89 $Y2=2.905
r102 29 40 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=11.805 $Y=2.99
+ $X2=11.155 $Y2=2.99
r103 28 39 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=9.725 $Y=2.99
+ $X2=10.8 $Y2=2.99
r104 21 36 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.72 $Y=1.175
+ $X2=9.72 $Y2=1.34
r105 21 23 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=9.72 $Y=1.175
+ $X2=9.72 $Y2=0.825
r106 18 28 8.97637 $w=1.7e-07 $l=2.74226e-07 $layer=LI1_cond $X=9.49 $Y=2.905
+ $X2=9.725 $Y2=2.99
r107 18 20 2.29036 $w=4.68e-07 $l=9e-08 $layer=LI1_cond $X=9.49 $Y=2.905
+ $X2=9.49 $Y2=2.815
r108 17 34 3.81727 $w=4.68e-07 $l=1.5e-07 $layer=LI1_cond $X=9.49 $Y=2.23
+ $X2=9.49 $Y2=2.08
r109 17 20 14.8874 $w=4.68e-07 $l=5.85e-07 $layer=LI1_cond $X=9.49 $Y=2.23
+ $X2=9.49 $Y2=2.815
r110 13 50 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=11.775 $Y=1.68
+ $X2=11.775 $Y2=1.515
r111 13 15 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=11.775 $Y=1.68
+ $X2=11.775 $Y2=2.34
r112 10 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.465 $Y=1.35
+ $X2=11.465 $Y2=1.515
r113 10 12 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=11.465 $Y=1.35
+ $X2=11.465 $Y2=0.92
r114 3 38 600 $w=1.7e-07 $l=1.09397e-06 $layer=licon1_PDIFF $count=1 $X=10.745
+ $Y=1.92 $X2=10.975 $Y2=2.905
r115 2 34 400 $w=1.7e-07 $l=3e-07 $layer=licon1_PDIFF $count=1 $X=9.285 $Y=1.84
+ $X2=9.42 $Y2=2.08
r116 2 20 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=9.285
+ $Y=1.84 $X2=9.42 $Y2=2.815
r117 1 23 91 $w=1.7e-07 $l=3.2078e-07 $layer=licon1_NDIFF $count=2 $X=9.545
+ $Y=0.58 $X2=9.72 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCIN_1%A_2004_136# 1 2 9 11 13 16 19 20 21 23 24
+ 25 28 35 40
r84 39 40 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=12.455 $Y=1.515
+ $X2=12.465 $Y2=1.515
r85 34 35 3.56523 $w=5.18e-07 $l=1.55e-07 $layer=LI1_cond $X=10.675 $Y=1
+ $X2=10.83 $Y2=1
r86 31 34 6.55543 $w=5.18e-07 $l=2.85e-07 $layer=LI1_cond $X=10.39 $Y=1
+ $X2=10.675 $Y2=1
r87 29 39 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=12.285 $Y=1.515
+ $X2=12.455 $Y2=1.515
r88 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.285
+ $Y=1.515 $X2=12.285 $Y2=1.515
r89 26 28 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=12.285 $Y=1.18
+ $X2=12.285 $Y2=1.515
r90 24 26 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=12.145 $Y=1.095
+ $X2=12.285 $Y2=1.18
r91 24 25 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=12.145 $Y=1.095
+ $X2=11.755 $Y2=1.095
r92 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.67 $Y=1.01
+ $X2=11.755 $Y2=1.095
r93 22 23 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=11.67 $Y=0.49
+ $X2=11.67 $Y2=1.01
r94 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.585 $Y=0.405
+ $X2=11.67 $Y2=0.49
r95 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=11.585 $Y=0.405
+ $X2=10.915 $Y2=0.405
r96 19 35 7.40362 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=10.83 $Y=0.74
+ $X2=10.83 $Y2=1
r97 18 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.83 $Y=0.49
+ $X2=10.915 $Y2=0.405
r98 18 19 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=10.83 $Y=0.49
+ $X2=10.83 $Y2=0.74
r99 14 31 5.03516 $w=2.5e-07 $l=2.6e-07 $layer=LI1_cond $X=10.39 $Y=1.26
+ $X2=10.39 $Y2=1
r100 14 16 37.1087 $w=2.48e-07 $l=8.05e-07 $layer=LI1_cond $X=10.39 $Y=1.26
+ $X2=10.39 $Y2=2.065
r101 11 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.465 $Y=1.35
+ $X2=12.465 $Y2=1.515
r102 11 13 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=12.465 $Y=1.35
+ $X2=12.465 $Y2=0.87
r103 7 39 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=12.455 $Y=1.68
+ $X2=12.455 $Y2=1.515
r104 7 9 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=12.455 $Y=1.68
+ $X2=12.455 $Y2=2.4
r105 2 16 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.295
+ $Y=1.92 $X2=10.43 $Y2=2.065
r106 1 34 45.5 $w=1.7e-07 $l=7.23878e-07 $layer=licon1_NDIFF $count=4 $X=10.02
+ $Y=0.68 $X2=10.675 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCIN_1%VPWR 1 2 3 4 15 21 25 29 34 35 36 38 43 58
+ 67 68 71 74 77
r101 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r102 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r103 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r104 68 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=12.24 $Y2=3.33
r105 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r106 65 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.395 $Y=3.33
+ $X2=12.27 $Y2=3.33
r107 65 67 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=12.395 $Y=3.33
+ $X2=12.72 $Y2=3.33
r108 64 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r109 63 64 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r110 61 64 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=11.76 $Y2=3.33
r111 60 63 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=9.36 $Y=3.33
+ $X2=11.76 $Y2=3.33
r112 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r113 58 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.145 $Y=3.33
+ $X2=12.27 $Y2=3.33
r114 58 63 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=12.145 $Y=3.33
+ $X2=11.76 $Y2=3.33
r115 57 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r116 56 57 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r117 54 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r118 53 56 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=8.88
+ $Y2=3.33
r119 53 54 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6 $Y=3.33
+ $X2=6 $Y2=3.33
r120 51 74 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=5.765 $Y=3.33
+ $X2=5.585 $Y2=3.33
r121 51 53 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.765 $Y=3.33
+ $X2=6 $Y2=3.33
r122 50 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r123 49 50 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r124 47 50 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=5.04 $Y2=3.33
r125 47 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r126 46 49 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=5.04 $Y2=3.33
r127 46 47 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r128 44 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.825 $Y=3.33
+ $X2=0.7 $Y2=3.33
r129 44 46 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.825 $Y=3.33
+ $X2=1.2 $Y2=3.33
r130 43 74 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=5.405 $Y=3.33
+ $X2=5.585 $Y2=3.33
r131 43 49 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.405 $Y=3.33
+ $X2=5.04 $Y2=3.33
r132 41 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r133 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r134 38 71 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.7 $Y2=3.33
r135 38 40 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.24 $Y2=3.33
r136 36 57 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=8.88 $Y2=3.33
r137 36 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r138 34 56 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=8.885 $Y=3.33
+ $X2=8.88 $Y2=3.33
r139 34 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.885 $Y=3.33
+ $X2=8.97 $Y2=3.33
r140 33 60 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.055 $Y=3.33
+ $X2=9.36 $Y2=3.33
r141 33 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.055 $Y=3.33
+ $X2=8.97 $Y2=3.33
r142 29 32 36.8782 $w=2.48e-07 $l=8e-07 $layer=LI1_cond $X=12.27 $Y=2.015
+ $X2=12.27 $Y2=2.815
r143 27 77 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.27 $Y=3.245
+ $X2=12.27 $Y2=3.33
r144 27 32 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=12.27 $Y=3.245
+ $X2=12.27 $Y2=2.815
r145 23 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.97 $Y=3.245
+ $X2=8.97 $Y2=3.33
r146 23 25 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=8.97 $Y=3.245
+ $X2=8.97 $Y2=2.16
r147 19 74 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.585 $Y=3.245
+ $X2=5.585 $Y2=3.33
r148 19 21 13.7653 $w=3.58e-07 $l=4.3e-07 $layer=LI1_cond $X=5.585 $Y=3.245
+ $X2=5.585 $Y2=2.815
r149 15 18 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=0.7 $Y=2.115 $X2=0.7
+ $Y2=2.815
r150 13 71 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=3.245
+ $X2=0.7 $Y2=3.33
r151 13 18 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.7 $Y=3.245 $X2=0.7
+ $Y2=2.815
r152 4 32 400 $w=1.7e-07 $l=1.14302e-06 $layer=licon1_PDIFF $count=1 $X=11.865
+ $Y=1.84 $X2=12.23 $Y2=2.815
r153 4 29 400 $w=1.7e-07 $l=4.43959e-07 $layer=licon1_PDIFF $count=1 $X=11.865
+ $Y=1.84 $X2=12.23 $Y2=2.015
r154 3 25 300 $w=1.7e-07 $l=5.26213e-07 $layer=licon1_PDIFF $count=2 $X=8.58
+ $Y=1.84 $X2=8.97 $Y2=2.16
r155 2 21 600 $w=1.7e-07 $l=1.04732e-06 $layer=licon1_PDIFF $count=1 $X=5.435
+ $Y=1.84 $X2=5.585 $Y2=2.815
r156 1 18 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.84 $X2=0.74 $Y2=2.815
r157 1 15 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.84 $X2=0.74 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCIN_1%A_259_368# 1 2 3 4 14 17 18 19 20 22 26 27
+ 28 31 34 35 39 41 46
c93 46 0 9.05624e-20 $X=3.09 $Y=1.005
c94 28 0 1.01566e-19 $X=3.175 $Y=0.34
c95 4 0 1.46093e-19 $X=2.64 $Y=2.09
r96 44 46 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.895 $Y=1.005
+ $X2=3.09 $Y2=1.005
r97 37 39 2.84554 $w=4.03e-07 $l=1e-07 $layer=LI1_cond $X=1.625 $Y=0.817
+ $X2=1.725 $Y2=0.817
r98 34 35 7.7063 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=1.59 $Y=1.985
+ $X2=1.59 $Y2=1.82
r99 29 31 21.8964 $w=2.48e-07 $l=4.75e-07 $layer=LI1_cond $X=3.82 $Y=0.425
+ $X2=3.82 $Y2=0.9
r100 27 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.695 $Y=0.34
+ $X2=3.82 $Y2=0.425
r101 27 28 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.695 $Y=0.34
+ $X2=3.175 $Y2=0.34
r102 26 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.09 $Y=0.92
+ $X2=3.09 $Y2=1.005
r103 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.09 $Y=0.425
+ $X2=3.175 $Y2=0.34
r104 25 26 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=3.09 $Y=0.425
+ $X2=3.09 $Y2=0.92
r105 23 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=1.09
+ $X2=2.895 $Y2=1.005
r106 23 41 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=2.895 $Y=1.09
+ $X2=2.895 $Y2=2.045
r107 20 43 2.65806 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=2.817 $Y=2.565
+ $X2=2.817 $Y2=2.65
r108 20 22 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=2.817 $Y=2.565
+ $X2=2.817 $Y2=2.225
r109 19 41 8.35379 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=2.817 $Y=2.207
+ $X2=2.817 $Y2=2.045
r110 19 22 0.638276 $w=3.23e-07 $l=1.8e-08 $layer=LI1_cond $X=2.817 $Y=2.207
+ $X2=2.817 $Y2=2.225
r111 17 43 5.06595 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=2.655 $Y=2.65
+ $X2=2.817 $Y2=2.65
r112 17 18 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=2.655 $Y=2.65
+ $X2=1.835 $Y2=2.65
r113 15 39 4.30998 $w=2.2e-07 $l=2.03e-07 $layer=LI1_cond $X=1.725 $Y=1.02
+ $X2=1.725 $Y2=0.817
r114 15 35 41.907 $w=2.18e-07 $l=8e-07 $layer=LI1_cond $X=1.725 $Y=1.02
+ $X2=1.725 $Y2=1.82
r115 14 18 9.14635 $w=1.7e-07 $l=2.84341e-07 $layer=LI1_cond $X=1.59 $Y=2.565
+ $X2=1.835 $Y2=2.65
r116 13 34 1.95278 $w=4.88e-07 $l=8e-08 $layer=LI1_cond $X=1.59 $Y=2.065
+ $X2=1.59 $Y2=1.985
r117 13 14 12.2049 $w=4.88e-07 $l=5e-07 $layer=LI1_cond $X=1.59 $Y=2.065
+ $X2=1.59 $Y2=2.565
r118 4 43 600 $w=1.7e-07 $l=6.41561e-07 $layer=licon1_PDIFF $count=1 $X=2.64
+ $Y=2.09 $X2=2.815 $Y2=2.65
r119 4 22 600 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=2.64
+ $Y=2.09 $X2=2.815 $Y2=2.225
r120 3 34 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.295
+ $Y=1.84 $X2=1.43 $Y2=1.985
r121 2 31 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=3.72
+ $Y=0.595 $X2=3.86 $Y2=0.9
r122 1 37 182 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.47 $X2=1.625 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCIN_1%A_1200_368# 1 2 9 14 15 17
r39 15 17 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=6.225 $Y=1.82
+ $X2=6.225 $Y2=1.065
r40 14 15 10.8446 $w=3.38e-07 $l=2.35e-07 $layer=LI1_cond $X=6.14 $Y=2.055
+ $X2=6.14 $Y2=1.82
r41 7 17 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.305 $Y=0.9
+ $X2=6.305 $Y2=1.065
r42 7 9 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=6.305 $Y=0.9 $X2=6.305
+ $Y2=0.55
r43 2 14 600 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=6 $Y=1.84
+ $X2=6.135 $Y2=2.055
r44 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.165
+ $Y=0.405 $X2=6.305 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCIN_1%COUT 1 2 8 11 14 21 22
c48 14 0 1.63318e-19 $X=6.805 $Y=0.56
r49 21 22 9.43695 $w=5.43e-07 $l=4.3e-07 $layer=LI1_cond $X=7.44 $Y=0.712
+ $X2=7.87 $Y2=0.712
r50 21 26 6.14499 $w=5.43e-07 $l=2.8e-07 $layer=LI1_cond $X=7.44 $Y=0.712
+ $X2=7.16 $Y2=0.712
r51 17 26 1.97518 $w=5.43e-07 $l=9e-08 $layer=LI1_cond $X=7.07 $Y=0.712 $X2=7.16
+ $Y2=0.712
r52 17 18 20.3897 $w=4.28e-07 $l=5.98e-07 $layer=LI1_cond $X=6.855 $Y=0.712
+ $X2=6.855 $Y2=1.31
r53 14 17 4.07375 $w=4.28e-07 $l=1.52e-07 $layer=LI1_cond $X=6.855 $Y=0.56
+ $X2=6.855 $Y2=0.712
r54 9 20 2.94173 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=7.07 $Y=2.5 $X2=6.945
+ $Y2=2.5
r55 9 11 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.07 $Y=2.5 $X2=7.5
+ $Y2=2.5
r56 8 20 4.82444 $w=1.7e-07 $l=1.83916e-07 $layer=LI1_cond $X=6.985 $Y=2.335
+ $X2=6.945 $Y2=2.5
r57 8 18 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=6.985 $Y=2.335
+ $X2=6.985 $Y2=1.31
r58 2 20 600 $w=1.7e-07 $l=6.46142e-07 $layer=licon1_PDIFF $count=1 $X=6.585
+ $Y=2 $X2=6.92 $Y2=2.5
r59 2 11 600 $w=1.7e-07 $l=1.13786e-06 $layer=licon1_PDIFF $count=1 $X=6.585
+ $Y=2 $X2=7.5 $Y2=2.5
r60 1 22 60.6667 $w=1.7e-07 $l=1.35028e-06 $layer=licon1_NDIFF $count=3 $X=6.595
+ $Y=0.405 $X2=7.87 $Y2=0.56
r61 1 26 60.6667 $w=1.7e-07 $l=6.37809e-07 $layer=licon1_NDIFF $count=3 $X=6.595
+ $Y=0.405 $X2=7.16 $Y2=0.56
r62 1 14 91 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_NDIFF $count=2 $X=6.595
+ $Y=0.405 $X2=6.805 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCIN_1%A_1598_400# 1 2 7 9 13 17 18
r29 17 18 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=8.29 $Y=1.82
+ $X2=8.29 $Y2=1.065
r30 11 18 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=8.37 $Y=0.9
+ $X2=8.37 $Y2=1.065
r31 11 13 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=8.37 $Y=0.9 $X2=8.37
+ $Y2=0.55
r32 7 17 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=8.25 $Y=1.945
+ $X2=8.25 $Y2=1.82
r33 7 9 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=8.25 $Y=1.945 $X2=8.25
+ $Y2=1.985
r34 2 9 300 $w=1.7e-07 $l=2.27376e-07 $layer=licon1_PDIFF $count=2 $X=7.99 $Y=2
+ $X2=8.21 $Y2=1.985
r35 1 13 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=8.16
+ $Y=0.405 $X2=8.37 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCIN_1%A_1967_384# 1 2 3 10 12 14 18 20 23 29 30
c48 20 0 8.64817e-20 $X=11.28 $Y=1.25
r49 29 30 8.83531 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=11.415 $Y=2.015
+ $X2=11.415 $Y2=1.85
r50 22 29 1.44055 $w=4.38e-07 $l=5.5e-08 $layer=LI1_cond $X=11.415 $Y=2.07
+ $X2=11.415 $Y2=2.015
r51 22 23 8.64332 $w=4.38e-07 $l=3.3e-07 $layer=LI1_cond $X=11.415 $Y=2.07
+ $X2=11.415 $Y2=2.4
r52 20 27 7.81924 $w=3.22e-07 $l=1.49248e-07 $layer=LI1_cond $X=11.28 $Y=1.25
+ $X2=11.25 $Y2=1.115
r53 20 30 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=11.28 $Y=1.25
+ $X2=11.28 $Y2=1.85
r54 16 27 2.21818 $w=3.3e-07 $l=6e-08 $layer=LI1_cond $X=11.25 $Y=1.055
+ $X2=11.25 $Y2=1.115
r55 16 18 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=11.25 $Y=1.055
+ $X2=11.25 $Y2=0.745
r56 15 25 3.40825 $w=1.7e-07 $l=1.19143e-07 $layer=LI1_cond $X=10.065 $Y=2.485
+ $X2=9.98 $Y2=2.567
r57 14 23 14.5445 $w=1.82e-07 $l=2.59037e-07 $layer=LI1_cond $X=11.195 $Y=2.485
+ $X2=11.415 $Y2=2.4
r58 14 15 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=11.195 $Y=2.485
+ $X2=10.065 $Y2=2.485
r59 10 25 3.40825 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=9.98 $Y=2.4 $X2=9.98
+ $Y2=2.567
r60 10 12 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.98 $Y=2.4
+ $X2=9.98 $Y2=2.065
r61 3 29 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=11.405
+ $Y=1.84 $X2=11.55 $Y2=2.015
r62 2 25 600 $w=1.7e-07 $l=7.18853e-07 $layer=licon1_PDIFF $count=1 $X=9.835
+ $Y=1.92 $X2=9.98 $Y2=2.57
r63 2 12 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=9.835
+ $Y=1.92 $X2=9.98 $Y2=2.065
r64 1 27 182 $w=1.7e-07 $l=5.59643e-07 $layer=licon1_NDIFF $count=1 $X=10.965
+ $Y=0.68 $X2=11.25 $Y2=1.115
r65 1 18 182 $w=1.7e-07 $l=3.15832e-07 $layer=licon1_NDIFF $count=1 $X=10.965
+ $Y=0.68 $X2=11.25 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCIN_1%SUM 1 2 7 8 9 10 11 12 13
r14 12 13 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=12.72 $Y=2.405
+ $X2=12.72 $Y2=2.775
r15 11 12 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=12.72 $Y=1.985
+ $X2=12.72 $Y2=2.405
r16 10 11 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=12.72 $Y=1.665
+ $X2=12.72 $Y2=1.985
r17 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=12.72 $Y=1.295
+ $X2=12.72 $Y2=1.665
r18 9 26 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=12.72 $Y=1.295
+ $X2=12.72 $Y2=1.095
r19 8 44 5.50001 $w=4.18e-07 $l=1.8e-07 $layer=LI1_cond $X=12.68 $Y=0.84
+ $X2=12.68 $Y2=0.66
r20 8 26 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=12.72 $Y=0.925
+ $X2=12.72 $Y2=1.095
r21 7 44 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=12.68 $Y=0.555
+ $X2=12.68 $Y2=0.66
r22 2 13 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=12.545
+ $Y=1.84 $X2=12.68 $Y2=2.815
r23 2 11 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=12.545
+ $Y=1.84 $X2=12.68 $Y2=1.985
r24 1 44 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=12.54
+ $Y=0.5 $X2=12.68 $Y2=0.66
r25 1 26 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=12.54
+ $Y=0.5 $X2=12.68 $Y2=1.095
.ends

.subckt PM_SKY130_FD_SC_MS__FAHCIN_1%VGND 1 2 3 4 15 19 23 27 29 31 36 41 49 59
+ 60 63 66 69 72
c116 19 0 1.27399e-19 $X=5.715 $Y=0.55
r117 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r118 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r119 66 67 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r120 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r121 60 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r122 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r123 57 72 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=12.345 $Y=0
+ $X2=12.135 $Y2=0
r124 57 59 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=12.345 $Y=0
+ $X2=12.72 $Y2=0
r125 56 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r126 55 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r127 53 56 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=11.76 $Y2=0
r128 53 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=8.88
+ $Y2=0
r129 52 55 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=9.36 $Y=0 $X2=11.76
+ $Y2=0
r130 52 53 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r131 50 69 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=9.045 $Y=0 $X2=8.875
+ $Y2=0
r132 50 52 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.045 $Y=0
+ $X2=9.36 $Y2=0
r133 49 72 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=11.925 $Y=0
+ $X2=12.135 $Y2=0
r134 49 55 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=11.925 $Y=0
+ $X2=11.76 $Y2=0
r135 48 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r136 47 48 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r137 45 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r138 44 47 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=6 $Y=0 $X2=8.4
+ $Y2=0
r139 44 45 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=0 $X2=6 $Y2=0
r140 42 66 11.3601 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=5.97 $Y=0 $X2=5.717
+ $Y2=0
r141 42 44 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=5.97 $Y=0 $X2=6 $Y2=0
r142 41 69 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=8.705 $Y=0 $X2=8.875
+ $Y2=0
r143 41 47 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.705 $Y=0 $X2=8.4
+ $Y2=0
r144 40 67 1.20413 $w=4.9e-07 $l=4.32e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=5.52
+ $Y2=0
r145 40 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r146 39 40 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r147 37 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.785
+ $Y2=0
r148 37 39 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.2
+ $Y2=0
r149 36 66 11.3601 $w=1.7e-07 $l=2.52e-07 $layer=LI1_cond $X=5.465 $Y=0
+ $X2=5.717 $Y2=0
r150 36 39 278.251 $w=1.68e-07 $l=4.265e-06 $layer=LI1_cond $X=5.465 $Y=0
+ $X2=1.2 $Y2=0
r151 34 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r152 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r153 31 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.785
+ $Y2=0
r154 31 33 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.24
+ $Y2=0
r155 29 48 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r156 29 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r157 25 72 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=12.135 $Y=0.085
+ $X2=12.135 $Y2=0
r158 25 27 15.3659 $w=4.18e-07 $l=5.6e-07 $layer=LI1_cond $X=12.135 $Y=0.085
+ $X2=12.135 $Y2=0.645
r159 21 69 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=8.875 $Y=0.085
+ $X2=8.875 $Y2=0
r160 21 23 15.7614 $w=3.38e-07 $l=4.65e-07 $layer=LI1_cond $X=8.875 $Y=0.085
+ $X2=8.875 $Y2=0.55
r161 17 66 2.09999 $w=5.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.717 $Y=0.085
+ $X2=5.717 $Y2=0
r162 17 19 11.0134 $w=5.03e-07 $l=4.65e-07 $layer=LI1_cond $X=5.717 $Y=0.085
+ $X2=5.717 $Y2=0.55
r163 13 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0
r164 13 15 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0.675
r165 4 27 182 $w=1.7e-07 $l=5.77062e-07 $layer=licon1_NDIFF $count=1 $X=11.54
+ $Y=0.6 $X2=12.095 $Y2=0.645
r166 3 23 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=8.66
+ $Y=0.405 $X2=8.875 $Y2=0.55
r167 2 19 182 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_NDIFF $count=1 $X=5.435
+ $Y=0.405 $X2=5.715 $Y2=0.55
r168 1 15 182 $w=1.7e-07 $l=3.96327e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.37 $X2=0.785 $Y2=0.675
.ends


* File: sky130_fd_sc_ms__o41a_4.spice
* Created: Wed Sep  2 12:27:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o41a_4.pex.spice"
.subckt sky130_fd_sc_ms__o41a_4  VNB VPB B1 A4 A3 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1010 N_X_M1010_d N_A_110_48#_M1010_g N_VGND_M1010_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2627 PD=1.02 PS=2.19 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75000.3
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1017 N_X_M1010_d N_A_110_48#_M1017_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.7
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1020 N_X_M1020_d N_A_110_48#_M1020_g N_VGND_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75001.2
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1024 N_X_M1020_d N_A_110_48#_M1024_g N_VGND_M1024_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.6
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1005 N_A_523_124#_M1005_d N_B1_M1005_g N_A_110_48#_M1005_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1824 AS=0.0896 PD=1.85 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75004.5 A=0.096 P=1.58 MULT=1
MM1016 N_A_523_124#_M1016_d N_B1_M1016_g N_A_110_48#_M1005_s VNB NLOWVT L=0.15
+ W=0.64 AD=0.1184 AS=0.0896 PD=1.01 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75004 A=0.096 P=1.58 MULT=1
MM1004 N_A_523_124#_M1016_d N_A3_M1004_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1184 AS=0.19135 PD=1.01 PS=1.26 NRD=16.872 NRS=60 M=1 R=4.26667
+ SA=75001.2 SB=75003.5 A=0.096 P=1.58 MULT=1
MM1000 N_A_523_124#_M1000_d N_A4_M1000_g N_VGND_M1004_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.19135 PD=0.92 PS=1.26 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.9
+ SB=75002.9 A=0.096 P=1.58 MULT=1
MM1027 N_A_523_124#_M1000_d N_A4_M1027_g N_VGND_M1027_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.3
+ SB=75002.4 A=0.096 P=1.58 MULT=1
MM1018 N_A_523_124#_M1018_d N_A3_M1018_g N_VGND_M1027_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0928 AS=0.0896 PD=0.93 PS=0.92 NRD=0.936 NRS=0 M=1 R=4.26667 SA=75002.7
+ SB=75002 A=0.096 P=1.58 MULT=1
MM1008 N_A_523_124#_M1018_d N_A2_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0928 AS=0.0896 PD=0.93 PS=0.92 NRD=0.936 NRS=0 M=1 R=4.26667 SA=75003.2
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1012 N_A_523_124#_M1012_d N_A1_M1012_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75003.6
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1013 N_A_523_124#_M1012_d N_A1_M1013_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.0896 AS=0.113125 PD=0.92 PS=1.005 NRD=0 NRS=0 M=1 R=4.26667 SA=75004
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1022 N_A_523_124#_M1022_d N_A2_M1022_g N_VGND_M1013_s VNB NLOWVT L=0.15 W=0.64
+ AD=0.1824 AS=0.113125 PD=1.85 PS=1.005 NRD=0 NRS=13.116 M=1 R=4.26667
+ SA=75004.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1003 N_X_M1003_d N_A_110_48#_M1003_g N_VPWR_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90002.3 A=0.2016 P=2.6 MULT=1
MM1006 N_X_M1003_d N_A_110_48#_M1006_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90001.8 A=0.2016 P=2.6 MULT=1
MM1007 N_X_M1007_d N_A_110_48#_M1007_g N_VPWR_M1006_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90001.4 A=0.2016 P=2.6 MULT=1
MM1009 N_X_M1007_d N_A_110_48#_M1009_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.211943 PD=1.39 PS=1.68571 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.5
+ SB=90000.9 A=0.2016 P=2.6 MULT=1
MM1011 N_A_110_48#_M1011_d N_B1_M1011_g N_VPWR_M1009_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.158957 PD=1.11 PS=1.26429 NRD=0 NRS=18.7544 M=1 R=4.66667
+ SA=90002.1 SB=90000.6 A=0.1512 P=2.04 MULT=1
MM1014 N_A_110_48#_M1011_d N_B1_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=0.84
+ AD=0.1134 AS=0.2352 PD=1.11 PS=2.24 NRD=0 NRS=0 M=1 R=4.66667 SA=90002.5
+ SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1015 N_A_854_368#_M1015_d N_A3_M1015_g N_A_762_368#_M1015_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90003.5 A=0.2016 P=2.6 MULT=1
MM1019 N_A_110_48#_M1019_d N_A4_M1019_g N_A_854_368#_M1015_d VPB PSHORT L=0.18
+ W=1.12 AD=0.1568 AS=0.1512 PD=1.4 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.6
+ SB=90003 A=0.2016 P=2.6 MULT=1
MM1021 N_A_110_48#_M1019_d N_A4_M1021_g N_A_854_368#_M1021_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1568 AS=0.1512 PD=1.4 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.1
+ SB=90002.6 A=0.2016 P=2.6 MULT=1
MM1023 N_A_854_368#_M1021_s N_A3_M1023_g N_A_762_368#_M1023_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90001.5 SB=90002.1 A=0.2016 P=2.6 MULT=1
MM1002 N_A_762_368#_M1023_s N_A2_M1002_g N_A_1216_368#_M1002_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90002
+ SB=90001.7 A=0.2016 P=2.6 MULT=1
MM1001 N_A_1216_368#_M1002_s N_A1_M1001_g N_VPWR_M1001_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1736 PD=1.39 PS=1.43 NRD=0 NRS=2.6201 M=1 R=6.22222
+ SA=90002.4 SB=90001.2 A=0.2016 P=2.6 MULT=1
MM1026 N_A_1216_368#_M1026_d N_A1_M1026_g N_VPWR_M1001_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1792 AS=0.1736 PD=1.44 PS=1.43 NRD=7.8997 NRS=2.6201 M=1 R=6.22222
+ SA=90002.9 SB=90000.7 A=0.2016 P=2.6 MULT=1
MM1025 N_A_762_368#_M1025_d N_A2_M1025_g N_A_1216_368#_M1026_d VPB PSHORT L=0.18
+ W=1.12 AD=0.3696 AS=0.1792 PD=2.9 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222
+ SA=90003.4 SB=90000.2 A=0.2016 P=2.6 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.8844 P=20.8
*
.include "sky130_fd_sc_ms__o41a_4.pxi.spice"
*
.ends
*
*

* NGSPICE file created from sky130_fd_sc_ms__sdfrbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_ms__sdfrbp_1 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 Q a_2513_424# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=2.912e+11p pd=2.76e+06u as=2.27097e+12p ps=1.957e+07u
M1001 VPWR SCD a_515_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=2.304e+11p ps=2e+06u
M1002 a_413_90# D a_312_90# VNB nlowvt w=420000u l=150000u
+  ad=3.26375e+11p pd=3.3e+06u as=1.491e+11p ps=1.55e+06u
M1003 VGND a_1747_74# a_2513_424# VNB nlowvt w=550000u l=150000u
+  ad=1.78918e+12p pd=1.476e+07u as=1.4575e+11p ps=1.63e+06u
M1004 a_1399_119# a_1369_93# a_1321_119# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.008e+11p ps=1.32e+06u
M1005 VGND a_2008_48# a_1966_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1006 VPWR a_1369_93# a_1331_463# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1007 a_1369_93# a_1235_119# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1008 VPWR a_1747_74# a_2513_424# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.184e+11p ps=2.2e+06u
M1009 a_2124_74# RESET_B VGND VNB nlowvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1010 Q_N a_1747_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1011 a_413_90# RESET_B VPWR VPB pshort w=640000u l=180000u
+  ad=4.654e+11p pd=5.04e+06u as=0p ps=0u
M1012 a_2008_48# a_1747_74# a_2124_74# VNB nlowvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1013 VGND CLK a_819_119# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.54e+11p ps=2.22e+06u
M1014 a_1037_119# a_819_119# VGND VNB nlowvt w=740000u l=150000u
+  ad=1.998e+11p pd=2.02e+06u as=0p ps=0u
M1015 a_1747_74# a_819_119# a_1369_93# VPB pshort w=1e+06u l=180000u
+  ad=3.9355e+11p pd=3.45e+06u as=0p ps=0u
M1016 a_1966_74# a_819_119# a_1747_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=4.519e+11p ps=3.17e+06u
M1017 a_341_464# SCE VPWR VPB pshort w=640000u l=180000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1018 VPWR SCE a_27_74# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=5.696e+11p ps=3.06e+06u
M1019 a_1235_119# a_1037_119# a_413_90# VPB pshort w=420000u l=180000u
+  ad=2.268e+11p pd=2.76e+06u as=0p ps=0u
M1020 a_2008_48# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1021 VPWR a_1747_74# a_2008_48# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_225_90# SCD a_545_97# VNB nlowvt w=420000u l=150000u
+  ad=2.64075e+11p pd=2.99e+06u as=8.82e+10p ps=1.26e+06u
M1023 a_312_90# a_27_74# a_225_90# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1331_463# a_819_119# a_1235_119# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR CLK a_819_119# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=3.136e+11p ps=2.8e+06u
M1026 Q_N a_1747_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1027 a_413_90# D a_341_464# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VGND RESET_B a_225_90# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1747_74# a_1037_119# a_1369_93# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=1.792e+11p ps=1.84e+06u
M1030 a_515_464# a_27_74# a_413_90# VPB pshort w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1235_119# a_819_119# a_413_90# VNB nlowvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1032 a_545_97# SCE a_413_90# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1972_489# a_1037_119# a_1747_74# VPB pshort w=420000u l=180000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1034 VGND RESET_B a_1399_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1037_119# a_819_119# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1036 a_1321_119# a_1037_119# a_1235_119# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 Q a_2513_424# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1038 VGND SCE a_27_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1039 VPWR a_2008_48# a_1972_489# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1235_119# RESET_B VPWR VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_1369_93# a_1235_119# VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


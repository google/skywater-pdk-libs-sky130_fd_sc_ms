* File: sky130_fd_sc_ms__o221ai_1.pex.spice
* Created: Wed Sep  2 12:23:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__O221AI_1%C1 3 7 9 13 14
r28 12 14 38.0526 $w=2.85e-07 $l=2.25e-07 $layer=POLY_cond $X=0.27 $Y=1.465
+ $X2=0.495 $Y2=1.465
r29 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.465 $X2=0.27 $Y2=1.465
r30 9 13 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.27 $Y=1.665 $X2=0.27
+ $Y2=1.465
r31 5 14 23.6772 $w=2.85e-07 $l=2.24332e-07 $layer=POLY_cond $X=0.635 $Y=1.63
+ $X2=0.495 $Y2=1.465
r32 5 7 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=0.635 $Y=1.63
+ $X2=0.635 $Y2=2.4
r33 1 14 17.7656 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=1.465
r34 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3 $X2=0.495
+ $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__O221AI_1%B1 5 9 11 14 15
r35 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.47
+ $Y=1.515 $X2=1.47 $Y2=1.515
r36 11 15 2.67779 $w=6.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.3 $Y=1.665 $X2=1.3
+ $Y2=1.515
r37 7 14 34.7346 $w=1.65e-07 $l=1.69926e-07 $layer=POLY_cond $X=1.555 $Y=1.35
+ $X2=1.545 $Y2=1.515
r38 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.555 $Y=1.35
+ $X2=1.555 $Y2=0.74
r39 3 14 34.7346 $w=1.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.545 $Y=1.68
+ $X2=1.545 $Y2=1.515
r40 3 5 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.545 $Y=1.68
+ $X2=1.545 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O221AI_1%B2 3 7 9 12 13
c39 7 0 6.24822e-20 $X=2.055 $Y=0.74
r40 12 15 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.04 $Y=1.515
+ $X2=2.04 $Y2=1.68
r41 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.04 $Y=1.515
+ $X2=2.04 $Y2=1.35
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.04
+ $Y=1.515 $X2=2.04 $Y2=1.515
r43 9 13 4.32166 $w=3.98e-07 $l=1.5e-07 $layer=LI1_cond $X=2.075 $Y=1.665
+ $X2=2.075 $Y2=1.515
r44 7 14 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.055 $Y=0.74
+ $X2=2.055 $Y2=1.35
r45 3 15 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=1.965 $Y=2.4
+ $X2=1.965 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O221AI_1%A2 3 7 9 10 11 12 19 20 36
c45 7 0 1.42066e-19 $X=2.555 $Y=0.74
r46 36 37 1.2285 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=1.68
r47 19 22 40.6903 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.61 $Y=1.515
+ $X2=2.61 $Y2=1.68
r48 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.61 $Y=1.515
+ $X2=2.61 $Y2=1.35
r49 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.515 $X2=2.61 $Y2=1.515
r50 11 12 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.65 $Y=2.405
+ $X2=2.65 $Y2=2.775
r51 10 11 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.65 $Y=2.035
+ $X2=2.65 $Y2=2.405
r52 9 36 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=2.61 $Y=1.63 $X2=2.61
+ $Y2=1.665
r53 9 20 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.61 $Y=1.63
+ $X2=2.61 $Y2=1.515
r54 9 10 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=2.65 $Y=1.715
+ $X2=2.65 $Y2=2.035
r55 9 37 1.61342 $w=2.48e-07 $l=3.5e-08 $layer=LI1_cond $X=2.65 $Y=1.715
+ $X2=2.65 $Y2=1.68
r56 7 21 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.555 $Y=0.74
+ $X2=2.555 $Y2=1.35
r57 3 22 279.871 $w=1.8e-07 $l=7.2e-07 $layer=POLY_cond $X=2.535 $Y=2.4
+ $X2=2.535 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_MS__O221AI_1%A1 3 7 9 10 17
r28 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.52
+ $Y=1.465 $X2=3.52 $Y2=1.465
r29 15 17 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=3.345 $Y=1.465
+ $X2=3.52 $Y2=1.465
r30 13 15 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=3.105 $Y=1.465
+ $X2=3.345 $Y2=1.465
r31 10 18 1.99346 $w=4.78e-07 $l=8e-08 $layer=LI1_cond $X=3.6 $Y=1.54 $X2=3.52
+ $Y2=1.54
r32 9 18 9.96732 $w=4.78e-07 $l=4e-07 $layer=LI1_cond $X=3.12 $Y=1.54 $X2=3.52
+ $Y2=1.54
r33 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.345 $Y=1.3
+ $X2=3.345 $Y2=1.465
r34 5 7 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.345 $Y=1.3 $X2=3.345
+ $Y2=0.74
r35 1 13 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.105 $Y=1.63
+ $X2=3.105 $Y2=1.465
r36 1 3 299.306 $w=1.8e-07 $l=7.7e-07 $layer=POLY_cond $X=3.105 $Y=1.63
+ $X2=3.105 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__O221AI_1%Y 1 2 3 12 15 16 17 18 20 28 29 40 44
r51 33 44 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=0.28 $Y=1.045
+ $X2=0.69 $Y2=1.045
r52 33 40 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.28 $Y=0.96
+ $X2=0.28 $Y2=0.925
r53 29 33 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=0.24 $Y=1.045 $X2=0.28
+ $Y2=1.045
r54 29 40 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.28 $Y=0.9
+ $X2=0.28 $Y2=0.925
r55 28 29 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.28 $Y=0.515
+ $X2=0.28 $Y2=0.9
r56 23 25 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.41 $Y=2.035
+ $X2=0.69 $Y2=2.035
r57 18 27 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=2.12 $X2=2.19
+ $Y2=2.035
r58 18 20 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.19 $Y=2.12
+ $X2=2.19 $Y2=2.815
r59 17 25 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=2.035
+ $X2=0.69 $Y2=2.035
r60 16 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=2.035
+ $X2=2.19 $Y2=2.035
r61 16 17 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=2.025 $Y=2.035
+ $X2=0.775 $Y2=2.035
r62 15 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.95
+ $X2=0.69 $Y2=2.035
r63 14 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.13
+ $X2=0.69 $Y2=1.045
r64 14 15 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=0.69 $Y=1.13
+ $X2=0.69 $Y2=1.95
r65 12 23 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=0.45 $Y=2.815
+ $X2=0.45 $Y2=2.12
r66 3 27 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=2.055
+ $Y=1.84 $X2=2.19 $Y2=2.115
r67 3 20 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.055
+ $Y=1.84 $X2=2.19 $Y2=2.815
r68 2 23 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.265
+ $Y=1.84 $X2=0.41 $Y2=2.115
r69 2 12 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.265
+ $Y=1.84 $X2=0.41 $Y2=2.815
r70 1 28 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__O221AI_1%VPWR 1 2 9 13 18 19 20 22 35 36 39
r37 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r38 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r39 33 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r40 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 30 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r42 29 32 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 27 39 14.7712 $w=1.7e-07 $l=4.08e-07 $layer=LI1_cond $X=1.56 $Y=3.33
+ $X2=1.152 $Y2=3.33
r45 27 29 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.56 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 22 39 14.7712 $w=1.7e-07 $l=4.07e-07 $layer=LI1_cond $X=0.745 $Y=3.33
+ $X2=1.152 $Y2=3.33
r49 22 24 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.745 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 20 33 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 20 30 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 18 32 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.165 $Y=3.33
+ $X2=3.12 $Y2=3.33
r53 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.165 $Y=3.33
+ $X2=3.33 $Y2=3.33
r54 17 35 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.495 $Y=3.33
+ $X2=3.6 $Y2=3.33
r55 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.495 $Y=3.33
+ $X2=3.33 $Y2=3.33
r56 13 16 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=3.33 $Y=2.115 $X2=3.33
+ $Y2=2.815
r57 11 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=3.245
+ $X2=3.33 $Y2=3.33
r58 11 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=3.33 $Y=3.245
+ $X2=3.33 $Y2=2.815
r59 7 39 3.16747 $w=8.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.152 $Y=3.245
+ $X2=1.152 $Y2=3.33
r60 7 9 12.768 $w=8.13e-07 $l=8.7e-07 $layer=LI1_cond $X=1.152 $Y=3.245
+ $X2=1.152 $Y2=2.375
r61 2 16 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.195
+ $Y=1.84 $X2=3.33 $Y2=2.815
r62 2 13 400 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=3.195
+ $Y=1.84 $X2=3.33 $Y2=2.115
r63 1 9 150 $w=1.7e-07 $l=8.19969e-07 $layer=licon1_PDIFF $count=4 $X=0.725
+ $Y=1.84 $X2=1.32 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_MS__O221AI_1%A_114_74# 1 2 7 9 14
c23 14 0 1.42066e-19 $X=1.84 $Y=0.435
c24 7 0 6.24822e-20 $X=1.675 $Y=0.435
r25 14 17 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=1.84 $Y=0.435
+ $X2=1.84 $Y2=0.63
r26 9 12 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=0.78 $Y=0.435
+ $X2=0.78 $Y2=0.605
r27 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0.435
+ $X2=0.78 $Y2=0.435
r28 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.675 $Y=0.435
+ $X2=1.84 $Y2=0.435
r29 7 8 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.675 $Y=0.435
+ $X2=0.945 $Y2=0.435
r30 2 17 182 $w=1.7e-07 $l=3.49571e-07 $layer=licon1_NDIFF $count=1 $X=1.63
+ $Y=0.37 $X2=1.84 $Y2=0.63
r31 1 12 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_MS__O221AI_1%A_239_74# 1 2 3 10 14 16 20 23 27
r46 23 25 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=1.34 $Y=0.965
+ $X2=1.34 $Y2=1.095
r47 18 20 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.56 $Y=0.96
+ $X2=3.56 $Y2=0.515
r48 17 27 8.61065 $w=1.7e-07 $l=1.77059e-07 $layer=LI1_cond $X=2.505 $Y=1.045
+ $X2=2.34 $Y2=1.07
r49 16 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.395 $Y=1.045
+ $X2=3.56 $Y2=0.96
r50 16 17 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=3.395 $Y=1.045
+ $X2=2.505 $Y2=1.045
r51 12 27 0.89609 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=2.34 $Y=0.96 $X2=2.34
+ $Y2=1.07
r52 12 14 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=2.34 $Y=0.96
+ $X2=2.34 $Y2=0.515
r53 11 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=1.095
+ $X2=1.34 $Y2=1.095
r54 10 27 8.61065 $w=1.7e-07 $l=1.77059e-07 $layer=LI1_cond $X=2.175 $Y=1.095
+ $X2=2.34 $Y2=1.07
r55 10 11 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.175 $Y=1.095
+ $X2=1.505 $Y2=1.095
r56 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.42
+ $Y=0.37 $X2=3.56 $Y2=0.515
r57 2 14 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=2.13
+ $Y=0.37 $X2=2.34 $Y2=0.515
r58 1 23 182 $w=1.7e-07 $l=6.63551e-07 $layer=licon1_NDIFF $count=1 $X=1.195
+ $Y=0.37 $X2=1.34 $Y2=0.965
.ends

.subckt PM_SKY130_FD_SC_MS__O221AI_1%VGND 1 6 8 10 20 21 24
r33 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r34 21 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r35 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r36 18 24 11.9488 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=3.225 $Y=0 $X2=2.95
+ $Y2=0
r37 18 20 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.225 $Y=0 $X2=3.6
+ $Y2=0
r38 17 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r39 16 17 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r40 12 16 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=2.64
+ $Y2=0
r41 12 13 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r42 10 24 11.9488 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.95
+ $Y2=0
r43 10 16 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.64
+ $Y2=0
r44 8 17 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r45 8 13 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=0.24
+ $Y2=0
r46 4 24 2.31338 $w=5.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.95 $Y=0.085 $X2=2.95
+ $Y2=0
r47 4 6 11.7433 $w=5.48e-07 $l=5.4e-07 $layer=LI1_cond $X=2.95 $Y=0.085 $X2=2.95
+ $Y2=0.625
r48 1 6 91 $w=1.7e-07 $l=6.1441e-07 $layer=licon1_NDIFF $count=2 $X=2.63 $Y=0.37
+ $X2=3.13 $Y2=0.625
.ends


* File: sky130_fd_sc_ms__o221ai_4.spice
* Created: Fri Aug 28 17:57:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_ms__o221ai_4.pex.spice"
.subckt sky130_fd_sc_ms__o221ai_4  VNB VPB C1 B1 B2 A1 A2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2	A2
* A1	A1
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1000 N_A_27_84#_M1000_d N_C1_M1000_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.2
+ SB=75001.5 A=0.111 P=1.78 MULT=1
MM1002 N_A_27_84#_M1002_d N_C1_M1002_g N_Y_M1000_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75000.6
+ SB=75001.1 A=0.111 P=1.78 MULT=1
MM1004 N_A_27_84#_M1002_d N_C1_M1004_g N_Y_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.1
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1018 N_A_27_84#_M1018_d N_C1_M1018_g N_Y_M1004_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75001.5
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1009 N_A_27_84#_M1009_d N_B1_M1009_g N_A_483_74#_M1009_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.2109 PD=1.02 PS=2.05 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.2 SB=75007 A=0.111 P=1.78 MULT=1
MM1011 N_A_27_84#_M1009_d N_B1_M1011_g N_A_483_74#_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75000.6 SB=75006.6 A=0.111 P=1.78 MULT=1
MM1030 N_A_27_84#_M1030_d N_B1_M1030_g N_A_483_74#_M1011_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.1 SB=75006.2 A=0.111 P=1.78 MULT=1
MM1006 N_A_483_74#_M1006_d N_B2_M1006_g N_A_27_84#_M1030_d VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.5 SB=75005.7 A=0.111 P=1.78 MULT=1
MM1015 N_A_483_74#_M1006_d N_B2_M1015_g N_A_27_84#_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75001.9 SB=75005.3 A=0.111 P=1.78 MULT=1
MM1016 N_A_483_74#_M1016_d N_B2_M1016_g N_A_27_84#_M1015_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.4 SB=75004.9 A=0.111 P=1.78 MULT=1
MM1026 N_A_483_74#_M1016_d N_B2_M1026_g N_A_27_84#_M1026_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1036 PD=1.02 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333
+ SA=75002.8 SB=75004.4 A=0.111 P=1.78 MULT=1
MM1037 N_A_27_84#_M1026_s N_B1_M1037_g N_A_483_74#_M1037_s VNB NLOWVT L=0.15
+ W=0.74 AD=0.1036 AS=0.1295 PD=1.02 PS=1.09 NRD=0 NRS=11.34 M=1 R=4.93333
+ SA=75003.2 SB=75004 A=0.111 P=1.78 MULT=1
MM1008 N_A_483_74#_M1037_s N_A1_M1008_g N_VGND_M1008_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1554 PD=1.09 PS=1.16 NRD=0 NRS=11.34 M=1 R=4.93333 SA=75003.7
+ SB=75003.5 A=0.111 P=1.78 MULT=1
MM1007 N_VGND_M1008_s N_A2_M1007_g N_A_483_74#_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1554 AS=0.1036 PD=1.16 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75004.3
+ SB=75002.9 A=0.111 P=1.78 MULT=1
MM1012 N_VGND_M1012_d N_A2_M1012_g N_A_483_74#_M1007_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75004.7
+ SB=75002.5 A=0.111 P=1.78 MULT=1
MM1017 N_VGND_M1012_d N_A2_M1017_g N_A_483_74#_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=11.34 NRS=0 M=1 R=4.93333 SA=75005.2
+ SB=75002 A=0.111 P=1.78 MULT=1
MM1019 N_VGND_M1019_d N_A2_M1019_g N_A_483_74#_M1017_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1073 AS=0.1036 PD=1.03 PS=1.02 NRD=0.804 NRS=0 M=1 R=4.93333 SA=75005.6
+ SB=75001.6 A=0.111 P=1.78 MULT=1
MM1027 N_A_483_74#_M1027_d N_A1_M1027_g N_VGND_M1019_d VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1073 PD=1.09 PS=1.03 NRD=11.34 NRS=0.804 M=1 R=4.93333
+ SA=75006.1 SB=75001.1 A=0.111 P=1.78 MULT=1
MM1031 N_A_483_74#_M1027_d N_A1_M1031_g N_VGND_M1031_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.1295 AS=0.1036 PD=1.09 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75006.6
+ SB=75000.6 A=0.111 P=1.78 MULT=1
MM1034 N_A_483_74#_M1034_d N_A1_M1034_g N_VGND_M1031_s VNB NLOWVT L=0.15 W=0.74
+ AD=0.2109 AS=0.1036 PD=2.05 PS=1.02 NRD=0 NRS=0 M=1 R=4.93333 SA=75007
+ SB=75000.2 A=0.111 P=1.78 MULT=1
MM1013 N_Y_M1013_d N_C1_M1013_g N_VPWR_M1013_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90000.2
+ SB=90009.3 A=0.2016 P=2.6 MULT=1
MM1014 N_Y_M1013_d N_C1_M1014_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1988 PD=1.39 PS=1.475 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90000.6
+ SB=90008.8 A=0.2016 P=2.6 MULT=1
MM1024 N_Y_M1024_d N_C1_M1024_g N_VPWR_M1014_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1652 AS=0.1988 PD=1.415 PS=1.475 NRD=3.5066 NRS=5.2599 M=1 R=6.22222
+ SA=90001.2 SB=90008.3 A=0.2016 P=2.6 MULT=1
MM1035 N_Y_M1024_d N_C1_M1035_g N_VPWR_M1035_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1652 AS=0.1792 PD=1.415 PS=1.44 NRD=0 NRS=0 M=1 R=6.22222 SA=90001.6
+ SB=90007.8 A=0.2016 P=2.6 MULT=1
MM1003 N_VPWR_M1035_s N_B1_M1003_g N_A_511_368#_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1512 PD=1.44 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90002.1
+ SB=90007.3 A=0.2016 P=2.6 MULT=1
MM1020 N_VPWR_M1020_d N_B1_M1020_g N_A_511_368#_M1003_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2072 AS=0.1512 PD=1.49 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90002.6
+ SB=90006.8 A=0.2016 P=2.6 MULT=1
MM1022 N_VPWR_M1020_d N_B1_M1022_g N_A_511_368#_M1022_s VPB PSHORT L=0.18 W=1.12
+ AD=0.2072 AS=0.1512 PD=1.49 PS=1.39 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90003.1
+ SB=90006.3 A=0.2016 P=2.6 MULT=1
MM1005 N_A_511_368#_M1022_s N_B2_M1005_g N_Y_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90003.6
+ SB=90005.8 A=0.2016 P=2.6 MULT=1
MM1025 N_A_511_368#_M1025_d N_B2_M1025_g N_Y_M1005_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90004
+ SB=90005.4 A=0.2016 P=2.6 MULT=1
MM1032 N_A_511_368#_M1025_d N_B2_M1032_g N_Y_M1032_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1792 PD=1.39 PS=1.44 NRD=0 NRS=7.8997 M=1 R=6.22222 SA=90004.5
+ SB=90004.9 A=0.2016 P=2.6 MULT=1
MM1036 N_A_511_368#_M1036_d N_B2_M1036_g N_Y_M1032_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1792 AS=0.1792 PD=1.44 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90005
+ SB=90004.4 A=0.2016 P=2.6 MULT=1
MM1028 N_VPWR_M1028_d N_B1_M1028_g N_A_511_368#_M1036_d VPB PSHORT L=0.18 W=1.12
+ AD=0.2072 AS=0.1792 PD=1.49 PS=1.44 NRD=7.8997 NRS=0 M=1 R=6.22222 SA=90005.5
+ SB=90003.9 A=0.2016 P=2.6 MULT=1
MM1001 N_A_1291_368#_M1001_d N_A1_M1001_g N_VPWR_M1028_d VPB PSHORT L=0.18
+ W=1.12 AD=0.182 AS=0.2072 PD=1.445 PS=1.49 NRD=0 NRS=7.8997 M=1 R=6.22222
+ SA=90006 SB=90003.4 A=0.2016 P=2.6 MULT=1
MM1021 N_Y_M1021_d N_A2_M1021_g N_A_1291_368#_M1001_d VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.182 PD=1.39 PS=1.445 NRD=0 NRS=8.7862 M=1 R=6.22222 SA=90006.6
+ SB=90002.9 A=0.2016 P=2.6 MULT=1
MM1023 N_Y_M1021_d N_A2_M1023_g N_A_1291_368#_M1023_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90007
+ SB=90002.4 A=0.2016 P=2.6 MULT=1
MM1029 N_Y_M1029_d N_A2_M1029_g N_A_1291_368#_M1023_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90007.5
+ SB=90002 A=0.2016 P=2.6 MULT=1
MM1033 N_Y_M1029_d N_A2_M1033_g N_A_1291_368#_M1033_s VPB PSHORT L=0.18 W=1.12
+ AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222 SA=90007.9
+ SB=90001.5 A=0.2016 P=2.6 MULT=1
MM1010 N_A_1291_368#_M1033_s N_A1_M1010_g N_VPWR_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90008.4 SB=90001.1 A=0.2016 P=2.6 MULT=1
MM1038 N_A_1291_368#_M1038_d N_A1_M1038_g N_VPWR_M1010_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.1512 PD=1.39 PS=1.39 NRD=0 NRS=0 M=1 R=6.22222
+ SA=90008.8 SB=90000.6 A=0.2016 P=2.6 MULT=1
MM1039 N_A_1291_368#_M1038_d N_A1_M1039_g N_VPWR_M1039_s VPB PSHORT L=0.18
+ W=1.12 AD=0.1512 AS=0.3136 PD=1.39 PS=2.8 NRD=0 NRS=0 M=1 R=6.22222 SA=90009.3
+ SB=90000.2 A=0.2016 P=2.6 MULT=1
DX40_noxref VNB VPB NWDIODE A=19.4556 P=24.64
*
.include "sky130_fd_sc_ms__o221ai_4.pxi.spice"
*
.ends
*
*

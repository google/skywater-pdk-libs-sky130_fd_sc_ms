# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__a2111oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__a2111oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.350000 4.675000 1.780000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.625200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.850000 1.350000 5.180000 1.780000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.514200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.180000 3.715000 1.550000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.514200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.505000 1.350000 2.755000 1.780000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  0.514200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.350000 1.315000 1.780000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  0.994300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.010000 2.500000 1.180000 ;
        RECT 0.125000 1.180000 0.355000 1.950000 ;
        RECT 0.125000 1.950000 1.085000 2.120000 ;
        RECT 0.755000 2.120000 1.085000 2.735000 ;
        RECT 1.160000 0.350000 1.490000 1.010000 ;
        RECT 2.170000 0.350000 2.500000 0.770000 ;
        RECT 2.170000 0.770000 4.330000 0.975000 ;
        RECT 2.170000 0.975000 2.500000 1.010000 ;
        RECT 4.000000 0.975000 4.330000 1.130000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.305000  2.290000 0.555000 2.905000 ;
      RECT 0.305000  2.905000 2.435000 3.075000 ;
      RECT 0.660000  0.085000 0.990000 0.840000 ;
      RECT 1.285000  1.950000 1.455000 2.905000 ;
      RECT 1.655000  1.950000 3.325000 2.120000 ;
      RECT 1.655000  2.120000 1.985000 2.735000 ;
      RECT 1.660000  0.085000 2.000000 0.840000 ;
      RECT 2.185000  2.290000 2.435000 2.905000 ;
      RECT 2.625000  2.290000 2.905000 2.905000 ;
      RECT 2.625000  2.905000 3.855000 3.075000 ;
      RECT 3.075000  1.820000 3.325000 1.950000 ;
      RECT 3.075000  2.120000 3.325000 2.735000 ;
      RECT 3.525000  1.950000 5.655000 2.120000 ;
      RECT 3.525000  2.120000 3.855000 2.905000 ;
      RECT 3.570000  0.350000 4.680000 0.600000 ;
      RECT 4.055000  2.290000 4.225000 3.245000 ;
      RECT 4.425000  2.120000 4.675000 2.980000 ;
      RECT 4.510000  0.600000 4.680000 1.010000 ;
      RECT 4.510000  1.010000 5.630000 1.180000 ;
      RECT 4.860000  0.085000 5.200000 0.840000 ;
      RECT 4.875000  2.290000 5.205000 3.245000 ;
      RECT 5.380000  0.350000 5.630000 1.010000 ;
      RECT 5.405000  1.820000 5.655000 1.950000 ;
      RECT 5.405000  2.120000 5.655000 2.980000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_ms__a2111oi_2
END LIBRARY

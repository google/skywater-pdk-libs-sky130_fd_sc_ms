* NGSPICE file created from sky130_fd_sc_ms__dlrbn_2.ext - technology: sky130A

.subckt sky130_fd_sc_ms__dlrbn_2 D GATE_N RESET_B VGND VNB VPB VPWR Q Q_N
M1000 VPWR a_838_48# Q VPB pshort w=1.12e+06u l=180000u
+  ad=2.6628e+12p pd=2.07e+07u as=3.024e+11p ps=2.78e+06u
M1001 a_1066_74# a_670_74# a_838_48# VNB nlowvt w=740000u l=150000u
+  ad=1.776e+11p pd=1.96e+06u as=2.109e+11p ps=2.05e+06u
M1002 VGND RESET_B a_1066_74# VNB nlowvt w=740000u l=150000u
+  ad=1.80345e+12p pd=1.499e+07u as=0p ps=0u
M1003 Q a_838_48# VGND VNB nlowvt w=740000u l=150000u
+  ad=2.072e+11p pd=2.04e+06u as=0p ps=0u
M1004 VPWR a_838_48# a_786_508# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=1.869e+11p ps=1.73e+06u
M1005 VPWR a_230_74# a_363_74# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=3.704e+11p ps=2.85e+06u
M1006 a_592_74# a_27_112# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.536e+11p pd=1.76e+06u as=0p ps=0u
M1007 a_670_74# a_230_74# a_592_74# VNB nlowvt w=640000u l=150000u
+  ad=2.44e+11p pd=2.18e+06u as=0p ps=0u
M1008 Q_N a_1448_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.024e+11p pd=2.78e+06u as=0p ps=0u
M1009 a_598_392# a_27_112# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.1e+11p pd=2.42e+06u as=0p ps=0u
M1010 VPWR a_1448_74# Q_N VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_838_48# a_670_74# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=3.136e+11p pd=2.8e+06u as=0p ps=0u
M1012 VPWR D a_27_112# VPB pshort w=840000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1013 a_230_74# GATE_N VGND VNB nlowvt w=740000u l=150000u
+  ad=2.109e+11p pd=2.05e+06u as=0p ps=0u
M1014 a_786_508# a_230_74# a_670_74# VPB pshort w=420000u l=180000u
+  ad=0p pd=0u as=3.265e+11p ps=2.74e+06u
M1015 a_230_74# GATE_N VPWR VPB pshort w=840000u l=180000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1016 VGND D a_27_112# VNB nlowvt w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1017 a_790_74# a_363_74# a_670_74# VNB nlowvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1018 a_1448_74# a_838_48# VGND VNB nlowvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1019 VGND a_838_48# Q VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_1448_74# Q_N VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.368e+11p ps=2.12e+06u
M1021 a_1448_74# a_838_48# VPWR VPB pshort w=1e+06u l=180000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1022 VGND a_230_74# a_363_74# VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=2.109e+11p ps=2.05e+06u
M1023 VGND a_838_48# a_790_74# VNB nlowvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_670_74# a_363_74# a_598_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Q a_838_48# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR RESET_B a_838_48# VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Q_N a_1448_74# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends


* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__dfbbp_1 CLK D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
X0 a_1318_119# a_214_74# a_1314_424# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X1 a_1474_446# a_1062_93# a_1708_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X2 a_1062_93# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8 w=640000u l=180000u
X3 VGND SET_B a_1708_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X4 VPWR D a_422_125# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X5 a_1020_379# a_1062_93# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X6 a_1421_508# a_1474_446# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X7 VPWR SET_B a_1474_446# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X8 VPWR SET_B a_671_93# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X9 a_2320_410# a_1474_446# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X10 a_716_379# a_671_93# VPWR VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X11 a_671_93# a_1062_93# a_872_119# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X12 a_2320_410# a_1474_446# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X13 a_1474_446# a_1314_424# a_1817_392# VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X14 a_872_119# a_520_87# a_671_93# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X15 a_1314_424# a_214_74# a_1421_508# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X16 a_1062_93# RESET_B VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X17 a_1314_424# a_27_74# a_1498_74# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X18 a_671_93# a_520_87# a_1020_379# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X19 a_606_87# a_671_93# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X20 VGND a_1474_446# Q_N VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X21 VPWR a_27_74# a_214_74# VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X22 VPWR a_671_93# a_1206_379# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X23 a_520_87# a_214_74# a_606_87# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X24 a_1498_74# a_1474_446# VGND VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X25 a_520_87# a_27_74# a_716_379# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X26 a_422_125# a_214_74# a_520_87# VPB sky130_fd_pr__pfet_01v8 w=420000u l=180000u
X27 a_422_125# a_27_74# a_520_87# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X28 VGND a_27_74# a_214_74# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X29 a_1817_392# a_1062_93# VPWR VPB sky130_fd_pr__pfet_01v8 w=1e+06u l=180000u
X30 VGND SET_B a_872_119# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X31 VGND a_671_93# a_1318_119# VNB sky130_fd_pr__nfet_01v8_lvt w=550000u l=150000u
X32 VPWR a_1474_446# Q_N VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X33 VGND a_2320_410# Q VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X34 a_27_74# CLK VPWR VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
X35 a_27_74# CLK VGND VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X36 a_1206_379# a_27_74# a_1314_424# VPB sky130_fd_pr__pfet_01v8 w=840000u l=180000u
X37 VGND D a_422_125# VNB sky130_fd_pr__nfet_01v8_lvt w=420000u l=150000u
X38 a_1708_74# a_1314_424# a_1474_446# VNB sky130_fd_pr__nfet_01v8_lvt w=740000u l=150000u
X39 VPWR a_2320_410# Q VPB sky130_fd_pr__pfet_01v8 w=1.12e+06u l=180000u
.ends

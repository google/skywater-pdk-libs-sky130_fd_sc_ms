# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_ms__ebufn_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.350000 3.865000 1.780000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.582000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.965000 1.180000 3.295000 1.650000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.599200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.615000 0.875000 1.130000 ;
        RECT 0.535000 1.130000 0.705000 1.800000 ;
        RECT 0.535000 1.800000 1.795000 1.970000 ;
        RECT 0.645000 1.970000 1.795000 2.150000 ;
        RECT 0.645000 2.150000 0.975000 2.735000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.250000 0.250000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.080000 0.250000 3.330000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.115000  0.255000 1.375000 0.425000 ;
      RECT 0.115000  0.425000 0.365000 1.130000 ;
      RECT 0.145000  2.140000 0.475000 2.905000 ;
      RECT 0.145000  2.905000 1.475000 3.075000 ;
      RECT 0.875000  1.300000 2.135000 1.630000 ;
      RECT 1.045000  0.425000 1.375000 0.960000 ;
      RECT 1.045000  0.960000 2.225000 1.130000 ;
      RECT 1.145000  2.320000 1.475000 2.580000 ;
      RECT 1.145000  2.580000 2.545000 2.750000 ;
      RECT 1.145000  2.750000 1.475000 2.905000 ;
      RECT 1.545000  0.085000 1.795000 0.790000 ;
      RECT 1.680000  2.920000 2.010000 3.245000 ;
      RECT 1.965000  1.630000 2.135000 2.240000 ;
      RECT 1.965000  2.240000 4.205000 2.410000 ;
      RECT 1.975000  0.350000 2.225000 0.960000 ;
      RECT 2.215000  2.750000 2.545000 2.980000 ;
      RECT 2.395000  0.325000 3.170000 1.010000 ;
      RECT 2.395000  1.010000 2.725000 1.820000 ;
      RECT 2.395000  1.820000 3.105000 2.070000 ;
      RECT 3.225000  2.610000 3.705000 3.245000 ;
      RECT 3.340000  0.085000 3.670000 1.010000 ;
      RECT 3.840000  0.350000 4.205000 1.030000 ;
      RECT 3.875000  1.950000 4.205000 2.240000 ;
      RECT 3.875000  2.410000 4.205000 2.860000 ;
      RECT 4.035000  1.030000 4.205000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_ms__ebufn_2
END LIBRARY

* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_ms__maj3_4 A B C VGND VNB VPB VPWR X
M1000 a_222_392# B a_504_125# VNB nlowvt w=640000u l=150000u
+  ad=5.376e+11p pd=5.52e+06u as=5.41775e+11p ps=4.6e+06u
M1001 X a_222_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=4.44e+11p pd=4.16e+06u as=1.2479e+12p ps=1.196e+07u
M1002 a_908_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=1.971e+12p ps=1.647e+07u
M1003 a_222_392# C a_906_78# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=4.45475e+11p ps=4.25e+06u
M1004 a_222_392# B a_122_392# VPB pshort w=1e+06u l=180000u
+  ad=8.6e+11p pd=7.72e+06u as=5.9e+11p ps=5.18e+06u
M1005 a_222_392# C a_908_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_906_78# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_122_392# A VPWR VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_122_392# B a_222_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A a_122_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND C a_504_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_906_78# C a_222_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A a_906_78# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_908_392# C a_222_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A a_908_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A a_114_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=5.7375e+11p ps=4.61e+06u
M1016 X a_222_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=6.048e+11p pd=5.56e+06u as=0p ps=0u
M1017 a_114_125# B a_222_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_504_125# C VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_222_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_222_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_114_125# A VGND VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 X a_222_392# VPWR VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND a_222_392# X VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_222_392# X VPB pshort w=1.12e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_222_392# B a_114_125# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_504_125# B a_222_392# VNB nlowvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 X a_222_392# VGND VNB nlowvt w=740000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_504_392# C VPWR VPB pshort w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=0p ps=0u
M1029 VPWR C a_504_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_504_392# B a_222_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_222_392# B a_504_392# VPB pshort w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_ms__and2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_ms__and2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.300000 0.435000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.291000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.300000 1.085000 1.780000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.509600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 0.350000 1.795000 0.790000 ;
        RECT 1.595000 1.720000 2.010000 1.890000 ;
        RECT 1.595000 1.890000 1.845000 2.980000 ;
        RECT 1.625000 0.790000 1.795000 0.850000 ;
        RECT 1.625000 0.850000 2.010000 1.020000 ;
        RECT 1.840000 1.020000 2.010000 1.720000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.400000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.245000 2.400000 3.415000 ;
      RECT 0.110000  1.950000 0.440000 3.245000 ;
      RECT 0.135000  0.350000 0.465000 0.960000 ;
      RECT 0.135000  0.960000 1.425000 1.130000 ;
      RECT 0.640000  1.950000 1.425000 2.120000 ;
      RECT 0.640000  2.120000 0.890000 2.980000 ;
      RECT 0.955000  0.085000 1.285000 0.790000 ;
      RECT 1.060000  2.290000 1.390000 3.245000 ;
      RECT 1.255000  1.130000 1.425000 1.220000 ;
      RECT 1.255000  1.220000 1.670000 1.550000 ;
      RECT 1.255000  1.550000 1.425000 1.950000 ;
      RECT 1.975000  0.085000 2.285000 0.680000 ;
      RECT 2.045000  2.060000 2.295000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
  END
END sky130_fd_sc_ms__and2_2
END LIBRARY

* File: sky130_fd_sc_ms__einvn_4.pex.spice
* Created: Fri Aug 28 17:33:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_MS__EINVN_4%TE_B 3 5 7 8 10 12 13 15 17 18 20 22 23 25
+ 27 28 29 30 31 35 39
c95 35 0 5.82364e-21 $X=0.29 $Y=1.465
c96 20 0 8.94367e-20 $X=2.475 $Y=1.725
c97 18 0 1.718e-19 $X=2.385 $Y=1.65
c98 8 0 1.6893e-19 $X=1.485 $Y=1.65
r99 38 39 36.463 $w=4.25e-07 $l=9e-08 $layer=POLY_cond $X=0.565 $Y=1.512
+ $X2=0.655 $Y2=1.512
r100 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.465 $X2=0.29 $Y2=1.465
r101 31 35 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.29 $Y=1.665 $X2=0.29
+ $Y2=1.465
r102 25 27 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=2.975 $Y=1.725
+ $X2=2.975 $Y2=2.4
r103 24 30 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.565 $Y=1.65
+ $X2=2.475 $Y2=1.65
r104 23 25 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.885 $Y=1.65
+ $X2=2.975 $Y2=1.725
r105 23 24 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.885 $Y=1.65
+ $X2=2.565 $Y2=1.65
r106 20 30 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.475 $Y=1.725
+ $X2=2.475 $Y2=1.65
r107 20 22 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=2.475 $Y=1.725
+ $X2=2.475 $Y2=2.4
r108 19 29 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.115 $Y=1.65
+ $X2=2.025 $Y2=1.65
r109 18 30 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.385 $Y=1.65
+ $X2=2.475 $Y2=1.65
r110 18 19 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.385 $Y=1.65
+ $X2=2.115 $Y2=1.65
r111 15 29 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.025 $Y=1.725
+ $X2=2.025 $Y2=1.65
r112 15 17 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=2.025 $Y=1.725
+ $X2=2.025 $Y2=2.4
r113 14 28 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.665 $Y=1.65
+ $X2=1.575 $Y2=1.65
r114 13 29 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.935 $Y=1.65
+ $X2=2.025 $Y2=1.65
r115 13 14 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.935 $Y=1.65
+ $X2=1.665 $Y2=1.65
r116 10 28 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=1.575 $Y=1.725
+ $X2=1.575 $Y2=1.65
r117 10 12 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=1.575 $Y=1.725
+ $X2=1.575 $Y2=2.4
r118 8 28 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.485 $Y=1.65
+ $X2=1.575 $Y2=1.65
r119 8 39 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=1.485 $Y=1.65
+ $X2=0.655 $Y2=1.65
r120 5 38 22.9127 $w=1.8e-07 $l=2.13e-07 $layer=POLY_cond $X=0.565 $Y=1.725
+ $X2=0.565 $Y2=1.512
r121 5 7 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=0.565 $Y=1.725
+ $X2=0.565 $Y2=2.4
r122 1 38 9.16018 $w=4.25e-07 $l=7e-08 $layer=POLY_cond $X=0.495 $Y=1.512
+ $X2=0.565 $Y2=1.512
r123 1 34 26.8262 $w=4.25e-07 $l=2.05e-07 $layer=POLY_cond $X=0.495 $Y=1.512
+ $X2=0.29 $Y2=1.512
r124 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.495 $Y=1.3
+ $X2=0.495 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_MS__EINVN_4%A_114_74# 1 2 7 8 9 11 12 14 16 17 19 21 22
+ 24 26 28 29 30 31 33 39
c89 39 0 3.83609e-19 $X=1.13 $Y=0.465
c90 22 0 1.82848e-19 $X=2.98 $Y=1.26
c91 8 0 5.82364e-21 $X=1.295 $Y=1.26
r92 43 44 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.145 $X2=1.13 $Y2=1.145
r93 41 43 10.4571 $w=7.35e-07 $l=6.3e-07 $layer=LI1_cond $X=0.92 $Y=0.515
+ $X2=0.92 $Y2=1.145
r94 39 44 118.906 $w=3.3e-07 $l=6.8e-07 $layer=POLY_cond $X=1.13 $Y=0.465
+ $X2=1.13 $Y2=1.145
r95 38 41 0.829932 $w=7.35e-07 $l=5e-08 $layer=LI1_cond $X=0.92 $Y=0.465
+ $X2=0.92 $Y2=0.515
r96 38 39 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=0.465 $X2=1.13 $Y2=0.465
r97 33 35 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.79 $Y=1.985
+ $X2=0.79 $Y2=2.815
r98 31 43 6.49103 $w=7.35e-07 $l=2.20624e-07 $layer=LI1_cond $X=0.79 $Y=1.31
+ $X2=0.92 $Y2=1.145
r99 31 33 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.79 $Y=1.31
+ $X2=0.79 $Y2=1.985
r100 27 44 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=1.13 $Y=1.185
+ $X2=1.13 $Y2=1.145
r101 24 26 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=3.055 $Y=1.185
+ $X2=3.055 $Y2=0.74
r102 23 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.26
+ $X2=2.625 $Y2=1.26
r103 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.98 $Y=1.26
+ $X2=3.055 $Y2=1.185
r104 22 23 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=1.26
+ $X2=2.7 $Y2=1.26
r105 19 30 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.625 $Y=1.185
+ $X2=2.625 $Y2=1.26
r106 19 21 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.625 $Y=1.185
+ $X2=2.625 $Y2=0.74
r107 18 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.27 $Y=1.26
+ $X2=2.195 $Y2=1.26
r108 17 30 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=1.26
+ $X2=2.625 $Y2=1.26
r109 17 18 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.26
+ $X2=2.27 $Y2=1.26
r110 14 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.195 $Y=1.185
+ $X2=2.195 $Y2=1.26
r111 14 16 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=2.195 $Y=1.185
+ $X2=2.195 $Y2=0.74
r112 13 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.84 $Y=1.26
+ $X2=1.765 $Y2=1.26
r113 12 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.12 $Y=1.26
+ $X2=2.195 $Y2=1.26
r114 12 13 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.12 $Y=1.26
+ $X2=1.84 $Y2=1.26
r115 9 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=1.185
+ $X2=1.765 $Y2=1.26
r116 9 11 142.993 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=1.765 $Y=1.185
+ $X2=1.765 $Y2=0.74
r117 8 27 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.295 $Y=1.26
+ $X2=1.13 $Y2=1.185
r118 7 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=1.26
+ $X2=1.765 $Y2=1.26
r119 7 8 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.69 $Y=1.26
+ $X2=1.295 $Y2=1.26
r120 2 35 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=0.655
+ $Y=1.84 $X2=0.79 $Y2=2.815
r121 2 33 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.655
+ $Y=1.84 $X2=0.79 $Y2=1.985
r122 1 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.37 $X2=0.71 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__EINVN_4%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 26 39
c84 1 0 6.80292e-20 $X=3.425 $Y=1.725
r85 41 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.88
+ $Y=1.385 $X2=4.88 $Y2=1.385
r86 39 41 9.36401 $w=4.89e-07 $l=9.5e-08 $layer=POLY_cond $X=4.785 $Y=1.472
+ $X2=4.88 $Y2=1.472
r87 38 39 0.985685 $w=4.89e-07 $l=1e-08 $layer=POLY_cond $X=4.775 $Y=1.472
+ $X2=4.785 $Y2=1.472
r88 37 38 41.3988 $w=4.89e-07 $l=4.2e-07 $layer=POLY_cond $X=4.355 $Y=1.472
+ $X2=4.775 $Y2=1.472
r89 36 37 2.95706 $w=4.89e-07 $l=3e-08 $layer=POLY_cond $X=4.325 $Y=1.472
+ $X2=4.355 $Y2=1.472
r90 34 36 12.3211 $w=4.89e-07 $l=1.25e-07 $layer=POLY_cond $X=4.2 $Y=1.472
+ $X2=4.325 $Y2=1.472
r91 34 35 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.2
+ $Y=1.385 $X2=4.2 $Y2=1.385
r92 32 34 28.092 $w=4.89e-07 $l=2.85e-07 $layer=POLY_cond $X=3.915 $Y=1.472
+ $X2=4.2 $Y2=1.472
r93 31 32 3.94274 $w=4.89e-07 $l=4e-08 $layer=POLY_cond $X=3.875 $Y=1.472
+ $X2=3.915 $Y2=1.472
r94 30 31 38.4417 $w=4.89e-07 $l=3.9e-07 $layer=POLY_cond $X=3.485 $Y=1.472
+ $X2=3.875 $Y2=1.472
r95 29 30 5.91411 $w=4.89e-07 $l=6e-08 $layer=POLY_cond $X=3.425 $Y=1.472
+ $X2=3.485 $Y2=1.472
r96 26 42 4.98354 $w=3.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.04 $Y=1.365
+ $X2=4.88 $Y2=1.365
r97 25 42 9.96707 $w=3.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.56 $Y=1.365
+ $X2=4.88 $Y2=1.365
r98 25 35 11.213 $w=3.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.56 $Y=1.365 $X2=4.2
+ $Y2=1.365
r99 22 39 30.8469 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=4.785 $Y=1.22
+ $X2=4.785 $Y2=1.472
r100 22 24 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.785 $Y=1.22
+ $X2=4.785 $Y2=0.74
r101 19 38 26.3167 $w=1.8e-07 $l=2.53e-07 $layer=POLY_cond $X=4.775 $Y=1.725
+ $X2=4.775 $Y2=1.472
r102 19 21 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=4.775 $Y=1.725
+ $X2=4.775 $Y2=2.4
r103 16 37 30.8469 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=4.355 $Y=1.22
+ $X2=4.355 $Y2=1.472
r104 16 18 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.355 $Y=1.22
+ $X2=4.355 $Y2=0.74
r105 13 36 26.3167 $w=1.8e-07 $l=2.53e-07 $layer=POLY_cond $X=4.325 $Y=1.725
+ $X2=4.325 $Y2=1.472
r106 13 15 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=4.325 $Y=1.725
+ $X2=4.325 $Y2=2.4
r107 10 32 30.8469 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=3.915 $Y=1.22
+ $X2=3.915 $Y2=1.472
r108 10 12 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.915 $Y=1.22
+ $X2=3.915 $Y2=0.74
r109 7 31 26.3167 $w=1.8e-07 $l=2.53e-07 $layer=POLY_cond $X=3.875 $Y=1.725
+ $X2=3.875 $Y2=1.472
r110 7 9 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.875 $Y=1.725
+ $X2=3.875 $Y2=2.4
r111 4 30 30.8469 $w=1.5e-07 $l=2.52e-07 $layer=POLY_cond $X=3.485 $Y=1.22
+ $X2=3.485 $Y2=1.472
r112 4 6 154.24 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.485 $Y=1.22
+ $X2=3.485 $Y2=0.74
r113 1 29 26.3167 $w=1.8e-07 $l=2.53e-07 $layer=POLY_cond $X=3.425 $Y=1.725
+ $X2=3.425 $Y2=1.472
r114 1 3 180.75 $w=1.8e-07 $l=6.75e-07 $layer=POLY_cond $X=3.425 $Y=1.725
+ $X2=3.425 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_MS__EINVN_4%VPWR 1 2 3 10 12 18 24 28 30 35 45 46 52 55
r61 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r63 45 46 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r64 43 46 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=5.04 $Y2=3.33
r65 42 45 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=5.04 $Y2=3.33
r66 42 43 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r67 40 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.865 $Y=3.33
+ $X2=2.7 $Y2=3.33
r68 40 42 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.865 $Y=3.33
+ $X2=3.12 $Y2=3.33
r69 39 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r71 36 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.885 $Y=3.33
+ $X2=1.76 $Y2=3.33
r72 36 38 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.885 $Y=3.33
+ $X2=2.16 $Y2=3.33
r73 35 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.535 $Y=3.33
+ $X2=2.7 $Y2=3.33
r74 35 38 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.535 $Y=3.33
+ $X2=2.16 $Y2=3.33
r75 34 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r76 34 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r77 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r78 31 49 3.94169 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r79 31 33 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r80 30 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.635 $Y=3.33
+ $X2=1.76 $Y2=3.33
r81 30 33 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=1.635 $Y=3.33
+ $X2=0.72 $Y2=3.33
r82 28 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r83 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r84 28 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r85 24 27 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=2.7 $Y=1.985 $X2=2.7
+ $Y2=2.815
r86 22 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.7 $Y=3.245 $X2=2.7
+ $Y2=3.33
r87 22 27 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.7 $Y=3.245 $X2=2.7
+ $Y2=2.815
r88 18 21 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=1.76 $Y=1.985
+ $X2=1.76 $Y2=2.815
r89 16 52 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.76 $Y=3.245
+ $X2=1.76 $Y2=3.33
r90 16 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=1.76 $Y=3.245
+ $X2=1.76 $Y2=2.815
r91 12 15 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=0.3 $Y=2.115 $X2=0.3
+ $Y2=2.815
r92 10 49 3.20147 $w=2.5e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.3 $Y=3.245
+ $X2=0.212 $Y2=3.33
r93 10 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.3 $Y=3.245 $X2=0.3
+ $Y2=2.815
r94 3 27 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.565
+ $Y=1.84 $X2=2.7 $Y2=2.815
r95 3 24 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.565
+ $Y=1.84 $X2=2.7 $Y2=1.985
r96 2 21 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=1.665
+ $Y=1.84 $X2=1.8 $Y2=2.815
r97 2 18 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.665
+ $Y=1.84 $X2=1.8 $Y2=1.985
r98 1 15 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.84 $X2=0.34 $Y2=2.815
r99 1 12 400 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.84 $X2=0.34 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_MS__EINVN_4%A_241_368# 1 2 3 4 5 18 22 23 26 30 35 38 39
+ 42 44 48 52 53
c88 39 0 8.94367e-20 $X=3.285 $Y=2.99
c89 35 0 6.80581e-20 $X=3.2 $Y=1.985
r90 48 51 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=5.04 $Y=1.985
+ $X2=5.04 $Y2=2.815
r91 46 51 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=5.04 $Y=2.905 $X2=5.04
+ $Y2=2.815
r92 45 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.185 $Y=2.99 $X2=4.1
+ $Y2=2.99
r93 44 46 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.915 $Y=2.99
+ $X2=5.04 $Y2=2.905
r94 44 45 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.915 $Y=2.99
+ $X2=4.185 $Y2=2.99
r95 40 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.1 $Y=2.905 $X2=4.1
+ $Y2=2.99
r96 40 42 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.1 $Y=2.905 $X2=4.1
+ $Y2=2.225
r97 38 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.015 $Y=2.99 $X2=4.1
+ $Y2=2.99
r98 38 39 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.015 $Y=2.99
+ $X2=3.285 $Y2=2.99
r99 35 37 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=3.16 $Y=1.985
+ $X2=3.16 $Y2=2.815
r100 33 39 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.16 $Y=2.905
+ $X2=3.285 $Y2=2.99
r101 33 37 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=3.16 $Y=2.905
+ $X2=3.16 $Y2=2.815
r102 32 35 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.16 $Y=1.65
+ $X2=3.16 $Y2=1.985
r103 31 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.335 $Y=1.565
+ $X2=2.21 $Y2=1.565
r104 30 32 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.035 $Y=1.565
+ $X2=3.16 $Y2=1.65
r105 30 31 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.035 $Y=1.565
+ $X2=2.335 $Y2=1.565
r106 26 28 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=2.21 $Y=1.985
+ $X2=2.21 $Y2=2.815
r107 24 52 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.21 $Y=1.65
+ $X2=2.21 $Y2=1.565
r108 24 26 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.21 $Y=1.65
+ $X2=2.21 $Y2=1.985
r109 22 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.085 $Y=1.565
+ $X2=2.21 $Y2=1.565
r110 22 23 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.085 $Y=1.565
+ $X2=1.435 $Y2=1.565
r111 18 20 38.2611 $w=2.48e-07 $l=8.3e-07 $layer=LI1_cond $X=1.31 $Y=1.985
+ $X2=1.31 $Y2=2.815
r112 16 23 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.31 $Y=1.65
+ $X2=1.435 $Y2=1.565
r113 16 18 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.31 $Y=1.65
+ $X2=1.31 $Y2=1.985
r114 5 51 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.84 $X2=5 $Y2=2.815
r115 5 48 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.84 $X2=5 $Y2=1.985
r116 4 42 300 $w=1.7e-07 $l=4.47437e-07 $layer=licon1_PDIFF $count=2 $X=3.965
+ $Y=1.84 $X2=4.1 $Y2=2.225
r117 3 37 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=3.065
+ $Y=1.84 $X2=3.2 $Y2=2.815
r118 3 35 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.065
+ $Y=1.84 $X2=3.2 $Y2=1.985
r119 2 28 400 $w=1.7e-07 $l=1.04031e-06 $layer=licon1_PDIFF $count=1 $X=2.115
+ $Y=1.84 $X2=2.25 $Y2=2.815
r120 2 26 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.115
+ $Y=1.84 $X2=2.25 $Y2=1.985
r121 1 20 400 $w=1.7e-07 $l=1.04499e-06 $layer=licon1_PDIFF $count=1 $X=1.205
+ $Y=1.84 $X2=1.35 $Y2=2.815
r122 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.205
+ $Y=1.84 $X2=1.35 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_MS__EINVN_4%Z 1 2 3 4 15 21 23 27 31 37 41 44
c49 44 0 1.82848e-19 $X=3.65 $Y=1.55
c50 21 0 6.80292e-20 $X=4.385 $Y=1.805
r51 41 46 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=3.65 $Y=1.665
+ $X2=3.65 $Y2=1.805
r52 41 44 5.79139 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.65 $Y=1.665
+ $X2=3.65 $Y2=1.55
r53 35 44 23.2909 $w=1.98e-07 $l=4.2e-07 $layer=LI1_cond $X=3.715 $Y=1.13
+ $X2=3.715 $Y2=1.55
r54 34 35 8.79174 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=3.74 $Y=0.95
+ $X2=3.74 $Y2=1.13
r55 31 34 2.76586 $w=2.48e-07 $l=6e-08 $layer=LI1_cond $X=3.74 $Y=0.89 $X2=3.74
+ $Y2=0.95
r56 27 29 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.55 $Y=1.97
+ $X2=4.55 $Y2=2.65
r57 25 27 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.55 $Y=1.89 $X2=4.55
+ $Y2=1.97
r58 24 31 0.964185 $w=2.4e-07 $l=1.25e-07 $layer=LI1_cond $X=3.865 $Y=0.89
+ $X2=3.74 $Y2=0.89
r59 23 37 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.57 $Y=0.89 $X2=4.57
+ $Y2=0.8
r60 23 24 29.7714 $w=2.38e-07 $l=6.2e-07 $layer=LI1_cond $X=4.485 $Y=0.89
+ $X2=3.865 $Y2=0.89
r61 22 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.815 $Y=1.805
+ $X2=3.65 $Y2=1.805
r62 21 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.385 $Y=1.805
+ $X2=4.55 $Y2=1.89
r63 21 22 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.385 $Y=1.805
+ $X2=3.815 $Y2=1.805
r64 15 17 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.65 $Y=1.97
+ $X2=3.65 $Y2=2.65
r65 13 46 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=3.65 $Y=1.89
+ $X2=3.65 $Y2=1.805
r66 13 15 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.65 $Y=1.89 $X2=3.65
+ $Y2=1.97
r67 4 29 400 $w=1.7e-07 $l=8.749e-07 $layer=licon1_PDIFF $count=1 $X=4.415
+ $Y=1.84 $X2=4.55 $Y2=2.65
r68 4 27 400 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_PDIFF $count=1 $X=4.415
+ $Y=1.84 $X2=4.55 $Y2=1.97
r69 3 17 400 $w=1.7e-07 $l=8.749e-07 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=1.84 $X2=3.65 $Y2=2.65
r70 3 15 400 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=1.84 $X2=3.65 $Y2=1.97
r71 2 37 182 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_NDIFF $count=1 $X=4.43
+ $Y=0.37 $X2=4.57 $Y2=0.8
r72 1 34 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.37 $X2=3.7 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_MS__EINVN_4%VGND 1 2 3 10 12 16 20 23 24 26 27 28 44 45
c61 16 0 1.89802e-19 $X=1.98 $Y=0.515
r62 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r63 44 45 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r64 42 45 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=5.04
+ $Y2=0
r65 41 44 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.12 $Y=0 $X2=5.04
+ $Y2=0
r66 41 42 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r67 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r68 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r69 33 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r70 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r71 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r72 30 48 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r73 30 32 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.72
+ $Y2=0
r74 28 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r75 28 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r76 28 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r77 26 38 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.64
+ $Y2=0
r78 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.675 $Y=0 $X2=2.84
+ $Y2=0
r79 25 41 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.005 $Y=0 $X2=3.12
+ $Y2=0
r80 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.005 $Y=0 $X2=2.84
+ $Y2=0
r81 23 35 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=1.68
+ $Y2=0
r82 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=1.98
+ $Y2=0
r83 22 38 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.145 $Y=0 $X2=2.64
+ $Y2=0
r84 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=0 $X2=1.98
+ $Y2=0
r85 18 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=0.085
+ $X2=2.84 $Y2=0
r86 18 20 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.84 $Y=0.085
+ $X2=2.84 $Y2=0.515
r87 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0
r88 14 16 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0.515
r89 10 48 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r90 10 12 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.515
r91 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.7
+ $Y=0.37 $X2=2.84 $Y2=0.515
r92 2 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.37 $X2=1.98 $Y2=0.515
r93 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.37 $X2=0.28 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_MS__EINVN_4%A_281_74# 1 2 3 4 5 18 20 21 24 26 28 29 30
+ 32 36 38 43
c82 38 0 1.718e-19 $X=2.41 $Y=1.225
c83 21 0 3.62737e-19 $X=1.635 $Y=1.225
r84 42 43 8.64642 $w=3.43e-07 $l=1.7e-07 $layer=LI1_cond $X=4.135 $Y=0.427
+ $X2=4.305 $Y2=0.427
r85 34 36 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5 $Y=0.425 $X2=5
+ $Y2=0.68
r86 32 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.835 $Y=0.34
+ $X2=5 $Y2=0.425
r87 32 43 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.835 $Y=0.34
+ $X2=4.305 $Y2=0.34
r88 31 40 2.9551 $w=3.45e-07 $l=1.25e-07 $layer=LI1_cond $X=3.435 $Y=0.427
+ $X2=3.31 $Y2=0.427
r89 30 42 0.0668083 $w=3.43e-07 $l=2e-09 $layer=LI1_cond $X=4.133 $Y=0.427
+ $X2=4.135 $Y2=0.427
r90 30 31 23.3161 $w=3.43e-07 $l=6.98e-07 $layer=LI1_cond $X=4.133 $Y=0.427
+ $X2=3.435 $Y2=0.427
r91 28 40 4.08986 $w=2.5e-07 $l=1.73e-07 $layer=LI1_cond $X=3.31 $Y=0.6 $X2=3.31
+ $Y2=0.427
r92 28 29 24.8928 $w=2.48e-07 $l=5.4e-07 $layer=LI1_cond $X=3.31 $Y=0.6 $X2=3.31
+ $Y2=1.14
r93 27 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.495 $Y=1.225
+ $X2=2.41 $Y2=1.225
r94 26 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.185 $Y=1.225
+ $X2=3.31 $Y2=1.14
r95 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.185 $Y=1.225
+ $X2=2.495 $Y2=1.225
r96 22 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=1.14 $X2=2.41
+ $Y2=1.225
r97 22 24 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.41 $Y=1.14
+ $X2=2.41 $Y2=0.515
r98 20 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.325 $Y=1.225
+ $X2=2.41 $Y2=1.225
r99 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.325 $Y=1.225
+ $X2=1.635 $Y2=1.225
r100 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.55 $Y=1.14
+ $X2=1.635 $Y2=1.225
r101 16 18 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.55 $Y=1.14
+ $X2=1.55 $Y2=0.515
r102 5 36 182 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_NDIFF $count=1 $X=4.86
+ $Y=0.37 $X2=5 $Y2=0.68
r103 4 42 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=3.99
+ $Y=0.37 $X2=4.135 $Y2=0.515
r104 3 40 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.13
+ $Y=0.37 $X2=3.27 $Y2=0.515
r105 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.37 $X2=2.41 $Y2=0.515
r106 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=1.405
+ $Y=0.37 $X2=1.55 $Y2=0.515
.ends

